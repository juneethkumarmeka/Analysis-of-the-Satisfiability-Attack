module basic_2500_25000_3000_8_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
and U0 (N_0,In_1603,In_370);
nor U1 (N_1,In_79,In_148);
nor U2 (N_2,In_896,In_544);
nor U3 (N_3,In_2258,In_2010);
nor U4 (N_4,In_1648,In_658);
nor U5 (N_5,In_1720,In_1500);
or U6 (N_6,In_1310,In_2484);
or U7 (N_7,In_1822,In_596);
xor U8 (N_8,In_1429,In_758);
and U9 (N_9,In_1768,In_1142);
and U10 (N_10,In_411,In_1981);
xnor U11 (N_11,In_2206,In_1431);
and U12 (N_12,In_1449,In_1138);
nand U13 (N_13,In_181,In_109);
nor U14 (N_14,In_2107,In_2271);
nor U15 (N_15,In_290,In_1908);
nor U16 (N_16,In_2468,In_1412);
xnor U17 (N_17,In_425,In_921);
nor U18 (N_18,In_473,In_1040);
nand U19 (N_19,In_1212,In_552);
and U20 (N_20,In_252,In_1240);
and U21 (N_21,In_764,In_219);
and U22 (N_22,In_2009,In_603);
and U23 (N_23,In_1417,In_832);
and U24 (N_24,In_1664,In_1752);
and U25 (N_25,In_114,In_840);
and U26 (N_26,In_1378,In_2116);
and U27 (N_27,In_1807,In_17);
and U28 (N_28,In_51,In_1242);
nor U29 (N_29,In_2238,In_2245);
or U30 (N_30,In_928,In_1344);
or U31 (N_31,In_2433,In_1070);
xnor U32 (N_32,In_1280,In_2353);
xor U33 (N_33,In_1734,In_377);
nor U34 (N_34,In_2007,In_1705);
or U35 (N_35,In_813,In_1639);
or U36 (N_36,In_1728,In_1395);
xor U37 (N_37,In_2482,In_1700);
and U38 (N_38,In_703,In_1208);
or U39 (N_39,In_2331,In_1420);
or U40 (N_40,In_1049,In_2413);
nor U41 (N_41,In_513,In_1007);
xor U42 (N_42,In_1003,In_1444);
nor U43 (N_43,In_1926,In_1618);
or U44 (N_44,In_2290,In_26);
nand U45 (N_45,In_830,In_716);
nand U46 (N_46,In_646,In_1349);
or U47 (N_47,In_1876,In_476);
or U48 (N_48,In_2099,In_1786);
nor U49 (N_49,In_890,In_1690);
and U50 (N_50,In_808,In_1505);
and U51 (N_51,In_167,In_2070);
or U52 (N_52,In_150,In_1064);
nor U53 (N_53,In_730,In_2430);
nor U54 (N_54,In_2462,In_2360);
nand U55 (N_55,In_2022,In_739);
or U56 (N_56,In_2244,In_756);
nand U57 (N_57,In_2459,In_136);
nand U58 (N_58,In_795,In_184);
xor U59 (N_59,In_523,In_296);
nor U60 (N_60,In_774,In_1462);
or U61 (N_61,In_452,In_2154);
nor U62 (N_62,In_271,In_2015);
nor U63 (N_63,In_2033,In_1388);
nor U64 (N_64,In_189,In_120);
nand U65 (N_65,In_1054,In_59);
nor U66 (N_66,In_1520,In_818);
nor U67 (N_67,In_2040,In_330);
and U68 (N_68,In_36,In_591);
nand U69 (N_69,In_230,In_2456);
nor U70 (N_70,In_933,In_21);
or U71 (N_71,In_18,In_1451);
or U72 (N_72,In_2112,In_785);
and U73 (N_73,In_888,In_2076);
nand U74 (N_74,In_563,In_45);
or U75 (N_75,In_710,In_1585);
or U76 (N_76,In_131,In_2182);
nor U77 (N_77,In_2374,In_1535);
or U78 (N_78,In_2348,In_626);
and U79 (N_79,In_328,In_958);
and U80 (N_80,In_2012,In_908);
xnor U81 (N_81,In_10,In_1352);
and U82 (N_82,In_153,In_1622);
or U83 (N_83,In_2043,In_2375);
nand U84 (N_84,In_2253,In_1816);
and U85 (N_85,In_485,In_164);
nand U86 (N_86,In_1011,In_175);
and U87 (N_87,In_227,In_1943);
and U88 (N_88,In_1989,In_418);
or U89 (N_89,In_2432,In_848);
and U90 (N_90,In_2094,In_266);
or U91 (N_91,In_2285,In_292);
nor U92 (N_92,In_2113,In_2442);
nor U93 (N_93,In_1925,In_2179);
and U94 (N_94,In_1909,In_2172);
nor U95 (N_95,In_1015,In_594);
and U96 (N_96,In_842,In_346);
or U97 (N_97,In_1404,In_1631);
and U98 (N_98,In_1961,In_2300);
or U99 (N_99,In_1386,In_963);
xor U100 (N_100,In_1406,In_1375);
or U101 (N_101,In_2342,In_535);
nor U102 (N_102,In_2226,In_500);
nor U103 (N_103,In_668,In_1591);
xnor U104 (N_104,In_1473,In_489);
nand U105 (N_105,In_58,In_639);
or U106 (N_106,In_877,In_2326);
and U107 (N_107,In_1584,In_321);
nand U108 (N_108,In_2307,In_1607);
or U109 (N_109,In_1521,In_715);
or U110 (N_110,In_1491,In_1014);
nand U111 (N_111,In_2277,In_2030);
nor U112 (N_112,In_636,In_422);
nand U113 (N_113,In_2026,In_1595);
nand U114 (N_114,In_1017,In_228);
nand U115 (N_115,In_2254,In_368);
xnor U116 (N_116,In_2117,In_341);
xor U117 (N_117,In_2448,In_1095);
nor U118 (N_118,In_1192,In_255);
xor U119 (N_119,In_681,In_1269);
or U120 (N_120,In_1725,In_1820);
or U121 (N_121,In_1793,In_235);
nor U122 (N_122,In_874,In_986);
and U123 (N_123,In_1244,In_1454);
and U124 (N_124,In_391,In_431);
or U125 (N_125,In_2287,In_1137);
nor U126 (N_126,In_530,In_2496);
nand U127 (N_127,In_53,In_2002);
xor U128 (N_128,In_1944,In_1243);
nor U129 (N_129,In_601,In_588);
and U130 (N_130,In_1812,In_1229);
or U131 (N_131,In_2155,In_168);
nor U132 (N_132,In_216,In_610);
xor U133 (N_133,In_950,In_1608);
or U134 (N_134,In_258,In_420);
nor U135 (N_135,In_772,In_1806);
nor U136 (N_136,In_1892,In_1744);
or U137 (N_137,In_1128,In_1995);
or U138 (N_138,In_738,In_638);
nand U139 (N_139,In_470,In_1588);
or U140 (N_140,In_2205,In_651);
and U141 (N_141,In_1048,In_30);
or U142 (N_142,In_1231,In_2);
and U143 (N_143,In_269,In_1047);
or U144 (N_144,In_1467,In_1679);
nand U145 (N_145,In_14,In_1319);
nor U146 (N_146,In_1029,In_2057);
and U147 (N_147,In_2443,In_2365);
and U148 (N_148,In_213,In_2261);
nor U149 (N_149,In_163,In_1790);
or U150 (N_150,In_2466,In_2233);
nand U151 (N_151,In_1547,In_1108);
nand U152 (N_152,In_358,In_946);
nand U153 (N_153,In_165,In_1996);
nand U154 (N_154,In_1264,In_1785);
and U155 (N_155,In_2477,In_1920);
nor U156 (N_156,In_1435,In_403);
nand U157 (N_157,In_2288,In_696);
nor U158 (N_158,In_43,In_985);
or U159 (N_159,In_860,In_735);
nor U160 (N_160,In_1067,In_171);
xor U161 (N_161,In_1899,In_1504);
or U162 (N_162,In_2311,In_966);
nand U163 (N_163,In_1125,In_1284);
nand U164 (N_164,In_1411,In_108);
and U165 (N_165,In_1617,In_333);
nand U166 (N_166,In_2207,In_1824);
nand U167 (N_167,In_1551,In_2252);
and U168 (N_168,In_1958,In_1202);
nand U169 (N_169,In_424,In_1030);
nand U170 (N_170,In_1236,In_1879);
or U171 (N_171,In_398,In_1298);
xor U172 (N_172,In_699,In_1488);
nor U173 (N_173,In_144,In_1219);
and U174 (N_174,In_1249,In_743);
or U175 (N_175,In_32,In_2495);
nor U176 (N_176,In_798,In_1536);
or U177 (N_177,In_1990,In_866);
and U178 (N_178,In_1457,In_520);
xnor U179 (N_179,In_1151,In_273);
nor U180 (N_180,In_1247,In_1537);
or U181 (N_181,In_1302,In_1530);
nor U182 (N_182,In_105,In_478);
nand U183 (N_183,In_99,In_1282);
nor U184 (N_184,In_2414,In_429);
nand U185 (N_185,In_644,In_1063);
nor U186 (N_186,In_508,In_769);
or U187 (N_187,In_1642,In_701);
xnor U188 (N_188,In_1153,In_2453);
or U189 (N_189,In_1200,In_2037);
or U190 (N_190,In_284,In_2256);
and U191 (N_191,In_1234,In_1238);
and U192 (N_192,In_1522,In_734);
and U193 (N_193,In_2279,In_487);
nand U194 (N_194,In_2020,In_2297);
or U195 (N_195,In_506,In_1938);
nor U196 (N_196,In_2354,In_616);
and U197 (N_197,In_1881,In_1992);
nand U198 (N_198,In_1563,In_1670);
and U199 (N_199,In_1795,In_631);
and U200 (N_200,In_443,In_2302);
nand U201 (N_201,In_1350,In_1903);
or U202 (N_202,In_1448,In_1901);
and U203 (N_203,In_731,In_2493);
or U204 (N_204,In_1727,In_834);
or U205 (N_205,In_1686,In_1321);
xor U206 (N_206,In_940,In_1136);
nor U207 (N_207,In_937,In_930);
or U208 (N_208,In_176,In_1983);
nand U209 (N_209,In_2161,In_750);
and U210 (N_210,In_1327,In_2235);
or U211 (N_211,In_903,In_1428);
nor U212 (N_212,In_1492,In_1283);
nor U213 (N_213,In_2321,In_1737);
or U214 (N_214,In_142,In_548);
and U215 (N_215,In_1760,In_2255);
nand U216 (N_216,In_1366,In_1916);
nor U217 (N_217,In_468,In_598);
or U218 (N_218,In_85,In_286);
xnor U219 (N_219,In_1432,In_1062);
nand U220 (N_220,In_1722,In_15);
nor U221 (N_221,In_1955,In_1154);
and U222 (N_222,In_1121,In_1866);
and U223 (N_223,In_1714,In_1098);
or U224 (N_224,In_1220,In_1484);
nand U225 (N_225,In_2283,In_1132);
nor U226 (N_226,In_1757,In_1114);
nand U227 (N_227,In_34,In_436);
and U228 (N_228,In_2134,In_1788);
nor U229 (N_229,In_1354,In_670);
or U230 (N_230,In_1849,In_2339);
and U231 (N_231,In_1178,In_2494);
nand U232 (N_232,In_2036,In_817);
xnor U233 (N_233,In_690,In_1074);
nand U234 (N_234,In_159,In_9);
or U235 (N_235,In_232,In_215);
or U236 (N_236,In_1754,In_697);
or U237 (N_237,In_349,In_304);
and U238 (N_238,In_637,In_1726);
nand U239 (N_239,In_179,In_1708);
or U240 (N_240,In_760,In_1365);
nand U241 (N_241,In_2332,In_2196);
and U242 (N_242,In_1037,In_684);
nor U243 (N_243,In_556,In_166);
nor U244 (N_244,In_2055,In_1345);
nor U245 (N_245,In_1322,In_177);
nor U246 (N_246,In_665,In_2014);
nand U247 (N_247,In_1106,In_479);
or U248 (N_248,In_231,In_1466);
nor U249 (N_249,In_2091,In_2352);
nor U250 (N_250,In_1965,In_983);
and U251 (N_251,In_540,In_674);
and U252 (N_252,In_2221,In_1079);
or U253 (N_253,In_852,In_2194);
nor U254 (N_254,In_335,In_1886);
nor U255 (N_255,In_1543,In_2241);
nand U256 (N_256,In_2188,In_1833);
nand U257 (N_257,In_1248,In_1994);
nand U258 (N_258,In_206,In_537);
nor U259 (N_259,In_2292,In_1842);
nor U260 (N_260,In_1532,In_766);
nor U261 (N_261,In_624,In_1443);
or U262 (N_262,In_1471,In_2262);
nand U263 (N_263,In_2324,In_1559);
nor U264 (N_264,In_2411,In_570);
nand U265 (N_265,In_2180,In_253);
nor U266 (N_266,In_1515,In_362);
and U267 (N_267,In_2282,In_880);
xnor U268 (N_268,In_1894,In_2230);
nand U269 (N_269,In_498,In_993);
nor U270 (N_270,In_158,In_851);
and U271 (N_271,In_2157,In_653);
and U272 (N_272,In_155,In_1534);
or U273 (N_273,In_2426,In_600);
or U274 (N_274,In_1698,In_1813);
nand U275 (N_275,In_753,In_1847);
and U276 (N_276,In_477,In_902);
and U277 (N_277,In_187,In_895);
or U278 (N_278,In_1256,In_1383);
xor U279 (N_279,In_384,In_115);
and U280 (N_280,In_931,In_495);
and U281 (N_281,In_1568,In_221);
nand U282 (N_282,In_975,In_1278);
nor U283 (N_283,In_2052,In_2425);
nor U284 (N_284,In_1258,In_2059);
xnor U285 (N_285,In_2195,In_2129);
nand U286 (N_286,In_143,In_1921);
and U287 (N_287,In_649,In_240);
and U288 (N_288,In_622,In_742);
and U289 (N_289,In_2387,In_1371);
or U290 (N_290,In_791,In_545);
nand U291 (N_291,In_1133,In_1170);
or U292 (N_292,In_1050,In_979);
xnor U293 (N_293,In_602,In_2485);
nand U294 (N_294,In_2431,In_2200);
nand U295 (N_295,In_320,In_2369);
or U296 (N_296,In_1835,In_1374);
xor U297 (N_297,In_1615,In_97);
nand U298 (N_298,In_133,In_1461);
xor U299 (N_299,In_1544,In_1748);
and U300 (N_300,In_2248,In_581);
xnor U301 (N_301,In_1272,In_1453);
nor U302 (N_302,In_2217,In_381);
or U303 (N_303,In_1102,In_771);
and U304 (N_304,In_2054,In_359);
nand U305 (N_305,In_765,In_347);
nand U306 (N_306,In_73,In_2388);
nand U307 (N_307,In_936,In_2489);
nand U308 (N_308,In_1541,In_1818);
nor U309 (N_309,In_1840,In_107);
nor U310 (N_310,In_233,In_1305);
nor U311 (N_311,In_2424,In_981);
and U312 (N_312,In_451,In_1742);
and U313 (N_313,In_679,In_2338);
or U314 (N_314,In_988,In_2275);
and U315 (N_315,In_723,In_1415);
and U316 (N_316,In_1006,In_1624);
or U317 (N_317,In_820,In_589);
and U318 (N_318,In_428,In_1948);
or U319 (N_319,In_1368,In_961);
nor U320 (N_320,In_1235,In_2164);
nor U321 (N_321,In_640,In_1335);
xnor U322 (N_322,In_1105,In_1086);
xor U323 (N_323,In_1896,In_906);
and U324 (N_324,In_1381,In_2240);
and U325 (N_325,In_74,In_2158);
and U326 (N_326,In_52,In_1499);
and U327 (N_327,In_19,In_2438);
nor U328 (N_328,In_1186,In_1286);
nor U329 (N_329,In_1171,In_1677);
or U330 (N_330,In_499,In_1394);
and U331 (N_331,In_1845,In_1507);
and U332 (N_332,In_305,In_7);
or U333 (N_333,In_827,In_1629);
or U334 (N_334,In_1287,In_247);
nand U335 (N_335,In_655,In_1041);
nand U336 (N_336,In_799,In_410);
and U337 (N_337,In_2165,In_1685);
or U338 (N_338,In_844,In_1158);
and U339 (N_339,In_1226,In_3);
and U340 (N_340,In_1065,In_2077);
and U341 (N_341,In_1330,In_1433);
and U342 (N_342,In_409,In_1023);
nand U343 (N_343,In_1717,In_641);
and U344 (N_344,In_1092,In_1191);
xnor U345 (N_345,In_666,In_1557);
and U346 (N_346,In_2122,In_920);
or U347 (N_347,In_900,In_2492);
and U348 (N_348,In_719,In_1377);
nand U349 (N_349,In_122,In_1055);
or U350 (N_350,In_343,In_1848);
nor U351 (N_351,In_406,In_2420);
nor U352 (N_352,In_2016,In_2347);
or U353 (N_353,In_2084,In_922);
or U354 (N_354,In_2296,In_50);
or U355 (N_355,In_1001,In_31);
and U356 (N_356,In_2111,In_1008);
and U357 (N_357,In_207,In_139);
nor U358 (N_358,In_486,In_426);
xor U359 (N_359,In_1085,In_2368);
nor U360 (N_360,In_2219,In_1638);
xnor U361 (N_361,In_483,In_1960);
nand U362 (N_362,In_2362,In_1463);
or U363 (N_363,In_2384,In_110);
nand U364 (N_364,In_512,In_1843);
nor U365 (N_365,In_1147,In_833);
or U366 (N_366,In_643,In_98);
xor U367 (N_367,In_1834,In_1398);
nor U368 (N_368,In_1456,In_1323);
nor U369 (N_369,In_664,In_84);
nor U370 (N_370,In_809,In_667);
nor U371 (N_371,In_62,In_259);
nor U372 (N_372,In_1068,In_557);
nand U373 (N_373,In_2104,In_127);
nand U374 (N_374,In_741,In_200);
or U375 (N_375,In_1204,In_1237);
xnor U376 (N_376,In_521,In_279);
xor U377 (N_377,In_1127,In_1019);
nor U378 (N_378,In_369,In_1980);
and U379 (N_379,In_1052,In_361);
nand U380 (N_380,In_2460,In_1392);
or U381 (N_381,In_1478,In_916);
nor U382 (N_382,In_1711,In_1773);
and U383 (N_383,In_2276,In_2062);
and U384 (N_384,In_198,In_492);
nor U385 (N_385,In_106,In_1416);
or U386 (N_386,In_2437,In_23);
or U387 (N_387,In_354,In_2467);
nand U388 (N_388,In_1749,In_2399);
nor U389 (N_389,In_1779,In_1567);
nand U390 (N_390,In_314,In_2146);
nand U391 (N_391,In_1299,In_609);
nand U392 (N_392,In_380,In_752);
and U393 (N_393,In_2303,In_1828);
nand U394 (N_394,In_1458,In_2457);
or U395 (N_395,In_1906,In_620);
and U396 (N_396,In_2143,In_2359);
or U397 (N_397,In_2102,In_821);
and U398 (N_398,In_22,In_1288);
or U399 (N_399,In_2449,In_2047);
nor U400 (N_400,In_590,In_660);
nor U401 (N_401,In_1599,In_2137);
nand U402 (N_402,In_1053,In_2476);
nand U403 (N_403,In_1671,In_308);
xnor U404 (N_404,In_415,In_1517);
nor U405 (N_405,In_515,In_1214);
nor U406 (N_406,In_287,In_1610);
and U407 (N_407,In_1391,In_300);
nand U408 (N_408,In_2228,In_718);
or U409 (N_409,In_1945,In_262);
and U410 (N_410,In_1823,In_1109);
or U411 (N_411,In_2395,In_137);
xor U412 (N_412,In_389,In_959);
or U413 (N_413,In_185,In_1946);
or U414 (N_414,In_1546,In_777);
nor U415 (N_415,In_342,In_773);
and U416 (N_416,In_1713,In_1611);
or U417 (N_417,In_299,In_1035);
nand U418 (N_418,In_494,In_2184);
nand U419 (N_419,In_397,In_1026);
nand U420 (N_420,In_663,In_151);
and U421 (N_421,In_83,In_319);
xor U422 (N_422,In_125,In_574);
xor U423 (N_423,In_732,In_1791);
nand U424 (N_424,In_1089,In_2396);
or U425 (N_425,In_2463,In_1940);
and U426 (N_426,In_547,In_1087);
or U427 (N_427,In_1018,In_1163);
nor U428 (N_428,In_1578,In_1738);
nor U429 (N_429,In_654,In_1117);
xnor U430 (N_430,In_2295,In_621);
and U431 (N_431,In_265,In_356);
and U432 (N_432,In_951,In_35);
xor U433 (N_433,In_1043,In_1772);
nand U434 (N_434,In_934,In_2092);
or U435 (N_435,In_650,In_2415);
or U436 (N_436,In_1941,In_623);
nand U437 (N_437,In_1157,In_2478);
and U438 (N_438,In_1852,In_1045);
or U439 (N_439,In_1558,In_1699);
nand U440 (N_440,In_2325,In_307);
nor U441 (N_441,In_438,In_283);
nor U442 (N_442,In_1424,In_2163);
or U443 (N_443,In_2142,In_587);
nor U444 (N_444,In_1873,In_126);
xor U445 (N_445,In_889,In_134);
nand U446 (N_446,In_571,In_1885);
or U447 (N_447,In_2141,In_2162);
nand U448 (N_448,In_1273,In_1739);
nand U449 (N_449,In_2066,In_2440);
nor U450 (N_450,In_1218,In_944);
or U451 (N_451,In_1553,In_671);
or U452 (N_452,In_432,In_463);
nor U453 (N_453,In_952,In_1183);
and U454 (N_454,In_980,In_1216);
nand U455 (N_455,In_1169,In_254);
xnor U456 (N_456,In_1704,In_1796);
or U457 (N_457,In_2061,In_416);
and U458 (N_458,In_1759,In_427);
or U459 (N_459,In_1645,In_1856);
and U460 (N_460,In_1985,In_1180);
xor U461 (N_461,In_2334,In_1403);
or U462 (N_462,In_824,In_178);
or U463 (N_463,In_1152,In_855);
or U464 (N_464,In_1933,In_1712);
nand U465 (N_465,In_712,In_1351);
or U466 (N_466,In_546,In_1575);
and U467 (N_467,In_1252,In_1110);
and U468 (N_468,In_2081,In_568);
nand U469 (N_469,In_2087,In_1215);
or U470 (N_470,In_2089,In_1819);
or U471 (N_471,In_135,In_1889);
nand U472 (N_472,In_1450,In_291);
nor U473 (N_473,In_1359,In_1576);
nand U474 (N_474,In_1592,In_285);
or U475 (N_475,In_1266,In_2082);
or U476 (N_476,In_1687,In_220);
or U477 (N_477,In_2109,In_2298);
xor U478 (N_478,In_659,In_2436);
nand U479 (N_479,In_272,In_2358);
or U480 (N_480,In_1957,In_1494);
or U481 (N_481,In_691,In_2259);
nand U482 (N_482,In_1002,In_2029);
or U483 (N_483,In_1174,In_1560);
nand U484 (N_484,In_1005,In_2427);
nand U485 (N_485,In_871,In_33);
xor U486 (N_486,In_965,In_706);
nand U487 (N_487,In_837,In_1732);
and U488 (N_488,In_1134,In_2377);
and U489 (N_489,In_978,In_1021);
nor U490 (N_490,In_1767,In_1389);
or U491 (N_491,In_1781,In_1486);
nand U492 (N_492,In_194,In_618);
nand U493 (N_493,In_1073,In_1988);
nor U494 (N_494,In_4,In_1666);
and U495 (N_495,In_350,In_1027);
nor U496 (N_496,In_2363,In_439);
or U497 (N_497,In_682,In_1213);
nand U498 (N_498,In_444,In_104);
nor U499 (N_499,In_1910,In_2380);
or U500 (N_500,In_72,In_413);
nand U501 (N_501,In_913,In_1844);
nand U502 (N_502,In_1402,In_2232);
and U503 (N_503,In_1195,In_1482);
or U504 (N_504,In_1259,In_997);
and U505 (N_505,In_904,In_1977);
or U506 (N_506,In_862,In_5);
nand U507 (N_507,In_2120,In_414);
xor U508 (N_508,In_1718,In_1929);
and U509 (N_509,In_1703,In_2312);
nor U510 (N_510,In_1755,In_1271);
and U511 (N_511,In_1827,In_911);
nand U512 (N_512,In_1328,In_214);
nor U513 (N_513,In_1285,In_536);
and U514 (N_514,In_686,In_113);
nor U515 (N_515,In_417,In_1851);
and U516 (N_516,In_1789,In_289);
or U517 (N_517,In_2058,In_1604);
nor U518 (N_518,In_46,In_1116);
or U519 (N_519,In_48,In_1295);
xnor U520 (N_520,In_2450,In_2171);
nand U521 (N_521,In_1953,In_1257);
or U522 (N_522,In_316,In_1605);
nand U523 (N_523,In_267,In_562);
and U524 (N_524,In_1654,In_49);
or U525 (N_525,In_982,In_2049);
nand U526 (N_526,In_223,In_355);
nor U527 (N_527,In_2193,In_1290);
xor U528 (N_528,In_1115,In_870);
and U529 (N_529,In_1656,In_90);
xnor U530 (N_530,In_504,In_2469);
or U531 (N_531,In_387,In_1337);
or U532 (N_532,In_1255,In_1614);
nor U533 (N_533,In_1915,In_2191);
and U534 (N_534,In_2491,In_327);
nand U535 (N_535,In_256,In_229);
nand U536 (N_536,In_1012,In_1877);
nand U537 (N_537,In_632,In_947);
and U538 (N_538,In_2257,In_241);
nor U539 (N_539,In_2045,In_2389);
xnor U540 (N_540,In_344,In_2383);
and U541 (N_541,In_2187,In_1724);
nand U542 (N_542,In_1164,In_124);
or U543 (N_543,In_2319,In_1710);
xor U544 (N_544,In_669,In_1071);
nand U545 (N_545,In_1692,In_974);
or U546 (N_546,In_1882,In_884);
or U547 (N_547,In_2034,In_1855);
and U548 (N_548,In_29,In_1223);
xnor U549 (N_549,In_1009,In_1805);
or U550 (N_550,In_1959,In_925);
nor U551 (N_551,In_2445,In_170);
nand U552 (N_552,In_2314,In_1735);
nand U553 (N_553,In_1609,In_2304);
nand U554 (N_554,In_720,In_779);
or U555 (N_555,In_2159,In_2323);
nor U556 (N_556,In_2222,In_2446);
nand U557 (N_557,In_1036,In_68);
nor U558 (N_558,In_138,In_806);
nor U559 (N_559,In_1556,In_1168);
nor U560 (N_560,In_239,In_2486);
nor U561 (N_561,In_1928,In_807);
or U562 (N_562,In_689,In_2273);
nand U563 (N_563,In_2067,In_2498);
or U564 (N_564,In_1746,In_672);
and U565 (N_565,In_2291,In_37);
nand U566 (N_566,In_2098,In_1911);
and U567 (N_567,In_502,In_1188);
or U568 (N_568,In_1438,In_1141);
and U569 (N_569,In_1838,In_1583);
nand U570 (N_570,In_2215,In_236);
and U571 (N_571,In_1890,In_329);
and U572 (N_572,In_605,In_2176);
xor U573 (N_573,In_858,In_280);
nand U574 (N_574,In_613,In_519);
nor U575 (N_575,In_27,In_1459);
nor U576 (N_576,In_1090,In_1401);
nor U577 (N_577,In_1628,In_1081);
and U578 (N_578,In_787,In_1436);
nand U579 (N_579,In_1148,In_0);
nor U580 (N_580,In_1221,In_915);
and U581 (N_581,In_2050,In_324);
nor U582 (N_582,In_2063,In_614);
or U583 (N_583,In_1172,In_317);
nor U584 (N_584,In_1691,In_2153);
or U585 (N_585,In_1093,In_69);
nor U586 (N_586,In_2447,In_203);
nand U587 (N_587,In_2133,In_615);
or U588 (N_588,In_2350,In_2421);
nand U589 (N_589,In_1028,In_678);
nor U590 (N_590,In_977,In_402);
nand U591 (N_591,In_191,In_2263);
or U592 (N_592,In_804,In_1301);
or U593 (N_593,In_1112,In_687);
nor U594 (N_594,In_94,In_174);
and U595 (N_595,In_16,In_1902);
nand U596 (N_596,In_2379,In_582);
and U597 (N_597,In_1821,In_2214);
or U598 (N_598,In_599,In_2328);
and U599 (N_599,In_1733,In_1753);
nand U600 (N_600,In_747,In_2381);
xor U601 (N_601,In_1801,In_1613);
or U602 (N_602,In_1808,In_6);
and U603 (N_603,In_318,In_24);
xor U604 (N_604,In_2422,In_825);
and U605 (N_605,In_1189,In_1419);
or U606 (N_606,In_1637,In_1487);
and U607 (N_607,In_1770,In_2105);
xor U608 (N_608,In_81,In_2470);
and U609 (N_609,In_676,In_210);
nand U610 (N_610,In_2372,In_340);
or U611 (N_611,In_1069,In_140);
xnor U612 (N_612,In_633,In_1783);
nand U613 (N_613,In_625,In_2183);
xnor U614 (N_614,In_1950,In_1156);
or U615 (N_615,In_2340,In_1279);
or U616 (N_616,In_918,In_1315);
nor U617 (N_617,In_2079,In_2173);
and U618 (N_618,In_2027,In_989);
or U619 (N_619,In_430,In_593);
and U620 (N_620,In_962,In_1696);
nand U621 (N_621,In_2246,In_2013);
and U622 (N_622,In_1442,In_763);
nand U623 (N_623,In_1190,In_1775);
nor U624 (N_624,In_160,In_1472);
and U625 (N_625,In_1425,In_882);
or U626 (N_626,In_169,In_1004);
or U627 (N_627,In_976,In_39);
nor U628 (N_628,In_1262,In_1144);
or U629 (N_629,In_2320,In_2074);
nand U630 (N_630,In_1393,In_183);
or U631 (N_631,In_310,In_1572);
nand U632 (N_632,In_2284,In_1644);
nand U633 (N_633,In_1832,In_1861);
and U634 (N_634,In_1730,In_584);
and U635 (N_635,In_2458,In_1715);
nor U636 (N_636,In_816,In_2028);
and U637 (N_637,In_1640,In_1379);
nand U638 (N_638,In_1160,In_1650);
nand U639 (N_639,In_1776,In_2023);
and U640 (N_640,In_859,In_2119);
nand U641 (N_641,In_802,In_388);
nand U642 (N_642,In_2386,In_2398);
and U643 (N_643,In_1799,In_364);
nor U644 (N_644,In_1673,In_2220);
nand U645 (N_645,In_2391,In_1951);
and U646 (N_646,In_1939,In_955);
and U647 (N_647,In_2202,In_2465);
and U648 (N_648,In_192,In_505);
and U649 (N_649,In_1974,In_395);
nand U650 (N_650,In_1721,In_209);
and U651 (N_651,In_149,In_1293);
or U652 (N_652,In_2224,In_1201);
and U653 (N_653,In_2305,In_237);
or U654 (N_654,In_2208,In_1542);
xor U655 (N_655,In_1874,In_553);
or U656 (N_656,In_2267,In_281);
and U657 (N_657,In_1803,In_1829);
nand U658 (N_658,In_943,In_401);
nor U659 (N_659,In_1421,In_607);
nor U660 (N_660,In_1013,In_80);
and U661 (N_661,In_2315,In_768);
nor U662 (N_662,In_996,In_1103);
and U663 (N_663,In_1331,In_1384);
or U664 (N_664,In_938,In_1225);
nor U665 (N_665,In_1145,In_784);
or U666 (N_666,In_490,In_1184);
nor U667 (N_667,In_1787,In_1993);
xnor U668 (N_668,In_2144,In_1306);
or U669 (N_669,In_386,In_685);
or U670 (N_670,In_1367,In_2021);
or U671 (N_671,In_1346,In_1590);
nand U672 (N_672,In_481,In_472);
xor U673 (N_673,In_1241,In_572);
and U674 (N_674,In_526,In_991);
nor U675 (N_675,In_1265,In_55);
xor U676 (N_676,In_268,In_1495);
nand U677 (N_677,In_251,In_1978);
and U678 (N_678,In_707,In_1122);
and U679 (N_679,In_87,In_385);
nand U680 (N_680,In_1826,In_186);
or U681 (N_681,In_1589,In_465);
nor U682 (N_682,In_1493,In_1632);
or U683 (N_683,In_1771,In_2210);
nand U684 (N_684,In_2345,In_932);
and U685 (N_685,In_2073,In_939);
or U686 (N_686,In_1082,In_1689);
nand U687 (N_687,In_2088,In_1232);
nand U688 (N_688,In_972,In_1777);
or U689 (N_689,In_1039,In_1475);
or U690 (N_690,In_1778,In_1080);
and U691 (N_691,In_2125,In_2402);
or U692 (N_692,In_1870,In_1347);
nand U693 (N_693,In_929,In_1490);
nand U694 (N_694,In_1927,In_948);
nor U695 (N_695,In_453,In_2250);
and U696 (N_696,In_1586,In_1762);
nor U697 (N_697,In_1177,In_1489);
and U698 (N_698,In_234,In_2211);
and U699 (N_699,In_224,In_1659);
nor U700 (N_700,In_790,In_1320);
nor U701 (N_701,In_128,In_2439);
and U702 (N_702,In_754,In_579);
xnor U703 (N_703,In_998,In_274);
nand U704 (N_704,In_1410,In_1905);
or U705 (N_705,In_1066,In_2095);
nand U706 (N_706,In_1869,In_2264);
nor U707 (N_707,In_1665,In_1326);
nor U708 (N_708,In_1853,In_897);
or U709 (N_709,In_796,In_1199);
or U710 (N_710,In_709,In_293);
or U711 (N_711,In_2203,In_257);
nand U712 (N_712,In_1859,In_459);
and U713 (N_713,In_2151,In_1268);
xor U714 (N_714,In_1782,In_1857);
or U715 (N_715,In_528,In_2370);
nor U716 (N_716,In_1313,In_1300);
or U717 (N_717,In_746,In_433);
and U718 (N_718,In_2428,In_375);
nand U719 (N_719,In_482,In_1736);
nand U720 (N_720,In_2167,In_1549);
nand U721 (N_721,In_1907,In_276);
and U722 (N_722,In_1975,In_1501);
nand U723 (N_723,In_1662,In_1124);
or U724 (N_724,In_129,In_910);
nor U725 (N_725,In_1647,In_1119);
xor U726 (N_726,In_767,In_154);
and U727 (N_727,In_2145,In_2064);
xor U728 (N_728,In_1860,In_1780);
xnor U729 (N_729,In_1895,In_2225);
nand U730 (N_730,In_1101,In_93);
or U731 (N_731,In_1477,In_1967);
nor U732 (N_732,In_2382,In_450);
and U733 (N_733,In_1088,In_531);
or U734 (N_734,In_2346,In_2131);
xor U735 (N_735,In_372,In_549);
or U736 (N_736,In_2025,In_1303);
nand U737 (N_737,In_1469,In_66);
nand U738 (N_738,In_1020,In_1952);
nand U739 (N_739,In_529,In_180);
nor U740 (N_740,In_2185,In_1511);
xor U741 (N_741,In_919,In_559);
and U742 (N_742,In_2227,In_1518);
nand U743 (N_743,In_1674,In_1669);
and U744 (N_744,In_111,In_1000);
nand U745 (N_745,In_1130,In_57);
or U746 (N_746,In_1470,In_1336);
nor U747 (N_747,In_1680,In_2132);
nor U748 (N_748,In_1548,In_1376);
or U749 (N_749,In_1937,In_2293);
or U750 (N_750,In_38,In_1176);
or U751 (N_751,In_872,In_1126);
nor U752 (N_752,In_2138,In_2174);
or U753 (N_753,In_1918,In_373);
xor U754 (N_754,In_576,In_509);
nand U755 (N_755,In_1513,In_1312);
nor U756 (N_756,In_2265,In_886);
and U757 (N_757,In_1593,In_2268);
and U758 (N_758,In_776,In_782);
nor U759 (N_759,In_1333,In_1099);
nand U760 (N_760,In_2170,In_803);
and U761 (N_761,In_899,In_2135);
or U762 (N_762,In_2306,In_1564);
nand U763 (N_763,In_1769,In_1516);
xnor U764 (N_764,In_1668,In_288);
nor U765 (N_765,In_1774,In_1797);
xnor U766 (N_766,In_1175,In_2101);
and U767 (N_767,In_2371,In_1574);
and U768 (N_768,In_627,In_2218);
nand U769 (N_769,In_243,In_1051);
or U770 (N_770,In_811,In_1620);
xor U771 (N_771,In_2213,In_1441);
nor U772 (N_772,In_525,In_102);
or U773 (N_773,In_322,In_2078);
or U774 (N_774,In_1527,In_2497);
nor U775 (N_775,In_1973,In_13);
or U776 (N_776,In_2190,In_733);
or U777 (N_777,In_1042,In_907);
or U778 (N_778,In_1625,In_990);
nand U779 (N_779,In_692,In_2429);
xor U780 (N_780,In_1701,In_2317);
or U781 (N_781,In_843,In_786);
nor U782 (N_782,In_2487,In_867);
nand U783 (N_783,In_1373,In_484);
nand U784 (N_784,In_604,In_680);
nor U785 (N_785,In_2110,In_41);
and U786 (N_786,In_1947,In_2086);
nor U787 (N_787,In_2106,In_475);
nor U788 (N_788,In_2483,In_1923);
nor U789 (N_789,In_1539,In_1135);
and U790 (N_790,In_1427,In_173);
and U791 (N_791,In_551,In_1962);
nor U792 (N_792,In_182,In_2404);
xor U793 (N_793,In_70,In_2071);
nand U794 (N_794,In_1526,In_2344);
and U795 (N_795,In_863,In_390);
and U796 (N_796,In_371,In_1930);
nor U797 (N_797,In_226,In_822);
nor U798 (N_798,In_2451,In_2318);
xnor U799 (N_799,In_96,In_1524);
or U800 (N_800,In_1514,In_847);
or U801 (N_801,In_1304,In_2005);
or U802 (N_802,In_583,In_2090);
nand U803 (N_803,In_1399,In_2299);
nor U804 (N_804,In_2140,In_2418);
nand U805 (N_805,In_797,In_1678);
or U806 (N_806,In_1653,In_1763);
or U807 (N_807,In_964,In_1914);
nor U808 (N_808,In_88,In_2280);
or U809 (N_809,In_801,In_1274);
nand U810 (N_810,In_1854,In_2199);
and U811 (N_811,In_748,In_1646);
and U812 (N_812,In_914,In_25);
nor U813 (N_813,In_2357,In_1538);
xor U814 (N_814,In_2364,In_901);
nor U815 (N_815,In_270,In_2351);
xor U816 (N_816,In_464,In_2011);
and U817 (N_817,In_2480,In_2243);
or U818 (N_818,In_841,In_1676);
and U819 (N_819,In_1107,In_1031);
nor U820 (N_820,In_2044,In_458);
or U821 (N_821,In_713,In_1123);
nor U822 (N_822,In_1131,In_1596);
or U823 (N_823,In_543,In_1512);
nor U824 (N_824,In_1033,In_1075);
nand U825 (N_825,In_1887,In_1196);
xnor U826 (N_826,In_1716,In_629);
and U827 (N_827,In_60,In_971);
and U828 (N_828,In_1942,In_561);
and U829 (N_829,In_700,In_1623);
nor U830 (N_830,In_770,In_2126);
nor U831 (N_831,In_331,In_1426);
or U832 (N_832,In_42,In_1032);
nor U833 (N_833,In_2069,In_1228);
and U834 (N_834,In_2096,In_737);
nor U835 (N_835,In_2006,In_1440);
and U836 (N_836,In_1332,In_442);
nand U837 (N_837,In_394,In_396);
nor U838 (N_838,In_1340,In_2473);
nand U839 (N_839,In_1100,In_145);
nor U840 (N_840,In_698,In_1372);
nor U841 (N_841,In_2423,In_2108);
nand U842 (N_842,In_1481,In_1418);
or U843 (N_843,In_1113,In_313);
xor U844 (N_844,In_1598,In_86);
nand U845 (N_845,In_1956,In_404);
nand U846 (N_846,In_1949,In_1969);
xnor U847 (N_847,In_474,In_1363);
nand U848 (N_848,In_1291,In_923);
nor U849 (N_849,In_1913,In_2065);
nand U850 (N_850,In_1275,In_1010);
nor U851 (N_851,In_44,In_728);
and U852 (N_852,In_130,In_54);
or U853 (N_853,In_1872,In_1550);
nand U854 (N_854,In_1723,In_2197);
and U855 (N_855,In_1276,In_2019);
xor U856 (N_856,In_2051,In_1307);
or U857 (N_857,In_1810,In_457);
and U858 (N_858,In_2053,In_1211);
or U859 (N_859,In_573,In_1764);
nand U860 (N_860,In_365,In_606);
and U861 (N_861,In_440,In_560);
and U862 (N_862,In_1206,In_63);
xor U863 (N_863,In_2266,In_2018);
nand U864 (N_864,In_1697,In_1966);
and U865 (N_865,In_408,In_2186);
nand U866 (N_866,In_724,In_2454);
nor U867 (N_867,In_2349,In_2366);
or U868 (N_868,In_673,In_2192);
nand U869 (N_869,In_987,In_1046);
or U870 (N_870,In_1525,In_711);
nor U871 (N_871,In_612,In_1447);
or U872 (N_872,In_2212,In_761);
or U873 (N_873,In_467,In_1839);
nor U874 (N_874,In_466,In_2416);
nand U875 (N_875,In_2083,In_2085);
nand U876 (N_876,In_554,In_1129);
nor U877 (N_877,In_942,In_2335);
or U878 (N_878,In_345,In_1658);
nand U879 (N_879,In_2269,In_1661);
or U880 (N_880,In_2128,In_496);
nor U881 (N_881,In_1750,In_100);
or U882 (N_882,In_1922,In_2475);
or U883 (N_883,In_1254,In_2166);
nand U884 (N_884,In_1334,In_1660);
xnor U885 (N_885,In_839,In_2000);
and U886 (N_886,In_968,In_1924);
nor U887 (N_887,In_337,In_1422);
nor U888 (N_888,In_1991,In_1187);
or U889 (N_889,In_1999,In_1239);
and U890 (N_890,In_2309,In_617);
nor U891 (N_891,In_662,In_275);
or U892 (N_892,In_2322,In_2123);
xnor U893 (N_893,In_1396,In_967);
nand U894 (N_894,In_2376,In_1672);
or U895 (N_895,In_211,In_2455);
and U896 (N_896,In_1875,In_510);
or U897 (N_897,In_2239,In_1528);
nand U898 (N_898,In_1883,In_1465);
xor U899 (N_899,In_261,In_311);
and U900 (N_900,In_103,In_683);
or U901 (N_901,In_2308,In_2032);
nor U902 (N_902,In_1510,In_1864);
xor U903 (N_903,In_249,In_469);
and U904 (N_904,In_278,In_1519);
nor U905 (N_905,In_2367,In_2336);
and U906 (N_906,In_56,In_1675);
or U907 (N_907,In_1800,In_1917);
and U908 (N_908,In_2406,In_2177);
xor U909 (N_909,In_2041,In_755);
nor U910 (N_910,In_2118,In_1695);
xnor U911 (N_911,In_1540,In_1709);
or U912 (N_912,In_694,In_1060);
xnor U913 (N_913,In_1863,In_1837);
nor U914 (N_914,In_778,In_1809);
and U915 (N_915,In_1165,In_1413);
and U916 (N_916,In_1203,In_956);
or U917 (N_917,In_471,In_1056);
and U918 (N_918,In_1059,In_1364);
or U919 (N_919,In_1260,In_172);
nand U920 (N_920,In_1635,In_2046);
nor U921 (N_921,In_1626,In_2394);
nand U922 (N_922,In_883,In_2100);
and U923 (N_923,In_1318,In_1606);
xor U924 (N_924,In_2042,In_1681);
nand U925 (N_925,In_729,In_162);
xor U926 (N_926,In_118,In_957);
nor U927 (N_927,In_2139,In_1719);
or U928 (N_928,In_1729,In_1579);
nor U929 (N_929,In_1731,In_1963);
nor U930 (N_930,In_1954,In_744);
and U931 (N_931,In_1562,In_2168);
and U932 (N_932,In_1224,In_794);
nand U933 (N_933,In_2390,In_2114);
nand U934 (N_934,In_2223,In_2189);
or U935 (N_935,In_1209,In_1360);
and U936 (N_936,In_92,In_294);
nor U937 (N_937,In_238,In_592);
xnor U938 (N_938,In_935,In_1566);
xor U939 (N_939,In_927,In_894);
or U940 (N_940,In_1057,In_1569);
or U941 (N_941,In_1747,In_1246);
nand U942 (N_942,In_857,In_8);
and U943 (N_943,In_960,In_1437);
nand U944 (N_944,In_1250,In_2169);
or U945 (N_945,In_575,In_656);
and U946 (N_946,In_1143,In_121);
and U947 (N_947,In_1968,In_2001);
or U948 (N_948,In_775,In_1479);
nand U949 (N_949,In_1545,In_1587);
nand U950 (N_950,In_1198,In_2278);
nor U951 (N_951,In_378,In_516);
and U952 (N_952,In_2274,In_945);
and U953 (N_953,In_1159,In_1167);
nor U954 (N_954,In_868,In_488);
nand U955 (N_955,In_2231,In_1508);
xor U956 (N_956,In_222,In_580);
nand U957 (N_957,In_823,In_864);
nor U958 (N_958,In_1904,In_28);
xnor U959 (N_959,In_1358,In_1496);
and U960 (N_960,In_435,In_1460);
nor U961 (N_961,In_363,In_1751);
nor U962 (N_962,In_2115,In_1222);
nand U963 (N_963,In_2435,In_217);
nand U964 (N_964,In_295,In_1097);
or U965 (N_965,In_1998,In_2361);
and U966 (N_966,In_1582,In_141);
or U967 (N_967,In_2160,In_82);
xor U968 (N_968,In_119,In_1292);
or U969 (N_969,In_1325,In_2039);
or U970 (N_970,In_2310,In_156);
and U971 (N_971,In_447,In_434);
nor U972 (N_972,In_1341,In_1324);
nand U973 (N_973,In_695,In_1245);
nand U974 (N_974,In_2479,In_1038);
nand U975 (N_975,In_708,In_412);
or U976 (N_976,In_999,In_2337);
or U977 (N_977,In_1652,In_393);
xnor U978 (N_978,In_348,In_260);
xor U979 (N_979,In_2378,In_1597);
and U980 (N_980,In_1140,In_493);
nand U981 (N_981,In_1408,In_65);
and U982 (N_982,In_1380,In_2461);
and U983 (N_983,In_419,In_642);
or U984 (N_984,In_829,In_1263);
or U985 (N_985,In_1024,In_1867);
xnor U986 (N_986,In_1972,In_2204);
and U987 (N_987,In_518,In_1155);
nand U988 (N_988,In_511,In_1498);
and U989 (N_989,In_2294,In_1227);
nor U990 (N_990,In_611,In_762);
xnor U991 (N_991,In_2035,In_11);
and U992 (N_992,In_196,In_1868);
nand U993 (N_993,In_1146,In_849);
or U994 (N_994,In_1446,In_212);
nand U995 (N_995,In_1483,In_1342);
or U996 (N_996,In_325,In_1636);
or U997 (N_997,In_1078,In_1745);
and U998 (N_998,In_1825,In_116);
nand U999 (N_999,In_89,In_244);
and U1000 (N_1000,In_1230,In_648);
and U1001 (N_1001,In_1841,In_1602);
and U1002 (N_1002,In_1817,In_647);
and U1003 (N_1003,In_652,In_2434);
and U1004 (N_1004,In_1405,In_887);
xnor U1005 (N_1005,In_195,In_828);
nand U1006 (N_1006,In_449,In_856);
nand U1007 (N_1007,In_2464,In_71);
nand U1008 (N_1008,In_2229,In_912);
or U1009 (N_1009,In_1792,In_1581);
or U1010 (N_1010,In_2403,In_845);
or U1011 (N_1011,In_1104,In_836);
or U1012 (N_1012,In_1912,In_353);
xnor U1013 (N_1013,In_199,In_2400);
and U1014 (N_1014,In_704,In_826);
or U1015 (N_1015,In_2373,In_608);
nand U1016 (N_1016,In_550,In_2286);
nand U1017 (N_1017,In_2003,In_1058);
xor U1018 (N_1018,In_970,In_1554);
or U1019 (N_1019,In_898,In_2341);
xnor U1020 (N_1020,In_2249,In_1702);
and U1021 (N_1021,In_745,In_360);
nand U1022 (N_1022,In_2289,In_1684);
xor U1023 (N_1023,In_1811,In_78);
nor U1024 (N_1024,In_892,In_1474);
or U1025 (N_1025,In_75,In_64);
nand U1026 (N_1026,In_2156,In_1356);
nand U1027 (N_1027,In_2130,In_1173);
and U1028 (N_1028,In_146,In_366);
and U1029 (N_1029,In_566,In_1503);
nor U1030 (N_1030,In_657,In_721);
or U1031 (N_1031,In_1756,In_1694);
xor U1032 (N_1032,In_76,In_1970);
nor U1033 (N_1033,In_1931,In_2356);
nand U1034 (N_1034,In_323,In_675);
or U1035 (N_1035,In_1016,In_382);
or U1036 (N_1036,In_2017,In_522);
nand U1037 (N_1037,In_1076,In_2343);
and U1038 (N_1038,In_1253,In_400);
nand U1039 (N_1039,In_1893,In_953);
and U1040 (N_1040,In_1083,In_1161);
xor U1041 (N_1041,In_619,In_2234);
and U1042 (N_1042,In_1641,In_245);
or U1043 (N_1043,In_188,In_445);
and U1044 (N_1044,In_2419,In_1627);
nand U1045 (N_1045,In_736,In_197);
nor U1046 (N_1046,In_1294,In_1118);
or U1047 (N_1047,In_873,In_1964);
xnor U1048 (N_1048,In_876,In_303);
xor U1049 (N_1049,In_1343,In_47);
nand U1050 (N_1050,In_1468,In_1934);
or U1051 (N_1051,In_423,In_2031);
nor U1052 (N_1052,In_1565,In_1369);
nand U1053 (N_1053,In_2072,In_2272);
nand U1054 (N_1054,In_1464,In_298);
xnor U1055 (N_1055,In_161,In_462);
and U1056 (N_1056,In_2488,In_1573);
nand U1057 (N_1057,In_208,In_1355);
nand U1058 (N_1058,In_969,In_853);
xor U1059 (N_1059,In_555,In_2410);
nand U1060 (N_1060,In_810,In_297);
nand U1061 (N_1061,In_780,In_645);
nor U1062 (N_1062,In_2327,In_2330);
or U1063 (N_1063,In_727,In_819);
or U1064 (N_1064,In_1523,In_1361);
nand U1065 (N_1065,In_1077,In_2150);
nand U1066 (N_1066,In_1570,In_861);
or U1067 (N_1067,In_1630,In_2481);
and U1068 (N_1068,In_20,In_1297);
nand U1069 (N_1069,In_514,In_1897);
xnor U1070 (N_1070,In_814,In_248);
nor U1071 (N_1071,In_480,In_2471);
nor U1072 (N_1072,In_1878,In_878);
and U1073 (N_1073,In_1194,In_2472);
or U1074 (N_1074,In_905,In_367);
or U1075 (N_1075,In_77,In_1682);
and U1076 (N_1076,In_1815,In_407);
and U1077 (N_1077,In_1657,In_538);
nand U1078 (N_1078,In_2201,In_1531);
or U1079 (N_1079,In_585,In_661);
nand U1080 (N_1080,In_2209,In_2038);
or U1081 (N_1081,In_1296,In_117);
and U1082 (N_1082,In_1400,In_1846);
or U1083 (N_1083,In_1111,In_2452);
and U1084 (N_1084,In_1338,In_2080);
xnor U1085 (N_1085,In_2237,In_1919);
nor U1086 (N_1086,In_677,In_524);
nor U1087 (N_1087,In_1979,In_2281);
and U1088 (N_1088,In_503,In_1308);
nand U1089 (N_1089,In_865,In_405);
nor U1090 (N_1090,In_190,In_448);
xnor U1091 (N_1091,In_1707,In_123);
nor U1092 (N_1092,In_501,In_630);
or U1093 (N_1093,In_1858,In_1600);
and U1094 (N_1094,In_2441,In_1162);
nand U1095 (N_1095,In_326,In_132);
nor U1096 (N_1096,In_357,In_2397);
and U1097 (N_1097,In_40,In_277);
or U1098 (N_1098,In_332,In_564);
xnor U1099 (N_1099,In_1149,In_2313);
nor U1100 (N_1100,In_246,In_1329);
nand U1101 (N_1101,In_850,In_1061);
nand U1102 (N_1102,In_815,In_941);
nor U1103 (N_1103,In_91,In_1476);
nor U1104 (N_1104,In_527,In_1207);
nor U1105 (N_1105,In_1452,In_67);
nor U1106 (N_1106,In_2216,In_1740);
xor U1107 (N_1107,In_1663,In_95);
xnor U1108 (N_1108,In_1758,In_875);
or U1109 (N_1109,In_1794,In_539);
nand U1110 (N_1110,In_1502,In_2097);
nor U1111 (N_1111,In_201,In_577);
nand U1112 (N_1112,In_460,In_2270);
nor U1113 (N_1113,In_2242,In_264);
nor U1114 (N_1114,In_1621,In_541);
nor U1115 (N_1115,In_1976,In_869);
and U1116 (N_1116,In_628,In_2251);
or U1117 (N_1117,In_2149,In_1094);
nand U1118 (N_1118,In_1580,In_693);
nand U1119 (N_1119,In_1182,In_1971);
or U1120 (N_1120,In_992,In_352);
nor U1121 (N_1121,In_218,In_1509);
nor U1122 (N_1122,In_759,In_336);
nor U1123 (N_1123,In_61,In_1743);
and U1124 (N_1124,In_1891,In_250);
xor U1125 (N_1125,In_1594,In_846);
nand U1126 (N_1126,In_491,In_1932);
nor U1127 (N_1127,In_1529,In_1423);
nand U1128 (N_1128,In_1289,In_1984);
nor U1129 (N_1129,In_2004,In_2236);
nand U1130 (N_1130,In_1643,In_1480);
or U1131 (N_1131,In_854,In_1485);
and U1132 (N_1132,In_1362,In_1044);
and U1133 (N_1133,In_2056,In_926);
nor U1134 (N_1134,In_705,In_446);
xnor U1135 (N_1135,In_800,In_2260);
nor U1136 (N_1136,In_881,In_2136);
xor U1137 (N_1137,In_792,In_2409);
nand U1138 (N_1138,In_2075,In_1836);
xnor U1139 (N_1139,In_2127,In_2068);
xnor U1140 (N_1140,In_567,In_338);
or U1141 (N_1141,In_534,In_2008);
nor U1142 (N_1142,In_725,In_1251);
nor U1143 (N_1143,In_2333,In_1561);
xnor U1144 (N_1144,In_517,In_376);
nor U1145 (N_1145,In_1982,In_793);
and U1146 (N_1146,In_1210,In_2301);
or U1147 (N_1147,In_1397,In_917);
and U1148 (N_1148,In_2355,In_533);
nand U1149 (N_1149,In_1741,In_565);
and U1150 (N_1150,In_12,In_1865);
or U1151 (N_1151,In_2103,In_1555);
or U1152 (N_1152,In_2060,In_1888);
nor U1153 (N_1153,In_2385,In_1577);
and U1154 (N_1154,In_421,In_2093);
nand U1155 (N_1155,In_383,In_597);
or U1156 (N_1156,In_1850,In_1804);
nand U1157 (N_1157,In_1025,In_740);
nor U1158 (N_1158,In_2412,In_1096);
nor U1159 (N_1159,In_1348,In_2316);
or U1160 (N_1160,In_1150,In_984);
and U1161 (N_1161,In_1571,In_586);
nand U1162 (N_1162,In_2499,In_225);
nand U1163 (N_1163,In_1034,In_1871);
nand U1164 (N_1164,In_634,In_339);
nand U1165 (N_1165,In_831,In_1409);
nor U1166 (N_1166,In_1612,In_994);
nand U1167 (N_1167,In_205,In_688);
nor U1168 (N_1168,In_1798,In_101);
and U1169 (N_1169,In_1309,In_1193);
nand U1170 (N_1170,In_2181,In_1179);
nor U1171 (N_1171,In_1651,In_392);
nor U1172 (N_1172,In_749,In_374);
or U1173 (N_1173,In_497,In_1997);
or U1174 (N_1174,In_885,In_893);
xor U1175 (N_1175,In_1205,In_751);
and U1176 (N_1176,In_1533,In_1655);
xor U1177 (N_1177,In_2124,In_2474);
nor U1178 (N_1178,In_1649,In_1166);
nand U1179 (N_1179,In_2198,In_954);
or U1180 (N_1180,In_1385,In_1693);
and U1181 (N_1181,In_1880,In_456);
or U1182 (N_1182,In_399,In_781);
and U1183 (N_1183,In_2148,In_2490);
and U1184 (N_1184,In_569,In_2405);
and U1185 (N_1185,In_1197,In_315);
nand U1186 (N_1186,In_812,In_1784);
and U1187 (N_1187,In_2175,In_334);
nor U1188 (N_1188,In_1139,In_2152);
and U1189 (N_1189,In_1862,In_726);
nand U1190 (N_1190,In_1814,In_1936);
and U1191 (N_1191,In_1281,In_995);
or U1192 (N_1192,In_1022,In_1766);
nor U1193 (N_1193,In_1497,In_1185);
nand U1194 (N_1194,In_1390,In_1091);
or U1195 (N_1195,In_351,In_1633);
nand U1196 (N_1196,In_1084,In_717);
nand U1197 (N_1197,In_1217,In_2444);
xor U1198 (N_1198,In_1314,In_2024);
or U1199 (N_1199,In_112,In_879);
nand U1200 (N_1200,In_157,In_1430);
and U1201 (N_1201,In_202,In_1072);
or U1202 (N_1202,In_1370,In_1765);
xor U1203 (N_1203,In_1619,In_1898);
and U1204 (N_1204,In_835,In_312);
nor U1205 (N_1205,In_757,In_789);
nor U1206 (N_1206,In_1987,In_1353);
nand U1207 (N_1207,In_1616,In_2247);
nand U1208 (N_1208,In_455,In_461);
nor U1209 (N_1209,In_454,In_1270);
nor U1210 (N_1210,In_891,In_302);
and U1211 (N_1211,In_2048,In_1267);
nand U1212 (N_1212,In_2408,In_1831);
and U1213 (N_1213,In_306,In_1986);
xor U1214 (N_1214,In_1277,In_1317);
and U1215 (N_1215,In_1445,In_1439);
xnor U1216 (N_1216,In_301,In_1802);
nand U1217 (N_1217,In_437,In_204);
nor U1218 (N_1218,In_532,In_1357);
nor U1219 (N_1219,In_2401,In_805);
or U1220 (N_1220,In_838,In_1884);
nand U1221 (N_1221,In_578,In_441);
or U1222 (N_1222,In_595,In_379);
or U1223 (N_1223,In_949,In_2178);
or U1224 (N_1224,In_722,In_1233);
and U1225 (N_1225,In_1339,In_2121);
xor U1226 (N_1226,In_924,In_1830);
or U1227 (N_1227,In_1120,In_147);
and U1228 (N_1228,In_1434,In_1311);
xnor U1229 (N_1229,In_263,In_635);
or U1230 (N_1230,In_193,In_909);
xnor U1231 (N_1231,In_542,In_2417);
or U1232 (N_1232,In_1900,In_1181);
or U1233 (N_1233,In_1683,In_1761);
xnor U1234 (N_1234,In_507,In_1316);
and U1235 (N_1235,In_309,In_1506);
nor U1236 (N_1236,In_2329,In_2392);
and U1237 (N_1237,In_973,In_2147);
and U1238 (N_1238,In_788,In_1706);
nor U1239 (N_1239,In_558,In_1688);
xor U1240 (N_1240,In_152,In_714);
or U1241 (N_1241,In_242,In_1601);
or U1242 (N_1242,In_1455,In_2407);
and U1243 (N_1243,In_1382,In_1667);
nor U1244 (N_1244,In_282,In_1552);
nand U1245 (N_1245,In_1935,In_1261);
nand U1246 (N_1246,In_1387,In_1414);
xor U1247 (N_1247,In_1634,In_1);
nand U1248 (N_1248,In_783,In_2393);
nor U1249 (N_1249,In_702,In_1407);
and U1250 (N_1250,In_1944,In_2003);
nor U1251 (N_1251,In_135,In_1603);
or U1252 (N_1252,In_886,In_1454);
nor U1253 (N_1253,In_1542,In_1701);
nor U1254 (N_1254,In_2136,In_2043);
and U1255 (N_1255,In_765,In_1676);
nor U1256 (N_1256,In_1733,In_418);
and U1257 (N_1257,In_2395,In_89);
nand U1258 (N_1258,In_1915,In_1560);
nor U1259 (N_1259,In_1509,In_991);
or U1260 (N_1260,In_1121,In_2279);
nor U1261 (N_1261,In_1148,In_792);
nand U1262 (N_1262,In_317,In_193);
nand U1263 (N_1263,In_52,In_2344);
xor U1264 (N_1264,In_317,In_980);
or U1265 (N_1265,In_191,In_511);
xor U1266 (N_1266,In_308,In_142);
nand U1267 (N_1267,In_2024,In_1721);
or U1268 (N_1268,In_916,In_726);
nor U1269 (N_1269,In_884,In_232);
nor U1270 (N_1270,In_1578,In_1096);
nor U1271 (N_1271,In_997,In_645);
nand U1272 (N_1272,In_677,In_2293);
nand U1273 (N_1273,In_1473,In_1885);
nor U1274 (N_1274,In_663,In_136);
nand U1275 (N_1275,In_2134,In_716);
nand U1276 (N_1276,In_1364,In_225);
or U1277 (N_1277,In_2240,In_445);
and U1278 (N_1278,In_2307,In_1391);
nand U1279 (N_1279,In_116,In_531);
nand U1280 (N_1280,In_1461,In_1623);
nand U1281 (N_1281,In_533,In_1583);
and U1282 (N_1282,In_2056,In_9);
and U1283 (N_1283,In_485,In_2343);
or U1284 (N_1284,In_1250,In_1231);
or U1285 (N_1285,In_285,In_221);
and U1286 (N_1286,In_236,In_499);
nor U1287 (N_1287,In_2282,In_1295);
and U1288 (N_1288,In_2401,In_1121);
nand U1289 (N_1289,In_2343,In_1363);
xor U1290 (N_1290,In_2359,In_106);
and U1291 (N_1291,In_1582,In_1366);
and U1292 (N_1292,In_938,In_801);
or U1293 (N_1293,In_1896,In_1217);
and U1294 (N_1294,In_1193,In_459);
and U1295 (N_1295,In_951,In_1924);
xor U1296 (N_1296,In_444,In_2189);
xor U1297 (N_1297,In_745,In_368);
and U1298 (N_1298,In_432,In_517);
nand U1299 (N_1299,In_978,In_96);
xor U1300 (N_1300,In_2468,In_1379);
nand U1301 (N_1301,In_1009,In_2053);
xor U1302 (N_1302,In_29,In_2100);
and U1303 (N_1303,In_1184,In_423);
nand U1304 (N_1304,In_1494,In_829);
or U1305 (N_1305,In_2264,In_1395);
and U1306 (N_1306,In_1482,In_532);
xnor U1307 (N_1307,In_730,In_831);
nor U1308 (N_1308,In_428,In_2336);
nor U1309 (N_1309,In_2107,In_590);
or U1310 (N_1310,In_1367,In_2442);
nand U1311 (N_1311,In_284,In_964);
and U1312 (N_1312,In_524,In_137);
nand U1313 (N_1313,In_2077,In_1116);
nor U1314 (N_1314,In_2455,In_1988);
and U1315 (N_1315,In_2273,In_1154);
xnor U1316 (N_1316,In_188,In_2156);
nand U1317 (N_1317,In_1032,In_216);
and U1318 (N_1318,In_2330,In_1950);
xor U1319 (N_1319,In_1711,In_1366);
nand U1320 (N_1320,In_2334,In_296);
and U1321 (N_1321,In_91,In_1946);
and U1322 (N_1322,In_2472,In_765);
nor U1323 (N_1323,In_411,In_1951);
nor U1324 (N_1324,In_102,In_2048);
nand U1325 (N_1325,In_2259,In_2200);
or U1326 (N_1326,In_484,In_603);
nand U1327 (N_1327,In_221,In_1959);
nand U1328 (N_1328,In_69,In_1817);
or U1329 (N_1329,In_2338,In_588);
nand U1330 (N_1330,In_77,In_354);
nor U1331 (N_1331,In_1863,In_2386);
xnor U1332 (N_1332,In_227,In_2010);
nor U1333 (N_1333,In_2355,In_26);
nand U1334 (N_1334,In_182,In_1989);
or U1335 (N_1335,In_936,In_963);
or U1336 (N_1336,In_882,In_1415);
nor U1337 (N_1337,In_717,In_910);
or U1338 (N_1338,In_796,In_258);
and U1339 (N_1339,In_2323,In_2083);
or U1340 (N_1340,In_1644,In_1434);
nand U1341 (N_1341,In_628,In_2263);
nand U1342 (N_1342,In_2109,In_1923);
nor U1343 (N_1343,In_2484,In_639);
or U1344 (N_1344,In_1281,In_1446);
nor U1345 (N_1345,In_1782,In_2433);
nand U1346 (N_1346,In_530,In_2292);
or U1347 (N_1347,In_1507,In_919);
nor U1348 (N_1348,In_1388,In_1207);
or U1349 (N_1349,In_2275,In_2377);
or U1350 (N_1350,In_1628,In_2014);
nor U1351 (N_1351,In_1608,In_2069);
and U1352 (N_1352,In_1554,In_2393);
nand U1353 (N_1353,In_1269,In_811);
xnor U1354 (N_1354,In_471,In_1164);
and U1355 (N_1355,In_1874,In_411);
nand U1356 (N_1356,In_140,In_815);
xor U1357 (N_1357,In_792,In_1796);
nor U1358 (N_1358,In_1612,In_1860);
nand U1359 (N_1359,In_1671,In_1851);
nor U1360 (N_1360,In_2178,In_231);
or U1361 (N_1361,In_1963,In_106);
and U1362 (N_1362,In_23,In_546);
or U1363 (N_1363,In_1378,In_1106);
xor U1364 (N_1364,In_672,In_1458);
and U1365 (N_1365,In_1288,In_613);
nor U1366 (N_1366,In_148,In_2017);
nor U1367 (N_1367,In_41,In_2388);
nand U1368 (N_1368,In_2075,In_1529);
or U1369 (N_1369,In_2184,In_1478);
nor U1370 (N_1370,In_248,In_301);
nand U1371 (N_1371,In_1918,In_1464);
nand U1372 (N_1372,In_867,In_570);
xnor U1373 (N_1373,In_106,In_2385);
or U1374 (N_1374,In_2338,In_513);
nand U1375 (N_1375,In_2073,In_1329);
nor U1376 (N_1376,In_638,In_1623);
nand U1377 (N_1377,In_552,In_1621);
and U1378 (N_1378,In_741,In_1135);
or U1379 (N_1379,In_2491,In_2019);
nand U1380 (N_1380,In_326,In_2159);
nand U1381 (N_1381,In_711,In_1643);
or U1382 (N_1382,In_1387,In_1314);
nor U1383 (N_1383,In_1934,In_597);
xor U1384 (N_1384,In_251,In_2145);
and U1385 (N_1385,In_1242,In_1358);
and U1386 (N_1386,In_264,In_571);
nand U1387 (N_1387,In_1474,In_2205);
or U1388 (N_1388,In_2477,In_1054);
nor U1389 (N_1389,In_908,In_416);
nand U1390 (N_1390,In_1501,In_52);
or U1391 (N_1391,In_194,In_1353);
nor U1392 (N_1392,In_118,In_2392);
and U1393 (N_1393,In_1699,In_125);
nor U1394 (N_1394,In_546,In_1347);
nor U1395 (N_1395,In_1437,In_2339);
or U1396 (N_1396,In_1486,In_547);
nor U1397 (N_1397,In_514,In_858);
nor U1398 (N_1398,In_1651,In_2232);
and U1399 (N_1399,In_932,In_2383);
or U1400 (N_1400,In_2087,In_1342);
nand U1401 (N_1401,In_1448,In_424);
and U1402 (N_1402,In_2299,In_1223);
or U1403 (N_1403,In_1422,In_920);
xor U1404 (N_1404,In_2290,In_937);
nand U1405 (N_1405,In_2296,In_2205);
and U1406 (N_1406,In_78,In_2490);
nand U1407 (N_1407,In_308,In_1970);
xnor U1408 (N_1408,In_1838,In_1413);
xor U1409 (N_1409,In_896,In_79);
and U1410 (N_1410,In_220,In_2062);
nor U1411 (N_1411,In_1404,In_14);
or U1412 (N_1412,In_1564,In_1227);
nor U1413 (N_1413,In_1065,In_1032);
or U1414 (N_1414,In_2156,In_517);
xnor U1415 (N_1415,In_1378,In_2020);
and U1416 (N_1416,In_1445,In_920);
or U1417 (N_1417,In_1956,In_2208);
nand U1418 (N_1418,In_541,In_344);
and U1419 (N_1419,In_1737,In_2399);
and U1420 (N_1420,In_1426,In_321);
or U1421 (N_1421,In_493,In_398);
xnor U1422 (N_1422,In_2159,In_1262);
or U1423 (N_1423,In_2423,In_1466);
or U1424 (N_1424,In_1882,In_90);
nand U1425 (N_1425,In_1045,In_291);
nand U1426 (N_1426,In_1689,In_1648);
nor U1427 (N_1427,In_268,In_13);
xnor U1428 (N_1428,In_1279,In_2309);
or U1429 (N_1429,In_2330,In_393);
nor U1430 (N_1430,In_1768,In_1959);
or U1431 (N_1431,In_1513,In_155);
nand U1432 (N_1432,In_1462,In_2491);
or U1433 (N_1433,In_1525,In_1231);
xnor U1434 (N_1434,In_646,In_398);
nor U1435 (N_1435,In_1926,In_521);
nand U1436 (N_1436,In_777,In_31);
nor U1437 (N_1437,In_895,In_1973);
nand U1438 (N_1438,In_2441,In_676);
nor U1439 (N_1439,In_2348,In_1257);
or U1440 (N_1440,In_141,In_118);
or U1441 (N_1441,In_819,In_2389);
or U1442 (N_1442,In_2364,In_1049);
nor U1443 (N_1443,In_1379,In_945);
xnor U1444 (N_1444,In_1202,In_1336);
nor U1445 (N_1445,In_283,In_427);
or U1446 (N_1446,In_1054,In_2363);
nand U1447 (N_1447,In_184,In_1740);
nand U1448 (N_1448,In_2367,In_1846);
nor U1449 (N_1449,In_2232,In_1150);
and U1450 (N_1450,In_841,In_2474);
or U1451 (N_1451,In_4,In_1909);
xnor U1452 (N_1452,In_1515,In_2087);
nand U1453 (N_1453,In_1868,In_1295);
xor U1454 (N_1454,In_2280,In_2265);
nor U1455 (N_1455,In_1802,In_1924);
or U1456 (N_1456,In_499,In_2186);
nor U1457 (N_1457,In_240,In_1651);
nor U1458 (N_1458,In_895,In_1414);
xor U1459 (N_1459,In_575,In_2004);
or U1460 (N_1460,In_2112,In_1235);
and U1461 (N_1461,In_275,In_1034);
and U1462 (N_1462,In_157,In_2414);
nor U1463 (N_1463,In_635,In_1215);
nand U1464 (N_1464,In_988,In_1793);
nor U1465 (N_1465,In_608,In_844);
nor U1466 (N_1466,In_2057,In_185);
and U1467 (N_1467,In_1084,In_863);
nand U1468 (N_1468,In_223,In_2023);
nor U1469 (N_1469,In_966,In_817);
or U1470 (N_1470,In_2285,In_1146);
or U1471 (N_1471,In_1186,In_1485);
or U1472 (N_1472,In_2296,In_1543);
or U1473 (N_1473,In_691,In_834);
nor U1474 (N_1474,In_551,In_2157);
or U1475 (N_1475,In_773,In_1787);
xnor U1476 (N_1476,In_172,In_380);
nor U1477 (N_1477,In_383,In_704);
and U1478 (N_1478,In_2495,In_1965);
nand U1479 (N_1479,In_37,In_1133);
nand U1480 (N_1480,In_1672,In_1497);
nor U1481 (N_1481,In_1219,In_289);
nor U1482 (N_1482,In_1606,In_225);
and U1483 (N_1483,In_2304,In_827);
xnor U1484 (N_1484,In_514,In_549);
and U1485 (N_1485,In_2418,In_1451);
and U1486 (N_1486,In_1479,In_1345);
nand U1487 (N_1487,In_880,In_1044);
and U1488 (N_1488,In_1781,In_1616);
nor U1489 (N_1489,In_2135,In_119);
nand U1490 (N_1490,In_70,In_1531);
and U1491 (N_1491,In_1187,In_1177);
nor U1492 (N_1492,In_42,In_319);
xor U1493 (N_1493,In_1288,In_1430);
or U1494 (N_1494,In_2096,In_249);
and U1495 (N_1495,In_1981,In_283);
and U1496 (N_1496,In_1791,In_1017);
nand U1497 (N_1497,In_2307,In_1530);
nand U1498 (N_1498,In_536,In_2265);
nor U1499 (N_1499,In_971,In_2436);
nor U1500 (N_1500,In_1533,In_1684);
nor U1501 (N_1501,In_1740,In_1058);
nor U1502 (N_1502,In_1960,In_603);
or U1503 (N_1503,In_409,In_2237);
and U1504 (N_1504,In_624,In_2152);
nand U1505 (N_1505,In_2489,In_141);
xor U1506 (N_1506,In_846,In_382);
nand U1507 (N_1507,In_2209,In_1609);
nand U1508 (N_1508,In_2452,In_1897);
nor U1509 (N_1509,In_1873,In_1296);
nor U1510 (N_1510,In_2093,In_1499);
nand U1511 (N_1511,In_2028,In_1759);
or U1512 (N_1512,In_378,In_2283);
nor U1513 (N_1513,In_2454,In_88);
and U1514 (N_1514,In_259,In_1933);
or U1515 (N_1515,In_1586,In_2478);
nand U1516 (N_1516,In_1644,In_1553);
nand U1517 (N_1517,In_1612,In_699);
nand U1518 (N_1518,In_1906,In_1972);
nand U1519 (N_1519,In_2146,In_2244);
nor U1520 (N_1520,In_1019,In_1221);
or U1521 (N_1521,In_2012,In_1510);
or U1522 (N_1522,In_1147,In_296);
nand U1523 (N_1523,In_1913,In_1520);
or U1524 (N_1524,In_2210,In_1638);
nand U1525 (N_1525,In_2103,In_1820);
nor U1526 (N_1526,In_2047,In_263);
nand U1527 (N_1527,In_2017,In_1300);
nor U1528 (N_1528,In_1696,In_2133);
and U1529 (N_1529,In_574,In_500);
nor U1530 (N_1530,In_522,In_286);
and U1531 (N_1531,In_899,In_684);
or U1532 (N_1532,In_1852,In_85);
and U1533 (N_1533,In_1918,In_1617);
nor U1534 (N_1534,In_139,In_1529);
nand U1535 (N_1535,In_754,In_1310);
or U1536 (N_1536,In_459,In_2);
or U1537 (N_1537,In_2014,In_1064);
nand U1538 (N_1538,In_1640,In_403);
or U1539 (N_1539,In_2148,In_196);
and U1540 (N_1540,In_495,In_2020);
xor U1541 (N_1541,In_1792,In_708);
nand U1542 (N_1542,In_923,In_2201);
nor U1543 (N_1543,In_965,In_483);
or U1544 (N_1544,In_287,In_1303);
nand U1545 (N_1545,In_1274,In_902);
or U1546 (N_1546,In_1595,In_1059);
and U1547 (N_1547,In_1170,In_376);
and U1548 (N_1548,In_1733,In_559);
nand U1549 (N_1549,In_264,In_680);
nor U1550 (N_1550,In_296,In_2007);
and U1551 (N_1551,In_1566,In_1745);
or U1552 (N_1552,In_943,In_1228);
nor U1553 (N_1553,In_118,In_1439);
nor U1554 (N_1554,In_2381,In_257);
nand U1555 (N_1555,In_1066,In_1901);
xnor U1556 (N_1556,In_693,In_1897);
nor U1557 (N_1557,In_839,In_2447);
or U1558 (N_1558,In_854,In_657);
and U1559 (N_1559,In_2449,In_661);
or U1560 (N_1560,In_1944,In_721);
nand U1561 (N_1561,In_239,In_3);
and U1562 (N_1562,In_1277,In_1305);
nor U1563 (N_1563,In_431,In_1766);
nor U1564 (N_1564,In_1006,In_978);
xor U1565 (N_1565,In_1442,In_548);
nor U1566 (N_1566,In_941,In_1301);
xnor U1567 (N_1567,In_2367,In_2418);
nor U1568 (N_1568,In_1901,In_2468);
and U1569 (N_1569,In_2067,In_898);
and U1570 (N_1570,In_1520,In_1761);
nor U1571 (N_1571,In_2024,In_2416);
xor U1572 (N_1572,In_510,In_898);
or U1573 (N_1573,In_1604,In_1711);
or U1574 (N_1574,In_1468,In_1931);
nand U1575 (N_1575,In_2031,In_1732);
and U1576 (N_1576,In_1722,In_1719);
and U1577 (N_1577,In_220,In_543);
and U1578 (N_1578,In_250,In_1113);
or U1579 (N_1579,In_684,In_1177);
and U1580 (N_1580,In_2111,In_1394);
nor U1581 (N_1581,In_87,In_772);
and U1582 (N_1582,In_1537,In_1115);
and U1583 (N_1583,In_1444,In_233);
nor U1584 (N_1584,In_1195,In_1278);
and U1585 (N_1585,In_2116,In_614);
and U1586 (N_1586,In_992,In_804);
nand U1587 (N_1587,In_1273,In_1177);
and U1588 (N_1588,In_2107,In_985);
and U1589 (N_1589,In_2498,In_1398);
and U1590 (N_1590,In_144,In_2416);
or U1591 (N_1591,In_772,In_567);
and U1592 (N_1592,In_1870,In_22);
xor U1593 (N_1593,In_2232,In_133);
or U1594 (N_1594,In_939,In_182);
and U1595 (N_1595,In_2142,In_1231);
nand U1596 (N_1596,In_2418,In_1278);
nand U1597 (N_1597,In_1009,In_1410);
nor U1598 (N_1598,In_2318,In_778);
xor U1599 (N_1599,In_1523,In_1488);
and U1600 (N_1600,In_785,In_1193);
and U1601 (N_1601,In_929,In_996);
and U1602 (N_1602,In_2352,In_1495);
and U1603 (N_1603,In_2451,In_537);
nand U1604 (N_1604,In_1728,In_2370);
nor U1605 (N_1605,In_1378,In_2435);
and U1606 (N_1606,In_2147,In_316);
nor U1607 (N_1607,In_1656,In_2063);
or U1608 (N_1608,In_367,In_1424);
nor U1609 (N_1609,In_355,In_575);
xor U1610 (N_1610,In_1756,In_569);
nand U1611 (N_1611,In_1579,In_872);
or U1612 (N_1612,In_2241,In_1801);
and U1613 (N_1613,In_554,In_1304);
or U1614 (N_1614,In_1188,In_2182);
or U1615 (N_1615,In_1075,In_309);
nand U1616 (N_1616,In_2179,In_2065);
and U1617 (N_1617,In_1890,In_1168);
nand U1618 (N_1618,In_2060,In_729);
and U1619 (N_1619,In_1806,In_324);
nor U1620 (N_1620,In_2249,In_2276);
nor U1621 (N_1621,In_440,In_2322);
or U1622 (N_1622,In_918,In_795);
and U1623 (N_1623,In_1861,In_855);
nor U1624 (N_1624,In_1629,In_1926);
or U1625 (N_1625,In_982,In_2048);
nor U1626 (N_1626,In_298,In_1703);
xor U1627 (N_1627,In_731,In_733);
and U1628 (N_1628,In_2344,In_2090);
nand U1629 (N_1629,In_2173,In_2123);
or U1630 (N_1630,In_835,In_2461);
nor U1631 (N_1631,In_2467,In_531);
nor U1632 (N_1632,In_496,In_826);
and U1633 (N_1633,In_1206,In_136);
nand U1634 (N_1634,In_176,In_114);
nor U1635 (N_1635,In_959,In_1408);
xnor U1636 (N_1636,In_89,In_1625);
and U1637 (N_1637,In_314,In_288);
and U1638 (N_1638,In_435,In_413);
or U1639 (N_1639,In_803,In_2141);
and U1640 (N_1640,In_1115,In_1634);
and U1641 (N_1641,In_1076,In_621);
nor U1642 (N_1642,In_184,In_139);
nand U1643 (N_1643,In_2134,In_1654);
or U1644 (N_1644,In_839,In_189);
nand U1645 (N_1645,In_765,In_1866);
or U1646 (N_1646,In_818,In_1334);
nor U1647 (N_1647,In_977,In_200);
xor U1648 (N_1648,In_1590,In_265);
and U1649 (N_1649,In_1770,In_1673);
and U1650 (N_1650,In_258,In_390);
and U1651 (N_1651,In_1147,In_435);
nand U1652 (N_1652,In_800,In_1088);
nor U1653 (N_1653,In_776,In_677);
nor U1654 (N_1654,In_245,In_1875);
nor U1655 (N_1655,In_2203,In_1762);
and U1656 (N_1656,In_2295,In_1802);
or U1657 (N_1657,In_1870,In_839);
nand U1658 (N_1658,In_1119,In_2302);
and U1659 (N_1659,In_1991,In_2362);
nor U1660 (N_1660,In_1794,In_1212);
xnor U1661 (N_1661,In_1648,In_47);
and U1662 (N_1662,In_361,In_993);
nand U1663 (N_1663,In_643,In_1561);
nor U1664 (N_1664,In_817,In_217);
or U1665 (N_1665,In_259,In_1467);
nor U1666 (N_1666,In_215,In_2154);
or U1667 (N_1667,In_2253,In_1730);
or U1668 (N_1668,In_40,In_2022);
and U1669 (N_1669,In_110,In_1562);
and U1670 (N_1670,In_434,In_139);
or U1671 (N_1671,In_2419,In_1244);
or U1672 (N_1672,In_864,In_167);
nand U1673 (N_1673,In_2027,In_1933);
or U1674 (N_1674,In_1526,In_1891);
nor U1675 (N_1675,In_1238,In_295);
or U1676 (N_1676,In_2111,In_2227);
nor U1677 (N_1677,In_1080,In_1228);
and U1678 (N_1678,In_1080,In_1092);
nand U1679 (N_1679,In_63,In_618);
or U1680 (N_1680,In_2053,In_2366);
nor U1681 (N_1681,In_1949,In_101);
nor U1682 (N_1682,In_2270,In_860);
or U1683 (N_1683,In_1977,In_1386);
nor U1684 (N_1684,In_340,In_712);
nand U1685 (N_1685,In_218,In_1950);
and U1686 (N_1686,In_631,In_2494);
and U1687 (N_1687,In_1568,In_1885);
or U1688 (N_1688,In_1855,In_615);
or U1689 (N_1689,In_1572,In_2356);
and U1690 (N_1690,In_817,In_1996);
xnor U1691 (N_1691,In_1901,In_788);
and U1692 (N_1692,In_1825,In_1419);
xnor U1693 (N_1693,In_2300,In_430);
nand U1694 (N_1694,In_66,In_501);
or U1695 (N_1695,In_2433,In_383);
nand U1696 (N_1696,In_1560,In_2353);
xnor U1697 (N_1697,In_2086,In_549);
nor U1698 (N_1698,In_1765,In_1973);
nand U1699 (N_1699,In_1752,In_708);
or U1700 (N_1700,In_157,In_560);
nor U1701 (N_1701,In_2298,In_524);
and U1702 (N_1702,In_679,In_711);
nor U1703 (N_1703,In_1499,In_1436);
xor U1704 (N_1704,In_1405,In_37);
or U1705 (N_1705,In_2285,In_1001);
nor U1706 (N_1706,In_278,In_2493);
xnor U1707 (N_1707,In_792,In_702);
or U1708 (N_1708,In_1775,In_576);
nand U1709 (N_1709,In_1451,In_386);
and U1710 (N_1710,In_1015,In_2390);
nor U1711 (N_1711,In_528,In_15);
nand U1712 (N_1712,In_1736,In_1656);
or U1713 (N_1713,In_1313,In_1894);
nand U1714 (N_1714,In_2238,In_2368);
or U1715 (N_1715,In_767,In_1389);
and U1716 (N_1716,In_1414,In_489);
nand U1717 (N_1717,In_948,In_1292);
and U1718 (N_1718,In_1809,In_65);
and U1719 (N_1719,In_1505,In_989);
or U1720 (N_1720,In_157,In_2087);
nand U1721 (N_1721,In_1568,In_525);
nand U1722 (N_1722,In_637,In_487);
nor U1723 (N_1723,In_1274,In_333);
or U1724 (N_1724,In_2194,In_1745);
and U1725 (N_1725,In_1756,In_1054);
nand U1726 (N_1726,In_1771,In_1227);
or U1727 (N_1727,In_2001,In_1834);
and U1728 (N_1728,In_677,In_260);
nor U1729 (N_1729,In_2081,In_2145);
nand U1730 (N_1730,In_1052,In_969);
xor U1731 (N_1731,In_2231,In_2440);
nor U1732 (N_1732,In_975,In_2121);
nand U1733 (N_1733,In_2001,In_2382);
nand U1734 (N_1734,In_1296,In_2048);
and U1735 (N_1735,In_745,In_2269);
and U1736 (N_1736,In_2364,In_747);
xor U1737 (N_1737,In_1834,In_1334);
nor U1738 (N_1738,In_4,In_1195);
or U1739 (N_1739,In_1881,In_2315);
and U1740 (N_1740,In_2192,In_742);
nand U1741 (N_1741,In_553,In_254);
nor U1742 (N_1742,In_1796,In_1395);
xor U1743 (N_1743,In_214,In_334);
xnor U1744 (N_1744,In_931,In_569);
nor U1745 (N_1745,In_71,In_18);
xor U1746 (N_1746,In_1189,In_552);
nand U1747 (N_1747,In_1354,In_2199);
nor U1748 (N_1748,In_377,In_2302);
xnor U1749 (N_1749,In_2289,In_2035);
and U1750 (N_1750,In_949,In_1018);
and U1751 (N_1751,In_234,In_1762);
nor U1752 (N_1752,In_133,In_811);
and U1753 (N_1753,In_474,In_1685);
or U1754 (N_1754,In_1594,In_945);
xnor U1755 (N_1755,In_470,In_1029);
nor U1756 (N_1756,In_1479,In_1315);
or U1757 (N_1757,In_2047,In_703);
nor U1758 (N_1758,In_1725,In_1324);
or U1759 (N_1759,In_1711,In_8);
nor U1760 (N_1760,In_853,In_1433);
nand U1761 (N_1761,In_491,In_788);
or U1762 (N_1762,In_710,In_47);
and U1763 (N_1763,In_1874,In_246);
nor U1764 (N_1764,In_246,In_1878);
nand U1765 (N_1765,In_1542,In_1331);
nand U1766 (N_1766,In_186,In_847);
or U1767 (N_1767,In_1275,In_1843);
and U1768 (N_1768,In_877,In_1572);
or U1769 (N_1769,In_2498,In_236);
nand U1770 (N_1770,In_276,In_1174);
or U1771 (N_1771,In_242,In_955);
nor U1772 (N_1772,In_895,In_234);
nor U1773 (N_1773,In_1496,In_57);
nand U1774 (N_1774,In_1215,In_225);
xor U1775 (N_1775,In_1509,In_1668);
nand U1776 (N_1776,In_2397,In_1132);
nand U1777 (N_1777,In_1142,In_2299);
nand U1778 (N_1778,In_2121,In_639);
nand U1779 (N_1779,In_2156,In_279);
and U1780 (N_1780,In_814,In_624);
or U1781 (N_1781,In_1728,In_1487);
nand U1782 (N_1782,In_2242,In_1881);
or U1783 (N_1783,In_1828,In_627);
nand U1784 (N_1784,In_958,In_2357);
nor U1785 (N_1785,In_2105,In_295);
or U1786 (N_1786,In_1880,In_181);
nand U1787 (N_1787,In_1715,In_976);
nor U1788 (N_1788,In_1597,In_760);
nor U1789 (N_1789,In_1065,In_838);
and U1790 (N_1790,In_1934,In_1500);
nor U1791 (N_1791,In_679,In_1370);
or U1792 (N_1792,In_2017,In_1745);
nand U1793 (N_1793,In_2055,In_1369);
nand U1794 (N_1794,In_1045,In_2334);
and U1795 (N_1795,In_2206,In_755);
nand U1796 (N_1796,In_2253,In_953);
xnor U1797 (N_1797,In_128,In_227);
xor U1798 (N_1798,In_1598,In_2369);
or U1799 (N_1799,In_411,In_2423);
nand U1800 (N_1800,In_2079,In_161);
or U1801 (N_1801,In_2464,In_2469);
and U1802 (N_1802,In_1297,In_1147);
nor U1803 (N_1803,In_7,In_162);
and U1804 (N_1804,In_251,In_1675);
nand U1805 (N_1805,In_2389,In_2468);
nor U1806 (N_1806,In_1656,In_1194);
nor U1807 (N_1807,In_177,In_2376);
nand U1808 (N_1808,In_1938,In_162);
and U1809 (N_1809,In_35,In_814);
nand U1810 (N_1810,In_1721,In_1339);
nand U1811 (N_1811,In_721,In_1095);
nand U1812 (N_1812,In_447,In_13);
and U1813 (N_1813,In_2225,In_702);
xnor U1814 (N_1814,In_2150,In_1142);
or U1815 (N_1815,In_2102,In_1253);
nand U1816 (N_1816,In_2487,In_1172);
nor U1817 (N_1817,In_1465,In_559);
and U1818 (N_1818,In_1573,In_2200);
xor U1819 (N_1819,In_1309,In_792);
nand U1820 (N_1820,In_1644,In_1213);
or U1821 (N_1821,In_1169,In_730);
nor U1822 (N_1822,In_1801,In_2193);
nor U1823 (N_1823,In_1749,In_165);
nand U1824 (N_1824,In_2309,In_1385);
nand U1825 (N_1825,In_622,In_1545);
nand U1826 (N_1826,In_269,In_1855);
and U1827 (N_1827,In_339,In_292);
or U1828 (N_1828,In_1686,In_783);
nand U1829 (N_1829,In_479,In_1840);
and U1830 (N_1830,In_425,In_495);
nor U1831 (N_1831,In_2485,In_2275);
and U1832 (N_1832,In_335,In_1247);
or U1833 (N_1833,In_1716,In_1345);
and U1834 (N_1834,In_1811,In_5);
or U1835 (N_1835,In_277,In_833);
nor U1836 (N_1836,In_1430,In_280);
nand U1837 (N_1837,In_1711,In_1013);
and U1838 (N_1838,In_1586,In_1432);
or U1839 (N_1839,In_271,In_1607);
nand U1840 (N_1840,In_1052,In_655);
or U1841 (N_1841,In_2015,In_2391);
nor U1842 (N_1842,In_2353,In_2137);
nor U1843 (N_1843,In_1894,In_1923);
or U1844 (N_1844,In_2037,In_1558);
nand U1845 (N_1845,In_944,In_123);
or U1846 (N_1846,In_1028,In_861);
or U1847 (N_1847,In_1813,In_1554);
nor U1848 (N_1848,In_1171,In_1565);
nand U1849 (N_1849,In_416,In_744);
or U1850 (N_1850,In_215,In_1096);
nor U1851 (N_1851,In_1915,In_2106);
xnor U1852 (N_1852,In_1494,In_608);
or U1853 (N_1853,In_528,In_1518);
or U1854 (N_1854,In_2216,In_1255);
or U1855 (N_1855,In_2086,In_2293);
and U1856 (N_1856,In_871,In_840);
nor U1857 (N_1857,In_979,In_1654);
or U1858 (N_1858,In_2302,In_638);
nor U1859 (N_1859,In_2187,In_1050);
and U1860 (N_1860,In_1802,In_1273);
nor U1861 (N_1861,In_1718,In_980);
xnor U1862 (N_1862,In_1649,In_2043);
xor U1863 (N_1863,In_1132,In_428);
nand U1864 (N_1864,In_426,In_824);
or U1865 (N_1865,In_2199,In_103);
or U1866 (N_1866,In_980,In_1996);
nand U1867 (N_1867,In_2206,In_60);
or U1868 (N_1868,In_1622,In_783);
nor U1869 (N_1869,In_985,In_870);
and U1870 (N_1870,In_319,In_1457);
and U1871 (N_1871,In_703,In_1836);
nand U1872 (N_1872,In_2468,In_1591);
xor U1873 (N_1873,In_414,In_620);
nor U1874 (N_1874,In_1610,In_163);
nor U1875 (N_1875,In_1784,In_755);
nor U1876 (N_1876,In_895,In_961);
nand U1877 (N_1877,In_713,In_1789);
xnor U1878 (N_1878,In_964,In_108);
xnor U1879 (N_1879,In_1530,In_275);
xnor U1880 (N_1880,In_1393,In_947);
xor U1881 (N_1881,In_2016,In_2035);
nand U1882 (N_1882,In_2439,In_1826);
or U1883 (N_1883,In_2270,In_1540);
and U1884 (N_1884,In_1442,In_544);
or U1885 (N_1885,In_1418,In_1763);
and U1886 (N_1886,In_1916,In_823);
and U1887 (N_1887,In_2053,In_1467);
and U1888 (N_1888,In_358,In_332);
nand U1889 (N_1889,In_984,In_1047);
and U1890 (N_1890,In_2448,In_1272);
nor U1891 (N_1891,In_386,In_1335);
nand U1892 (N_1892,In_2341,In_469);
and U1893 (N_1893,In_1193,In_630);
and U1894 (N_1894,In_1819,In_1045);
xnor U1895 (N_1895,In_190,In_1359);
or U1896 (N_1896,In_472,In_1943);
or U1897 (N_1897,In_2054,In_1562);
and U1898 (N_1898,In_2172,In_432);
and U1899 (N_1899,In_819,In_30);
and U1900 (N_1900,In_1787,In_1910);
or U1901 (N_1901,In_2058,In_554);
and U1902 (N_1902,In_2365,In_1700);
and U1903 (N_1903,In_895,In_2000);
nor U1904 (N_1904,In_286,In_2025);
and U1905 (N_1905,In_405,In_967);
and U1906 (N_1906,In_878,In_656);
or U1907 (N_1907,In_2409,In_981);
xor U1908 (N_1908,In_48,In_1879);
or U1909 (N_1909,In_331,In_2200);
nor U1910 (N_1910,In_261,In_1440);
nand U1911 (N_1911,In_289,In_2208);
nor U1912 (N_1912,In_1530,In_4);
and U1913 (N_1913,In_1515,In_2293);
or U1914 (N_1914,In_209,In_1962);
nor U1915 (N_1915,In_1198,In_1709);
or U1916 (N_1916,In_948,In_576);
and U1917 (N_1917,In_2440,In_488);
nand U1918 (N_1918,In_1302,In_636);
nand U1919 (N_1919,In_4,In_1382);
or U1920 (N_1920,In_832,In_2013);
nand U1921 (N_1921,In_1101,In_2184);
or U1922 (N_1922,In_934,In_1350);
nor U1923 (N_1923,In_949,In_1099);
and U1924 (N_1924,In_942,In_210);
or U1925 (N_1925,In_1569,In_296);
xnor U1926 (N_1926,In_1483,In_2391);
or U1927 (N_1927,In_1860,In_180);
nor U1928 (N_1928,In_1451,In_712);
xnor U1929 (N_1929,In_977,In_2143);
nand U1930 (N_1930,In_1403,In_1799);
or U1931 (N_1931,In_986,In_1599);
nor U1932 (N_1932,In_762,In_2226);
xnor U1933 (N_1933,In_1199,In_113);
and U1934 (N_1934,In_1047,In_1584);
or U1935 (N_1935,In_16,In_1185);
or U1936 (N_1936,In_1528,In_1013);
or U1937 (N_1937,In_2223,In_1953);
nand U1938 (N_1938,In_1199,In_1128);
and U1939 (N_1939,In_661,In_1958);
nor U1940 (N_1940,In_121,In_970);
nor U1941 (N_1941,In_980,In_13);
xnor U1942 (N_1942,In_2289,In_572);
or U1943 (N_1943,In_1116,In_184);
or U1944 (N_1944,In_556,In_527);
or U1945 (N_1945,In_1344,In_79);
or U1946 (N_1946,In_2073,In_866);
and U1947 (N_1947,In_1587,In_1487);
xor U1948 (N_1948,In_2295,In_1807);
nor U1949 (N_1949,In_1921,In_1342);
and U1950 (N_1950,In_2421,In_254);
nand U1951 (N_1951,In_1626,In_115);
and U1952 (N_1952,In_1331,In_1323);
and U1953 (N_1953,In_1802,In_738);
xor U1954 (N_1954,In_1087,In_1088);
nand U1955 (N_1955,In_1928,In_1932);
nand U1956 (N_1956,In_1265,In_125);
nand U1957 (N_1957,In_655,In_2354);
and U1958 (N_1958,In_1491,In_617);
nor U1959 (N_1959,In_2412,In_974);
nand U1960 (N_1960,In_1859,In_1040);
nor U1961 (N_1961,In_173,In_1526);
xnor U1962 (N_1962,In_589,In_1805);
or U1963 (N_1963,In_968,In_2035);
nor U1964 (N_1964,In_2107,In_1718);
xnor U1965 (N_1965,In_1715,In_1840);
nand U1966 (N_1966,In_340,In_799);
or U1967 (N_1967,In_347,In_1125);
and U1968 (N_1968,In_1251,In_1362);
xnor U1969 (N_1969,In_1570,In_200);
or U1970 (N_1970,In_1012,In_1690);
xor U1971 (N_1971,In_1259,In_2147);
xor U1972 (N_1972,In_2294,In_868);
nor U1973 (N_1973,In_1057,In_1034);
xor U1974 (N_1974,In_791,In_624);
nand U1975 (N_1975,In_210,In_2251);
or U1976 (N_1976,In_1168,In_2478);
nand U1977 (N_1977,In_524,In_2373);
or U1978 (N_1978,In_1716,In_2480);
or U1979 (N_1979,In_475,In_1519);
nand U1980 (N_1980,In_26,In_1817);
or U1981 (N_1981,In_2012,In_1857);
or U1982 (N_1982,In_56,In_1066);
nand U1983 (N_1983,In_1047,In_2180);
nor U1984 (N_1984,In_531,In_2396);
xor U1985 (N_1985,In_70,In_1381);
nand U1986 (N_1986,In_127,In_1585);
or U1987 (N_1987,In_435,In_1523);
and U1988 (N_1988,In_2113,In_617);
or U1989 (N_1989,In_920,In_258);
nand U1990 (N_1990,In_2410,In_742);
nor U1991 (N_1991,In_965,In_1384);
nor U1992 (N_1992,In_2419,In_2478);
or U1993 (N_1993,In_2288,In_2074);
or U1994 (N_1994,In_766,In_1549);
nand U1995 (N_1995,In_1740,In_1457);
nand U1996 (N_1996,In_952,In_349);
nand U1997 (N_1997,In_1910,In_1683);
nor U1998 (N_1998,In_2273,In_264);
and U1999 (N_1999,In_510,In_108);
and U2000 (N_2000,In_2470,In_739);
nand U2001 (N_2001,In_1300,In_1325);
and U2002 (N_2002,In_999,In_1640);
nand U2003 (N_2003,In_1830,In_2067);
nand U2004 (N_2004,In_1794,In_440);
or U2005 (N_2005,In_1438,In_2490);
nand U2006 (N_2006,In_865,In_1497);
or U2007 (N_2007,In_1783,In_2056);
or U2008 (N_2008,In_114,In_475);
xor U2009 (N_2009,In_2261,In_2430);
nor U2010 (N_2010,In_457,In_2334);
and U2011 (N_2011,In_248,In_1912);
or U2012 (N_2012,In_291,In_925);
nand U2013 (N_2013,In_1451,In_1744);
and U2014 (N_2014,In_323,In_634);
and U2015 (N_2015,In_241,In_1363);
xor U2016 (N_2016,In_2059,In_202);
or U2017 (N_2017,In_1333,In_2285);
or U2018 (N_2018,In_1108,In_378);
nor U2019 (N_2019,In_1119,In_841);
nor U2020 (N_2020,In_2270,In_782);
nand U2021 (N_2021,In_625,In_996);
and U2022 (N_2022,In_1404,In_2456);
and U2023 (N_2023,In_661,In_221);
and U2024 (N_2024,In_1693,In_2404);
or U2025 (N_2025,In_1869,In_88);
nor U2026 (N_2026,In_2018,In_1531);
nor U2027 (N_2027,In_516,In_719);
nor U2028 (N_2028,In_1058,In_1580);
or U2029 (N_2029,In_557,In_1043);
nand U2030 (N_2030,In_1807,In_182);
and U2031 (N_2031,In_191,In_2207);
xor U2032 (N_2032,In_2085,In_528);
and U2033 (N_2033,In_2319,In_418);
nor U2034 (N_2034,In_2397,In_933);
xnor U2035 (N_2035,In_314,In_1775);
or U2036 (N_2036,In_1572,In_1533);
nor U2037 (N_2037,In_963,In_1429);
or U2038 (N_2038,In_1810,In_506);
nor U2039 (N_2039,In_624,In_2210);
nand U2040 (N_2040,In_327,In_147);
or U2041 (N_2041,In_138,In_2263);
and U2042 (N_2042,In_48,In_1866);
and U2043 (N_2043,In_1040,In_1403);
nor U2044 (N_2044,In_29,In_1229);
and U2045 (N_2045,In_1950,In_48);
xor U2046 (N_2046,In_1987,In_944);
nand U2047 (N_2047,In_173,In_1059);
nor U2048 (N_2048,In_1211,In_2398);
xor U2049 (N_2049,In_654,In_1549);
nor U2050 (N_2050,In_1684,In_2156);
or U2051 (N_2051,In_39,In_420);
and U2052 (N_2052,In_660,In_871);
xnor U2053 (N_2053,In_1841,In_1036);
and U2054 (N_2054,In_2391,In_1214);
nand U2055 (N_2055,In_1902,In_855);
nand U2056 (N_2056,In_2392,In_1466);
nor U2057 (N_2057,In_69,In_1488);
or U2058 (N_2058,In_1648,In_428);
nor U2059 (N_2059,In_1450,In_1927);
and U2060 (N_2060,In_532,In_663);
or U2061 (N_2061,In_367,In_2325);
and U2062 (N_2062,In_2425,In_1575);
nand U2063 (N_2063,In_2354,In_1399);
or U2064 (N_2064,In_753,In_998);
nand U2065 (N_2065,In_378,In_2491);
nand U2066 (N_2066,In_923,In_2331);
and U2067 (N_2067,In_165,In_1831);
and U2068 (N_2068,In_1208,In_969);
or U2069 (N_2069,In_2143,In_676);
nor U2070 (N_2070,In_224,In_1939);
or U2071 (N_2071,In_1298,In_2222);
xor U2072 (N_2072,In_682,In_782);
and U2073 (N_2073,In_1386,In_18);
nand U2074 (N_2074,In_1059,In_2205);
nand U2075 (N_2075,In_414,In_2081);
nand U2076 (N_2076,In_1088,In_57);
nor U2077 (N_2077,In_881,In_635);
or U2078 (N_2078,In_1325,In_1516);
nand U2079 (N_2079,In_1621,In_547);
xor U2080 (N_2080,In_578,In_1909);
or U2081 (N_2081,In_1116,In_466);
or U2082 (N_2082,In_799,In_72);
nor U2083 (N_2083,In_1489,In_807);
nand U2084 (N_2084,In_12,In_2010);
and U2085 (N_2085,In_1139,In_2010);
nor U2086 (N_2086,In_2174,In_169);
nand U2087 (N_2087,In_418,In_1913);
nor U2088 (N_2088,In_1775,In_2238);
nor U2089 (N_2089,In_1085,In_959);
and U2090 (N_2090,In_1474,In_2434);
and U2091 (N_2091,In_618,In_1672);
xnor U2092 (N_2092,In_712,In_1879);
and U2093 (N_2093,In_1907,In_919);
and U2094 (N_2094,In_446,In_762);
nand U2095 (N_2095,In_1081,In_569);
xnor U2096 (N_2096,In_1376,In_1401);
xnor U2097 (N_2097,In_539,In_1012);
and U2098 (N_2098,In_1590,In_1444);
nand U2099 (N_2099,In_501,In_1370);
or U2100 (N_2100,In_2275,In_1736);
and U2101 (N_2101,In_1452,In_1496);
and U2102 (N_2102,In_735,In_2344);
nand U2103 (N_2103,In_532,In_1230);
nor U2104 (N_2104,In_426,In_1887);
or U2105 (N_2105,In_1421,In_1598);
or U2106 (N_2106,In_1319,In_1909);
nor U2107 (N_2107,In_1432,In_2413);
nor U2108 (N_2108,In_980,In_2195);
and U2109 (N_2109,In_1561,In_676);
or U2110 (N_2110,In_994,In_1001);
or U2111 (N_2111,In_1,In_334);
or U2112 (N_2112,In_173,In_671);
or U2113 (N_2113,In_1104,In_864);
nor U2114 (N_2114,In_1023,In_3);
or U2115 (N_2115,In_1820,In_2238);
and U2116 (N_2116,In_989,In_588);
nand U2117 (N_2117,In_367,In_2432);
or U2118 (N_2118,In_1511,In_588);
or U2119 (N_2119,In_2132,In_2332);
nor U2120 (N_2120,In_1993,In_58);
xor U2121 (N_2121,In_1540,In_1943);
nand U2122 (N_2122,In_1089,In_69);
nand U2123 (N_2123,In_399,In_112);
nand U2124 (N_2124,In_1547,In_2410);
or U2125 (N_2125,In_1220,In_2285);
nor U2126 (N_2126,In_97,In_1271);
nor U2127 (N_2127,In_1531,In_196);
nor U2128 (N_2128,In_1357,In_818);
or U2129 (N_2129,In_1417,In_2032);
or U2130 (N_2130,In_1084,In_1388);
nand U2131 (N_2131,In_834,In_1081);
and U2132 (N_2132,In_2224,In_1260);
nor U2133 (N_2133,In_1924,In_1778);
or U2134 (N_2134,In_1125,In_1101);
or U2135 (N_2135,In_572,In_529);
xnor U2136 (N_2136,In_2350,In_740);
or U2137 (N_2137,In_382,In_2291);
nor U2138 (N_2138,In_1842,In_1882);
and U2139 (N_2139,In_657,In_2485);
or U2140 (N_2140,In_1476,In_2273);
or U2141 (N_2141,In_1863,In_2342);
nor U2142 (N_2142,In_1754,In_1707);
and U2143 (N_2143,In_2202,In_800);
nor U2144 (N_2144,In_421,In_883);
or U2145 (N_2145,In_1894,In_2364);
and U2146 (N_2146,In_2301,In_1980);
nand U2147 (N_2147,In_2468,In_844);
or U2148 (N_2148,In_953,In_53);
nand U2149 (N_2149,In_1566,In_1008);
and U2150 (N_2150,In_184,In_804);
or U2151 (N_2151,In_383,In_1929);
nand U2152 (N_2152,In_152,In_549);
xnor U2153 (N_2153,In_1862,In_1444);
nand U2154 (N_2154,In_433,In_1248);
nor U2155 (N_2155,In_1921,In_1134);
and U2156 (N_2156,In_134,In_1558);
and U2157 (N_2157,In_770,In_1297);
and U2158 (N_2158,In_1372,In_918);
nand U2159 (N_2159,In_419,In_2447);
or U2160 (N_2160,In_1850,In_2484);
nor U2161 (N_2161,In_551,In_1589);
or U2162 (N_2162,In_1996,In_912);
xnor U2163 (N_2163,In_1873,In_1584);
and U2164 (N_2164,In_1719,In_973);
nor U2165 (N_2165,In_346,In_1906);
or U2166 (N_2166,In_2451,In_189);
nand U2167 (N_2167,In_181,In_72);
nor U2168 (N_2168,In_672,In_755);
or U2169 (N_2169,In_1387,In_2254);
nand U2170 (N_2170,In_1684,In_170);
nor U2171 (N_2171,In_739,In_215);
and U2172 (N_2172,In_1501,In_280);
xor U2173 (N_2173,In_185,In_1665);
nor U2174 (N_2174,In_1037,In_1102);
nand U2175 (N_2175,In_1964,In_1908);
and U2176 (N_2176,In_2496,In_1949);
or U2177 (N_2177,In_1695,In_2048);
and U2178 (N_2178,In_1960,In_253);
nor U2179 (N_2179,In_2430,In_214);
nor U2180 (N_2180,In_1382,In_749);
nor U2181 (N_2181,In_2016,In_867);
or U2182 (N_2182,In_846,In_756);
xor U2183 (N_2183,In_2283,In_1238);
nor U2184 (N_2184,In_1238,In_1499);
or U2185 (N_2185,In_1368,In_1177);
nand U2186 (N_2186,In_561,In_470);
and U2187 (N_2187,In_1127,In_2164);
or U2188 (N_2188,In_1245,In_138);
and U2189 (N_2189,In_1336,In_138);
and U2190 (N_2190,In_1560,In_1765);
nand U2191 (N_2191,In_131,In_2463);
or U2192 (N_2192,In_1295,In_558);
nor U2193 (N_2193,In_197,In_1522);
or U2194 (N_2194,In_412,In_997);
and U2195 (N_2195,In_715,In_2264);
nand U2196 (N_2196,In_663,In_1520);
nand U2197 (N_2197,In_2057,In_686);
xor U2198 (N_2198,In_2098,In_2204);
nor U2199 (N_2199,In_2288,In_489);
nor U2200 (N_2200,In_1994,In_1354);
or U2201 (N_2201,In_2316,In_2417);
nand U2202 (N_2202,In_723,In_1987);
xnor U2203 (N_2203,In_205,In_2245);
and U2204 (N_2204,In_2452,In_153);
nor U2205 (N_2205,In_2042,In_329);
and U2206 (N_2206,In_331,In_554);
or U2207 (N_2207,In_18,In_2316);
or U2208 (N_2208,In_77,In_1200);
or U2209 (N_2209,In_1268,In_1685);
nand U2210 (N_2210,In_2257,In_1244);
and U2211 (N_2211,In_1787,In_2435);
nand U2212 (N_2212,In_1191,In_2273);
or U2213 (N_2213,In_912,In_264);
and U2214 (N_2214,In_1301,In_1183);
nand U2215 (N_2215,In_2419,In_1969);
nor U2216 (N_2216,In_1999,In_1686);
or U2217 (N_2217,In_631,In_2343);
or U2218 (N_2218,In_2348,In_1237);
and U2219 (N_2219,In_807,In_2301);
nor U2220 (N_2220,In_1923,In_1420);
or U2221 (N_2221,In_168,In_938);
nor U2222 (N_2222,In_844,In_1008);
or U2223 (N_2223,In_1889,In_228);
and U2224 (N_2224,In_1922,In_1118);
nand U2225 (N_2225,In_1690,In_2499);
nand U2226 (N_2226,In_1576,In_958);
and U2227 (N_2227,In_1613,In_1635);
and U2228 (N_2228,In_977,In_2465);
or U2229 (N_2229,In_2098,In_1725);
nor U2230 (N_2230,In_999,In_137);
nand U2231 (N_2231,In_1050,In_2404);
or U2232 (N_2232,In_2092,In_2436);
and U2233 (N_2233,In_1501,In_128);
or U2234 (N_2234,In_1945,In_1223);
or U2235 (N_2235,In_1187,In_117);
nor U2236 (N_2236,In_1412,In_590);
nor U2237 (N_2237,In_1102,In_1752);
nand U2238 (N_2238,In_1481,In_477);
nor U2239 (N_2239,In_382,In_828);
nand U2240 (N_2240,In_1773,In_1230);
and U2241 (N_2241,In_2234,In_2073);
and U2242 (N_2242,In_438,In_1024);
or U2243 (N_2243,In_371,In_1550);
or U2244 (N_2244,In_1927,In_968);
or U2245 (N_2245,In_2199,In_1569);
and U2246 (N_2246,In_1092,In_2057);
and U2247 (N_2247,In_162,In_31);
and U2248 (N_2248,In_2398,In_2206);
xor U2249 (N_2249,In_2244,In_136);
nor U2250 (N_2250,In_2015,In_64);
or U2251 (N_2251,In_255,In_1408);
or U2252 (N_2252,In_1254,In_904);
and U2253 (N_2253,In_1425,In_723);
or U2254 (N_2254,In_609,In_1939);
xnor U2255 (N_2255,In_806,In_1941);
nand U2256 (N_2256,In_2437,In_75);
nor U2257 (N_2257,In_314,In_246);
nor U2258 (N_2258,In_1089,In_2194);
or U2259 (N_2259,In_1083,In_113);
and U2260 (N_2260,In_998,In_2440);
and U2261 (N_2261,In_1431,In_953);
nor U2262 (N_2262,In_1739,In_1406);
and U2263 (N_2263,In_293,In_2076);
xnor U2264 (N_2264,In_1606,In_1842);
nor U2265 (N_2265,In_1830,In_850);
nand U2266 (N_2266,In_576,In_2006);
and U2267 (N_2267,In_2483,In_727);
xor U2268 (N_2268,In_96,In_2095);
or U2269 (N_2269,In_751,In_1858);
xor U2270 (N_2270,In_528,In_1830);
nor U2271 (N_2271,In_142,In_997);
nand U2272 (N_2272,In_1864,In_838);
nand U2273 (N_2273,In_188,In_48);
xor U2274 (N_2274,In_688,In_201);
and U2275 (N_2275,In_1508,In_1639);
or U2276 (N_2276,In_588,In_640);
or U2277 (N_2277,In_2131,In_2494);
nor U2278 (N_2278,In_402,In_835);
nand U2279 (N_2279,In_1116,In_2114);
and U2280 (N_2280,In_304,In_2136);
nor U2281 (N_2281,In_550,In_2262);
and U2282 (N_2282,In_1601,In_269);
or U2283 (N_2283,In_936,In_2047);
and U2284 (N_2284,In_1141,In_1855);
or U2285 (N_2285,In_1649,In_482);
nand U2286 (N_2286,In_387,In_1407);
nand U2287 (N_2287,In_1698,In_705);
or U2288 (N_2288,In_364,In_448);
and U2289 (N_2289,In_278,In_173);
and U2290 (N_2290,In_165,In_2379);
and U2291 (N_2291,In_2333,In_698);
nand U2292 (N_2292,In_876,In_2305);
or U2293 (N_2293,In_1740,In_991);
nand U2294 (N_2294,In_2043,In_1827);
nor U2295 (N_2295,In_2194,In_979);
or U2296 (N_2296,In_2004,In_854);
nand U2297 (N_2297,In_1862,In_1575);
xnor U2298 (N_2298,In_677,In_1974);
and U2299 (N_2299,In_1536,In_717);
and U2300 (N_2300,In_263,In_1028);
nor U2301 (N_2301,In_949,In_496);
or U2302 (N_2302,In_1019,In_1085);
nor U2303 (N_2303,In_1960,In_2333);
or U2304 (N_2304,In_399,In_1203);
or U2305 (N_2305,In_201,In_34);
or U2306 (N_2306,In_2293,In_803);
nand U2307 (N_2307,In_228,In_2439);
nor U2308 (N_2308,In_452,In_1151);
nand U2309 (N_2309,In_466,In_310);
nor U2310 (N_2310,In_1306,In_2458);
and U2311 (N_2311,In_2185,In_1025);
and U2312 (N_2312,In_548,In_1817);
nor U2313 (N_2313,In_1306,In_1945);
or U2314 (N_2314,In_1401,In_2088);
or U2315 (N_2315,In_190,In_1856);
xnor U2316 (N_2316,In_632,In_1648);
or U2317 (N_2317,In_1494,In_2043);
and U2318 (N_2318,In_2475,In_794);
and U2319 (N_2319,In_2388,In_1357);
or U2320 (N_2320,In_1028,In_345);
or U2321 (N_2321,In_1901,In_2454);
nor U2322 (N_2322,In_1897,In_1501);
nor U2323 (N_2323,In_794,In_157);
nand U2324 (N_2324,In_693,In_1519);
or U2325 (N_2325,In_133,In_233);
nand U2326 (N_2326,In_936,In_2412);
and U2327 (N_2327,In_911,In_1260);
or U2328 (N_2328,In_1152,In_1731);
xor U2329 (N_2329,In_8,In_318);
nor U2330 (N_2330,In_2230,In_1585);
nand U2331 (N_2331,In_66,In_2421);
and U2332 (N_2332,In_2384,In_940);
or U2333 (N_2333,In_1732,In_2094);
nor U2334 (N_2334,In_595,In_2091);
or U2335 (N_2335,In_2129,In_2178);
or U2336 (N_2336,In_1833,In_116);
and U2337 (N_2337,In_44,In_2205);
nand U2338 (N_2338,In_2075,In_1045);
and U2339 (N_2339,In_1549,In_2450);
nand U2340 (N_2340,In_1435,In_1042);
or U2341 (N_2341,In_2393,In_914);
nor U2342 (N_2342,In_1743,In_140);
or U2343 (N_2343,In_401,In_2445);
nor U2344 (N_2344,In_688,In_2048);
xnor U2345 (N_2345,In_1294,In_1558);
nand U2346 (N_2346,In_1867,In_356);
or U2347 (N_2347,In_1293,In_1748);
xnor U2348 (N_2348,In_2244,In_1900);
xor U2349 (N_2349,In_378,In_1145);
or U2350 (N_2350,In_297,In_2047);
or U2351 (N_2351,In_2096,In_1884);
and U2352 (N_2352,In_1000,In_1371);
xor U2353 (N_2353,In_2344,In_1776);
nand U2354 (N_2354,In_1284,In_2217);
and U2355 (N_2355,In_580,In_1678);
nor U2356 (N_2356,In_1025,In_1650);
and U2357 (N_2357,In_2082,In_1053);
nand U2358 (N_2358,In_1481,In_2126);
nand U2359 (N_2359,In_894,In_1127);
and U2360 (N_2360,In_122,In_215);
and U2361 (N_2361,In_1777,In_1957);
nand U2362 (N_2362,In_2177,In_1577);
and U2363 (N_2363,In_166,In_478);
or U2364 (N_2364,In_158,In_2030);
nor U2365 (N_2365,In_1892,In_574);
xor U2366 (N_2366,In_271,In_1175);
xor U2367 (N_2367,In_1711,In_396);
nand U2368 (N_2368,In_2375,In_1521);
and U2369 (N_2369,In_1516,In_1915);
nand U2370 (N_2370,In_1443,In_1057);
and U2371 (N_2371,In_2122,In_2035);
nor U2372 (N_2372,In_1360,In_1439);
nor U2373 (N_2373,In_1192,In_797);
and U2374 (N_2374,In_1772,In_2352);
nand U2375 (N_2375,In_2296,In_2079);
xnor U2376 (N_2376,In_1073,In_420);
and U2377 (N_2377,In_2331,In_564);
and U2378 (N_2378,In_735,In_2273);
or U2379 (N_2379,In_643,In_1569);
and U2380 (N_2380,In_1185,In_1777);
and U2381 (N_2381,In_452,In_1606);
nor U2382 (N_2382,In_253,In_1152);
or U2383 (N_2383,In_215,In_1993);
nor U2384 (N_2384,In_1973,In_442);
and U2385 (N_2385,In_1947,In_68);
and U2386 (N_2386,In_113,In_954);
xor U2387 (N_2387,In_268,In_1132);
and U2388 (N_2388,In_1830,In_1350);
and U2389 (N_2389,In_1474,In_2211);
nor U2390 (N_2390,In_1864,In_388);
or U2391 (N_2391,In_2295,In_498);
nand U2392 (N_2392,In_1602,In_346);
or U2393 (N_2393,In_1001,In_2346);
nor U2394 (N_2394,In_1406,In_2213);
nand U2395 (N_2395,In_1486,In_880);
and U2396 (N_2396,In_928,In_735);
or U2397 (N_2397,In_2442,In_34);
nand U2398 (N_2398,In_183,In_714);
or U2399 (N_2399,In_423,In_2028);
xor U2400 (N_2400,In_1719,In_2016);
nand U2401 (N_2401,In_1012,In_791);
or U2402 (N_2402,In_291,In_335);
or U2403 (N_2403,In_1191,In_2379);
nand U2404 (N_2404,In_1179,In_2357);
and U2405 (N_2405,In_606,In_2379);
or U2406 (N_2406,In_507,In_689);
nand U2407 (N_2407,In_484,In_938);
nor U2408 (N_2408,In_5,In_1667);
xnor U2409 (N_2409,In_2162,In_1273);
and U2410 (N_2410,In_1283,In_1658);
xor U2411 (N_2411,In_1158,In_1495);
and U2412 (N_2412,In_2291,In_1742);
nor U2413 (N_2413,In_1855,In_2172);
nand U2414 (N_2414,In_2390,In_674);
and U2415 (N_2415,In_1201,In_766);
or U2416 (N_2416,In_97,In_1441);
and U2417 (N_2417,In_249,In_1887);
and U2418 (N_2418,In_2453,In_1886);
or U2419 (N_2419,In_2090,In_390);
or U2420 (N_2420,In_1717,In_1442);
nand U2421 (N_2421,In_2276,In_616);
or U2422 (N_2422,In_1097,In_1616);
xnor U2423 (N_2423,In_1055,In_192);
nand U2424 (N_2424,In_662,In_1991);
xnor U2425 (N_2425,In_154,In_1172);
and U2426 (N_2426,In_1284,In_443);
nand U2427 (N_2427,In_445,In_2059);
nand U2428 (N_2428,In_2295,In_510);
and U2429 (N_2429,In_2056,In_1396);
nand U2430 (N_2430,In_1530,In_273);
xor U2431 (N_2431,In_1176,In_279);
nor U2432 (N_2432,In_52,In_1133);
nor U2433 (N_2433,In_489,In_976);
and U2434 (N_2434,In_1900,In_957);
nor U2435 (N_2435,In_1770,In_1874);
and U2436 (N_2436,In_634,In_1491);
xor U2437 (N_2437,In_1876,In_8);
xnor U2438 (N_2438,In_2197,In_503);
nand U2439 (N_2439,In_228,In_2082);
and U2440 (N_2440,In_2439,In_680);
nor U2441 (N_2441,In_2413,In_743);
nor U2442 (N_2442,In_660,In_189);
and U2443 (N_2443,In_95,In_812);
nor U2444 (N_2444,In_1342,In_2195);
nand U2445 (N_2445,In_59,In_581);
and U2446 (N_2446,In_2485,In_1526);
nor U2447 (N_2447,In_2080,In_509);
or U2448 (N_2448,In_436,In_2199);
nand U2449 (N_2449,In_571,In_490);
nor U2450 (N_2450,In_1976,In_31);
and U2451 (N_2451,In_2201,In_523);
nor U2452 (N_2452,In_1683,In_461);
nor U2453 (N_2453,In_59,In_1659);
nand U2454 (N_2454,In_768,In_1946);
nor U2455 (N_2455,In_1925,In_1895);
and U2456 (N_2456,In_2450,In_175);
nand U2457 (N_2457,In_1624,In_1190);
nand U2458 (N_2458,In_1042,In_151);
or U2459 (N_2459,In_394,In_1542);
and U2460 (N_2460,In_923,In_1716);
nand U2461 (N_2461,In_1237,In_1720);
nor U2462 (N_2462,In_478,In_1646);
or U2463 (N_2463,In_1337,In_1415);
nand U2464 (N_2464,In_2262,In_1975);
nor U2465 (N_2465,In_384,In_1540);
or U2466 (N_2466,In_2308,In_128);
and U2467 (N_2467,In_1418,In_1841);
and U2468 (N_2468,In_1643,In_1701);
and U2469 (N_2469,In_442,In_2210);
and U2470 (N_2470,In_1282,In_61);
nor U2471 (N_2471,In_2165,In_1560);
nand U2472 (N_2472,In_2066,In_1158);
or U2473 (N_2473,In_1530,In_620);
and U2474 (N_2474,In_1130,In_620);
and U2475 (N_2475,In_2091,In_362);
xnor U2476 (N_2476,In_2494,In_2072);
or U2477 (N_2477,In_2302,In_1917);
nor U2478 (N_2478,In_111,In_2267);
nor U2479 (N_2479,In_1655,In_1396);
and U2480 (N_2480,In_1565,In_91);
or U2481 (N_2481,In_1304,In_814);
xor U2482 (N_2482,In_1452,In_2081);
nor U2483 (N_2483,In_2413,In_499);
or U2484 (N_2484,In_1989,In_1532);
nor U2485 (N_2485,In_1913,In_1089);
nor U2486 (N_2486,In_940,In_2215);
or U2487 (N_2487,In_1058,In_914);
or U2488 (N_2488,In_1430,In_531);
or U2489 (N_2489,In_1990,In_1913);
and U2490 (N_2490,In_1176,In_1117);
xor U2491 (N_2491,In_837,In_1094);
nand U2492 (N_2492,In_2098,In_1803);
nand U2493 (N_2493,In_1656,In_812);
and U2494 (N_2494,In_807,In_465);
xor U2495 (N_2495,In_1812,In_1861);
and U2496 (N_2496,In_1867,In_273);
nand U2497 (N_2497,In_152,In_2269);
nand U2498 (N_2498,In_1773,In_1440);
or U2499 (N_2499,In_1096,In_2160);
and U2500 (N_2500,In_1598,In_1794);
nand U2501 (N_2501,In_516,In_1279);
and U2502 (N_2502,In_2244,In_2323);
xor U2503 (N_2503,In_827,In_20);
nand U2504 (N_2504,In_1436,In_1086);
and U2505 (N_2505,In_1804,In_1462);
and U2506 (N_2506,In_2377,In_274);
and U2507 (N_2507,In_1978,In_2026);
or U2508 (N_2508,In_468,In_1752);
nand U2509 (N_2509,In_894,In_1445);
nor U2510 (N_2510,In_329,In_968);
nor U2511 (N_2511,In_1734,In_1008);
nor U2512 (N_2512,In_2083,In_1536);
nand U2513 (N_2513,In_2073,In_1530);
nor U2514 (N_2514,In_354,In_944);
nand U2515 (N_2515,In_615,In_774);
nand U2516 (N_2516,In_837,In_1861);
and U2517 (N_2517,In_1089,In_782);
nor U2518 (N_2518,In_744,In_1932);
and U2519 (N_2519,In_2341,In_1441);
or U2520 (N_2520,In_1626,In_2047);
nor U2521 (N_2521,In_204,In_118);
and U2522 (N_2522,In_1661,In_2070);
xor U2523 (N_2523,In_827,In_1080);
and U2524 (N_2524,In_1447,In_1615);
and U2525 (N_2525,In_174,In_1172);
and U2526 (N_2526,In_2270,In_1360);
or U2527 (N_2527,In_460,In_1149);
and U2528 (N_2528,In_1815,In_798);
nand U2529 (N_2529,In_267,In_186);
nand U2530 (N_2530,In_1604,In_2179);
xor U2531 (N_2531,In_608,In_2353);
or U2532 (N_2532,In_224,In_2401);
nor U2533 (N_2533,In_815,In_443);
nand U2534 (N_2534,In_1159,In_2317);
nand U2535 (N_2535,In_1343,In_1729);
and U2536 (N_2536,In_954,In_97);
nor U2537 (N_2537,In_1067,In_722);
nor U2538 (N_2538,In_1732,In_741);
or U2539 (N_2539,In_1510,In_2455);
and U2540 (N_2540,In_1508,In_2131);
or U2541 (N_2541,In_1322,In_579);
xor U2542 (N_2542,In_1779,In_2208);
and U2543 (N_2543,In_1520,In_1800);
and U2544 (N_2544,In_2350,In_1511);
or U2545 (N_2545,In_21,In_1108);
nand U2546 (N_2546,In_1975,In_834);
xor U2547 (N_2547,In_1031,In_269);
and U2548 (N_2548,In_2058,In_1788);
or U2549 (N_2549,In_1771,In_1816);
or U2550 (N_2550,In_1855,In_1991);
nand U2551 (N_2551,In_1722,In_60);
nor U2552 (N_2552,In_2380,In_1238);
and U2553 (N_2553,In_2491,In_1362);
nand U2554 (N_2554,In_944,In_1213);
or U2555 (N_2555,In_1849,In_136);
xnor U2556 (N_2556,In_1003,In_381);
and U2557 (N_2557,In_2325,In_408);
and U2558 (N_2558,In_2482,In_1107);
nand U2559 (N_2559,In_2205,In_1119);
nor U2560 (N_2560,In_2191,In_1296);
xnor U2561 (N_2561,In_76,In_898);
or U2562 (N_2562,In_1735,In_1561);
nand U2563 (N_2563,In_1897,In_1552);
and U2564 (N_2564,In_359,In_1632);
and U2565 (N_2565,In_1712,In_2013);
xor U2566 (N_2566,In_458,In_1284);
nand U2567 (N_2567,In_1212,In_1606);
and U2568 (N_2568,In_778,In_2450);
xor U2569 (N_2569,In_1161,In_1215);
nand U2570 (N_2570,In_1478,In_1091);
and U2571 (N_2571,In_2010,In_536);
and U2572 (N_2572,In_927,In_2114);
xor U2573 (N_2573,In_1443,In_169);
or U2574 (N_2574,In_1240,In_2167);
and U2575 (N_2575,In_1611,In_2478);
or U2576 (N_2576,In_2449,In_1060);
or U2577 (N_2577,In_2155,In_2400);
nor U2578 (N_2578,In_166,In_2453);
and U2579 (N_2579,In_1392,In_1068);
nor U2580 (N_2580,In_2157,In_1597);
and U2581 (N_2581,In_1944,In_1754);
or U2582 (N_2582,In_1729,In_889);
and U2583 (N_2583,In_2018,In_1847);
nand U2584 (N_2584,In_1584,In_609);
nor U2585 (N_2585,In_788,In_2053);
or U2586 (N_2586,In_24,In_545);
or U2587 (N_2587,In_2187,In_1438);
nor U2588 (N_2588,In_778,In_1240);
and U2589 (N_2589,In_1979,In_1202);
or U2590 (N_2590,In_343,In_2293);
xor U2591 (N_2591,In_182,In_449);
and U2592 (N_2592,In_2446,In_1034);
and U2593 (N_2593,In_981,In_2252);
or U2594 (N_2594,In_799,In_670);
nand U2595 (N_2595,In_341,In_272);
xnor U2596 (N_2596,In_663,In_148);
nand U2597 (N_2597,In_1342,In_2231);
nand U2598 (N_2598,In_1280,In_2042);
xnor U2599 (N_2599,In_640,In_1685);
nand U2600 (N_2600,In_837,In_289);
nor U2601 (N_2601,In_506,In_572);
and U2602 (N_2602,In_1649,In_1693);
and U2603 (N_2603,In_2328,In_788);
nor U2604 (N_2604,In_1432,In_1064);
or U2605 (N_2605,In_2472,In_140);
nand U2606 (N_2606,In_948,In_1814);
or U2607 (N_2607,In_924,In_1428);
or U2608 (N_2608,In_1667,In_1548);
nor U2609 (N_2609,In_659,In_1946);
nand U2610 (N_2610,In_2102,In_370);
or U2611 (N_2611,In_457,In_701);
and U2612 (N_2612,In_902,In_764);
xor U2613 (N_2613,In_709,In_617);
and U2614 (N_2614,In_1281,In_1089);
nand U2615 (N_2615,In_2430,In_2170);
nor U2616 (N_2616,In_498,In_354);
nand U2617 (N_2617,In_1383,In_2439);
nor U2618 (N_2618,In_522,In_368);
nand U2619 (N_2619,In_452,In_694);
or U2620 (N_2620,In_2235,In_2260);
or U2621 (N_2621,In_2161,In_2376);
nor U2622 (N_2622,In_787,In_1322);
nand U2623 (N_2623,In_198,In_1918);
nor U2624 (N_2624,In_2322,In_2297);
xnor U2625 (N_2625,In_2066,In_186);
nor U2626 (N_2626,In_1846,In_905);
or U2627 (N_2627,In_2211,In_2288);
nor U2628 (N_2628,In_1269,In_1542);
nand U2629 (N_2629,In_372,In_560);
nand U2630 (N_2630,In_930,In_1549);
nand U2631 (N_2631,In_656,In_407);
and U2632 (N_2632,In_2119,In_1935);
or U2633 (N_2633,In_893,In_1913);
and U2634 (N_2634,In_512,In_1461);
or U2635 (N_2635,In_2081,In_1782);
nand U2636 (N_2636,In_2034,In_1819);
nor U2637 (N_2637,In_1904,In_1860);
nor U2638 (N_2638,In_1985,In_1458);
nand U2639 (N_2639,In_1754,In_2014);
or U2640 (N_2640,In_2164,In_1078);
and U2641 (N_2641,In_494,In_1786);
or U2642 (N_2642,In_373,In_1815);
and U2643 (N_2643,In_1751,In_1328);
or U2644 (N_2644,In_30,In_470);
nor U2645 (N_2645,In_1594,In_720);
nand U2646 (N_2646,In_2442,In_445);
nor U2647 (N_2647,In_2437,In_1015);
nor U2648 (N_2648,In_749,In_300);
nand U2649 (N_2649,In_94,In_242);
and U2650 (N_2650,In_756,In_1695);
nand U2651 (N_2651,In_2348,In_664);
and U2652 (N_2652,In_1297,In_2316);
xnor U2653 (N_2653,In_95,In_1185);
or U2654 (N_2654,In_888,In_2174);
or U2655 (N_2655,In_2458,In_1893);
or U2656 (N_2656,In_1222,In_61);
nor U2657 (N_2657,In_319,In_1674);
nor U2658 (N_2658,In_1755,In_2309);
nand U2659 (N_2659,In_2069,In_1735);
and U2660 (N_2660,In_389,In_446);
or U2661 (N_2661,In_1590,In_1588);
nor U2662 (N_2662,In_45,In_2081);
nor U2663 (N_2663,In_1070,In_1950);
nor U2664 (N_2664,In_2030,In_362);
xor U2665 (N_2665,In_1519,In_384);
and U2666 (N_2666,In_1964,In_846);
or U2667 (N_2667,In_160,In_95);
nand U2668 (N_2668,In_574,In_999);
nor U2669 (N_2669,In_2360,In_1524);
nand U2670 (N_2670,In_422,In_279);
or U2671 (N_2671,In_1316,In_1430);
nand U2672 (N_2672,In_1935,In_1707);
nor U2673 (N_2673,In_2150,In_107);
or U2674 (N_2674,In_1810,In_1688);
or U2675 (N_2675,In_752,In_1180);
nand U2676 (N_2676,In_426,In_2193);
or U2677 (N_2677,In_45,In_769);
nand U2678 (N_2678,In_766,In_1464);
xor U2679 (N_2679,In_2044,In_1880);
xor U2680 (N_2680,In_203,In_795);
or U2681 (N_2681,In_651,In_1363);
nor U2682 (N_2682,In_1955,In_201);
or U2683 (N_2683,In_248,In_1260);
or U2684 (N_2684,In_696,In_1896);
and U2685 (N_2685,In_481,In_2360);
or U2686 (N_2686,In_1608,In_615);
and U2687 (N_2687,In_2300,In_774);
nor U2688 (N_2688,In_2318,In_2144);
and U2689 (N_2689,In_884,In_1495);
nand U2690 (N_2690,In_1759,In_256);
and U2691 (N_2691,In_2235,In_293);
xor U2692 (N_2692,In_1154,In_2245);
nor U2693 (N_2693,In_1600,In_1465);
or U2694 (N_2694,In_1615,In_920);
and U2695 (N_2695,In_638,In_74);
nor U2696 (N_2696,In_693,In_1817);
or U2697 (N_2697,In_2076,In_1046);
nor U2698 (N_2698,In_2087,In_1057);
xnor U2699 (N_2699,In_1832,In_22);
or U2700 (N_2700,In_185,In_2032);
or U2701 (N_2701,In_888,In_498);
nand U2702 (N_2702,In_1268,In_1868);
and U2703 (N_2703,In_418,In_164);
and U2704 (N_2704,In_1897,In_754);
nor U2705 (N_2705,In_847,In_1401);
or U2706 (N_2706,In_1251,In_1454);
nor U2707 (N_2707,In_1327,In_12);
and U2708 (N_2708,In_570,In_164);
or U2709 (N_2709,In_1132,In_501);
or U2710 (N_2710,In_878,In_1935);
xnor U2711 (N_2711,In_2147,In_2292);
and U2712 (N_2712,In_1629,In_2167);
or U2713 (N_2713,In_327,In_2312);
nor U2714 (N_2714,In_1959,In_1761);
nor U2715 (N_2715,In_1102,In_1542);
nand U2716 (N_2716,In_906,In_168);
nor U2717 (N_2717,In_138,In_2374);
and U2718 (N_2718,In_2255,In_24);
xnor U2719 (N_2719,In_286,In_520);
nor U2720 (N_2720,In_552,In_1512);
or U2721 (N_2721,In_1102,In_1835);
or U2722 (N_2722,In_1463,In_170);
or U2723 (N_2723,In_562,In_1241);
or U2724 (N_2724,In_813,In_752);
nand U2725 (N_2725,In_1496,In_2355);
and U2726 (N_2726,In_666,In_791);
xnor U2727 (N_2727,In_1851,In_2271);
or U2728 (N_2728,In_321,In_2047);
or U2729 (N_2729,In_995,In_27);
nand U2730 (N_2730,In_1285,In_11);
nor U2731 (N_2731,In_2394,In_2461);
nand U2732 (N_2732,In_1614,In_1922);
nand U2733 (N_2733,In_1980,In_1164);
xnor U2734 (N_2734,In_1144,In_1052);
nand U2735 (N_2735,In_228,In_2206);
and U2736 (N_2736,In_1824,In_485);
nand U2737 (N_2737,In_2466,In_2005);
nand U2738 (N_2738,In_181,In_1424);
or U2739 (N_2739,In_2381,In_819);
nand U2740 (N_2740,In_1289,In_2265);
nand U2741 (N_2741,In_815,In_1955);
or U2742 (N_2742,In_754,In_285);
and U2743 (N_2743,In_1320,In_1148);
nor U2744 (N_2744,In_785,In_622);
or U2745 (N_2745,In_1294,In_90);
xor U2746 (N_2746,In_35,In_123);
nor U2747 (N_2747,In_1002,In_157);
nand U2748 (N_2748,In_2412,In_990);
nor U2749 (N_2749,In_548,In_1112);
nor U2750 (N_2750,In_360,In_1186);
and U2751 (N_2751,In_2034,In_1142);
nand U2752 (N_2752,In_394,In_1835);
nand U2753 (N_2753,In_1372,In_2056);
and U2754 (N_2754,In_1093,In_919);
nor U2755 (N_2755,In_1208,In_2195);
nor U2756 (N_2756,In_480,In_238);
and U2757 (N_2757,In_1092,In_25);
nor U2758 (N_2758,In_2316,In_1186);
and U2759 (N_2759,In_2258,In_2424);
xnor U2760 (N_2760,In_782,In_805);
or U2761 (N_2761,In_1769,In_910);
nand U2762 (N_2762,In_2356,In_936);
nor U2763 (N_2763,In_267,In_2016);
nor U2764 (N_2764,In_2343,In_78);
xnor U2765 (N_2765,In_760,In_1747);
nand U2766 (N_2766,In_1953,In_596);
or U2767 (N_2767,In_710,In_324);
nand U2768 (N_2768,In_1672,In_2236);
xor U2769 (N_2769,In_487,In_105);
nor U2770 (N_2770,In_848,In_1097);
nor U2771 (N_2771,In_1605,In_110);
and U2772 (N_2772,In_1304,In_606);
nor U2773 (N_2773,In_660,In_1908);
and U2774 (N_2774,In_817,In_90);
and U2775 (N_2775,In_668,In_1028);
xnor U2776 (N_2776,In_804,In_1569);
xor U2777 (N_2777,In_583,In_1311);
nand U2778 (N_2778,In_1145,In_1511);
or U2779 (N_2779,In_1023,In_2420);
or U2780 (N_2780,In_102,In_1434);
and U2781 (N_2781,In_1463,In_88);
nor U2782 (N_2782,In_184,In_300);
and U2783 (N_2783,In_1170,In_1979);
nand U2784 (N_2784,In_889,In_1911);
or U2785 (N_2785,In_1184,In_1578);
nand U2786 (N_2786,In_1928,In_2350);
nand U2787 (N_2787,In_6,In_966);
and U2788 (N_2788,In_2041,In_332);
nor U2789 (N_2789,In_916,In_573);
xnor U2790 (N_2790,In_659,In_1390);
nand U2791 (N_2791,In_1528,In_694);
nand U2792 (N_2792,In_1122,In_1279);
nand U2793 (N_2793,In_1792,In_2211);
nor U2794 (N_2794,In_1301,In_2119);
nand U2795 (N_2795,In_1115,In_1201);
nand U2796 (N_2796,In_1575,In_1726);
nor U2797 (N_2797,In_826,In_1570);
nor U2798 (N_2798,In_997,In_948);
or U2799 (N_2799,In_1872,In_1640);
nor U2800 (N_2800,In_1159,In_1724);
xnor U2801 (N_2801,In_2098,In_2449);
nor U2802 (N_2802,In_257,In_1232);
nor U2803 (N_2803,In_1577,In_1771);
nand U2804 (N_2804,In_328,In_554);
and U2805 (N_2805,In_1953,In_1269);
and U2806 (N_2806,In_1450,In_45);
nand U2807 (N_2807,In_1512,In_1812);
xnor U2808 (N_2808,In_1807,In_1247);
or U2809 (N_2809,In_606,In_858);
nor U2810 (N_2810,In_1194,In_981);
nand U2811 (N_2811,In_1982,In_1474);
xnor U2812 (N_2812,In_1670,In_486);
nand U2813 (N_2813,In_885,In_1815);
or U2814 (N_2814,In_2290,In_608);
nand U2815 (N_2815,In_1482,In_1346);
nor U2816 (N_2816,In_1024,In_300);
nand U2817 (N_2817,In_1185,In_1558);
nand U2818 (N_2818,In_881,In_1902);
or U2819 (N_2819,In_514,In_167);
xor U2820 (N_2820,In_658,In_2417);
nor U2821 (N_2821,In_2186,In_898);
and U2822 (N_2822,In_1859,In_1067);
nor U2823 (N_2823,In_2157,In_1779);
nor U2824 (N_2824,In_1902,In_1781);
and U2825 (N_2825,In_1172,In_2155);
nand U2826 (N_2826,In_632,In_256);
nand U2827 (N_2827,In_728,In_1318);
nand U2828 (N_2828,In_1960,In_997);
xnor U2829 (N_2829,In_1323,In_1185);
and U2830 (N_2830,In_482,In_112);
or U2831 (N_2831,In_2,In_534);
and U2832 (N_2832,In_1068,In_1424);
nand U2833 (N_2833,In_2358,In_729);
xor U2834 (N_2834,In_2407,In_80);
nor U2835 (N_2835,In_1201,In_454);
nand U2836 (N_2836,In_1681,In_2486);
xnor U2837 (N_2837,In_411,In_376);
or U2838 (N_2838,In_2460,In_243);
and U2839 (N_2839,In_1963,In_654);
nand U2840 (N_2840,In_1078,In_1319);
xor U2841 (N_2841,In_23,In_2353);
and U2842 (N_2842,In_474,In_747);
nor U2843 (N_2843,In_1048,In_2386);
and U2844 (N_2844,In_527,In_620);
and U2845 (N_2845,In_2131,In_412);
nor U2846 (N_2846,In_1925,In_1821);
nor U2847 (N_2847,In_1683,In_664);
or U2848 (N_2848,In_1784,In_1686);
or U2849 (N_2849,In_955,In_816);
nand U2850 (N_2850,In_462,In_471);
nor U2851 (N_2851,In_382,In_524);
nor U2852 (N_2852,In_197,In_2066);
nor U2853 (N_2853,In_937,In_1845);
nor U2854 (N_2854,In_1022,In_645);
xor U2855 (N_2855,In_2412,In_2396);
or U2856 (N_2856,In_921,In_1293);
nand U2857 (N_2857,In_954,In_2429);
or U2858 (N_2858,In_941,In_2007);
and U2859 (N_2859,In_1686,In_36);
and U2860 (N_2860,In_1135,In_1448);
or U2861 (N_2861,In_2322,In_2233);
xor U2862 (N_2862,In_2309,In_648);
or U2863 (N_2863,In_2030,In_1999);
nand U2864 (N_2864,In_2087,In_1232);
nor U2865 (N_2865,In_2088,In_438);
nor U2866 (N_2866,In_2454,In_99);
or U2867 (N_2867,In_1602,In_114);
nand U2868 (N_2868,In_1242,In_391);
or U2869 (N_2869,In_155,In_172);
nor U2870 (N_2870,In_2341,In_933);
nand U2871 (N_2871,In_1748,In_1367);
nand U2872 (N_2872,In_110,In_2081);
and U2873 (N_2873,In_2291,In_792);
and U2874 (N_2874,In_1980,In_1265);
or U2875 (N_2875,In_1742,In_1197);
or U2876 (N_2876,In_1976,In_1653);
nor U2877 (N_2877,In_2405,In_665);
and U2878 (N_2878,In_1567,In_2093);
nand U2879 (N_2879,In_2272,In_2057);
or U2880 (N_2880,In_2054,In_2477);
nand U2881 (N_2881,In_1934,In_1635);
xnor U2882 (N_2882,In_1822,In_1296);
nor U2883 (N_2883,In_944,In_419);
and U2884 (N_2884,In_1999,In_624);
nor U2885 (N_2885,In_981,In_1501);
nor U2886 (N_2886,In_2128,In_75);
nand U2887 (N_2887,In_384,In_707);
or U2888 (N_2888,In_2385,In_933);
nand U2889 (N_2889,In_1168,In_1626);
xnor U2890 (N_2890,In_2046,In_435);
xor U2891 (N_2891,In_502,In_1755);
nor U2892 (N_2892,In_288,In_1697);
or U2893 (N_2893,In_1779,In_243);
or U2894 (N_2894,In_1268,In_942);
nand U2895 (N_2895,In_1612,In_104);
or U2896 (N_2896,In_1508,In_2087);
or U2897 (N_2897,In_1519,In_671);
nand U2898 (N_2898,In_1497,In_2134);
nor U2899 (N_2899,In_210,In_978);
and U2900 (N_2900,In_1911,In_476);
nand U2901 (N_2901,In_66,In_1573);
nand U2902 (N_2902,In_2293,In_2306);
and U2903 (N_2903,In_607,In_2101);
xnor U2904 (N_2904,In_2332,In_472);
nand U2905 (N_2905,In_577,In_1015);
nor U2906 (N_2906,In_1798,In_1743);
and U2907 (N_2907,In_199,In_1238);
and U2908 (N_2908,In_864,In_305);
or U2909 (N_2909,In_1470,In_1855);
nor U2910 (N_2910,In_2300,In_1113);
or U2911 (N_2911,In_32,In_1850);
and U2912 (N_2912,In_1089,In_1531);
and U2913 (N_2913,In_1110,In_1050);
or U2914 (N_2914,In_1659,In_1107);
nor U2915 (N_2915,In_60,In_287);
and U2916 (N_2916,In_1755,In_728);
nor U2917 (N_2917,In_356,In_1004);
and U2918 (N_2918,In_2121,In_1434);
or U2919 (N_2919,In_1113,In_1308);
nand U2920 (N_2920,In_1165,In_626);
and U2921 (N_2921,In_397,In_1895);
nand U2922 (N_2922,In_1402,In_2121);
or U2923 (N_2923,In_2138,In_1071);
xnor U2924 (N_2924,In_1564,In_1517);
and U2925 (N_2925,In_1942,In_835);
and U2926 (N_2926,In_1480,In_2195);
nor U2927 (N_2927,In_102,In_1678);
or U2928 (N_2928,In_1982,In_915);
and U2929 (N_2929,In_2120,In_2233);
nand U2930 (N_2930,In_613,In_369);
nand U2931 (N_2931,In_2071,In_860);
nor U2932 (N_2932,In_40,In_1291);
nand U2933 (N_2933,In_248,In_742);
nor U2934 (N_2934,In_2461,In_113);
or U2935 (N_2935,In_431,In_441);
nor U2936 (N_2936,In_977,In_1593);
or U2937 (N_2937,In_749,In_154);
nor U2938 (N_2938,In_1509,In_1386);
nand U2939 (N_2939,In_736,In_1678);
nand U2940 (N_2940,In_1543,In_1837);
xor U2941 (N_2941,In_1297,In_2058);
nor U2942 (N_2942,In_1994,In_1730);
nand U2943 (N_2943,In_1481,In_838);
nand U2944 (N_2944,In_2006,In_1749);
nor U2945 (N_2945,In_1778,In_1722);
xnor U2946 (N_2946,In_1801,In_1748);
nor U2947 (N_2947,In_2273,In_2498);
and U2948 (N_2948,In_849,In_34);
xnor U2949 (N_2949,In_1568,In_2031);
or U2950 (N_2950,In_1514,In_1466);
nor U2951 (N_2951,In_1436,In_1365);
nor U2952 (N_2952,In_966,In_2049);
or U2953 (N_2953,In_321,In_1388);
nor U2954 (N_2954,In_1600,In_1890);
and U2955 (N_2955,In_2382,In_1159);
nand U2956 (N_2956,In_18,In_2076);
nor U2957 (N_2957,In_701,In_1498);
nor U2958 (N_2958,In_585,In_1679);
and U2959 (N_2959,In_730,In_1878);
xor U2960 (N_2960,In_1092,In_140);
or U2961 (N_2961,In_322,In_484);
nand U2962 (N_2962,In_1881,In_688);
and U2963 (N_2963,In_2252,In_2262);
or U2964 (N_2964,In_1090,In_1878);
and U2965 (N_2965,In_160,In_683);
or U2966 (N_2966,In_2254,In_2388);
and U2967 (N_2967,In_1470,In_795);
and U2968 (N_2968,In_2188,In_1232);
nand U2969 (N_2969,In_1430,In_2468);
or U2970 (N_2970,In_1487,In_101);
or U2971 (N_2971,In_1499,In_1073);
and U2972 (N_2972,In_1323,In_1352);
and U2973 (N_2973,In_2109,In_96);
nand U2974 (N_2974,In_1631,In_221);
nor U2975 (N_2975,In_1971,In_663);
nor U2976 (N_2976,In_211,In_2292);
or U2977 (N_2977,In_1335,In_1393);
nor U2978 (N_2978,In_1392,In_1737);
or U2979 (N_2979,In_1891,In_2108);
or U2980 (N_2980,In_1355,In_39);
nand U2981 (N_2981,In_1655,In_1838);
or U2982 (N_2982,In_1657,In_2231);
or U2983 (N_2983,In_790,In_198);
or U2984 (N_2984,In_519,In_1787);
nor U2985 (N_2985,In_1142,In_2084);
nand U2986 (N_2986,In_1961,In_483);
and U2987 (N_2987,In_1180,In_1286);
and U2988 (N_2988,In_1314,In_1219);
and U2989 (N_2989,In_1982,In_698);
or U2990 (N_2990,In_2298,In_785);
xnor U2991 (N_2991,In_755,In_526);
nand U2992 (N_2992,In_247,In_137);
nor U2993 (N_2993,In_167,In_781);
xor U2994 (N_2994,In_718,In_689);
or U2995 (N_2995,In_2165,In_1479);
and U2996 (N_2996,In_1007,In_730);
or U2997 (N_2997,In_305,In_1251);
or U2998 (N_2998,In_1599,In_1913);
nor U2999 (N_2999,In_1491,In_1918);
nor U3000 (N_3000,In_1823,In_2496);
or U3001 (N_3001,In_1370,In_412);
nand U3002 (N_3002,In_386,In_1009);
and U3003 (N_3003,In_395,In_1935);
xor U3004 (N_3004,In_2108,In_2470);
and U3005 (N_3005,In_663,In_1712);
or U3006 (N_3006,In_1134,In_1404);
nor U3007 (N_3007,In_1126,In_1236);
or U3008 (N_3008,In_930,In_2231);
nor U3009 (N_3009,In_2469,In_2057);
nor U3010 (N_3010,In_433,In_666);
or U3011 (N_3011,In_974,In_2100);
and U3012 (N_3012,In_638,In_1712);
or U3013 (N_3013,In_2006,In_1932);
xor U3014 (N_3014,In_2139,In_2123);
nor U3015 (N_3015,In_314,In_1599);
nand U3016 (N_3016,In_2129,In_712);
or U3017 (N_3017,In_1025,In_636);
nand U3018 (N_3018,In_1200,In_317);
nor U3019 (N_3019,In_806,In_1550);
nor U3020 (N_3020,In_871,In_1363);
xnor U3021 (N_3021,In_2175,In_37);
and U3022 (N_3022,In_310,In_1244);
nor U3023 (N_3023,In_2303,In_928);
or U3024 (N_3024,In_1516,In_730);
or U3025 (N_3025,In_1405,In_1814);
nor U3026 (N_3026,In_2159,In_1272);
nand U3027 (N_3027,In_588,In_1445);
xnor U3028 (N_3028,In_570,In_608);
or U3029 (N_3029,In_2334,In_2102);
xnor U3030 (N_3030,In_280,In_542);
or U3031 (N_3031,In_1973,In_2490);
nand U3032 (N_3032,In_1587,In_1771);
nor U3033 (N_3033,In_674,In_1191);
and U3034 (N_3034,In_230,In_487);
and U3035 (N_3035,In_1350,In_902);
nor U3036 (N_3036,In_2233,In_2084);
and U3037 (N_3037,In_2375,In_713);
and U3038 (N_3038,In_1596,In_4);
xor U3039 (N_3039,In_1477,In_573);
or U3040 (N_3040,In_1651,In_335);
nor U3041 (N_3041,In_1734,In_333);
or U3042 (N_3042,In_1537,In_833);
or U3043 (N_3043,In_1464,In_1356);
nor U3044 (N_3044,In_1640,In_1873);
nor U3045 (N_3045,In_810,In_1645);
and U3046 (N_3046,In_365,In_663);
nand U3047 (N_3047,In_2332,In_127);
and U3048 (N_3048,In_301,In_2079);
nand U3049 (N_3049,In_8,In_511);
nor U3050 (N_3050,In_1726,In_2317);
nand U3051 (N_3051,In_2144,In_1992);
nand U3052 (N_3052,In_1814,In_501);
and U3053 (N_3053,In_260,In_2362);
or U3054 (N_3054,In_917,In_249);
nand U3055 (N_3055,In_1319,In_1419);
nand U3056 (N_3056,In_2128,In_838);
or U3057 (N_3057,In_2215,In_599);
nor U3058 (N_3058,In_1934,In_279);
or U3059 (N_3059,In_855,In_1915);
nor U3060 (N_3060,In_1570,In_1696);
nand U3061 (N_3061,In_659,In_1906);
or U3062 (N_3062,In_259,In_1938);
nor U3063 (N_3063,In_802,In_806);
and U3064 (N_3064,In_762,In_1932);
and U3065 (N_3065,In_432,In_475);
nand U3066 (N_3066,In_2280,In_520);
nand U3067 (N_3067,In_97,In_302);
xnor U3068 (N_3068,In_664,In_485);
or U3069 (N_3069,In_1712,In_565);
and U3070 (N_3070,In_2437,In_2065);
nor U3071 (N_3071,In_1680,In_1994);
and U3072 (N_3072,In_2053,In_1341);
nor U3073 (N_3073,In_1766,In_1949);
nor U3074 (N_3074,In_447,In_713);
nor U3075 (N_3075,In_837,In_2139);
nor U3076 (N_3076,In_1671,In_1663);
xor U3077 (N_3077,In_2160,In_1696);
and U3078 (N_3078,In_932,In_1737);
nor U3079 (N_3079,In_759,In_714);
or U3080 (N_3080,In_1254,In_542);
and U3081 (N_3081,In_189,In_1302);
and U3082 (N_3082,In_1920,In_378);
nor U3083 (N_3083,In_1223,In_1422);
nand U3084 (N_3084,In_1308,In_1430);
nor U3085 (N_3085,In_1394,In_220);
nand U3086 (N_3086,In_1537,In_2066);
xnor U3087 (N_3087,In_2140,In_2358);
and U3088 (N_3088,In_1875,In_808);
or U3089 (N_3089,In_1736,In_798);
and U3090 (N_3090,In_1403,In_1410);
xnor U3091 (N_3091,In_1410,In_139);
nor U3092 (N_3092,In_1753,In_1975);
nand U3093 (N_3093,In_2415,In_2307);
nor U3094 (N_3094,In_607,In_513);
nand U3095 (N_3095,In_804,In_1861);
and U3096 (N_3096,In_1208,In_1273);
xnor U3097 (N_3097,In_1035,In_1011);
nor U3098 (N_3098,In_360,In_1591);
nor U3099 (N_3099,In_1908,In_1207);
nor U3100 (N_3100,In_2352,In_1043);
and U3101 (N_3101,In_337,In_1938);
or U3102 (N_3102,In_2258,In_573);
nor U3103 (N_3103,In_1046,In_2290);
nor U3104 (N_3104,In_408,In_36);
and U3105 (N_3105,In_836,In_1162);
or U3106 (N_3106,In_859,In_1351);
and U3107 (N_3107,In_1539,In_1379);
xor U3108 (N_3108,In_1352,In_1907);
and U3109 (N_3109,In_371,In_1699);
nand U3110 (N_3110,In_708,In_370);
nor U3111 (N_3111,In_669,In_1257);
nand U3112 (N_3112,In_368,In_2178);
nor U3113 (N_3113,In_330,In_1833);
xor U3114 (N_3114,In_2245,In_186);
xnor U3115 (N_3115,In_412,In_817);
xnor U3116 (N_3116,In_1464,In_1185);
nor U3117 (N_3117,In_1795,In_1686);
nand U3118 (N_3118,In_1296,In_1925);
or U3119 (N_3119,In_2100,In_830);
nor U3120 (N_3120,In_1197,In_1852);
nor U3121 (N_3121,In_2357,In_2276);
nor U3122 (N_3122,In_673,In_2272);
and U3123 (N_3123,In_567,In_1519);
or U3124 (N_3124,In_1994,In_256);
nand U3125 (N_3125,N_945,N_2625);
or U3126 (N_3126,N_1910,N_2457);
or U3127 (N_3127,N_771,N_385);
and U3128 (N_3128,N_1208,N_1893);
nor U3129 (N_3129,N_1666,N_1495);
nand U3130 (N_3130,N_3057,N_151);
nand U3131 (N_3131,N_2251,N_2581);
nor U3132 (N_3132,N_1009,N_737);
and U3133 (N_3133,N_2160,N_2245);
nor U3134 (N_3134,N_40,N_336);
and U3135 (N_3135,N_280,N_637);
xnor U3136 (N_3136,N_1076,N_1891);
nand U3137 (N_3137,N_2173,N_1122);
nand U3138 (N_3138,N_2656,N_332);
xor U3139 (N_3139,N_784,N_2159);
or U3140 (N_3140,N_1583,N_342);
and U3141 (N_3141,N_1657,N_2341);
and U3142 (N_3142,N_1106,N_1873);
nor U3143 (N_3143,N_2229,N_1280);
nand U3144 (N_3144,N_2301,N_2793);
nor U3145 (N_3145,N_2682,N_3053);
nand U3146 (N_3146,N_1047,N_1257);
xnor U3147 (N_3147,N_965,N_113);
and U3148 (N_3148,N_2823,N_193);
or U3149 (N_3149,N_2769,N_1236);
or U3150 (N_3150,N_2700,N_532);
nor U3151 (N_3151,N_2056,N_2760);
or U3152 (N_3152,N_2427,N_1648);
or U3153 (N_3153,N_772,N_2322);
and U3154 (N_3154,N_2943,N_2630);
nand U3155 (N_3155,N_182,N_1405);
nand U3156 (N_3156,N_2189,N_2812);
xor U3157 (N_3157,N_2932,N_1478);
and U3158 (N_3158,N_1718,N_844);
or U3159 (N_3159,N_1810,N_821);
and U3160 (N_3160,N_155,N_2207);
nand U3161 (N_3161,N_1414,N_73);
or U3162 (N_3162,N_3113,N_1744);
and U3163 (N_3163,N_243,N_2406);
nand U3164 (N_3164,N_222,N_1113);
nand U3165 (N_3165,N_1221,N_998);
nor U3166 (N_3166,N_934,N_223);
nor U3167 (N_3167,N_2255,N_261);
or U3168 (N_3168,N_2277,N_761);
and U3169 (N_3169,N_443,N_1282);
and U3170 (N_3170,N_160,N_747);
nand U3171 (N_3171,N_2551,N_87);
or U3172 (N_3172,N_136,N_529);
or U3173 (N_3173,N_2832,N_2208);
xnor U3174 (N_3174,N_1838,N_1289);
nor U3175 (N_3175,N_1929,N_1480);
xor U3176 (N_3176,N_0,N_403);
or U3177 (N_3177,N_1402,N_1259);
and U3178 (N_3178,N_76,N_1630);
or U3179 (N_3179,N_835,N_2090);
and U3180 (N_3180,N_2980,N_179);
xnor U3181 (N_3181,N_2047,N_1541);
nor U3182 (N_3182,N_2120,N_1870);
xnor U3183 (N_3183,N_1256,N_690);
and U3184 (N_3184,N_834,N_1129);
nor U3185 (N_3185,N_18,N_3118);
nor U3186 (N_3186,N_1748,N_1918);
nand U3187 (N_3187,N_440,N_1215);
and U3188 (N_3188,N_1363,N_1501);
nand U3189 (N_3189,N_1439,N_477);
xor U3190 (N_3190,N_3007,N_1373);
or U3191 (N_3191,N_399,N_1375);
nor U3192 (N_3192,N_1885,N_1612);
or U3193 (N_3193,N_2535,N_1070);
nor U3194 (N_3194,N_1824,N_409);
nand U3195 (N_3195,N_3115,N_2973);
nand U3196 (N_3196,N_2006,N_2580);
nor U3197 (N_3197,N_1120,N_2368);
nor U3198 (N_3198,N_2717,N_2830);
nor U3199 (N_3199,N_2051,N_2136);
nor U3200 (N_3200,N_1174,N_513);
or U3201 (N_3201,N_871,N_1328);
nand U3202 (N_3202,N_2171,N_928);
and U3203 (N_3203,N_1258,N_338);
and U3204 (N_3204,N_1344,N_2305);
nor U3205 (N_3205,N_2704,N_1287);
xor U3206 (N_3206,N_273,N_1529);
and U3207 (N_3207,N_517,N_561);
nor U3208 (N_3208,N_2519,N_1551);
and U3209 (N_3209,N_1493,N_3055);
xor U3210 (N_3210,N_674,N_2435);
xnor U3211 (N_3211,N_398,N_1710);
nand U3212 (N_3212,N_1720,N_382);
nand U3213 (N_3213,N_2963,N_2058);
and U3214 (N_3214,N_226,N_150);
nor U3215 (N_3215,N_363,N_670);
and U3216 (N_3216,N_1051,N_1762);
and U3217 (N_3217,N_1865,N_1845);
or U3218 (N_3218,N_2706,N_2050);
nand U3219 (N_3219,N_1152,N_446);
or U3220 (N_3220,N_1453,N_1996);
nor U3221 (N_3221,N_251,N_2137);
nand U3222 (N_3222,N_2312,N_2602);
or U3223 (N_3223,N_2903,N_2228);
and U3224 (N_3224,N_705,N_476);
and U3225 (N_3225,N_1068,N_2086);
nor U3226 (N_3226,N_3033,N_2697);
nor U3227 (N_3227,N_717,N_2773);
nor U3228 (N_3228,N_990,N_2079);
nand U3229 (N_3229,N_2088,N_754);
or U3230 (N_3230,N_1823,N_692);
xor U3231 (N_3231,N_2799,N_1192);
nand U3232 (N_3232,N_3059,N_1341);
and U3233 (N_3233,N_1046,N_2092);
or U3234 (N_3234,N_1950,N_2397);
or U3235 (N_3235,N_269,N_495);
and U3236 (N_3236,N_2095,N_1124);
nand U3237 (N_3237,N_1981,N_1568);
or U3238 (N_3238,N_1246,N_2611);
or U3239 (N_3239,N_3048,N_842);
nor U3240 (N_3240,N_1136,N_2779);
nor U3241 (N_3241,N_1456,N_101);
or U3242 (N_3242,N_2357,N_1254);
nor U3243 (N_3243,N_1677,N_2867);
and U3244 (N_3244,N_1734,N_833);
and U3245 (N_3245,N_882,N_1274);
or U3246 (N_3246,N_819,N_1108);
nor U3247 (N_3247,N_2100,N_572);
and U3248 (N_3248,N_662,N_171);
xor U3249 (N_3249,N_2096,N_2216);
and U3250 (N_3250,N_704,N_2895);
or U3251 (N_3251,N_1735,N_2547);
xnor U3252 (N_3252,N_1085,N_1242);
or U3253 (N_3253,N_1639,N_2371);
and U3254 (N_3254,N_907,N_2914);
nor U3255 (N_3255,N_2673,N_130);
nor U3256 (N_3256,N_1022,N_324);
nor U3257 (N_3257,N_1105,N_797);
xor U3258 (N_3258,N_1925,N_1755);
or U3259 (N_3259,N_2787,N_2707);
nand U3260 (N_3260,N_327,N_1275);
xor U3261 (N_3261,N_1017,N_1978);
and U3262 (N_3262,N_836,N_144);
or U3263 (N_3263,N_299,N_1010);
or U3264 (N_3264,N_330,N_2569);
nor U3265 (N_3265,N_210,N_2178);
and U3266 (N_3266,N_2885,N_1489);
or U3267 (N_3267,N_59,N_1969);
nand U3268 (N_3268,N_2572,N_2545);
nor U3269 (N_3269,N_1071,N_2174);
nand U3270 (N_3270,N_2621,N_1708);
or U3271 (N_3271,N_633,N_2113);
nor U3272 (N_3272,N_2157,N_500);
nand U3273 (N_3273,N_271,N_1768);
nand U3274 (N_3274,N_1619,N_1594);
and U3275 (N_3275,N_1695,N_693);
nand U3276 (N_3276,N_1315,N_2380);
and U3277 (N_3277,N_1726,N_1798);
or U3278 (N_3278,N_2195,N_3001);
nor U3279 (N_3279,N_663,N_287);
nor U3280 (N_3280,N_1880,N_1386);
nand U3281 (N_3281,N_2784,N_743);
or U3282 (N_3282,N_2664,N_1743);
or U3283 (N_3283,N_951,N_2453);
nand U3284 (N_3284,N_541,N_3109);
or U3285 (N_3285,N_511,N_1988);
and U3286 (N_3286,N_460,N_539);
nor U3287 (N_3287,N_1625,N_3079);
nor U3288 (N_3288,N_1788,N_1055);
and U3289 (N_3289,N_2484,N_388);
and U3290 (N_3290,N_1252,N_3008);
or U3291 (N_3291,N_2358,N_163);
xnor U3292 (N_3292,N_368,N_329);
or U3293 (N_3293,N_1939,N_1214);
xor U3294 (N_3294,N_2996,N_466);
or U3295 (N_3295,N_2951,N_2643);
or U3296 (N_3296,N_3060,N_1596);
nor U3297 (N_3297,N_2893,N_2711);
and U3298 (N_3298,N_570,N_2199);
or U3299 (N_3299,N_11,N_2953);
or U3300 (N_3300,N_28,N_2532);
nand U3301 (N_3301,N_1526,N_228);
nor U3302 (N_3302,N_1787,N_926);
nor U3303 (N_3303,N_1503,N_1652);
or U3304 (N_3304,N_864,N_830);
nor U3305 (N_3305,N_1818,N_2029);
or U3306 (N_3306,N_1429,N_2510);
and U3307 (N_3307,N_1904,N_499);
and U3308 (N_3308,N_818,N_3010);
nor U3309 (N_3309,N_555,N_581);
nand U3310 (N_3310,N_1466,N_2946);
and U3311 (N_3311,N_1595,N_1806);
nor U3312 (N_3312,N_321,N_34);
nor U3313 (N_3313,N_162,N_1143);
nor U3314 (N_3314,N_2858,N_2729);
xor U3315 (N_3315,N_1107,N_2655);
nor U3316 (N_3316,N_2472,N_9);
nor U3317 (N_3317,N_141,N_783);
and U3318 (N_3318,N_2814,N_3051);
nand U3319 (N_3319,N_3075,N_765);
or U3320 (N_3320,N_758,N_1669);
and U3321 (N_3321,N_413,N_1723);
nand U3322 (N_3322,N_571,N_120);
or U3323 (N_3323,N_2109,N_291);
xor U3324 (N_3324,N_69,N_849);
or U3325 (N_3325,N_2504,N_2940);
xor U3326 (N_3326,N_964,N_573);
and U3327 (N_3327,N_2078,N_1977);
nor U3328 (N_3328,N_929,N_2146);
and U3329 (N_3329,N_1922,N_2891);
or U3330 (N_3330,N_2233,N_183);
and U3331 (N_3331,N_25,N_974);
and U3332 (N_3332,N_1229,N_1211);
and U3333 (N_3333,N_445,N_1767);
nand U3334 (N_3334,N_1225,N_1029);
xor U3335 (N_3335,N_127,N_2181);
nand U3336 (N_3336,N_2278,N_2298);
or U3337 (N_3337,N_2281,N_2549);
xnor U3338 (N_3338,N_1004,N_568);
nor U3339 (N_3339,N_2937,N_2169);
or U3340 (N_3340,N_153,N_1623);
or U3341 (N_3341,N_1294,N_1430);
nand U3342 (N_3342,N_841,N_1878);
nor U3343 (N_3343,N_795,N_2496);
and U3344 (N_3344,N_1682,N_488);
and U3345 (N_3345,N_682,N_905);
nand U3346 (N_3346,N_1314,N_1464);
or U3347 (N_3347,N_256,N_458);
nand U3348 (N_3348,N_1005,N_3000);
nor U3349 (N_3349,N_126,N_2520);
nand U3350 (N_3350,N_139,N_230);
and U3351 (N_3351,N_2000,N_2220);
xor U3352 (N_3352,N_1799,N_2498);
nor U3353 (N_3353,N_2486,N_2360);
nor U3354 (N_3354,N_2663,N_2796);
nand U3355 (N_3355,N_756,N_2437);
and U3356 (N_3356,N_975,N_991);
and U3357 (N_3357,N_190,N_790);
nand U3358 (N_3358,N_2600,N_1839);
nand U3359 (N_3359,N_2882,N_2884);
and U3360 (N_3360,N_198,N_240);
and U3361 (N_3361,N_1132,N_2023);
nand U3362 (N_3362,N_421,N_563);
xor U3363 (N_3363,N_52,N_3088);
xnor U3364 (N_3364,N_1813,N_2657);
nand U3365 (N_3365,N_1853,N_2124);
nand U3366 (N_3366,N_1597,N_31);
nand U3367 (N_3367,N_1423,N_1329);
nor U3368 (N_3368,N_1976,N_132);
nand U3369 (N_3369,N_2755,N_938);
nor U3370 (N_3370,N_2046,N_1616);
nand U3371 (N_3371,N_669,N_2751);
or U3372 (N_3372,N_1425,N_1559);
or U3373 (N_3373,N_3030,N_644);
or U3374 (N_3374,N_97,N_265);
and U3375 (N_3375,N_195,N_2405);
nand U3376 (N_3376,N_1002,N_897);
nand U3377 (N_3377,N_931,N_673);
xnor U3378 (N_3378,N_2501,N_3083);
and U3379 (N_3379,N_2014,N_184);
nor U3380 (N_3380,N_253,N_392);
nor U3381 (N_3381,N_1808,N_2919);
or U3382 (N_3382,N_2587,N_1069);
and U3383 (N_3383,N_400,N_1760);
and U3384 (N_3384,N_595,N_2622);
and U3385 (N_3385,N_1779,N_1956);
nand U3386 (N_3386,N_918,N_481);
xor U3387 (N_3387,N_1674,N_254);
or U3388 (N_3388,N_507,N_293);
nand U3389 (N_3389,N_2708,N_2552);
nor U3390 (N_3390,N_2144,N_1027);
nor U3391 (N_3391,N_2333,N_1484);
nor U3392 (N_3392,N_1947,N_394);
or U3393 (N_3393,N_1602,N_5);
and U3394 (N_3394,N_1585,N_1292);
nor U3395 (N_3395,N_1919,N_107);
or U3396 (N_3396,N_903,N_736);
or U3397 (N_3397,N_351,N_1131);
nor U3398 (N_3398,N_20,N_1795);
and U3399 (N_3399,N_920,N_828);
or U3400 (N_3400,N_1512,N_2597);
or U3401 (N_3401,N_815,N_623);
nor U3402 (N_3402,N_1745,N_1620);
xnor U3403 (N_3403,N_2458,N_2723);
or U3404 (N_3404,N_2346,N_2045);
and U3405 (N_3405,N_2138,N_1569);
xnor U3406 (N_3406,N_1097,N_285);
nor U3407 (N_3407,N_1624,N_764);
or U3408 (N_3408,N_1383,N_2410);
xor U3409 (N_3409,N_1531,N_2791);
nand U3410 (N_3410,N_339,N_1575);
xor U3411 (N_3411,N_755,N_1058);
or U3412 (N_3412,N_542,N_237);
nand U3413 (N_3413,N_560,N_1213);
xor U3414 (N_3414,N_1738,N_1642);
or U3415 (N_3415,N_2969,N_909);
nor U3416 (N_3416,N_2645,N_2678);
and U3417 (N_3417,N_2020,N_3114);
or U3418 (N_3418,N_2082,N_2741);
xor U3419 (N_3419,N_2221,N_1933);
or U3420 (N_3420,N_1586,N_427);
or U3421 (N_3421,N_346,N_1632);
and U3422 (N_3422,N_799,N_64);
xnor U3423 (N_3423,N_1992,N_1295);
xnor U3424 (N_3424,N_1794,N_2637);
nor U3425 (N_3425,N_1509,N_1308);
xnor U3426 (N_3426,N_534,N_2147);
and U3427 (N_3427,N_2231,N_2854);
nand U3428 (N_3428,N_483,N_364);
xnor U3429 (N_3429,N_2263,N_565);
nor U3430 (N_3430,N_1693,N_2703);
and U3431 (N_3431,N_1067,N_714);
nor U3432 (N_3432,N_2665,N_1158);
and U3433 (N_3433,N_1442,N_464);
nand U3434 (N_3434,N_703,N_391);
or U3435 (N_3435,N_1326,N_1157);
nand U3436 (N_3436,N_2289,N_2977);
or U3437 (N_3437,N_1944,N_2343);
nand U3438 (N_3438,N_328,N_412);
nor U3439 (N_3439,N_2469,N_2713);
and U3440 (N_3440,N_2190,N_829);
and U3441 (N_3441,N_2167,N_143);
nand U3442 (N_3442,N_3061,N_88);
and U3443 (N_3443,N_2531,N_985);
or U3444 (N_3444,N_42,N_2459);
nand U3445 (N_3445,N_2815,N_583);
nor U3446 (N_3446,N_967,N_1077);
or U3447 (N_3447,N_2982,N_1212);
and U3448 (N_3448,N_1321,N_191);
or U3449 (N_3449,N_677,N_875);
and U3450 (N_3450,N_1955,N_1990);
nand U3451 (N_3451,N_2944,N_404);
or U3452 (N_3452,N_232,N_2487);
or U3453 (N_3453,N_2164,N_2808);
nor U3454 (N_3454,N_2202,N_607);
and U3455 (N_3455,N_994,N_1921);
or U3456 (N_3456,N_2155,N_1222);
nor U3457 (N_3457,N_2416,N_2876);
and U3458 (N_3458,N_2337,N_1181);
xor U3459 (N_3459,N_58,N_3035);
and U3460 (N_3460,N_2064,N_1931);
and U3461 (N_3461,N_402,N_2870);
nor U3462 (N_3462,N_2910,N_2240);
or U3463 (N_3463,N_778,N_489);
nand U3464 (N_3464,N_879,N_2544);
nand U3465 (N_3465,N_2479,N_1886);
or U3466 (N_3466,N_2131,N_6);
nor U3467 (N_3467,N_2241,N_691);
xor U3468 (N_3468,N_196,N_1296);
nand U3469 (N_3469,N_2266,N_1237);
and U3470 (N_3470,N_1961,N_1892);
or U3471 (N_3471,N_1672,N_1604);
nor U3472 (N_3472,N_549,N_200);
xor U3473 (N_3473,N_2701,N_2502);
or U3474 (N_3474,N_667,N_1975);
or U3475 (N_3475,N_2950,N_1443);
nand U3476 (N_3476,N_2809,N_1364);
or U3477 (N_3477,N_56,N_621);
and U3478 (N_3478,N_231,N_2690);
nor U3479 (N_3479,N_2675,N_1418);
nor U3480 (N_3480,N_1075,N_1727);
or U3481 (N_3481,N_3023,N_3068);
and U3482 (N_3482,N_759,N_422);
and U3483 (N_3483,N_1087,N_393);
or U3484 (N_3484,N_1283,N_229);
or U3485 (N_3485,N_405,N_824);
nand U3486 (N_3486,N_2871,N_2738);
nor U3487 (N_3487,N_1338,N_2512);
xor U3488 (N_3488,N_1916,N_2260);
nand U3489 (N_3489,N_1888,N_1054);
or U3490 (N_3490,N_2603,N_3081);
or U3491 (N_3491,N_55,N_1525);
nand U3492 (N_3492,N_2440,N_554);
or U3493 (N_3493,N_2348,N_1902);
xor U3494 (N_3494,N_843,N_1716);
nor U3495 (N_3495,N_629,N_1681);
xor U3496 (N_3496,N_377,N_935);
nor U3497 (N_3497,N_2835,N_1532);
nand U3498 (N_3498,N_587,N_1769);
nor U3499 (N_3499,N_2890,N_2237);
and U3500 (N_3500,N_696,N_1820);
nor U3501 (N_3501,N_2062,N_438);
and U3502 (N_3502,N_1177,N_1465);
xnor U3503 (N_3503,N_17,N_335);
and U3504 (N_3504,N_1679,N_956);
nor U3505 (N_3505,N_2279,N_283);
nand U3506 (N_3506,N_2788,N_810);
nor U3507 (N_3507,N_2620,N_2444);
and U3508 (N_3508,N_2686,N_490);
or U3509 (N_3509,N_559,N_3112);
or U3510 (N_3510,N_1251,N_433);
nor U3511 (N_3511,N_2275,N_2243);
or U3512 (N_3512,N_1180,N_77);
nand U3513 (N_3513,N_2129,N_2745);
nand U3514 (N_3514,N_2771,N_1093);
nor U3515 (N_3515,N_1359,N_1731);
or U3516 (N_3516,N_1685,N_2877);
nor U3517 (N_3517,N_214,N_1590);
nand U3518 (N_3518,N_1062,N_2483);
or U3519 (N_3519,N_2500,N_1217);
or U3520 (N_3520,N_1766,N_2834);
or U3521 (N_3521,N_2443,N_376);
nand U3522 (N_3522,N_1370,N_2269);
nor U3523 (N_3523,N_1717,N_1654);
nand U3524 (N_3524,N_1757,N_2456);
nand U3525 (N_3525,N_2554,N_719);
nor U3526 (N_3526,N_248,N_426);
nor U3527 (N_3527,N_2546,N_480);
nor U3528 (N_3528,N_2777,N_683);
or U3529 (N_3529,N_2669,N_1451);
nor U3530 (N_3530,N_26,N_1118);
and U3531 (N_3531,N_249,N_2414);
and U3532 (N_3532,N_618,N_1034);
nand U3533 (N_3533,N_1833,N_2271);
and U3534 (N_3534,N_1895,N_2803);
and U3535 (N_3535,N_1842,N_1923);
nor U3536 (N_3536,N_766,N_2238);
or U3537 (N_3537,N_2857,N_744);
and U3538 (N_3538,N_774,N_167);
nand U3539 (N_3539,N_1968,N_1516);
nor U3540 (N_3540,N_128,N_2094);
xnor U3541 (N_3541,N_732,N_1140);
nor U3542 (N_3542,N_728,N_2819);
and U3543 (N_3543,N_1063,N_2753);
nor U3544 (N_3544,N_1574,N_1603);
or U3545 (N_3545,N_1518,N_798);
or U3546 (N_3546,N_1638,N_2034);
and U3547 (N_3547,N_1875,N_1013);
or U3548 (N_3548,N_2756,N_812);
nand U3549 (N_3549,N_2356,N_2370);
and U3550 (N_3550,N_2608,N_67);
xor U3551 (N_3551,N_2126,N_699);
and U3552 (N_3552,N_1154,N_3085);
nor U3553 (N_3553,N_2219,N_1410);
nor U3554 (N_3554,N_1235,N_1688);
and U3555 (N_3555,N_1534,N_2244);
and U3556 (N_3556,N_3024,N_1450);
nand U3557 (N_3557,N_207,N_2191);
nor U3558 (N_3558,N_1234,N_2567);
nand U3559 (N_3559,N_1345,N_2404);
nor U3560 (N_3560,N_1663,N_2909);
nand U3561 (N_3561,N_1894,N_2720);
and U3562 (N_3562,N_2748,N_3034);
nand U3563 (N_3563,N_1467,N_158);
or U3564 (N_3564,N_2077,N_2618);
nor U3565 (N_3565,N_1194,N_486);
or U3566 (N_3566,N_2460,N_1094);
and U3567 (N_3567,N_1378,N_2956);
and U3568 (N_3568,N_1216,N_334);
nand U3569 (N_3569,N_2846,N_145);
or U3570 (N_3570,N_2254,N_823);
xnor U3571 (N_3571,N_861,N_2605);
and U3572 (N_3572,N_910,N_2362);
nand U3573 (N_3573,N_2441,N_1340);
xnor U3574 (N_3574,N_1006,N_2206);
or U3575 (N_3575,N_1629,N_2344);
nor U3576 (N_3576,N_2847,N_1631);
and U3577 (N_3577,N_2172,N_2896);
and U3578 (N_3578,N_1288,N_550);
xor U3579 (N_3579,N_2941,N_2999);
nor U3580 (N_3580,N_1301,N_1371);
nor U3581 (N_3581,N_366,N_1736);
nand U3582 (N_3582,N_1872,N_2115);
nor U3583 (N_3583,N_1539,N_2792);
xor U3584 (N_3584,N_2538,N_2610);
nor U3585 (N_3585,N_2292,N_1200);
and U3586 (N_3586,N_2695,N_1601);
nor U3587 (N_3587,N_501,N_2227);
and U3588 (N_3588,N_3009,N_2259);
nor U3589 (N_3589,N_3005,N_2097);
nand U3590 (N_3590,N_2872,N_2525);
or U3591 (N_3591,N_2482,N_741);
and U3592 (N_3592,N_591,N_187);
xor U3593 (N_3593,N_937,N_2040);
nand U3594 (N_3594,N_3069,N_1561);
xnor U3595 (N_3595,N_264,N_2217);
and U3596 (N_3596,N_1230,N_1271);
xnor U3597 (N_3597,N_551,N_2252);
or U3598 (N_3598,N_1098,N_2421);
or U3599 (N_3599,N_2617,N_630);
or U3600 (N_3600,N_2762,N_2253);
and U3601 (N_3601,N_2452,N_1724);
nor U3602 (N_3602,N_14,N_2372);
or U3603 (N_3603,N_33,N_2661);
and U3604 (N_3604,N_2873,N_235);
and U3605 (N_3605,N_1860,N_415);
and U3606 (N_3606,N_1827,N_360);
or U3607 (N_3607,N_1206,N_424);
nor U3608 (N_3608,N_652,N_688);
and U3609 (N_3609,N_2672,N_2148);
nor U3610 (N_3610,N_1172,N_19);
and U3611 (N_3611,N_1020,N_260);
nor U3612 (N_3612,N_2627,N_117);
or U3613 (N_3613,N_2623,N_4);
nand U3614 (N_3614,N_1700,N_2736);
nand U3615 (N_3615,N_2691,N_2994);
or U3616 (N_3616,N_1519,N_2429);
nor U3617 (N_3617,N_3003,N_2447);
nand U3618 (N_3618,N_289,N_3031);
or U3619 (N_3619,N_2740,N_49);
nand U3620 (N_3620,N_471,N_131);
or U3621 (N_3621,N_1538,N_2248);
nor U3622 (N_3622,N_1809,N_85);
or U3623 (N_3623,N_562,N_1426);
or U3624 (N_3624,N_1633,N_1517);
nor U3625 (N_3625,N_1957,N_955);
nand U3626 (N_3626,N_2752,N_685);
and U3627 (N_3627,N_2288,N_3011);
nor U3628 (N_3628,N_1441,N_1249);
nor U3629 (N_3629,N_60,N_1021);
nand U3630 (N_3630,N_577,N_411);
nor U3631 (N_3631,N_1095,N_866);
and U3632 (N_3632,N_140,N_1896);
nand U3633 (N_3633,N_1658,N_2754);
nor U3634 (N_3634,N_2257,N_611);
nand U3635 (N_3635,N_651,N_2647);
nand U3636 (N_3636,N_1038,N_281);
and U3637 (N_3637,N_723,N_2382);
or U3638 (N_3638,N_2373,N_726);
and U3639 (N_3639,N_1406,N_567);
or U3640 (N_3640,N_370,N_872);
or U3641 (N_3641,N_1356,N_1404);
nand U3642 (N_3642,N_1928,N_2391);
or U3643 (N_3643,N_953,N_531);
nor U3644 (N_3644,N_2615,N_36);
nor U3645 (N_3645,N_1039,N_2070);
or U3646 (N_3646,N_2465,N_2879);
or U3647 (N_3647,N_1472,N_1764);
or U3648 (N_3648,N_2636,N_2067);
nor U3649 (N_3649,N_2574,N_1759);
xor U3650 (N_3650,N_2526,N_516);
nand U3651 (N_3651,N_1683,N_915);
nor U3652 (N_3652,N_2582,N_2924);
nand U3653 (N_3653,N_1765,N_615);
or U3654 (N_3654,N_1191,N_2401);
nor U3655 (N_3655,N_2295,N_1041);
and U3656 (N_3656,N_2677,N_762);
nand U3657 (N_3657,N_1134,N_3100);
nand U3658 (N_3658,N_1111,N_2003);
nor U3659 (N_3659,N_1876,N_3066);
nand U3660 (N_3660,N_356,N_2624);
nand U3661 (N_3661,N_1655,N_3006);
nor U3662 (N_3662,N_3121,N_1459);
or U3663 (N_3663,N_972,N_1562);
nor U3664 (N_3664,N_2749,N_890);
nand U3665 (N_3665,N_585,N_1807);
and U3666 (N_3666,N_851,N_2031);
nor U3667 (N_3667,N_2381,N_1437);
xor U3668 (N_3668,N_1830,N_1994);
nand U3669 (N_3669,N_1709,N_169);
or U3670 (N_3670,N_1974,N_2030);
and U3671 (N_3671,N_2230,N_3078);
nand U3672 (N_3672,N_625,N_2766);
or U3673 (N_3673,N_447,N_697);
nand U3674 (N_3674,N_10,N_1550);
nand U3675 (N_3675,N_2638,N_1649);
nor U3676 (N_3676,N_3028,N_1121);
nor U3677 (N_3677,N_1846,N_494);
nor U3678 (N_3678,N_1995,N_2210);
or U3679 (N_3679,N_2493,N_1758);
or U3680 (N_3680,N_2007,N_2721);
nor U3681 (N_3681,N_1312,N_2436);
nor U3682 (N_3682,N_1514,N_2415);
or U3683 (N_3683,N_1395,N_2598);
nor U3684 (N_3684,N_2820,N_430);
or U3685 (N_3685,N_1463,N_35);
and U3686 (N_3686,N_2746,N_2466);
or U3687 (N_3687,N_1115,N_1161);
and U3688 (N_3688,N_2590,N_977);
nand U3689 (N_3689,N_3016,N_3038);
and U3690 (N_3690,N_2066,N_1198);
or U3691 (N_3691,N_3067,N_1399);
or U3692 (N_3692,N_148,N_2922);
nor U3693 (N_3693,N_1515,N_1828);
and U3694 (N_3694,N_1791,N_2105);
xor U3695 (N_3695,N_2162,N_209);
nor U3696 (N_3696,N_149,N_1634);
and U3697 (N_3697,N_2511,N_2261);
nor U3698 (N_3698,N_96,N_344);
nand U3699 (N_3699,N_13,N_2595);
nor U3700 (N_3700,N_1431,N_987);
nand U3701 (N_3701,N_961,N_1913);
nand U3702 (N_3702,N_1149,N_315);
and U3703 (N_3703,N_676,N_1417);
xnor U3704 (N_3704,N_2845,N_545);
and U3705 (N_3705,N_2018,N_99);
nor U3706 (N_3706,N_1863,N_1324);
and U3707 (N_3707,N_852,N_245);
nor U3708 (N_3708,N_2196,N_410);
xnor U3709 (N_3709,N_1626,N_1366);
nand U3710 (N_3710,N_2462,N_1117);
nand U3711 (N_3711,N_1684,N_3101);
or U3712 (N_3712,N_313,N_1422);
or U3713 (N_3713,N_2781,N_2958);
and U3714 (N_3714,N_2899,N_2490);
nand U3715 (N_3715,N_1887,N_3056);
or U3716 (N_3716,N_1231,N_147);
nor U3717 (N_3717,N_2203,N_1025);
nand U3718 (N_3718,N_2232,N_301);
or U3719 (N_3719,N_452,N_3012);
and U3720 (N_3720,N_2426,N_354);
or U3721 (N_3721,N_1789,N_1028);
and U3722 (N_3722,N_712,N_68);
xor U3723 (N_3723,N_2838,N_3082);
and U3724 (N_3724,N_2601,N_401);
nor U3725 (N_3725,N_518,N_453);
nor U3726 (N_3726,N_2829,N_661);
or U3727 (N_3727,N_609,N_2329);
nor U3728 (N_3728,N_2307,N_2828);
nor U3729 (N_3729,N_361,N_2294);
nor U3730 (N_3730,N_988,N_1621);
nand U3731 (N_3731,N_22,N_1999);
nand U3732 (N_3732,N_2768,N_932);
nand U3733 (N_3733,N_2389,N_1197);
or U3734 (N_3734,N_989,N_2270);
nand U3735 (N_3735,N_432,N_1448);
xor U3736 (N_3736,N_3070,N_2361);
nand U3737 (N_3737,N_2084,N_175);
nor U3738 (N_3738,N_1722,N_456);
and U3739 (N_3739,N_1133,N_46);
nor U3740 (N_3740,N_2223,N_178);
nand U3741 (N_3741,N_1148,N_1946);
nor U3742 (N_3742,N_700,N_602);
xnor U3743 (N_3743,N_1546,N_2087);
xor U3744 (N_3744,N_3095,N_157);
or U3745 (N_3745,N_2743,N_1952);
or U3746 (N_3746,N_1365,N_161);
or U3747 (N_3747,N_707,N_1050);
nand U3748 (N_3748,N_862,N_1060);
nand U3749 (N_3749,N_913,N_2353);
and U3750 (N_3750,N_2722,N_1327);
and U3751 (N_3751,N_1742,N_110);
nand U3752 (N_3752,N_1449,N_297);
or U3753 (N_3753,N_2528,N_1413);
xnor U3754 (N_3754,N_2366,N_1018);
and U3755 (N_3755,N_1661,N_2974);
or U3756 (N_3756,N_444,N_108);
xnor U3757 (N_3757,N_2267,N_973);
nand U3758 (N_3758,N_2836,N_146);
or U3759 (N_3759,N_1874,N_1703);
nand U3760 (N_3760,N_1290,N_1384);
or U3761 (N_3761,N_679,N_1352);
or U3762 (N_3762,N_2107,N_3014);
and U3763 (N_3763,N_1647,N_70);
or U3764 (N_3764,N_1549,N_1877);
nor U3765 (N_3765,N_2102,N_1385);
nor U3766 (N_3766,N_1353,N_1866);
nor U3767 (N_3767,N_2824,N_1687);
nand U3768 (N_3768,N_1869,N_104);
xnor U3769 (N_3769,N_3027,N_1281);
nand U3770 (N_3770,N_984,N_2359);
nor U3771 (N_3771,N_465,N_406);
nand U3772 (N_3772,N_1186,N_1016);
nand U3773 (N_3773,N_362,N_1084);
and U3774 (N_3774,N_176,N_944);
and U3775 (N_3775,N_2354,N_337);
or U3776 (N_3776,N_1,N_1024);
nand U3777 (N_3777,N_2908,N_1424);
nor U3778 (N_3778,N_1219,N_2942);
or U3779 (N_3779,N_1754,N_1556);
xnor U3780 (N_3780,N_2399,N_2168);
nor U3781 (N_3781,N_2987,N_1109);
nand U3782 (N_3782,N_689,N_2135);
nor U3783 (N_3783,N_2689,N_2390);
nor U3784 (N_3784,N_941,N_1250);
or U3785 (N_3785,N_2523,N_94);
or U3786 (N_3786,N_2264,N_709);
and U3787 (N_3787,N_1110,N_2599);
and U3788 (N_3788,N_238,N_2417);
nand U3789 (N_3789,N_503,N_1775);
xnor U3790 (N_3790,N_2628,N_298);
nor U3791 (N_3791,N_725,N_659);
nor U3792 (N_3792,N_3116,N_1379);
nor U3793 (N_3793,N_2907,N_262);
nand U3794 (N_3794,N_917,N_1205);
nor U3795 (N_3795,N_420,N_1455);
or U3796 (N_3796,N_2127,N_2635);
nor U3797 (N_3797,N_845,N_889);
nand U3798 (N_3798,N_912,N_1091);
nand U3799 (N_3799,N_1160,N_2506);
and U3800 (N_3800,N_1169,N_1857);
and U3801 (N_3801,N_2327,N_1325);
and U3802 (N_3802,N_450,N_1199);
nor U3803 (N_3803,N_1232,N_3072);
or U3804 (N_3804,N_2025,N_1543);
nor U3805 (N_3805,N_2556,N_246);
nand U3806 (N_3806,N_1350,N_2296);
and U3807 (N_3807,N_1622,N_3094);
and U3808 (N_3808,N_1542,N_1577);
or U3809 (N_3809,N_1890,N_827);
nand U3810 (N_3810,N_2335,N_2995);
nor U3811 (N_3811,N_2521,N_701);
nor U3812 (N_3812,N_1797,N_2492);
nand U3813 (N_3813,N_900,N_2560);
nand U3814 (N_3814,N_2163,N_1267);
xor U3815 (N_3815,N_1741,N_154);
nor U3816 (N_3816,N_3018,N_39);
nor U3817 (N_3817,N_2536,N_1528);
nor U3818 (N_3818,N_2565,N_2376);
and U3819 (N_3819,N_2694,N_2825);
nor U3820 (N_3820,N_1427,N_168);
or U3821 (N_3821,N_2304,N_1840);
xnor U3822 (N_3822,N_2586,N_268);
and U3823 (N_3823,N_1485,N_2114);
nor U3824 (N_3824,N_1481,N_1690);
nand U3825 (N_3825,N_867,N_2328);
or U3826 (N_3826,N_2902,N_2962);
nor U3827 (N_3827,N_603,N_807);
nor U3828 (N_3828,N_2387,N_2132);
or U3829 (N_3829,N_2929,N_2222);
nand U3830 (N_3830,N_2609,N_1128);
nand U3831 (N_3831,N_2142,N_1914);
or U3832 (N_3832,N_2499,N_613);
and U3833 (N_3833,N_957,N_1447);
or U3834 (N_3834,N_2015,N_853);
nand U3835 (N_3835,N_124,N_1991);
nor U3836 (N_3836,N_2986,N_1773);
nand U3837 (N_3837,N_1960,N_1273);
nor U3838 (N_3838,N_2063,N_2968);
and U3839 (N_3839,N_2433,N_1433);
nand U3840 (N_3840,N_2964,N_1244);
or U3841 (N_3841,N_2215,N_1336);
nor U3842 (N_3842,N_259,N_2491);
nand U3843 (N_3843,N_1446,N_569);
nor U3844 (N_3844,N_2101,N_1119);
or U3845 (N_3845,N_2365,N_1293);
nor U3846 (N_3846,N_2331,N_2211);
xor U3847 (N_3847,N_2575,N_267);
or U3848 (N_3848,N_1829,N_2325);
nand U3849 (N_3849,N_2727,N_854);
and U3850 (N_3850,N_84,N_1176);
and U3851 (N_3851,N_436,N_1854);
and U3852 (N_3852,N_2235,N_1530);
xor U3853 (N_3853,N_785,N_1008);
nand U3854 (N_3854,N_2059,N_272);
xor U3855 (N_3855,N_2774,N_901);
and U3856 (N_3856,N_1276,N_1305);
and U3857 (N_3857,N_860,N_202);
or U3858 (N_3858,N_2821,N_2911);
nor U3859 (N_3859,N_203,N_79);
and U3860 (N_3860,N_1003,N_1438);
or U3861 (N_3861,N_2640,N_996);
and U3862 (N_3862,N_2844,N_2053);
nor U3863 (N_3863,N_2398,N_1592);
or U3864 (N_3864,N_2916,N_933);
nor U3865 (N_3865,N_1740,N_1476);
and U3866 (N_3866,N_1061,N_914);
or U3867 (N_3867,N_457,N_1535);
nor U3868 (N_3868,N_3042,N_2900);
or U3869 (N_3869,N_1505,N_2038);
xor U3870 (N_3870,N_1776,N_733);
and U3871 (N_3871,N_1676,N_2856);
and U3872 (N_3872,N_1973,N_2930);
and U3873 (N_3873,N_746,N_1588);
or U3874 (N_3874,N_2851,N_2110);
nor U3875 (N_3875,N_216,N_1811);
nor U3876 (N_3876,N_687,N_1403);
nor U3877 (N_3877,N_2315,N_90);
nand U3878 (N_3878,N_2481,N_536);
or U3879 (N_3879,N_982,N_1390);
nor U3880 (N_3880,N_2765,N_1591);
or U3881 (N_3881,N_2776,N_2542);
nand U3882 (N_3882,N_2103,N_1123);
nand U3883 (N_3883,N_24,N_48);
and U3884 (N_3884,N_2985,N_638);
nand U3885 (N_3885,N_616,N_2468);
or U3886 (N_3886,N_102,N_2364);
nor U3887 (N_3887,N_817,N_2175);
and U3888 (N_3888,N_1048,N_2291);
nand U3889 (N_3889,N_418,N_2300);
nor U3890 (N_3890,N_2048,N_2543);
nor U3891 (N_3891,N_2374,N_1209);
nor U3892 (N_3892,N_1335,N_2612);
nor U3893 (N_3893,N_2562,N_2297);
nor U3894 (N_3894,N_596,N_491);
and U3895 (N_3895,N_384,N_2674);
nor U3896 (N_3896,N_706,N_2226);
and U3897 (N_3897,N_1303,N_564);
nor U3898 (N_3898,N_2949,N_1367);
xnor U3899 (N_3899,N_2927,N_227);
nor U3900 (N_3900,N_2939,N_1646);
and U3901 (N_3901,N_1011,N_884);
nand U3902 (N_3902,N_1504,N_1469);
nor U3903 (N_3903,N_1477,N_1468);
nor U3904 (N_3904,N_2476,N_2651);
or U3905 (N_3905,N_2386,N_1387);
nor U3906 (N_3906,N_809,N_2177);
and U3907 (N_3907,N_3124,N_1330);
nor U3908 (N_3908,N_2170,N_2522);
xor U3909 (N_3909,N_119,N_1159);
xnor U3910 (N_3910,N_2917,N_1589);
and U3911 (N_3911,N_952,N_57);
nand U3912 (N_3912,N_2688,N_748);
and U3913 (N_3913,N_2450,N_1203);
nor U3914 (N_3914,N_1822,N_713);
and U3915 (N_3915,N_1962,N_2438);
and U3916 (N_3916,N_185,N_718);
nor U3917 (N_3917,N_3087,N_942);
and U3918 (N_3918,N_949,N_671);
nand U3919 (N_3919,N_2965,N_2377);
or U3920 (N_3920,N_1635,N_442);
and U3921 (N_3921,N_2853,N_2125);
and U3922 (N_3922,N_296,N_2757);
or U3923 (N_3923,N_2280,N_2971);
nor U3924 (N_3924,N_1460,N_367);
or U3925 (N_3925,N_2790,N_1332);
or U3926 (N_3926,N_1268,N_1670);
nand U3927 (N_3927,N_2739,N_858);
nor U3928 (N_3928,N_3020,N_1320);
nand U3929 (N_3929,N_78,N_622);
nand U3930 (N_3930,N_2878,N_38);
nor U3931 (N_3931,N_3117,N_2273);
and U3932 (N_3932,N_1560,N_2548);
or U3933 (N_3933,N_2967,N_787);
or U3934 (N_3934,N_2888,N_1023);
nand U3935 (N_3935,N_2385,N_1761);
or U3936 (N_3936,N_3098,N_2840);
and U3937 (N_3937,N_1989,N_792);
nand U3938 (N_3938,N_1705,N_612);
or U3939 (N_3939,N_658,N_159);
nand U3940 (N_3940,N_2709,N_1033);
or U3941 (N_3941,N_2576,N_540);
nand U3942 (N_3942,N_1605,N_2607);
or U3943 (N_3943,N_3047,N_1362);
nand U3944 (N_3944,N_2393,N_1196);
nand U3945 (N_3945,N_1949,N_2778);
nor U3946 (N_3946,N_1317,N_255);
nand U3947 (N_3947,N_1150,N_2679);
nand U3948 (N_3948,N_2646,N_1307);
nand U3949 (N_3949,N_553,N_927);
nor U3950 (N_3950,N_588,N_472);
and U3951 (N_3951,N_839,N_112);
and U3952 (N_3952,N_3096,N_801);
or U3953 (N_3953,N_218,N_2733);
nor U3954 (N_3954,N_1563,N_2010);
nor U3955 (N_3955,N_576,N_2471);
or U3956 (N_3956,N_1243,N_1388);
nor U3957 (N_3957,N_2886,N_311);
or U3958 (N_3958,N_1627,N_1707);
or U3959 (N_3959,N_995,N_2489);
nor U3960 (N_3960,N_891,N_30);
xor U3961 (N_3961,N_1462,N_2782);
xor U3962 (N_3962,N_1357,N_654);
nor U3963 (N_3963,N_624,N_1096);
or U3964 (N_3964,N_381,N_1730);
or U3965 (N_3965,N_1343,N_1226);
xor U3966 (N_3966,N_1600,N_434);
xor U3967 (N_3967,N_2324,N_2290);
or U3968 (N_3968,N_1671,N_1397);
and U3969 (N_3969,N_2692,N_2032);
and U3970 (N_3970,N_2898,N_2702);
or U3971 (N_3971,N_2118,N_1073);
and U3972 (N_3972,N_1696,N_1486);
nand U3973 (N_3973,N_1610,N_1571);
nand U3974 (N_3974,N_396,N_2152);
and U3975 (N_3975,N_181,N_2188);
nor U3976 (N_3976,N_1407,N_2043);
nor U3977 (N_3977,N_2375,N_1342);
or U3978 (N_3978,N_1261,N_474);
and U3979 (N_3979,N_2938,N_379);
nor U3980 (N_3980,N_1537,N_535);
nor U3981 (N_3981,N_288,N_2649);
or U3982 (N_3982,N_1239,N_848);
xor U3983 (N_3983,N_898,N_74);
or U3984 (N_3984,N_1987,N_199);
nor U3985 (N_3985,N_2687,N_454);
or U3986 (N_3986,N_2140,N_111);
and U3987 (N_3987,N_2883,N_1499);
nand U3988 (N_3988,N_1576,N_1943);
nor U3989 (N_3989,N_558,N_1668);
nand U3990 (N_3990,N_2578,N_924);
nor U3991 (N_3991,N_2422,N_720);
and U3992 (N_3992,N_1524,N_284);
xnor U3993 (N_3993,N_2505,N_1190);
nand U3994 (N_3994,N_1434,N_347);
or U3995 (N_3995,N_2413,N_646);
and U3996 (N_3996,N_2249,N_244);
nor U3997 (N_3997,N_2961,N_1747);
or U3998 (N_3998,N_962,N_1168);
xnor U3999 (N_3999,N_2764,N_2837);
xor U4000 (N_4000,N_752,N_1637);
nand U4001 (N_4001,N_2179,N_1907);
nor U4002 (N_4002,N_1558,N_1897);
xnor U4003 (N_4003,N_2396,N_525);
nand U4004 (N_4004,N_515,N_1358);
xnor U4005 (N_4005,N_2991,N_2983);
nor U4006 (N_4006,N_2514,N_2418);
or U4007 (N_4007,N_1909,N_2947);
nand U4008 (N_4008,N_3108,N_1178);
nand U4009 (N_4009,N_665,N_727);
xor U4010 (N_4010,N_478,N_632);
and U4011 (N_4011,N_2997,N_350);
nor U4012 (N_4012,N_686,N_225);
xor U4013 (N_4013,N_83,N_1868);
nand U4014 (N_4014,N_2874,N_2035);
nor U4015 (N_4015,N_1511,N_1015);
or U4016 (N_4016,N_2193,N_217);
and U4017 (N_4017,N_2204,N_1573);
nand U4018 (N_4018,N_2467,N_2284);
xor U4019 (N_4019,N_1572,N_2698);
and U4020 (N_4020,N_2533,N_204);
nor U4021 (N_4021,N_2826,N_417);
nand U4022 (N_4022,N_1617,N_2897);
or U4023 (N_4023,N_1889,N_469);
xor U4024 (N_4024,N_2785,N_3050);
or U4025 (N_4025,N_1848,N_414);
and U4026 (N_4026,N_1770,N_300);
nor U4027 (N_4027,N_1392,N_2806);
nand U4028 (N_4028,N_2816,N_597);
nand U4029 (N_4029,N_1488,N_416);
and U4030 (N_4030,N_479,N_1053);
and U4031 (N_4031,N_1905,N_2306);
or U4032 (N_4032,N_1494,N_731);
and U4033 (N_4033,N_27,N_2205);
nand U4034 (N_4034,N_2798,N_822);
nor U4035 (N_4035,N_80,N_3084);
nand U4036 (N_4036,N_711,N_514);
and U4037 (N_4037,N_2309,N_1983);
and U4038 (N_4038,N_2864,N_1471);
nor U4039 (N_4039,N_1938,N_1900);
and U4040 (N_4040,N_2,N_3073);
nand U4041 (N_4041,N_1253,N_832);
nor U4042 (N_4042,N_1971,N_341);
and U4043 (N_4043,N_2054,N_2049);
nand U4044 (N_4044,N_2928,N_1581);
nor U4045 (N_4045,N_1825,N_1316);
nor U4046 (N_4046,N_2811,N_1269);
or U4047 (N_4047,N_574,N_322);
nor U4048 (N_4048,N_2494,N_1932);
nor U4049 (N_4049,N_2022,N_1043);
nor U4050 (N_4050,N_1100,N_2654);
nor U4051 (N_4051,N_2336,N_523);
nor U4052 (N_4052,N_2461,N_2589);
xnor U4053 (N_4053,N_3025,N_302);
or U4054 (N_4054,N_664,N_2121);
and U4055 (N_4055,N_2218,N_1185);
nor U4056 (N_4056,N_2464,N_1712);
xor U4057 (N_4057,N_2213,N_2775);
nand U4058 (N_4058,N_2478,N_1871);
nand U4059 (N_4059,N_352,N_2239);
nand U4060 (N_4060,N_2419,N_462);
nor U4061 (N_4061,N_1771,N_1507);
and U4062 (N_4062,N_1153,N_114);
nor U4063 (N_4063,N_1721,N_608);
nor U4064 (N_4064,N_2080,N_2130);
nand U4065 (N_4065,N_2524,N_3026);
nand U4066 (N_4066,N_856,N_1382);
xnor U4067 (N_4067,N_2931,N_3120);
or U4068 (N_4068,N_2192,N_142);
nand U4069 (N_4069,N_2831,N_2614);
or U4070 (N_4070,N_2553,N_340);
nor U4071 (N_4071,N_1260,N_1997);
and U4072 (N_4072,N_451,N_1608);
nand U4073 (N_4073,N_528,N_1567);
nor U4074 (N_4074,N_794,N_348);
nor U4075 (N_4075,N_3106,N_1318);
or U4076 (N_4076,N_378,N_286);
or U4077 (N_4077,N_1945,N_213);
and U4078 (N_4078,N_2742,N_2061);
nor U4079 (N_4079,N_976,N_197);
or U4080 (N_4080,N_1302,N_1533);
nor U4081 (N_4081,N_1521,N_1030);
or U4082 (N_4082,N_916,N_129);
nand U4083 (N_4083,N_1012,N_3090);
and U4084 (N_4084,N_971,N_1941);
and U4085 (N_4085,N_3097,N_397);
or U4086 (N_4086,N_266,N_1165);
nand U4087 (N_4087,N_2887,N_648);
nand U4088 (N_4088,N_371,N_2041);
xor U4089 (N_4089,N_745,N_1936);
nor U4090 (N_4090,N_123,N_2842);
xnor U4091 (N_4091,N_1394,N_1272);
and U4092 (N_4092,N_1566,N_2993);
or U4093 (N_4093,N_1240,N_1954);
and U4094 (N_4094,N_2534,N_939);
and U4095 (N_4095,N_1680,N_2128);
nor U4096 (N_4096,N_610,N_1245);
or U4097 (N_4097,N_1965,N_2894);
and U4098 (N_4098,N_2807,N_2379);
or U4099 (N_4099,N_189,N_2750);
xor U4100 (N_4100,N_782,N_326);
nor U4101 (N_4101,N_1660,N_2988);
and U4102 (N_4102,N_1299,N_1915);
or U4103 (N_4103,N_1856,N_2286);
nor U4104 (N_4104,N_640,N_2394);
xor U4105 (N_4105,N_653,N_2861);
nor U4106 (N_4106,N_1408,N_604);
or U4107 (N_4107,N_2108,N_796);
and U4108 (N_4108,N_2176,N_2737);
or U4109 (N_4109,N_3022,N_2936);
nand U4110 (N_4110,N_1640,N_786);
nor U4111 (N_4111,N_1065,N_734);
nor U4112 (N_4112,N_15,N_2075);
and U4113 (N_4113,N_1368,N_601);
or U4114 (N_4114,N_1189,N_3054);
and U4115 (N_4115,N_1544,N_2566);
nor U4116 (N_4116,N_2818,N_1599);
or U4117 (N_4117,N_1337,N_672);
and U4118 (N_4118,N_2724,N_125);
nand U4119 (N_4119,N_383,N_1233);
and U4120 (N_4120,N_2153,N_2106);
nand U4121 (N_4121,N_636,N_1565);
or U4122 (N_4122,N_221,N_2420);
and U4123 (N_4123,N_2540,N_2104);
and U4124 (N_4124,N_1490,N_1339);
nand U4125 (N_4125,N_1112,N_2833);
nand U4126 (N_4126,N_2550,N_2445);
nand U4127 (N_4127,N_2004,N_1031);
nor U4128 (N_4128,N_3111,N_2272);
nand U4129 (N_4129,N_594,N_21);
nor U4130 (N_4130,N_605,N_3017);
xor U4131 (N_4131,N_2904,N_695);
and U4132 (N_4132,N_2923,N_118);
nand U4133 (N_4133,N_1934,N_2921);
or U4134 (N_4134,N_963,N_2761);
or U4135 (N_4135,N_1926,N_2772);
nor U4136 (N_4136,N_2002,N_252);
nand U4137 (N_4137,N_1906,N_103);
nor U4138 (N_4138,N_837,N_1858);
nand U4139 (N_4139,N_1618,N_1953);
nor U4140 (N_4140,N_2055,N_435);
or U4141 (N_4141,N_1224,N_2726);
nand U4142 (N_4142,N_702,N_3052);
nor U4143 (N_4143,N_2133,N_2588);
and U4144 (N_4144,N_2016,N_1461);
nor U4145 (N_4145,N_2412,N_645);
and U4146 (N_4146,N_1421,N_2859);
and U4147 (N_4147,N_1912,N_1547);
nor U4148 (N_4148,N_475,N_537);
nor U4149 (N_4149,N_1347,N_642);
nand U4150 (N_4150,N_2593,N_1920);
or U4151 (N_4151,N_1665,N_2954);
nand U4152 (N_4152,N_2313,N_502);
or U4153 (N_4153,N_1279,N_72);
nand U4154 (N_4154,N_493,N_1080);
nand U4155 (N_4155,N_1103,N_2276);
nor U4156 (N_4156,N_1187,N_1554);
nor U4157 (N_4157,N_470,N_2959);
nor U4158 (N_4158,N_239,N_1440);
nor U4159 (N_4159,N_1202,N_2074);
and U4160 (N_4160,N_3105,N_429);
nor U4161 (N_4161,N_1125,N_2008);
nand U4162 (N_4162,N_1428,N_2283);
nand U4163 (N_4163,N_194,N_2880);
or U4164 (N_4164,N_2585,N_387);
and U4165 (N_4165,N_1964,N_730);
or U4166 (N_4166,N_1615,N_1291);
nor U4167 (N_4167,N_2513,N_2978);
nand U4168 (N_4168,N_186,N_966);
and U4169 (N_4169,N_1445,N_333);
or U4170 (N_4170,N_37,N_1796);
xor U4171 (N_4171,N_45,N_7);
nand U4172 (N_4172,N_16,N_2274);
nor U4173 (N_4173,N_826,N_2920);
and U4174 (N_4174,N_643,N_1783);
and U4175 (N_4175,N_592,N_2011);
or U4176 (N_4176,N_1979,N_2156);
nand U4177 (N_4177,N_983,N_2434);
and U4178 (N_4178,N_2571,N_3062);
and U4179 (N_4179,N_408,N_992);
or U4180 (N_4180,N_2952,N_859);
or U4181 (N_4181,N_1814,N_66);
or U4182 (N_4182,N_2299,N_2889);
or U4183 (N_4183,N_1297,N_2905);
or U4184 (N_4184,N_32,N_1785);
and U4185 (N_4185,N_1804,N_2027);
or U4186 (N_4186,N_1482,N_2839);
or U4187 (N_4187,N_1774,N_1998);
nor U4188 (N_4188,N_847,N_1419);
xor U4189 (N_4189,N_911,N_895);
nor U4190 (N_4190,N_2183,N_1175);
and U4191 (N_4191,N_2242,N_1985);
nor U4192 (N_4192,N_770,N_1713);
nand U4193 (N_4193,N_1927,N_1081);
and U4194 (N_4194,N_1948,N_1114);
nor U4195 (N_4195,N_2141,N_881);
nand U4196 (N_4196,N_1416,N_1170);
or U4197 (N_4197,N_923,N_2568);
and U4198 (N_4198,N_873,N_2619);
nor U4199 (N_4199,N_773,N_1400);
nand U4200 (N_4200,N_887,N_2503);
and U4201 (N_4201,N_109,N_215);
or U4202 (N_4202,N_2081,N_95);
xnor U4203 (N_4203,N_2728,N_655);
nor U4204 (N_4204,N_979,N_582);
nand U4205 (N_4205,N_919,N_2068);
xor U4206 (N_4206,N_2639,N_250);
and U4207 (N_4207,N_1644,N_277);
nor U4208 (N_4208,N_86,N_1102);
or U4209 (N_4209,N_547,N_275);
xnor U4210 (N_4210,N_3071,N_678);
and U4211 (N_4211,N_2497,N_2480);
or U4212 (N_4212,N_310,N_82);
or U4213 (N_4213,N_2659,N_3077);
and U4214 (N_4214,N_2735,N_524);
or U4215 (N_4215,N_1300,N_3122);
and U4216 (N_4216,N_2005,N_1951);
nand U4217 (N_4217,N_1753,N_2093);
nor U4218 (N_4218,N_386,N_1587);
nand U4219 (N_4219,N_498,N_2392);
and U4220 (N_4220,N_2320,N_2145);
or U4221 (N_4221,N_1035,N_2933);
nand U4222 (N_4222,N_369,N_2881);
and U4223 (N_4223,N_2577,N_98);
or U4224 (N_4224,N_2653,N_584);
and U4225 (N_4225,N_1986,N_1673);
xor U4226 (N_4226,N_3037,N_3080);
nand U4227 (N_4227,N_1262,N_825);
or U4228 (N_4228,N_1126,N_2805);
nand U4229 (N_4229,N_2981,N_1570);
and U4230 (N_4230,N_2425,N_1746);
nand U4231 (N_4231,N_1458,N_2990);
nand U4232 (N_4232,N_1847,N_2402);
nand U4233 (N_4233,N_212,N_2326);
or U4234 (N_4234,N_71,N_1510);
nand U4235 (N_4235,N_1780,N_2813);
nor U4236 (N_4236,N_2225,N_2555);
nor U4237 (N_4237,N_1284,N_278);
and U4238 (N_4238,N_1127,N_777);
nor U4239 (N_4239,N_1884,N_1911);
nand U4240 (N_4240,N_2579,N_91);
or U4241 (N_4241,N_781,N_2648);
nor U4242 (N_4242,N_1940,N_2979);
and U4243 (N_4243,N_89,N_878);
nand U4244 (N_4244,N_1763,N_936);
or U4245 (N_4245,N_800,N_2342);
nand U4246 (N_4246,N_508,N_1584);
and U4247 (N_4247,N_389,N_2212);
nor U4248 (N_4248,N_2431,N_2347);
and U4249 (N_4249,N_544,N_2868);
xnor U4250 (N_4250,N_461,N_981);
and U4251 (N_4251,N_2558,N_2714);
nor U4252 (N_4252,N_270,N_1607);
nor U4253 (N_4253,N_1286,N_2680);
or U4254 (N_4254,N_1389,N_1377);
nand U4255 (N_4255,N_482,N_428);
nand U4256 (N_4256,N_1349,N_3036);
nand U4257 (N_4257,N_1444,N_1506);
or U4258 (N_4258,N_617,N_2875);
or U4259 (N_4259,N_1309,N_1201);
nand U4260 (N_4260,N_2039,N_1733);
and U4261 (N_4261,N_279,N_2071);
nand U4262 (N_4262,N_627,N_3029);
nor U4263 (N_4263,N_1334,N_753);
nor U4264 (N_4264,N_1101,N_2363);
nor U4265 (N_4265,N_619,N_776);
xor U4266 (N_4266,N_2563,N_2403);
nor U4267 (N_4267,N_1545,N_1164);
nand U4268 (N_4268,N_656,N_2632);
nand U4269 (N_4269,N_1210,N_2794);
nand U4270 (N_4270,N_586,N_135);
nand U4271 (N_4271,N_869,N_742);
or U4272 (N_4272,N_138,N_1801);
or U4273 (N_4273,N_2850,N_2009);
nand U4274 (N_4274,N_359,N_959);
or U4275 (N_4275,N_274,N_2065);
and U4276 (N_4276,N_2463,N_1137);
or U4277 (N_4277,N_1298,N_201);
nor U4278 (N_4278,N_1037,N_2182);
nor U4279 (N_4279,N_863,N_2662);
or U4280 (N_4280,N_325,N_2789);
or U4281 (N_4281,N_1130,N_1651);
or U4282 (N_4282,N_1372,N_2119);
or U4283 (N_4283,N_2671,N_708);
nor U4284 (N_4284,N_2180,N_1044);
nor U4285 (N_4285,N_1739,N_459);
nand U4286 (N_4286,N_2712,N_395);
nor U4287 (N_4287,N_3049,N_3032);
nor U4288 (N_4288,N_1319,N_2310);
nand U4289 (N_4289,N_814,N_92);
nor U4290 (N_4290,N_893,N_641);
or U4291 (N_4291,N_2918,N_902);
nor U4292 (N_4292,N_188,N_106);
nor U4293 (N_4293,N_2400,N_165);
and U4294 (N_4294,N_2236,N_950);
nor U4295 (N_4295,N_308,N_1835);
or U4296 (N_4296,N_3064,N_751);
nand U4297 (N_4297,N_3002,N_1984);
nor U4298 (N_4298,N_2314,N_2186);
or U4299 (N_4299,N_2758,N_419);
nand U4300 (N_4300,N_1864,N_2098);
nand U4301 (N_4301,N_1074,N_1263);
and U4302 (N_4302,N_543,N_1935);
nand U4303 (N_4303,N_2187,N_1821);
or U4304 (N_4304,N_788,N_960);
and U4305 (N_4305,N_1852,N_50);
nor U4306 (N_4306,N_2631,N_2287);
and U4307 (N_4307,N_316,N_1698);
nand U4308 (N_4308,N_1664,N_2250);
xnor U4309 (N_4309,N_811,N_1266);
nand U4310 (N_4310,N_1145,N_2935);
nor U4311 (N_4311,N_2408,N_2209);
or U4312 (N_4312,N_2705,N_578);
and U4313 (N_4313,N_721,N_2584);
and U4314 (N_4314,N_1207,N_1089);
nor U4315 (N_4315,N_208,N_986);
or U4316 (N_4316,N_3045,N_2017);
nand U4317 (N_4317,N_172,N_769);
or U4318 (N_4318,N_2488,N_1844);
nor U4319 (N_4319,N_1714,N_519);
nor U4320 (N_4320,N_1728,N_2256);
or U4321 (N_4321,N_538,N_2718);
nor U4322 (N_4322,N_505,N_520);
nor U4323 (N_4323,N_857,N_1285);
nand U4324 (N_4324,N_2670,N_1697);
nand U4325 (N_4325,N_1147,N_2975);
nand U4326 (N_4326,N_1401,N_2591);
nand U4327 (N_4327,N_2258,N_2860);
nand U4328 (N_4328,N_1659,N_93);
xnor U4329 (N_4329,N_724,N_306);
and U4330 (N_4330,N_1083,N_304);
nand U4331 (N_4331,N_2613,N_2763);
or U4332 (N_4332,N_3015,N_1223);
nor U4333 (N_4333,N_51,N_242);
or U4334 (N_4334,N_211,N_1432);
or U4335 (N_4335,N_3058,N_883);
nor U4336 (N_4336,N_1641,N_775);
nand U4337 (N_4337,N_43,N_2797);
xor U4338 (N_4338,N_1817,N_1042);
nor U4339 (N_4339,N_1522,N_1454);
xnor U4340 (N_4340,N_1826,N_1220);
or U4341 (N_4341,N_2508,N_318);
nand U4342 (N_4342,N_2912,N_1917);
nor U4343 (N_4343,N_1167,N_1470);
or U4344 (N_4344,N_954,N_1138);
and U4345 (N_4345,N_2507,N_1474);
nor U4346 (N_4346,N_1415,N_997);
nor U4347 (N_4347,N_2185,N_1849);
or U4348 (N_4348,N_487,N_2154);
nor U4349 (N_4349,N_1862,N_1255);
or U4350 (N_4350,N_241,N_425);
xor U4351 (N_4351,N_1527,N_2683);
nor U4352 (N_4352,N_1816,N_816);
and U4353 (N_4353,N_2234,N_740);
and U4354 (N_4354,N_448,N_2451);
and U4355 (N_4355,N_1553,N_789);
and U4356 (N_4356,N_2955,N_2321);
or U4357 (N_4357,N_2428,N_3104);
xnor U4358 (N_4358,N_958,N_1694);
or U4359 (N_4359,N_2224,N_2557);
or U4360 (N_4360,N_1699,N_649);
nor U4361 (N_4361,N_886,N_2841);
nand U4362 (N_4362,N_1151,N_2802);
nor U4363 (N_4363,N_2369,N_1851);
nor U4364 (N_4364,N_2527,N_2285);
and U4365 (N_4365,N_276,N_1966);
nand U4366 (N_4366,N_3021,N_2442);
nor U4367 (N_4367,N_806,N_1883);
or U4368 (N_4368,N_1007,N_2594);
or U4369 (N_4369,N_2606,N_234);
and U4370 (N_4370,N_3046,N_1473);
nor U4371 (N_4371,N_1812,N_1580);
or U4372 (N_4372,N_380,N_166);
nor U4373 (N_4373,N_1475,N_2795);
nand U4374 (N_4374,N_358,N_1879);
nor U4375 (N_4375,N_2474,N_1861);
or U4376 (N_4376,N_2184,N_224);
nor U4377 (N_4377,N_1072,N_2616);
nor U4378 (N_4378,N_1086,N_2340);
nor U4379 (N_4379,N_2069,N_1781);
and U4380 (N_4380,N_1578,N_156);
and U4381 (N_4381,N_763,N_1898);
nand U4382 (N_4382,N_2780,N_1564);
nor U4383 (N_4383,N_2699,N_2021);
nor U4384 (N_4384,N_1141,N_2111);
nor U4385 (N_4385,N_497,N_220);
nor U4386 (N_4386,N_2383,N_192);
and U4387 (N_4387,N_2515,N_1306);
xor U4388 (N_4388,N_1719,N_1715);
and U4389 (N_4389,N_2906,N_2367);
and U4390 (N_4390,N_1803,N_2351);
or U4391 (N_4391,N_1304,N_512);
and U4392 (N_4392,N_2710,N_750);
nor U4393 (N_4393,N_2112,N_437);
and U4394 (N_4394,N_593,N_439);
xor U4395 (N_4395,N_2744,N_1675);
and U4396 (N_4396,N_2564,N_2913);
and U4397 (N_4397,N_353,N_1701);
or U4398 (N_4398,N_1737,N_2073);
nand U4399 (N_4399,N_1045,N_1520);
nand U4400 (N_4400,N_2123,N_760);
and U4401 (N_4401,N_1834,N_2455);
or U4402 (N_4402,N_3110,N_2570);
nor U4403 (N_4403,N_2865,N_152);
nand U4404 (N_4404,N_666,N_390);
and U4405 (N_4405,N_1972,N_1540);
nor U4406 (N_4406,N_2134,N_2477);
nand U4407 (N_4407,N_1678,N_2517);
and U4408 (N_4408,N_2866,N_63);
nor U4409 (N_4409,N_876,N_1643);
and U4410 (N_4410,N_3107,N_1435);
and U4411 (N_4411,N_2345,N_3123);
nand U4412 (N_4412,N_1800,N_1881);
nor U4413 (N_4413,N_1348,N_3004);
or U4414 (N_4414,N_802,N_868);
or U4415 (N_4415,N_496,N_1204);
and U4416 (N_4416,N_1026,N_530);
nand U4417 (N_4417,N_2970,N_1614);
nand U4418 (N_4418,N_485,N_1241);
nor U4419 (N_4419,N_2658,N_1729);
nor U4420 (N_4420,N_2470,N_2378);
nor U4421 (N_4421,N_1502,N_1523);
nand U4422 (N_4422,N_1193,N_729);
or U4423 (N_4423,N_600,N_1899);
or U4424 (N_4424,N_2731,N_2783);
and U4425 (N_4425,N_2666,N_606);
nand U4426 (N_4426,N_1354,N_2037);
and U4427 (N_4427,N_1040,N_263);
xnor U4428 (N_4428,N_509,N_2439);
and U4429 (N_4429,N_993,N_133);
and U4430 (N_4430,N_2161,N_628);
nor U4431 (N_4431,N_2076,N_75);
nand U4432 (N_4432,N_1351,N_3044);
and U4433 (N_4433,N_855,N_647);
or U4434 (N_4434,N_1398,N_290);
nand U4435 (N_4435,N_2262,N_372);
and U4436 (N_4436,N_657,N_2303);
nand U4437 (N_4437,N_698,N_137);
and U4438 (N_4438,N_320,N_3013);
nor U4439 (N_4439,N_1139,N_1993);
nor U4440 (N_4440,N_1000,N_1057);
nor U4441 (N_4441,N_1228,N_946);
nand U4442 (N_4442,N_295,N_940);
nor U4443 (N_4443,N_970,N_2759);
and U4444 (N_4444,N_1970,N_803);
or U4445 (N_4445,N_2633,N_1802);
and U4446 (N_4446,N_675,N_715);
or U4447 (N_4447,N_948,N_164);
xor U4448 (N_4448,N_846,N_53);
and U4449 (N_4449,N_54,N_2214);
nor U4450 (N_4450,N_681,N_2767);
nor U4451 (N_4451,N_2349,N_1756);
or U4452 (N_4452,N_1238,N_2122);
or U4453 (N_4453,N_1381,N_546);
or U4454 (N_4454,N_1323,N_1457);
nor U4455 (N_4455,N_2151,N_1732);
and U4456 (N_4456,N_3103,N_904);
nand U4457 (N_4457,N_2454,N_1452);
nor U4458 (N_4458,N_1166,N_23);
and U4459 (N_4459,N_2311,N_2862);
nand U4460 (N_4460,N_2827,N_105);
nand U4461 (N_4461,N_2592,N_1144);
or U4462 (N_4462,N_2317,N_1750);
nor U4463 (N_4463,N_41,N_2992);
nor U4464 (N_4464,N_1784,N_431);
or U4465 (N_4465,N_1322,N_1171);
or U4466 (N_4466,N_1500,N_2732);
or U4467 (N_4467,N_894,N_1967);
xnor U4468 (N_4468,N_1393,N_1116);
or U4469 (N_4469,N_468,N_3091);
nand U4470 (N_4470,N_1492,N_2852);
or U4471 (N_4471,N_1369,N_2676);
nand U4472 (N_4472,N_1702,N_484);
and U4473 (N_4473,N_1924,N_1513);
and U4474 (N_4474,N_2539,N_1958);
nor U4475 (N_4475,N_2057,N_1227);
nor U4476 (N_4476,N_838,N_2810);
xor U4477 (N_4477,N_373,N_1850);
nor U4478 (N_4478,N_2855,N_12);
and U4479 (N_4479,N_365,N_1611);
nand U4480 (N_4480,N_2957,N_1772);
or U4481 (N_4481,N_635,N_1982);
and U4482 (N_4482,N_219,N_906);
nand U4483 (N_4483,N_2384,N_3063);
or U4484 (N_4484,N_1593,N_1361);
xnor U4485 (N_4485,N_831,N_749);
nand U4486 (N_4486,N_473,N_1598);
or U4487 (N_4487,N_870,N_1396);
nor U4488 (N_4488,N_2013,N_1092);
nand U4489 (N_4489,N_2044,N_1146);
or U4490 (N_4490,N_2200,N_2925);
and U4491 (N_4491,N_180,N_1656);
nand U4492 (N_4492,N_61,N_121);
nor U4493 (N_4493,N_2323,N_2388);
nor U4494 (N_4494,N_1156,N_2626);
nor U4495 (N_4495,N_2028,N_374);
nand U4496 (N_4496,N_943,N_1725);
or U4497 (N_4497,N_2650,N_1479);
and U4498 (N_4498,N_2559,N_2473);
xor U4499 (N_4499,N_2561,N_1636);
nor U4500 (N_4500,N_1173,N_1487);
xnor U4501 (N_4501,N_1609,N_1667);
nor U4502 (N_4502,N_589,N_1815);
xnor U4503 (N_4503,N_2318,N_1247);
xor U4504 (N_4504,N_1497,N_908);
nand U4505 (N_4505,N_2863,N_840);
and U4506 (N_4506,N_874,N_556);
xor U4507 (N_4507,N_3092,N_2786);
or U4508 (N_4508,N_738,N_1711);
xnor U4509 (N_4509,N_1270,N_2530);
and U4510 (N_4510,N_808,N_3074);
nand U4511 (N_4511,N_1786,N_1836);
nor U4512 (N_4512,N_2667,N_1355);
nand U4513 (N_4513,N_1841,N_2644);
xor U4514 (N_4514,N_2116,N_1805);
nand U4515 (N_4515,N_3,N_2024);
or U4516 (N_4516,N_2989,N_3099);
nand U4517 (N_4517,N_634,N_804);
xor U4518 (N_4518,N_1855,N_1195);
and U4519 (N_4519,N_2800,N_233);
or U4520 (N_4520,N_1496,N_1163);
xnor U4521 (N_4521,N_1088,N_1380);
nor U4522 (N_4522,N_2583,N_2642);
nor U4523 (N_4523,N_2033,N_791);
and U4524 (N_4524,N_768,N_2604);
nor U4525 (N_4525,N_2198,N_650);
or U4526 (N_4526,N_323,N_620);
or U4527 (N_4527,N_2685,N_2293);
nor U4528 (N_4528,N_735,N_1079);
or U4529 (N_4529,N_1311,N_526);
and U4530 (N_4530,N_100,N_1142);
or U4531 (N_4531,N_2165,N_885);
xor U4532 (N_4532,N_626,N_3089);
nor U4533 (N_4533,N_1059,N_580);
and U4534 (N_4534,N_1310,N_2734);
and U4535 (N_4535,N_1662,N_2423);
or U4536 (N_4536,N_2012,N_2149);
or U4537 (N_4537,N_1582,N_548);
nand U4538 (N_4538,N_680,N_1483);
and U4539 (N_4539,N_206,N_2166);
and U4540 (N_4540,N_1837,N_1313);
nor U4541 (N_4541,N_3086,N_1831);
nor U4542 (N_4542,N_1056,N_449);
nand U4543 (N_4543,N_355,N_3119);
or U4544 (N_4544,N_793,N_1792);
nand U4545 (N_4545,N_2901,N_2430);
or U4546 (N_4546,N_65,N_463);
or U4547 (N_4547,N_1333,N_247);
or U4548 (N_4548,N_1066,N_1188);
or U4549 (N_4549,N_1749,N_1179);
nand U4550 (N_4550,N_407,N_1653);
or U4551 (N_4551,N_510,N_1331);
nand U4552 (N_4552,N_930,N_716);
and U4553 (N_4553,N_319,N_2268);
or U4554 (N_4554,N_116,N_1182);
or U4555 (N_4555,N_896,N_767);
nand U4556 (N_4556,N_2641,N_1790);
nand U4557 (N_4557,N_1052,N_533);
nor U4558 (N_4558,N_2804,N_2019);
or U4559 (N_4559,N_899,N_134);
nor U4560 (N_4560,N_566,N_850);
nor U4561 (N_4561,N_2892,N_2725);
nor U4562 (N_4562,N_1606,N_1014);
nand U4563 (N_4563,N_1706,N_2449);
nor U4564 (N_4564,N_2926,N_1135);
or U4565 (N_4565,N_1930,N_1001);
and U4566 (N_4566,N_1412,N_375);
xnor U4567 (N_4567,N_2668,N_2817);
or U4568 (N_4568,N_29,N_1436);
nand U4569 (N_4569,N_2060,N_1277);
and U4570 (N_4570,N_999,N_3093);
nor U4571 (N_4571,N_590,N_2395);
and U4572 (N_4572,N_2355,N_2848);
xnor U4573 (N_4573,N_1751,N_292);
xor U4574 (N_4574,N_62,N_2537);
nor U4575 (N_4575,N_2495,N_739);
or U4576 (N_4576,N_2541,N_1548);
nand U4577 (N_4577,N_2339,N_170);
or U4578 (N_4578,N_888,N_3039);
and U4579 (N_4579,N_1963,N_2083);
nand U4580 (N_4580,N_947,N_1778);
nor U4581 (N_4581,N_969,N_757);
and U4582 (N_4582,N_1278,N_2001);
or U4583 (N_4583,N_1689,N_877);
nand U4584 (N_4584,N_2629,N_1498);
nand U4585 (N_4585,N_1218,N_174);
xor U4586 (N_4586,N_1078,N_2282);
nand U4587 (N_4587,N_2948,N_122);
nor U4588 (N_4588,N_575,N_1555);
or U4589 (N_4589,N_880,N_2747);
or U4590 (N_4590,N_1183,N_441);
or U4591 (N_4591,N_305,N_1090);
nor U4592 (N_4592,N_1691,N_2158);
or U4593 (N_4593,N_2302,N_2596);
or U4594 (N_4594,N_1793,N_282);
nor U4595 (N_4595,N_1832,N_805);
and U4596 (N_4596,N_81,N_2976);
nand U4597 (N_4597,N_3102,N_2407);
nand U4598 (N_4598,N_2042,N_2770);
nor U4599 (N_4599,N_2934,N_2246);
nand U4600 (N_4600,N_1162,N_2099);
nand U4601 (N_4601,N_1155,N_660);
and U4602 (N_4602,N_1184,N_314);
nand U4603 (N_4603,N_2915,N_1908);
xnor U4604 (N_4604,N_177,N_115);
nor U4605 (N_4605,N_1536,N_357);
and U4606 (N_4606,N_2338,N_1937);
or U4607 (N_4607,N_865,N_2984);
nor U4608 (N_4608,N_779,N_2197);
nor U4609 (N_4609,N_2350,N_2573);
xnor U4610 (N_4610,N_467,N_1411);
nor U4611 (N_4611,N_1980,N_1064);
nor U4612 (N_4612,N_294,N_1374);
and U4613 (N_4613,N_2089,N_631);
xnor U4614 (N_4614,N_1346,N_2485);
nand U4615 (N_4615,N_694,N_2681);
xnor U4616 (N_4616,N_978,N_2409);
and U4617 (N_4617,N_423,N_2966);
nor U4618 (N_4618,N_2822,N_2448);
and U4619 (N_4619,N_2715,N_1082);
nor U4620 (N_4620,N_2843,N_1686);
or U4621 (N_4621,N_2849,N_925);
nor U4622 (N_4622,N_2660,N_2330);
or U4623 (N_4623,N_2696,N_257);
or U4624 (N_4624,N_1420,N_1019);
xnor U4625 (N_4625,N_2316,N_1032);
nor U4626 (N_4626,N_1491,N_8);
or U4627 (N_4627,N_2693,N_504);
nand U4628 (N_4628,N_2201,N_2085);
and U4629 (N_4629,N_2719,N_236);
nand U4630 (N_4630,N_1104,N_922);
xnor U4631 (N_4631,N_1409,N_2972);
nand U4632 (N_4632,N_3043,N_2945);
and U4633 (N_4633,N_1752,N_921);
nand U4634 (N_4634,N_3041,N_639);
or U4635 (N_4635,N_2117,N_1628);
nand U4636 (N_4636,N_980,N_1777);
xor U4637 (N_4637,N_579,N_1819);
and U4638 (N_4638,N_1903,N_2194);
nand U4639 (N_4639,N_1508,N_820);
xnor U4640 (N_4640,N_892,N_3076);
nand U4641 (N_4641,N_2424,N_1959);
or U4642 (N_4642,N_1942,N_205);
and U4643 (N_4643,N_527,N_2652);
or U4644 (N_4644,N_1613,N_47);
or U4645 (N_4645,N_1264,N_968);
or U4646 (N_4646,N_2509,N_1376);
xnor U4647 (N_4647,N_2143,N_710);
nand U4648 (N_4648,N_522,N_3065);
nor U4649 (N_4649,N_684,N_2052);
nand U4650 (N_4650,N_2716,N_2869);
nor U4651 (N_4651,N_2319,N_3040);
or U4652 (N_4652,N_780,N_2518);
and U4653 (N_4653,N_2072,N_2529);
and U4654 (N_4654,N_2139,N_309);
nand U4655 (N_4655,N_2332,N_2446);
nor U4656 (N_4656,N_307,N_345);
nand U4657 (N_4657,N_1704,N_2308);
or U4658 (N_4658,N_44,N_2801);
nand U4659 (N_4659,N_2150,N_2475);
or U4660 (N_4660,N_668,N_1650);
or U4661 (N_4661,N_1248,N_1882);
nor U4662 (N_4662,N_506,N_2730);
and U4663 (N_4663,N_2352,N_2684);
nor U4664 (N_4664,N_492,N_1557);
nor U4665 (N_4665,N_2411,N_455);
nor U4666 (N_4666,N_349,N_1859);
and U4667 (N_4667,N_2091,N_1901);
nor U4668 (N_4668,N_1360,N_1099);
nor U4669 (N_4669,N_1579,N_173);
nand U4670 (N_4670,N_557,N_1692);
nor U4671 (N_4671,N_1049,N_1782);
nor U4672 (N_4672,N_312,N_331);
and U4673 (N_4673,N_521,N_813);
xnor U4674 (N_4674,N_258,N_614);
nor U4675 (N_4675,N_1036,N_317);
nor U4676 (N_4676,N_2334,N_1843);
nand U4677 (N_4677,N_343,N_2026);
nor U4678 (N_4678,N_599,N_2036);
xnor U4679 (N_4679,N_2634,N_1645);
or U4680 (N_4680,N_2516,N_3019);
nand U4681 (N_4681,N_1391,N_2265);
or U4682 (N_4682,N_303,N_2998);
nand U4683 (N_4683,N_552,N_1867);
nand U4684 (N_4684,N_2247,N_2432);
nand U4685 (N_4685,N_1552,N_722);
xor U4686 (N_4686,N_2960,N_1265);
or U4687 (N_4687,N_598,N_2405);
xnor U4688 (N_4688,N_1281,N_1580);
and U4689 (N_4689,N_1790,N_2655);
nor U4690 (N_4690,N_2683,N_794);
nor U4691 (N_4691,N_733,N_947);
and U4692 (N_4692,N_2845,N_2103);
nand U4693 (N_4693,N_2920,N_2984);
xnor U4694 (N_4694,N_1967,N_3103);
nand U4695 (N_4695,N_822,N_1673);
or U4696 (N_4696,N_482,N_2217);
xnor U4697 (N_4697,N_2353,N_2530);
or U4698 (N_4698,N_2283,N_2694);
nor U4699 (N_4699,N_2360,N_917);
nand U4700 (N_4700,N_266,N_267);
and U4701 (N_4701,N_3078,N_2055);
nor U4702 (N_4702,N_202,N_288);
or U4703 (N_4703,N_2899,N_243);
xnor U4704 (N_4704,N_2641,N_1594);
nand U4705 (N_4705,N_2251,N_1524);
nand U4706 (N_4706,N_1738,N_365);
and U4707 (N_4707,N_1189,N_748);
or U4708 (N_4708,N_1645,N_520);
and U4709 (N_4709,N_2744,N_1162);
nand U4710 (N_4710,N_767,N_1480);
and U4711 (N_4711,N_952,N_995);
or U4712 (N_4712,N_1721,N_2317);
or U4713 (N_4713,N_1068,N_2054);
or U4714 (N_4714,N_142,N_2348);
nor U4715 (N_4715,N_790,N_1410);
nor U4716 (N_4716,N_142,N_2964);
and U4717 (N_4717,N_2423,N_3071);
nor U4718 (N_4718,N_2500,N_1329);
and U4719 (N_4719,N_589,N_1254);
nand U4720 (N_4720,N_2946,N_2709);
or U4721 (N_4721,N_2692,N_2753);
xnor U4722 (N_4722,N_980,N_3007);
nand U4723 (N_4723,N_226,N_1422);
nor U4724 (N_4724,N_935,N_2957);
nor U4725 (N_4725,N_853,N_2417);
nand U4726 (N_4726,N_2225,N_384);
or U4727 (N_4727,N_3024,N_2115);
nor U4728 (N_4728,N_1060,N_592);
and U4729 (N_4729,N_11,N_236);
or U4730 (N_4730,N_1936,N_2584);
or U4731 (N_4731,N_2634,N_2529);
nand U4732 (N_4732,N_168,N_2849);
nor U4733 (N_4733,N_237,N_990);
and U4734 (N_4734,N_1817,N_877);
and U4735 (N_4735,N_19,N_2061);
and U4736 (N_4736,N_3055,N_980);
nor U4737 (N_4737,N_454,N_1476);
nor U4738 (N_4738,N_1812,N_3121);
nor U4739 (N_4739,N_2783,N_623);
or U4740 (N_4740,N_1528,N_2811);
or U4741 (N_4741,N_1270,N_428);
or U4742 (N_4742,N_170,N_1452);
nand U4743 (N_4743,N_816,N_2918);
nor U4744 (N_4744,N_971,N_2152);
and U4745 (N_4745,N_171,N_534);
and U4746 (N_4746,N_274,N_1346);
and U4747 (N_4747,N_2420,N_2653);
xnor U4748 (N_4748,N_2104,N_2709);
or U4749 (N_4749,N_1420,N_1360);
nand U4750 (N_4750,N_1004,N_2375);
nand U4751 (N_4751,N_751,N_2133);
and U4752 (N_4752,N_1353,N_304);
and U4753 (N_4753,N_2135,N_1982);
and U4754 (N_4754,N_1914,N_726);
xor U4755 (N_4755,N_1975,N_931);
and U4756 (N_4756,N_1733,N_2571);
or U4757 (N_4757,N_3060,N_1199);
or U4758 (N_4758,N_2967,N_2842);
or U4759 (N_4759,N_1456,N_182);
or U4760 (N_4760,N_1004,N_2507);
nand U4761 (N_4761,N_2780,N_3109);
nor U4762 (N_4762,N_2291,N_2854);
nand U4763 (N_4763,N_2835,N_2305);
nor U4764 (N_4764,N_2993,N_612);
nand U4765 (N_4765,N_2163,N_645);
and U4766 (N_4766,N_2231,N_2078);
xnor U4767 (N_4767,N_2933,N_563);
nor U4768 (N_4768,N_1637,N_2855);
or U4769 (N_4769,N_408,N_1366);
and U4770 (N_4770,N_342,N_1112);
nand U4771 (N_4771,N_1762,N_2745);
or U4772 (N_4772,N_2638,N_2036);
or U4773 (N_4773,N_1187,N_2702);
or U4774 (N_4774,N_2623,N_1555);
nor U4775 (N_4775,N_1286,N_690);
and U4776 (N_4776,N_2492,N_2977);
and U4777 (N_4777,N_1430,N_1478);
nand U4778 (N_4778,N_550,N_1016);
or U4779 (N_4779,N_114,N_2495);
or U4780 (N_4780,N_1609,N_2529);
and U4781 (N_4781,N_149,N_1990);
and U4782 (N_4782,N_500,N_398);
nand U4783 (N_4783,N_645,N_262);
and U4784 (N_4784,N_2428,N_587);
nor U4785 (N_4785,N_2382,N_2717);
xnor U4786 (N_4786,N_2732,N_400);
or U4787 (N_4787,N_1053,N_2608);
nand U4788 (N_4788,N_2897,N_709);
xor U4789 (N_4789,N_678,N_83);
or U4790 (N_4790,N_1805,N_1030);
nand U4791 (N_4791,N_1883,N_2591);
or U4792 (N_4792,N_305,N_1169);
nor U4793 (N_4793,N_1140,N_1563);
nand U4794 (N_4794,N_1573,N_1535);
nand U4795 (N_4795,N_2629,N_607);
or U4796 (N_4796,N_943,N_3096);
or U4797 (N_4797,N_2385,N_1640);
nand U4798 (N_4798,N_862,N_286);
nor U4799 (N_4799,N_1352,N_860);
nor U4800 (N_4800,N_2718,N_2608);
and U4801 (N_4801,N_1774,N_1968);
and U4802 (N_4802,N_2072,N_746);
and U4803 (N_4803,N_2704,N_1563);
nor U4804 (N_4804,N_1417,N_1301);
nor U4805 (N_4805,N_2013,N_1493);
or U4806 (N_4806,N_1974,N_312);
or U4807 (N_4807,N_1483,N_1924);
nand U4808 (N_4808,N_1643,N_1942);
xor U4809 (N_4809,N_48,N_1634);
nand U4810 (N_4810,N_1188,N_1959);
nor U4811 (N_4811,N_1294,N_1819);
nand U4812 (N_4812,N_2579,N_2164);
nand U4813 (N_4813,N_261,N_1137);
or U4814 (N_4814,N_2060,N_2933);
nor U4815 (N_4815,N_1542,N_378);
or U4816 (N_4816,N_2411,N_2085);
or U4817 (N_4817,N_2154,N_1847);
xor U4818 (N_4818,N_2019,N_492);
nand U4819 (N_4819,N_1832,N_22);
nand U4820 (N_4820,N_1648,N_2904);
nand U4821 (N_4821,N_1927,N_2030);
and U4822 (N_4822,N_1299,N_1725);
and U4823 (N_4823,N_360,N_761);
xnor U4824 (N_4824,N_372,N_235);
nand U4825 (N_4825,N_383,N_2287);
or U4826 (N_4826,N_1139,N_2144);
nand U4827 (N_4827,N_126,N_113);
or U4828 (N_4828,N_1092,N_279);
and U4829 (N_4829,N_349,N_41);
nor U4830 (N_4830,N_860,N_710);
nand U4831 (N_4831,N_1332,N_1335);
or U4832 (N_4832,N_1576,N_1478);
and U4833 (N_4833,N_887,N_2886);
nor U4834 (N_4834,N_1248,N_76);
and U4835 (N_4835,N_510,N_1416);
or U4836 (N_4836,N_174,N_1906);
or U4837 (N_4837,N_2081,N_1270);
and U4838 (N_4838,N_1285,N_2842);
and U4839 (N_4839,N_2274,N_2926);
nor U4840 (N_4840,N_1306,N_501);
or U4841 (N_4841,N_545,N_3082);
and U4842 (N_4842,N_859,N_2958);
or U4843 (N_4843,N_417,N_1769);
and U4844 (N_4844,N_2064,N_854);
xor U4845 (N_4845,N_2955,N_1424);
nand U4846 (N_4846,N_1419,N_869);
xnor U4847 (N_4847,N_73,N_2391);
nor U4848 (N_4848,N_306,N_995);
nand U4849 (N_4849,N_2362,N_3080);
nand U4850 (N_4850,N_2606,N_2366);
and U4851 (N_4851,N_2801,N_1060);
nor U4852 (N_4852,N_2307,N_2168);
and U4853 (N_4853,N_2772,N_1321);
or U4854 (N_4854,N_2664,N_1920);
and U4855 (N_4855,N_2506,N_109);
and U4856 (N_4856,N_2335,N_1728);
or U4857 (N_4857,N_163,N_2670);
nor U4858 (N_4858,N_2437,N_1890);
and U4859 (N_4859,N_2372,N_211);
or U4860 (N_4860,N_338,N_3006);
nand U4861 (N_4861,N_2762,N_1226);
and U4862 (N_4862,N_2655,N_2325);
or U4863 (N_4863,N_757,N_1347);
and U4864 (N_4864,N_462,N_1488);
nor U4865 (N_4865,N_3102,N_2735);
and U4866 (N_4866,N_3081,N_1104);
nand U4867 (N_4867,N_3026,N_2393);
nor U4868 (N_4868,N_1682,N_1435);
and U4869 (N_4869,N_2896,N_2026);
and U4870 (N_4870,N_1872,N_761);
xnor U4871 (N_4871,N_2096,N_2411);
and U4872 (N_4872,N_2861,N_912);
and U4873 (N_4873,N_221,N_2983);
xor U4874 (N_4874,N_207,N_514);
and U4875 (N_4875,N_558,N_2248);
nand U4876 (N_4876,N_2053,N_1887);
nor U4877 (N_4877,N_984,N_1521);
or U4878 (N_4878,N_2074,N_2764);
or U4879 (N_4879,N_2446,N_1030);
and U4880 (N_4880,N_2024,N_622);
nand U4881 (N_4881,N_2527,N_742);
nor U4882 (N_4882,N_2269,N_1674);
nand U4883 (N_4883,N_1066,N_1453);
and U4884 (N_4884,N_1906,N_1548);
nand U4885 (N_4885,N_2981,N_733);
nand U4886 (N_4886,N_575,N_2272);
and U4887 (N_4887,N_1481,N_1480);
xor U4888 (N_4888,N_1256,N_1476);
nand U4889 (N_4889,N_2065,N_1460);
nand U4890 (N_4890,N_426,N_2662);
and U4891 (N_4891,N_1082,N_1975);
nand U4892 (N_4892,N_452,N_923);
xor U4893 (N_4893,N_633,N_1516);
nor U4894 (N_4894,N_1031,N_2542);
xnor U4895 (N_4895,N_1367,N_2311);
nor U4896 (N_4896,N_2523,N_2899);
nor U4897 (N_4897,N_1786,N_468);
nand U4898 (N_4898,N_2143,N_2701);
or U4899 (N_4899,N_816,N_1300);
xor U4900 (N_4900,N_2223,N_2313);
and U4901 (N_4901,N_2620,N_586);
or U4902 (N_4902,N_2892,N_2510);
and U4903 (N_4903,N_1655,N_2966);
nand U4904 (N_4904,N_2415,N_2963);
nor U4905 (N_4905,N_1727,N_1219);
nand U4906 (N_4906,N_803,N_2786);
nor U4907 (N_4907,N_1172,N_766);
xor U4908 (N_4908,N_3101,N_2212);
nand U4909 (N_4909,N_1112,N_1183);
or U4910 (N_4910,N_2287,N_2042);
nor U4911 (N_4911,N_1889,N_1461);
nor U4912 (N_4912,N_2737,N_2118);
nand U4913 (N_4913,N_1327,N_110);
nand U4914 (N_4914,N_2735,N_1606);
nor U4915 (N_4915,N_2365,N_2544);
nand U4916 (N_4916,N_2959,N_2997);
nor U4917 (N_4917,N_597,N_739);
or U4918 (N_4918,N_789,N_2542);
xor U4919 (N_4919,N_1326,N_1456);
or U4920 (N_4920,N_113,N_2996);
and U4921 (N_4921,N_1400,N_700);
nand U4922 (N_4922,N_590,N_2727);
nand U4923 (N_4923,N_1467,N_2486);
and U4924 (N_4924,N_1433,N_2789);
nand U4925 (N_4925,N_1522,N_1181);
and U4926 (N_4926,N_1140,N_11);
and U4927 (N_4927,N_3013,N_891);
nor U4928 (N_4928,N_918,N_1304);
nand U4929 (N_4929,N_2392,N_2709);
and U4930 (N_4930,N_798,N_1825);
nand U4931 (N_4931,N_1378,N_2827);
nor U4932 (N_4932,N_2610,N_2751);
nor U4933 (N_4933,N_396,N_104);
and U4934 (N_4934,N_561,N_1308);
xor U4935 (N_4935,N_2963,N_791);
xnor U4936 (N_4936,N_1260,N_324);
and U4937 (N_4937,N_2452,N_2584);
xor U4938 (N_4938,N_2032,N_617);
and U4939 (N_4939,N_410,N_663);
or U4940 (N_4940,N_1755,N_2589);
or U4941 (N_4941,N_2610,N_1144);
and U4942 (N_4942,N_2064,N_1475);
and U4943 (N_4943,N_866,N_1522);
and U4944 (N_4944,N_2265,N_223);
or U4945 (N_4945,N_814,N_2928);
and U4946 (N_4946,N_2531,N_2083);
nor U4947 (N_4947,N_205,N_537);
and U4948 (N_4948,N_967,N_2874);
xnor U4949 (N_4949,N_2003,N_324);
and U4950 (N_4950,N_646,N_1503);
xnor U4951 (N_4951,N_615,N_705);
nor U4952 (N_4952,N_374,N_445);
or U4953 (N_4953,N_2348,N_812);
nand U4954 (N_4954,N_1384,N_1363);
or U4955 (N_4955,N_2659,N_2877);
or U4956 (N_4956,N_2361,N_2064);
or U4957 (N_4957,N_1488,N_1038);
nand U4958 (N_4958,N_3073,N_2471);
or U4959 (N_4959,N_965,N_2585);
nor U4960 (N_4960,N_302,N_1079);
or U4961 (N_4961,N_2811,N_3062);
nand U4962 (N_4962,N_580,N_2103);
nor U4963 (N_4963,N_1186,N_961);
and U4964 (N_4964,N_2055,N_330);
or U4965 (N_4965,N_528,N_1501);
nor U4966 (N_4966,N_236,N_1977);
nand U4967 (N_4967,N_2323,N_1301);
nor U4968 (N_4968,N_697,N_1758);
or U4969 (N_4969,N_36,N_551);
xor U4970 (N_4970,N_186,N_1991);
nor U4971 (N_4971,N_753,N_1494);
and U4972 (N_4972,N_1123,N_1003);
or U4973 (N_4973,N_183,N_3089);
nand U4974 (N_4974,N_1471,N_2589);
nand U4975 (N_4975,N_2923,N_2843);
or U4976 (N_4976,N_278,N_953);
nand U4977 (N_4977,N_434,N_580);
nor U4978 (N_4978,N_63,N_1409);
and U4979 (N_4979,N_1387,N_341);
or U4980 (N_4980,N_907,N_1547);
and U4981 (N_4981,N_593,N_117);
or U4982 (N_4982,N_2700,N_2396);
or U4983 (N_4983,N_604,N_2689);
nand U4984 (N_4984,N_1303,N_1570);
and U4985 (N_4985,N_1455,N_2034);
nor U4986 (N_4986,N_1096,N_1247);
nor U4987 (N_4987,N_882,N_2978);
xor U4988 (N_4988,N_475,N_1048);
nand U4989 (N_4989,N_744,N_2489);
and U4990 (N_4990,N_1063,N_1304);
nand U4991 (N_4991,N_750,N_2029);
nor U4992 (N_4992,N_2008,N_2140);
and U4993 (N_4993,N_1420,N_306);
nor U4994 (N_4994,N_161,N_1400);
nor U4995 (N_4995,N_1630,N_882);
nand U4996 (N_4996,N_3011,N_2026);
and U4997 (N_4997,N_1725,N_1228);
nor U4998 (N_4998,N_2686,N_2558);
and U4999 (N_4999,N_205,N_697);
nor U5000 (N_5000,N_555,N_362);
and U5001 (N_5001,N_1851,N_1937);
or U5002 (N_5002,N_406,N_2491);
or U5003 (N_5003,N_1615,N_792);
nand U5004 (N_5004,N_1373,N_835);
and U5005 (N_5005,N_340,N_2667);
xnor U5006 (N_5006,N_108,N_2032);
and U5007 (N_5007,N_2205,N_2281);
or U5008 (N_5008,N_2611,N_967);
xnor U5009 (N_5009,N_2558,N_49);
xor U5010 (N_5010,N_2062,N_560);
nand U5011 (N_5011,N_945,N_887);
and U5012 (N_5012,N_2436,N_1139);
and U5013 (N_5013,N_2351,N_1610);
nor U5014 (N_5014,N_58,N_79);
nor U5015 (N_5015,N_9,N_2868);
nand U5016 (N_5016,N_1980,N_1368);
nor U5017 (N_5017,N_1396,N_1079);
or U5018 (N_5018,N_1545,N_1759);
nor U5019 (N_5019,N_2807,N_716);
nor U5020 (N_5020,N_2512,N_113);
nor U5021 (N_5021,N_2167,N_2934);
or U5022 (N_5022,N_1674,N_2276);
nand U5023 (N_5023,N_1429,N_1453);
nand U5024 (N_5024,N_758,N_3028);
and U5025 (N_5025,N_1470,N_728);
or U5026 (N_5026,N_3008,N_456);
xnor U5027 (N_5027,N_12,N_942);
or U5028 (N_5028,N_689,N_374);
xor U5029 (N_5029,N_1413,N_1833);
and U5030 (N_5030,N_456,N_324);
nand U5031 (N_5031,N_809,N_2787);
and U5032 (N_5032,N_673,N_1070);
nor U5033 (N_5033,N_2330,N_621);
nor U5034 (N_5034,N_434,N_2937);
or U5035 (N_5035,N_1806,N_497);
xor U5036 (N_5036,N_923,N_2500);
xor U5037 (N_5037,N_1097,N_1831);
nor U5038 (N_5038,N_1155,N_594);
nor U5039 (N_5039,N_2553,N_8);
nor U5040 (N_5040,N_1568,N_2093);
or U5041 (N_5041,N_55,N_2838);
xor U5042 (N_5042,N_731,N_1561);
nor U5043 (N_5043,N_1279,N_2555);
and U5044 (N_5044,N_1926,N_644);
or U5045 (N_5045,N_2245,N_1000);
nand U5046 (N_5046,N_1596,N_638);
or U5047 (N_5047,N_814,N_640);
and U5048 (N_5048,N_2183,N_202);
and U5049 (N_5049,N_1721,N_2085);
or U5050 (N_5050,N_1780,N_2378);
nor U5051 (N_5051,N_1788,N_149);
or U5052 (N_5052,N_1978,N_2909);
or U5053 (N_5053,N_2039,N_1709);
nor U5054 (N_5054,N_2894,N_744);
or U5055 (N_5055,N_1048,N_1521);
xor U5056 (N_5056,N_1492,N_2167);
nand U5057 (N_5057,N_340,N_2653);
nand U5058 (N_5058,N_2293,N_2611);
or U5059 (N_5059,N_1691,N_1985);
nor U5060 (N_5060,N_1632,N_1683);
and U5061 (N_5061,N_1576,N_2756);
nor U5062 (N_5062,N_1087,N_482);
or U5063 (N_5063,N_1128,N_2321);
or U5064 (N_5064,N_264,N_2357);
nand U5065 (N_5065,N_561,N_1118);
nand U5066 (N_5066,N_947,N_2240);
nand U5067 (N_5067,N_3110,N_1506);
xnor U5068 (N_5068,N_2215,N_1627);
nand U5069 (N_5069,N_1268,N_1421);
or U5070 (N_5070,N_489,N_2506);
and U5071 (N_5071,N_1460,N_438);
and U5072 (N_5072,N_2813,N_739);
or U5073 (N_5073,N_1842,N_1647);
and U5074 (N_5074,N_871,N_595);
xor U5075 (N_5075,N_1213,N_492);
nor U5076 (N_5076,N_600,N_2103);
nor U5077 (N_5077,N_805,N_2434);
and U5078 (N_5078,N_1162,N_2871);
and U5079 (N_5079,N_1571,N_1579);
nor U5080 (N_5080,N_2618,N_769);
xnor U5081 (N_5081,N_1644,N_1978);
or U5082 (N_5082,N_843,N_3053);
nand U5083 (N_5083,N_2210,N_1603);
nand U5084 (N_5084,N_2661,N_1589);
xnor U5085 (N_5085,N_3062,N_2047);
xnor U5086 (N_5086,N_1962,N_1189);
and U5087 (N_5087,N_1110,N_2024);
or U5088 (N_5088,N_2581,N_41);
xnor U5089 (N_5089,N_1447,N_2796);
nand U5090 (N_5090,N_86,N_737);
and U5091 (N_5091,N_740,N_2658);
xor U5092 (N_5092,N_1159,N_3085);
nor U5093 (N_5093,N_1056,N_1766);
nand U5094 (N_5094,N_2600,N_2978);
and U5095 (N_5095,N_394,N_1905);
or U5096 (N_5096,N_330,N_857);
nor U5097 (N_5097,N_2856,N_788);
nand U5098 (N_5098,N_1587,N_999);
xnor U5099 (N_5099,N_1270,N_215);
nand U5100 (N_5100,N_2178,N_3013);
nor U5101 (N_5101,N_1606,N_2750);
xor U5102 (N_5102,N_1305,N_2381);
or U5103 (N_5103,N_1089,N_1199);
and U5104 (N_5104,N_1826,N_956);
nand U5105 (N_5105,N_2412,N_385);
nand U5106 (N_5106,N_2757,N_2704);
or U5107 (N_5107,N_1914,N_1063);
xor U5108 (N_5108,N_1097,N_2296);
or U5109 (N_5109,N_1138,N_1792);
or U5110 (N_5110,N_1461,N_1207);
nand U5111 (N_5111,N_2783,N_3035);
and U5112 (N_5112,N_103,N_1266);
and U5113 (N_5113,N_737,N_2393);
nand U5114 (N_5114,N_1518,N_54);
and U5115 (N_5115,N_477,N_2968);
and U5116 (N_5116,N_168,N_2809);
and U5117 (N_5117,N_1437,N_567);
nor U5118 (N_5118,N_2848,N_1166);
nor U5119 (N_5119,N_114,N_130);
nand U5120 (N_5120,N_2633,N_1092);
nand U5121 (N_5121,N_2997,N_536);
or U5122 (N_5122,N_1865,N_2935);
nor U5123 (N_5123,N_1894,N_751);
and U5124 (N_5124,N_1519,N_896);
or U5125 (N_5125,N_2656,N_2738);
nor U5126 (N_5126,N_1430,N_626);
nand U5127 (N_5127,N_2380,N_1945);
and U5128 (N_5128,N_1336,N_2744);
and U5129 (N_5129,N_2291,N_1618);
and U5130 (N_5130,N_2575,N_1451);
nand U5131 (N_5131,N_1294,N_74);
nand U5132 (N_5132,N_1466,N_1474);
nor U5133 (N_5133,N_509,N_1946);
or U5134 (N_5134,N_1527,N_2712);
nor U5135 (N_5135,N_1535,N_902);
and U5136 (N_5136,N_379,N_1398);
xor U5137 (N_5137,N_1942,N_2169);
and U5138 (N_5138,N_2202,N_1183);
or U5139 (N_5139,N_2888,N_652);
and U5140 (N_5140,N_1783,N_1430);
nor U5141 (N_5141,N_456,N_2610);
nor U5142 (N_5142,N_2997,N_2910);
nor U5143 (N_5143,N_1082,N_1398);
nor U5144 (N_5144,N_337,N_984);
and U5145 (N_5145,N_416,N_1077);
xor U5146 (N_5146,N_2248,N_1423);
xor U5147 (N_5147,N_2464,N_132);
xor U5148 (N_5148,N_2924,N_2029);
and U5149 (N_5149,N_2334,N_2876);
and U5150 (N_5150,N_2276,N_1691);
and U5151 (N_5151,N_3019,N_695);
and U5152 (N_5152,N_176,N_2912);
nor U5153 (N_5153,N_2609,N_225);
and U5154 (N_5154,N_2623,N_380);
nand U5155 (N_5155,N_1530,N_228);
nor U5156 (N_5156,N_1664,N_3023);
nand U5157 (N_5157,N_2800,N_1013);
nor U5158 (N_5158,N_1036,N_2764);
xor U5159 (N_5159,N_477,N_2885);
nand U5160 (N_5160,N_166,N_927);
or U5161 (N_5161,N_991,N_2227);
or U5162 (N_5162,N_1361,N_2532);
or U5163 (N_5163,N_2365,N_2019);
or U5164 (N_5164,N_817,N_2306);
or U5165 (N_5165,N_4,N_193);
and U5166 (N_5166,N_412,N_370);
and U5167 (N_5167,N_2221,N_1045);
and U5168 (N_5168,N_795,N_2828);
and U5169 (N_5169,N_2364,N_428);
nand U5170 (N_5170,N_524,N_1332);
nand U5171 (N_5171,N_2264,N_1315);
nand U5172 (N_5172,N_1512,N_1982);
and U5173 (N_5173,N_1692,N_1889);
nor U5174 (N_5174,N_615,N_1440);
nand U5175 (N_5175,N_624,N_2476);
nand U5176 (N_5176,N_2356,N_2877);
or U5177 (N_5177,N_25,N_1747);
nor U5178 (N_5178,N_2424,N_1923);
nand U5179 (N_5179,N_2922,N_1880);
nor U5180 (N_5180,N_1351,N_2167);
nand U5181 (N_5181,N_574,N_2151);
or U5182 (N_5182,N_1519,N_2003);
or U5183 (N_5183,N_834,N_1151);
or U5184 (N_5184,N_2604,N_814);
nand U5185 (N_5185,N_930,N_1296);
or U5186 (N_5186,N_191,N_740);
and U5187 (N_5187,N_1326,N_49);
or U5188 (N_5188,N_891,N_1989);
or U5189 (N_5189,N_532,N_960);
nor U5190 (N_5190,N_54,N_2631);
nor U5191 (N_5191,N_2581,N_2739);
or U5192 (N_5192,N_2741,N_386);
xnor U5193 (N_5193,N_1360,N_606);
xor U5194 (N_5194,N_1870,N_564);
and U5195 (N_5195,N_2604,N_2985);
or U5196 (N_5196,N_1799,N_1248);
and U5197 (N_5197,N_706,N_779);
and U5198 (N_5198,N_847,N_997);
xor U5199 (N_5199,N_612,N_2718);
and U5200 (N_5200,N_610,N_1052);
and U5201 (N_5201,N_1724,N_321);
or U5202 (N_5202,N_2001,N_2259);
and U5203 (N_5203,N_59,N_2888);
and U5204 (N_5204,N_1553,N_2141);
or U5205 (N_5205,N_532,N_1519);
and U5206 (N_5206,N_734,N_2675);
nand U5207 (N_5207,N_1693,N_564);
nor U5208 (N_5208,N_1643,N_2460);
or U5209 (N_5209,N_242,N_2991);
and U5210 (N_5210,N_1341,N_2052);
or U5211 (N_5211,N_1269,N_1257);
and U5212 (N_5212,N_2759,N_1133);
or U5213 (N_5213,N_2846,N_2117);
nand U5214 (N_5214,N_1947,N_101);
or U5215 (N_5215,N_31,N_1643);
or U5216 (N_5216,N_1223,N_1271);
nor U5217 (N_5217,N_2066,N_89);
and U5218 (N_5218,N_1440,N_2237);
nor U5219 (N_5219,N_2758,N_2053);
nand U5220 (N_5220,N_1426,N_2948);
and U5221 (N_5221,N_808,N_2047);
nand U5222 (N_5222,N_2554,N_2563);
nor U5223 (N_5223,N_433,N_2522);
and U5224 (N_5224,N_1178,N_2588);
and U5225 (N_5225,N_874,N_699);
and U5226 (N_5226,N_3011,N_727);
nor U5227 (N_5227,N_3050,N_2828);
nor U5228 (N_5228,N_1425,N_1009);
and U5229 (N_5229,N_2927,N_2816);
nor U5230 (N_5230,N_436,N_2914);
or U5231 (N_5231,N_2542,N_2891);
and U5232 (N_5232,N_1473,N_2671);
nand U5233 (N_5233,N_2198,N_2734);
and U5234 (N_5234,N_1317,N_1308);
nand U5235 (N_5235,N_470,N_2624);
and U5236 (N_5236,N_2356,N_3068);
nor U5237 (N_5237,N_1852,N_2721);
or U5238 (N_5238,N_691,N_1330);
or U5239 (N_5239,N_2777,N_106);
nand U5240 (N_5240,N_2270,N_880);
nand U5241 (N_5241,N_2996,N_1448);
nor U5242 (N_5242,N_17,N_2880);
and U5243 (N_5243,N_199,N_2220);
or U5244 (N_5244,N_274,N_2663);
nand U5245 (N_5245,N_1807,N_886);
nor U5246 (N_5246,N_1585,N_870);
nor U5247 (N_5247,N_1426,N_2228);
nand U5248 (N_5248,N_670,N_1904);
or U5249 (N_5249,N_1208,N_2738);
or U5250 (N_5250,N_419,N_1813);
and U5251 (N_5251,N_2586,N_2082);
nand U5252 (N_5252,N_865,N_814);
and U5253 (N_5253,N_1367,N_487);
or U5254 (N_5254,N_1014,N_2529);
nand U5255 (N_5255,N_537,N_581);
xor U5256 (N_5256,N_399,N_2209);
and U5257 (N_5257,N_1696,N_2964);
nor U5258 (N_5258,N_1043,N_1469);
nor U5259 (N_5259,N_1651,N_426);
or U5260 (N_5260,N_3124,N_2110);
nor U5261 (N_5261,N_2719,N_751);
nand U5262 (N_5262,N_2070,N_1311);
xnor U5263 (N_5263,N_2748,N_2181);
nor U5264 (N_5264,N_2899,N_820);
nand U5265 (N_5265,N_1303,N_2826);
nor U5266 (N_5266,N_2635,N_232);
or U5267 (N_5267,N_2150,N_858);
and U5268 (N_5268,N_1966,N_3111);
or U5269 (N_5269,N_883,N_323);
nand U5270 (N_5270,N_2861,N_469);
nor U5271 (N_5271,N_2614,N_1052);
nand U5272 (N_5272,N_1159,N_2666);
nand U5273 (N_5273,N_2236,N_1324);
nor U5274 (N_5274,N_2729,N_1330);
nand U5275 (N_5275,N_881,N_2552);
and U5276 (N_5276,N_1517,N_960);
nor U5277 (N_5277,N_2809,N_3081);
and U5278 (N_5278,N_2002,N_2898);
xor U5279 (N_5279,N_255,N_417);
nand U5280 (N_5280,N_658,N_472);
nor U5281 (N_5281,N_880,N_584);
or U5282 (N_5282,N_2212,N_1143);
nor U5283 (N_5283,N_1815,N_3);
nand U5284 (N_5284,N_468,N_1249);
or U5285 (N_5285,N_3109,N_936);
or U5286 (N_5286,N_2901,N_2841);
nor U5287 (N_5287,N_909,N_886);
or U5288 (N_5288,N_1834,N_2228);
and U5289 (N_5289,N_2064,N_84);
and U5290 (N_5290,N_451,N_1529);
nand U5291 (N_5291,N_1431,N_332);
nand U5292 (N_5292,N_231,N_3079);
nand U5293 (N_5293,N_1872,N_104);
nand U5294 (N_5294,N_2562,N_1850);
nand U5295 (N_5295,N_1036,N_2257);
nor U5296 (N_5296,N_798,N_398);
or U5297 (N_5297,N_2536,N_41);
nand U5298 (N_5298,N_3010,N_2868);
nand U5299 (N_5299,N_1730,N_3039);
nand U5300 (N_5300,N_120,N_2200);
nor U5301 (N_5301,N_2103,N_2748);
or U5302 (N_5302,N_1752,N_204);
or U5303 (N_5303,N_2712,N_406);
nand U5304 (N_5304,N_370,N_2983);
or U5305 (N_5305,N_1529,N_2190);
xnor U5306 (N_5306,N_303,N_1850);
nand U5307 (N_5307,N_449,N_2004);
nor U5308 (N_5308,N_1607,N_2327);
xnor U5309 (N_5309,N_131,N_836);
and U5310 (N_5310,N_592,N_1711);
or U5311 (N_5311,N_2737,N_1461);
nor U5312 (N_5312,N_1931,N_231);
nor U5313 (N_5313,N_298,N_1523);
nand U5314 (N_5314,N_993,N_2217);
or U5315 (N_5315,N_2091,N_1873);
nand U5316 (N_5316,N_1618,N_2404);
nand U5317 (N_5317,N_1119,N_2681);
and U5318 (N_5318,N_403,N_1550);
and U5319 (N_5319,N_2130,N_2823);
xor U5320 (N_5320,N_2940,N_1140);
nand U5321 (N_5321,N_3076,N_980);
nor U5322 (N_5322,N_1273,N_1131);
xor U5323 (N_5323,N_606,N_3104);
nor U5324 (N_5324,N_1155,N_637);
and U5325 (N_5325,N_1376,N_568);
or U5326 (N_5326,N_3080,N_950);
xor U5327 (N_5327,N_1396,N_2650);
nor U5328 (N_5328,N_2036,N_2919);
and U5329 (N_5329,N_1519,N_396);
nand U5330 (N_5330,N_2860,N_1073);
nand U5331 (N_5331,N_2483,N_1645);
nand U5332 (N_5332,N_708,N_1196);
and U5333 (N_5333,N_2708,N_2623);
and U5334 (N_5334,N_2279,N_3072);
nand U5335 (N_5335,N_2335,N_173);
and U5336 (N_5336,N_1072,N_524);
nor U5337 (N_5337,N_1523,N_1317);
xnor U5338 (N_5338,N_1858,N_1513);
or U5339 (N_5339,N_3112,N_1153);
nand U5340 (N_5340,N_582,N_2188);
and U5341 (N_5341,N_2419,N_1462);
xor U5342 (N_5342,N_1121,N_209);
nand U5343 (N_5343,N_1867,N_3042);
nand U5344 (N_5344,N_2751,N_1749);
nor U5345 (N_5345,N_2411,N_97);
or U5346 (N_5346,N_3116,N_664);
or U5347 (N_5347,N_2805,N_2483);
nor U5348 (N_5348,N_2235,N_500);
nand U5349 (N_5349,N_2627,N_1566);
nor U5350 (N_5350,N_2477,N_2773);
or U5351 (N_5351,N_2667,N_1913);
nand U5352 (N_5352,N_1757,N_1673);
nand U5353 (N_5353,N_2290,N_1735);
nor U5354 (N_5354,N_2985,N_1459);
and U5355 (N_5355,N_113,N_1437);
xnor U5356 (N_5356,N_2844,N_96);
nor U5357 (N_5357,N_2937,N_2970);
nand U5358 (N_5358,N_1383,N_965);
and U5359 (N_5359,N_1332,N_129);
nor U5360 (N_5360,N_1860,N_905);
nor U5361 (N_5361,N_117,N_2439);
or U5362 (N_5362,N_1422,N_1065);
nand U5363 (N_5363,N_1096,N_288);
or U5364 (N_5364,N_1364,N_2895);
nor U5365 (N_5365,N_953,N_2009);
nand U5366 (N_5366,N_1959,N_1255);
xor U5367 (N_5367,N_2350,N_1056);
nand U5368 (N_5368,N_3071,N_2530);
nor U5369 (N_5369,N_2686,N_2353);
nor U5370 (N_5370,N_2131,N_1058);
nand U5371 (N_5371,N_2665,N_2119);
xor U5372 (N_5372,N_1990,N_1977);
and U5373 (N_5373,N_2699,N_861);
or U5374 (N_5374,N_965,N_869);
nand U5375 (N_5375,N_154,N_1036);
nor U5376 (N_5376,N_1441,N_293);
nor U5377 (N_5377,N_751,N_1775);
and U5378 (N_5378,N_2996,N_2385);
xnor U5379 (N_5379,N_920,N_433);
or U5380 (N_5380,N_216,N_194);
nand U5381 (N_5381,N_437,N_1352);
nor U5382 (N_5382,N_1252,N_1012);
nand U5383 (N_5383,N_2498,N_2111);
and U5384 (N_5384,N_712,N_351);
or U5385 (N_5385,N_2033,N_844);
nor U5386 (N_5386,N_1510,N_767);
nand U5387 (N_5387,N_2925,N_1209);
nor U5388 (N_5388,N_1595,N_1471);
nand U5389 (N_5389,N_2541,N_1141);
or U5390 (N_5390,N_1426,N_567);
and U5391 (N_5391,N_3069,N_2077);
and U5392 (N_5392,N_1766,N_112);
or U5393 (N_5393,N_1866,N_646);
and U5394 (N_5394,N_896,N_1023);
or U5395 (N_5395,N_1100,N_2196);
and U5396 (N_5396,N_488,N_1936);
or U5397 (N_5397,N_1729,N_1332);
nand U5398 (N_5398,N_518,N_1295);
nor U5399 (N_5399,N_2189,N_2308);
nor U5400 (N_5400,N_926,N_328);
nand U5401 (N_5401,N_571,N_781);
nand U5402 (N_5402,N_107,N_397);
or U5403 (N_5403,N_1594,N_2368);
nor U5404 (N_5404,N_506,N_513);
nor U5405 (N_5405,N_398,N_1476);
and U5406 (N_5406,N_446,N_946);
xnor U5407 (N_5407,N_936,N_2114);
and U5408 (N_5408,N_691,N_2644);
or U5409 (N_5409,N_748,N_765);
xor U5410 (N_5410,N_2222,N_158);
nand U5411 (N_5411,N_1551,N_1595);
nand U5412 (N_5412,N_1850,N_89);
nor U5413 (N_5413,N_1489,N_2999);
or U5414 (N_5414,N_2541,N_2288);
and U5415 (N_5415,N_358,N_2745);
or U5416 (N_5416,N_1523,N_599);
or U5417 (N_5417,N_231,N_2817);
nand U5418 (N_5418,N_1654,N_553);
nor U5419 (N_5419,N_2008,N_1120);
nor U5420 (N_5420,N_150,N_3049);
nand U5421 (N_5421,N_1429,N_1519);
nor U5422 (N_5422,N_1114,N_719);
and U5423 (N_5423,N_2213,N_1808);
xnor U5424 (N_5424,N_2649,N_2345);
nand U5425 (N_5425,N_1899,N_232);
nor U5426 (N_5426,N_1512,N_3067);
nor U5427 (N_5427,N_3024,N_2117);
and U5428 (N_5428,N_900,N_635);
nor U5429 (N_5429,N_1718,N_410);
nor U5430 (N_5430,N_2474,N_2282);
and U5431 (N_5431,N_1321,N_2468);
nand U5432 (N_5432,N_30,N_938);
and U5433 (N_5433,N_461,N_592);
nand U5434 (N_5434,N_752,N_2917);
and U5435 (N_5435,N_1681,N_2653);
or U5436 (N_5436,N_2937,N_87);
and U5437 (N_5437,N_182,N_993);
nor U5438 (N_5438,N_2738,N_564);
and U5439 (N_5439,N_2588,N_2722);
or U5440 (N_5440,N_1323,N_2322);
and U5441 (N_5441,N_1678,N_1702);
nor U5442 (N_5442,N_2831,N_2731);
nand U5443 (N_5443,N_464,N_2872);
nand U5444 (N_5444,N_598,N_831);
xor U5445 (N_5445,N_2411,N_606);
and U5446 (N_5446,N_1998,N_2529);
and U5447 (N_5447,N_2018,N_2595);
nand U5448 (N_5448,N_237,N_198);
and U5449 (N_5449,N_208,N_1412);
nor U5450 (N_5450,N_2838,N_3110);
or U5451 (N_5451,N_961,N_2573);
or U5452 (N_5452,N_2476,N_1738);
nor U5453 (N_5453,N_7,N_627);
or U5454 (N_5454,N_1292,N_1094);
xnor U5455 (N_5455,N_980,N_1098);
xor U5456 (N_5456,N_310,N_392);
and U5457 (N_5457,N_1932,N_2985);
xor U5458 (N_5458,N_2509,N_2206);
nor U5459 (N_5459,N_2958,N_1826);
nor U5460 (N_5460,N_458,N_1838);
or U5461 (N_5461,N_826,N_36);
and U5462 (N_5462,N_2580,N_2515);
nor U5463 (N_5463,N_1436,N_205);
or U5464 (N_5464,N_1231,N_2126);
xnor U5465 (N_5465,N_505,N_573);
or U5466 (N_5466,N_2725,N_2434);
nor U5467 (N_5467,N_645,N_1996);
nor U5468 (N_5468,N_225,N_2158);
nor U5469 (N_5469,N_2183,N_2468);
or U5470 (N_5470,N_646,N_3011);
and U5471 (N_5471,N_2876,N_1182);
nor U5472 (N_5472,N_2598,N_2147);
xnor U5473 (N_5473,N_1630,N_2072);
nor U5474 (N_5474,N_2117,N_2929);
nor U5475 (N_5475,N_2657,N_3094);
and U5476 (N_5476,N_912,N_300);
nand U5477 (N_5477,N_429,N_2293);
nand U5478 (N_5478,N_7,N_1008);
or U5479 (N_5479,N_2895,N_840);
or U5480 (N_5480,N_2863,N_221);
nand U5481 (N_5481,N_1225,N_1915);
nand U5482 (N_5482,N_556,N_2188);
nor U5483 (N_5483,N_2964,N_1031);
nor U5484 (N_5484,N_197,N_2783);
nor U5485 (N_5485,N_1424,N_1579);
or U5486 (N_5486,N_235,N_1494);
and U5487 (N_5487,N_3116,N_688);
xnor U5488 (N_5488,N_623,N_1621);
nand U5489 (N_5489,N_2774,N_1411);
and U5490 (N_5490,N_371,N_1298);
xnor U5491 (N_5491,N_2649,N_1124);
and U5492 (N_5492,N_1566,N_247);
nand U5493 (N_5493,N_1569,N_2939);
or U5494 (N_5494,N_339,N_214);
nand U5495 (N_5495,N_2490,N_1611);
or U5496 (N_5496,N_870,N_1277);
xnor U5497 (N_5497,N_2364,N_2354);
and U5498 (N_5498,N_1312,N_2044);
nor U5499 (N_5499,N_234,N_1732);
nor U5500 (N_5500,N_2074,N_258);
nor U5501 (N_5501,N_2281,N_2785);
or U5502 (N_5502,N_992,N_191);
xor U5503 (N_5503,N_622,N_502);
nor U5504 (N_5504,N_1422,N_1167);
and U5505 (N_5505,N_84,N_2375);
or U5506 (N_5506,N_366,N_345);
and U5507 (N_5507,N_2632,N_29);
nor U5508 (N_5508,N_2031,N_1932);
nand U5509 (N_5509,N_2235,N_3035);
nand U5510 (N_5510,N_1154,N_799);
and U5511 (N_5511,N_516,N_661);
and U5512 (N_5512,N_1794,N_1340);
or U5513 (N_5513,N_1528,N_1679);
and U5514 (N_5514,N_2129,N_2456);
nor U5515 (N_5515,N_2495,N_879);
xor U5516 (N_5516,N_2691,N_139);
or U5517 (N_5517,N_803,N_2388);
nand U5518 (N_5518,N_2605,N_1378);
xor U5519 (N_5519,N_1903,N_1714);
nand U5520 (N_5520,N_1313,N_2782);
or U5521 (N_5521,N_91,N_2042);
nand U5522 (N_5522,N_1348,N_140);
or U5523 (N_5523,N_574,N_1937);
nor U5524 (N_5524,N_1757,N_1913);
or U5525 (N_5525,N_1505,N_2122);
xor U5526 (N_5526,N_2513,N_91);
and U5527 (N_5527,N_1821,N_1807);
nand U5528 (N_5528,N_112,N_2301);
nor U5529 (N_5529,N_2343,N_576);
nand U5530 (N_5530,N_449,N_610);
nand U5531 (N_5531,N_2695,N_2867);
xor U5532 (N_5532,N_3089,N_1939);
and U5533 (N_5533,N_2304,N_1552);
nand U5534 (N_5534,N_2541,N_1360);
xor U5535 (N_5535,N_1790,N_2153);
and U5536 (N_5536,N_3053,N_2121);
nor U5537 (N_5537,N_2659,N_267);
nand U5538 (N_5538,N_2660,N_1354);
nor U5539 (N_5539,N_1618,N_1981);
and U5540 (N_5540,N_2584,N_2629);
nand U5541 (N_5541,N_2778,N_1439);
nor U5542 (N_5542,N_2498,N_1957);
nand U5543 (N_5543,N_1729,N_2446);
nor U5544 (N_5544,N_2415,N_1708);
nand U5545 (N_5545,N_400,N_123);
and U5546 (N_5546,N_1617,N_2377);
or U5547 (N_5547,N_409,N_580);
nand U5548 (N_5548,N_691,N_1542);
and U5549 (N_5549,N_2962,N_2832);
nand U5550 (N_5550,N_2956,N_2614);
nand U5551 (N_5551,N_2653,N_2424);
and U5552 (N_5552,N_1556,N_1110);
and U5553 (N_5553,N_2104,N_2842);
and U5554 (N_5554,N_1049,N_561);
nand U5555 (N_5555,N_631,N_2071);
nor U5556 (N_5556,N_649,N_453);
nor U5557 (N_5557,N_2149,N_2055);
and U5558 (N_5558,N_219,N_3002);
xor U5559 (N_5559,N_3039,N_1626);
or U5560 (N_5560,N_1376,N_2538);
nor U5561 (N_5561,N_2010,N_752);
nor U5562 (N_5562,N_793,N_1120);
nor U5563 (N_5563,N_3018,N_3094);
nor U5564 (N_5564,N_866,N_677);
nor U5565 (N_5565,N_1335,N_125);
nor U5566 (N_5566,N_1985,N_212);
and U5567 (N_5567,N_942,N_1887);
xnor U5568 (N_5568,N_758,N_3109);
xnor U5569 (N_5569,N_1108,N_1769);
or U5570 (N_5570,N_2751,N_412);
and U5571 (N_5571,N_2629,N_2920);
nand U5572 (N_5572,N_3008,N_1476);
and U5573 (N_5573,N_2390,N_1918);
or U5574 (N_5574,N_2051,N_545);
nand U5575 (N_5575,N_2430,N_983);
and U5576 (N_5576,N_1412,N_2013);
xor U5577 (N_5577,N_158,N_843);
or U5578 (N_5578,N_576,N_927);
nand U5579 (N_5579,N_1793,N_512);
and U5580 (N_5580,N_1590,N_1755);
nand U5581 (N_5581,N_2500,N_1093);
xnor U5582 (N_5582,N_1517,N_2944);
nand U5583 (N_5583,N_1940,N_814);
nand U5584 (N_5584,N_2428,N_1317);
xnor U5585 (N_5585,N_2058,N_409);
nand U5586 (N_5586,N_2339,N_2705);
or U5587 (N_5587,N_277,N_2682);
nand U5588 (N_5588,N_592,N_2796);
nor U5589 (N_5589,N_2713,N_2493);
or U5590 (N_5590,N_1193,N_1396);
nor U5591 (N_5591,N_12,N_2513);
and U5592 (N_5592,N_2736,N_926);
nand U5593 (N_5593,N_3066,N_1284);
or U5594 (N_5594,N_2371,N_1738);
and U5595 (N_5595,N_1122,N_1438);
nand U5596 (N_5596,N_3014,N_1420);
nor U5597 (N_5597,N_2149,N_605);
nor U5598 (N_5598,N_2216,N_1255);
and U5599 (N_5599,N_427,N_2348);
and U5600 (N_5600,N_1349,N_2156);
or U5601 (N_5601,N_582,N_2621);
or U5602 (N_5602,N_1851,N_627);
nand U5603 (N_5603,N_1243,N_920);
xor U5604 (N_5604,N_253,N_132);
nor U5605 (N_5605,N_1485,N_2625);
nand U5606 (N_5606,N_3078,N_660);
nor U5607 (N_5607,N_1354,N_2776);
and U5608 (N_5608,N_1163,N_1370);
or U5609 (N_5609,N_793,N_2782);
nor U5610 (N_5610,N_2525,N_1939);
nand U5611 (N_5611,N_2632,N_1074);
or U5612 (N_5612,N_1546,N_2503);
and U5613 (N_5613,N_545,N_225);
nand U5614 (N_5614,N_804,N_2279);
nand U5615 (N_5615,N_2873,N_788);
and U5616 (N_5616,N_480,N_2008);
nor U5617 (N_5617,N_2212,N_253);
and U5618 (N_5618,N_2642,N_2802);
nor U5619 (N_5619,N_435,N_2384);
or U5620 (N_5620,N_1340,N_1242);
or U5621 (N_5621,N_939,N_923);
and U5622 (N_5622,N_1378,N_2021);
and U5623 (N_5623,N_3115,N_1658);
nor U5624 (N_5624,N_1257,N_849);
nor U5625 (N_5625,N_444,N_1004);
or U5626 (N_5626,N_2031,N_623);
nand U5627 (N_5627,N_2014,N_364);
xnor U5628 (N_5628,N_421,N_789);
nand U5629 (N_5629,N_17,N_2267);
nor U5630 (N_5630,N_1095,N_333);
and U5631 (N_5631,N_387,N_1638);
and U5632 (N_5632,N_2027,N_1865);
or U5633 (N_5633,N_577,N_123);
and U5634 (N_5634,N_787,N_612);
nand U5635 (N_5635,N_3124,N_1846);
and U5636 (N_5636,N_1285,N_1470);
and U5637 (N_5637,N_1055,N_989);
nor U5638 (N_5638,N_1983,N_2196);
or U5639 (N_5639,N_1909,N_83);
nor U5640 (N_5640,N_3091,N_2314);
nor U5641 (N_5641,N_82,N_2663);
and U5642 (N_5642,N_552,N_2535);
xor U5643 (N_5643,N_385,N_1237);
nor U5644 (N_5644,N_1130,N_2673);
and U5645 (N_5645,N_3071,N_2859);
nand U5646 (N_5646,N_983,N_205);
or U5647 (N_5647,N_142,N_2353);
and U5648 (N_5648,N_612,N_2127);
and U5649 (N_5649,N_2773,N_443);
and U5650 (N_5650,N_3086,N_1237);
and U5651 (N_5651,N_1337,N_2406);
nor U5652 (N_5652,N_2606,N_2667);
and U5653 (N_5653,N_918,N_2444);
nor U5654 (N_5654,N_38,N_1970);
xnor U5655 (N_5655,N_325,N_1934);
nand U5656 (N_5656,N_2652,N_1218);
or U5657 (N_5657,N_501,N_221);
nor U5658 (N_5658,N_2113,N_2287);
or U5659 (N_5659,N_1943,N_1178);
and U5660 (N_5660,N_1209,N_2115);
xor U5661 (N_5661,N_1371,N_2517);
nor U5662 (N_5662,N_764,N_863);
and U5663 (N_5663,N_214,N_2715);
nand U5664 (N_5664,N_2585,N_263);
or U5665 (N_5665,N_3122,N_2871);
or U5666 (N_5666,N_2838,N_2199);
or U5667 (N_5667,N_268,N_568);
or U5668 (N_5668,N_655,N_916);
or U5669 (N_5669,N_2161,N_1568);
nand U5670 (N_5670,N_2252,N_2955);
nand U5671 (N_5671,N_1748,N_1712);
and U5672 (N_5672,N_2101,N_2445);
and U5673 (N_5673,N_2664,N_717);
and U5674 (N_5674,N_991,N_3048);
xor U5675 (N_5675,N_818,N_2072);
and U5676 (N_5676,N_1318,N_3122);
nand U5677 (N_5677,N_945,N_1101);
or U5678 (N_5678,N_1611,N_1598);
nor U5679 (N_5679,N_2643,N_464);
and U5680 (N_5680,N_881,N_2085);
and U5681 (N_5681,N_1674,N_1283);
nor U5682 (N_5682,N_934,N_739);
nor U5683 (N_5683,N_165,N_394);
or U5684 (N_5684,N_2881,N_2617);
nand U5685 (N_5685,N_1716,N_239);
or U5686 (N_5686,N_1006,N_2011);
and U5687 (N_5687,N_1936,N_2745);
nand U5688 (N_5688,N_2861,N_2405);
and U5689 (N_5689,N_714,N_467);
and U5690 (N_5690,N_2671,N_1378);
nand U5691 (N_5691,N_910,N_1033);
nor U5692 (N_5692,N_315,N_2681);
or U5693 (N_5693,N_2821,N_699);
nor U5694 (N_5694,N_562,N_258);
xor U5695 (N_5695,N_2583,N_662);
or U5696 (N_5696,N_2372,N_205);
nor U5697 (N_5697,N_1150,N_2354);
xnor U5698 (N_5698,N_347,N_1755);
nand U5699 (N_5699,N_507,N_2365);
nand U5700 (N_5700,N_2567,N_1002);
nand U5701 (N_5701,N_1279,N_2724);
nand U5702 (N_5702,N_757,N_1431);
and U5703 (N_5703,N_396,N_3049);
and U5704 (N_5704,N_2283,N_336);
xor U5705 (N_5705,N_1360,N_2671);
nand U5706 (N_5706,N_3033,N_1928);
nor U5707 (N_5707,N_2685,N_2309);
or U5708 (N_5708,N_1753,N_2936);
nor U5709 (N_5709,N_1667,N_3042);
or U5710 (N_5710,N_2572,N_1992);
or U5711 (N_5711,N_798,N_2060);
nor U5712 (N_5712,N_1702,N_1971);
and U5713 (N_5713,N_1717,N_2426);
and U5714 (N_5714,N_2025,N_1086);
nor U5715 (N_5715,N_794,N_2039);
nand U5716 (N_5716,N_2538,N_2712);
nor U5717 (N_5717,N_221,N_1373);
xor U5718 (N_5718,N_2315,N_1867);
nand U5719 (N_5719,N_2208,N_2350);
or U5720 (N_5720,N_1680,N_855);
nand U5721 (N_5721,N_1664,N_1155);
or U5722 (N_5722,N_490,N_1546);
or U5723 (N_5723,N_308,N_2547);
or U5724 (N_5724,N_2178,N_633);
xnor U5725 (N_5725,N_1466,N_1085);
xnor U5726 (N_5726,N_3097,N_781);
and U5727 (N_5727,N_2811,N_452);
nand U5728 (N_5728,N_2697,N_2079);
or U5729 (N_5729,N_2417,N_636);
nand U5730 (N_5730,N_1854,N_360);
nor U5731 (N_5731,N_504,N_2125);
nor U5732 (N_5732,N_1481,N_204);
and U5733 (N_5733,N_2086,N_750);
or U5734 (N_5734,N_1827,N_1872);
and U5735 (N_5735,N_2699,N_1470);
and U5736 (N_5736,N_1417,N_1536);
xor U5737 (N_5737,N_2064,N_828);
or U5738 (N_5738,N_2681,N_3119);
xor U5739 (N_5739,N_1892,N_750);
nor U5740 (N_5740,N_1887,N_1561);
nor U5741 (N_5741,N_1078,N_2517);
or U5742 (N_5742,N_247,N_2513);
nor U5743 (N_5743,N_1675,N_695);
nor U5744 (N_5744,N_3049,N_1433);
nor U5745 (N_5745,N_590,N_2038);
and U5746 (N_5746,N_2523,N_2305);
and U5747 (N_5747,N_1441,N_2057);
and U5748 (N_5748,N_514,N_1729);
or U5749 (N_5749,N_1021,N_1019);
and U5750 (N_5750,N_2052,N_1465);
nor U5751 (N_5751,N_2569,N_685);
or U5752 (N_5752,N_1173,N_489);
or U5753 (N_5753,N_217,N_502);
nand U5754 (N_5754,N_2833,N_2447);
nor U5755 (N_5755,N_482,N_1734);
and U5756 (N_5756,N_1614,N_541);
xnor U5757 (N_5757,N_1088,N_1446);
nor U5758 (N_5758,N_38,N_3014);
nor U5759 (N_5759,N_1193,N_1737);
and U5760 (N_5760,N_775,N_3121);
nor U5761 (N_5761,N_2840,N_2928);
and U5762 (N_5762,N_2540,N_462);
or U5763 (N_5763,N_2519,N_124);
nand U5764 (N_5764,N_1804,N_1945);
nand U5765 (N_5765,N_1332,N_2477);
or U5766 (N_5766,N_2279,N_543);
xor U5767 (N_5767,N_1377,N_1787);
nand U5768 (N_5768,N_817,N_1710);
or U5769 (N_5769,N_2587,N_2451);
and U5770 (N_5770,N_1663,N_1618);
or U5771 (N_5771,N_3050,N_39);
and U5772 (N_5772,N_3008,N_2111);
or U5773 (N_5773,N_1543,N_2847);
and U5774 (N_5774,N_1676,N_476);
nand U5775 (N_5775,N_1857,N_1957);
nor U5776 (N_5776,N_487,N_1540);
xor U5777 (N_5777,N_644,N_1462);
or U5778 (N_5778,N_767,N_2818);
nand U5779 (N_5779,N_1582,N_2953);
or U5780 (N_5780,N_635,N_658);
or U5781 (N_5781,N_2863,N_1999);
nor U5782 (N_5782,N_1118,N_1433);
nand U5783 (N_5783,N_1577,N_140);
or U5784 (N_5784,N_392,N_881);
and U5785 (N_5785,N_779,N_2775);
nor U5786 (N_5786,N_1103,N_44);
and U5787 (N_5787,N_1437,N_168);
nor U5788 (N_5788,N_1924,N_452);
nand U5789 (N_5789,N_2270,N_1755);
and U5790 (N_5790,N_988,N_1838);
and U5791 (N_5791,N_1537,N_2310);
nand U5792 (N_5792,N_2189,N_773);
and U5793 (N_5793,N_2124,N_2666);
and U5794 (N_5794,N_2130,N_222);
or U5795 (N_5795,N_214,N_205);
nand U5796 (N_5796,N_622,N_244);
or U5797 (N_5797,N_2990,N_143);
or U5798 (N_5798,N_2978,N_2402);
xnor U5799 (N_5799,N_1708,N_2351);
or U5800 (N_5800,N_1026,N_2674);
nand U5801 (N_5801,N_619,N_293);
nor U5802 (N_5802,N_1506,N_1452);
nor U5803 (N_5803,N_1963,N_1561);
or U5804 (N_5804,N_1620,N_368);
nand U5805 (N_5805,N_2101,N_256);
and U5806 (N_5806,N_296,N_1832);
or U5807 (N_5807,N_2780,N_1485);
nor U5808 (N_5808,N_214,N_1914);
nor U5809 (N_5809,N_1887,N_106);
nand U5810 (N_5810,N_1207,N_1929);
nor U5811 (N_5811,N_2029,N_1140);
nor U5812 (N_5812,N_758,N_223);
and U5813 (N_5813,N_1554,N_1289);
nand U5814 (N_5814,N_1076,N_127);
and U5815 (N_5815,N_2809,N_2779);
nor U5816 (N_5816,N_3056,N_861);
nand U5817 (N_5817,N_3009,N_2581);
and U5818 (N_5818,N_1008,N_1399);
nor U5819 (N_5819,N_1244,N_1216);
nor U5820 (N_5820,N_1591,N_1370);
xnor U5821 (N_5821,N_1407,N_834);
nor U5822 (N_5822,N_1019,N_2345);
xnor U5823 (N_5823,N_1872,N_1927);
nand U5824 (N_5824,N_1812,N_2493);
and U5825 (N_5825,N_1683,N_463);
nor U5826 (N_5826,N_900,N_510);
nor U5827 (N_5827,N_2314,N_489);
nand U5828 (N_5828,N_2338,N_1814);
nand U5829 (N_5829,N_2910,N_2283);
nand U5830 (N_5830,N_255,N_250);
nand U5831 (N_5831,N_2231,N_954);
xor U5832 (N_5832,N_864,N_1636);
nor U5833 (N_5833,N_1676,N_2594);
and U5834 (N_5834,N_3007,N_1484);
nand U5835 (N_5835,N_1326,N_520);
nor U5836 (N_5836,N_1339,N_3074);
nand U5837 (N_5837,N_2403,N_801);
and U5838 (N_5838,N_1885,N_1737);
and U5839 (N_5839,N_629,N_363);
nor U5840 (N_5840,N_1429,N_2328);
or U5841 (N_5841,N_749,N_2693);
nor U5842 (N_5842,N_1011,N_71);
nor U5843 (N_5843,N_2202,N_2071);
nor U5844 (N_5844,N_661,N_2782);
and U5845 (N_5845,N_379,N_1393);
nor U5846 (N_5846,N_1575,N_218);
or U5847 (N_5847,N_1084,N_513);
nand U5848 (N_5848,N_1184,N_3029);
or U5849 (N_5849,N_1344,N_2540);
or U5850 (N_5850,N_1709,N_1820);
or U5851 (N_5851,N_2574,N_1832);
nor U5852 (N_5852,N_2308,N_1418);
or U5853 (N_5853,N_1783,N_1690);
and U5854 (N_5854,N_240,N_2385);
and U5855 (N_5855,N_653,N_1887);
and U5856 (N_5856,N_593,N_2519);
and U5857 (N_5857,N_2173,N_207);
and U5858 (N_5858,N_2398,N_2587);
xor U5859 (N_5859,N_1334,N_704);
xnor U5860 (N_5860,N_637,N_1439);
nand U5861 (N_5861,N_485,N_395);
and U5862 (N_5862,N_2832,N_970);
nand U5863 (N_5863,N_740,N_1273);
or U5864 (N_5864,N_2154,N_2305);
xnor U5865 (N_5865,N_1484,N_1221);
or U5866 (N_5866,N_2642,N_671);
or U5867 (N_5867,N_430,N_1644);
or U5868 (N_5868,N_1178,N_266);
or U5869 (N_5869,N_513,N_910);
and U5870 (N_5870,N_1438,N_1129);
or U5871 (N_5871,N_1476,N_438);
or U5872 (N_5872,N_303,N_12);
nand U5873 (N_5873,N_2448,N_629);
nand U5874 (N_5874,N_1811,N_872);
or U5875 (N_5875,N_424,N_3039);
or U5876 (N_5876,N_1334,N_1010);
and U5877 (N_5877,N_1228,N_2095);
or U5878 (N_5878,N_1056,N_583);
or U5879 (N_5879,N_3034,N_1149);
or U5880 (N_5880,N_1373,N_1712);
or U5881 (N_5881,N_2501,N_623);
nand U5882 (N_5882,N_2548,N_541);
and U5883 (N_5883,N_754,N_741);
or U5884 (N_5884,N_2208,N_2885);
xor U5885 (N_5885,N_2974,N_354);
xnor U5886 (N_5886,N_3082,N_1350);
nand U5887 (N_5887,N_2103,N_56);
nand U5888 (N_5888,N_2469,N_1906);
and U5889 (N_5889,N_847,N_3117);
xnor U5890 (N_5890,N_874,N_2405);
and U5891 (N_5891,N_2503,N_2367);
nand U5892 (N_5892,N_2789,N_1423);
and U5893 (N_5893,N_3087,N_1745);
and U5894 (N_5894,N_2068,N_1521);
xor U5895 (N_5895,N_2279,N_1722);
xor U5896 (N_5896,N_1465,N_2633);
nand U5897 (N_5897,N_1905,N_1197);
nand U5898 (N_5898,N_195,N_1516);
nand U5899 (N_5899,N_2708,N_2099);
and U5900 (N_5900,N_2003,N_2101);
xor U5901 (N_5901,N_2332,N_2362);
and U5902 (N_5902,N_2443,N_2594);
nor U5903 (N_5903,N_1495,N_2529);
nand U5904 (N_5904,N_111,N_1797);
and U5905 (N_5905,N_2887,N_803);
and U5906 (N_5906,N_368,N_1296);
or U5907 (N_5907,N_1162,N_1440);
xnor U5908 (N_5908,N_973,N_982);
nor U5909 (N_5909,N_458,N_895);
nand U5910 (N_5910,N_2372,N_1181);
nand U5911 (N_5911,N_1470,N_2701);
and U5912 (N_5912,N_237,N_2599);
xor U5913 (N_5913,N_2357,N_594);
or U5914 (N_5914,N_1901,N_773);
or U5915 (N_5915,N_661,N_1725);
nand U5916 (N_5916,N_721,N_43);
nand U5917 (N_5917,N_2454,N_2255);
nor U5918 (N_5918,N_2931,N_2895);
and U5919 (N_5919,N_272,N_164);
nor U5920 (N_5920,N_2122,N_1375);
nor U5921 (N_5921,N_1174,N_2950);
xor U5922 (N_5922,N_549,N_2496);
nor U5923 (N_5923,N_776,N_1179);
nand U5924 (N_5924,N_3070,N_1205);
and U5925 (N_5925,N_2330,N_856);
or U5926 (N_5926,N_2485,N_1262);
and U5927 (N_5927,N_1896,N_1960);
xnor U5928 (N_5928,N_1502,N_1189);
or U5929 (N_5929,N_2043,N_1031);
and U5930 (N_5930,N_64,N_2228);
nand U5931 (N_5931,N_157,N_890);
or U5932 (N_5932,N_37,N_241);
nand U5933 (N_5933,N_1157,N_2308);
nand U5934 (N_5934,N_2720,N_3098);
nand U5935 (N_5935,N_2280,N_2340);
nor U5936 (N_5936,N_1659,N_2028);
nand U5937 (N_5937,N_2161,N_1588);
or U5938 (N_5938,N_464,N_1177);
or U5939 (N_5939,N_2639,N_1818);
nor U5940 (N_5940,N_2647,N_74);
nand U5941 (N_5941,N_2566,N_2008);
and U5942 (N_5942,N_535,N_3008);
or U5943 (N_5943,N_1151,N_3035);
and U5944 (N_5944,N_1611,N_1834);
xnor U5945 (N_5945,N_1252,N_868);
nand U5946 (N_5946,N_1536,N_1105);
and U5947 (N_5947,N_709,N_1287);
nor U5948 (N_5948,N_1747,N_437);
and U5949 (N_5949,N_2407,N_1601);
or U5950 (N_5950,N_766,N_894);
and U5951 (N_5951,N_2548,N_1027);
or U5952 (N_5952,N_1698,N_1449);
nor U5953 (N_5953,N_274,N_1653);
nor U5954 (N_5954,N_2699,N_2105);
xor U5955 (N_5955,N_1806,N_2346);
nand U5956 (N_5956,N_735,N_2295);
nand U5957 (N_5957,N_2202,N_1523);
nor U5958 (N_5958,N_866,N_2824);
nor U5959 (N_5959,N_1312,N_846);
and U5960 (N_5960,N_2145,N_2778);
nand U5961 (N_5961,N_146,N_861);
and U5962 (N_5962,N_1627,N_2369);
xnor U5963 (N_5963,N_265,N_1421);
nor U5964 (N_5964,N_2740,N_510);
and U5965 (N_5965,N_1007,N_2921);
nor U5966 (N_5966,N_880,N_1788);
and U5967 (N_5967,N_2651,N_2949);
xor U5968 (N_5968,N_2756,N_1900);
and U5969 (N_5969,N_1290,N_562);
nor U5970 (N_5970,N_1368,N_73);
or U5971 (N_5971,N_1295,N_2357);
nor U5972 (N_5972,N_155,N_1723);
and U5973 (N_5973,N_187,N_1188);
or U5974 (N_5974,N_2173,N_2002);
and U5975 (N_5975,N_991,N_729);
and U5976 (N_5976,N_297,N_2166);
nor U5977 (N_5977,N_1015,N_2499);
nand U5978 (N_5978,N_2019,N_1386);
and U5979 (N_5979,N_788,N_1559);
and U5980 (N_5980,N_2347,N_2372);
nor U5981 (N_5981,N_2460,N_486);
or U5982 (N_5982,N_1480,N_1073);
xor U5983 (N_5983,N_2854,N_1956);
nor U5984 (N_5984,N_2345,N_2456);
nor U5985 (N_5985,N_525,N_2512);
xnor U5986 (N_5986,N_1460,N_266);
and U5987 (N_5987,N_1224,N_1938);
and U5988 (N_5988,N_785,N_1245);
nor U5989 (N_5989,N_773,N_847);
or U5990 (N_5990,N_687,N_2830);
nand U5991 (N_5991,N_1530,N_1188);
or U5992 (N_5992,N_2539,N_310);
or U5993 (N_5993,N_1186,N_1923);
xnor U5994 (N_5994,N_867,N_181);
or U5995 (N_5995,N_636,N_631);
or U5996 (N_5996,N_2190,N_793);
or U5997 (N_5997,N_1355,N_1486);
and U5998 (N_5998,N_301,N_938);
nor U5999 (N_5999,N_2220,N_87);
nor U6000 (N_6000,N_2134,N_2943);
xnor U6001 (N_6001,N_2581,N_136);
nor U6002 (N_6002,N_1803,N_656);
and U6003 (N_6003,N_2930,N_1353);
nand U6004 (N_6004,N_2480,N_1292);
and U6005 (N_6005,N_2120,N_1443);
or U6006 (N_6006,N_1148,N_22);
and U6007 (N_6007,N_1000,N_1414);
xor U6008 (N_6008,N_1713,N_233);
and U6009 (N_6009,N_1683,N_1355);
and U6010 (N_6010,N_492,N_2775);
xor U6011 (N_6011,N_237,N_70);
nand U6012 (N_6012,N_482,N_978);
nor U6013 (N_6013,N_1536,N_2369);
or U6014 (N_6014,N_1298,N_2115);
nor U6015 (N_6015,N_1161,N_916);
or U6016 (N_6016,N_1766,N_1072);
and U6017 (N_6017,N_784,N_742);
or U6018 (N_6018,N_2430,N_2332);
and U6019 (N_6019,N_352,N_1626);
or U6020 (N_6020,N_1786,N_484);
nor U6021 (N_6021,N_1823,N_612);
xnor U6022 (N_6022,N_322,N_1592);
nor U6023 (N_6023,N_1515,N_2005);
and U6024 (N_6024,N_2810,N_2519);
nor U6025 (N_6025,N_1196,N_1402);
nand U6026 (N_6026,N_864,N_1187);
or U6027 (N_6027,N_2624,N_2973);
nand U6028 (N_6028,N_2633,N_732);
nand U6029 (N_6029,N_845,N_853);
or U6030 (N_6030,N_2682,N_1941);
and U6031 (N_6031,N_2251,N_1274);
nor U6032 (N_6032,N_2232,N_1934);
or U6033 (N_6033,N_1284,N_881);
nor U6034 (N_6034,N_2646,N_2536);
nand U6035 (N_6035,N_1612,N_1083);
or U6036 (N_6036,N_367,N_684);
and U6037 (N_6037,N_2374,N_1913);
nor U6038 (N_6038,N_2837,N_458);
xnor U6039 (N_6039,N_1458,N_3085);
nand U6040 (N_6040,N_1738,N_893);
nand U6041 (N_6041,N_259,N_982);
and U6042 (N_6042,N_953,N_2623);
and U6043 (N_6043,N_1652,N_2690);
nand U6044 (N_6044,N_2149,N_433);
and U6045 (N_6045,N_1529,N_961);
or U6046 (N_6046,N_2966,N_2382);
or U6047 (N_6047,N_1361,N_631);
xor U6048 (N_6048,N_2945,N_1193);
or U6049 (N_6049,N_1404,N_914);
or U6050 (N_6050,N_1227,N_2446);
nor U6051 (N_6051,N_1092,N_1568);
and U6052 (N_6052,N_105,N_2767);
nand U6053 (N_6053,N_1492,N_1337);
nand U6054 (N_6054,N_3012,N_2294);
and U6055 (N_6055,N_1297,N_2668);
nand U6056 (N_6056,N_1322,N_3112);
or U6057 (N_6057,N_1137,N_2473);
nor U6058 (N_6058,N_964,N_2393);
or U6059 (N_6059,N_1775,N_2005);
nor U6060 (N_6060,N_1311,N_1133);
or U6061 (N_6061,N_2869,N_933);
and U6062 (N_6062,N_3095,N_325);
xor U6063 (N_6063,N_2115,N_1239);
nor U6064 (N_6064,N_35,N_1074);
nand U6065 (N_6065,N_2037,N_834);
or U6066 (N_6066,N_2822,N_696);
nand U6067 (N_6067,N_1839,N_1695);
nand U6068 (N_6068,N_497,N_1542);
or U6069 (N_6069,N_221,N_1525);
and U6070 (N_6070,N_2676,N_903);
or U6071 (N_6071,N_2740,N_139);
nor U6072 (N_6072,N_2905,N_763);
nand U6073 (N_6073,N_190,N_87);
or U6074 (N_6074,N_935,N_2400);
nor U6075 (N_6075,N_1698,N_724);
and U6076 (N_6076,N_2627,N_2666);
xor U6077 (N_6077,N_3122,N_2569);
or U6078 (N_6078,N_625,N_2027);
nand U6079 (N_6079,N_810,N_1214);
nand U6080 (N_6080,N_42,N_68);
and U6081 (N_6081,N_1760,N_2580);
xnor U6082 (N_6082,N_3116,N_268);
nor U6083 (N_6083,N_2074,N_22);
and U6084 (N_6084,N_448,N_2526);
nor U6085 (N_6085,N_1808,N_193);
or U6086 (N_6086,N_2506,N_1774);
nor U6087 (N_6087,N_1715,N_1762);
nand U6088 (N_6088,N_1844,N_2794);
nor U6089 (N_6089,N_2769,N_2763);
or U6090 (N_6090,N_1131,N_2663);
nand U6091 (N_6091,N_2633,N_2638);
nand U6092 (N_6092,N_2741,N_1249);
nor U6093 (N_6093,N_2448,N_1429);
and U6094 (N_6094,N_1664,N_3119);
xnor U6095 (N_6095,N_1386,N_964);
xor U6096 (N_6096,N_2206,N_292);
or U6097 (N_6097,N_914,N_531);
and U6098 (N_6098,N_2358,N_156);
nand U6099 (N_6099,N_236,N_1761);
and U6100 (N_6100,N_1268,N_2877);
nor U6101 (N_6101,N_1787,N_1280);
and U6102 (N_6102,N_2018,N_2296);
or U6103 (N_6103,N_357,N_1149);
nor U6104 (N_6104,N_557,N_2640);
or U6105 (N_6105,N_2015,N_2645);
xnor U6106 (N_6106,N_1764,N_1495);
nor U6107 (N_6107,N_2967,N_2222);
nand U6108 (N_6108,N_1801,N_864);
or U6109 (N_6109,N_2843,N_210);
nor U6110 (N_6110,N_2594,N_2607);
or U6111 (N_6111,N_2712,N_2931);
nand U6112 (N_6112,N_3021,N_1204);
nand U6113 (N_6113,N_1803,N_902);
nor U6114 (N_6114,N_1949,N_1666);
nor U6115 (N_6115,N_115,N_1940);
nor U6116 (N_6116,N_2845,N_2857);
nor U6117 (N_6117,N_1017,N_1353);
nand U6118 (N_6118,N_3076,N_3107);
xor U6119 (N_6119,N_2176,N_884);
or U6120 (N_6120,N_947,N_1285);
nor U6121 (N_6121,N_1404,N_781);
nand U6122 (N_6122,N_394,N_1224);
or U6123 (N_6123,N_3039,N_3026);
nor U6124 (N_6124,N_2533,N_2157);
and U6125 (N_6125,N_2406,N_2435);
nand U6126 (N_6126,N_1347,N_627);
nand U6127 (N_6127,N_895,N_367);
or U6128 (N_6128,N_2337,N_1189);
or U6129 (N_6129,N_2041,N_2721);
nor U6130 (N_6130,N_1335,N_949);
or U6131 (N_6131,N_2178,N_2511);
xnor U6132 (N_6132,N_1068,N_480);
or U6133 (N_6133,N_1268,N_1494);
nor U6134 (N_6134,N_3112,N_2610);
xnor U6135 (N_6135,N_2018,N_105);
nand U6136 (N_6136,N_1820,N_2947);
nor U6137 (N_6137,N_2791,N_1743);
and U6138 (N_6138,N_2686,N_425);
xor U6139 (N_6139,N_806,N_1704);
nand U6140 (N_6140,N_2509,N_14);
nor U6141 (N_6141,N_1952,N_3037);
nand U6142 (N_6142,N_864,N_415);
nor U6143 (N_6143,N_579,N_329);
or U6144 (N_6144,N_988,N_1195);
nand U6145 (N_6145,N_2433,N_106);
nor U6146 (N_6146,N_2842,N_1374);
and U6147 (N_6147,N_2407,N_447);
nor U6148 (N_6148,N_1982,N_2097);
or U6149 (N_6149,N_1809,N_2598);
nand U6150 (N_6150,N_1409,N_355);
or U6151 (N_6151,N_2801,N_167);
or U6152 (N_6152,N_269,N_829);
or U6153 (N_6153,N_2884,N_2819);
or U6154 (N_6154,N_1949,N_1751);
nor U6155 (N_6155,N_260,N_495);
nand U6156 (N_6156,N_2001,N_1108);
and U6157 (N_6157,N_1725,N_969);
or U6158 (N_6158,N_1533,N_1269);
nand U6159 (N_6159,N_149,N_1008);
nor U6160 (N_6160,N_3059,N_2353);
or U6161 (N_6161,N_2642,N_1021);
xor U6162 (N_6162,N_2729,N_1570);
nor U6163 (N_6163,N_595,N_2056);
nor U6164 (N_6164,N_2547,N_2413);
nand U6165 (N_6165,N_3120,N_2231);
or U6166 (N_6166,N_2339,N_3042);
or U6167 (N_6167,N_1133,N_3041);
or U6168 (N_6168,N_3073,N_988);
nand U6169 (N_6169,N_1906,N_682);
xor U6170 (N_6170,N_238,N_286);
nor U6171 (N_6171,N_654,N_2636);
and U6172 (N_6172,N_2905,N_1506);
nand U6173 (N_6173,N_1901,N_519);
or U6174 (N_6174,N_2181,N_2092);
nand U6175 (N_6175,N_2867,N_2973);
nand U6176 (N_6176,N_2937,N_936);
nand U6177 (N_6177,N_2052,N_2601);
or U6178 (N_6178,N_2562,N_2383);
nor U6179 (N_6179,N_2085,N_167);
nand U6180 (N_6180,N_1425,N_2962);
or U6181 (N_6181,N_1500,N_2619);
nor U6182 (N_6182,N_889,N_2210);
and U6183 (N_6183,N_2284,N_1401);
nor U6184 (N_6184,N_1913,N_1793);
or U6185 (N_6185,N_1091,N_294);
and U6186 (N_6186,N_1822,N_1798);
and U6187 (N_6187,N_1893,N_1973);
xor U6188 (N_6188,N_871,N_2111);
nor U6189 (N_6189,N_1641,N_961);
and U6190 (N_6190,N_290,N_924);
or U6191 (N_6191,N_2432,N_1162);
or U6192 (N_6192,N_2176,N_543);
and U6193 (N_6193,N_487,N_1768);
and U6194 (N_6194,N_2085,N_515);
nand U6195 (N_6195,N_2352,N_2343);
nand U6196 (N_6196,N_1949,N_1038);
nor U6197 (N_6197,N_1779,N_2629);
nor U6198 (N_6198,N_1014,N_2139);
and U6199 (N_6199,N_2235,N_489);
or U6200 (N_6200,N_2158,N_1363);
and U6201 (N_6201,N_1425,N_810);
nand U6202 (N_6202,N_2010,N_1960);
and U6203 (N_6203,N_2980,N_2418);
or U6204 (N_6204,N_1096,N_2296);
or U6205 (N_6205,N_2448,N_962);
xor U6206 (N_6206,N_2071,N_983);
and U6207 (N_6207,N_2338,N_3056);
and U6208 (N_6208,N_2725,N_3108);
nor U6209 (N_6209,N_217,N_547);
nand U6210 (N_6210,N_548,N_2550);
or U6211 (N_6211,N_2093,N_1037);
and U6212 (N_6212,N_801,N_2684);
and U6213 (N_6213,N_2222,N_1056);
nor U6214 (N_6214,N_2813,N_1439);
nor U6215 (N_6215,N_2657,N_2964);
nor U6216 (N_6216,N_399,N_2282);
or U6217 (N_6217,N_2210,N_670);
xnor U6218 (N_6218,N_2946,N_1092);
or U6219 (N_6219,N_2692,N_724);
nand U6220 (N_6220,N_243,N_2047);
and U6221 (N_6221,N_1550,N_554);
nand U6222 (N_6222,N_10,N_1691);
nor U6223 (N_6223,N_2422,N_1874);
or U6224 (N_6224,N_320,N_2178);
or U6225 (N_6225,N_1834,N_2047);
or U6226 (N_6226,N_1604,N_548);
and U6227 (N_6227,N_345,N_2643);
nand U6228 (N_6228,N_1865,N_1499);
and U6229 (N_6229,N_1399,N_954);
nand U6230 (N_6230,N_1948,N_2474);
or U6231 (N_6231,N_1922,N_3062);
or U6232 (N_6232,N_823,N_2170);
or U6233 (N_6233,N_1384,N_1716);
nand U6234 (N_6234,N_667,N_428);
xnor U6235 (N_6235,N_2953,N_2154);
nand U6236 (N_6236,N_1870,N_1587);
nor U6237 (N_6237,N_1627,N_890);
and U6238 (N_6238,N_1374,N_3064);
and U6239 (N_6239,N_1626,N_2537);
nand U6240 (N_6240,N_2670,N_1405);
nor U6241 (N_6241,N_273,N_2560);
and U6242 (N_6242,N_2073,N_1898);
and U6243 (N_6243,N_3083,N_921);
or U6244 (N_6244,N_615,N_1966);
nor U6245 (N_6245,N_2794,N_514);
and U6246 (N_6246,N_2073,N_1441);
or U6247 (N_6247,N_2442,N_977);
nor U6248 (N_6248,N_265,N_2204);
and U6249 (N_6249,N_2540,N_1920);
or U6250 (N_6250,N_4582,N_3630);
or U6251 (N_6251,N_5417,N_5766);
xnor U6252 (N_6252,N_3718,N_4701);
nor U6253 (N_6253,N_5716,N_4261);
nand U6254 (N_6254,N_5252,N_5150);
and U6255 (N_6255,N_5874,N_4783);
and U6256 (N_6256,N_6064,N_3629);
and U6257 (N_6257,N_3563,N_5425);
or U6258 (N_6258,N_5688,N_5893);
or U6259 (N_6259,N_6096,N_5611);
xnor U6260 (N_6260,N_3374,N_4080);
nor U6261 (N_6261,N_5929,N_3517);
or U6262 (N_6262,N_3420,N_5603);
nand U6263 (N_6263,N_5123,N_5590);
and U6264 (N_6264,N_5151,N_4415);
or U6265 (N_6265,N_5178,N_6032);
nand U6266 (N_6266,N_4916,N_4336);
or U6267 (N_6267,N_4233,N_5259);
xor U6268 (N_6268,N_5880,N_3156);
xnor U6269 (N_6269,N_5206,N_6238);
or U6270 (N_6270,N_5555,N_4899);
nor U6271 (N_6271,N_5162,N_4073);
nand U6272 (N_6272,N_4104,N_4259);
or U6273 (N_6273,N_5952,N_5209);
nand U6274 (N_6274,N_5888,N_3645);
and U6275 (N_6275,N_6118,N_3611);
nand U6276 (N_6276,N_4269,N_5413);
or U6277 (N_6277,N_3881,N_4043);
or U6278 (N_6278,N_5018,N_5816);
nor U6279 (N_6279,N_4301,N_4372);
nand U6280 (N_6280,N_5633,N_4252);
and U6281 (N_6281,N_5400,N_4587);
xnor U6282 (N_6282,N_5433,N_5134);
or U6283 (N_6283,N_5853,N_3448);
and U6284 (N_6284,N_4721,N_3543);
nor U6285 (N_6285,N_5080,N_4975);
or U6286 (N_6286,N_5357,N_3759);
or U6287 (N_6287,N_5600,N_5075);
nor U6288 (N_6288,N_4921,N_4468);
nand U6289 (N_6289,N_5138,N_5619);
nand U6290 (N_6290,N_3796,N_4840);
or U6291 (N_6291,N_5765,N_5902);
and U6292 (N_6292,N_3421,N_3625);
nand U6293 (N_6293,N_5191,N_5673);
nand U6294 (N_6294,N_5937,N_3486);
or U6295 (N_6295,N_3904,N_3149);
or U6296 (N_6296,N_5658,N_6139);
nor U6297 (N_6297,N_4948,N_4149);
or U6298 (N_6298,N_5592,N_3685);
nor U6299 (N_6299,N_4941,N_4381);
nand U6300 (N_6300,N_4809,N_4369);
nor U6301 (N_6301,N_4284,N_6062);
and U6302 (N_6302,N_6068,N_5833);
xor U6303 (N_6303,N_5015,N_3129);
nor U6304 (N_6304,N_4793,N_4990);
nor U6305 (N_6305,N_4691,N_5041);
and U6306 (N_6306,N_4098,N_5239);
xnor U6307 (N_6307,N_4495,N_5675);
and U6308 (N_6308,N_4623,N_4483);
nand U6309 (N_6309,N_3622,N_5589);
or U6310 (N_6310,N_4481,N_5728);
and U6311 (N_6311,N_6150,N_4199);
nand U6312 (N_6312,N_3277,N_4583);
or U6313 (N_6313,N_5900,N_4973);
and U6314 (N_6314,N_5883,N_3975);
or U6315 (N_6315,N_5468,N_4643);
nor U6316 (N_6316,N_5768,N_3273);
nor U6317 (N_6317,N_5480,N_3832);
and U6318 (N_6318,N_4334,N_5449);
or U6319 (N_6319,N_5612,N_3360);
nor U6320 (N_6320,N_5062,N_5756);
and U6321 (N_6321,N_4452,N_5793);
nand U6322 (N_6322,N_3481,N_3213);
nor U6323 (N_6323,N_3197,N_3280);
and U6324 (N_6324,N_6225,N_5613);
or U6325 (N_6325,N_6074,N_3690);
nor U6326 (N_6326,N_6015,N_5530);
nor U6327 (N_6327,N_4907,N_4477);
nor U6328 (N_6328,N_3684,N_5081);
nor U6329 (N_6329,N_5471,N_3480);
nand U6330 (N_6330,N_4656,N_4471);
nand U6331 (N_6331,N_3494,N_4548);
and U6332 (N_6332,N_6080,N_5367);
nand U6333 (N_6333,N_4472,N_6167);
or U6334 (N_6334,N_4271,N_3766);
or U6335 (N_6335,N_4052,N_5091);
nor U6336 (N_6336,N_6035,N_3815);
nand U6337 (N_6337,N_5634,N_5927);
nor U6338 (N_6338,N_4089,N_3900);
or U6339 (N_6339,N_5679,N_5414);
xor U6340 (N_6340,N_3362,N_5222);
and U6341 (N_6341,N_5648,N_6195);
nor U6342 (N_6342,N_3820,N_3949);
xor U6343 (N_6343,N_4242,N_4355);
nand U6344 (N_6344,N_5656,N_5050);
and U6345 (N_6345,N_6115,N_4824);
or U6346 (N_6346,N_3447,N_4856);
or U6347 (N_6347,N_4131,N_5840);
nor U6348 (N_6348,N_3653,N_4880);
or U6349 (N_6349,N_5059,N_3935);
xor U6350 (N_6350,N_5109,N_5243);
and U6351 (N_6351,N_5186,N_6149);
nor U6352 (N_6352,N_5052,N_5096);
nor U6353 (N_6353,N_4204,N_3222);
nand U6354 (N_6354,N_3206,N_5384);
nand U6355 (N_6355,N_3315,N_5821);
nor U6356 (N_6356,N_4298,N_4276);
nor U6357 (N_6357,N_5264,N_3751);
or U6358 (N_6358,N_3638,N_3310);
nor U6359 (N_6359,N_4039,N_4407);
and U6360 (N_6360,N_5415,N_3391);
nor U6361 (N_6361,N_6141,N_4597);
nand U6362 (N_6362,N_4215,N_6021);
nor U6363 (N_6363,N_5971,N_4771);
and U6364 (N_6364,N_3394,N_3670);
nor U6365 (N_6365,N_5301,N_4116);
nor U6366 (N_6366,N_5376,N_3999);
or U6367 (N_6367,N_5005,N_4475);
nand U6368 (N_6368,N_3363,N_3793);
and U6369 (N_6369,N_3728,N_4992);
and U6370 (N_6370,N_4041,N_4718);
and U6371 (N_6371,N_5334,N_4959);
or U6372 (N_6372,N_6114,N_5213);
or U6373 (N_6373,N_4685,N_5877);
nor U6374 (N_6374,N_3553,N_4222);
or U6375 (N_6375,N_5926,N_5175);
and U6376 (N_6376,N_4096,N_5047);
nor U6377 (N_6377,N_4191,N_4090);
or U6378 (N_6378,N_5056,N_5549);
or U6379 (N_6379,N_5529,N_3603);
nor U6380 (N_6380,N_3619,N_6174);
and U6381 (N_6381,N_4891,N_5278);
and U6382 (N_6382,N_4987,N_5390);
and U6383 (N_6383,N_5604,N_5408);
xnor U6384 (N_6384,N_5789,N_4711);
nand U6385 (N_6385,N_4379,N_6089);
xnor U6386 (N_6386,N_5636,N_5616);
nand U6387 (N_6387,N_5389,N_4885);
nor U6388 (N_6388,N_5442,N_4955);
and U6389 (N_6389,N_4665,N_3328);
nand U6390 (N_6390,N_4595,N_4779);
xnor U6391 (N_6391,N_6069,N_4217);
nor U6392 (N_6392,N_4561,N_3986);
xor U6393 (N_6393,N_5709,N_4299);
nor U6394 (N_6394,N_3242,N_4784);
nor U6395 (N_6395,N_6176,N_3381);
nand U6396 (N_6396,N_4945,N_5418);
nor U6397 (N_6397,N_4786,N_3926);
and U6398 (N_6398,N_3569,N_3698);
nand U6399 (N_6399,N_4974,N_5176);
nor U6400 (N_6400,N_4757,N_5446);
xnor U6401 (N_6401,N_5295,N_4581);
nor U6402 (N_6402,N_5095,N_3680);
or U6403 (N_6403,N_5657,N_5274);
and U6404 (N_6404,N_3623,N_6196);
or U6405 (N_6405,N_4105,N_4198);
nand U6406 (N_6406,N_4433,N_4040);
and U6407 (N_6407,N_3178,N_5492);
nor U6408 (N_6408,N_3706,N_6000);
or U6409 (N_6409,N_4487,N_6082);
nor U6410 (N_6410,N_4835,N_3595);
nand U6411 (N_6411,N_3550,N_3261);
nand U6412 (N_6412,N_5942,N_4063);
and U6413 (N_6413,N_5819,N_4796);
xor U6414 (N_6414,N_4730,N_5116);
or U6415 (N_6415,N_4640,N_3988);
nand U6416 (N_6416,N_4932,N_5683);
and U6417 (N_6417,N_5597,N_3584);
and U6418 (N_6418,N_4687,N_3410);
and U6419 (N_6419,N_3295,N_4056);
nand U6420 (N_6420,N_5411,N_3483);
and U6421 (N_6421,N_5375,N_3503);
xnor U6422 (N_6422,N_4200,N_4127);
xnor U6423 (N_6423,N_4702,N_5621);
nand U6424 (N_6424,N_5855,N_4659);
nor U6425 (N_6425,N_3231,N_5484);
nand U6426 (N_6426,N_3979,N_5294);
nand U6427 (N_6427,N_5806,N_5285);
and U6428 (N_6428,N_3216,N_4577);
nor U6429 (N_6429,N_3687,N_4494);
or U6430 (N_6430,N_3202,N_5614);
or U6431 (N_6431,N_5823,N_5280);
and U6432 (N_6432,N_3895,N_4270);
and U6433 (N_6433,N_4050,N_3225);
or U6434 (N_6434,N_3589,N_4406);
nor U6435 (N_6435,N_4574,N_5832);
nand U6436 (N_6436,N_6019,N_5824);
nand U6437 (N_6437,N_3604,N_5079);
and U6438 (N_6438,N_5754,N_5953);
or U6439 (N_6439,N_4862,N_4717);
and U6440 (N_6440,N_3205,N_5714);
nor U6441 (N_6441,N_3300,N_4123);
nor U6442 (N_6442,N_5216,N_5977);
nor U6443 (N_6443,N_4542,N_5579);
nor U6444 (N_6444,N_4906,N_4989);
or U6445 (N_6445,N_5131,N_3676);
nor U6446 (N_6446,N_4311,N_4257);
nand U6447 (N_6447,N_3914,N_4812);
nor U6448 (N_6448,N_3825,N_4136);
or U6449 (N_6449,N_3586,N_6065);
and U6450 (N_6450,N_3664,N_3554);
and U6451 (N_6451,N_5536,N_3739);
nor U6452 (N_6452,N_4053,N_4744);
or U6453 (N_6453,N_3239,N_3160);
xor U6454 (N_6454,N_4345,N_5179);
nand U6455 (N_6455,N_3588,N_4354);
and U6456 (N_6456,N_4283,N_3341);
xor U6457 (N_6457,N_4462,N_6144);
nor U6458 (N_6458,N_5758,N_4716);
and U6459 (N_6459,N_6148,N_5727);
or U6460 (N_6460,N_4174,N_4165);
xor U6461 (N_6461,N_5328,N_5598);
nand U6462 (N_6462,N_4361,N_5847);
nand U6463 (N_6463,N_3181,N_3865);
xor U6464 (N_6464,N_5525,N_3734);
or U6465 (N_6465,N_4003,N_3897);
nand U6466 (N_6466,N_5924,N_4175);
or U6467 (N_6467,N_3144,N_3972);
or U6468 (N_6468,N_6230,N_3203);
or U6469 (N_6469,N_4535,N_3937);
nand U6470 (N_6470,N_6161,N_5837);
or U6471 (N_6471,N_4129,N_3911);
nand U6472 (N_6472,N_3422,N_5201);
and U6473 (N_6473,N_3322,N_5661);
nor U6474 (N_6474,N_4814,N_4085);
nor U6475 (N_6475,N_5055,N_3722);
and U6476 (N_6476,N_4375,N_4313);
nand U6477 (N_6477,N_5784,N_3753);
and U6478 (N_6478,N_3971,N_5867);
xnor U6479 (N_6479,N_5310,N_4780);
nor U6480 (N_6480,N_4947,N_4344);
nor U6481 (N_6481,N_4450,N_3218);
xor U6482 (N_6482,N_5548,N_5732);
or U6483 (N_6483,N_3965,N_4719);
nand U6484 (N_6484,N_5583,N_6140);
or U6485 (N_6485,N_3343,N_4209);
nor U6486 (N_6486,N_3940,N_5996);
or U6487 (N_6487,N_3870,N_5038);
and U6488 (N_6488,N_3373,N_4273);
nor U6489 (N_6489,N_4310,N_5662);
and U6490 (N_6490,N_5368,N_4754);
or U6491 (N_6491,N_5354,N_4103);
nand U6492 (N_6492,N_4706,N_3204);
nor U6493 (N_6493,N_5308,N_3727);
and U6494 (N_6494,N_5042,N_5782);
nand U6495 (N_6495,N_5256,N_4571);
and U6496 (N_6496,N_3736,N_5581);
xnor U6497 (N_6497,N_4410,N_4739);
nand U6498 (N_6498,N_4058,N_4042);
or U6499 (N_6499,N_4759,N_3414);
nor U6500 (N_6500,N_5183,N_5118);
or U6501 (N_6501,N_4999,N_4338);
nor U6502 (N_6502,N_3590,N_6247);
nand U6503 (N_6503,N_4076,N_4505);
nor U6504 (N_6504,N_3379,N_4480);
and U6505 (N_6505,N_5298,N_4421);
xor U6506 (N_6506,N_6075,N_5170);
and U6507 (N_6507,N_3652,N_6116);
nor U6508 (N_6508,N_5469,N_3336);
and U6509 (N_6509,N_5448,N_5998);
nor U6510 (N_6510,N_4445,N_5940);
nor U6511 (N_6511,N_4950,N_5092);
nand U6512 (N_6512,N_5540,N_5029);
xnor U6513 (N_6513,N_4146,N_3763);
and U6514 (N_6514,N_5647,N_4876);
xor U6515 (N_6515,N_3529,N_6145);
nor U6516 (N_6516,N_5342,N_4898);
nand U6517 (N_6517,N_6037,N_4296);
or U6518 (N_6518,N_5521,N_4667);
and U6519 (N_6519,N_5761,N_5773);
nand U6520 (N_6520,N_3268,N_3806);
or U6521 (N_6521,N_5524,N_5211);
nor U6522 (N_6522,N_5160,N_5316);
and U6523 (N_6523,N_3839,N_5396);
xor U6524 (N_6524,N_4111,N_6111);
and U6525 (N_6525,N_3325,N_5801);
or U6526 (N_6526,N_4893,N_3666);
and U6527 (N_6527,N_3299,N_3817);
xor U6528 (N_6528,N_5775,N_4949);
xor U6529 (N_6529,N_5169,N_4446);
nand U6530 (N_6530,N_5786,N_3134);
xor U6531 (N_6531,N_4235,N_5273);
and U6532 (N_6532,N_4742,N_4680);
or U6533 (N_6533,N_6209,N_4061);
nand U6534 (N_6534,N_5866,N_3741);
or U6535 (N_6535,N_4015,N_5698);
nor U6536 (N_6536,N_3179,N_5682);
nor U6537 (N_6537,N_5393,N_4325);
nand U6538 (N_6538,N_3671,N_4476);
nand U6539 (N_6539,N_5649,N_5276);
nand U6540 (N_6540,N_4622,N_4218);
nand U6541 (N_6541,N_4486,N_4037);
nor U6542 (N_6542,N_4833,N_4021);
xnor U6543 (N_6543,N_6220,N_4887);
and U6544 (N_6544,N_4182,N_4456);
or U6545 (N_6545,N_4097,N_3473);
or U6546 (N_6546,N_4069,N_4618);
nand U6547 (N_6547,N_3318,N_4422);
nor U6548 (N_6548,N_5947,N_4335);
nor U6549 (N_6549,N_3861,N_4376);
and U6550 (N_6550,N_4006,N_6232);
and U6551 (N_6551,N_4366,N_5460);
nand U6552 (N_6552,N_4424,N_3397);
nor U6553 (N_6553,N_5102,N_3158);
and U6554 (N_6554,N_5128,N_3615);
nand U6555 (N_6555,N_5970,N_5802);
nand U6556 (N_6556,N_5043,N_5918);
nand U6557 (N_6557,N_6070,N_4557);
or U6558 (N_6558,N_5282,N_3361);
nand U6559 (N_6559,N_5496,N_5547);
and U6560 (N_6560,N_5190,N_3351);
and U6561 (N_6561,N_4364,N_6224);
nor U6562 (N_6562,N_3555,N_3678);
nor U6563 (N_6563,N_5336,N_4628);
xnor U6564 (N_6564,N_6119,N_4180);
xnor U6565 (N_6565,N_3393,N_4447);
or U6566 (N_6566,N_4638,N_3885);
nor U6567 (N_6567,N_6152,N_5810);
xor U6568 (N_6568,N_3518,N_4081);
and U6569 (N_6569,N_6029,N_3308);
or U6570 (N_6570,N_6007,N_3883);
nor U6571 (N_6571,N_3298,N_5572);
xor U6572 (N_6572,N_5622,N_5836);
or U6573 (N_6573,N_3462,N_5660);
nand U6574 (N_6574,N_3834,N_5518);
nor U6575 (N_6575,N_4135,N_3587);
or U6576 (N_6576,N_3848,N_3748);
or U6577 (N_6577,N_4297,N_5564);
xor U6578 (N_6578,N_6156,N_3335);
or U6579 (N_6579,N_3715,N_3990);
and U6580 (N_6580,N_5421,N_6242);
nand U6581 (N_6581,N_5694,N_4474);
and U6582 (N_6582,N_3235,N_4093);
nand U6583 (N_6583,N_3945,N_3578);
nand U6584 (N_6584,N_4869,N_4314);
nand U6585 (N_6585,N_6108,N_3176);
xnor U6586 (N_6586,N_5508,N_4842);
and U6587 (N_6587,N_4412,N_5987);
and U6588 (N_6588,N_4889,N_4092);
or U6589 (N_6589,N_6157,N_3211);
xor U6590 (N_6590,N_3974,N_3219);
or U6591 (N_6591,N_3789,N_5046);
and U6592 (N_6592,N_3531,N_6235);
and U6593 (N_6593,N_4646,N_5129);
nand U6594 (N_6594,N_4137,N_4114);
xor U6595 (N_6595,N_3628,N_4781);
and U6596 (N_6596,N_3783,N_5585);
and U6597 (N_6597,N_6077,N_5678);
and U6598 (N_6598,N_5881,N_5167);
and U6599 (N_6599,N_4629,N_3309);
and U6600 (N_6600,N_3755,N_3484);
nand U6601 (N_6601,N_5717,N_4892);
or U6602 (N_6602,N_3514,N_4119);
nand U6603 (N_6603,N_4747,N_3375);
nand U6604 (N_6604,N_3174,N_3857);
nor U6605 (N_6605,N_3286,N_5687);
xor U6606 (N_6606,N_3469,N_6155);
or U6607 (N_6607,N_5045,N_4173);
nand U6608 (N_6608,N_4288,N_3384);
or U6609 (N_6609,N_3145,N_3499);
nor U6610 (N_6610,N_5378,N_3417);
nand U6611 (N_6611,N_3632,N_4340);
xnor U6612 (N_6612,N_4225,N_3866);
nand U6613 (N_6613,N_4825,N_5692);
and U6614 (N_6614,N_4290,N_5260);
and U6615 (N_6615,N_4183,N_5083);
or U6616 (N_6616,N_6097,N_5182);
nor U6617 (N_6617,N_5475,N_3925);
or U6618 (N_6618,N_4491,N_3304);
xor U6619 (N_6619,N_3505,N_5197);
or U6620 (N_6620,N_4306,N_5731);
and U6621 (N_6621,N_3463,N_5035);
and U6622 (N_6622,N_3532,N_5110);
or U6623 (N_6623,N_3530,N_5820);
nor U6624 (N_6624,N_3657,N_6177);
and U6625 (N_6625,N_4467,N_4339);
nand U6626 (N_6626,N_4565,N_4749);
and U6627 (N_6627,N_4584,N_5556);
nand U6628 (N_6628,N_3407,N_5337);
nand U6629 (N_6629,N_3702,N_5204);
xnor U6630 (N_6630,N_3791,N_4304);
nor U6631 (N_6631,N_5745,N_3612);
and U6632 (N_6632,N_4437,N_5982);
nor U6633 (N_6633,N_3294,N_3616);
nor U6634 (N_6634,N_5371,N_4001);
and U6635 (N_6635,N_6214,N_5507);
nor U6636 (N_6636,N_5435,N_5355);
and U6637 (N_6637,N_4018,N_4509);
nor U6638 (N_6638,N_4260,N_5910);
nor U6639 (N_6639,N_3223,N_4291);
and U6640 (N_6640,N_4503,N_3468);
nor U6641 (N_6641,N_3608,N_3686);
nor U6642 (N_6642,N_5771,N_6244);
nor U6643 (N_6643,N_4884,N_4821);
or U6644 (N_6644,N_3559,N_4074);
or U6645 (N_6645,N_4351,N_5774);
xnor U6646 (N_6646,N_6004,N_3166);
and U6647 (N_6647,N_5168,N_4546);
and U6648 (N_6648,N_4036,N_5203);
and U6649 (N_6649,N_4167,N_4559);
xor U6650 (N_6650,N_3380,N_4024);
or U6651 (N_6651,N_5374,N_4541);
nor U6652 (N_6652,N_3512,N_4122);
nor U6653 (N_6653,N_4696,N_4926);
and U6654 (N_6654,N_4463,N_3187);
or U6655 (N_6655,N_5467,N_3546);
nand U6656 (N_6656,N_5114,N_3449);
or U6657 (N_6657,N_4172,N_4693);
nor U6658 (N_6658,N_5193,N_4432);
nand U6659 (N_6659,N_5778,N_5637);
and U6660 (N_6660,N_6093,N_3472);
nor U6661 (N_6661,N_3545,N_5711);
nor U6662 (N_6662,N_5314,N_3575);
nand U6663 (N_6663,N_4416,N_5356);
and U6664 (N_6664,N_5323,N_5088);
xnor U6665 (N_6665,N_5350,N_4930);
nand U6666 (N_6666,N_4874,N_4348);
and U6667 (N_6667,N_4658,N_5401);
or U6668 (N_6668,N_4620,N_4139);
xor U6669 (N_6669,N_5552,N_3436);
and U6670 (N_6670,N_5625,N_5788);
nand U6671 (N_6671,N_4594,N_4830);
nand U6672 (N_6672,N_4184,N_4820);
or U6673 (N_6673,N_5125,N_4212);
nor U6674 (N_6674,N_4019,N_6142);
or U6675 (N_6675,N_6005,N_4767);
xor U6676 (N_6676,N_5185,N_5228);
nand U6677 (N_6677,N_5930,N_4828);
nand U6678 (N_6678,N_3740,N_4777);
or U6679 (N_6679,N_5058,N_5398);
or U6680 (N_6680,N_4435,N_5587);
nor U6681 (N_6681,N_3229,N_5632);
nand U6682 (N_6682,N_3359,N_4841);
nor U6683 (N_6683,N_4329,N_3388);
or U6684 (N_6684,N_4698,N_3795);
xor U6685 (N_6685,N_5164,N_3913);
xnor U6686 (N_6686,N_5242,N_5751);
or U6687 (N_6687,N_3143,N_4797);
nor U6688 (N_6688,N_3833,N_5718);
nor U6689 (N_6689,N_3571,N_4558);
or U6690 (N_6690,N_5850,N_4357);
and U6691 (N_6691,N_5057,N_3334);
nand U6692 (N_6692,N_6044,N_3992);
nand U6693 (N_6693,N_6128,N_5137);
nand U6694 (N_6694,N_4872,N_4722);
nand U6695 (N_6695,N_5188,N_5764);
nor U6696 (N_6696,N_3402,N_5283);
or U6697 (N_6697,N_3398,N_3183);
or U6698 (N_6698,N_5886,N_5967);
or U6699 (N_6699,N_3989,N_4047);
and U6700 (N_6700,N_5112,N_5174);
nand U6701 (N_6701,N_5805,N_5962);
or U6702 (N_6702,N_5233,N_3226);
and U6703 (N_6703,N_5857,N_4922);
nand U6704 (N_6704,N_3390,N_3889);
nand U6705 (N_6705,N_3502,N_4265);
nor U6706 (N_6706,N_6010,N_4611);
and U6707 (N_6707,N_5030,N_3634);
nor U6708 (N_6708,N_4179,N_3962);
and U6709 (N_6709,N_4909,N_3928);
nor U6710 (N_6710,N_4489,N_5828);
nor U6711 (N_6711,N_4591,N_5245);
nor U6712 (N_6712,N_4946,N_5708);
and U6713 (N_6713,N_4258,N_4787);
and U6714 (N_6714,N_6090,N_5602);
and U6715 (N_6715,N_4312,N_3746);
or U6716 (N_6716,N_4762,N_4300);
or U6717 (N_6717,N_4391,N_6125);
nor U6718 (N_6718,N_4453,N_5402);
nor U6719 (N_6719,N_5346,N_5566);
or U6720 (N_6720,N_4378,N_5457);
nor U6721 (N_6721,N_3807,N_5723);
nor U6722 (N_6722,N_5307,N_6178);
or U6723 (N_6723,N_5325,N_3396);
nand U6724 (N_6724,N_4029,N_6181);
nor U6725 (N_6725,N_3279,N_3303);
xor U6726 (N_6726,N_3136,N_4399);
nor U6727 (N_6727,N_4838,N_3916);
nand U6728 (N_6728,N_4478,N_5423);
and U6729 (N_6729,N_4110,N_3663);
nor U6730 (N_6730,N_5726,N_3976);
or U6731 (N_6731,N_3830,N_4563);
nor U6732 (N_6732,N_5528,N_4633);
and U6733 (N_6733,N_4289,N_4617);
nand U6734 (N_6734,N_4025,N_3581);
xnor U6735 (N_6735,N_3408,N_3973);
nand U6736 (N_6736,N_4112,N_6016);
or U6737 (N_6737,N_5012,N_4550);
nor U6738 (N_6738,N_5236,N_5958);
nor U6739 (N_6739,N_3842,N_4991);
xor U6740 (N_6740,N_3931,N_3981);
and U6741 (N_6741,N_4804,N_3128);
or U6742 (N_6742,N_6135,N_4517);
xor U6743 (N_6743,N_5219,N_5997);
nand U6744 (N_6744,N_6237,N_5752);
or U6745 (N_6745,N_4536,N_3329);
nand U6746 (N_6746,N_5792,N_5905);
or U6747 (N_6747,N_3573,N_3159);
nor U6748 (N_6748,N_4692,N_4208);
or U6749 (N_6749,N_3301,N_5912);
and U6750 (N_6750,N_4836,N_5428);
and U6751 (N_6751,N_4769,N_5086);
or U6752 (N_6752,N_5734,N_5757);
and U6753 (N_6753,N_4728,N_4385);
xnor U6754 (N_6754,N_3557,N_6184);
or U6755 (N_6755,N_5101,N_3934);
or U6756 (N_6756,N_3260,N_5620);
or U6757 (N_6757,N_3535,N_3954);
nand U6758 (N_6758,N_4580,N_3327);
and U6759 (N_6759,N_4734,N_4621);
nand U6760 (N_6760,N_5434,N_4937);
nor U6761 (N_6761,N_6009,N_4908);
and U6762 (N_6762,N_5515,N_5161);
and U6763 (N_6763,N_4055,N_3923);
nand U6764 (N_6764,N_5322,N_5436);
nor U6765 (N_6765,N_4263,N_5842);
nand U6766 (N_6766,N_3765,N_5781);
nand U6767 (N_6767,N_5493,N_3792);
and U6768 (N_6768,N_5479,N_5399);
xnor U6769 (N_6769,N_3168,N_4928);
nand U6770 (N_6770,N_5104,N_6236);
nand U6771 (N_6771,N_4791,N_5385);
and U6772 (N_6772,N_3737,N_4349);
nand U6773 (N_6773,N_5016,N_5366);
nand U6774 (N_6774,N_3228,N_5247);
and U6775 (N_6775,N_4413,N_3906);
nand U6776 (N_6776,N_4046,N_6041);
nor U6777 (N_6777,N_5238,N_3192);
xor U6778 (N_6778,N_4171,N_3495);
nor U6779 (N_6779,N_4187,N_3233);
nor U6780 (N_6780,N_6109,N_4455);
or U6781 (N_6781,N_4652,N_5994);
nor U6782 (N_6782,N_4682,N_3844);
and U6783 (N_6783,N_5643,N_6223);
nor U6784 (N_6784,N_4178,N_4294);
nand U6785 (N_6785,N_5068,N_5753);
or U6786 (N_6786,N_5060,N_5935);
nor U6787 (N_6787,N_5192,N_3403);
xnor U6788 (N_6788,N_5652,N_4551);
and U6789 (N_6789,N_5955,N_3921);
nor U6790 (N_6790,N_3852,N_5470);
or U6791 (N_6791,N_3491,N_3292);
and U6792 (N_6792,N_4250,N_3266);
or U6793 (N_6793,N_4256,N_4027);
nor U6794 (N_6794,N_3246,N_6104);
nor U6795 (N_6795,N_5650,N_4126);
nand U6796 (N_6796,N_3501,N_5318);
and U6797 (N_6797,N_3668,N_3259);
or U6798 (N_6798,N_4134,N_4902);
nand U6799 (N_6799,N_4847,N_4493);
nor U6800 (N_6800,N_5826,N_5037);
and U6801 (N_6801,N_5576,N_6056);
nand U6802 (N_6802,N_4639,N_4157);
or U6803 (N_6803,N_6098,N_3406);
xor U6804 (N_6804,N_4868,N_4848);
or U6805 (N_6805,N_4210,N_5154);
or U6806 (N_6806,N_6205,N_5815);
or U6807 (N_6807,N_5706,N_4277);
or U6808 (N_6808,N_4619,N_3660);
nor U6809 (N_6809,N_6023,N_6031);
and U6810 (N_6810,N_6083,N_3465);
xor U6811 (N_6811,N_6239,N_3526);
nor U6812 (N_6812,N_4994,N_5431);
nor U6813 (N_6813,N_5527,N_5340);
nand U6814 (N_6814,N_3790,N_5214);
nand U6815 (N_6815,N_5606,N_4590);
nor U6816 (N_6816,N_5800,N_5416);
or U6817 (N_6817,N_3441,N_4935);
nand U6818 (N_6818,N_3855,N_3860);
nand U6819 (N_6819,N_4913,N_4470);
nand U6820 (N_6820,N_4274,N_5105);
or U6821 (N_6821,N_3283,N_4578);
nand U6822 (N_6822,N_4850,N_5149);
nand U6823 (N_6823,N_5920,N_4206);
and U6824 (N_6824,N_5562,N_5184);
or U6825 (N_6825,N_5713,N_3661);
nand U6826 (N_6826,N_5007,N_6162);
nand U6827 (N_6827,N_4384,N_3551);
and U6828 (N_6828,N_3528,N_5710);
nand U6829 (N_6829,N_4293,N_5253);
xor U6830 (N_6830,N_3797,N_5651);
nand U6831 (N_6831,N_4464,N_3428);
and U6832 (N_6832,N_4013,N_5729);
nand U6833 (N_6833,N_3800,N_4323);
nand U6834 (N_6834,N_5873,N_5404);
nand U6835 (N_6835,N_3679,N_5427);
nor U6836 (N_6836,N_6231,N_3370);
xor U6837 (N_6837,N_5946,N_4512);
nor U6838 (N_6838,N_3324,N_5825);
or U6839 (N_6839,N_5309,N_3966);
nor U6840 (N_6840,N_5473,N_4995);
nand U6841 (N_6841,N_5780,N_3750);
nor U6842 (N_6842,N_5258,N_4726);
or U6843 (N_6843,N_3803,N_3352);
nand U6844 (N_6844,N_4863,N_3274);
nand U6845 (N_6845,N_5671,N_4390);
and U6846 (N_6846,N_4854,N_5142);
nor U6847 (N_6847,N_3568,N_4967);
and U6848 (N_6848,N_3654,N_5730);
or U6849 (N_6849,N_5372,N_5445);
and U6850 (N_6850,N_3756,N_4065);
nand U6851 (N_6851,N_6129,N_3243);
and U6852 (N_6852,N_5133,N_4855);
nand U6853 (N_6853,N_4799,N_4570);
nor U6854 (N_6854,N_4121,N_4232);
and U6855 (N_6855,N_4094,N_4164);
nand U6856 (N_6856,N_5653,N_4608);
xnor U6857 (N_6857,N_5856,N_3726);
nor U6858 (N_6858,N_5290,N_5969);
xor U6859 (N_6859,N_5028,N_3354);
and U6860 (N_6860,N_5237,N_4158);
nor U6861 (N_6861,N_5573,N_4226);
xor U6862 (N_6862,N_4508,N_6011);
and U6863 (N_6863,N_3985,N_4418);
xor U6864 (N_6864,N_5317,N_5218);
and U6865 (N_6865,N_4156,N_6147);
and U6866 (N_6866,N_3620,N_3998);
and U6867 (N_6867,N_5642,N_4520);
and U6868 (N_6868,N_5699,N_3907);
or U6869 (N_6869,N_4923,N_3153);
nand U6870 (N_6870,N_4244,N_3614);
or U6871 (N_6871,N_5458,N_3271);
and U6872 (N_6872,N_5979,N_6226);
nor U6873 (N_6873,N_5070,N_4572);
and U6874 (N_6874,N_4484,N_5440);
xor U6875 (N_6875,N_6133,N_3709);
xnor U6876 (N_6876,N_3689,N_3644);
nor U6877 (N_6877,N_6246,N_4279);
nand U6878 (N_6878,N_5235,N_4202);
nor U6879 (N_6879,N_4560,N_4353);
and U6880 (N_6880,N_3459,N_3650);
or U6881 (N_6881,N_3513,N_5158);
xor U6882 (N_6882,N_5501,N_4579);
or U6883 (N_6883,N_4246,N_5978);
and U6884 (N_6884,N_5797,N_5510);
and U6885 (N_6885,N_4924,N_4568);
and U6886 (N_6886,N_4857,N_4588);
nand U6887 (N_6887,N_3943,N_4940);
xnor U6888 (N_6888,N_3701,N_3488);
and U6889 (N_6889,N_4161,N_3209);
or U6890 (N_6890,N_5522,N_3314);
nand U6891 (N_6891,N_3941,N_5439);
and U6892 (N_6892,N_6165,N_4573);
nor U6893 (N_6893,N_4753,N_4943);
or U6894 (N_6894,N_3912,N_5450);
nor U6895 (N_6895,N_6216,N_4231);
or U6896 (N_6896,N_5831,N_5738);
nor U6897 (N_6897,N_4197,N_5438);
and U6898 (N_6898,N_3383,N_4883);
nand U6899 (N_6899,N_4441,N_5747);
nor U6900 (N_6900,N_6057,N_5351);
nand U6901 (N_6901,N_6197,N_3533);
and U6902 (N_6902,N_4811,N_3932);
xor U6903 (N_6903,N_5869,N_4326);
or U6904 (N_6904,N_6169,N_6143);
xnor U6905 (N_6905,N_4816,N_3665);
xnor U6906 (N_6906,N_6101,N_5755);
and U6907 (N_6907,N_4374,N_3157);
xor U6908 (N_6908,N_5224,N_6212);
or U6909 (N_6909,N_3576,N_5004);
and U6910 (N_6910,N_5759,N_5147);
and U6911 (N_6911,N_5139,N_5495);
and U6912 (N_6912,N_4014,N_4895);
nand U6913 (N_6913,N_5380,N_6079);
and U6914 (N_6914,N_5938,N_5365);
nand U6915 (N_6915,N_3592,N_4566);
nor U6916 (N_6916,N_5406,N_5945);
nand U6917 (N_6917,N_3577,N_5344);
nand U6918 (N_6918,N_5181,N_3313);
or U6919 (N_6919,N_3182,N_4914);
nand U6920 (N_6920,N_4382,N_4095);
nand U6921 (N_6921,N_4818,N_4528);
nor U6922 (N_6922,N_3321,N_3667);
and U6923 (N_6923,N_4223,N_3593);
or U6924 (N_6924,N_3582,N_5506);
or U6925 (N_6925,N_4020,N_4253);
xor U6926 (N_6926,N_5791,N_3700);
or U6927 (N_6927,N_5610,N_3311);
or U6928 (N_6928,N_4772,N_5361);
xnor U6929 (N_6929,N_5770,N_5878);
nand U6930 (N_6930,N_5230,N_6027);
xnor U6931 (N_6931,N_3710,N_5550);
xnor U6932 (N_6932,N_6240,N_3720);
nor U6933 (N_6933,N_5574,N_3154);
nor U6934 (N_6934,N_6110,N_4449);
or U6935 (N_6935,N_3996,N_3511);
xnor U6936 (N_6936,N_3255,N_4125);
or U6937 (N_6937,N_5956,N_4031);
and U6938 (N_6938,N_3640,N_5577);
xnor U6939 (N_6939,N_6172,N_4281);
nor U6940 (N_6940,N_3598,N_5922);
nor U6941 (N_6941,N_4538,N_5036);
nand U6942 (N_6942,N_3438,N_5386);
xor U6943 (N_6943,N_5321,N_4091);
or U6944 (N_6944,N_5943,N_4396);
nor U6945 (N_6945,N_4534,N_4832);
and U6946 (N_6946,N_5639,N_4066);
nand U6947 (N_6947,N_4341,N_5627);
nor U6948 (N_6948,N_5631,N_5082);
or U6949 (N_6949,N_3682,N_5512);
xor U6950 (N_6950,N_5672,N_5394);
and U6951 (N_6951,N_6086,N_4363);
and U6952 (N_6952,N_4613,N_4873);
or U6953 (N_6953,N_5067,N_3331);
or U6954 (N_6954,N_3752,N_5241);
or U6955 (N_6955,N_4980,N_3357);
nand U6956 (N_6956,N_4272,N_6248);
and U6957 (N_6957,N_6036,N_4022);
nand U6958 (N_6958,N_5272,N_4752);
nor U6959 (N_6959,N_5093,N_3958);
and U6960 (N_6960,N_6117,N_5240);
nor U6961 (N_6961,N_4634,N_4106);
and U6962 (N_6962,N_5119,N_5960);
or U6963 (N_6963,N_5255,N_3782);
and U6964 (N_6964,N_4589,N_4330);
or U6965 (N_6965,N_5595,N_5951);
nand U6966 (N_6966,N_5868,N_5249);
nand U6967 (N_6967,N_4844,N_4423);
or U6968 (N_6968,N_3627,N_4084);
and U6969 (N_6969,N_5335,N_4420);
nand U6970 (N_6970,N_5397,N_5263);
or U6971 (N_6971,N_4181,N_5049);
or U6972 (N_6972,N_3867,N_3544);
or U6973 (N_6973,N_6229,N_6055);
nand U6974 (N_6974,N_3135,N_3610);
and U6975 (N_6975,N_5305,N_3489);
nor U6976 (N_6976,N_6121,N_5807);
or U6977 (N_6977,N_5884,N_4782);
xor U6978 (N_6978,N_3355,N_3658);
nand U6979 (N_6979,N_4768,N_6207);
nand U6980 (N_6980,N_3345,N_3193);
nand U6981 (N_6981,N_4683,N_5663);
nor U6982 (N_6982,N_3950,N_5303);
xnor U6983 (N_6983,N_5670,N_4359);
nand U6984 (N_6984,N_4641,N_4408);
nand U6985 (N_6985,N_3836,N_4562);
nor U6986 (N_6986,N_5388,N_5968);
nand U6987 (N_6987,N_5538,N_6073);
or U6988 (N_6988,N_5106,N_6175);
nand U6989 (N_6989,N_3453,N_3471);
or U6990 (N_6990,N_4676,N_4033);
nand U6991 (N_6991,N_5039,N_3778);
nor U6992 (N_6992,N_3942,N_4115);
nor U6993 (N_6993,N_5363,N_4030);
xnor U6994 (N_6994,N_6025,N_5911);
nor U6995 (N_6995,N_5795,N_4498);
nand U6996 (N_6996,N_5531,N_3522);
nor U6997 (N_6997,N_4800,N_4649);
nor U6998 (N_6998,N_3147,N_3460);
nor U6999 (N_6999,N_5014,N_5292);
or U7000 (N_7000,N_5140,N_5013);
nand U7001 (N_7001,N_5229,N_4278);
nor U7002 (N_7002,N_5261,N_6017);
nor U7003 (N_7003,N_5914,N_5432);
xnor U7004 (N_7004,N_5769,N_5127);
or U7005 (N_7005,N_3856,N_5596);
nand U7006 (N_7006,N_5299,N_5934);
nand U7007 (N_7007,N_4079,N_3880);
or U7008 (N_7008,N_6053,N_3850);
and U7009 (N_7009,N_5410,N_3146);
or U7010 (N_7010,N_5580,N_3170);
or U7011 (N_7011,N_4712,N_5568);
and U7012 (N_7012,N_4107,N_4805);
or U7013 (N_7013,N_3378,N_3464);
nor U7014 (N_7014,N_3191,N_3419);
nand U7015 (N_7015,N_4317,N_5347);
nor U7016 (N_7016,N_4228,N_3186);
and U7017 (N_7017,N_4624,N_5132);
or U7018 (N_7018,N_4988,N_4078);
xor U7019 (N_7019,N_3199,N_3892);
xor U7020 (N_7020,N_3415,N_3184);
nand U7021 (N_7021,N_5000,N_4694);
and U7022 (N_7022,N_5875,N_5919);
or U7023 (N_7023,N_5921,N_3493);
nand U7024 (N_7024,N_3548,N_3626);
nand U7025 (N_7025,N_3201,N_4688);
or U7026 (N_7026,N_5684,N_3977);
nand U7027 (N_7027,N_4343,N_4843);
and U7028 (N_7028,N_6188,N_4650);
nand U7029 (N_7029,N_5700,N_3456);
and U7030 (N_7030,N_5514,N_6200);
or U7031 (N_7031,N_4370,N_5407);
or U7032 (N_7032,N_5560,N_3691);
or U7033 (N_7033,N_5477,N_6233);
or U7034 (N_7034,N_3240,N_4230);
nor U7035 (N_7035,N_4601,N_4120);
nand U7036 (N_7036,N_5094,N_3779);
or U7037 (N_7037,N_4068,N_4501);
and U7038 (N_7038,N_3258,N_4707);
nand U7039 (N_7039,N_5664,N_3429);
nor U7040 (N_7040,N_4743,N_4846);
or U7041 (N_7041,N_3878,N_5895);
or U7042 (N_7042,N_3358,N_5849);
nor U7043 (N_7043,N_5453,N_4077);
nor U7044 (N_7044,N_4829,N_3451);
and U7045 (N_7045,N_5811,N_4185);
and U7046 (N_7046,N_3542,N_5145);
nor U7047 (N_7047,N_4996,N_6151);
xor U7048 (N_7048,N_5640,N_3677);
nor U7049 (N_7049,N_6189,N_3859);
xor U7050 (N_7050,N_4545,N_5787);
xor U7051 (N_7051,N_6076,N_3655);
or U7052 (N_7052,N_3194,N_4813);
nand U7053 (N_7053,N_3828,N_4496);
nor U7054 (N_7054,N_3829,N_3326);
nand U7055 (N_7055,N_5084,N_3561);
xnor U7056 (N_7056,N_5377,N_5459);
nand U7057 (N_7057,N_3450,N_3580);
and U7058 (N_7058,N_6186,N_4933);
xnor U7059 (N_7059,N_4879,N_4083);
and U7060 (N_7060,N_5845,N_3173);
or U7061 (N_7061,N_3647,N_4012);
nand U7062 (N_7062,N_4352,N_5776);
nand U7063 (N_7063,N_3635,N_3694);
or U7064 (N_7064,N_5227,N_4411);
xnor U7065 (N_7065,N_4839,N_4555);
and U7066 (N_7066,N_4637,N_4993);
nor U7067 (N_7067,N_4731,N_5157);
and U7068 (N_7068,N_3487,N_5899);
nor U7069 (N_7069,N_5383,N_5744);
nand U7070 (N_7070,N_3431,N_4117);
and U7071 (N_7071,N_3552,N_4100);
and U7072 (N_7072,N_3939,N_3307);
nor U7073 (N_7073,N_6249,N_5983);
nand U7074 (N_7074,N_3845,N_3401);
and U7075 (N_7075,N_5879,N_4044);
xnor U7076 (N_7076,N_3920,N_4492);
xor U7077 (N_7077,N_5557,N_3248);
and U7078 (N_7078,N_3411,N_4166);
or U7079 (N_7079,N_4715,N_5011);
nor U7080 (N_7080,N_3337,N_3320);
nor U7081 (N_7081,N_3887,N_3585);
nor U7082 (N_7082,N_5628,N_3781);
nor U7083 (N_7083,N_3346,N_4750);
and U7084 (N_7084,N_3479,N_4466);
and U7085 (N_7085,N_4521,N_5171);
xnor U7086 (N_7086,N_6112,N_5194);
nor U7087 (N_7087,N_6078,N_3400);
or U7088 (N_7088,N_4513,N_3523);
nor U7089 (N_7089,N_4194,N_5499);
and U7090 (N_7090,N_3762,N_6061);
xor U7091 (N_7091,N_3492,N_5291);
and U7092 (N_7092,N_5689,N_3980);
and U7093 (N_7093,N_4602,N_4826);
nor U7094 (N_7094,N_3637,N_4064);
nand U7095 (N_7095,N_6173,N_3284);
and U7096 (N_7096,N_3922,N_4510);
nand U7097 (N_7097,N_5593,N_3938);
nand U7098 (N_7098,N_4404,N_3822);
or U7099 (N_7099,N_5455,N_3873);
nor U7100 (N_7100,N_5313,N_4490);
and U7101 (N_7101,N_3963,N_5044);
nor U7102 (N_7102,N_4245,N_3607);
nand U7103 (N_7103,N_5017,N_4795);
nand U7104 (N_7104,N_3217,N_4237);
and U7105 (N_7105,N_4007,N_3412);
nor U7106 (N_7106,N_4853,N_5767);
nand U7107 (N_7107,N_3386,N_6132);
or U7108 (N_7108,N_4927,N_4275);
nor U7109 (N_7109,N_3744,N_3843);
or U7110 (N_7110,N_3387,N_6183);
or U7111 (N_7111,N_3238,N_5870);
nor U7112 (N_7112,N_4051,N_3621);
and U7113 (N_7113,N_3167,N_6067);
or U7114 (N_7114,N_3455,N_5533);
or U7115 (N_7115,N_3743,N_3814);
nand U7116 (N_7116,N_3951,N_6159);
nand U7117 (N_7117,N_5992,N_3399);
nor U7118 (N_7118,N_5338,N_3810);
and U7119 (N_7119,N_3264,N_5205);
nor U7120 (N_7120,N_6234,N_4049);
nand U7121 (N_7121,N_6038,N_3639);
xnor U7122 (N_7122,N_4234,N_5288);
xnor U7123 (N_7123,N_3899,N_5494);
nand U7124 (N_7124,N_5424,N_3983);
nand U7125 (N_7125,N_5463,N_3567);
or U7126 (N_7126,N_6095,N_5520);
or U7127 (N_7127,N_4738,N_5069);
xnor U7128 (N_7128,N_6024,N_3696);
and U7129 (N_7129,N_4302,N_5327);
nand U7130 (N_7130,N_3767,N_4801);
xnor U7131 (N_7131,N_3827,N_5854);
nand U7132 (N_7132,N_4674,N_3253);
and U7133 (N_7133,N_3440,N_4009);
and U7134 (N_7134,N_5173,N_3267);
nand U7135 (N_7135,N_5076,N_3991);
xor U7136 (N_7136,N_5511,N_3754);
nor U7137 (N_7137,N_3884,N_4207);
nand U7138 (N_7138,N_5545,N_3742);
xor U7139 (N_7139,N_3995,N_5490);
nor U7140 (N_7140,N_4356,N_5936);
nand U7141 (N_7141,N_4666,N_6099);
nand U7142 (N_7142,N_5554,N_3212);
or U7143 (N_7143,N_6217,N_4867);
xnor U7144 (N_7144,N_5244,N_5108);
or U7145 (N_7145,N_5601,N_4729);
nand U7146 (N_7146,N_5324,N_3365);
nor U7147 (N_7147,N_3385,N_5443);
and U7148 (N_7148,N_3214,N_4377);
and U7149 (N_7149,N_3882,N_4479);
and U7150 (N_7150,N_4960,N_4875);
and U7151 (N_7151,N_4699,N_4155);
and U7152 (N_7152,N_5733,N_4186);
nor U7153 (N_7153,N_5551,N_5326);
or U7154 (N_7154,N_5712,N_4526);
nor U7155 (N_7155,N_4038,N_3705);
and U7156 (N_7156,N_3692,N_6071);
nor U7157 (N_7157,N_6127,N_4414);
nand U7158 (N_7158,N_3443,N_5482);
nor U7159 (N_7159,N_4213,N_5217);
and U7160 (N_7160,N_5973,N_4647);
xor U7161 (N_7161,N_5674,N_3224);
or U7162 (N_7162,N_5491,N_3139);
or U7163 (N_7163,N_5741,N_4956);
nand U7164 (N_7164,N_5208,N_5097);
nand U7165 (N_7165,N_5991,N_4248);
nor U7166 (N_7166,N_4319,N_3729);
nand U7167 (N_7167,N_4789,N_3858);
nand U7168 (N_7168,N_5705,N_5743);
nor U7169 (N_7169,N_3747,N_4522);
nand U7170 (N_7170,N_3252,N_5523);
and U7171 (N_7171,N_4169,N_3367);
or U7172 (N_7172,N_5472,N_4671);
and U7173 (N_7173,N_3872,N_5841);
nand U7174 (N_7174,N_5629,N_5680);
xnor U7175 (N_7175,N_6012,N_3446);
and U7176 (N_7176,N_5961,N_5333);
nor U7177 (N_7177,N_3190,N_5681);
nand U7178 (N_7178,N_6126,N_3583);
and U7179 (N_7179,N_3774,N_6058);
nand U7180 (N_7180,N_3846,N_3952);
nor U7181 (N_7181,N_4434,N_3776);
and U7182 (N_7182,N_5202,N_3161);
and U7183 (N_7183,N_4392,N_5882);
nor U7184 (N_7184,N_5859,N_5267);
and U7185 (N_7185,N_3738,N_3894);
nand U7186 (N_7186,N_3293,N_3933);
or U7187 (N_7187,N_4890,N_3785);
nand U7188 (N_7188,N_3376,N_6008);
and U7189 (N_7189,N_5198,N_4219);
or U7190 (N_7190,N_4221,N_3725);
and U7191 (N_7191,N_3982,N_5546);
and U7192 (N_7192,N_5231,N_4417);
nand U7193 (N_7193,N_4901,N_5265);
and U7194 (N_7194,N_4845,N_4554);
and U7195 (N_7195,N_4144,N_4439);
or U7196 (N_7196,N_4894,N_3348);
and U7197 (N_7197,N_3272,N_6138);
nand U7198 (N_7198,N_3338,N_5465);
and U7199 (N_7199,N_4976,N_4985);
nor U7200 (N_7200,N_5563,N_6107);
or U7201 (N_7201,N_4151,N_4625);
or U7202 (N_7202,N_4075,N_5829);
nand U7203 (N_7203,N_4241,N_4262);
nand U7204 (N_7204,N_6120,N_5685);
and U7205 (N_7205,N_4997,N_4032);
and U7206 (N_7206,N_3564,N_5925);
or U7207 (N_7207,N_6094,N_5848);
nor U7208 (N_7208,N_4350,N_3648);
or U7209 (N_7209,N_4761,N_4939);
nand U7210 (N_7210,N_4017,N_3306);
nand U7211 (N_7211,N_4748,N_5122);
xor U7212 (N_7212,N_6154,N_4429);
nand U7213 (N_7213,N_5107,N_4977);
and U7214 (N_7214,N_5159,N_4428);
or U7215 (N_7215,N_4607,N_5437);
and U7216 (N_7216,N_6194,N_5027);
nor U7217 (N_7217,N_5395,N_4827);
or U7218 (N_7218,N_5248,N_4109);
or U7219 (N_7219,N_4383,N_4224);
and U7220 (N_7220,N_4653,N_4942);
and U7221 (N_7221,N_6003,N_4442);
or U7222 (N_7222,N_4807,N_5901);
and U7223 (N_7223,N_3142,N_6215);
nand U7224 (N_7224,N_4147,N_4604);
and U7225 (N_7225,N_5024,N_3478);
nor U7226 (N_7226,N_6245,N_6203);
or U7227 (N_7227,N_5691,N_3200);
and U7228 (N_7228,N_4168,N_4527);
or U7229 (N_7229,N_6124,N_3642);
and U7230 (N_7230,N_4368,N_3333);
or U7231 (N_7231,N_4938,N_5115);
nor U7232 (N_7232,N_4765,N_4426);
nand U7233 (N_7233,N_4405,N_5071);
nand U7234 (N_7234,N_6213,N_6081);
nand U7235 (N_7235,N_6063,N_6088);
nand U7236 (N_7236,N_5485,N_4531);
and U7237 (N_7237,N_4860,N_5422);
and U7238 (N_7238,N_5320,N_3175);
or U7239 (N_7239,N_5279,N_4708);
or U7240 (N_7240,N_3234,N_3432);
or U7241 (N_7241,N_4267,N_3801);
nor U7242 (N_7242,N_5074,N_3330);
and U7243 (N_7243,N_4929,N_3656);
nand U7244 (N_7244,N_5739,N_4523);
xor U7245 (N_7245,N_4529,N_5655);
xor U7246 (N_7246,N_4981,N_3955);
nor U7247 (N_7247,N_5999,N_3509);
nor U7248 (N_7248,N_5266,N_3994);
and U7249 (N_7249,N_3141,N_4430);
nor U7250 (N_7250,N_4148,N_4254);
nor U7251 (N_7251,N_4953,N_5897);
or U7252 (N_7252,N_4143,N_3901);
or U7253 (N_7253,N_5117,N_5737);
or U7254 (N_7254,N_4240,N_5623);
and U7255 (N_7255,N_5087,N_3461);
or U7256 (N_7256,N_4704,N_5257);
or U7257 (N_7257,N_4684,N_4870);
nand U7258 (N_7258,N_3269,N_4910);
nor U7259 (N_7259,N_3208,N_3675);
or U7260 (N_7260,N_4530,N_5827);
or U7261 (N_7261,N_4287,N_3853);
nand U7262 (N_7262,N_4905,N_6046);
nand U7263 (N_7263,N_6166,N_6048);
nand U7264 (N_7264,N_5331,N_3319);
xnor U7265 (N_7265,N_5503,N_4227);
nor U7266 (N_7266,N_4725,N_6028);
and U7267 (N_7267,N_4861,N_4865);
or U7268 (N_7268,N_3445,N_5539);
and U7269 (N_7269,N_6227,N_4010);
nor U7270 (N_7270,N_6072,N_5441);
xor U7271 (N_7271,N_4458,N_4745);
nand U7272 (N_7272,N_3875,N_4788);
and U7273 (N_7273,N_5349,N_3948);
and U7274 (N_7274,N_3804,N_5165);
and U7275 (N_7275,N_5502,N_3171);
nor U7276 (N_7276,N_5690,N_5779);
or U7277 (N_7277,N_4539,N_3257);
nor U7278 (N_7278,N_3256,N_3188);
nand U7279 (N_7279,N_4142,N_3332);
nand U7280 (N_7280,N_3305,N_3716);
nor U7281 (N_7281,N_5760,N_5941);
or U7282 (N_7282,N_6164,N_5607);
nor U7283 (N_7283,N_4454,N_4766);
nand U7284 (N_7284,N_5669,N_4651);
nor U7285 (N_7285,N_4236,N_4598);
and U7286 (N_7286,N_3594,N_5565);
or U7287 (N_7287,N_5156,N_4386);
and U7288 (N_7288,N_4059,N_3347);
or U7289 (N_7289,N_5569,N_3944);
and U7290 (N_7290,N_5269,N_4709);
xnor U7291 (N_7291,N_5409,N_4362);
nor U7292 (N_7292,N_3405,N_5293);
or U7293 (N_7293,N_3717,N_6199);
and U7294 (N_7294,N_3960,N_6171);
nand U7295 (N_7295,N_6187,N_5250);
or U7296 (N_7296,N_4984,N_3643);
and U7297 (N_7297,N_5099,N_5234);
xnor U7298 (N_7298,N_5120,N_4177);
nand U7299 (N_7299,N_3703,N_5898);
nor U7300 (N_7300,N_5950,N_5025);
nand U7301 (N_7301,N_4954,N_3162);
or U7302 (N_7302,N_5861,N_4163);
and U7303 (N_7303,N_6168,N_4400);
nor U7304 (N_7304,N_5750,N_3968);
xor U7305 (N_7305,N_4307,N_3624);
and U7306 (N_7306,N_6052,N_4778);
and U7307 (N_7307,N_3835,N_6087);
and U7308 (N_7308,N_4626,N_3547);
nand U7309 (N_7309,N_4264,N_3771);
nand U7310 (N_7310,N_3163,N_3477);
and U7311 (N_7311,N_4575,N_4342);
nor U7312 (N_7312,N_5858,N_5270);
nor U7313 (N_7313,N_5630,N_3831);
and U7314 (N_7314,N_5894,N_3254);
xor U7315 (N_7315,N_4596,N_4331);
and U7316 (N_7316,N_3597,N_4964);
nand U7317 (N_7317,N_3132,N_3249);
xor U7318 (N_7318,N_4803,N_4918);
or U7319 (N_7319,N_5146,N_5887);
or U7320 (N_7320,N_5818,N_3787);
nor U7321 (N_7321,N_4387,N_4661);
and U7322 (N_7322,N_5537,N_4153);
nor U7323 (N_7323,N_3424,N_5817);
and U7324 (N_7324,N_5065,N_6211);
nand U7325 (N_7325,N_5839,N_5382);
and U7326 (N_7326,N_5666,N_4903);
nor U7327 (N_7327,N_3673,N_4866);
xnor U7328 (N_7328,N_3435,N_4741);
nand U7329 (N_7329,N_5803,N_4859);
nor U7330 (N_7330,N_3371,N_4002);
xnor U7331 (N_7331,N_4798,N_3265);
nand U7332 (N_7332,N_5989,N_4713);
or U7333 (N_7333,N_3282,N_3695);
and U7334 (N_7334,N_4150,N_3601);
nand U7335 (N_7335,N_4328,N_4070);
nor U7336 (N_7336,N_4720,N_5909);
and U7337 (N_7337,N_5917,N_6002);
and U7338 (N_7338,N_6084,N_4308);
nand U7339 (N_7339,N_5799,N_5659);
nand U7340 (N_7340,N_4425,N_6163);
nor U7341 (N_7341,N_5031,N_4504);
nor U7342 (N_7342,N_4118,N_5364);
and U7343 (N_7343,N_5852,N_4499);
xor U7344 (N_7344,N_3641,N_4965);
nor U7345 (N_7345,N_5772,N_3148);
nand U7346 (N_7346,N_6130,N_5500);
nand U7347 (N_7347,N_5452,N_5923);
nor U7348 (N_7348,N_5246,N_4071);
nand U7349 (N_7349,N_3427,N_4631);
nand U7350 (N_7350,N_5053,N_6179);
nor U7351 (N_7351,N_5605,N_3476);
nor U7352 (N_7352,N_5906,N_4897);
nand U7353 (N_7353,N_5358,N_3799);
nor U7354 (N_7354,N_4877,N_4249);
and U7355 (N_7355,N_3659,N_4785);
and U7356 (N_7356,N_4642,N_4280);
nand U7357 (N_7357,N_4016,N_4705);
or U7358 (N_7358,N_5641,N_3470);
nand U7359 (N_7359,N_5519,N_5834);
nor U7360 (N_7360,N_4309,N_6020);
nand U7361 (N_7361,N_3442,N_3155);
or U7362 (N_7362,N_3674,N_3276);
nand U7363 (N_7363,N_4686,N_5040);
or U7364 (N_7364,N_6160,N_4794);
or U7365 (N_7365,N_4878,N_3350);
and U7366 (N_7366,N_3823,N_3871);
and U7367 (N_7367,N_3777,N_4681);
nor U7368 (N_7368,N_4968,N_6039);
or U7369 (N_7369,N_4654,N_4403);
and U7370 (N_7370,N_4630,N_3693);
or U7371 (N_7371,N_3927,N_5974);
nor U7372 (N_7372,N_5890,N_3930);
nor U7373 (N_7373,N_4635,N_4834);
nor U7374 (N_7374,N_3416,N_4755);
xnor U7375 (N_7375,N_5702,N_4533);
or U7376 (N_7376,N_5762,N_5221);
nand U7377 (N_7377,N_3967,N_4966);
nor U7378 (N_7378,N_5462,N_4102);
or U7379 (N_7379,N_5715,N_5988);
or U7380 (N_7380,N_4082,N_3527);
xnor U7381 (N_7381,N_6060,N_4627);
or U7382 (N_7382,N_3697,N_3430);
or U7383 (N_7383,N_4140,N_4888);
nand U7384 (N_7384,N_4190,N_5019);
or U7385 (N_7385,N_6040,N_4663);
and U7386 (N_7386,N_5359,N_4460);
nand U7387 (N_7387,N_5089,N_3903);
or U7388 (N_7388,N_3506,N_4011);
and U7389 (N_7389,N_5412,N_4660);
xnor U7390 (N_7390,N_4507,N_5959);
nand U7391 (N_7391,N_5939,N_4035);
nor U7392 (N_7392,N_4970,N_5391);
or U7393 (N_7393,N_3185,N_3317);
nand U7394 (N_7394,N_3784,N_5152);
nand U7395 (N_7395,N_5200,N_5985);
nand U7396 (N_7396,N_5251,N_3540);
and U7397 (N_7397,N_5281,N_5586);
or U7398 (N_7398,N_3426,N_5990);
or U7399 (N_7399,N_5725,N_4367);
nor U7400 (N_7400,N_5090,N_4427);
and U7401 (N_7401,N_4664,N_4333);
or U7402 (N_7402,N_3485,N_4969);
or U7403 (N_7403,N_6100,N_3602);
and U7404 (N_7404,N_6182,N_5646);
or U7405 (N_7405,N_4000,N_4912);
and U7406 (N_7406,N_3250,N_4189);
or U7407 (N_7407,N_5695,N_4864);
nand U7408 (N_7408,N_3409,N_3245);
nand U7409 (N_7409,N_5486,N_5136);
nand U7410 (N_7410,N_4775,N_3127);
nand U7411 (N_7411,N_4958,N_3237);
xor U7412 (N_7412,N_4518,N_5722);
or U7413 (N_7413,N_6123,N_4609);
or U7414 (N_7414,N_5509,N_4585);
or U7415 (N_7415,N_4540,N_3711);
xor U7416 (N_7416,N_3770,N_4188);
or U7417 (N_7417,N_6102,N_4770);
nor U7418 (N_7418,N_5348,N_5262);
and U7419 (N_7419,N_5668,N_3681);
or U7420 (N_7420,N_4057,N_5008);
nand U7421 (N_7421,N_5736,N_4465);
or U7422 (N_7422,N_3556,N_5794);
and U7423 (N_7423,N_3369,N_5907);
or U7424 (N_7424,N_3721,N_4152);
or U7425 (N_7425,N_5742,N_3773);
or U7426 (N_7426,N_4819,N_4346);
nand U7427 (N_7427,N_3524,N_5559);
or U7428 (N_7428,N_3368,N_5001);
nor U7429 (N_7429,N_3775,N_5635);
nand U7430 (N_7430,N_3490,N_5916);
and U7431 (N_7431,N_5966,N_4360);
and U7432 (N_7432,N_3730,N_4849);
nor U7433 (N_7433,N_3247,N_3172);
and U7434 (N_7434,N_6026,N_3786);
or U7435 (N_7435,N_3893,N_3137);
and U7436 (N_7436,N_5813,N_3562);
nor U7437 (N_7437,N_4655,N_5429);
and U7438 (N_7438,N_4592,N_4983);
nand U7439 (N_7439,N_3993,N_5553);
and U7440 (N_7440,N_6106,N_3372);
nor U7441 (N_7441,N_5405,N_5215);
or U7442 (N_7442,N_4485,N_4515);
nand U7443 (N_7443,N_3708,N_3500);
and U7444 (N_7444,N_4286,N_6180);
nor U7445 (N_7445,N_3467,N_3364);
nand U7446 (N_7446,N_3344,N_5300);
and U7447 (N_7447,N_4451,N_3510);
or U7448 (N_7448,N_5461,N_3969);
and U7449 (N_7449,N_3395,N_3824);
nand U7450 (N_7450,N_4320,N_3961);
nand U7451 (N_7451,N_3196,N_4858);
xnor U7452 (N_7452,N_5993,N_3498);
nor U7453 (N_7453,N_4979,N_4808);
or U7454 (N_7454,N_4961,N_5319);
nand U7455 (N_7455,N_3816,N_6219);
nand U7456 (N_7456,N_3957,N_6206);
nand U7457 (N_7457,N_4255,N_3574);
and U7458 (N_7458,N_3288,N_4514);
or U7459 (N_7459,N_6158,N_5707);
and U7460 (N_7460,N_4318,N_4203);
or U7461 (N_7461,N_5360,N_3507);
and U7462 (N_7462,N_3342,N_5505);
and U7463 (N_7463,N_4108,N_4593);
and U7464 (N_7464,N_6105,N_3457);
nor U7465 (N_7465,N_5720,N_5748);
nor U7466 (N_7466,N_5526,N_6153);
and U7467 (N_7467,N_5931,N_3195);
and U7468 (N_7468,N_3389,N_3287);
or U7469 (N_7469,N_6059,N_5872);
or U7470 (N_7470,N_5885,N_5498);
and U7471 (N_7471,N_3227,N_3618);
nand U7472 (N_7472,N_3164,N_3864);
and U7473 (N_7473,N_5353,N_4689);
nand U7474 (N_7474,N_3886,N_6191);
nand U7475 (N_7475,N_4675,N_4305);
xor U7476 (N_7476,N_4678,N_5860);
and U7477 (N_7477,N_4506,N_4397);
and U7478 (N_7478,N_3497,N_5143);
nor U7479 (N_7479,N_5976,N_3805);
xor U7480 (N_7480,N_4657,N_5226);
or U7481 (N_7481,N_3339,N_4072);
and U7482 (N_7482,N_5172,N_4124);
and U7483 (N_7483,N_5009,N_5489);
nor U7484 (N_7484,N_4438,N_5312);
or U7485 (N_7485,N_5542,N_5166);
nor U7486 (N_7486,N_6047,N_3475);
and U7487 (N_7487,N_3840,N_4760);
and U7488 (N_7488,N_5419,N_6049);
and U7489 (N_7489,N_4444,N_5032);
nand U7490 (N_7490,N_6045,N_3366);
xor U7491 (N_7491,N_4295,N_4303);
or U7492 (N_7492,N_3606,N_3285);
or U7493 (N_7493,N_5077,N_3232);
or U7494 (N_7494,N_6022,N_5148);
nand U7495 (N_7495,N_5048,N_3534);
xor U7496 (N_7496,N_3537,N_5864);
nor U7497 (N_7497,N_4239,N_5676);
and U7498 (N_7498,N_5387,N_6190);
xor U7499 (N_7499,N_5862,N_3854);
or U7500 (N_7500,N_5740,N_6014);
nor U7501 (N_7501,N_5516,N_4920);
and U7502 (N_7502,N_5006,N_5403);
or U7503 (N_7503,N_4243,N_5582);
and U7504 (N_7504,N_6050,N_3565);
nor U7505 (N_7505,N_4516,N_3382);
xnor U7506 (N_7506,N_3596,N_5871);
and U7507 (N_7507,N_6210,N_4238);
nor U7508 (N_7508,N_4815,N_6006);
xnor U7509 (N_7509,N_5844,N_3599);
xor U7510 (N_7510,N_4461,N_4831);
nor U7511 (N_7511,N_4004,N_3946);
or U7512 (N_7512,N_5232,N_4322);
nand U7513 (N_7513,N_3521,N_3539);
or U7514 (N_7514,N_5561,N_5980);
or U7515 (N_7515,N_5981,N_4457);
and U7516 (N_7516,N_4915,N_5487);
xor U7517 (N_7517,N_4576,N_4371);
nand U7518 (N_7518,N_4886,N_4196);
xnor U7519 (N_7519,N_3896,N_3278);
and U7520 (N_7520,N_5061,N_4567);
xnor U7521 (N_7521,N_4211,N_3508);
nand U7522 (N_7522,N_5933,N_4431);
nand U7523 (N_7523,N_3649,N_5835);
and U7524 (N_7524,N_4138,N_6034);
and U7525 (N_7525,N_3987,N_4028);
nor U7526 (N_7526,N_5693,N_3466);
or U7527 (N_7527,N_3210,N_3997);
xor U7528 (N_7528,N_5289,N_3482);
xor U7529 (N_7529,N_4543,N_3633);
or U7530 (N_7530,N_3458,N_4919);
or U7531 (N_7531,N_4673,N_4205);
or U7532 (N_7532,N_3519,N_5304);
nor U7533 (N_7533,N_5021,N_5763);
or U7534 (N_7534,N_5570,N_6221);
nor U7535 (N_7535,N_4154,N_5796);
nor U7536 (N_7536,N_6103,N_4060);
nor U7537 (N_7537,N_3570,N_3520);
or U7538 (N_7538,N_3712,N_5957);
and U7539 (N_7539,N_3207,N_6198);
and U7540 (N_7540,N_5963,N_5696);
nor U7541 (N_7541,N_5638,N_3910);
and U7542 (N_7542,N_3579,N_5701);
or U7543 (N_7543,N_5023,N_4101);
nand U7544 (N_7544,N_3423,N_5126);
nand U7545 (N_7545,N_3891,N_5464);
and U7546 (N_7546,N_6204,N_4672);
and U7547 (N_7547,N_4401,N_5454);
nor U7548 (N_7548,N_3275,N_4380);
nand U7549 (N_7549,N_5315,N_3549);
nand U7550 (N_7550,N_4321,N_3898);
nand U7551 (N_7551,N_4648,N_6091);
or U7552 (N_7552,N_4564,N_3516);
nor U7553 (N_7553,N_5578,N_3915);
nand U7554 (N_7554,N_3669,N_5903);
and U7555 (N_7555,N_4837,N_4502);
nor U7556 (N_7556,N_3909,N_5352);
nor U7557 (N_7557,N_4365,N_3688);
or U7558 (N_7558,N_5392,N_5798);
nor U7559 (N_7559,N_4251,N_5654);
and U7560 (N_7560,N_3672,N_5078);
nand U7561 (N_7561,N_4045,N_4740);
or U7562 (N_7562,N_4247,N_3761);
or U7563 (N_7563,N_3704,N_6192);
and U7564 (N_7564,N_4141,N_5370);
nand U7565 (N_7565,N_4553,N_4746);
xor U7566 (N_7566,N_5381,N_4603);
and U7567 (N_7567,N_4882,N_5098);
or U7568 (N_7568,N_3813,N_3732);
xor U7569 (N_7569,N_4936,N_5617);
and U7570 (N_7570,N_4176,N_5271);
or U7571 (N_7571,N_5481,N_5513);
nor U7572 (N_7572,N_5483,N_5456);
or U7573 (N_7573,N_5889,N_4737);
nor U7574 (N_7574,N_4519,N_5153);
nand U7575 (N_7575,N_5584,N_3140);
or U7576 (N_7576,N_3772,N_5020);
and U7577 (N_7577,N_4951,N_5124);
nand U7578 (N_7578,N_4723,N_6085);
or U7579 (N_7579,N_3241,N_5624);
or U7580 (N_7580,N_3515,N_5223);
or U7581 (N_7581,N_3496,N_6122);
nand U7582 (N_7582,N_3413,N_4733);
nor U7583 (N_7583,N_3126,N_4679);
nand U7584 (N_7584,N_5220,N_4500);
or U7585 (N_7585,N_4586,N_3683);
or U7586 (N_7586,N_4026,N_3745);
or U7587 (N_7587,N_5196,N_5476);
nor U7588 (N_7588,N_4332,N_5721);
nor U7589 (N_7589,N_5618,N_5343);
and U7590 (N_7590,N_3847,N_4911);
nand U7591 (N_7591,N_5155,N_3918);
or U7592 (N_7592,N_3525,N_5615);
nor U7593 (N_7593,N_4823,N_3863);
xor U7594 (N_7594,N_4710,N_5187);
nor U7595 (N_7595,N_5287,N_3591);
nand U7596 (N_7596,N_4972,N_4347);
nand U7597 (N_7597,N_4537,N_5534);
or U7598 (N_7598,N_3811,N_5010);
and U7599 (N_7599,N_4670,N_4971);
and U7600 (N_7600,N_3959,N_4159);
nand U7601 (N_7601,N_3769,N_5063);
nor U7602 (N_7602,N_6018,N_5488);
or U7603 (N_7603,N_5296,N_3760);
xor U7604 (N_7604,N_5599,N_3713);
nor U7605 (N_7605,N_4690,N_4448);
nand U7606 (N_7606,N_4881,N_4034);
or U7607 (N_7607,N_5135,N_4459);
and U7608 (N_7608,N_4616,N_6185);
nor U7609 (N_7609,N_3504,N_3818);
and U7610 (N_7610,N_3572,N_5002);
and U7611 (N_7611,N_5704,N_4170);
nand U7612 (N_7612,N_4606,N_5544);
and U7613 (N_7613,N_3349,N_5451);
nand U7614 (N_7614,N_6051,N_5644);
or U7615 (N_7615,N_3125,N_5904);
xor U7616 (N_7616,N_3617,N_6146);
or U7617 (N_7617,N_4005,N_4552);
nand U7618 (N_7618,N_4764,N_4790);
nor U7619 (N_7619,N_3536,N_5163);
and U7620 (N_7620,N_4398,N_5830);
and U7621 (N_7621,N_5783,N_4952);
and U7622 (N_7622,N_3838,N_5330);
or U7623 (N_7623,N_5735,N_5932);
and U7624 (N_7624,N_3768,N_3323);
nand U7625 (N_7625,N_3437,N_4285);
nand U7626 (N_7626,N_5785,N_4934);
nand U7627 (N_7627,N_5609,N_5749);
and U7628 (N_7628,N_5003,N_3919);
or U7629 (N_7629,N_4394,N_3353);
nor U7630 (N_7630,N_3600,N_4373);
nor U7631 (N_7631,N_3780,N_3841);
xor U7632 (N_7632,N_3757,N_3874);
or U7633 (N_7633,N_3151,N_5703);
and U7634 (N_7634,N_5286,N_3538);
xnor U7635 (N_7635,N_3905,N_3707);
xor U7636 (N_7636,N_5995,N_4732);
nor U7637 (N_7637,N_4852,N_5790);
nor U7638 (N_7638,N_4316,N_3917);
nand U7639 (N_7639,N_3433,N_3749);
nand U7640 (N_7640,N_6054,N_3613);
or U7641 (N_7641,N_4806,N_3877);
nor U7642 (N_7642,N_4282,N_5892);
xor U7643 (N_7643,N_4544,N_5667);
and U7644 (N_7644,N_5575,N_5567);
nand U7645 (N_7645,N_3152,N_5072);
nand U7646 (N_7646,N_4758,N_3924);
or U7647 (N_7647,N_3947,N_4440);
or U7648 (N_7648,N_5843,N_6241);
nand U7649 (N_7649,N_5846,N_5876);
nand U7650 (N_7650,N_4773,N_3251);
nor U7651 (N_7651,N_3230,N_4962);
and U7652 (N_7652,N_3798,N_4644);
and U7653 (N_7653,N_3302,N_5225);
nand U7654 (N_7654,N_5195,N_5329);
nand U7655 (N_7655,N_5965,N_6222);
xnor U7656 (N_7656,N_3802,N_4266);
nor U7657 (N_7657,N_5113,N_3609);
nor U7658 (N_7658,N_3876,N_3888);
and U7659 (N_7659,N_5212,N_6218);
and U7660 (N_7660,N_3377,N_4851);
nand U7661 (N_7661,N_5341,N_4697);
nor U7662 (N_7662,N_5777,N_4615);
and U7663 (N_7663,N_4402,N_5275);
or U7664 (N_7664,N_6170,N_6134);
nand U7665 (N_7665,N_3984,N_6228);
nand U7666 (N_7666,N_4904,N_5954);
xor U7667 (N_7667,N_3719,N_4668);
nor U7668 (N_7668,N_4062,N_5891);
nor U7669 (N_7669,N_5306,N_4917);
nor U7670 (N_7670,N_4419,N_5177);
and U7671 (N_7671,N_5033,N_4048);
xor U7672 (N_7672,N_3812,N_3290);
or U7673 (N_7673,N_5054,N_4703);
nand U7674 (N_7674,N_3340,N_5311);
nand U7675 (N_7675,N_4067,N_3169);
nand U7676 (N_7676,N_3189,N_4482);
and U7677 (N_7677,N_6043,N_4677);
or U7678 (N_7678,N_4998,N_3890);
or U7679 (N_7679,N_5588,N_5865);
or U7680 (N_7680,N_6030,N_4327);
nor U7681 (N_7681,N_4532,N_5822);
and U7682 (N_7682,N_5944,N_4896);
nand U7683 (N_7683,N_3138,N_5189);
and U7684 (N_7684,N_4008,N_4193);
or U7685 (N_7685,N_4645,N_4524);
and U7686 (N_7686,N_3474,N_6131);
and U7687 (N_7687,N_5103,N_3316);
or U7688 (N_7688,N_4409,N_4393);
nand U7689 (N_7689,N_6243,N_4569);
nand U7690 (N_7690,N_3929,N_6193);
nor U7691 (N_7691,N_4735,N_5838);
or U7692 (N_7692,N_5665,N_4511);
and U7693 (N_7693,N_4160,N_5949);
and U7694 (N_7694,N_3646,N_3699);
nor U7695 (N_7695,N_5207,N_5332);
or U7696 (N_7696,N_3936,N_4871);
nand U7697 (N_7697,N_3978,N_5064);
or U7698 (N_7698,N_3560,N_5430);
and U7699 (N_7699,N_4054,N_4756);
nand U7700 (N_7700,N_3868,N_3130);
or U7701 (N_7701,N_6208,N_6013);
nand U7702 (N_7702,N_4614,N_4292);
nand U7703 (N_7703,N_4669,N_5277);
and U7704 (N_7704,N_3788,N_4195);
and U7705 (N_7705,N_5268,N_3636);
or U7706 (N_7706,N_6042,N_5180);
or U7707 (N_7707,N_4087,N_5497);
nand U7708 (N_7708,N_5812,N_3221);
and U7709 (N_7709,N_5591,N_5724);
nand U7710 (N_7710,N_3418,N_3862);
or U7711 (N_7711,N_5444,N_5645);
xnor U7712 (N_7712,N_5066,N_5297);
nor U7713 (N_7713,N_4636,N_3605);
or U7714 (N_7714,N_5254,N_4315);
nand U7715 (N_7715,N_5051,N_3851);
xnor U7716 (N_7716,N_5130,N_3439);
and U7717 (N_7717,N_5284,N_4802);
nor U7718 (N_7718,N_3558,N_6136);
and U7719 (N_7719,N_4388,N_3724);
nor U7720 (N_7720,N_4229,N_3794);
and U7721 (N_7721,N_6201,N_3956);
nand U7722 (N_7722,N_5535,N_3165);
nor U7723 (N_7723,N_5100,N_3809);
or U7724 (N_7724,N_3404,N_5532);
nor U7725 (N_7725,N_4547,N_5948);
nand U7726 (N_7726,N_3908,N_3356);
and U7727 (N_7727,N_4337,N_3849);
and U7728 (N_7728,N_3454,N_5804);
or U7729 (N_7729,N_4358,N_5210);
nand U7730 (N_7730,N_4113,N_5541);
or U7731 (N_7731,N_5144,N_3291);
and U7732 (N_7732,N_5677,N_5121);
nand U7733 (N_7733,N_5073,N_3970);
nand U7734 (N_7734,N_5808,N_4900);
or U7735 (N_7735,N_3198,N_5746);
xor U7736 (N_7736,N_5915,N_4023);
or U7737 (N_7737,N_4556,N_3289);
or U7738 (N_7738,N_3869,N_4610);
and U7739 (N_7739,N_5986,N_5626);
or U7740 (N_7740,N_5302,N_3541);
or U7741 (N_7741,N_5373,N_4549);
nand U7742 (N_7742,N_3764,N_6202);
nor U7743 (N_7743,N_3281,N_4695);
nand U7744 (N_7744,N_5964,N_3953);
xnor U7745 (N_7745,N_3731,N_4792);
xnor U7746 (N_7746,N_3236,N_5851);
nand U7747 (N_7747,N_5420,N_3434);
and U7748 (N_7748,N_4662,N_3215);
nand U7749 (N_7749,N_4099,N_3821);
and U7750 (N_7750,N_5504,N_4957);
nand U7751 (N_7751,N_3263,N_5896);
nor U7752 (N_7752,N_5085,N_5022);
and U7753 (N_7753,N_3902,N_3819);
and U7754 (N_7754,N_5719,N_3758);
xor U7755 (N_7755,N_4220,N_4525);
and U7756 (N_7756,N_4128,N_4944);
nand U7757 (N_7757,N_4192,N_4724);
or U7758 (N_7758,N_3131,N_5558);
and U7759 (N_7759,N_6092,N_6137);
nand U7760 (N_7760,N_5908,N_5426);
and U7761 (N_7761,N_4488,N_5345);
nand U7762 (N_7762,N_4632,N_5913);
and U7763 (N_7763,N_4130,N_4436);
and U7764 (N_7764,N_4132,N_4931);
nor U7765 (N_7765,N_4612,N_3714);
or U7766 (N_7766,N_5686,N_3826);
or U7767 (N_7767,N_4443,N_4145);
xnor U7768 (N_7768,N_4088,N_4714);
nor U7769 (N_7769,N_3808,N_4978);
nor U7770 (N_7770,N_4963,N_3452);
or U7771 (N_7771,N_5697,N_5026);
nor U7772 (N_7772,N_4469,N_5369);
nor U7773 (N_7773,N_4763,N_5571);
and U7774 (N_7774,N_5517,N_4751);
and U7775 (N_7775,N_3735,N_3879);
nand U7776 (N_7776,N_3133,N_4925);
or U7777 (N_7777,N_4736,N_3964);
xnor U7778 (N_7778,N_3312,N_3220);
and U7779 (N_7779,N_5928,N_4086);
nand U7780 (N_7780,N_6113,N_3180);
or U7781 (N_7781,N_4214,N_4389);
and U7782 (N_7782,N_5111,N_5972);
xnor U7783 (N_7783,N_4268,N_4822);
nand U7784 (N_7784,N_5594,N_3262);
xor U7785 (N_7785,N_3270,N_5543);
nand U7786 (N_7786,N_5362,N_4133);
nand U7787 (N_7787,N_4162,N_4201);
and U7788 (N_7788,N_3177,N_3631);
xor U7789 (N_7789,N_5809,N_6001);
and U7790 (N_7790,N_4986,N_5474);
or U7791 (N_7791,N_3425,N_3723);
and U7792 (N_7792,N_5379,N_5863);
nor U7793 (N_7793,N_3651,N_5199);
nor U7794 (N_7794,N_5608,N_3733);
nor U7795 (N_7795,N_5984,N_3150);
and U7796 (N_7796,N_4216,N_3244);
nand U7797 (N_7797,N_4497,N_4776);
nand U7798 (N_7798,N_4982,N_5466);
or U7799 (N_7799,N_5141,N_4817);
and U7800 (N_7800,N_5478,N_4700);
nor U7801 (N_7801,N_5447,N_4605);
and U7802 (N_7802,N_3566,N_5339);
and U7803 (N_7803,N_4599,N_6066);
nor U7804 (N_7804,N_3392,N_5975);
and U7805 (N_7805,N_3296,N_6033);
nor U7806 (N_7806,N_5034,N_3444);
and U7807 (N_7807,N_3837,N_4600);
nand U7808 (N_7808,N_4727,N_3662);
nand U7809 (N_7809,N_5814,N_4395);
and U7810 (N_7810,N_4774,N_4473);
or U7811 (N_7811,N_4324,N_4810);
and U7812 (N_7812,N_3297,N_5889);
and U7813 (N_7813,N_4048,N_6225);
nor U7814 (N_7814,N_4636,N_5049);
and U7815 (N_7815,N_3804,N_3202);
or U7816 (N_7816,N_3789,N_5536);
and U7817 (N_7817,N_3467,N_5994);
nor U7818 (N_7818,N_3331,N_5349);
or U7819 (N_7819,N_4549,N_5970);
xnor U7820 (N_7820,N_5639,N_4698);
nand U7821 (N_7821,N_4032,N_6057);
nand U7822 (N_7822,N_5726,N_5792);
or U7823 (N_7823,N_5945,N_5384);
and U7824 (N_7824,N_4806,N_5162);
nor U7825 (N_7825,N_4666,N_5447);
nand U7826 (N_7826,N_5551,N_5859);
or U7827 (N_7827,N_3271,N_4199);
nor U7828 (N_7828,N_5473,N_3525);
nand U7829 (N_7829,N_4156,N_4511);
or U7830 (N_7830,N_5031,N_3367);
and U7831 (N_7831,N_5717,N_4646);
nand U7832 (N_7832,N_5979,N_6110);
nor U7833 (N_7833,N_4204,N_3546);
and U7834 (N_7834,N_3168,N_4724);
and U7835 (N_7835,N_3410,N_5279);
nor U7836 (N_7836,N_3382,N_4502);
nor U7837 (N_7837,N_5266,N_5627);
or U7838 (N_7838,N_6105,N_4138);
or U7839 (N_7839,N_5564,N_3934);
nor U7840 (N_7840,N_4491,N_4271);
xnor U7841 (N_7841,N_5678,N_4236);
or U7842 (N_7842,N_5752,N_5669);
nand U7843 (N_7843,N_3793,N_3823);
nor U7844 (N_7844,N_4911,N_5879);
and U7845 (N_7845,N_4150,N_3430);
and U7846 (N_7846,N_4167,N_4659);
and U7847 (N_7847,N_4489,N_3798);
nor U7848 (N_7848,N_4693,N_5823);
nand U7849 (N_7849,N_4808,N_5927);
and U7850 (N_7850,N_3682,N_5821);
and U7851 (N_7851,N_5263,N_4622);
nor U7852 (N_7852,N_4854,N_5112);
xor U7853 (N_7853,N_6032,N_3311);
xnor U7854 (N_7854,N_4159,N_4890);
nor U7855 (N_7855,N_3297,N_5540);
and U7856 (N_7856,N_4830,N_5438);
nand U7857 (N_7857,N_3902,N_3532);
and U7858 (N_7858,N_4006,N_5253);
nand U7859 (N_7859,N_3908,N_6056);
and U7860 (N_7860,N_4373,N_6051);
and U7861 (N_7861,N_3682,N_6100);
nand U7862 (N_7862,N_3991,N_6132);
nand U7863 (N_7863,N_5118,N_4858);
and U7864 (N_7864,N_4372,N_3859);
and U7865 (N_7865,N_3348,N_5281);
and U7866 (N_7866,N_4817,N_4244);
or U7867 (N_7867,N_4433,N_3995);
xor U7868 (N_7868,N_4480,N_6249);
and U7869 (N_7869,N_4092,N_4558);
nor U7870 (N_7870,N_3845,N_3417);
or U7871 (N_7871,N_4589,N_3968);
nor U7872 (N_7872,N_5128,N_4240);
and U7873 (N_7873,N_4364,N_5619);
xnor U7874 (N_7874,N_4293,N_3577);
nor U7875 (N_7875,N_5451,N_6088);
or U7876 (N_7876,N_5568,N_5501);
xor U7877 (N_7877,N_5357,N_3351);
nand U7878 (N_7878,N_3552,N_4195);
nand U7879 (N_7879,N_3915,N_3312);
nor U7880 (N_7880,N_3915,N_3804);
nor U7881 (N_7881,N_5901,N_4667);
nor U7882 (N_7882,N_5048,N_4062);
and U7883 (N_7883,N_5285,N_5544);
nor U7884 (N_7884,N_4225,N_3334);
nand U7885 (N_7885,N_6198,N_5308);
or U7886 (N_7886,N_4905,N_4908);
nand U7887 (N_7887,N_5894,N_4515);
nor U7888 (N_7888,N_5531,N_3152);
or U7889 (N_7889,N_5651,N_6005);
and U7890 (N_7890,N_5280,N_4321);
nor U7891 (N_7891,N_4740,N_5470);
nand U7892 (N_7892,N_3294,N_3631);
or U7893 (N_7893,N_4725,N_3411);
nand U7894 (N_7894,N_4060,N_5583);
nand U7895 (N_7895,N_5516,N_4119);
nor U7896 (N_7896,N_5756,N_6215);
or U7897 (N_7897,N_4642,N_4051);
or U7898 (N_7898,N_5648,N_5170);
nand U7899 (N_7899,N_3862,N_5298);
nand U7900 (N_7900,N_4607,N_5931);
nor U7901 (N_7901,N_3613,N_5888);
nand U7902 (N_7902,N_5928,N_3847);
nand U7903 (N_7903,N_4797,N_4138);
and U7904 (N_7904,N_3607,N_5475);
nand U7905 (N_7905,N_5607,N_4648);
nand U7906 (N_7906,N_6042,N_4604);
nor U7907 (N_7907,N_4198,N_3662);
nand U7908 (N_7908,N_3767,N_4449);
and U7909 (N_7909,N_6038,N_5106);
and U7910 (N_7910,N_4090,N_4999);
xnor U7911 (N_7911,N_5699,N_4165);
nand U7912 (N_7912,N_4467,N_5047);
nand U7913 (N_7913,N_5969,N_3494);
xor U7914 (N_7914,N_5886,N_5411);
nor U7915 (N_7915,N_6114,N_5284);
or U7916 (N_7916,N_4547,N_5445);
nand U7917 (N_7917,N_4520,N_6069);
nor U7918 (N_7918,N_5579,N_3950);
nand U7919 (N_7919,N_3468,N_4215);
or U7920 (N_7920,N_4579,N_5902);
nor U7921 (N_7921,N_4777,N_4728);
or U7922 (N_7922,N_4383,N_5729);
nand U7923 (N_7923,N_5673,N_4609);
or U7924 (N_7924,N_5516,N_3882);
nand U7925 (N_7925,N_4303,N_3733);
or U7926 (N_7926,N_4977,N_4422);
and U7927 (N_7927,N_4493,N_6232);
and U7928 (N_7928,N_3949,N_3714);
nor U7929 (N_7929,N_3867,N_3213);
nor U7930 (N_7930,N_3195,N_5264);
or U7931 (N_7931,N_4026,N_3860);
nand U7932 (N_7932,N_5414,N_5387);
or U7933 (N_7933,N_5158,N_4780);
nor U7934 (N_7934,N_5563,N_4590);
and U7935 (N_7935,N_5254,N_5773);
nor U7936 (N_7936,N_3249,N_3160);
or U7937 (N_7937,N_5046,N_4924);
nand U7938 (N_7938,N_4164,N_5768);
or U7939 (N_7939,N_5654,N_4475);
nand U7940 (N_7940,N_5914,N_6101);
and U7941 (N_7941,N_4359,N_4966);
or U7942 (N_7942,N_3552,N_5357);
nor U7943 (N_7943,N_5458,N_4171);
or U7944 (N_7944,N_4342,N_3763);
or U7945 (N_7945,N_4538,N_3438);
nor U7946 (N_7946,N_5060,N_5480);
and U7947 (N_7947,N_5806,N_3155);
and U7948 (N_7948,N_5910,N_3621);
and U7949 (N_7949,N_5722,N_5427);
nand U7950 (N_7950,N_3830,N_3569);
nand U7951 (N_7951,N_4115,N_3505);
nand U7952 (N_7952,N_4030,N_4536);
nor U7953 (N_7953,N_5758,N_4027);
nor U7954 (N_7954,N_4122,N_5633);
nand U7955 (N_7955,N_3956,N_5157);
nand U7956 (N_7956,N_5189,N_5557);
and U7957 (N_7957,N_6151,N_4025);
and U7958 (N_7958,N_4694,N_5978);
and U7959 (N_7959,N_4014,N_5235);
and U7960 (N_7960,N_3962,N_5404);
and U7961 (N_7961,N_5691,N_4956);
or U7962 (N_7962,N_3260,N_6118);
or U7963 (N_7963,N_5790,N_5942);
xnor U7964 (N_7964,N_5398,N_3254);
nor U7965 (N_7965,N_5126,N_5113);
nand U7966 (N_7966,N_4065,N_4839);
nor U7967 (N_7967,N_3774,N_6015);
nor U7968 (N_7968,N_4139,N_5539);
nand U7969 (N_7969,N_3979,N_4103);
nand U7970 (N_7970,N_3573,N_4739);
nand U7971 (N_7971,N_3794,N_4792);
nor U7972 (N_7972,N_5571,N_6244);
xor U7973 (N_7973,N_5555,N_3908);
and U7974 (N_7974,N_5184,N_3779);
or U7975 (N_7975,N_3471,N_5322);
nor U7976 (N_7976,N_5868,N_4325);
nand U7977 (N_7977,N_4234,N_4721);
or U7978 (N_7978,N_4623,N_5391);
and U7979 (N_7979,N_4580,N_3568);
and U7980 (N_7980,N_5396,N_3447);
and U7981 (N_7981,N_3456,N_4626);
nor U7982 (N_7982,N_4243,N_4458);
nor U7983 (N_7983,N_6197,N_4080);
or U7984 (N_7984,N_3582,N_3702);
nor U7985 (N_7985,N_3499,N_5662);
and U7986 (N_7986,N_4000,N_3949);
and U7987 (N_7987,N_5559,N_3500);
xnor U7988 (N_7988,N_5105,N_6162);
nand U7989 (N_7989,N_4516,N_3780);
nand U7990 (N_7990,N_3704,N_5629);
nand U7991 (N_7991,N_3565,N_3944);
and U7992 (N_7992,N_3732,N_5699);
and U7993 (N_7993,N_4667,N_5236);
and U7994 (N_7994,N_4242,N_4467);
nand U7995 (N_7995,N_5962,N_5544);
and U7996 (N_7996,N_3860,N_5042);
nor U7997 (N_7997,N_3983,N_6127);
nand U7998 (N_7998,N_6102,N_5004);
xor U7999 (N_7999,N_4328,N_4464);
nor U8000 (N_8000,N_4923,N_3902);
and U8001 (N_8001,N_4820,N_5508);
nor U8002 (N_8002,N_5091,N_3507);
nor U8003 (N_8003,N_5483,N_3363);
or U8004 (N_8004,N_4399,N_4375);
and U8005 (N_8005,N_3367,N_5440);
nor U8006 (N_8006,N_5151,N_6129);
and U8007 (N_8007,N_5792,N_5836);
nor U8008 (N_8008,N_6021,N_6089);
and U8009 (N_8009,N_6145,N_3439);
nor U8010 (N_8010,N_4008,N_4068);
nand U8011 (N_8011,N_5576,N_3249);
nand U8012 (N_8012,N_5092,N_6016);
nand U8013 (N_8013,N_6133,N_4979);
nand U8014 (N_8014,N_5245,N_6207);
nand U8015 (N_8015,N_4629,N_5681);
nand U8016 (N_8016,N_3614,N_3320);
xnor U8017 (N_8017,N_3224,N_5433);
or U8018 (N_8018,N_6091,N_3637);
and U8019 (N_8019,N_4202,N_5228);
and U8020 (N_8020,N_5538,N_4691);
nand U8021 (N_8021,N_4231,N_5694);
and U8022 (N_8022,N_5801,N_4340);
and U8023 (N_8023,N_4975,N_3267);
or U8024 (N_8024,N_6151,N_5425);
or U8025 (N_8025,N_3618,N_5154);
and U8026 (N_8026,N_5642,N_6241);
xnor U8027 (N_8027,N_4101,N_4341);
nand U8028 (N_8028,N_5543,N_5877);
and U8029 (N_8029,N_5396,N_5617);
nor U8030 (N_8030,N_3885,N_5523);
or U8031 (N_8031,N_4418,N_4071);
nand U8032 (N_8032,N_4965,N_3651);
and U8033 (N_8033,N_3226,N_3679);
or U8034 (N_8034,N_5373,N_4007);
nor U8035 (N_8035,N_4374,N_3635);
nand U8036 (N_8036,N_4207,N_3930);
and U8037 (N_8037,N_4167,N_3844);
or U8038 (N_8038,N_5931,N_3565);
or U8039 (N_8039,N_4718,N_4841);
nor U8040 (N_8040,N_5872,N_3212);
xnor U8041 (N_8041,N_5370,N_5654);
and U8042 (N_8042,N_3796,N_5413);
nand U8043 (N_8043,N_5622,N_3587);
nand U8044 (N_8044,N_3960,N_5085);
nand U8045 (N_8045,N_3767,N_4514);
and U8046 (N_8046,N_5476,N_5329);
or U8047 (N_8047,N_4537,N_4392);
nand U8048 (N_8048,N_4232,N_5639);
or U8049 (N_8049,N_5246,N_5122);
and U8050 (N_8050,N_3330,N_3302);
or U8051 (N_8051,N_3224,N_4061);
or U8052 (N_8052,N_3683,N_5747);
xor U8053 (N_8053,N_4965,N_5150);
or U8054 (N_8054,N_3197,N_5404);
nor U8055 (N_8055,N_3154,N_4006);
or U8056 (N_8056,N_5109,N_3439);
nor U8057 (N_8057,N_4071,N_3458);
nor U8058 (N_8058,N_6219,N_3332);
xor U8059 (N_8059,N_4498,N_3948);
xor U8060 (N_8060,N_3551,N_3505);
nand U8061 (N_8061,N_3818,N_4708);
or U8062 (N_8062,N_5100,N_5738);
nand U8063 (N_8063,N_4118,N_5543);
nor U8064 (N_8064,N_5488,N_3949);
nor U8065 (N_8065,N_5950,N_5942);
and U8066 (N_8066,N_4437,N_6073);
nor U8067 (N_8067,N_4709,N_4744);
nand U8068 (N_8068,N_4394,N_4196);
and U8069 (N_8069,N_3392,N_3435);
nor U8070 (N_8070,N_3147,N_4961);
nor U8071 (N_8071,N_5941,N_5572);
xnor U8072 (N_8072,N_6079,N_3699);
or U8073 (N_8073,N_5795,N_3553);
nand U8074 (N_8074,N_3305,N_3138);
or U8075 (N_8075,N_5440,N_4232);
nor U8076 (N_8076,N_6049,N_4833);
or U8077 (N_8077,N_4580,N_5511);
and U8078 (N_8078,N_4263,N_4115);
or U8079 (N_8079,N_5132,N_4483);
nand U8080 (N_8080,N_3895,N_4722);
or U8081 (N_8081,N_6121,N_6123);
nand U8082 (N_8082,N_5849,N_6158);
and U8083 (N_8083,N_5565,N_3325);
or U8084 (N_8084,N_6244,N_5007);
nor U8085 (N_8085,N_5927,N_3894);
nand U8086 (N_8086,N_5493,N_4551);
nor U8087 (N_8087,N_3179,N_5483);
and U8088 (N_8088,N_4130,N_4581);
nor U8089 (N_8089,N_4357,N_5489);
and U8090 (N_8090,N_4896,N_5666);
xor U8091 (N_8091,N_3222,N_3542);
or U8092 (N_8092,N_4509,N_4666);
nand U8093 (N_8093,N_4854,N_3991);
nand U8094 (N_8094,N_4448,N_5015);
and U8095 (N_8095,N_5887,N_5513);
xnor U8096 (N_8096,N_3304,N_5870);
or U8097 (N_8097,N_5381,N_3495);
or U8098 (N_8098,N_3258,N_6163);
xor U8099 (N_8099,N_5298,N_5530);
nor U8100 (N_8100,N_5282,N_6150);
and U8101 (N_8101,N_5069,N_5459);
xnor U8102 (N_8102,N_3197,N_4877);
and U8103 (N_8103,N_4726,N_4196);
nand U8104 (N_8104,N_5201,N_4604);
and U8105 (N_8105,N_3261,N_3463);
and U8106 (N_8106,N_4768,N_5790);
nand U8107 (N_8107,N_4335,N_5475);
or U8108 (N_8108,N_4883,N_5818);
and U8109 (N_8109,N_4443,N_6231);
or U8110 (N_8110,N_3284,N_4803);
nor U8111 (N_8111,N_5156,N_5784);
nand U8112 (N_8112,N_5786,N_5980);
nor U8113 (N_8113,N_5504,N_5217);
or U8114 (N_8114,N_4368,N_5875);
xor U8115 (N_8115,N_4954,N_4982);
nor U8116 (N_8116,N_4070,N_3566);
nor U8117 (N_8117,N_4687,N_3807);
nand U8118 (N_8118,N_4662,N_4958);
and U8119 (N_8119,N_4371,N_5378);
and U8120 (N_8120,N_3845,N_4498);
and U8121 (N_8121,N_3151,N_5218);
and U8122 (N_8122,N_4229,N_5514);
nor U8123 (N_8123,N_6171,N_5448);
and U8124 (N_8124,N_4610,N_3430);
nor U8125 (N_8125,N_4812,N_5364);
or U8126 (N_8126,N_3268,N_3809);
or U8127 (N_8127,N_4192,N_4250);
nor U8128 (N_8128,N_4998,N_5875);
and U8129 (N_8129,N_5772,N_4373);
nand U8130 (N_8130,N_6006,N_4420);
or U8131 (N_8131,N_4647,N_3881);
nand U8132 (N_8132,N_5739,N_4580);
and U8133 (N_8133,N_6205,N_4073);
or U8134 (N_8134,N_5636,N_4449);
and U8135 (N_8135,N_6050,N_4502);
nand U8136 (N_8136,N_6222,N_3515);
nor U8137 (N_8137,N_5732,N_4817);
xor U8138 (N_8138,N_5375,N_4103);
nor U8139 (N_8139,N_3679,N_4379);
or U8140 (N_8140,N_5398,N_3158);
or U8141 (N_8141,N_3430,N_3660);
nor U8142 (N_8142,N_4264,N_5515);
and U8143 (N_8143,N_3818,N_5491);
or U8144 (N_8144,N_4762,N_4633);
and U8145 (N_8145,N_3940,N_6185);
or U8146 (N_8146,N_5376,N_3476);
and U8147 (N_8147,N_4881,N_6191);
xor U8148 (N_8148,N_4859,N_5680);
or U8149 (N_8149,N_5682,N_4457);
nor U8150 (N_8150,N_3641,N_5285);
nand U8151 (N_8151,N_5028,N_3885);
or U8152 (N_8152,N_4375,N_3752);
and U8153 (N_8153,N_3464,N_5177);
nor U8154 (N_8154,N_4839,N_4658);
nand U8155 (N_8155,N_4262,N_5840);
nor U8156 (N_8156,N_5292,N_3563);
nand U8157 (N_8157,N_4674,N_5993);
nor U8158 (N_8158,N_5605,N_3455);
nand U8159 (N_8159,N_5292,N_5291);
xnor U8160 (N_8160,N_4594,N_5235);
nand U8161 (N_8161,N_5244,N_6004);
and U8162 (N_8162,N_5997,N_6031);
or U8163 (N_8163,N_6179,N_5445);
xor U8164 (N_8164,N_6123,N_3190);
nor U8165 (N_8165,N_3866,N_4484);
and U8166 (N_8166,N_5107,N_4776);
or U8167 (N_8167,N_5584,N_5324);
or U8168 (N_8168,N_5626,N_5790);
nor U8169 (N_8169,N_5336,N_5098);
and U8170 (N_8170,N_5913,N_6232);
xnor U8171 (N_8171,N_5865,N_4802);
nor U8172 (N_8172,N_5325,N_4364);
and U8173 (N_8173,N_4710,N_3719);
nand U8174 (N_8174,N_5815,N_3357);
nand U8175 (N_8175,N_4514,N_3971);
nor U8176 (N_8176,N_3351,N_3358);
and U8177 (N_8177,N_3157,N_5246);
xor U8178 (N_8178,N_3823,N_5955);
nand U8179 (N_8179,N_4907,N_5074);
nand U8180 (N_8180,N_3856,N_4604);
nor U8181 (N_8181,N_4073,N_5424);
nand U8182 (N_8182,N_5524,N_3197);
and U8183 (N_8183,N_4384,N_5054);
nor U8184 (N_8184,N_3817,N_5633);
xor U8185 (N_8185,N_3841,N_3696);
nor U8186 (N_8186,N_3571,N_3713);
nand U8187 (N_8187,N_3630,N_3697);
or U8188 (N_8188,N_5257,N_6055);
xnor U8189 (N_8189,N_3275,N_4895);
nand U8190 (N_8190,N_4079,N_6115);
xnor U8191 (N_8191,N_4388,N_5938);
nor U8192 (N_8192,N_3850,N_5048);
nand U8193 (N_8193,N_6143,N_3807);
nor U8194 (N_8194,N_4000,N_5427);
nand U8195 (N_8195,N_5182,N_3353);
or U8196 (N_8196,N_4266,N_5998);
or U8197 (N_8197,N_4460,N_5296);
xor U8198 (N_8198,N_4610,N_5220);
and U8199 (N_8199,N_3589,N_4291);
nand U8200 (N_8200,N_4054,N_6120);
nor U8201 (N_8201,N_5563,N_4042);
nor U8202 (N_8202,N_4951,N_4947);
and U8203 (N_8203,N_4524,N_5014);
or U8204 (N_8204,N_3197,N_5936);
nor U8205 (N_8205,N_4535,N_4484);
nor U8206 (N_8206,N_4985,N_4605);
or U8207 (N_8207,N_3418,N_3180);
xnor U8208 (N_8208,N_4890,N_3207);
xnor U8209 (N_8209,N_4279,N_5507);
nand U8210 (N_8210,N_3758,N_5805);
and U8211 (N_8211,N_4783,N_5251);
nand U8212 (N_8212,N_4309,N_4322);
or U8213 (N_8213,N_4439,N_3293);
xor U8214 (N_8214,N_3318,N_6075);
and U8215 (N_8215,N_3231,N_6055);
and U8216 (N_8216,N_4227,N_4555);
nor U8217 (N_8217,N_4554,N_3541);
nand U8218 (N_8218,N_4299,N_4504);
xnor U8219 (N_8219,N_5964,N_4631);
and U8220 (N_8220,N_3856,N_5607);
nor U8221 (N_8221,N_4944,N_3850);
or U8222 (N_8222,N_5282,N_5060);
nand U8223 (N_8223,N_4062,N_6175);
nand U8224 (N_8224,N_5556,N_3738);
nor U8225 (N_8225,N_3652,N_5125);
or U8226 (N_8226,N_5082,N_3200);
or U8227 (N_8227,N_6059,N_5511);
or U8228 (N_8228,N_3454,N_5427);
nand U8229 (N_8229,N_3369,N_6229);
nand U8230 (N_8230,N_6082,N_3870);
nor U8231 (N_8231,N_3875,N_5031);
or U8232 (N_8232,N_3310,N_4262);
nand U8233 (N_8233,N_3436,N_5310);
nand U8234 (N_8234,N_5035,N_3438);
and U8235 (N_8235,N_4261,N_3893);
nor U8236 (N_8236,N_5155,N_3669);
nor U8237 (N_8237,N_5264,N_5165);
nand U8238 (N_8238,N_6009,N_5957);
and U8239 (N_8239,N_4442,N_4538);
nand U8240 (N_8240,N_6135,N_5266);
nand U8241 (N_8241,N_4914,N_5383);
xnor U8242 (N_8242,N_3554,N_4820);
and U8243 (N_8243,N_3196,N_5897);
or U8244 (N_8244,N_5929,N_3494);
xnor U8245 (N_8245,N_4647,N_5924);
or U8246 (N_8246,N_4336,N_5927);
xor U8247 (N_8247,N_4165,N_3982);
or U8248 (N_8248,N_4541,N_3987);
and U8249 (N_8249,N_4424,N_5581);
nand U8250 (N_8250,N_5888,N_6178);
nor U8251 (N_8251,N_4227,N_3728);
nand U8252 (N_8252,N_3599,N_4555);
and U8253 (N_8253,N_3404,N_5726);
and U8254 (N_8254,N_5703,N_3558);
or U8255 (N_8255,N_3420,N_4475);
or U8256 (N_8256,N_3937,N_5302);
or U8257 (N_8257,N_4564,N_3938);
or U8258 (N_8258,N_5582,N_4437);
nand U8259 (N_8259,N_4862,N_3307);
nor U8260 (N_8260,N_5014,N_3642);
nand U8261 (N_8261,N_5895,N_5508);
or U8262 (N_8262,N_4685,N_5482);
xnor U8263 (N_8263,N_5127,N_4679);
nand U8264 (N_8264,N_6138,N_4155);
and U8265 (N_8265,N_5768,N_5540);
xnor U8266 (N_8266,N_3729,N_4316);
nand U8267 (N_8267,N_5238,N_6160);
and U8268 (N_8268,N_3689,N_3935);
and U8269 (N_8269,N_3759,N_3685);
nor U8270 (N_8270,N_5663,N_5591);
and U8271 (N_8271,N_3903,N_4247);
nand U8272 (N_8272,N_4339,N_4409);
nand U8273 (N_8273,N_4832,N_3951);
nor U8274 (N_8274,N_5159,N_3931);
or U8275 (N_8275,N_5556,N_3631);
and U8276 (N_8276,N_4482,N_3304);
nand U8277 (N_8277,N_6055,N_3854);
and U8278 (N_8278,N_5671,N_4258);
nor U8279 (N_8279,N_4191,N_4841);
xor U8280 (N_8280,N_4307,N_4555);
nor U8281 (N_8281,N_6047,N_5118);
xor U8282 (N_8282,N_4369,N_5425);
xor U8283 (N_8283,N_5390,N_4048);
xor U8284 (N_8284,N_5969,N_6042);
nor U8285 (N_8285,N_3341,N_4466);
or U8286 (N_8286,N_4936,N_3809);
and U8287 (N_8287,N_5873,N_4636);
and U8288 (N_8288,N_3609,N_3150);
or U8289 (N_8289,N_5641,N_3181);
and U8290 (N_8290,N_3555,N_5631);
nor U8291 (N_8291,N_4234,N_6151);
nand U8292 (N_8292,N_3305,N_5008);
nor U8293 (N_8293,N_5102,N_5173);
nor U8294 (N_8294,N_5045,N_4094);
and U8295 (N_8295,N_5098,N_5166);
and U8296 (N_8296,N_5592,N_4855);
nand U8297 (N_8297,N_3724,N_5859);
xor U8298 (N_8298,N_3316,N_3450);
nor U8299 (N_8299,N_5065,N_5064);
nor U8300 (N_8300,N_3741,N_6163);
and U8301 (N_8301,N_6083,N_5041);
or U8302 (N_8302,N_3701,N_5046);
nand U8303 (N_8303,N_5597,N_5804);
xor U8304 (N_8304,N_5967,N_4188);
nand U8305 (N_8305,N_4746,N_4667);
or U8306 (N_8306,N_5035,N_4664);
and U8307 (N_8307,N_3705,N_4440);
nor U8308 (N_8308,N_3507,N_3577);
nor U8309 (N_8309,N_4057,N_4444);
xnor U8310 (N_8310,N_3301,N_5751);
nand U8311 (N_8311,N_4749,N_5428);
and U8312 (N_8312,N_4024,N_4606);
and U8313 (N_8313,N_4955,N_3834);
or U8314 (N_8314,N_5703,N_4888);
or U8315 (N_8315,N_4661,N_5212);
nor U8316 (N_8316,N_5352,N_5105);
or U8317 (N_8317,N_3472,N_5892);
or U8318 (N_8318,N_5648,N_3414);
or U8319 (N_8319,N_4885,N_3410);
nand U8320 (N_8320,N_6103,N_4540);
and U8321 (N_8321,N_4048,N_3647);
nor U8322 (N_8322,N_5381,N_3630);
and U8323 (N_8323,N_4844,N_3186);
xnor U8324 (N_8324,N_5122,N_4903);
nand U8325 (N_8325,N_4893,N_6225);
and U8326 (N_8326,N_3760,N_3962);
and U8327 (N_8327,N_5316,N_6145);
nor U8328 (N_8328,N_4076,N_3877);
nor U8329 (N_8329,N_4653,N_3170);
or U8330 (N_8330,N_5622,N_4165);
or U8331 (N_8331,N_6065,N_4025);
nor U8332 (N_8332,N_3179,N_5059);
and U8333 (N_8333,N_3457,N_3129);
or U8334 (N_8334,N_5684,N_4133);
and U8335 (N_8335,N_4436,N_4433);
or U8336 (N_8336,N_3991,N_3473);
nor U8337 (N_8337,N_3349,N_4869);
or U8338 (N_8338,N_6099,N_4661);
or U8339 (N_8339,N_3732,N_4174);
nor U8340 (N_8340,N_3316,N_4678);
or U8341 (N_8341,N_5245,N_5910);
and U8342 (N_8342,N_5185,N_4725);
and U8343 (N_8343,N_3411,N_4253);
or U8344 (N_8344,N_5039,N_4297);
nor U8345 (N_8345,N_4737,N_5838);
nor U8346 (N_8346,N_5069,N_5457);
or U8347 (N_8347,N_3814,N_3564);
nand U8348 (N_8348,N_6239,N_3245);
nor U8349 (N_8349,N_3538,N_5052);
nor U8350 (N_8350,N_3303,N_4195);
or U8351 (N_8351,N_4594,N_4484);
and U8352 (N_8352,N_4666,N_6051);
and U8353 (N_8353,N_6246,N_5948);
or U8354 (N_8354,N_3781,N_3139);
and U8355 (N_8355,N_4524,N_5643);
xnor U8356 (N_8356,N_5398,N_5426);
nand U8357 (N_8357,N_4052,N_6247);
nor U8358 (N_8358,N_5677,N_3200);
and U8359 (N_8359,N_3691,N_5478);
nand U8360 (N_8360,N_4929,N_5832);
or U8361 (N_8361,N_3320,N_5285);
nand U8362 (N_8362,N_5774,N_3902);
nor U8363 (N_8363,N_4483,N_3383);
or U8364 (N_8364,N_3798,N_3377);
and U8365 (N_8365,N_5708,N_3188);
nor U8366 (N_8366,N_4906,N_3607);
nand U8367 (N_8367,N_5482,N_3693);
nor U8368 (N_8368,N_3273,N_4758);
nand U8369 (N_8369,N_5734,N_6126);
and U8370 (N_8370,N_3655,N_3978);
nor U8371 (N_8371,N_5210,N_5932);
or U8372 (N_8372,N_4432,N_5210);
nand U8373 (N_8373,N_6075,N_4636);
nand U8374 (N_8374,N_5509,N_3552);
nor U8375 (N_8375,N_3577,N_4201);
or U8376 (N_8376,N_6128,N_4007);
or U8377 (N_8377,N_5278,N_6092);
nand U8378 (N_8378,N_4991,N_4986);
nand U8379 (N_8379,N_5595,N_5988);
and U8380 (N_8380,N_4735,N_5182);
xor U8381 (N_8381,N_5441,N_3172);
or U8382 (N_8382,N_4004,N_3186);
xor U8383 (N_8383,N_5610,N_6089);
nor U8384 (N_8384,N_3757,N_6115);
xnor U8385 (N_8385,N_5393,N_5492);
nand U8386 (N_8386,N_4946,N_5069);
nor U8387 (N_8387,N_4288,N_5072);
nor U8388 (N_8388,N_5423,N_3483);
and U8389 (N_8389,N_3499,N_6117);
xnor U8390 (N_8390,N_4700,N_4273);
and U8391 (N_8391,N_6163,N_5653);
nor U8392 (N_8392,N_3363,N_5084);
nand U8393 (N_8393,N_3554,N_4713);
nor U8394 (N_8394,N_3126,N_4514);
nor U8395 (N_8395,N_5940,N_5052);
nor U8396 (N_8396,N_3321,N_5900);
nand U8397 (N_8397,N_5244,N_3858);
or U8398 (N_8398,N_6062,N_4441);
or U8399 (N_8399,N_4339,N_5898);
nor U8400 (N_8400,N_4848,N_4717);
and U8401 (N_8401,N_4335,N_3885);
xnor U8402 (N_8402,N_5069,N_5582);
nand U8403 (N_8403,N_3616,N_5279);
xnor U8404 (N_8404,N_3463,N_3867);
or U8405 (N_8405,N_3975,N_6198);
or U8406 (N_8406,N_4254,N_4342);
nand U8407 (N_8407,N_5786,N_3195);
and U8408 (N_8408,N_5603,N_5477);
nor U8409 (N_8409,N_4424,N_5058);
nor U8410 (N_8410,N_3162,N_4942);
nand U8411 (N_8411,N_4107,N_5798);
xnor U8412 (N_8412,N_3781,N_5007);
and U8413 (N_8413,N_5519,N_6083);
xnor U8414 (N_8414,N_4123,N_3713);
or U8415 (N_8415,N_6143,N_3559);
nand U8416 (N_8416,N_5209,N_5299);
and U8417 (N_8417,N_3370,N_4938);
and U8418 (N_8418,N_3822,N_3995);
or U8419 (N_8419,N_6074,N_5725);
nand U8420 (N_8420,N_3194,N_3146);
or U8421 (N_8421,N_5335,N_4102);
nand U8422 (N_8422,N_4750,N_4948);
and U8423 (N_8423,N_5414,N_3573);
or U8424 (N_8424,N_5981,N_4857);
nand U8425 (N_8425,N_4118,N_5086);
nand U8426 (N_8426,N_4188,N_3465);
nor U8427 (N_8427,N_4522,N_4235);
and U8428 (N_8428,N_5398,N_3942);
nand U8429 (N_8429,N_5719,N_4168);
nor U8430 (N_8430,N_4416,N_6242);
and U8431 (N_8431,N_4645,N_5580);
or U8432 (N_8432,N_4168,N_6159);
nand U8433 (N_8433,N_4694,N_5119);
nand U8434 (N_8434,N_3561,N_6055);
nor U8435 (N_8435,N_5707,N_4871);
nand U8436 (N_8436,N_5296,N_4185);
xor U8437 (N_8437,N_4299,N_5782);
nand U8438 (N_8438,N_5426,N_5852);
nor U8439 (N_8439,N_3953,N_3538);
nor U8440 (N_8440,N_4518,N_3713);
nand U8441 (N_8441,N_5671,N_4580);
nand U8442 (N_8442,N_4175,N_5407);
and U8443 (N_8443,N_4200,N_5606);
nand U8444 (N_8444,N_4629,N_3616);
or U8445 (N_8445,N_5230,N_4993);
nand U8446 (N_8446,N_3180,N_5749);
nand U8447 (N_8447,N_4411,N_3954);
nor U8448 (N_8448,N_3523,N_3291);
nand U8449 (N_8449,N_6036,N_5778);
nor U8450 (N_8450,N_4266,N_4904);
xor U8451 (N_8451,N_4933,N_5826);
nand U8452 (N_8452,N_3547,N_3397);
and U8453 (N_8453,N_5746,N_4040);
xnor U8454 (N_8454,N_5897,N_4285);
nand U8455 (N_8455,N_4712,N_4288);
nor U8456 (N_8456,N_3709,N_5314);
and U8457 (N_8457,N_5092,N_4674);
and U8458 (N_8458,N_4656,N_6102);
and U8459 (N_8459,N_5295,N_5783);
and U8460 (N_8460,N_6089,N_5103);
nor U8461 (N_8461,N_5190,N_5147);
and U8462 (N_8462,N_5596,N_3527);
or U8463 (N_8463,N_5287,N_4839);
or U8464 (N_8464,N_3954,N_4891);
and U8465 (N_8465,N_3375,N_6216);
and U8466 (N_8466,N_3153,N_3214);
nand U8467 (N_8467,N_3569,N_5965);
nand U8468 (N_8468,N_4061,N_5323);
nand U8469 (N_8469,N_3534,N_5694);
nand U8470 (N_8470,N_3142,N_6007);
nor U8471 (N_8471,N_4560,N_5235);
nand U8472 (N_8472,N_3274,N_3625);
xor U8473 (N_8473,N_3778,N_4376);
nor U8474 (N_8474,N_5906,N_5377);
nand U8475 (N_8475,N_3163,N_5648);
and U8476 (N_8476,N_3953,N_4874);
and U8477 (N_8477,N_4234,N_5096);
and U8478 (N_8478,N_5183,N_5679);
xor U8479 (N_8479,N_4984,N_5106);
nand U8480 (N_8480,N_6122,N_6030);
nor U8481 (N_8481,N_3222,N_6102);
nand U8482 (N_8482,N_3392,N_3608);
xor U8483 (N_8483,N_3852,N_6113);
and U8484 (N_8484,N_5069,N_5948);
nand U8485 (N_8485,N_6169,N_4201);
nand U8486 (N_8486,N_5341,N_5838);
nor U8487 (N_8487,N_4916,N_4672);
xnor U8488 (N_8488,N_3641,N_6244);
or U8489 (N_8489,N_6215,N_4027);
or U8490 (N_8490,N_3301,N_4710);
or U8491 (N_8491,N_4279,N_4850);
or U8492 (N_8492,N_3279,N_3169);
or U8493 (N_8493,N_5784,N_3718);
nand U8494 (N_8494,N_5932,N_3338);
or U8495 (N_8495,N_3322,N_4044);
nor U8496 (N_8496,N_5076,N_3747);
nand U8497 (N_8497,N_4385,N_5404);
and U8498 (N_8498,N_3528,N_4617);
nor U8499 (N_8499,N_5323,N_3758);
nand U8500 (N_8500,N_5335,N_5636);
nor U8501 (N_8501,N_3147,N_3580);
nand U8502 (N_8502,N_6081,N_5162);
and U8503 (N_8503,N_5553,N_3906);
nand U8504 (N_8504,N_4369,N_5086);
xnor U8505 (N_8505,N_6221,N_5564);
and U8506 (N_8506,N_5056,N_5812);
nor U8507 (N_8507,N_3167,N_6030);
or U8508 (N_8508,N_5325,N_3854);
nor U8509 (N_8509,N_4284,N_3484);
or U8510 (N_8510,N_6080,N_4296);
nor U8511 (N_8511,N_3853,N_4549);
or U8512 (N_8512,N_5584,N_5549);
nor U8513 (N_8513,N_6244,N_5591);
and U8514 (N_8514,N_6201,N_3463);
and U8515 (N_8515,N_3481,N_4443);
or U8516 (N_8516,N_4165,N_4730);
or U8517 (N_8517,N_4723,N_4775);
nor U8518 (N_8518,N_4591,N_5048);
nand U8519 (N_8519,N_4845,N_6084);
and U8520 (N_8520,N_5458,N_5779);
xor U8521 (N_8521,N_4628,N_4678);
nor U8522 (N_8522,N_4082,N_5736);
nand U8523 (N_8523,N_4677,N_4083);
and U8524 (N_8524,N_4904,N_4100);
or U8525 (N_8525,N_6089,N_4372);
or U8526 (N_8526,N_5015,N_3915);
nor U8527 (N_8527,N_6124,N_3557);
or U8528 (N_8528,N_3346,N_3786);
or U8529 (N_8529,N_5212,N_5665);
nor U8530 (N_8530,N_5716,N_4731);
and U8531 (N_8531,N_4672,N_5126);
or U8532 (N_8532,N_5861,N_4735);
and U8533 (N_8533,N_3311,N_5956);
and U8534 (N_8534,N_4627,N_6080);
and U8535 (N_8535,N_4725,N_4116);
nand U8536 (N_8536,N_5675,N_4595);
and U8537 (N_8537,N_4942,N_3475);
and U8538 (N_8538,N_5119,N_3915);
xor U8539 (N_8539,N_3628,N_3307);
xor U8540 (N_8540,N_5104,N_4052);
nand U8541 (N_8541,N_5366,N_4407);
xnor U8542 (N_8542,N_5941,N_3736);
nor U8543 (N_8543,N_5394,N_3561);
nand U8544 (N_8544,N_5905,N_6182);
nor U8545 (N_8545,N_4304,N_5196);
or U8546 (N_8546,N_6141,N_3309);
nand U8547 (N_8547,N_5942,N_6244);
xor U8548 (N_8548,N_4557,N_6196);
nand U8549 (N_8549,N_4463,N_4772);
or U8550 (N_8550,N_5809,N_4850);
nand U8551 (N_8551,N_3402,N_3894);
or U8552 (N_8552,N_3859,N_5193);
xnor U8553 (N_8553,N_3757,N_5732);
or U8554 (N_8554,N_3741,N_4419);
or U8555 (N_8555,N_3898,N_4521);
and U8556 (N_8556,N_3751,N_6113);
xor U8557 (N_8557,N_6083,N_5596);
nor U8558 (N_8558,N_5721,N_5817);
xnor U8559 (N_8559,N_4686,N_5008);
nand U8560 (N_8560,N_3886,N_3650);
or U8561 (N_8561,N_5456,N_4681);
and U8562 (N_8562,N_4913,N_4296);
nand U8563 (N_8563,N_4750,N_3157);
and U8564 (N_8564,N_3622,N_5770);
nor U8565 (N_8565,N_4148,N_3288);
and U8566 (N_8566,N_5856,N_4572);
and U8567 (N_8567,N_4656,N_3168);
xnor U8568 (N_8568,N_5303,N_4866);
nor U8569 (N_8569,N_5188,N_3418);
and U8570 (N_8570,N_3197,N_5779);
or U8571 (N_8571,N_5933,N_4219);
nor U8572 (N_8572,N_5097,N_6080);
and U8573 (N_8573,N_3621,N_3464);
or U8574 (N_8574,N_4012,N_4768);
or U8575 (N_8575,N_3519,N_4435);
xnor U8576 (N_8576,N_5322,N_5398);
or U8577 (N_8577,N_4211,N_4159);
nand U8578 (N_8578,N_3704,N_6226);
or U8579 (N_8579,N_4225,N_5382);
nand U8580 (N_8580,N_5814,N_5579);
and U8581 (N_8581,N_5194,N_4457);
nor U8582 (N_8582,N_5485,N_3781);
or U8583 (N_8583,N_3610,N_5528);
or U8584 (N_8584,N_3591,N_4170);
or U8585 (N_8585,N_3343,N_3565);
nand U8586 (N_8586,N_3407,N_3590);
nand U8587 (N_8587,N_4950,N_5056);
nor U8588 (N_8588,N_3125,N_4829);
or U8589 (N_8589,N_4376,N_5451);
and U8590 (N_8590,N_5560,N_4823);
or U8591 (N_8591,N_6132,N_4434);
and U8592 (N_8592,N_3231,N_5726);
nor U8593 (N_8593,N_3445,N_5291);
or U8594 (N_8594,N_4616,N_4718);
nand U8595 (N_8595,N_5278,N_5270);
or U8596 (N_8596,N_6228,N_4884);
or U8597 (N_8597,N_4025,N_4060);
and U8598 (N_8598,N_3492,N_3141);
nor U8599 (N_8599,N_5908,N_5272);
or U8600 (N_8600,N_4185,N_4258);
xnor U8601 (N_8601,N_5014,N_3360);
xnor U8602 (N_8602,N_5415,N_3225);
and U8603 (N_8603,N_5972,N_6056);
nor U8604 (N_8604,N_4129,N_3770);
and U8605 (N_8605,N_5563,N_3711);
and U8606 (N_8606,N_4338,N_6060);
nor U8607 (N_8607,N_3589,N_5067);
nor U8608 (N_8608,N_6148,N_5361);
and U8609 (N_8609,N_3791,N_3599);
nand U8610 (N_8610,N_5152,N_4798);
nand U8611 (N_8611,N_4301,N_4683);
nor U8612 (N_8612,N_4468,N_5595);
and U8613 (N_8613,N_4095,N_3512);
and U8614 (N_8614,N_5871,N_3797);
nand U8615 (N_8615,N_4862,N_5081);
or U8616 (N_8616,N_3231,N_4586);
nor U8617 (N_8617,N_5710,N_3499);
nand U8618 (N_8618,N_3979,N_5711);
or U8619 (N_8619,N_3543,N_3889);
nand U8620 (N_8620,N_6088,N_6065);
xnor U8621 (N_8621,N_3861,N_5739);
or U8622 (N_8622,N_5082,N_4934);
nor U8623 (N_8623,N_4366,N_4701);
or U8624 (N_8624,N_3285,N_3137);
nand U8625 (N_8625,N_5924,N_3895);
nor U8626 (N_8626,N_3693,N_5081);
or U8627 (N_8627,N_4022,N_3204);
or U8628 (N_8628,N_5466,N_3300);
nor U8629 (N_8629,N_4528,N_4272);
or U8630 (N_8630,N_4989,N_5724);
nand U8631 (N_8631,N_4613,N_5581);
nor U8632 (N_8632,N_5506,N_5656);
or U8633 (N_8633,N_5623,N_5939);
and U8634 (N_8634,N_3881,N_5182);
or U8635 (N_8635,N_3227,N_6169);
xnor U8636 (N_8636,N_5505,N_5370);
nand U8637 (N_8637,N_3872,N_3877);
and U8638 (N_8638,N_5641,N_4097);
and U8639 (N_8639,N_3566,N_3270);
and U8640 (N_8640,N_3802,N_5931);
nand U8641 (N_8641,N_6213,N_5681);
and U8642 (N_8642,N_3350,N_5792);
nor U8643 (N_8643,N_3587,N_4037);
and U8644 (N_8644,N_5445,N_5516);
xnor U8645 (N_8645,N_5438,N_5456);
xnor U8646 (N_8646,N_5273,N_6044);
xor U8647 (N_8647,N_4264,N_5650);
nor U8648 (N_8648,N_5223,N_5130);
nor U8649 (N_8649,N_5524,N_4854);
nand U8650 (N_8650,N_4886,N_3185);
nand U8651 (N_8651,N_4504,N_5428);
and U8652 (N_8652,N_5793,N_5339);
nand U8653 (N_8653,N_3490,N_5552);
or U8654 (N_8654,N_3254,N_4162);
or U8655 (N_8655,N_3363,N_4472);
and U8656 (N_8656,N_4948,N_3373);
nor U8657 (N_8657,N_4500,N_6126);
and U8658 (N_8658,N_5441,N_4494);
and U8659 (N_8659,N_3602,N_5121);
nand U8660 (N_8660,N_3808,N_4538);
nor U8661 (N_8661,N_5219,N_5774);
xor U8662 (N_8662,N_5650,N_5473);
nand U8663 (N_8663,N_4807,N_5305);
nand U8664 (N_8664,N_6097,N_3918);
nor U8665 (N_8665,N_3409,N_3437);
nand U8666 (N_8666,N_3653,N_5461);
nand U8667 (N_8667,N_6122,N_3129);
or U8668 (N_8668,N_3669,N_4257);
nor U8669 (N_8669,N_3405,N_5925);
or U8670 (N_8670,N_5321,N_4385);
and U8671 (N_8671,N_3384,N_3225);
nand U8672 (N_8672,N_4693,N_4304);
nor U8673 (N_8673,N_3846,N_4104);
and U8674 (N_8674,N_5447,N_5633);
xnor U8675 (N_8675,N_4613,N_5112);
and U8676 (N_8676,N_3604,N_3188);
nand U8677 (N_8677,N_3298,N_3727);
nor U8678 (N_8678,N_4706,N_5613);
xor U8679 (N_8679,N_5821,N_5144);
nor U8680 (N_8680,N_4208,N_4315);
nand U8681 (N_8681,N_3208,N_5024);
and U8682 (N_8682,N_5009,N_4964);
nor U8683 (N_8683,N_4088,N_6230);
and U8684 (N_8684,N_3883,N_5430);
or U8685 (N_8685,N_5421,N_5453);
nor U8686 (N_8686,N_3721,N_4213);
and U8687 (N_8687,N_4727,N_5555);
xnor U8688 (N_8688,N_4282,N_4829);
nor U8689 (N_8689,N_4968,N_3323);
nor U8690 (N_8690,N_3941,N_4913);
xnor U8691 (N_8691,N_6112,N_4306);
nand U8692 (N_8692,N_4858,N_3349);
and U8693 (N_8693,N_4702,N_5368);
xnor U8694 (N_8694,N_4905,N_3341);
nand U8695 (N_8695,N_6117,N_6153);
nor U8696 (N_8696,N_5633,N_4404);
nand U8697 (N_8697,N_6082,N_4043);
nand U8698 (N_8698,N_5952,N_3842);
and U8699 (N_8699,N_6045,N_3695);
nand U8700 (N_8700,N_5938,N_3957);
and U8701 (N_8701,N_5790,N_4733);
nor U8702 (N_8702,N_5670,N_5778);
or U8703 (N_8703,N_3546,N_3631);
nand U8704 (N_8704,N_5354,N_3715);
nor U8705 (N_8705,N_6160,N_5078);
nor U8706 (N_8706,N_5410,N_3354);
or U8707 (N_8707,N_6186,N_3538);
nand U8708 (N_8708,N_4849,N_3635);
nor U8709 (N_8709,N_4660,N_4563);
nor U8710 (N_8710,N_6084,N_6206);
xor U8711 (N_8711,N_3605,N_4017);
nand U8712 (N_8712,N_3708,N_3306);
xnor U8713 (N_8713,N_5896,N_3836);
nand U8714 (N_8714,N_3557,N_5849);
xor U8715 (N_8715,N_5137,N_4160);
xnor U8716 (N_8716,N_5357,N_3894);
nor U8717 (N_8717,N_5433,N_4923);
or U8718 (N_8718,N_5460,N_4485);
nand U8719 (N_8719,N_3681,N_3373);
or U8720 (N_8720,N_5332,N_6232);
nand U8721 (N_8721,N_3393,N_4290);
nor U8722 (N_8722,N_4943,N_4733);
nor U8723 (N_8723,N_3361,N_5984);
and U8724 (N_8724,N_4861,N_4498);
nand U8725 (N_8725,N_6135,N_3578);
nor U8726 (N_8726,N_3797,N_3979);
or U8727 (N_8727,N_4002,N_5350);
and U8728 (N_8728,N_4158,N_5176);
nand U8729 (N_8729,N_5685,N_4677);
or U8730 (N_8730,N_4426,N_3509);
or U8731 (N_8731,N_4505,N_3225);
xor U8732 (N_8732,N_4424,N_3936);
nand U8733 (N_8733,N_3368,N_4663);
nand U8734 (N_8734,N_3149,N_5839);
xor U8735 (N_8735,N_5675,N_5373);
nor U8736 (N_8736,N_4904,N_3322);
nand U8737 (N_8737,N_5994,N_4367);
nand U8738 (N_8738,N_4075,N_4414);
nor U8739 (N_8739,N_3581,N_3858);
nand U8740 (N_8740,N_5905,N_3702);
or U8741 (N_8741,N_5926,N_3365);
and U8742 (N_8742,N_5224,N_3626);
or U8743 (N_8743,N_5025,N_5537);
nand U8744 (N_8744,N_5166,N_3610);
and U8745 (N_8745,N_4219,N_4527);
nand U8746 (N_8746,N_4383,N_5485);
nand U8747 (N_8747,N_5897,N_5605);
nand U8748 (N_8748,N_6058,N_5538);
xor U8749 (N_8749,N_5027,N_4013);
nand U8750 (N_8750,N_5799,N_5605);
or U8751 (N_8751,N_5379,N_5193);
nor U8752 (N_8752,N_4437,N_3676);
nor U8753 (N_8753,N_5796,N_5017);
or U8754 (N_8754,N_6238,N_3482);
nor U8755 (N_8755,N_4507,N_4508);
nand U8756 (N_8756,N_3885,N_4912);
xnor U8757 (N_8757,N_4182,N_4046);
or U8758 (N_8758,N_3418,N_6052);
and U8759 (N_8759,N_5225,N_4286);
or U8760 (N_8760,N_5764,N_5677);
xor U8761 (N_8761,N_3535,N_5957);
and U8762 (N_8762,N_4994,N_4431);
or U8763 (N_8763,N_4717,N_4368);
or U8764 (N_8764,N_3579,N_4868);
xnor U8765 (N_8765,N_4072,N_3170);
or U8766 (N_8766,N_3428,N_4039);
nand U8767 (N_8767,N_4147,N_3657);
and U8768 (N_8768,N_3292,N_4544);
xnor U8769 (N_8769,N_3475,N_4620);
or U8770 (N_8770,N_6235,N_4343);
nand U8771 (N_8771,N_6028,N_5298);
nand U8772 (N_8772,N_4518,N_5698);
nand U8773 (N_8773,N_4101,N_6080);
and U8774 (N_8774,N_5246,N_4227);
xnor U8775 (N_8775,N_5791,N_4643);
or U8776 (N_8776,N_4856,N_5782);
or U8777 (N_8777,N_6145,N_3635);
nor U8778 (N_8778,N_5624,N_6224);
and U8779 (N_8779,N_5879,N_3694);
nor U8780 (N_8780,N_5748,N_3962);
nor U8781 (N_8781,N_6216,N_4482);
or U8782 (N_8782,N_4432,N_3623);
nor U8783 (N_8783,N_5922,N_3339);
or U8784 (N_8784,N_4042,N_5095);
or U8785 (N_8785,N_3295,N_4730);
and U8786 (N_8786,N_5804,N_3283);
nand U8787 (N_8787,N_3519,N_5711);
or U8788 (N_8788,N_4664,N_3537);
or U8789 (N_8789,N_5720,N_5159);
and U8790 (N_8790,N_4646,N_4692);
or U8791 (N_8791,N_4943,N_4854);
nand U8792 (N_8792,N_4083,N_3450);
or U8793 (N_8793,N_3651,N_5150);
nor U8794 (N_8794,N_4195,N_4021);
and U8795 (N_8795,N_4998,N_3255);
nand U8796 (N_8796,N_4489,N_3648);
and U8797 (N_8797,N_6010,N_4635);
or U8798 (N_8798,N_3872,N_4031);
and U8799 (N_8799,N_4261,N_5016);
xor U8800 (N_8800,N_5063,N_4151);
xor U8801 (N_8801,N_3611,N_4713);
nor U8802 (N_8802,N_6089,N_5713);
or U8803 (N_8803,N_4781,N_3156);
xnor U8804 (N_8804,N_3696,N_5905);
nand U8805 (N_8805,N_3952,N_5359);
xor U8806 (N_8806,N_6152,N_3554);
xor U8807 (N_8807,N_5821,N_4733);
nor U8808 (N_8808,N_4403,N_6077);
xnor U8809 (N_8809,N_4898,N_5978);
nor U8810 (N_8810,N_5523,N_4311);
and U8811 (N_8811,N_4996,N_5997);
xor U8812 (N_8812,N_5803,N_4531);
and U8813 (N_8813,N_4502,N_4718);
or U8814 (N_8814,N_5806,N_4102);
or U8815 (N_8815,N_5493,N_3701);
nand U8816 (N_8816,N_4054,N_4580);
xor U8817 (N_8817,N_5067,N_3963);
nor U8818 (N_8818,N_4189,N_6033);
nand U8819 (N_8819,N_4179,N_4472);
and U8820 (N_8820,N_5549,N_3254);
or U8821 (N_8821,N_5086,N_3406);
or U8822 (N_8822,N_5908,N_3620);
or U8823 (N_8823,N_3825,N_6014);
and U8824 (N_8824,N_5774,N_5972);
xor U8825 (N_8825,N_4255,N_3293);
nor U8826 (N_8826,N_4426,N_4865);
and U8827 (N_8827,N_5142,N_6000);
nand U8828 (N_8828,N_3731,N_3889);
and U8829 (N_8829,N_4289,N_5082);
nor U8830 (N_8830,N_4003,N_5514);
and U8831 (N_8831,N_3752,N_5735);
xnor U8832 (N_8832,N_3569,N_3336);
nand U8833 (N_8833,N_5329,N_3978);
or U8834 (N_8834,N_3133,N_4360);
and U8835 (N_8835,N_4003,N_6016);
or U8836 (N_8836,N_5889,N_5599);
nand U8837 (N_8837,N_4179,N_5272);
or U8838 (N_8838,N_3861,N_5220);
nand U8839 (N_8839,N_4738,N_5673);
nand U8840 (N_8840,N_3803,N_4180);
and U8841 (N_8841,N_4765,N_3741);
or U8842 (N_8842,N_3253,N_4852);
and U8843 (N_8843,N_4029,N_5111);
or U8844 (N_8844,N_4309,N_3329);
or U8845 (N_8845,N_4655,N_3427);
or U8846 (N_8846,N_3949,N_6211);
or U8847 (N_8847,N_4594,N_4244);
and U8848 (N_8848,N_5021,N_4546);
or U8849 (N_8849,N_5136,N_6169);
nand U8850 (N_8850,N_5610,N_3500);
nand U8851 (N_8851,N_3471,N_5618);
nand U8852 (N_8852,N_4083,N_4840);
or U8853 (N_8853,N_4411,N_5049);
nor U8854 (N_8854,N_4827,N_4678);
nand U8855 (N_8855,N_4841,N_5236);
nand U8856 (N_8856,N_3324,N_4493);
nand U8857 (N_8857,N_5068,N_4667);
or U8858 (N_8858,N_4638,N_4490);
or U8859 (N_8859,N_3465,N_4845);
or U8860 (N_8860,N_4228,N_3846);
nand U8861 (N_8861,N_4856,N_4316);
and U8862 (N_8862,N_5183,N_4205);
or U8863 (N_8863,N_6020,N_5031);
xor U8864 (N_8864,N_3796,N_4815);
nor U8865 (N_8865,N_5682,N_5844);
nand U8866 (N_8866,N_5045,N_3935);
xnor U8867 (N_8867,N_4971,N_4126);
nor U8868 (N_8868,N_4170,N_6185);
nor U8869 (N_8869,N_5778,N_6168);
and U8870 (N_8870,N_3798,N_4286);
nor U8871 (N_8871,N_5675,N_6240);
nor U8872 (N_8872,N_3733,N_4224);
and U8873 (N_8873,N_3263,N_3790);
nor U8874 (N_8874,N_3743,N_4988);
nand U8875 (N_8875,N_4067,N_4734);
or U8876 (N_8876,N_4051,N_6208);
nand U8877 (N_8877,N_3487,N_5533);
and U8878 (N_8878,N_6038,N_3565);
nand U8879 (N_8879,N_4697,N_4764);
or U8880 (N_8880,N_5170,N_5821);
and U8881 (N_8881,N_4077,N_3640);
nand U8882 (N_8882,N_5831,N_3408);
nand U8883 (N_8883,N_4055,N_5926);
or U8884 (N_8884,N_5511,N_6177);
nand U8885 (N_8885,N_5768,N_3771);
nor U8886 (N_8886,N_4151,N_3829);
xor U8887 (N_8887,N_5551,N_3326);
nor U8888 (N_8888,N_5261,N_5826);
and U8889 (N_8889,N_4474,N_4581);
nor U8890 (N_8890,N_3319,N_4159);
nor U8891 (N_8891,N_3629,N_3248);
nor U8892 (N_8892,N_4695,N_4495);
nor U8893 (N_8893,N_4684,N_5311);
or U8894 (N_8894,N_3246,N_5482);
or U8895 (N_8895,N_3875,N_5842);
nor U8896 (N_8896,N_5754,N_5818);
nand U8897 (N_8897,N_5885,N_4927);
nand U8898 (N_8898,N_6189,N_6112);
xnor U8899 (N_8899,N_3288,N_4552);
and U8900 (N_8900,N_5622,N_4983);
and U8901 (N_8901,N_3801,N_5447);
or U8902 (N_8902,N_3416,N_5321);
nand U8903 (N_8903,N_5094,N_3858);
or U8904 (N_8904,N_5395,N_5101);
and U8905 (N_8905,N_5191,N_3369);
nand U8906 (N_8906,N_5569,N_5280);
nand U8907 (N_8907,N_5681,N_5904);
nand U8908 (N_8908,N_3166,N_4093);
and U8909 (N_8909,N_6235,N_5272);
xnor U8910 (N_8910,N_5094,N_3153);
nor U8911 (N_8911,N_5791,N_4986);
or U8912 (N_8912,N_4851,N_4536);
nor U8913 (N_8913,N_5734,N_5184);
and U8914 (N_8914,N_6086,N_5176);
nor U8915 (N_8915,N_5744,N_4767);
xor U8916 (N_8916,N_3544,N_3479);
nor U8917 (N_8917,N_4839,N_3538);
and U8918 (N_8918,N_3796,N_3248);
nand U8919 (N_8919,N_5449,N_5233);
or U8920 (N_8920,N_5542,N_5160);
and U8921 (N_8921,N_6032,N_3608);
xor U8922 (N_8922,N_5280,N_4551);
nor U8923 (N_8923,N_3581,N_4933);
nand U8924 (N_8924,N_5069,N_3532);
nor U8925 (N_8925,N_3126,N_6249);
nor U8926 (N_8926,N_5135,N_3812);
nand U8927 (N_8927,N_3268,N_4194);
nor U8928 (N_8928,N_4830,N_4453);
and U8929 (N_8929,N_4676,N_6177);
and U8930 (N_8930,N_4145,N_3827);
nor U8931 (N_8931,N_5749,N_3452);
nor U8932 (N_8932,N_4970,N_6037);
nor U8933 (N_8933,N_6121,N_4409);
nor U8934 (N_8934,N_5319,N_5979);
or U8935 (N_8935,N_4872,N_5796);
nand U8936 (N_8936,N_3152,N_3519);
nor U8937 (N_8937,N_4908,N_5349);
nand U8938 (N_8938,N_3615,N_4670);
and U8939 (N_8939,N_3232,N_6014);
or U8940 (N_8940,N_5057,N_4089);
or U8941 (N_8941,N_6094,N_4313);
or U8942 (N_8942,N_4611,N_3607);
or U8943 (N_8943,N_4871,N_5974);
nand U8944 (N_8944,N_3442,N_5072);
or U8945 (N_8945,N_6243,N_3644);
nor U8946 (N_8946,N_3643,N_5932);
nand U8947 (N_8947,N_5991,N_5747);
or U8948 (N_8948,N_4929,N_3629);
or U8949 (N_8949,N_5282,N_3323);
nor U8950 (N_8950,N_3275,N_3568);
and U8951 (N_8951,N_4651,N_4839);
and U8952 (N_8952,N_5728,N_5987);
nor U8953 (N_8953,N_3235,N_5067);
and U8954 (N_8954,N_5575,N_5077);
xor U8955 (N_8955,N_5640,N_3159);
nor U8956 (N_8956,N_3518,N_6148);
and U8957 (N_8957,N_5552,N_5731);
or U8958 (N_8958,N_3518,N_4766);
or U8959 (N_8959,N_5394,N_3892);
nor U8960 (N_8960,N_4257,N_4597);
nor U8961 (N_8961,N_6078,N_4729);
nand U8962 (N_8962,N_4059,N_4330);
nand U8963 (N_8963,N_6190,N_4986);
or U8964 (N_8964,N_3692,N_3902);
nor U8965 (N_8965,N_5971,N_6133);
nand U8966 (N_8966,N_6033,N_5541);
or U8967 (N_8967,N_3621,N_6216);
or U8968 (N_8968,N_4510,N_5479);
nand U8969 (N_8969,N_5285,N_3213);
and U8970 (N_8970,N_3649,N_6174);
and U8971 (N_8971,N_5768,N_5371);
nor U8972 (N_8972,N_4227,N_4367);
nand U8973 (N_8973,N_3535,N_4262);
nor U8974 (N_8974,N_3695,N_4301);
nand U8975 (N_8975,N_5605,N_3338);
and U8976 (N_8976,N_5963,N_5434);
or U8977 (N_8977,N_3740,N_4271);
or U8978 (N_8978,N_6094,N_3556);
nand U8979 (N_8979,N_5664,N_4046);
nand U8980 (N_8980,N_4790,N_4082);
and U8981 (N_8981,N_5638,N_4116);
or U8982 (N_8982,N_6171,N_3932);
and U8983 (N_8983,N_5965,N_5920);
and U8984 (N_8984,N_5050,N_5175);
or U8985 (N_8985,N_6184,N_4698);
and U8986 (N_8986,N_3893,N_5591);
and U8987 (N_8987,N_5952,N_4005);
nor U8988 (N_8988,N_5198,N_4954);
and U8989 (N_8989,N_5384,N_5314);
nand U8990 (N_8990,N_5595,N_6111);
and U8991 (N_8991,N_4359,N_5143);
and U8992 (N_8992,N_3861,N_4938);
nor U8993 (N_8993,N_5396,N_6041);
nor U8994 (N_8994,N_3328,N_3921);
nand U8995 (N_8995,N_3633,N_4145);
nand U8996 (N_8996,N_3572,N_3995);
nor U8997 (N_8997,N_4982,N_5159);
nand U8998 (N_8998,N_4632,N_5627);
xor U8999 (N_8999,N_5221,N_5824);
and U9000 (N_9000,N_6050,N_5764);
or U9001 (N_9001,N_5663,N_4893);
or U9002 (N_9002,N_5467,N_4490);
nand U9003 (N_9003,N_3570,N_6122);
nand U9004 (N_9004,N_3863,N_5693);
or U9005 (N_9005,N_3573,N_3493);
and U9006 (N_9006,N_5621,N_4346);
xnor U9007 (N_9007,N_4863,N_5631);
nor U9008 (N_9008,N_3384,N_4166);
nand U9009 (N_9009,N_6014,N_3333);
nor U9010 (N_9010,N_4784,N_4551);
and U9011 (N_9011,N_4977,N_3511);
or U9012 (N_9012,N_4153,N_3667);
or U9013 (N_9013,N_4605,N_5819);
nand U9014 (N_9014,N_6067,N_5630);
or U9015 (N_9015,N_5202,N_4669);
or U9016 (N_9016,N_4772,N_4512);
nand U9017 (N_9017,N_3887,N_3724);
and U9018 (N_9018,N_5185,N_5914);
and U9019 (N_9019,N_4794,N_3130);
or U9020 (N_9020,N_3838,N_4723);
xor U9021 (N_9021,N_6026,N_6216);
or U9022 (N_9022,N_3988,N_5342);
nand U9023 (N_9023,N_5183,N_4470);
nor U9024 (N_9024,N_3529,N_3924);
nand U9025 (N_9025,N_4658,N_6074);
nand U9026 (N_9026,N_4555,N_4605);
and U9027 (N_9027,N_5805,N_5494);
nor U9028 (N_9028,N_4376,N_5904);
nor U9029 (N_9029,N_5671,N_4445);
nor U9030 (N_9030,N_5045,N_5718);
and U9031 (N_9031,N_5439,N_6081);
or U9032 (N_9032,N_5638,N_5035);
nor U9033 (N_9033,N_4564,N_3979);
or U9034 (N_9034,N_4757,N_4957);
or U9035 (N_9035,N_3186,N_3773);
nor U9036 (N_9036,N_4103,N_4869);
or U9037 (N_9037,N_3262,N_5998);
nand U9038 (N_9038,N_4865,N_5983);
or U9039 (N_9039,N_5758,N_5105);
and U9040 (N_9040,N_3451,N_3423);
or U9041 (N_9041,N_5240,N_3200);
nor U9042 (N_9042,N_3614,N_6200);
nor U9043 (N_9043,N_4778,N_5974);
nor U9044 (N_9044,N_5435,N_6022);
xnor U9045 (N_9045,N_3435,N_3504);
or U9046 (N_9046,N_3955,N_3370);
nor U9047 (N_9047,N_3350,N_5210);
nor U9048 (N_9048,N_5541,N_4469);
xor U9049 (N_9049,N_6189,N_4467);
or U9050 (N_9050,N_5952,N_5018);
or U9051 (N_9051,N_3984,N_6197);
nand U9052 (N_9052,N_5931,N_3405);
nand U9053 (N_9053,N_4888,N_5853);
nor U9054 (N_9054,N_4676,N_5144);
or U9055 (N_9055,N_4176,N_5859);
nand U9056 (N_9056,N_6039,N_3179);
or U9057 (N_9057,N_3284,N_4865);
nor U9058 (N_9058,N_3315,N_5661);
and U9059 (N_9059,N_4689,N_4345);
nor U9060 (N_9060,N_4958,N_5021);
or U9061 (N_9061,N_4870,N_3605);
nand U9062 (N_9062,N_3347,N_3920);
or U9063 (N_9063,N_4077,N_4348);
nand U9064 (N_9064,N_5552,N_6107);
nand U9065 (N_9065,N_5032,N_3333);
and U9066 (N_9066,N_6044,N_4688);
or U9067 (N_9067,N_3137,N_4982);
nand U9068 (N_9068,N_4175,N_3455);
or U9069 (N_9069,N_5462,N_5117);
nor U9070 (N_9070,N_5636,N_4404);
xnor U9071 (N_9071,N_3654,N_3756);
nand U9072 (N_9072,N_5809,N_3990);
nor U9073 (N_9073,N_3435,N_5602);
nand U9074 (N_9074,N_4727,N_4706);
nor U9075 (N_9075,N_5802,N_5672);
and U9076 (N_9076,N_5956,N_4865);
nor U9077 (N_9077,N_3734,N_3386);
nand U9078 (N_9078,N_3807,N_5855);
xor U9079 (N_9079,N_5331,N_3199);
and U9080 (N_9080,N_4789,N_3648);
and U9081 (N_9081,N_5938,N_6058);
and U9082 (N_9082,N_4782,N_4445);
and U9083 (N_9083,N_5050,N_4823);
and U9084 (N_9084,N_4783,N_4991);
and U9085 (N_9085,N_4977,N_3209);
nand U9086 (N_9086,N_5227,N_3527);
or U9087 (N_9087,N_5419,N_5635);
and U9088 (N_9088,N_5958,N_3858);
nand U9089 (N_9089,N_4398,N_3842);
nor U9090 (N_9090,N_3698,N_6091);
nor U9091 (N_9091,N_4620,N_4854);
and U9092 (N_9092,N_6003,N_5099);
nor U9093 (N_9093,N_5696,N_3130);
or U9094 (N_9094,N_4459,N_4401);
and U9095 (N_9095,N_5567,N_3205);
xor U9096 (N_9096,N_5471,N_3904);
nand U9097 (N_9097,N_4260,N_4136);
and U9098 (N_9098,N_5386,N_5330);
and U9099 (N_9099,N_5893,N_3354);
nor U9100 (N_9100,N_5628,N_5438);
nor U9101 (N_9101,N_4924,N_4482);
nor U9102 (N_9102,N_5153,N_4101);
and U9103 (N_9103,N_4188,N_6219);
and U9104 (N_9104,N_4550,N_3910);
or U9105 (N_9105,N_4105,N_3198);
or U9106 (N_9106,N_4770,N_3673);
and U9107 (N_9107,N_4742,N_5692);
and U9108 (N_9108,N_3660,N_5511);
or U9109 (N_9109,N_5585,N_5430);
and U9110 (N_9110,N_5499,N_5460);
nor U9111 (N_9111,N_4747,N_4946);
and U9112 (N_9112,N_5510,N_6245);
or U9113 (N_9113,N_4578,N_5641);
and U9114 (N_9114,N_4241,N_3867);
xor U9115 (N_9115,N_4257,N_4858);
nand U9116 (N_9116,N_6001,N_4361);
nor U9117 (N_9117,N_5081,N_3137);
and U9118 (N_9118,N_3937,N_3660);
nand U9119 (N_9119,N_3741,N_5246);
nand U9120 (N_9120,N_4373,N_4122);
nor U9121 (N_9121,N_3653,N_4514);
and U9122 (N_9122,N_4999,N_3774);
nor U9123 (N_9123,N_4424,N_5715);
nor U9124 (N_9124,N_4440,N_3157);
nand U9125 (N_9125,N_3541,N_3949);
nor U9126 (N_9126,N_5029,N_5022);
and U9127 (N_9127,N_6205,N_5579);
or U9128 (N_9128,N_4345,N_3899);
nor U9129 (N_9129,N_4333,N_3844);
and U9130 (N_9130,N_5811,N_3555);
or U9131 (N_9131,N_4244,N_5487);
nand U9132 (N_9132,N_4376,N_6088);
nor U9133 (N_9133,N_5981,N_5995);
nand U9134 (N_9134,N_5135,N_5575);
and U9135 (N_9135,N_4897,N_5878);
and U9136 (N_9136,N_3274,N_5455);
xnor U9137 (N_9137,N_3601,N_4800);
or U9138 (N_9138,N_4804,N_3587);
nand U9139 (N_9139,N_4447,N_4572);
and U9140 (N_9140,N_4516,N_3548);
nor U9141 (N_9141,N_5085,N_5317);
nor U9142 (N_9142,N_4023,N_4841);
nand U9143 (N_9143,N_3670,N_5189);
nor U9144 (N_9144,N_3807,N_3727);
nor U9145 (N_9145,N_5606,N_5066);
or U9146 (N_9146,N_5133,N_4924);
nor U9147 (N_9147,N_6207,N_6128);
xor U9148 (N_9148,N_5189,N_6000);
or U9149 (N_9149,N_3907,N_4849);
nand U9150 (N_9150,N_5959,N_3885);
xnor U9151 (N_9151,N_4067,N_5077);
and U9152 (N_9152,N_3921,N_6150);
nor U9153 (N_9153,N_4838,N_6240);
and U9154 (N_9154,N_5329,N_5585);
xnor U9155 (N_9155,N_5906,N_5927);
nor U9156 (N_9156,N_4831,N_6035);
or U9157 (N_9157,N_5261,N_5323);
and U9158 (N_9158,N_3195,N_6191);
or U9159 (N_9159,N_3354,N_3931);
nand U9160 (N_9160,N_4400,N_4853);
and U9161 (N_9161,N_4598,N_6037);
nand U9162 (N_9162,N_3869,N_4014);
nor U9163 (N_9163,N_4724,N_3943);
nor U9164 (N_9164,N_4851,N_5549);
and U9165 (N_9165,N_6010,N_3376);
or U9166 (N_9166,N_5522,N_4254);
or U9167 (N_9167,N_5754,N_4437);
xnor U9168 (N_9168,N_3708,N_3990);
nor U9169 (N_9169,N_5080,N_4262);
and U9170 (N_9170,N_3971,N_3981);
or U9171 (N_9171,N_3204,N_5393);
nor U9172 (N_9172,N_5439,N_3586);
nor U9173 (N_9173,N_3863,N_5283);
and U9174 (N_9174,N_4573,N_5814);
or U9175 (N_9175,N_3189,N_4383);
or U9176 (N_9176,N_4998,N_4416);
nor U9177 (N_9177,N_3825,N_4335);
nor U9178 (N_9178,N_5014,N_5414);
and U9179 (N_9179,N_3284,N_5353);
and U9180 (N_9180,N_5411,N_5006);
and U9181 (N_9181,N_5467,N_3948);
or U9182 (N_9182,N_4868,N_5403);
or U9183 (N_9183,N_4364,N_5826);
nor U9184 (N_9184,N_4410,N_4324);
and U9185 (N_9185,N_6194,N_3372);
nand U9186 (N_9186,N_5599,N_5909);
nor U9187 (N_9187,N_3828,N_5131);
and U9188 (N_9188,N_5495,N_3159);
or U9189 (N_9189,N_4594,N_5125);
or U9190 (N_9190,N_4790,N_3900);
or U9191 (N_9191,N_4974,N_5436);
nand U9192 (N_9192,N_4881,N_4096);
nor U9193 (N_9193,N_5608,N_6208);
nand U9194 (N_9194,N_3898,N_4600);
nand U9195 (N_9195,N_4666,N_4907);
xor U9196 (N_9196,N_4229,N_5747);
or U9197 (N_9197,N_4385,N_3395);
nor U9198 (N_9198,N_5076,N_4288);
nor U9199 (N_9199,N_5728,N_5606);
nand U9200 (N_9200,N_3946,N_4626);
or U9201 (N_9201,N_6190,N_3669);
xor U9202 (N_9202,N_3560,N_5814);
and U9203 (N_9203,N_5529,N_4351);
nand U9204 (N_9204,N_4557,N_5666);
and U9205 (N_9205,N_3453,N_3902);
nand U9206 (N_9206,N_4138,N_4588);
xnor U9207 (N_9207,N_3549,N_6216);
xor U9208 (N_9208,N_5289,N_5263);
or U9209 (N_9209,N_3334,N_5646);
nand U9210 (N_9210,N_4344,N_5792);
and U9211 (N_9211,N_4660,N_4359);
nand U9212 (N_9212,N_5106,N_3126);
nor U9213 (N_9213,N_6130,N_4362);
or U9214 (N_9214,N_6174,N_4423);
xnor U9215 (N_9215,N_4587,N_3599);
nor U9216 (N_9216,N_6160,N_3713);
or U9217 (N_9217,N_4745,N_5609);
and U9218 (N_9218,N_5416,N_5891);
and U9219 (N_9219,N_6209,N_5617);
nand U9220 (N_9220,N_3356,N_3899);
or U9221 (N_9221,N_3349,N_3855);
nor U9222 (N_9222,N_3645,N_5801);
nand U9223 (N_9223,N_5811,N_3285);
and U9224 (N_9224,N_4637,N_5014);
or U9225 (N_9225,N_4724,N_4831);
or U9226 (N_9226,N_5356,N_3859);
and U9227 (N_9227,N_6008,N_3174);
and U9228 (N_9228,N_3776,N_4450);
nand U9229 (N_9229,N_6050,N_4767);
or U9230 (N_9230,N_5511,N_3130);
and U9231 (N_9231,N_4007,N_4929);
nand U9232 (N_9232,N_5605,N_3961);
nand U9233 (N_9233,N_3156,N_4320);
xor U9234 (N_9234,N_3228,N_4098);
or U9235 (N_9235,N_5608,N_3596);
nand U9236 (N_9236,N_3993,N_3386);
and U9237 (N_9237,N_5586,N_5804);
nor U9238 (N_9238,N_6166,N_5419);
or U9239 (N_9239,N_3146,N_5544);
or U9240 (N_9240,N_5614,N_5766);
or U9241 (N_9241,N_5659,N_3148);
and U9242 (N_9242,N_5706,N_5347);
nor U9243 (N_9243,N_3337,N_4926);
nor U9244 (N_9244,N_6245,N_4917);
nor U9245 (N_9245,N_3687,N_4738);
nor U9246 (N_9246,N_4692,N_5117);
nor U9247 (N_9247,N_4925,N_3148);
xor U9248 (N_9248,N_4016,N_5373);
nand U9249 (N_9249,N_6023,N_6107);
nand U9250 (N_9250,N_5488,N_5616);
nand U9251 (N_9251,N_5225,N_6184);
nor U9252 (N_9252,N_5035,N_4088);
nand U9253 (N_9253,N_5369,N_3588);
and U9254 (N_9254,N_3942,N_4302);
nand U9255 (N_9255,N_3663,N_4882);
nor U9256 (N_9256,N_3561,N_6039);
nor U9257 (N_9257,N_6193,N_3778);
nand U9258 (N_9258,N_4490,N_6177);
and U9259 (N_9259,N_5414,N_4006);
and U9260 (N_9260,N_5391,N_5654);
and U9261 (N_9261,N_5242,N_5009);
nor U9262 (N_9262,N_5699,N_4887);
xnor U9263 (N_9263,N_6069,N_5893);
xor U9264 (N_9264,N_5846,N_5655);
and U9265 (N_9265,N_6000,N_5621);
nor U9266 (N_9266,N_3236,N_5847);
and U9267 (N_9267,N_6102,N_6174);
or U9268 (N_9268,N_4267,N_3589);
and U9269 (N_9269,N_3883,N_5112);
nor U9270 (N_9270,N_6210,N_4604);
and U9271 (N_9271,N_4824,N_3405);
and U9272 (N_9272,N_4437,N_3696);
and U9273 (N_9273,N_3896,N_4059);
nand U9274 (N_9274,N_6193,N_5691);
and U9275 (N_9275,N_6103,N_3981);
nor U9276 (N_9276,N_3709,N_4198);
nand U9277 (N_9277,N_5454,N_5053);
and U9278 (N_9278,N_5267,N_6220);
and U9279 (N_9279,N_6156,N_5077);
and U9280 (N_9280,N_5006,N_4519);
or U9281 (N_9281,N_5189,N_4074);
nor U9282 (N_9282,N_5860,N_3444);
and U9283 (N_9283,N_3797,N_3281);
nor U9284 (N_9284,N_4126,N_5868);
xor U9285 (N_9285,N_5312,N_6225);
nand U9286 (N_9286,N_5207,N_3414);
nand U9287 (N_9287,N_5693,N_4813);
and U9288 (N_9288,N_5663,N_4715);
nand U9289 (N_9289,N_3656,N_3497);
and U9290 (N_9290,N_4063,N_3530);
or U9291 (N_9291,N_3954,N_4170);
nor U9292 (N_9292,N_3284,N_3551);
nor U9293 (N_9293,N_4745,N_4655);
xor U9294 (N_9294,N_5228,N_3129);
nor U9295 (N_9295,N_4562,N_3511);
or U9296 (N_9296,N_5492,N_5687);
nand U9297 (N_9297,N_4351,N_5076);
nand U9298 (N_9298,N_4952,N_3932);
and U9299 (N_9299,N_5742,N_4778);
nand U9300 (N_9300,N_4927,N_5244);
nand U9301 (N_9301,N_3360,N_3183);
or U9302 (N_9302,N_6187,N_6047);
nand U9303 (N_9303,N_3734,N_4214);
and U9304 (N_9304,N_4926,N_3493);
xnor U9305 (N_9305,N_5592,N_6151);
nand U9306 (N_9306,N_6048,N_4140);
or U9307 (N_9307,N_3681,N_5829);
and U9308 (N_9308,N_4133,N_5088);
xor U9309 (N_9309,N_3431,N_5517);
or U9310 (N_9310,N_5503,N_5029);
and U9311 (N_9311,N_4977,N_4954);
or U9312 (N_9312,N_5117,N_5548);
or U9313 (N_9313,N_4738,N_3919);
or U9314 (N_9314,N_5313,N_6098);
nor U9315 (N_9315,N_4842,N_4386);
or U9316 (N_9316,N_3561,N_6179);
and U9317 (N_9317,N_6104,N_5867);
and U9318 (N_9318,N_4802,N_5879);
nor U9319 (N_9319,N_5126,N_3992);
xor U9320 (N_9320,N_4558,N_4493);
nor U9321 (N_9321,N_3956,N_5262);
nor U9322 (N_9322,N_3188,N_5511);
nor U9323 (N_9323,N_5081,N_4021);
or U9324 (N_9324,N_5866,N_4441);
nand U9325 (N_9325,N_4773,N_5363);
and U9326 (N_9326,N_3453,N_3480);
nor U9327 (N_9327,N_3621,N_4166);
nor U9328 (N_9328,N_5586,N_3347);
nor U9329 (N_9329,N_3258,N_3660);
nand U9330 (N_9330,N_3380,N_5907);
and U9331 (N_9331,N_5876,N_4328);
or U9332 (N_9332,N_5459,N_3240);
and U9333 (N_9333,N_3240,N_4859);
nand U9334 (N_9334,N_4717,N_5661);
xor U9335 (N_9335,N_5032,N_5526);
or U9336 (N_9336,N_5192,N_3341);
or U9337 (N_9337,N_3342,N_4764);
nor U9338 (N_9338,N_5821,N_4026);
nand U9339 (N_9339,N_4375,N_4181);
nand U9340 (N_9340,N_3411,N_5590);
xor U9341 (N_9341,N_4430,N_3212);
xor U9342 (N_9342,N_3797,N_5977);
xnor U9343 (N_9343,N_4605,N_3358);
and U9344 (N_9344,N_4803,N_4579);
and U9345 (N_9345,N_4150,N_4071);
xor U9346 (N_9346,N_5448,N_4523);
nor U9347 (N_9347,N_5578,N_3822);
nand U9348 (N_9348,N_3792,N_5497);
and U9349 (N_9349,N_6224,N_5065);
nor U9350 (N_9350,N_4003,N_5590);
nor U9351 (N_9351,N_4294,N_6189);
or U9352 (N_9352,N_3834,N_6027);
and U9353 (N_9353,N_5879,N_3408);
and U9354 (N_9354,N_5756,N_4065);
nand U9355 (N_9355,N_5578,N_5820);
or U9356 (N_9356,N_5248,N_5881);
and U9357 (N_9357,N_4617,N_6021);
and U9358 (N_9358,N_3877,N_4083);
xnor U9359 (N_9359,N_5490,N_5866);
nor U9360 (N_9360,N_5663,N_4981);
nand U9361 (N_9361,N_3876,N_3510);
nand U9362 (N_9362,N_3995,N_4576);
and U9363 (N_9363,N_5893,N_3343);
or U9364 (N_9364,N_5517,N_5563);
nand U9365 (N_9365,N_4509,N_5209);
nor U9366 (N_9366,N_5908,N_3807);
and U9367 (N_9367,N_5912,N_5577);
nor U9368 (N_9368,N_6179,N_6140);
xor U9369 (N_9369,N_3221,N_4837);
nor U9370 (N_9370,N_3912,N_3890);
nor U9371 (N_9371,N_4972,N_5051);
nor U9372 (N_9372,N_4597,N_5427);
nor U9373 (N_9373,N_4396,N_4683);
and U9374 (N_9374,N_3892,N_4782);
nand U9375 (N_9375,N_8254,N_8773);
or U9376 (N_9376,N_8082,N_8504);
xor U9377 (N_9377,N_9252,N_8041);
or U9378 (N_9378,N_6836,N_7930);
nor U9379 (N_9379,N_6995,N_7178);
or U9380 (N_9380,N_8793,N_7459);
nor U9381 (N_9381,N_8664,N_6280);
xor U9382 (N_9382,N_6657,N_8111);
nand U9383 (N_9383,N_8234,N_8830);
and U9384 (N_9384,N_8565,N_7355);
and U9385 (N_9385,N_9098,N_8892);
nand U9386 (N_9386,N_6669,N_7221);
and U9387 (N_9387,N_6962,N_8846);
and U9388 (N_9388,N_9031,N_6360);
or U9389 (N_9389,N_8491,N_6472);
and U9390 (N_9390,N_8095,N_7324);
nor U9391 (N_9391,N_7339,N_8995);
nor U9392 (N_9392,N_8979,N_6679);
nor U9393 (N_9393,N_7928,N_7916);
or U9394 (N_9394,N_7761,N_7822);
nor U9395 (N_9395,N_8774,N_7931);
and U9396 (N_9396,N_7310,N_6477);
nor U9397 (N_9397,N_8197,N_6466);
nor U9398 (N_9398,N_8649,N_6674);
or U9399 (N_9399,N_6482,N_6361);
or U9400 (N_9400,N_7697,N_8354);
nand U9401 (N_9401,N_8477,N_7535);
xnor U9402 (N_9402,N_8984,N_7924);
nand U9403 (N_9403,N_8790,N_8896);
nor U9404 (N_9404,N_9042,N_7584);
or U9405 (N_9405,N_8445,N_8609);
nand U9406 (N_9406,N_6831,N_8463);
or U9407 (N_9407,N_8129,N_7439);
nor U9408 (N_9408,N_7001,N_6368);
or U9409 (N_9409,N_9317,N_9193);
and U9410 (N_9410,N_8211,N_7243);
nor U9411 (N_9411,N_6964,N_8507);
nand U9412 (N_9412,N_7283,N_8668);
nor U9413 (N_9413,N_7389,N_7403);
nand U9414 (N_9414,N_8809,N_7060);
and U9415 (N_9415,N_9188,N_8673);
xnor U9416 (N_9416,N_7009,N_6814);
nor U9417 (N_9417,N_9244,N_8711);
and U9418 (N_9418,N_6906,N_8933);
or U9419 (N_9419,N_7643,N_7300);
xor U9420 (N_9420,N_7046,N_7981);
and U9421 (N_9421,N_6927,N_7621);
and U9422 (N_9422,N_8467,N_6733);
nand U9423 (N_9423,N_7586,N_8479);
xnor U9424 (N_9424,N_9243,N_8627);
or U9425 (N_9425,N_7017,N_6261);
nor U9426 (N_9426,N_8901,N_8065);
nand U9427 (N_9427,N_8781,N_7135);
nand U9428 (N_9428,N_6933,N_9358);
and U9429 (N_9429,N_6292,N_7566);
or U9430 (N_9430,N_6256,N_8575);
or U9431 (N_9431,N_7756,N_6849);
and U9432 (N_9432,N_8546,N_9223);
xnor U9433 (N_9433,N_7508,N_9204);
nor U9434 (N_9434,N_7190,N_8990);
or U9435 (N_9435,N_7932,N_9249);
and U9436 (N_9436,N_7701,N_8614);
or U9437 (N_9437,N_7502,N_6535);
nor U9438 (N_9438,N_9310,N_7296);
nor U9439 (N_9439,N_7679,N_8151);
and U9440 (N_9440,N_7765,N_7984);
xor U9441 (N_9441,N_6810,N_8561);
and U9442 (N_9442,N_8251,N_8438);
nor U9443 (N_9443,N_6608,N_6720);
and U9444 (N_9444,N_8223,N_7831);
xor U9445 (N_9445,N_6603,N_8114);
nand U9446 (N_9446,N_6808,N_8891);
nor U9447 (N_9447,N_8369,N_9112);
xor U9448 (N_9448,N_8521,N_8391);
nand U9449 (N_9449,N_9183,N_7220);
and U9450 (N_9450,N_7239,N_7342);
nor U9451 (N_9451,N_6526,N_7636);
xor U9452 (N_9452,N_8954,N_7742);
nand U9453 (N_9453,N_7232,N_7289);
nand U9454 (N_9454,N_6598,N_6834);
and U9455 (N_9455,N_7503,N_8998);
xnor U9456 (N_9456,N_7795,N_7019);
and U9457 (N_9457,N_8416,N_6916);
nand U9458 (N_9458,N_6681,N_7091);
nand U9459 (N_9459,N_7381,N_8124);
and U9460 (N_9460,N_8777,N_6764);
or U9461 (N_9461,N_8652,N_8909);
and U9462 (N_9462,N_8820,N_6485);
nor U9463 (N_9463,N_8838,N_7690);
nand U9464 (N_9464,N_9199,N_7315);
nand U9465 (N_9465,N_8269,N_8674);
and U9466 (N_9466,N_8178,N_9079);
nand U9467 (N_9467,N_7383,N_9116);
nor U9468 (N_9468,N_9080,N_6708);
xnor U9469 (N_9469,N_6353,N_7896);
or U9470 (N_9470,N_8196,N_8259);
or U9471 (N_9471,N_9076,N_7422);
nor U9472 (N_9472,N_8286,N_6787);
xnor U9473 (N_9473,N_7694,N_7734);
nand U9474 (N_9474,N_6772,N_7406);
or U9475 (N_9475,N_8028,N_7320);
nand U9476 (N_9476,N_6621,N_6542);
nand U9477 (N_9477,N_6401,N_7118);
nor U9478 (N_9478,N_6788,N_7732);
and U9479 (N_9479,N_9187,N_8572);
nor U9480 (N_9480,N_7787,N_8441);
nand U9481 (N_9481,N_7428,N_7707);
or U9482 (N_9482,N_6845,N_7559);
xnor U9483 (N_9483,N_6451,N_6682);
nand U9484 (N_9484,N_7337,N_9104);
nand U9485 (N_9485,N_9032,N_6832);
or U9486 (N_9486,N_8958,N_6464);
nand U9487 (N_9487,N_7969,N_7978);
and U9488 (N_9488,N_7045,N_8378);
nand U9489 (N_9489,N_6771,N_7730);
nor U9490 (N_9490,N_9304,N_7042);
or U9491 (N_9491,N_9290,N_8074);
and U9492 (N_9492,N_7581,N_8700);
nor U9493 (N_9493,N_9351,N_7868);
and U9494 (N_9494,N_9131,N_9364);
or U9495 (N_9495,N_6806,N_8540);
nor U9496 (N_9496,N_6984,N_9093);
and U9497 (N_9497,N_6650,N_7311);
xor U9498 (N_9498,N_7224,N_8358);
nor U9499 (N_9499,N_8603,N_7833);
and U9500 (N_9500,N_7478,N_6253);
and U9501 (N_9501,N_9040,N_7134);
or U9502 (N_9502,N_6884,N_8198);
and U9503 (N_9503,N_7014,N_8917);
nand U9504 (N_9504,N_7470,N_6615);
or U9505 (N_9505,N_6877,N_7915);
or U9506 (N_9506,N_6555,N_7628);
and U9507 (N_9507,N_7692,N_6308);
nor U9508 (N_9508,N_6726,N_6533);
nor U9509 (N_9509,N_8293,N_8537);
or U9510 (N_9510,N_7100,N_7211);
nand U9511 (N_9511,N_7662,N_6638);
or U9512 (N_9512,N_6700,N_8545);
and U9513 (N_9513,N_9319,N_6908);
and U9514 (N_9514,N_9258,N_8796);
and U9515 (N_9515,N_8877,N_8659);
or U9516 (N_9516,N_6851,N_8425);
nand U9517 (N_9517,N_7711,N_8621);
and U9518 (N_9518,N_6975,N_7321);
nor U9519 (N_9519,N_8840,N_7665);
or U9520 (N_9520,N_6564,N_7667);
nor U9521 (N_9521,N_7455,N_8771);
nand U9522 (N_9522,N_7480,N_7369);
xnor U9523 (N_9523,N_8133,N_6839);
nor U9524 (N_9524,N_8488,N_7361);
nor U9525 (N_9525,N_9232,N_8408);
or U9526 (N_9526,N_8157,N_8000);
and U9527 (N_9527,N_8719,N_6701);
and U9528 (N_9528,N_6854,N_6340);
and U9529 (N_9529,N_8233,N_9118);
or U9530 (N_9530,N_7533,N_8106);
xor U9531 (N_9531,N_7008,N_8138);
nor U9532 (N_9532,N_6479,N_7704);
xor U9533 (N_9533,N_7912,N_6795);
or U9534 (N_9534,N_8109,N_7033);
nor U9535 (N_9535,N_7563,N_6909);
or U9536 (N_9536,N_7805,N_6871);
nor U9537 (N_9537,N_7025,N_7929);
nor U9538 (N_9538,N_7029,N_6942);
nor U9539 (N_9539,N_6758,N_8505);
nand U9540 (N_9540,N_6568,N_6950);
nand U9541 (N_9541,N_9090,N_9009);
nand U9542 (N_9542,N_6566,N_9352);
and U9543 (N_9543,N_7316,N_6433);
nand U9544 (N_9544,N_7784,N_7307);
nand U9545 (N_9545,N_8515,N_8115);
nand U9546 (N_9546,N_7957,N_6958);
and U9547 (N_9547,N_7150,N_7780);
nand U9548 (N_9548,N_8553,N_8192);
nand U9549 (N_9549,N_6561,N_9006);
nand U9550 (N_9550,N_8769,N_8849);
and U9551 (N_9551,N_6302,N_7249);
nor U9552 (N_9552,N_7070,N_8193);
or U9553 (N_9553,N_6627,N_8583);
or U9554 (N_9554,N_7292,N_7467);
nor U9555 (N_9555,N_6548,N_6799);
xor U9556 (N_9556,N_7096,N_8607);
xor U9557 (N_9557,N_6362,N_6966);
and U9558 (N_9558,N_7461,N_6623);
xor U9559 (N_9559,N_7404,N_7479);
nor U9560 (N_9560,N_7652,N_8804);
nor U9561 (N_9561,N_8420,N_9095);
nor U9562 (N_9562,N_6759,N_8835);
nor U9563 (N_9563,N_7849,N_8025);
or U9564 (N_9564,N_8387,N_7565);
nor U9565 (N_9565,N_7631,N_8461);
nor U9566 (N_9566,N_6968,N_7672);
nand U9567 (N_9567,N_8271,N_9289);
nor U9568 (N_9568,N_7699,N_7886);
and U9569 (N_9569,N_7836,N_6949);
and U9570 (N_9570,N_6894,N_8883);
nor U9571 (N_9571,N_8320,N_9338);
nor U9572 (N_9572,N_7801,N_6296);
nand U9573 (N_9573,N_9221,N_7956);
nor U9574 (N_9574,N_8860,N_8745);
and U9575 (N_9575,N_7201,N_7858);
and U9576 (N_9576,N_7464,N_7166);
and U9577 (N_9577,N_9102,N_9019);
and U9578 (N_9578,N_8740,N_7917);
and U9579 (N_9579,N_6835,N_7774);
nor U9580 (N_9580,N_7641,N_8119);
nand U9581 (N_9581,N_6637,N_8520);
xnor U9582 (N_9582,N_8534,N_6318);
nor U9583 (N_9583,N_7154,N_6571);
nand U9584 (N_9584,N_8353,N_6811);
xor U9585 (N_9585,N_9328,N_7791);
and U9586 (N_9586,N_7825,N_7106);
and U9587 (N_9587,N_7673,N_7866);
or U9588 (N_9588,N_7781,N_7510);
nor U9589 (N_9589,N_9343,N_6605);
nand U9590 (N_9590,N_6889,N_6418);
and U9591 (N_9591,N_6512,N_7299);
nand U9592 (N_9592,N_8448,N_9302);
and U9593 (N_9593,N_7813,N_7645);
and U9594 (N_9594,N_7173,N_7995);
nand U9595 (N_9595,N_6519,N_6596);
or U9596 (N_9596,N_8924,N_7907);
or U9597 (N_9597,N_6928,N_7577);
or U9598 (N_9598,N_8871,N_6945);
or U9599 (N_9599,N_6746,N_9155);
xor U9600 (N_9600,N_7233,N_6738);
nand U9601 (N_9601,N_6915,N_8310);
and U9602 (N_9602,N_8619,N_7192);
nand U9603 (N_9603,N_7326,N_7855);
xor U9604 (N_9604,N_8303,N_8181);
and U9605 (N_9605,N_6996,N_6595);
nand U9606 (N_9606,N_6777,N_8201);
nor U9607 (N_9607,N_6973,N_8688);
nor U9608 (N_9608,N_8337,N_9146);
nor U9609 (N_9609,N_8007,N_7823);
and U9610 (N_9610,N_9354,N_7397);
or U9611 (N_9611,N_6475,N_6752);
nand U9612 (N_9612,N_6429,N_7020);
nor U9613 (N_9613,N_7696,N_8362);
xnor U9614 (N_9614,N_8004,N_9371);
nor U9615 (N_9615,N_7132,N_8168);
and U9616 (N_9616,N_8383,N_6689);
nor U9617 (N_9617,N_7513,N_6807);
nor U9618 (N_9618,N_9287,N_7114);
or U9619 (N_9619,N_7927,N_8380);
nor U9620 (N_9620,N_9194,N_7555);
or U9621 (N_9621,N_7773,N_9361);
nor U9622 (N_9622,N_6287,N_8925);
and U9623 (N_9623,N_7741,N_7890);
and U9624 (N_9624,N_7517,N_7380);
and U9625 (N_9625,N_9096,N_8724);
nand U9626 (N_9626,N_6597,N_7658);
and U9627 (N_9627,N_8921,N_9129);
xnor U9628 (N_9628,N_6447,N_6270);
or U9629 (N_9629,N_7259,N_9094);
nor U9630 (N_9630,N_7573,N_8356);
nand U9631 (N_9631,N_6502,N_7015);
nand U9632 (N_9632,N_8913,N_8024);
nand U9633 (N_9633,N_7514,N_7094);
or U9634 (N_9634,N_6667,N_9219);
nand U9635 (N_9635,N_7184,N_8512);
and U9636 (N_9636,N_7427,N_8890);
nand U9637 (N_9637,N_6794,N_9333);
and U9638 (N_9638,N_6747,N_7706);
nor U9639 (N_9639,N_7038,N_8381);
nand U9640 (N_9640,N_9298,N_8671);
or U9641 (N_9641,N_9058,N_6986);
nor U9642 (N_9642,N_9119,N_7417);
and U9643 (N_9643,N_9161,N_8847);
nor U9644 (N_9644,N_7893,N_7494);
or U9645 (N_9645,N_8173,N_6873);
and U9646 (N_9646,N_7169,N_9253);
nor U9647 (N_9647,N_7052,N_8685);
or U9648 (N_9648,N_6969,N_7269);
nor U9649 (N_9649,N_6818,N_7497);
nand U9650 (N_9650,N_9245,N_9332);
nand U9651 (N_9651,N_7241,N_7161);
nor U9652 (N_9652,N_9149,N_7608);
nand U9653 (N_9653,N_9173,N_7772);
or U9654 (N_9654,N_9145,N_7605);
nand U9655 (N_9655,N_7212,N_7953);
nor U9656 (N_9656,N_7343,N_8529);
xor U9657 (N_9657,N_6768,N_6357);
and U9658 (N_9658,N_8312,N_6396);
nand U9659 (N_9659,N_7465,N_8524);
and U9660 (N_9660,N_8910,N_6859);
xnor U9661 (N_9661,N_7314,N_7804);
or U9662 (N_9662,N_7340,N_6328);
xnor U9663 (N_9663,N_8655,N_9097);
nand U9664 (N_9664,N_8404,N_8350);
and U9665 (N_9665,N_6983,N_8042);
and U9666 (N_9666,N_7058,N_8606);
nand U9667 (N_9667,N_8828,N_7487);
or U9668 (N_9668,N_6640,N_7590);
or U9669 (N_9669,N_8530,N_8329);
and U9670 (N_9670,N_9089,N_8516);
nand U9671 (N_9671,N_9336,N_7705);
nor U9672 (N_9672,N_6351,N_6952);
nor U9673 (N_9673,N_7377,N_7121);
nor U9674 (N_9674,N_9132,N_8451);
and U9675 (N_9675,N_7031,N_7585);
nand U9676 (N_9676,N_9138,N_6581);
nor U9677 (N_9677,N_8807,N_7285);
nor U9678 (N_9678,N_8142,N_6293);
and U9679 (N_9679,N_7944,N_7724);
and U9680 (N_9680,N_6670,N_7685);
xor U9681 (N_9681,N_8699,N_9053);
nor U9682 (N_9682,N_8429,N_6522);
nand U9683 (N_9683,N_7830,N_8826);
nor U9684 (N_9684,N_7098,N_8570);
and U9685 (N_9685,N_6792,N_9108);
xor U9686 (N_9686,N_9197,N_7575);
and U9687 (N_9687,N_7204,N_9350);
nor U9688 (N_9688,N_6658,N_8418);
and U9689 (N_9689,N_8940,N_6900);
xor U9690 (N_9690,N_7264,N_7617);
nor U9691 (N_9691,N_7670,N_7053);
nand U9692 (N_9692,N_7208,N_8812);
and U9693 (N_9693,N_8704,N_7452);
and U9694 (N_9694,N_7133,N_9230);
and U9695 (N_9695,N_7165,N_7681);
or U9696 (N_9696,N_7758,N_8856);
and U9697 (N_9697,N_9224,N_6523);
and U9698 (N_9698,N_7542,N_7153);
nor U9699 (N_9699,N_7164,N_7295);
nand U9700 (N_9700,N_6745,N_9140);
nor U9701 (N_9701,N_8236,N_8815);
and U9702 (N_9702,N_8803,N_8047);
and U9703 (N_9703,N_6826,N_6599);
xnor U9704 (N_9704,N_6677,N_9265);
nor U9705 (N_9705,N_6718,N_8935);
nand U9706 (N_9706,N_7217,N_7576);
nand U9707 (N_9707,N_9251,N_7659);
or U9708 (N_9708,N_8968,N_7602);
and U9709 (N_9709,N_6407,N_9022);
xor U9710 (N_9710,N_6980,N_8229);
nor U9711 (N_9711,N_8278,N_8772);
nor U9712 (N_9712,N_7237,N_8411);
nor U9713 (N_9713,N_8283,N_7867);
nand U9714 (N_9714,N_8232,N_6757);
and U9715 (N_9715,N_6749,N_7941);
and U9716 (N_9716,N_8205,N_8795);
nor U9717 (N_9717,N_8373,N_7595);
nor U9718 (N_9718,N_7401,N_8348);
and U9719 (N_9719,N_9303,N_8499);
nand U9720 (N_9720,N_6532,N_8349);
and U9721 (N_9721,N_6487,N_7789);
or U9722 (N_9722,N_7994,N_8122);
or U9723 (N_9723,N_7888,N_6730);
nand U9724 (N_9724,N_7538,N_7609);
nor U9725 (N_9725,N_8919,N_9068);
nor U9726 (N_9726,N_6323,N_8947);
or U9727 (N_9727,N_7828,N_6629);
nand U9728 (N_9728,N_7446,N_9267);
or U9729 (N_9729,N_8611,N_8069);
nor U9730 (N_9730,N_6993,N_7368);
and U9731 (N_9731,N_8599,N_9105);
nand U9732 (N_9732,N_8029,N_8675);
nor U9733 (N_9733,N_6886,N_7272);
nand U9734 (N_9734,N_8666,N_8296);
xnor U9735 (N_9735,N_9099,N_7733);
or U9736 (N_9736,N_7718,N_7829);
nor U9737 (N_9737,N_9296,N_6506);
nand U9738 (N_9738,N_8249,N_7714);
xor U9739 (N_9739,N_8975,N_7796);
and U9740 (N_9740,N_9218,N_9003);
nand U9741 (N_9741,N_7883,N_6286);
or U9742 (N_9742,N_9142,N_9266);
and U9743 (N_9743,N_7005,N_9020);
nand U9744 (N_9744,N_9049,N_7587);
and U9745 (N_9745,N_7968,N_8426);
nand U9746 (N_9746,N_8336,N_7543);
or U9747 (N_9747,N_8153,N_7751);
nand U9748 (N_9748,N_8123,N_6661);
or U9749 (N_9749,N_9081,N_7122);
and U9750 (N_9750,N_6630,N_6279);
nand U9751 (N_9751,N_8727,N_8757);
and U9752 (N_9752,N_6940,N_7443);
or U9753 (N_9753,N_6514,N_6520);
nor U9754 (N_9754,N_8118,N_9348);
nor U9755 (N_9755,N_8893,N_6529);
or U9756 (N_9756,N_7350,N_8839);
and U9757 (N_9757,N_7170,N_7640);
nand U9758 (N_9758,N_7878,N_8152);
or U9759 (N_9759,N_8385,N_8459);
or U9760 (N_9760,N_9167,N_8942);
nand U9761 (N_9761,N_8698,N_7261);
or U9762 (N_9762,N_8615,N_8055);
nand U9763 (N_9763,N_7485,N_6312);
or U9764 (N_9764,N_8985,N_8214);
or U9765 (N_9765,N_8261,N_9181);
or U9766 (N_9766,N_6705,N_8932);
nand U9767 (N_9767,N_6363,N_7319);
and U9768 (N_9768,N_6699,N_8315);
nor U9769 (N_9769,N_9176,N_8334);
nor U9770 (N_9770,N_8552,N_7421);
nor U9771 (N_9771,N_8147,N_6865);
nor U9772 (N_9772,N_6815,N_8183);
or U9773 (N_9773,N_7140,N_6303);
nor U9774 (N_9774,N_7936,N_7660);
or U9775 (N_9775,N_7372,N_9048);
and U9776 (N_9776,N_7356,N_9226);
nor U9777 (N_9777,N_6731,N_8368);
nand U9778 (N_9778,N_6271,N_6925);
nand U9779 (N_9779,N_7528,N_9077);
xnor U9780 (N_9780,N_6741,N_9008);
xnor U9781 (N_9781,N_6707,N_7909);
and U9782 (N_9782,N_8978,N_7144);
nand U9783 (N_9783,N_7007,N_7861);
nor U9784 (N_9784,N_7024,N_7882);
or U9785 (N_9785,N_7352,N_6493);
or U9786 (N_9786,N_6591,N_9311);
and U9787 (N_9787,N_6497,N_7934);
nand U9788 (N_9788,N_7599,N_9247);
or U9789 (N_9789,N_8616,N_7477);
nand U9790 (N_9790,N_7183,N_8590);
and U9791 (N_9791,N_6546,N_7719);
and U9792 (N_9792,N_7899,N_7998);
or U9793 (N_9793,N_6467,N_7203);
nand U9794 (N_9794,N_7120,N_6651);
nor U9795 (N_9795,N_7838,N_6724);
xor U9796 (N_9796,N_7580,N_7702);
xor U9797 (N_9797,N_7454,N_9050);
nand U9798 (N_9798,N_7540,N_8658);
xor U9799 (N_9799,N_6635,N_8983);
nor U9800 (N_9800,N_6306,N_7364);
and U9801 (N_9801,N_8228,N_9016);
nor U9802 (N_9802,N_7398,N_6920);
and U9803 (N_9803,N_8339,N_6305);
and U9804 (N_9804,N_9214,N_6498);
and U9805 (N_9805,N_8474,N_8372);
nor U9806 (N_9806,N_8185,N_6450);
or U9807 (N_9807,N_8881,N_7630);
nor U9808 (N_9808,N_6404,N_6486);
nand U9809 (N_9809,N_7971,N_6489);
or U9810 (N_9810,N_9257,N_8920);
and U9811 (N_9811,N_6402,N_8478);
and U9812 (N_9812,N_8766,N_8367);
or U9813 (N_9813,N_9159,N_6592);
nor U9814 (N_9814,N_8876,N_7095);
nand U9815 (N_9815,N_7044,N_9270);
and U9816 (N_9816,N_7954,N_8021);
xnor U9817 (N_9817,N_7149,N_8440);
or U9818 (N_9818,N_8470,N_6926);
or U9819 (N_9819,N_8117,N_8725);
nor U9820 (N_9820,N_7466,N_7570);
nand U9821 (N_9821,N_8579,N_8916);
and U9822 (N_9822,N_8489,N_6510);
nor U9823 (N_9823,N_7414,N_9337);
nor U9824 (N_9824,N_6773,N_9010);
and U9825 (N_9825,N_9153,N_8464);
nand U9826 (N_9826,N_7457,N_8255);
and U9827 (N_9827,N_8882,N_8669);
or U9828 (N_9828,N_7552,N_7088);
and U9829 (N_9829,N_8798,N_9029);
and U9830 (N_9830,N_6391,N_8842);
and U9831 (N_9831,N_6255,N_8297);
and U9832 (N_9832,N_8389,N_7554);
and U9833 (N_9833,N_6524,N_7275);
nor U9834 (N_9834,N_6992,N_7843);
nand U9835 (N_9835,N_8172,N_7418);
and U9836 (N_9836,N_9217,N_7683);
nand U9837 (N_9837,N_9373,N_8285);
nor U9838 (N_9838,N_7491,N_6505);
nor U9839 (N_9839,N_8639,N_9115);
or U9840 (N_9840,N_6999,N_6582);
or U9841 (N_9841,N_8080,N_7752);
nor U9842 (N_9842,N_6517,N_8099);
nand U9843 (N_9843,N_7354,N_9255);
xor U9844 (N_9844,N_7964,N_8326);
or U9845 (N_9845,N_8816,N_7755);
and U9846 (N_9846,N_6342,N_7877);
xnor U9847 (N_9847,N_7923,N_9201);
nand U9848 (N_9848,N_8098,N_8006);
xor U9849 (N_9849,N_8038,N_9154);
or U9850 (N_9850,N_7816,N_7400);
or U9851 (N_9851,N_6266,N_7790);
xor U9852 (N_9852,N_8146,N_8061);
nand U9853 (N_9853,N_7175,N_9300);
or U9854 (N_9854,N_7327,N_6574);
and U9855 (N_9855,N_6567,N_8805);
xor U9856 (N_9856,N_7030,N_8050);
or U9857 (N_9857,N_7278,N_6725);
xnor U9858 (N_9858,N_8309,N_6899);
nor U9859 (N_9859,N_9122,N_7198);
or U9860 (N_9860,N_8075,N_6508);
or U9861 (N_9861,N_8056,N_6366);
and U9862 (N_9862,N_8783,N_6763);
or U9863 (N_9863,N_9178,N_8643);
or U9864 (N_9864,N_8057,N_9370);
and U9865 (N_9865,N_6994,N_6437);
nand U9866 (N_9866,N_6878,N_8681);
and U9867 (N_9867,N_6300,N_7903);
nor U9868 (N_9868,N_8895,N_6501);
or U9869 (N_9869,N_9242,N_6837);
and U9870 (N_9870,N_7073,N_6728);
and U9871 (N_9871,N_6495,N_7210);
nor U9872 (N_9872,N_8810,N_9210);
or U9873 (N_9873,N_7983,N_9086);
nor U9874 (N_9874,N_8403,N_7181);
or U9875 (N_9875,N_6552,N_9134);
nand U9876 (N_9876,N_6272,N_9241);
nand U9877 (N_9877,N_7783,N_8247);
and U9878 (N_9878,N_6978,N_7688);
and U9879 (N_9879,N_8102,N_6632);
nand U9880 (N_9880,N_9164,N_7469);
nand U9881 (N_9881,N_8903,N_6710);
and U9882 (N_9882,N_8299,N_7196);
or U9883 (N_9883,N_8511,N_8015);
nor U9884 (N_9884,N_7193,N_8600);
nor U9885 (N_9885,N_7474,N_6696);
or U9886 (N_9886,N_7553,N_7200);
or U9887 (N_9887,N_8508,N_8227);
or U9888 (N_9888,N_8322,N_7698);
and U9889 (N_9889,N_7571,N_9260);
nand U9890 (N_9890,N_9182,N_8898);
and U9891 (N_9891,N_6919,N_8087);
or U9892 (N_9892,N_8595,N_8884);
xor U9893 (N_9893,N_9309,N_6676);
and U9894 (N_9894,N_8419,N_7809);
nor U9895 (N_9895,N_7386,N_8313);
and U9896 (N_9896,N_9240,N_8116);
and U9897 (N_9897,N_6860,N_8394);
and U9898 (N_9898,N_7146,N_6671);
nand U9899 (N_9899,N_6833,N_6703);
or U9900 (N_9900,N_7256,N_7139);
nor U9901 (N_9901,N_7126,N_7717);
or U9902 (N_9902,N_8889,N_8813);
nand U9903 (N_9903,N_8242,N_8557);
and U9904 (N_9904,N_6584,N_9367);
nor U9905 (N_9905,N_7441,N_7358);
nor U9906 (N_9906,N_7982,N_6324);
or U9907 (N_9907,N_7509,N_9206);
nand U9908 (N_9908,N_9281,N_6686);
and U9909 (N_9909,N_9314,N_9141);
nand U9910 (N_9910,N_7876,N_9156);
and U9911 (N_9911,N_8638,N_8585);
xnor U9912 (N_9912,N_8861,N_9121);
xor U9913 (N_9913,N_7650,N_8376);
nand U9914 (N_9914,N_8494,N_6488);
xor U9915 (N_9915,N_7786,N_8415);
nand U9916 (N_9916,N_7384,N_6715);
nand U9917 (N_9917,N_9023,N_9360);
and U9918 (N_9918,N_9035,N_6939);
and U9919 (N_9919,N_8154,N_6379);
and U9920 (N_9920,N_8714,N_8171);
nor U9921 (N_9921,N_7817,N_8780);
nand U9922 (N_9922,N_8991,N_6456);
or U9923 (N_9923,N_9363,N_6770);
nand U9924 (N_9924,N_6905,N_7056);
nor U9925 (N_9925,N_6327,N_7715);
and U9926 (N_9926,N_7062,N_7304);
or U9927 (N_9927,N_7639,N_8741);
nor U9928 (N_9928,N_8155,N_9174);
xor U9929 (N_9929,N_6371,N_7202);
or U9930 (N_9930,N_6652,N_6822);
and U9931 (N_9931,N_8295,N_7280);
nand U9932 (N_9932,N_7946,N_8943);
and U9933 (N_9933,N_9374,N_9372);
nor U9934 (N_9934,N_6453,N_8718);
xnor U9935 (N_9935,N_9238,N_7504);
or U9936 (N_9936,N_9101,N_8905);
nand U9937 (N_9937,N_7048,N_7392);
nand U9938 (N_9938,N_6449,N_7567);
and U9939 (N_9939,N_9128,N_8260);
and U9940 (N_9940,N_8684,N_6474);
nand U9941 (N_9941,N_7856,N_9045);
xnor U9942 (N_9942,N_8859,N_8879);
nor U9943 (N_9943,N_7996,N_6979);
nor U9944 (N_9944,N_7837,N_6283);
or U9945 (N_9945,N_8974,N_6706);
nand U9946 (N_9946,N_7716,N_6572);
and U9947 (N_9947,N_7875,N_9269);
or U9948 (N_9948,N_7616,N_9066);
nand U9949 (N_9949,N_7764,N_7709);
or U9950 (N_9950,N_7000,N_8645);
and U9951 (N_9951,N_7874,N_8928);
xor U9952 (N_9952,N_6478,N_8164);
nand U9953 (N_9953,N_7760,N_8219);
nor U9954 (N_9954,N_7558,N_7093);
or U9955 (N_9955,N_9120,N_6876);
nand U9956 (N_9956,N_7735,N_9323);
nor U9957 (N_9957,N_6672,N_7090);
or U9958 (N_9958,N_7408,N_7853);
xor U9959 (N_9959,N_9166,N_8215);
and U9960 (N_9960,N_9327,N_8574);
xor U9961 (N_9961,N_6325,N_8706);
nor U9962 (N_9962,N_8651,N_7537);
or U9963 (N_9963,N_7505,N_8314);
nand U9964 (N_9964,N_8970,N_8735);
and U9965 (N_9965,N_6589,N_6298);
nor U9966 (N_9966,N_7530,N_7574);
and U9967 (N_9967,N_6816,N_9114);
nor U9968 (N_9968,N_7610,N_8043);
nand U9969 (N_9969,N_8641,N_8982);
nor U9970 (N_9970,N_9005,N_7227);
and U9971 (N_9971,N_7965,N_6365);
nand U9972 (N_9972,N_6403,N_9286);
xor U9973 (N_9973,N_7824,N_8137);
nor U9974 (N_9974,N_7745,N_7661);
nor U9975 (N_9975,N_7177,N_7821);
nand U9976 (N_9976,N_9228,N_7238);
or U9977 (N_9977,N_7152,N_8680);
xnor U9978 (N_9978,N_6307,N_8981);
and U9979 (N_9979,N_8068,N_6330);
nand U9980 (N_9980,N_9069,N_7394);
nor U9981 (N_9981,N_7865,N_7050);
and U9982 (N_9982,N_6395,N_7591);
and U9983 (N_9983,N_8731,N_7747);
nand U9984 (N_9984,N_8190,N_9231);
or U9985 (N_9985,N_8127,N_8654);
nand U9986 (N_9986,N_9106,N_7156);
or U9987 (N_9987,N_7128,N_7666);
and U9988 (N_9988,N_9170,N_9339);
and U9989 (N_9989,N_6499,N_9103);
and U9990 (N_9990,N_6269,N_9130);
nor U9991 (N_9991,N_8571,N_8084);
nor U9992 (N_9992,N_7379,N_7107);
and U9993 (N_9993,N_7894,N_9057);
and U9994 (N_9994,N_6294,N_7084);
or U9995 (N_9995,N_8836,N_7960);
xor U9996 (N_9996,N_8132,N_8092);
nor U9997 (N_9997,N_6709,N_6694);
nor U9998 (N_9998,N_7619,N_8258);
nand U9999 (N_9999,N_7881,N_7648);
or U10000 (N_10000,N_9250,N_7072);
or U10001 (N_10001,N_7099,N_7157);
or U10002 (N_10002,N_8677,N_7473);
or U10003 (N_10003,N_8993,N_7112);
xor U10004 (N_10004,N_7080,N_7318);
nand U10005 (N_10005,N_8063,N_6869);
xnor U10006 (N_10006,N_7252,N_6735);
and U10007 (N_10007,N_7075,N_8811);
xnor U10008 (N_10008,N_8687,N_7351);
xnor U10009 (N_10009,N_8656,N_6610);
nand U10010 (N_10010,N_8434,N_6431);
nand U10011 (N_10011,N_7950,N_8427);
nand U10012 (N_10012,N_7832,N_7972);
and U10013 (N_10013,N_8591,N_9222);
nand U10014 (N_10014,N_8272,N_7897);
nor U10015 (N_10015,N_9148,N_6419);
nor U10016 (N_10016,N_6383,N_8179);
nor U10017 (N_10017,N_9212,N_7642);
xnor U10018 (N_10018,N_8386,N_8855);
nor U10019 (N_10019,N_6974,N_8778);
nor U10020 (N_10020,N_7271,N_6793);
nand U10021 (N_10021,N_8421,N_8747);
or U10022 (N_10022,N_8203,N_6740);
nand U10023 (N_10023,N_8160,N_7245);
or U10024 (N_10024,N_8238,N_6753);
or U10025 (N_10025,N_7782,N_6847);
nand U10026 (N_10026,N_7651,N_6516);
or U10027 (N_10027,N_6855,N_8103);
or U10028 (N_10028,N_8276,N_6617);
and U10029 (N_10029,N_8189,N_9144);
and U10030 (N_10030,N_9056,N_6825);
nand U10031 (N_10031,N_9011,N_8829);
or U10032 (N_10032,N_6476,N_9043);
nand U10033 (N_10033,N_8485,N_8325);
nand U10034 (N_10034,N_8946,N_8857);
or U10035 (N_10035,N_7250,N_7163);
nand U10036 (N_10036,N_7626,N_8869);
nand U10037 (N_10037,N_6461,N_8945);
nor U10038 (N_10038,N_7810,N_8141);
or U10039 (N_10039,N_8904,N_7223);
or U10040 (N_10040,N_8163,N_8662);
nand U10041 (N_10041,N_9021,N_8246);
nand U10042 (N_10042,N_7738,N_7199);
xnor U10043 (N_10043,N_8010,N_8934);
nor U10044 (N_10044,N_6415,N_6620);
and U10045 (N_10045,N_7597,N_9111);
or U10046 (N_10046,N_6742,N_7004);
nor U10047 (N_10047,N_7914,N_6848);
or U10048 (N_10048,N_7815,N_8832);
and U10049 (N_10049,N_9185,N_8513);
and U10050 (N_10050,N_8469,N_6693);
or U10051 (N_10051,N_7607,N_6444);
nor U10052 (N_10052,N_7197,N_6463);
nand U10053 (N_10053,N_7850,N_7247);
nand U10054 (N_10054,N_7059,N_9365);
nand U10055 (N_10055,N_7942,N_6883);
and U10056 (N_10056,N_9263,N_6755);
nand U10057 (N_10057,N_7357,N_7536);
and U10058 (N_10058,N_6424,N_6767);
nand U10059 (N_10059,N_8967,N_6989);
nand U10060 (N_10060,N_7425,N_7130);
nand U10061 (N_10061,N_7812,N_7412);
and U10062 (N_10062,N_6769,N_6583);
and U10063 (N_10063,N_9294,N_6697);
nand U10064 (N_10064,N_8049,N_9073);
nor U10065 (N_10065,N_7449,N_8927);
nor U10066 (N_10066,N_8617,N_7328);
nand U10067 (N_10067,N_8475,N_6376);
or U10068 (N_10068,N_8424,N_7794);
nand U10069 (N_10069,N_6304,N_7424);
xnor U10070 (N_10070,N_6911,N_7159);
and U10071 (N_10071,N_6954,N_7490);
xnor U10072 (N_10072,N_7129,N_8188);
or U10073 (N_10073,N_7647,N_8961);
or U10074 (N_10074,N_6783,N_7797);
nor U10075 (N_10075,N_8723,N_9124);
nand U10076 (N_10076,N_7322,N_8333);
or U10077 (N_10077,N_7363,N_6500);
nand U10078 (N_10078,N_7689,N_6665);
nand U10079 (N_10079,N_8751,N_8094);
nor U10080 (N_10080,N_9236,N_7294);
and U10081 (N_10081,N_6496,N_8756);
or U10082 (N_10082,N_9297,N_7979);
nand U10083 (N_10083,N_7993,N_9059);
nor U10084 (N_10084,N_9334,N_6471);
or U10085 (N_10085,N_8490,N_9172);
and U10086 (N_10086,N_9109,N_9169);
xnor U10087 (N_10087,N_7228,N_6341);
nand U10088 (N_10088,N_8789,N_9345);
nand U10089 (N_10089,N_7977,N_6369);
xor U10090 (N_10090,N_8739,N_8208);
and U10091 (N_10091,N_8046,N_8779);
nand U10092 (N_10092,N_8289,N_8212);
or U10093 (N_10093,N_6577,N_7123);
or U10094 (N_10094,N_6963,N_8560);
nor U10095 (N_10095,N_8060,N_6872);
nor U10096 (N_10096,N_9271,N_9203);
nand U10097 (N_10097,N_7240,N_6554);
or U10098 (N_10098,N_8863,N_7989);
and U10099 (N_10099,N_9133,N_6675);
nand U10100 (N_10100,N_8519,N_6609);
xor U10101 (N_10101,N_6481,N_9028);
and U10102 (N_10102,N_6530,N_8317);
nand U10103 (N_10103,N_6455,N_8964);
and U10104 (N_10104,N_7393,N_6800);
nand U10105 (N_10105,N_8800,N_6299);
nor U10106 (N_10106,N_6712,N_7757);
or U10107 (N_10107,N_7303,N_7612);
xnor U10108 (N_10108,N_8096,N_7880);
or U10109 (N_10109,N_7803,N_8407);
and U10110 (N_10110,N_7305,N_9051);
nor U10111 (N_10111,N_7918,N_8417);
xor U10112 (N_10112,N_8527,N_8013);
and U10113 (N_10113,N_7986,N_8626);
or U10114 (N_10114,N_8506,N_8589);
nand U10115 (N_10115,N_7776,N_6587);
nand U10116 (N_10116,N_8447,N_6515);
and U10117 (N_10117,N_6547,N_7744);
or U10118 (N_10118,N_9279,N_7174);
nor U10119 (N_10119,N_8086,N_8678);
nand U10120 (N_10120,N_7426,N_9233);
nor U10121 (N_10121,N_6662,N_6852);
xor U10122 (N_10122,N_8253,N_6887);
nor U10123 (N_10123,N_8323,N_9330);
or U10124 (N_10124,N_6985,N_8392);
or U10125 (N_10125,N_8690,N_7353);
xor U10126 (N_10126,N_7396,N_6760);
nor U10127 (N_10127,N_7472,N_8413);
and U10128 (N_10128,N_8493,N_8401);
nand U10129 (N_10129,N_8868,N_7185);
nor U10130 (N_10130,N_7625,N_7677);
xor U10131 (N_10131,N_8097,N_8598);
and U10132 (N_10132,N_6879,N_7460);
or U10133 (N_10133,N_8722,N_8539);
and U10134 (N_10134,N_8709,N_9284);
nand U10135 (N_10135,N_6678,N_6684);
and U10136 (N_10136,N_6277,N_7545);
xor U10137 (N_10137,N_9034,N_7468);
nor U10138 (N_10138,N_8629,N_8280);
and U10139 (N_10139,N_7276,N_9313);
or U10140 (N_10140,N_7622,N_8548);
nor U10141 (N_10141,N_7057,N_8195);
or U10142 (N_10142,N_7298,N_7101);
xnor U10143 (N_10143,N_6727,N_8184);
or U10144 (N_10144,N_8263,N_7458);
nor U10145 (N_10145,N_8547,N_8170);
xor U10146 (N_10146,N_9225,N_7655);
xnor U10147 (N_10147,N_8582,N_7870);
nor U10148 (N_10148,N_6440,N_8498);
nor U10149 (N_10149,N_7365,N_6698);
and U10150 (N_10150,N_9200,N_9085);
nand U10151 (N_10151,N_7451,N_8937);
or U10152 (N_10152,N_8588,N_8344);
or U10153 (N_10153,N_9190,N_7507);
or U10154 (N_10154,N_7518,N_8931);
nand U10155 (N_10155,N_8300,N_8977);
xor U10156 (N_10156,N_6990,N_9292);
and U10157 (N_10157,N_6938,N_7671);
xor U10158 (N_10158,N_9002,N_7726);
nor U10159 (N_10159,N_8737,N_8594);
nor U10160 (N_10160,N_6624,N_6893);
xor U10161 (N_10161,N_8031,N_8858);
nor U10162 (N_10162,N_9301,N_7061);
or U10163 (N_10163,N_9322,N_7959);
nand U10164 (N_10164,N_7919,N_8457);
or U10165 (N_10165,N_6625,N_6820);
and U10166 (N_10166,N_9033,N_7205);
and U10167 (N_10167,N_7656,N_6976);
and U10168 (N_10168,N_9283,N_8483);
or U10169 (N_10169,N_7047,N_6690);
nor U10170 (N_10170,N_8532,N_7043);
nand U10171 (N_10171,N_8481,N_8471);
or U10172 (N_10172,N_6531,N_6646);
nand U10173 (N_10173,N_8083,N_9060);
nor U10174 (N_10174,N_8637,N_7325);
nor U10175 (N_10175,N_9036,N_7862);
nor U10176 (N_10176,N_8555,N_8576);
nor U10177 (N_10177,N_6483,N_8156);
nand U10178 (N_10178,N_7022,N_8235);
and U10179 (N_10179,N_7785,N_8566);
nor U10180 (N_10180,N_6673,N_8237);
or U10181 (N_10181,N_7119,N_9039);
nand U10182 (N_10182,N_7219,N_6405);
and U10183 (N_10183,N_7889,N_6882);
or U10184 (N_10184,N_7207,N_6411);
or U10185 (N_10185,N_7432,N_7945);
or U10186 (N_10186,N_7527,N_7871);
or U10187 (N_10187,N_7054,N_7270);
nor U10188 (N_10188,N_9084,N_7708);
nand U10189 (N_10189,N_8134,N_6441);
nand U10190 (N_10190,N_7799,N_9278);
nand U10191 (N_10191,N_8100,N_7712);
or U10192 (N_10192,N_8697,N_6917);
or U10193 (N_10193,N_7967,N_8437);
nor U10194 (N_10194,N_8186,N_8768);
and U10195 (N_10195,N_6413,N_6830);
nand U10196 (N_10196,N_7814,N_6864);
nand U10197 (N_10197,N_8587,N_6473);
nand U10198 (N_10198,N_7431,N_8672);
nor U10199 (N_10199,N_9165,N_6394);
nand U10200 (N_10200,N_6563,N_7811);
nor U10201 (N_10201,N_7083,N_8482);
nor U10202 (N_10202,N_8039,N_8716);
or U10203 (N_10203,N_6345,N_6784);
or U10204 (N_10204,N_8396,N_7568);
xor U10205 (N_10205,N_7331,N_7179);
nand U10206 (N_10206,N_8694,N_6704);
xor U10207 (N_10207,N_7669,N_9237);
xor U10208 (N_10208,N_9065,N_6812);
xnor U10209 (N_10209,N_9100,N_6503);
nand U10210 (N_10210,N_7332,N_6936);
or U10211 (N_10211,N_7087,N_7973);
nor U10212 (N_10212,N_8110,N_7333);
and U10213 (N_10213,N_7359,N_6842);
nor U10214 (N_10214,N_8433,N_8077);
and U10215 (N_10215,N_7988,N_6492);
and U10216 (N_10216,N_6998,N_9234);
or U10217 (N_10217,N_7006,N_7182);
nor U10218 (N_10218,N_7023,N_7063);
nor U10219 (N_10219,N_7230,N_6649);
nor U10220 (N_10220,N_9012,N_7347);
or U10221 (N_10221,N_8085,N_7703);
or U10222 (N_10222,N_7792,N_6354);
nand U10223 (N_10223,N_8128,N_6774);
nor U10224 (N_10224,N_7036,N_6525);
nand U10225 (N_10225,N_6438,N_7588);
and U10226 (N_10226,N_8107,N_7103);
and U10227 (N_10227,N_7693,N_7556);
and U10228 (N_10228,N_8355,N_6721);
nand U10229 (N_10229,N_8562,N_7255);
nor U10230 (N_10230,N_6813,N_8026);
and U10231 (N_10231,N_7113,N_6902);
and U10232 (N_10232,N_7955,N_6372);
and U10233 (N_10233,N_8878,N_7990);
nor U10234 (N_10234,N_8708,N_7547);
nor U10235 (N_10235,N_7160,N_8872);
and U10236 (N_10236,N_8176,N_8833);
nor U10237 (N_10237,N_7137,N_8536);
and U10238 (N_10238,N_8458,N_7700);
nor U10239 (N_10239,N_6853,N_7102);
nand U10240 (N_10240,N_6732,N_8120);
or U10241 (N_10241,N_8902,N_8343);
xnor U10242 (N_10242,N_7390,N_7262);
or U10243 (N_10243,N_9329,N_9189);
nand U10244 (N_10244,N_9213,N_7729);
and U10245 (N_10245,N_8266,N_9062);
nor U10246 (N_10246,N_9075,N_7887);
nor U10247 (N_10247,N_8218,N_8748);
or U10248 (N_10248,N_9064,N_7263);
and U10249 (N_10249,N_8341,N_7578);
or U10250 (N_10250,N_8202,N_8758);
nor U10251 (N_10251,N_7842,N_8973);
nand U10252 (N_10252,N_6317,N_8165);
nor U10253 (N_10253,N_7512,N_6948);
and U10254 (N_10254,N_9152,N_7447);
or U10255 (N_10255,N_8759,N_7367);
and U10256 (N_10256,N_7873,N_7346);
and U10257 (N_10257,N_6970,N_6459);
nand U10258 (N_10258,N_8199,N_9366);
nand U10259 (N_10259,N_6462,N_6480);
nor U10260 (N_10260,N_6897,N_7922);
nor U10261 (N_10261,N_7958,N_8365);
and U10262 (N_10262,N_6426,N_7495);
and U10263 (N_10263,N_7407,N_7234);
and U10264 (N_10264,N_7317,N_8667);
nand U10265 (N_10265,N_7040,N_7759);
and U10266 (N_10266,N_8754,N_8182);
or U10267 (N_10267,N_7531,N_8359);
nor U10268 (N_10268,N_8302,N_7550);
xor U10269 (N_10269,N_9272,N_7071);
or U10270 (N_10270,N_8166,N_7532);
and U10271 (N_10271,N_8533,N_8542);
and U10272 (N_10272,N_7746,N_9180);
nor U10273 (N_10273,N_8635,N_8862);
nor U10274 (N_10274,N_7949,N_8052);
nor U10275 (N_10275,N_8244,N_8017);
nor U10276 (N_10276,N_8556,N_9198);
nand U10277 (N_10277,N_6569,N_7674);
or U10278 (N_10278,N_9305,N_8692);
and U10279 (N_10279,N_8808,N_9264);
nand U10280 (N_10280,N_7051,N_6291);
and U10281 (N_10281,N_7766,N_9063);
and U10282 (N_10282,N_9274,N_8398);
or U10283 (N_10283,N_9175,N_6484);
nor U10284 (N_10284,N_7301,N_6778);
nor U10285 (N_10285,N_7859,N_7975);
or U10286 (N_10286,N_6373,N_8377);
and U10287 (N_10287,N_8762,N_6729);
or U10288 (N_10288,N_6841,N_7731);
xnor U10289 (N_10289,N_6867,N_8241);
or U10290 (N_10290,N_6761,N_7167);
nand U10291 (N_10291,N_7411,N_9229);
xnor U10292 (N_10292,N_8252,N_8818);
nor U10293 (N_10293,N_7231,N_8371);
or U10294 (N_10294,N_6924,N_8020);
or U10295 (N_10295,N_7037,N_8728);
nor U10296 (N_10296,N_8854,N_6386);
nor U10297 (N_10297,N_8509,N_7341);
nand U10298 (N_10298,N_7970,N_8535);
nand U10299 (N_10299,N_6914,N_7596);
nor U10300 (N_10300,N_6861,N_6284);
or U10301 (N_10301,N_7611,N_8374);
or U10302 (N_10302,N_9318,N_8347);
nor U10303 (N_10303,N_7549,N_8169);
nand U10304 (N_10304,N_6252,N_8340);
or U10305 (N_10305,N_6573,N_7395);
or U10306 (N_10306,N_8305,N_6468);
nand U10307 (N_10307,N_8206,N_7405);
nand U10308 (N_10308,N_6344,N_7653);
and U10309 (N_10309,N_7116,N_6780);
or U10310 (N_10310,N_8503,N_7362);
nand U10311 (N_10311,N_8971,N_8525);
and U10312 (N_10312,N_7235,N_6334);
nand U10313 (N_10313,N_7589,N_6465);
xor U10314 (N_10314,N_6626,N_8008);
and U10315 (N_10315,N_6918,N_8953);
nand U10316 (N_10316,N_7499,N_6762);
nand U10317 (N_10317,N_6604,N_8853);
nand U10318 (N_10318,N_8538,N_6295);
nand U10319 (N_10319,N_7448,N_8518);
and U10320 (N_10320,N_6723,N_7375);
and U10321 (N_10321,N_8379,N_7615);
nand U10322 (N_10322,N_8011,N_9007);
nor U10323 (N_10323,N_6585,N_7086);
and U10324 (N_10324,N_7435,N_8647);
nor U10325 (N_10325,N_6874,N_8726);
nand U10326 (N_10326,N_8908,N_7409);
and U10327 (N_10327,N_7189,N_8760);
and U10328 (N_10328,N_6846,N_6639);
xor U10329 (N_10329,N_9110,N_8161);
nor U10330 (N_10330,N_8761,N_7191);
nor U10331 (N_10331,N_8517,N_9055);
or U10332 (N_10332,N_6590,N_8480);
nor U10333 (N_10333,N_8135,N_6448);
nand U10334 (N_10334,N_6370,N_6602);
xnor U10335 (N_10335,N_7297,N_8414);
nor U10336 (N_10336,N_7721,N_8402);
and U10337 (N_10337,N_7722,N_6659);
nor U10338 (N_10338,N_9321,N_8814);
nand U10339 (N_10339,N_7710,N_6910);
xnor U10340 (N_10340,N_7430,N_9184);
or U10341 (N_10341,N_7668,N_7078);
nor U10342 (N_10342,N_6904,N_6310);
nand U10343 (N_10343,N_6262,N_8915);
nand U10344 (N_10344,N_7623,N_8121);
nand U10345 (N_10345,N_7104,N_7376);
or U10346 (N_10346,N_7905,N_6289);
or U10347 (N_10347,N_7725,N_6643);
or U10348 (N_10348,N_8665,N_7511);
or U10349 (N_10349,N_7345,N_7770);
or U10350 (N_10350,N_7728,N_9137);
xnor U10351 (N_10351,N_8957,N_7806);
and U10352 (N_10352,N_6457,N_8636);
and U10353 (N_10353,N_6288,N_7281);
nor U10354 (N_10354,N_6281,N_7743);
and U10355 (N_10355,N_6335,N_8604);
xor U10356 (N_10356,N_6537,N_8550);
xor U10357 (N_10357,N_7644,N_7963);
and U10358 (N_10358,N_8848,N_6888);
and U10359 (N_10359,N_6858,N_7382);
nor U10360 (N_10360,N_9018,N_9061);
nand U10361 (N_10361,N_7516,N_6558);
or U10362 (N_10362,N_8370,N_7762);
and U10363 (N_10363,N_8794,N_6856);
nor U10364 (N_10364,N_7634,N_6491);
and U10365 (N_10365,N_7541,N_7003);
and U10366 (N_10366,N_8788,N_7306);
and U10367 (N_10367,N_9160,N_7145);
nor U10368 (N_10368,N_7436,N_6944);
or U10369 (N_10369,N_9220,N_8586);
or U10370 (N_10370,N_8112,N_7680);
nor U10371 (N_10371,N_8695,N_8996);
xnor U10372 (N_10372,N_8143,N_6406);
nand U10373 (N_10373,N_7476,N_9324);
nand U10374 (N_10374,N_6967,N_8073);
or U10375 (N_10375,N_8755,N_7489);
or U10376 (N_10376,N_6398,N_9139);
nand U10377 (N_10377,N_6660,N_6666);
nor U10378 (N_10378,N_8851,N_6367);
nand U10379 (N_10379,N_8375,N_8742);
xnor U10380 (N_10380,N_7277,N_6410);
xor U10381 (N_10381,N_7750,N_7564);
or U10382 (N_10382,N_8455,N_6560);
and U10383 (N_10383,N_7273,N_6436);
or U10384 (N_10384,N_9261,N_7433);
xnor U10385 (N_10385,N_8633,N_7845);
and U10386 (N_10386,N_8568,N_7947);
nand U10387 (N_10387,N_8792,N_8733);
or U10388 (N_10388,N_9186,N_7748);
and U10389 (N_10389,N_6521,N_9088);
and U10390 (N_10390,N_9135,N_8472);
or U10391 (N_10391,N_8549,N_8693);
nand U10392 (N_10392,N_7713,N_8079);
or U10393 (N_10393,N_9291,N_7582);
nor U10394 (N_10394,N_7013,N_8250);
nand U10395 (N_10395,N_6775,N_6358);
nor U10396 (N_10396,N_7068,N_8443);
and U10397 (N_10397,N_8360,N_7329);
nand U10398 (N_10398,N_8948,N_8799);
and U10399 (N_10399,N_7450,N_6586);
or U10400 (N_10400,N_7188,N_8630);
nand U10401 (N_10401,N_8363,N_9143);
xnor U10402 (N_10402,N_8140,N_6748);
nor U10403 (N_10403,N_6653,N_8712);
nor U10404 (N_10404,N_6685,N_7216);
and U10405 (N_10405,N_8914,N_6443);
nand U10406 (N_10406,N_7613,N_7592);
xnor U10407 (N_10407,N_8824,N_6434);
nor U10408 (N_10408,N_7901,N_6951);
or U10409 (N_10409,N_8526,N_8976);
xor U10410 (N_10410,N_8382,N_9171);
nor U10411 (N_10411,N_8081,N_9046);
nand U10412 (N_10412,N_7148,N_6425);
or U10413 (N_10413,N_8022,N_9315);
nand U10414 (N_10414,N_9208,N_6719);
and U10415 (N_10415,N_6580,N_8435);
or U10416 (N_10416,N_8887,N_7251);
nor U10417 (N_10417,N_9052,N_7606);
or U10418 (N_10418,N_7840,N_7141);
or U10419 (N_10419,N_6956,N_8177);
nand U10420 (N_10420,N_6562,N_8486);
or U10421 (N_10421,N_6663,N_8352);
or U10422 (N_10422,N_6321,N_8710);
or U10423 (N_10423,N_6965,N_9307);
nor U10424 (N_10424,N_9353,N_6716);
nand U10425 (N_10425,N_6739,N_6423);
nand U10426 (N_10426,N_9123,N_8845);
nand U10427 (N_10427,N_9276,N_6301);
or U10428 (N_10428,N_8104,N_7818);
nor U10429 (N_10429,N_7105,N_8131);
xor U10430 (N_10430,N_7839,N_8393);
or U10431 (N_10431,N_8551,N_6565);
and U10432 (N_10432,N_8051,N_8602);
nand U10433 (N_10433,N_8256,N_8944);
or U10434 (N_10434,N_8514,N_7520);
nand U10435 (N_10435,N_7284,N_8460);
or U10436 (N_10436,N_8734,N_9038);
nand U10437 (N_10437,N_8554,N_7028);
and U10438 (N_10438,N_8613,N_9117);
and U10439 (N_10439,N_6575,N_6931);
nor U10440 (N_10440,N_7416,N_6356);
nand U10441 (N_10441,N_8290,N_8784);
or U10442 (N_10442,N_7854,N_6267);
and U10443 (N_10443,N_9326,N_7974);
xor U10444 (N_10444,N_8776,N_8988);
nor U10445 (N_10445,N_7961,N_7026);
or U10446 (N_10446,N_8150,N_6390);
nor U10447 (N_10447,N_8319,N_7391);
nand U10448 (N_10448,N_6539,N_6273);
and U10449 (N_10449,N_9227,N_6875);
and U10450 (N_10450,N_7999,N_7336);
nand U10451 (N_10451,N_7069,N_9177);
or U10452 (N_10452,N_7125,N_7898);
nand U10453 (N_10453,N_8366,N_8717);
nand U10454 (N_10454,N_8867,N_7186);
nand U10455 (N_10455,N_8384,N_6798);
nor U10456 (N_10456,N_8462,N_8949);
nor U10457 (N_10457,N_6961,N_7632);
and U10458 (N_10458,N_8569,N_7214);
nor U10459 (N_10459,N_6801,N_7921);
nor U10460 (N_10460,N_8660,N_6439);
or U10461 (N_10461,N_6957,N_7360);
or U10462 (N_10462,N_9280,N_6634);
nand U10463 (N_10463,N_8450,N_7438);
nor U10464 (N_10464,N_8044,N_8732);
or U10465 (N_10465,N_7664,N_8071);
nor U10466 (N_10466,N_7206,N_8345);
and U10467 (N_10467,N_7777,N_6412);
nor U10468 (N_10468,N_8573,N_7413);
nor U10469 (N_10469,N_6923,N_9030);
nor U10470 (N_10470,N_7291,N_7027);
nor U10471 (N_10471,N_7723,N_7158);
xor U10472 (N_10472,N_9192,N_8113);
nand U10473 (N_10473,N_6290,N_7820);
nand U10474 (N_10474,N_7857,N_6432);
or U10475 (N_10475,N_7115,N_7976);
nand U10476 (N_10476,N_7771,N_8495);
xnor U10477 (N_10477,N_7884,N_7635);
nand U10478 (N_10478,N_7010,N_8955);
nor U10479 (N_10479,N_8819,N_7598);
nand U10480 (N_10480,N_8019,N_7254);
nand U10481 (N_10481,N_8175,N_6717);
nor U10482 (N_10482,N_7195,N_8101);
or U10483 (N_10483,N_8400,N_8736);
xor U10484 (N_10484,N_8888,N_7779);
nand U10485 (N_10485,N_7055,N_6556);
nand U10486 (N_10486,N_6259,N_8584);
nand U10487 (N_10487,N_8268,N_6442);
nor U10488 (N_10488,N_8648,N_7074);
and U10489 (N_10489,N_8997,N_8596);
or U10490 (N_10490,N_6454,N_8321);
or U10491 (N_10491,N_6430,N_7583);
nor U10492 (N_10492,N_6601,N_6528);
or U10493 (N_10493,N_8642,N_7415);
or U10494 (N_10494,N_7891,N_6385);
nand U10495 (N_10495,N_7180,N_6545);
xor U10496 (N_10496,N_8578,N_8484);
or U10497 (N_10497,N_6378,N_7529);
and U10498 (N_10498,N_8048,N_6534);
xnor U10499 (N_10499,N_6445,N_8012);
xnor U10500 (N_10500,N_6348,N_9091);
nand U10501 (N_10501,N_9356,N_6896);
and U10502 (N_10502,N_7171,N_8906);
and U10503 (N_10503,N_9014,N_7997);
or U10504 (N_10504,N_7420,N_8610);
or U10505 (N_10505,N_6903,N_7481);
nand U10506 (N_10506,N_7366,N_9288);
or U10507 (N_10507,N_6350,N_6278);
xor U10508 (N_10508,N_8986,N_7778);
or U10509 (N_10509,N_8650,N_8559);
and U10510 (N_10510,N_8224,N_6921);
xnor U10511 (N_10511,N_7378,N_8032);
or U10512 (N_10512,N_8764,N_8139);
nand U10513 (N_10513,N_9001,N_8053);
xnor U10514 (N_10514,N_7082,N_6988);
or U10515 (N_10515,N_7864,N_7085);
or U10516 (N_10516,N_7562,N_6891);
and U10517 (N_10517,N_7290,N_7551);
nor U10518 (N_10518,N_6460,N_6687);
nor U10519 (N_10519,N_8070,N_8428);
xor U10520 (N_10520,N_8632,N_7737);
nand U10521 (N_10521,N_8930,N_7966);
or U10522 (N_10522,N_8497,N_8306);
nor U10523 (N_10523,N_9136,N_7980);
and U10524 (N_10524,N_6343,N_6409);
or U10525 (N_10525,N_8091,N_7385);
xnor U10526 (N_10526,N_8158,N_6868);
or U10527 (N_10527,N_6250,N_6336);
xnor U10528 (N_10528,N_6688,N_6955);
and U10529 (N_10529,N_7471,N_8852);
nand U10530 (N_10530,N_7248,N_9158);
nand U10531 (N_10531,N_7526,N_8501);
nor U10532 (N_10532,N_7768,N_7939);
or U10533 (N_10533,N_8797,N_9147);
and U10534 (N_10534,N_8390,N_7498);
and U10535 (N_10535,N_8405,N_7265);
xor U10536 (N_10536,N_6427,N_8279);
nor U10537 (N_10537,N_8966,N_6953);
and U10538 (N_10538,N_7323,N_9083);
nand U10539 (N_10539,N_8822,N_9107);
nor U10540 (N_10540,N_7016,N_6536);
and U10541 (N_10541,N_8899,N_7288);
nand U10542 (N_10542,N_8500,N_7904);
and U10543 (N_10543,N_6981,N_8144);
or U10544 (N_10544,N_8844,N_8054);
and U10545 (N_10545,N_6885,N_8316);
or U10546 (N_10546,N_7187,N_7638);
nor U10547 (N_10547,N_8265,N_6791);
or U10548 (N_10548,N_6866,N_8691);
or U10549 (N_10549,N_6946,N_9126);
xor U10550 (N_10550,N_6421,N_6470);
xor U10551 (N_10551,N_6668,N_6870);
nor U10552 (N_10552,N_9092,N_8866);
or U10553 (N_10553,N_7951,N_8361);
or U10554 (N_10554,N_8577,N_8825);
or U10555 (N_10555,N_8581,N_8880);
nor U10556 (N_10556,N_6809,N_6416);
nand U10557 (N_10557,N_9027,N_6789);
or U10558 (N_10558,N_8770,N_6641);
or U10559 (N_10559,N_6754,N_8062);
or U10560 (N_10560,N_8264,N_9299);
nand U10561 (N_10561,N_6388,N_9357);
and U10562 (N_10562,N_6618,N_7827);
or U10563 (N_10563,N_8220,N_6850);
or U10564 (N_10564,N_7834,N_6930);
or U10565 (N_10565,N_7110,N_6260);
or U10566 (N_10566,N_6781,N_8002);
nor U10567 (N_10567,N_9306,N_7089);
or U10568 (N_10568,N_6782,N_6349);
nor U10569 (N_10569,N_7131,N_6346);
and U10570 (N_10570,N_8148,N_8624);
nor U10571 (N_10571,N_6722,N_8466);
and U10572 (N_10572,N_8058,N_8187);
nor U10573 (N_10573,N_8628,N_8487);
nand U10574 (N_10574,N_6352,N_9282);
and U10575 (N_10575,N_8226,N_8653);
nand U10576 (N_10576,N_6593,N_7011);
and U10577 (N_10577,N_7900,N_6691);
or U10578 (N_10578,N_6971,N_7604);
and U10579 (N_10579,N_7618,N_6817);
nor U10580 (N_10580,N_7614,N_8744);
or U10581 (N_10581,N_7663,N_8338);
and U10582 (N_10582,N_9216,N_7260);
nand U10583 (N_10583,N_8541,N_6907);
nor U10584 (N_10584,N_8951,N_8827);
or U10585 (N_10585,N_6509,N_8753);
nand U10586 (N_10586,N_8231,N_9331);
and U10587 (N_10587,N_6737,N_7109);
and U10588 (N_10588,N_7560,N_6251);
or U10589 (N_10589,N_8980,N_7142);
and U10590 (N_10590,N_8194,N_6316);
nand U10591 (N_10591,N_8531,N_7012);
or U10592 (N_10592,N_9273,N_6823);
nor U10593 (N_10593,N_8037,N_8230);
nor U10594 (N_10594,N_9074,N_7910);
or U10595 (N_10595,N_8911,N_8397);
xor U10596 (N_10596,N_7720,N_6374);
nand U10597 (N_10597,N_8701,N_8870);
nor U10598 (N_10598,N_7800,N_8388);
and U10599 (N_10599,N_6932,N_6713);
or U10600 (N_10600,N_6458,N_8167);
or U10601 (N_10601,N_8939,N_8330);
and U10602 (N_10602,N_8775,N_7222);
xnor U10603 (N_10603,N_7309,N_8005);
or U10604 (N_10604,N_6314,N_8510);
nand U10605 (N_10605,N_9196,N_6380);
xnor U10606 (N_10606,N_8018,N_6654);
nand U10607 (N_10607,N_7434,N_7633);
and U10608 (N_10608,N_6557,N_7399);
nor U10609 (N_10609,N_8713,N_8623);
nor U10610 (N_10610,N_6647,N_7767);
nor U10611 (N_10611,N_8960,N_7691);
or U10612 (N_10612,N_6382,N_6803);
nor U10613 (N_10613,N_6527,N_8035);
nand U10614 (N_10614,N_8332,N_8875);
and U10615 (N_10615,N_8631,N_7136);
and U10616 (N_10616,N_7138,N_8918);
nor U10617 (N_10617,N_7500,N_8752);
nor U10618 (N_10618,N_6400,N_8749);
nor U10619 (N_10619,N_7525,N_8743);
nand U10620 (N_10620,N_8159,N_8922);
nor U10621 (N_10621,N_7419,N_8207);
or U10622 (N_10622,N_8894,N_6549);
and U10623 (N_10623,N_7846,N_9340);
nand U10624 (N_10624,N_7863,N_8410);
or U10625 (N_10625,N_7453,N_7620);
nand U10626 (N_10626,N_8817,N_7079);
and U10627 (N_10627,N_7860,N_6744);
and U10628 (N_10628,N_9037,N_6614);
or U10629 (N_10629,N_9179,N_6766);
xnor U10630 (N_10630,N_6714,N_6550);
and U10631 (N_10631,N_7736,N_6588);
nand U10632 (N_10632,N_7268,N_7601);
nor U10633 (N_10633,N_9349,N_6422);
xor U10634 (N_10634,N_6319,N_6543);
xnor U10635 (N_10635,N_9295,N_6297);
xor U10636 (N_10636,N_9151,N_6960);
xor U10637 (N_10637,N_7410,N_8304);
nor U10638 (N_10638,N_7334,N_8999);
xor U10639 (N_10639,N_7194,N_9047);
nor U10640 (N_10640,N_7124,N_6642);
nand U10641 (N_10641,N_6494,N_6347);
nand U10642 (N_10642,N_7002,N_8834);
nor U10643 (N_10643,N_9209,N_7274);
nor U10644 (N_10644,N_6389,N_6263);
nor U10645 (N_10645,N_9067,N_8294);
and U10646 (N_10646,N_8301,N_7826);
nor U10647 (N_10647,N_8823,N_8729);
xor U10648 (N_10648,N_6890,N_6258);
or U10649 (N_10649,N_6452,N_8787);
nand U10650 (N_10650,N_6633,N_6309);
nand U10651 (N_10651,N_7872,N_7754);
or U10652 (N_10652,N_7242,N_7926);
nand U10653 (N_10653,N_8439,N_8962);
nand U10654 (N_10654,N_8034,N_8746);
xor U10655 (N_10655,N_6507,N_6446);
xnor U10656 (N_10656,N_8622,N_6504);
and U10657 (N_10657,N_8136,N_8522);
or U10658 (N_10658,N_8696,N_8267);
nor U10659 (N_10659,N_7097,N_7279);
nor U10660 (N_10660,N_7943,N_8806);
nor U10661 (N_10661,N_7908,N_8331);
xor U10662 (N_10662,N_6511,N_8720);
nor U10663 (N_10663,N_9015,N_9004);
or U10664 (N_10664,N_8248,N_8686);
and U10665 (N_10665,N_7444,N_9125);
and U10666 (N_10666,N_8989,N_8191);
nand U10667 (N_10667,N_6736,N_8040);
nand U10668 (N_10668,N_9191,N_7257);
nand U10669 (N_10669,N_7572,N_8926);
nor U10670 (N_10670,N_7493,N_6972);
or U10671 (N_10671,N_7749,N_8929);
and U10672 (N_10672,N_7646,N_8221);
and U10673 (N_10673,N_8281,N_6695);
nor U10674 (N_10674,N_8204,N_6315);
and U10675 (N_10675,N_7371,N_8431);
and U10676 (N_10676,N_8449,N_8657);
and U10677 (N_10677,N_6399,N_9195);
nand U10678 (N_10678,N_8162,N_6417);
and U10679 (N_10679,N_8543,N_9202);
and U10680 (N_10680,N_6282,N_9127);
nand U10681 (N_10681,N_6311,N_7032);
nand U10682 (N_10682,N_8406,N_9026);
nor U10683 (N_10683,N_9013,N_8090);
and U10684 (N_10684,N_7209,N_6544);
and U10685 (N_10685,N_8821,N_6645);
xnor U10686 (N_10686,N_8210,N_7127);
or U10687 (N_10687,N_6393,N_6843);
nand U10688 (N_10688,N_6756,N_8088);
nand U10689 (N_10689,N_7282,N_6765);
nand U10690 (N_10690,N_7727,N_8750);
nand U10691 (N_10691,N_7769,N_7649);
nand U10692 (N_10692,N_7920,N_6274);
or U10693 (N_10693,N_7579,N_8217);
nand U10694 (N_10694,N_6844,N_7678);
and U10695 (N_10695,N_7349,N_9041);
nand U10696 (N_10696,N_8963,N_8634);
nand U10697 (N_10697,N_8275,N_8676);
nand U10698 (N_10698,N_8767,N_7266);
or U10699 (N_10699,N_7475,N_7302);
nor U10700 (N_10700,N_8492,N_8952);
xor U10701 (N_10701,N_8936,N_7462);
xnor U10702 (N_10702,N_7049,N_7387);
and U10703 (N_10703,N_8444,N_7267);
or U10704 (N_10704,N_6613,N_8873);
nor U10705 (N_10705,N_7066,N_8432);
nand U10706 (N_10706,N_6991,N_6913);
or U10707 (N_10707,N_7521,N_8528);
xnor U10708 (N_10708,N_8036,N_7985);
nand U10709 (N_10709,N_6656,N_7229);
nand U10710 (N_10710,N_7293,N_9325);
nor U10711 (N_10711,N_9000,N_7076);
and U10712 (N_10712,N_8409,N_8446);
and U10713 (N_10713,N_6797,N_7092);
and U10714 (N_10714,N_6863,N_6355);
nor U10715 (N_10715,N_6551,N_8023);
and U10716 (N_10716,N_8452,N_6702);
nand U10717 (N_10717,N_7687,N_8801);
nand U10718 (N_10718,N_7763,N_6790);
or U10719 (N_10719,N_7534,N_6880);
nand U10720 (N_10720,N_7151,N_8045);
and U10721 (N_10721,N_7213,N_6786);
nand U10722 (N_10722,N_7287,N_9259);
nor U10723 (N_10723,N_6612,N_6384);
or U10724 (N_10724,N_7548,N_8679);
nor U10725 (N_10725,N_8108,N_7176);
nor U10726 (N_10726,N_9293,N_8430);
nand U10727 (N_10727,N_9211,N_6265);
and U10728 (N_10728,N_7034,N_7935);
nand U10729 (N_10729,N_7522,N_6898);
and U10730 (N_10730,N_7081,N_6375);
and U10731 (N_10731,N_7962,N_8213);
xnor U10732 (N_10732,N_7686,N_9150);
nand U10733 (N_10733,N_8078,N_7374);
xor U10734 (N_10734,N_7902,N_6622);
nor U10735 (N_10735,N_7111,N_8454);
nor U10736 (N_10736,N_7286,N_9205);
or U10737 (N_10737,N_8298,N_8262);
and U10738 (N_10738,N_8436,N_7523);
xnor U10739 (N_10739,N_6333,N_9368);
xnor U10740 (N_10740,N_8683,N_8850);
and U10741 (N_10741,N_6594,N_8597);
xnor U10742 (N_10742,N_6785,N_6776);
and U10743 (N_10743,N_8663,N_8180);
nand U10744 (N_10744,N_7067,N_8291);
or U10745 (N_10745,N_6387,N_7624);
or U10746 (N_10746,N_7593,N_7852);
nand U10747 (N_10747,N_8009,N_7308);
and U10748 (N_10748,N_7885,N_6912);
nand U10749 (N_10749,N_6268,N_8130);
nor U10750 (N_10750,N_8791,N_8730);
nand U10751 (N_10751,N_7496,N_9235);
xnor U10752 (N_10752,N_7684,N_8245);
nor U10753 (N_10753,N_7654,N_6579);
nand U10754 (N_10754,N_8282,N_8277);
or U10755 (N_10755,N_7501,N_7155);
and U10756 (N_10756,N_8782,N_6636);
and U10757 (N_10757,N_8064,N_9024);
xor U10758 (N_10758,N_7808,N_6734);
and U10759 (N_10759,N_6648,N_8763);
and U10760 (N_10760,N_8423,N_8468);
and U10761 (N_10761,N_6276,N_9168);
or U10762 (N_10762,N_7236,N_7258);
and U10763 (N_10763,N_8456,N_6934);
nor U10764 (N_10764,N_6840,N_8502);
xnor U10765 (N_10765,N_9157,N_8174);
or U10766 (N_10766,N_8802,N_7244);
or U10767 (N_10767,N_7429,N_8969);
or U10768 (N_10768,N_6397,N_8292);
nand U10769 (N_10769,N_6796,N_8335);
or U10770 (N_10770,N_7041,N_7952);
nor U10771 (N_10771,N_8689,N_8721);
or U10772 (N_10772,N_7594,N_7948);
and U10773 (N_10773,N_8066,N_6750);
nand U10774 (N_10774,N_8923,N_6683);
and U10775 (N_10775,N_8987,N_8442);
xnor U10776 (N_10776,N_7215,N_8067);
and U10777 (N_10777,N_6824,N_9078);
and U10778 (N_10778,N_6359,N_7506);
or U10779 (N_10779,N_8625,N_7940);
xor U10780 (N_10780,N_7065,N_7933);
nand U10781 (N_10781,N_9071,N_7911);
nand U10782 (N_10782,N_8965,N_7740);
or U10783 (N_10783,N_9256,N_8014);
or U10784 (N_10784,N_6779,N_6606);
nand U10785 (N_10785,N_8601,N_8580);
nand U10786 (N_10786,N_8324,N_7108);
nor U10787 (N_10787,N_9275,N_8453);
or U10788 (N_10788,N_9335,N_6935);
and U10789 (N_10789,N_6381,N_9268);
or U10790 (N_10790,N_8646,N_8209);
or U10791 (N_10791,N_8785,N_8558);
nand U10792 (N_10792,N_8564,N_9025);
nand U10793 (N_10793,N_8089,N_6628);
and U10794 (N_10794,N_9207,N_7064);
xor U10795 (N_10795,N_8105,N_8476);
nand U10796 (N_10796,N_6513,N_7445);
and U10797 (N_10797,N_7440,N_9044);
or U10798 (N_10798,N_7519,N_8357);
xor U10799 (N_10799,N_6518,N_8307);
and U10800 (N_10800,N_7676,N_9369);
nor U10801 (N_10801,N_7627,N_6804);
nor U10802 (N_10802,N_8912,N_6329);
and U10803 (N_10803,N_8837,N_7482);
or U10804 (N_10804,N_9342,N_6541);
nand U10805 (N_10805,N_7925,N_7835);
and U10806 (N_10806,N_6857,N_6377);
nor U10807 (N_10807,N_6664,N_6490);
or U10808 (N_10808,N_8992,N_6326);
or U10809 (N_10809,N_7077,N_6331);
nand U10810 (N_10810,N_6578,N_7848);
nand U10811 (N_10811,N_8145,N_6631);
and U10812 (N_10812,N_7892,N_8273);
nand U10813 (N_10813,N_8342,N_6881);
and U10814 (N_10814,N_8072,N_6264);
xor U10815 (N_10815,N_6408,N_8682);
or U10816 (N_10816,N_6827,N_6819);
and U10817 (N_10817,N_7218,N_7246);
nor U10818 (N_10818,N_8897,N_8308);
or U10819 (N_10819,N_7515,N_8001);
and U10820 (N_10820,N_8612,N_6254);
or U10821 (N_10821,N_8605,N_8216);
and U10822 (N_10822,N_8149,N_6987);
and U10823 (N_10823,N_7172,N_8567);
nor U10824 (N_10824,N_7569,N_8994);
nor U10825 (N_10825,N_7370,N_7807);
nor U10826 (N_10826,N_7544,N_8707);
nand U10827 (N_10827,N_7312,N_8620);
or U10828 (N_10828,N_6611,N_7484);
nand U10829 (N_10829,N_8257,N_7629);
nor U10830 (N_10830,N_9082,N_6332);
and U10831 (N_10831,N_7147,N_7793);
nand U10832 (N_10832,N_9163,N_8274);
nand U10833 (N_10833,N_9248,N_7488);
nand U10834 (N_10834,N_7987,N_8956);
nor U10835 (N_10835,N_8592,N_8030);
nor U10836 (N_10836,N_6619,N_9347);
nand U10837 (N_10837,N_6644,N_6414);
or U10838 (N_10838,N_7035,N_6977);
or U10839 (N_10839,N_6428,N_7938);
and U10840 (N_10840,N_6751,N_7895);
and U10841 (N_10841,N_7600,N_8523);
and U10842 (N_10842,N_8843,N_6322);
or U10843 (N_10843,N_7802,N_7442);
or U10844 (N_10844,N_9017,N_9285);
and U10845 (N_10845,N_8287,N_8364);
nor U10846 (N_10846,N_8422,N_8705);
nand U10847 (N_10847,N_6862,N_8864);
and U10848 (N_10848,N_8240,N_6559);
or U10849 (N_10849,N_8239,N_8618);
nor U10850 (N_10850,N_6364,N_7603);
or U10851 (N_10851,N_6892,N_8288);
and U10852 (N_10852,N_7851,N_8670);
and U10853 (N_10853,N_8346,N_8640);
nand U10854 (N_10854,N_9346,N_6743);
and U10855 (N_10855,N_8033,N_6937);
and U10856 (N_10856,N_7168,N_7788);
nand U10857 (N_10857,N_7847,N_9362);
and U10858 (N_10858,N_6275,N_6941);
nand U10859 (N_10859,N_6392,N_6435);
or U10860 (N_10860,N_8003,N_8874);
nand U10861 (N_10861,N_7330,N_7483);
and U10862 (N_10862,N_6680,N_8593);
and U10863 (N_10863,N_6829,N_8059);
and U10864 (N_10864,N_8563,N_6600);
xor U10865 (N_10865,N_6922,N_7335);
nand U10866 (N_10866,N_8644,N_7841);
nor U10867 (N_10867,N_8399,N_6257);
or U10868 (N_10868,N_8465,N_8941);
nand U10869 (N_10869,N_7423,N_6901);
or U10870 (N_10870,N_9312,N_7021);
xor U10871 (N_10871,N_7775,N_7313);
nor U10872 (N_10872,N_6339,N_8076);
xnor U10873 (N_10873,N_6607,N_7682);
or U10874 (N_10874,N_8938,N_7906);
or U10875 (N_10875,N_9341,N_8831);
nor U10876 (N_10876,N_6828,N_8765);
and U10877 (N_10877,N_7388,N_8093);
and U10878 (N_10878,N_7253,N_8318);
or U10879 (N_10879,N_6692,N_8395);
nor U10880 (N_10880,N_8661,N_6313);
xor U10881 (N_10881,N_6338,N_7557);
or U10882 (N_10882,N_8328,N_9072);
and U10883 (N_10883,N_6929,N_8703);
nand U10884 (N_10884,N_7879,N_7637);
xor U10885 (N_10885,N_9070,N_8200);
or U10886 (N_10886,N_8786,N_9344);
nor U10887 (N_10887,N_9308,N_9254);
xor U10888 (N_10888,N_7226,N_7437);
xor U10889 (N_10889,N_7117,N_8865);
nand U10890 (N_10890,N_8496,N_8284);
and U10891 (N_10891,N_8126,N_7344);
nand U10892 (N_10892,N_7991,N_7143);
xor U10893 (N_10893,N_6959,N_8907);
or U10894 (N_10894,N_8886,N_9359);
or U10895 (N_10895,N_6982,N_7913);
nor U10896 (N_10896,N_9215,N_6947);
or U10897 (N_10897,N_8125,N_8608);
and U10898 (N_10898,N_6320,N_8222);
or U10899 (N_10899,N_7486,N_7798);
nand U10900 (N_10900,N_8327,N_9316);
nor U10901 (N_10901,N_9162,N_6576);
xnor U10902 (N_10902,N_7338,N_8950);
and U10903 (N_10903,N_7456,N_9054);
or U10904 (N_10904,N_7753,N_7492);
xor U10905 (N_10905,N_9246,N_6895);
xnor U10906 (N_10906,N_7348,N_8702);
nor U10907 (N_10907,N_6337,N_7675);
or U10908 (N_10908,N_7463,N_8715);
nand U10909 (N_10909,N_8473,N_8885);
xnor U10910 (N_10910,N_6553,N_6805);
xor U10911 (N_10911,N_8311,N_9262);
nand U10912 (N_10912,N_6838,N_6997);
nor U10913 (N_10913,N_7819,N_6420);
nor U10914 (N_10914,N_8900,N_7018);
and U10915 (N_10915,N_6469,N_6711);
nand U10916 (N_10916,N_6943,N_7992);
nor U10917 (N_10917,N_6285,N_7657);
or U10918 (N_10918,N_8351,N_7844);
and U10919 (N_10919,N_7739,N_8972);
and U10920 (N_10920,N_8841,N_6821);
and U10921 (N_10921,N_8270,N_7546);
or U10922 (N_10922,N_8225,N_7162);
nand U10923 (N_10923,N_9355,N_8243);
nand U10924 (N_10924,N_9113,N_8738);
or U10925 (N_10925,N_7695,N_7373);
nor U10926 (N_10926,N_9239,N_7937);
nand U10927 (N_10927,N_7524,N_6540);
xnor U10928 (N_10928,N_8412,N_6802);
and U10929 (N_10929,N_6538,N_8959);
nor U10930 (N_10930,N_9320,N_7561);
nor U10931 (N_10931,N_7039,N_9087);
nor U10932 (N_10932,N_8544,N_7869);
nand U10933 (N_10933,N_8027,N_8016);
and U10934 (N_10934,N_6570,N_7539);
and U10935 (N_10935,N_6655,N_7402);
or U10936 (N_10936,N_7225,N_6616);
nor U10937 (N_10937,N_9277,N_6256);
and U10938 (N_10938,N_9262,N_8612);
and U10939 (N_10939,N_6287,N_9226);
and U10940 (N_10940,N_8128,N_7152);
nor U10941 (N_10941,N_7006,N_7081);
nor U10942 (N_10942,N_6733,N_7990);
nor U10943 (N_10943,N_7286,N_6971);
and U10944 (N_10944,N_7420,N_7963);
or U10945 (N_10945,N_8785,N_8680);
and U10946 (N_10946,N_9249,N_8918);
nand U10947 (N_10947,N_7721,N_8180);
xor U10948 (N_10948,N_9084,N_8495);
and U10949 (N_10949,N_7014,N_8045);
or U10950 (N_10950,N_9177,N_9195);
nand U10951 (N_10951,N_7178,N_7128);
nand U10952 (N_10952,N_8463,N_7377);
nor U10953 (N_10953,N_8354,N_7818);
nand U10954 (N_10954,N_9032,N_6437);
xnor U10955 (N_10955,N_6900,N_8002);
nand U10956 (N_10956,N_8214,N_8618);
or U10957 (N_10957,N_9345,N_8668);
nand U10958 (N_10958,N_6318,N_8697);
or U10959 (N_10959,N_8028,N_6565);
nand U10960 (N_10960,N_6580,N_6346);
nand U10961 (N_10961,N_7118,N_7525);
xor U10962 (N_10962,N_8776,N_6317);
nor U10963 (N_10963,N_8510,N_7016);
or U10964 (N_10964,N_9117,N_8357);
or U10965 (N_10965,N_6414,N_8515);
xnor U10966 (N_10966,N_8695,N_7467);
or U10967 (N_10967,N_8602,N_8003);
nand U10968 (N_10968,N_8491,N_6995);
and U10969 (N_10969,N_7660,N_8659);
and U10970 (N_10970,N_6879,N_8754);
and U10971 (N_10971,N_7079,N_8106);
or U10972 (N_10972,N_9106,N_6670);
and U10973 (N_10973,N_7444,N_9351);
nand U10974 (N_10974,N_8931,N_7331);
nand U10975 (N_10975,N_7847,N_8660);
or U10976 (N_10976,N_8631,N_7883);
nand U10977 (N_10977,N_9250,N_8811);
nand U10978 (N_10978,N_6608,N_7753);
nor U10979 (N_10979,N_7897,N_9299);
nor U10980 (N_10980,N_8970,N_8119);
or U10981 (N_10981,N_8543,N_9107);
or U10982 (N_10982,N_6799,N_8370);
and U10983 (N_10983,N_8536,N_6618);
nor U10984 (N_10984,N_6363,N_7113);
or U10985 (N_10985,N_7017,N_9066);
and U10986 (N_10986,N_7119,N_8502);
or U10987 (N_10987,N_7080,N_9310);
or U10988 (N_10988,N_7563,N_6429);
nor U10989 (N_10989,N_8466,N_7242);
nand U10990 (N_10990,N_9227,N_7573);
or U10991 (N_10991,N_9136,N_7574);
or U10992 (N_10992,N_6647,N_8687);
nand U10993 (N_10993,N_6573,N_8580);
and U10994 (N_10994,N_7236,N_8478);
or U10995 (N_10995,N_6327,N_6873);
or U10996 (N_10996,N_6720,N_6972);
nor U10997 (N_10997,N_6902,N_7725);
and U10998 (N_10998,N_9022,N_6852);
nand U10999 (N_10999,N_6623,N_7501);
or U11000 (N_11000,N_8026,N_8619);
nand U11001 (N_11001,N_7159,N_9022);
nor U11002 (N_11002,N_7547,N_6519);
or U11003 (N_11003,N_7035,N_7791);
nor U11004 (N_11004,N_8051,N_6896);
or U11005 (N_11005,N_8357,N_7946);
and U11006 (N_11006,N_7652,N_7362);
nand U11007 (N_11007,N_6789,N_8871);
nor U11008 (N_11008,N_6896,N_8883);
nand U11009 (N_11009,N_9275,N_7556);
nor U11010 (N_11010,N_8391,N_6989);
or U11011 (N_11011,N_7680,N_8064);
or U11012 (N_11012,N_6762,N_8689);
or U11013 (N_11013,N_6509,N_6823);
nor U11014 (N_11014,N_6595,N_6903);
xnor U11015 (N_11015,N_7978,N_7968);
nand U11016 (N_11016,N_7886,N_8581);
nand U11017 (N_11017,N_9127,N_9170);
nand U11018 (N_11018,N_8815,N_6363);
or U11019 (N_11019,N_6268,N_7040);
nor U11020 (N_11020,N_8634,N_8215);
nand U11021 (N_11021,N_9247,N_8828);
nor U11022 (N_11022,N_8535,N_6958);
or U11023 (N_11023,N_8884,N_7368);
or U11024 (N_11024,N_6920,N_8931);
xor U11025 (N_11025,N_6635,N_6612);
nor U11026 (N_11026,N_8320,N_8793);
or U11027 (N_11027,N_8637,N_8289);
nor U11028 (N_11028,N_7851,N_8029);
and U11029 (N_11029,N_7309,N_8582);
xnor U11030 (N_11030,N_7636,N_8639);
or U11031 (N_11031,N_7543,N_7097);
xnor U11032 (N_11032,N_7411,N_7770);
or U11033 (N_11033,N_8103,N_8966);
nand U11034 (N_11034,N_6384,N_8306);
or U11035 (N_11035,N_7436,N_6680);
and U11036 (N_11036,N_7981,N_8981);
nor U11037 (N_11037,N_8673,N_6797);
nand U11038 (N_11038,N_7893,N_7404);
xor U11039 (N_11039,N_8490,N_7886);
or U11040 (N_11040,N_6796,N_6463);
nand U11041 (N_11041,N_8043,N_8938);
and U11042 (N_11042,N_6630,N_8303);
nand U11043 (N_11043,N_8048,N_8570);
xnor U11044 (N_11044,N_7100,N_6323);
nand U11045 (N_11045,N_8217,N_6595);
or U11046 (N_11046,N_9363,N_6693);
nor U11047 (N_11047,N_8868,N_8258);
nand U11048 (N_11048,N_6668,N_6497);
and U11049 (N_11049,N_8837,N_6873);
xnor U11050 (N_11050,N_8528,N_8580);
nor U11051 (N_11051,N_9290,N_8190);
or U11052 (N_11052,N_7164,N_8244);
and U11053 (N_11053,N_9343,N_8608);
or U11054 (N_11054,N_7191,N_7964);
and U11055 (N_11055,N_7886,N_6928);
nor U11056 (N_11056,N_9323,N_6494);
xor U11057 (N_11057,N_8512,N_8233);
or U11058 (N_11058,N_8488,N_6335);
or U11059 (N_11059,N_7555,N_6500);
nor U11060 (N_11060,N_8260,N_7966);
and U11061 (N_11061,N_7385,N_9199);
or U11062 (N_11062,N_8703,N_8321);
nor U11063 (N_11063,N_6973,N_6377);
nand U11064 (N_11064,N_8866,N_9373);
or U11065 (N_11065,N_8482,N_9286);
nor U11066 (N_11066,N_6475,N_6762);
nand U11067 (N_11067,N_9283,N_8468);
or U11068 (N_11068,N_8847,N_6273);
and U11069 (N_11069,N_8820,N_8494);
and U11070 (N_11070,N_7694,N_8579);
nand U11071 (N_11071,N_7611,N_6568);
nand U11072 (N_11072,N_7278,N_8184);
nor U11073 (N_11073,N_7639,N_8007);
or U11074 (N_11074,N_7541,N_8330);
or U11075 (N_11075,N_7263,N_6700);
and U11076 (N_11076,N_8678,N_7758);
or U11077 (N_11077,N_7536,N_9342);
or U11078 (N_11078,N_6471,N_9266);
nand U11079 (N_11079,N_8478,N_6400);
and U11080 (N_11080,N_6971,N_8009);
and U11081 (N_11081,N_6696,N_9173);
or U11082 (N_11082,N_6266,N_6846);
and U11083 (N_11083,N_7668,N_7152);
nor U11084 (N_11084,N_9186,N_9308);
nand U11085 (N_11085,N_7459,N_8965);
or U11086 (N_11086,N_8876,N_6253);
and U11087 (N_11087,N_7045,N_6824);
nand U11088 (N_11088,N_6748,N_7367);
and U11089 (N_11089,N_8823,N_6910);
nand U11090 (N_11090,N_8377,N_8931);
or U11091 (N_11091,N_8632,N_8675);
or U11092 (N_11092,N_6851,N_7080);
nand U11093 (N_11093,N_9294,N_8866);
and U11094 (N_11094,N_9029,N_6549);
or U11095 (N_11095,N_6632,N_8167);
xnor U11096 (N_11096,N_8724,N_6963);
nor U11097 (N_11097,N_6984,N_7327);
or U11098 (N_11098,N_6619,N_7587);
nor U11099 (N_11099,N_6780,N_7933);
nand U11100 (N_11100,N_7136,N_6285);
xor U11101 (N_11101,N_9110,N_7748);
nor U11102 (N_11102,N_8698,N_6970);
nand U11103 (N_11103,N_7590,N_7717);
or U11104 (N_11104,N_7751,N_7297);
or U11105 (N_11105,N_6592,N_8799);
and U11106 (N_11106,N_6366,N_7846);
and U11107 (N_11107,N_9064,N_7583);
nor U11108 (N_11108,N_8391,N_7676);
nor U11109 (N_11109,N_7744,N_8481);
nor U11110 (N_11110,N_7137,N_8530);
nand U11111 (N_11111,N_7462,N_6768);
xor U11112 (N_11112,N_8560,N_7827);
nand U11113 (N_11113,N_8411,N_8398);
or U11114 (N_11114,N_7959,N_8463);
or U11115 (N_11115,N_7422,N_7125);
nand U11116 (N_11116,N_8777,N_7430);
or U11117 (N_11117,N_6422,N_7134);
or U11118 (N_11118,N_8314,N_7254);
nand U11119 (N_11119,N_8781,N_9291);
or U11120 (N_11120,N_8900,N_9078);
nand U11121 (N_11121,N_6783,N_8241);
nor U11122 (N_11122,N_7071,N_6737);
nor U11123 (N_11123,N_6889,N_8824);
nor U11124 (N_11124,N_7694,N_8901);
nor U11125 (N_11125,N_8460,N_8808);
nor U11126 (N_11126,N_9116,N_9203);
xnor U11127 (N_11127,N_8968,N_7399);
or U11128 (N_11128,N_6744,N_8826);
and U11129 (N_11129,N_6343,N_7047);
nand U11130 (N_11130,N_7198,N_7134);
and U11131 (N_11131,N_6282,N_9370);
xnor U11132 (N_11132,N_7294,N_9046);
and U11133 (N_11133,N_7854,N_7699);
and U11134 (N_11134,N_6767,N_6822);
and U11135 (N_11135,N_6857,N_9335);
and U11136 (N_11136,N_7984,N_7745);
and U11137 (N_11137,N_6663,N_7524);
xnor U11138 (N_11138,N_9002,N_8715);
and U11139 (N_11139,N_8792,N_7883);
nor U11140 (N_11140,N_9054,N_6460);
and U11141 (N_11141,N_8985,N_8396);
nand U11142 (N_11142,N_7166,N_6368);
or U11143 (N_11143,N_7779,N_9182);
nor U11144 (N_11144,N_9126,N_7513);
nand U11145 (N_11145,N_8942,N_8361);
xor U11146 (N_11146,N_8126,N_7938);
xnor U11147 (N_11147,N_8270,N_6323);
xnor U11148 (N_11148,N_6388,N_9255);
and U11149 (N_11149,N_9141,N_7767);
and U11150 (N_11150,N_8771,N_7414);
and U11151 (N_11151,N_8162,N_6749);
nand U11152 (N_11152,N_8414,N_8812);
or U11153 (N_11153,N_7339,N_7854);
or U11154 (N_11154,N_7105,N_6806);
xor U11155 (N_11155,N_7399,N_7327);
nand U11156 (N_11156,N_8207,N_9312);
or U11157 (N_11157,N_7956,N_6549);
nor U11158 (N_11158,N_9014,N_7692);
or U11159 (N_11159,N_9159,N_8622);
and U11160 (N_11160,N_7738,N_8960);
or U11161 (N_11161,N_7607,N_7560);
nor U11162 (N_11162,N_8441,N_7151);
nand U11163 (N_11163,N_6620,N_7246);
nand U11164 (N_11164,N_7541,N_8395);
and U11165 (N_11165,N_6942,N_9361);
and U11166 (N_11166,N_7155,N_6570);
nand U11167 (N_11167,N_7808,N_7997);
nand U11168 (N_11168,N_9373,N_6368);
nand U11169 (N_11169,N_7815,N_8777);
nand U11170 (N_11170,N_9299,N_7540);
or U11171 (N_11171,N_8749,N_7713);
and U11172 (N_11172,N_8757,N_7052);
or U11173 (N_11173,N_7832,N_7801);
nor U11174 (N_11174,N_8770,N_6592);
nor U11175 (N_11175,N_7636,N_7029);
nor U11176 (N_11176,N_6430,N_6845);
or U11177 (N_11177,N_8031,N_6969);
nor U11178 (N_11178,N_7309,N_8378);
nand U11179 (N_11179,N_7044,N_7741);
nor U11180 (N_11180,N_6489,N_6630);
and U11181 (N_11181,N_9028,N_6456);
and U11182 (N_11182,N_6330,N_6924);
and U11183 (N_11183,N_6877,N_9335);
nand U11184 (N_11184,N_8215,N_6974);
or U11185 (N_11185,N_8120,N_7886);
nand U11186 (N_11186,N_8954,N_8213);
nand U11187 (N_11187,N_7190,N_9369);
nand U11188 (N_11188,N_7943,N_6427);
nor U11189 (N_11189,N_8928,N_7368);
xor U11190 (N_11190,N_7557,N_8839);
nand U11191 (N_11191,N_7469,N_7301);
nand U11192 (N_11192,N_7829,N_8307);
nand U11193 (N_11193,N_7649,N_6536);
or U11194 (N_11194,N_8978,N_6367);
and U11195 (N_11195,N_8078,N_7418);
nor U11196 (N_11196,N_7053,N_8618);
and U11197 (N_11197,N_9082,N_7709);
nand U11198 (N_11198,N_9006,N_7352);
nor U11199 (N_11199,N_9268,N_9092);
nand U11200 (N_11200,N_6479,N_6461);
and U11201 (N_11201,N_7680,N_7340);
and U11202 (N_11202,N_7172,N_6595);
nor U11203 (N_11203,N_9165,N_7011);
nor U11204 (N_11204,N_7785,N_9285);
or U11205 (N_11205,N_6411,N_9355);
or U11206 (N_11206,N_6672,N_6580);
or U11207 (N_11207,N_8337,N_6389);
nor U11208 (N_11208,N_8014,N_6669);
xnor U11209 (N_11209,N_8299,N_6400);
xnor U11210 (N_11210,N_7196,N_6779);
and U11211 (N_11211,N_7419,N_6346);
and U11212 (N_11212,N_8001,N_9108);
nor U11213 (N_11213,N_8284,N_8478);
xor U11214 (N_11214,N_6321,N_7939);
nor U11215 (N_11215,N_8654,N_7146);
and U11216 (N_11216,N_9226,N_6970);
nand U11217 (N_11217,N_8957,N_8938);
and U11218 (N_11218,N_7525,N_7137);
xor U11219 (N_11219,N_7263,N_6553);
nor U11220 (N_11220,N_9166,N_6549);
xnor U11221 (N_11221,N_6349,N_6888);
nand U11222 (N_11222,N_9023,N_6374);
nand U11223 (N_11223,N_7542,N_8420);
and U11224 (N_11224,N_6564,N_7696);
or U11225 (N_11225,N_8038,N_9237);
xor U11226 (N_11226,N_8200,N_8085);
or U11227 (N_11227,N_7981,N_7408);
nand U11228 (N_11228,N_8871,N_8446);
nand U11229 (N_11229,N_8615,N_8203);
nand U11230 (N_11230,N_7402,N_7081);
nor U11231 (N_11231,N_7397,N_7563);
and U11232 (N_11232,N_7587,N_8608);
xor U11233 (N_11233,N_7275,N_7314);
and U11234 (N_11234,N_7698,N_8049);
and U11235 (N_11235,N_7551,N_8982);
or U11236 (N_11236,N_8523,N_8098);
or U11237 (N_11237,N_6743,N_6827);
nor U11238 (N_11238,N_7041,N_9185);
nor U11239 (N_11239,N_7983,N_6463);
or U11240 (N_11240,N_8848,N_6384);
nand U11241 (N_11241,N_9054,N_8073);
nand U11242 (N_11242,N_8437,N_7263);
and U11243 (N_11243,N_7946,N_6314);
xnor U11244 (N_11244,N_7071,N_7711);
or U11245 (N_11245,N_7858,N_8905);
nor U11246 (N_11246,N_9256,N_7469);
or U11247 (N_11247,N_7706,N_9035);
nand U11248 (N_11248,N_9196,N_6930);
nand U11249 (N_11249,N_8156,N_9287);
xor U11250 (N_11250,N_9136,N_6766);
or U11251 (N_11251,N_6405,N_8815);
nor U11252 (N_11252,N_7040,N_8613);
nand U11253 (N_11253,N_7981,N_8831);
or U11254 (N_11254,N_6977,N_8297);
nand U11255 (N_11255,N_8908,N_6518);
and U11256 (N_11256,N_7556,N_7859);
xnor U11257 (N_11257,N_7566,N_9360);
or U11258 (N_11258,N_8979,N_7103);
xnor U11259 (N_11259,N_7588,N_8593);
nor U11260 (N_11260,N_8747,N_6798);
nand U11261 (N_11261,N_7469,N_6724);
or U11262 (N_11262,N_8578,N_8267);
and U11263 (N_11263,N_9181,N_8585);
or U11264 (N_11264,N_7416,N_6721);
xor U11265 (N_11265,N_6344,N_7197);
xnor U11266 (N_11266,N_7343,N_6426);
nand U11267 (N_11267,N_8674,N_7622);
nor U11268 (N_11268,N_8338,N_7647);
or U11269 (N_11269,N_9081,N_6480);
nor U11270 (N_11270,N_8449,N_6707);
nand U11271 (N_11271,N_7685,N_7526);
or U11272 (N_11272,N_6946,N_6809);
or U11273 (N_11273,N_8965,N_9370);
nand U11274 (N_11274,N_8046,N_8435);
nor U11275 (N_11275,N_9357,N_8946);
nand U11276 (N_11276,N_6702,N_8642);
xor U11277 (N_11277,N_8021,N_9316);
xor U11278 (N_11278,N_6768,N_8349);
nor U11279 (N_11279,N_7228,N_8915);
nand U11280 (N_11280,N_7487,N_9039);
and U11281 (N_11281,N_7125,N_6658);
and U11282 (N_11282,N_7353,N_8739);
nand U11283 (N_11283,N_6536,N_8551);
nand U11284 (N_11284,N_6891,N_8260);
or U11285 (N_11285,N_8874,N_7841);
or U11286 (N_11286,N_8830,N_7893);
nand U11287 (N_11287,N_9131,N_8007);
nor U11288 (N_11288,N_8070,N_7406);
xor U11289 (N_11289,N_8160,N_7449);
or U11290 (N_11290,N_8162,N_6579);
nand U11291 (N_11291,N_9273,N_6912);
nand U11292 (N_11292,N_6956,N_8248);
nor U11293 (N_11293,N_8922,N_7654);
xor U11294 (N_11294,N_7060,N_7670);
or U11295 (N_11295,N_9080,N_7981);
nand U11296 (N_11296,N_7380,N_6756);
nand U11297 (N_11297,N_8998,N_7803);
and U11298 (N_11298,N_7921,N_7481);
nand U11299 (N_11299,N_8493,N_9356);
or U11300 (N_11300,N_8561,N_9054);
nor U11301 (N_11301,N_8642,N_7895);
and U11302 (N_11302,N_7816,N_9215);
nor U11303 (N_11303,N_6778,N_6633);
nor U11304 (N_11304,N_7186,N_8603);
and U11305 (N_11305,N_7793,N_7512);
nor U11306 (N_11306,N_6931,N_8963);
or U11307 (N_11307,N_7665,N_8208);
nand U11308 (N_11308,N_8625,N_9290);
and U11309 (N_11309,N_8119,N_8195);
and U11310 (N_11310,N_7187,N_6779);
nor U11311 (N_11311,N_6796,N_8377);
and U11312 (N_11312,N_6421,N_9328);
xor U11313 (N_11313,N_9077,N_8222);
and U11314 (N_11314,N_9006,N_7729);
nor U11315 (N_11315,N_7303,N_6900);
and U11316 (N_11316,N_6976,N_6777);
and U11317 (N_11317,N_6976,N_9330);
and U11318 (N_11318,N_8845,N_8623);
nand U11319 (N_11319,N_8919,N_7921);
and U11320 (N_11320,N_6777,N_8168);
and U11321 (N_11321,N_9035,N_8686);
nand U11322 (N_11322,N_6473,N_7664);
or U11323 (N_11323,N_8732,N_8196);
and U11324 (N_11324,N_7750,N_9367);
nor U11325 (N_11325,N_9179,N_6747);
nor U11326 (N_11326,N_9006,N_7706);
nor U11327 (N_11327,N_8784,N_7547);
and U11328 (N_11328,N_6254,N_8698);
or U11329 (N_11329,N_6467,N_6375);
and U11330 (N_11330,N_8001,N_9164);
xnor U11331 (N_11331,N_8100,N_9013);
nor U11332 (N_11332,N_9085,N_8949);
nor U11333 (N_11333,N_6441,N_6871);
and U11334 (N_11334,N_7500,N_6797);
nor U11335 (N_11335,N_8946,N_7542);
nor U11336 (N_11336,N_7199,N_7009);
nand U11337 (N_11337,N_7206,N_8212);
xnor U11338 (N_11338,N_7278,N_7685);
and U11339 (N_11339,N_7743,N_8322);
and U11340 (N_11340,N_7186,N_9115);
or U11341 (N_11341,N_6939,N_6348);
and U11342 (N_11342,N_7705,N_6702);
and U11343 (N_11343,N_8531,N_8360);
or U11344 (N_11344,N_9307,N_7452);
nor U11345 (N_11345,N_8423,N_6699);
nor U11346 (N_11346,N_7404,N_8420);
nand U11347 (N_11347,N_7899,N_9093);
and U11348 (N_11348,N_7291,N_8237);
or U11349 (N_11349,N_8317,N_7974);
or U11350 (N_11350,N_8203,N_8467);
and U11351 (N_11351,N_7321,N_8973);
or U11352 (N_11352,N_8543,N_6352);
xnor U11353 (N_11353,N_8687,N_6375);
and U11354 (N_11354,N_7522,N_6950);
and U11355 (N_11355,N_7853,N_6400);
nand U11356 (N_11356,N_6881,N_7665);
nor U11357 (N_11357,N_8484,N_7995);
xnor U11358 (N_11358,N_7084,N_8301);
xor U11359 (N_11359,N_8765,N_7936);
or U11360 (N_11360,N_7761,N_9116);
nand U11361 (N_11361,N_8787,N_8529);
and U11362 (N_11362,N_7400,N_8545);
nor U11363 (N_11363,N_6937,N_8437);
or U11364 (N_11364,N_7770,N_7497);
xor U11365 (N_11365,N_7615,N_8698);
xor U11366 (N_11366,N_8260,N_8938);
or U11367 (N_11367,N_6845,N_6271);
nand U11368 (N_11368,N_9204,N_9025);
or U11369 (N_11369,N_7265,N_8617);
nand U11370 (N_11370,N_8447,N_8245);
nor U11371 (N_11371,N_7701,N_7865);
nand U11372 (N_11372,N_8962,N_7229);
or U11373 (N_11373,N_6816,N_7514);
xnor U11374 (N_11374,N_7984,N_8660);
nor U11375 (N_11375,N_7044,N_6804);
and U11376 (N_11376,N_7397,N_6403);
nand U11377 (N_11377,N_8157,N_7889);
or U11378 (N_11378,N_9312,N_7336);
nand U11379 (N_11379,N_8749,N_8043);
nand U11380 (N_11380,N_6784,N_8440);
or U11381 (N_11381,N_7712,N_8931);
nand U11382 (N_11382,N_7639,N_9282);
and U11383 (N_11383,N_7011,N_8607);
and U11384 (N_11384,N_6427,N_6769);
and U11385 (N_11385,N_6524,N_8116);
nand U11386 (N_11386,N_7272,N_8081);
nand U11387 (N_11387,N_8513,N_9115);
nor U11388 (N_11388,N_6456,N_6878);
nor U11389 (N_11389,N_8424,N_6689);
and U11390 (N_11390,N_8148,N_8931);
xor U11391 (N_11391,N_7476,N_9058);
nand U11392 (N_11392,N_8947,N_8063);
or U11393 (N_11393,N_7309,N_7544);
or U11394 (N_11394,N_6987,N_8377);
nand U11395 (N_11395,N_7072,N_9033);
or U11396 (N_11396,N_8474,N_7539);
xor U11397 (N_11397,N_9188,N_8169);
nor U11398 (N_11398,N_6736,N_8442);
xnor U11399 (N_11399,N_8113,N_6587);
or U11400 (N_11400,N_7278,N_6471);
nand U11401 (N_11401,N_6842,N_7529);
nand U11402 (N_11402,N_8133,N_7557);
or U11403 (N_11403,N_8378,N_9174);
xnor U11404 (N_11404,N_7122,N_7860);
and U11405 (N_11405,N_7795,N_8275);
xnor U11406 (N_11406,N_7139,N_8569);
and U11407 (N_11407,N_9297,N_8779);
xor U11408 (N_11408,N_8324,N_7339);
and U11409 (N_11409,N_9127,N_6694);
nand U11410 (N_11410,N_7195,N_6727);
or U11411 (N_11411,N_8057,N_8461);
nor U11412 (N_11412,N_8055,N_9208);
nor U11413 (N_11413,N_7519,N_9108);
nand U11414 (N_11414,N_8080,N_8376);
or U11415 (N_11415,N_8699,N_7392);
and U11416 (N_11416,N_6810,N_6693);
nand U11417 (N_11417,N_8617,N_6614);
xor U11418 (N_11418,N_7351,N_6830);
nand U11419 (N_11419,N_7150,N_7732);
and U11420 (N_11420,N_8026,N_6305);
nor U11421 (N_11421,N_8264,N_9219);
nor U11422 (N_11422,N_8609,N_7106);
or U11423 (N_11423,N_7519,N_7854);
or U11424 (N_11424,N_8614,N_8280);
nor U11425 (N_11425,N_8304,N_8881);
nor U11426 (N_11426,N_8578,N_7212);
or U11427 (N_11427,N_6283,N_6439);
and U11428 (N_11428,N_8483,N_7257);
or U11429 (N_11429,N_8001,N_8306);
nor U11430 (N_11430,N_7373,N_6464);
nand U11431 (N_11431,N_8663,N_8985);
nand U11432 (N_11432,N_6735,N_7290);
nand U11433 (N_11433,N_7132,N_8961);
or U11434 (N_11434,N_6772,N_7595);
nor U11435 (N_11435,N_6680,N_8125);
nor U11436 (N_11436,N_8063,N_7096);
nand U11437 (N_11437,N_6448,N_8194);
xnor U11438 (N_11438,N_7775,N_7040);
nand U11439 (N_11439,N_6450,N_7433);
or U11440 (N_11440,N_8928,N_7366);
nor U11441 (N_11441,N_9097,N_8065);
nor U11442 (N_11442,N_7839,N_7286);
nand U11443 (N_11443,N_8450,N_8362);
nor U11444 (N_11444,N_8012,N_7705);
and U11445 (N_11445,N_7446,N_8250);
or U11446 (N_11446,N_9004,N_7680);
or U11447 (N_11447,N_6361,N_6605);
nand U11448 (N_11448,N_8665,N_8933);
or U11449 (N_11449,N_8060,N_7101);
xor U11450 (N_11450,N_7308,N_7835);
and U11451 (N_11451,N_8225,N_7363);
nand U11452 (N_11452,N_6303,N_8328);
and U11453 (N_11453,N_8432,N_7545);
nor U11454 (N_11454,N_7981,N_7652);
nor U11455 (N_11455,N_7891,N_7950);
nand U11456 (N_11456,N_9095,N_6375);
nor U11457 (N_11457,N_9115,N_8057);
nor U11458 (N_11458,N_8538,N_7464);
and U11459 (N_11459,N_8825,N_7786);
or U11460 (N_11460,N_8041,N_7546);
and U11461 (N_11461,N_6660,N_9270);
and U11462 (N_11462,N_7578,N_6395);
nor U11463 (N_11463,N_7783,N_8771);
or U11464 (N_11464,N_8706,N_7097);
nand U11465 (N_11465,N_8429,N_7356);
and U11466 (N_11466,N_8992,N_7759);
and U11467 (N_11467,N_8270,N_7623);
and U11468 (N_11468,N_7048,N_8555);
xor U11469 (N_11469,N_9145,N_6741);
or U11470 (N_11470,N_9247,N_8783);
nand U11471 (N_11471,N_9311,N_9327);
xor U11472 (N_11472,N_6560,N_8531);
and U11473 (N_11473,N_8967,N_6288);
or U11474 (N_11474,N_7191,N_8440);
nor U11475 (N_11475,N_8839,N_7685);
and U11476 (N_11476,N_6743,N_6549);
and U11477 (N_11477,N_8406,N_8630);
and U11478 (N_11478,N_8133,N_9341);
or U11479 (N_11479,N_7160,N_6440);
xor U11480 (N_11480,N_6564,N_8118);
or U11481 (N_11481,N_8239,N_9000);
nor U11482 (N_11482,N_7699,N_8517);
and U11483 (N_11483,N_6665,N_7137);
nand U11484 (N_11484,N_9047,N_7461);
nand U11485 (N_11485,N_7277,N_8894);
nor U11486 (N_11486,N_8376,N_6434);
nor U11487 (N_11487,N_8729,N_8290);
and U11488 (N_11488,N_6714,N_8256);
and U11489 (N_11489,N_8262,N_8535);
and U11490 (N_11490,N_8568,N_9309);
and U11491 (N_11491,N_7463,N_8883);
xnor U11492 (N_11492,N_6944,N_6760);
nand U11493 (N_11493,N_8302,N_8008);
or U11494 (N_11494,N_6400,N_6519);
xnor U11495 (N_11495,N_7964,N_7893);
nand U11496 (N_11496,N_9197,N_7423);
or U11497 (N_11497,N_9118,N_6598);
nor U11498 (N_11498,N_6352,N_7590);
or U11499 (N_11499,N_7233,N_7073);
or U11500 (N_11500,N_7737,N_8095);
or U11501 (N_11501,N_7964,N_7900);
and U11502 (N_11502,N_8713,N_8871);
and U11503 (N_11503,N_8139,N_7808);
nor U11504 (N_11504,N_6949,N_7215);
nor U11505 (N_11505,N_7989,N_8779);
nor U11506 (N_11506,N_9350,N_9229);
or U11507 (N_11507,N_8657,N_9303);
and U11508 (N_11508,N_6909,N_7037);
and U11509 (N_11509,N_8533,N_8558);
nor U11510 (N_11510,N_8453,N_8116);
or U11511 (N_11511,N_7943,N_8991);
nor U11512 (N_11512,N_6336,N_8737);
and U11513 (N_11513,N_7696,N_7438);
or U11514 (N_11514,N_8258,N_7775);
nand U11515 (N_11515,N_7381,N_6830);
and U11516 (N_11516,N_7337,N_8418);
or U11517 (N_11517,N_8137,N_7206);
nor U11518 (N_11518,N_8640,N_6395);
or U11519 (N_11519,N_7746,N_6809);
nand U11520 (N_11520,N_8904,N_7770);
nand U11521 (N_11521,N_9270,N_8260);
nor U11522 (N_11522,N_8206,N_6493);
and U11523 (N_11523,N_7927,N_6565);
or U11524 (N_11524,N_7946,N_7907);
and U11525 (N_11525,N_6684,N_6634);
nand U11526 (N_11526,N_9137,N_8371);
or U11527 (N_11527,N_6764,N_6362);
nor U11528 (N_11528,N_8428,N_9028);
or U11529 (N_11529,N_7719,N_7880);
nor U11530 (N_11530,N_8980,N_9262);
or U11531 (N_11531,N_8615,N_7314);
and U11532 (N_11532,N_7781,N_6698);
or U11533 (N_11533,N_8341,N_8833);
nand U11534 (N_11534,N_7330,N_8463);
and U11535 (N_11535,N_7060,N_8827);
nand U11536 (N_11536,N_9352,N_7962);
and U11537 (N_11537,N_7041,N_8655);
nand U11538 (N_11538,N_8257,N_6856);
xor U11539 (N_11539,N_7271,N_7421);
and U11540 (N_11540,N_7198,N_7885);
or U11541 (N_11541,N_9075,N_8871);
or U11542 (N_11542,N_6844,N_8218);
nand U11543 (N_11543,N_8411,N_6419);
and U11544 (N_11544,N_7001,N_8985);
or U11545 (N_11545,N_6893,N_6759);
nand U11546 (N_11546,N_6972,N_8610);
or U11547 (N_11547,N_6872,N_6301);
and U11548 (N_11548,N_7605,N_9213);
nor U11549 (N_11549,N_9072,N_7462);
nand U11550 (N_11550,N_7100,N_7782);
xnor U11551 (N_11551,N_7526,N_7128);
and U11552 (N_11552,N_7376,N_7859);
nor U11553 (N_11553,N_8089,N_6672);
nor U11554 (N_11554,N_7060,N_8166);
and U11555 (N_11555,N_6383,N_6520);
and U11556 (N_11556,N_7869,N_8784);
nand U11557 (N_11557,N_7606,N_8286);
and U11558 (N_11558,N_7757,N_7286);
or U11559 (N_11559,N_6415,N_7065);
or U11560 (N_11560,N_6260,N_7339);
or U11561 (N_11561,N_9186,N_8922);
or U11562 (N_11562,N_8691,N_7087);
or U11563 (N_11563,N_7018,N_7721);
and U11564 (N_11564,N_8373,N_7826);
and U11565 (N_11565,N_8727,N_8092);
and U11566 (N_11566,N_6843,N_8248);
and U11567 (N_11567,N_7760,N_9275);
and U11568 (N_11568,N_8142,N_6948);
nor U11569 (N_11569,N_7084,N_8024);
nand U11570 (N_11570,N_7730,N_8130);
and U11571 (N_11571,N_8478,N_7866);
or U11572 (N_11572,N_6309,N_6318);
and U11573 (N_11573,N_6258,N_6278);
and U11574 (N_11574,N_7850,N_9162);
xnor U11575 (N_11575,N_7603,N_7831);
and U11576 (N_11576,N_8291,N_8612);
and U11577 (N_11577,N_8531,N_8323);
and U11578 (N_11578,N_7810,N_7455);
xor U11579 (N_11579,N_7874,N_6778);
or U11580 (N_11580,N_8438,N_8620);
nor U11581 (N_11581,N_6936,N_8392);
nand U11582 (N_11582,N_9042,N_6549);
or U11583 (N_11583,N_8691,N_8904);
nand U11584 (N_11584,N_7689,N_9045);
or U11585 (N_11585,N_8753,N_8026);
nor U11586 (N_11586,N_7565,N_7913);
or U11587 (N_11587,N_6792,N_6272);
and U11588 (N_11588,N_8195,N_8400);
and U11589 (N_11589,N_9284,N_6445);
and U11590 (N_11590,N_6280,N_6587);
nor U11591 (N_11591,N_9265,N_8507);
nand U11592 (N_11592,N_9031,N_6611);
nand U11593 (N_11593,N_6752,N_7105);
nor U11594 (N_11594,N_6661,N_7794);
or U11595 (N_11595,N_8348,N_8887);
nor U11596 (N_11596,N_6409,N_8005);
and U11597 (N_11597,N_8816,N_8965);
nor U11598 (N_11598,N_7023,N_7605);
and U11599 (N_11599,N_6647,N_6549);
or U11600 (N_11600,N_8340,N_8267);
nor U11601 (N_11601,N_8555,N_6651);
nand U11602 (N_11602,N_8811,N_8547);
nand U11603 (N_11603,N_8172,N_7562);
nor U11604 (N_11604,N_7406,N_9094);
and U11605 (N_11605,N_6927,N_6503);
and U11606 (N_11606,N_6604,N_6390);
or U11607 (N_11607,N_8382,N_6557);
xnor U11608 (N_11608,N_8678,N_7424);
nand U11609 (N_11609,N_8948,N_8539);
nor U11610 (N_11610,N_8998,N_7317);
nand U11611 (N_11611,N_7197,N_6279);
nand U11612 (N_11612,N_7637,N_6385);
and U11613 (N_11613,N_7456,N_8277);
nand U11614 (N_11614,N_6596,N_7775);
nand U11615 (N_11615,N_9066,N_6275);
and U11616 (N_11616,N_9041,N_6895);
or U11617 (N_11617,N_7898,N_7677);
xor U11618 (N_11618,N_8924,N_6845);
nor U11619 (N_11619,N_8744,N_9066);
nand U11620 (N_11620,N_8687,N_8588);
nand U11621 (N_11621,N_8537,N_7761);
nor U11622 (N_11622,N_8956,N_7872);
nor U11623 (N_11623,N_9029,N_7039);
nor U11624 (N_11624,N_6932,N_6780);
and U11625 (N_11625,N_7660,N_6668);
and U11626 (N_11626,N_8120,N_9291);
and U11627 (N_11627,N_6760,N_6303);
nor U11628 (N_11628,N_6461,N_6658);
or U11629 (N_11629,N_9289,N_8721);
nor U11630 (N_11630,N_9048,N_7361);
or U11631 (N_11631,N_9170,N_7346);
nor U11632 (N_11632,N_8461,N_8380);
nand U11633 (N_11633,N_9004,N_6737);
or U11634 (N_11634,N_8278,N_6645);
nor U11635 (N_11635,N_8634,N_9373);
nor U11636 (N_11636,N_7559,N_9361);
nor U11637 (N_11637,N_8744,N_6283);
nand U11638 (N_11638,N_7307,N_6621);
and U11639 (N_11639,N_8705,N_7655);
and U11640 (N_11640,N_9306,N_8011);
xnor U11641 (N_11641,N_8172,N_8328);
or U11642 (N_11642,N_8764,N_6772);
and U11643 (N_11643,N_8847,N_8685);
and U11644 (N_11644,N_7937,N_7593);
nor U11645 (N_11645,N_7266,N_8962);
xnor U11646 (N_11646,N_6837,N_6652);
nand U11647 (N_11647,N_6427,N_8679);
or U11648 (N_11648,N_7043,N_8975);
xor U11649 (N_11649,N_7941,N_7276);
and U11650 (N_11650,N_8132,N_6417);
nand U11651 (N_11651,N_6800,N_7297);
and U11652 (N_11652,N_8920,N_7899);
nor U11653 (N_11653,N_6766,N_8532);
nor U11654 (N_11654,N_8991,N_8733);
nand U11655 (N_11655,N_8942,N_6373);
or U11656 (N_11656,N_8231,N_8432);
and U11657 (N_11657,N_7119,N_6578);
nor U11658 (N_11658,N_8722,N_8689);
nor U11659 (N_11659,N_9087,N_8976);
xor U11660 (N_11660,N_9017,N_8814);
nor U11661 (N_11661,N_8137,N_8822);
and U11662 (N_11662,N_6665,N_8972);
nand U11663 (N_11663,N_8543,N_8369);
nor U11664 (N_11664,N_8601,N_8547);
nor U11665 (N_11665,N_8992,N_8040);
nand U11666 (N_11666,N_7857,N_8038);
xnor U11667 (N_11667,N_7676,N_8811);
or U11668 (N_11668,N_6294,N_8684);
or U11669 (N_11669,N_6250,N_6561);
nor U11670 (N_11670,N_7276,N_7690);
nor U11671 (N_11671,N_7524,N_9308);
or U11672 (N_11672,N_6367,N_7716);
nor U11673 (N_11673,N_8910,N_8198);
nor U11674 (N_11674,N_6476,N_7398);
and U11675 (N_11675,N_9353,N_8568);
nor U11676 (N_11676,N_8567,N_8272);
nand U11677 (N_11677,N_8776,N_8230);
nand U11678 (N_11678,N_6954,N_6905);
nor U11679 (N_11679,N_9190,N_7845);
or U11680 (N_11680,N_8053,N_7244);
xor U11681 (N_11681,N_7547,N_7062);
nor U11682 (N_11682,N_6997,N_8296);
nand U11683 (N_11683,N_7766,N_8524);
or U11684 (N_11684,N_8416,N_6880);
xor U11685 (N_11685,N_8428,N_8170);
nand U11686 (N_11686,N_8437,N_7085);
and U11687 (N_11687,N_7214,N_7313);
nor U11688 (N_11688,N_8812,N_7344);
or U11689 (N_11689,N_8270,N_6421);
or U11690 (N_11690,N_7080,N_8268);
or U11691 (N_11691,N_8871,N_7987);
or U11692 (N_11692,N_8139,N_7664);
nand U11693 (N_11693,N_9088,N_6561);
and U11694 (N_11694,N_7414,N_6605);
or U11695 (N_11695,N_6792,N_7164);
nor U11696 (N_11696,N_8418,N_6463);
nand U11697 (N_11697,N_6755,N_7520);
nand U11698 (N_11698,N_9238,N_6294);
nor U11699 (N_11699,N_8484,N_7965);
nand U11700 (N_11700,N_6623,N_6417);
and U11701 (N_11701,N_8984,N_9332);
nand U11702 (N_11702,N_7193,N_8998);
nor U11703 (N_11703,N_6526,N_9281);
xnor U11704 (N_11704,N_6694,N_8536);
and U11705 (N_11705,N_8037,N_8766);
xor U11706 (N_11706,N_6816,N_6541);
xor U11707 (N_11707,N_7020,N_8121);
or U11708 (N_11708,N_7844,N_9321);
or U11709 (N_11709,N_8598,N_6920);
and U11710 (N_11710,N_6376,N_9044);
nand U11711 (N_11711,N_8876,N_9284);
nand U11712 (N_11712,N_6287,N_6318);
nor U11713 (N_11713,N_6734,N_8134);
or U11714 (N_11714,N_9269,N_6559);
nor U11715 (N_11715,N_8902,N_7696);
xnor U11716 (N_11716,N_7954,N_8750);
nor U11717 (N_11717,N_6679,N_6516);
and U11718 (N_11718,N_7471,N_6639);
and U11719 (N_11719,N_7461,N_9087);
or U11720 (N_11720,N_8561,N_7251);
or U11721 (N_11721,N_8104,N_8930);
xnor U11722 (N_11722,N_8753,N_6683);
xnor U11723 (N_11723,N_8099,N_7546);
nand U11724 (N_11724,N_7601,N_8458);
nor U11725 (N_11725,N_7167,N_6924);
nor U11726 (N_11726,N_6321,N_7662);
nor U11727 (N_11727,N_8870,N_6934);
nand U11728 (N_11728,N_7573,N_6789);
nor U11729 (N_11729,N_6906,N_9216);
or U11730 (N_11730,N_9286,N_7081);
and U11731 (N_11731,N_7251,N_6520);
nand U11732 (N_11732,N_7027,N_6455);
or U11733 (N_11733,N_7604,N_6373);
or U11734 (N_11734,N_8212,N_8792);
and U11735 (N_11735,N_6643,N_6392);
and U11736 (N_11736,N_8309,N_8089);
or U11737 (N_11737,N_8035,N_9087);
nor U11738 (N_11738,N_8284,N_6488);
or U11739 (N_11739,N_8279,N_6944);
and U11740 (N_11740,N_7955,N_8798);
xor U11741 (N_11741,N_7066,N_6973);
or U11742 (N_11742,N_8930,N_9289);
nor U11743 (N_11743,N_6651,N_8030);
nor U11744 (N_11744,N_8471,N_7390);
nand U11745 (N_11745,N_8627,N_8507);
and U11746 (N_11746,N_7248,N_9131);
or U11747 (N_11747,N_9333,N_7207);
nand U11748 (N_11748,N_6437,N_6458);
nand U11749 (N_11749,N_7185,N_8497);
and U11750 (N_11750,N_9071,N_8375);
xnor U11751 (N_11751,N_6676,N_8112);
or U11752 (N_11752,N_9369,N_7663);
and U11753 (N_11753,N_7041,N_9017);
nand U11754 (N_11754,N_9146,N_7022);
xnor U11755 (N_11755,N_7134,N_8647);
nand U11756 (N_11756,N_8645,N_6812);
or U11757 (N_11757,N_7934,N_7747);
nor U11758 (N_11758,N_8100,N_8865);
nand U11759 (N_11759,N_9210,N_6823);
nor U11760 (N_11760,N_6513,N_7093);
nor U11761 (N_11761,N_7934,N_8699);
and U11762 (N_11762,N_7848,N_6865);
and U11763 (N_11763,N_8777,N_7239);
and U11764 (N_11764,N_6971,N_8814);
nor U11765 (N_11765,N_7488,N_8967);
nand U11766 (N_11766,N_8543,N_8613);
nand U11767 (N_11767,N_9081,N_8529);
nor U11768 (N_11768,N_8636,N_7509);
nor U11769 (N_11769,N_8589,N_9050);
and U11770 (N_11770,N_7263,N_9245);
nor U11771 (N_11771,N_9292,N_7701);
and U11772 (N_11772,N_7632,N_8761);
or U11773 (N_11773,N_8020,N_9068);
and U11774 (N_11774,N_6422,N_8620);
or U11775 (N_11775,N_7726,N_7111);
nand U11776 (N_11776,N_7369,N_9299);
and U11777 (N_11777,N_9359,N_7871);
nor U11778 (N_11778,N_8914,N_6973);
or U11779 (N_11779,N_8620,N_7652);
nor U11780 (N_11780,N_7204,N_9009);
or U11781 (N_11781,N_9212,N_9250);
nand U11782 (N_11782,N_9107,N_7814);
xor U11783 (N_11783,N_8426,N_6652);
and U11784 (N_11784,N_9118,N_6458);
nand U11785 (N_11785,N_9166,N_7293);
or U11786 (N_11786,N_6802,N_7844);
nor U11787 (N_11787,N_7332,N_7818);
nand U11788 (N_11788,N_8858,N_7347);
and U11789 (N_11789,N_9238,N_8979);
and U11790 (N_11790,N_6438,N_6716);
and U11791 (N_11791,N_8686,N_8482);
and U11792 (N_11792,N_8516,N_6744);
or U11793 (N_11793,N_6932,N_7404);
nor U11794 (N_11794,N_8079,N_6854);
nor U11795 (N_11795,N_6742,N_8638);
and U11796 (N_11796,N_7745,N_6842);
or U11797 (N_11797,N_8892,N_8454);
and U11798 (N_11798,N_6956,N_8159);
and U11799 (N_11799,N_6805,N_8331);
nor U11800 (N_11800,N_8821,N_6747);
or U11801 (N_11801,N_6735,N_9306);
nand U11802 (N_11802,N_9354,N_6615);
nand U11803 (N_11803,N_8799,N_6333);
and U11804 (N_11804,N_6744,N_6509);
or U11805 (N_11805,N_6785,N_8640);
or U11806 (N_11806,N_8435,N_9213);
and U11807 (N_11807,N_8890,N_7943);
and U11808 (N_11808,N_8584,N_8933);
and U11809 (N_11809,N_8885,N_6420);
nand U11810 (N_11810,N_8932,N_9293);
nand U11811 (N_11811,N_7061,N_8293);
nand U11812 (N_11812,N_6902,N_7570);
or U11813 (N_11813,N_7178,N_6411);
nor U11814 (N_11814,N_6365,N_9171);
nand U11815 (N_11815,N_7083,N_6995);
nand U11816 (N_11816,N_8127,N_8740);
nand U11817 (N_11817,N_8531,N_9143);
nor U11818 (N_11818,N_9253,N_9335);
nand U11819 (N_11819,N_8710,N_8833);
nand U11820 (N_11820,N_8809,N_7322);
and U11821 (N_11821,N_8043,N_7379);
xor U11822 (N_11822,N_7561,N_8051);
nand U11823 (N_11823,N_7761,N_6865);
or U11824 (N_11824,N_9023,N_6618);
and U11825 (N_11825,N_9146,N_8912);
nand U11826 (N_11826,N_7231,N_7894);
nand U11827 (N_11827,N_7960,N_9212);
or U11828 (N_11828,N_6658,N_7220);
nand U11829 (N_11829,N_7524,N_7704);
or U11830 (N_11830,N_8447,N_7856);
nand U11831 (N_11831,N_8524,N_9219);
xnor U11832 (N_11832,N_7473,N_9154);
and U11833 (N_11833,N_8360,N_6951);
and U11834 (N_11834,N_7930,N_6483);
and U11835 (N_11835,N_9335,N_9220);
or U11836 (N_11836,N_7263,N_8302);
nor U11837 (N_11837,N_6278,N_7084);
and U11838 (N_11838,N_6857,N_6682);
and U11839 (N_11839,N_7940,N_7283);
nand U11840 (N_11840,N_8643,N_6475);
nor U11841 (N_11841,N_7991,N_6272);
or U11842 (N_11842,N_9289,N_7383);
or U11843 (N_11843,N_9131,N_8244);
nor U11844 (N_11844,N_7601,N_8947);
nor U11845 (N_11845,N_7448,N_8014);
and U11846 (N_11846,N_7188,N_7322);
and U11847 (N_11847,N_8646,N_6832);
xor U11848 (N_11848,N_8495,N_7137);
nand U11849 (N_11849,N_8406,N_8370);
or U11850 (N_11850,N_7198,N_7304);
nand U11851 (N_11851,N_7608,N_7460);
nor U11852 (N_11852,N_7579,N_6816);
nor U11853 (N_11853,N_9335,N_6273);
and U11854 (N_11854,N_8854,N_7870);
nor U11855 (N_11855,N_8331,N_8059);
or U11856 (N_11856,N_6359,N_9189);
nor U11857 (N_11857,N_6609,N_7607);
nor U11858 (N_11858,N_7380,N_8216);
or U11859 (N_11859,N_7292,N_9261);
nand U11860 (N_11860,N_7971,N_7783);
nand U11861 (N_11861,N_7584,N_8870);
and U11862 (N_11862,N_8448,N_8190);
or U11863 (N_11863,N_7758,N_8693);
nand U11864 (N_11864,N_9009,N_6308);
nor U11865 (N_11865,N_7248,N_9243);
nor U11866 (N_11866,N_6294,N_8311);
nand U11867 (N_11867,N_8858,N_6395);
xnor U11868 (N_11868,N_8539,N_6802);
nor U11869 (N_11869,N_7984,N_6539);
nor U11870 (N_11870,N_8362,N_7327);
or U11871 (N_11871,N_9217,N_6916);
nand U11872 (N_11872,N_8887,N_7292);
and U11873 (N_11873,N_8673,N_6613);
nand U11874 (N_11874,N_6666,N_6867);
nor U11875 (N_11875,N_7665,N_8947);
or U11876 (N_11876,N_7855,N_7504);
nand U11877 (N_11877,N_9273,N_9316);
nor U11878 (N_11878,N_8363,N_6876);
nand U11879 (N_11879,N_6297,N_7472);
and U11880 (N_11880,N_7796,N_8736);
nor U11881 (N_11881,N_6289,N_6953);
nand U11882 (N_11882,N_7621,N_7200);
nor U11883 (N_11883,N_9092,N_8553);
nor U11884 (N_11884,N_7487,N_6585);
nand U11885 (N_11885,N_7455,N_7988);
nor U11886 (N_11886,N_6420,N_8926);
or U11887 (N_11887,N_7731,N_8987);
nor U11888 (N_11888,N_7478,N_6443);
nand U11889 (N_11889,N_9300,N_7254);
and U11890 (N_11890,N_8416,N_8534);
and U11891 (N_11891,N_8953,N_8210);
nor U11892 (N_11892,N_6266,N_7191);
and U11893 (N_11893,N_8024,N_7279);
or U11894 (N_11894,N_6853,N_6929);
nor U11895 (N_11895,N_6378,N_6274);
and U11896 (N_11896,N_7788,N_8264);
nor U11897 (N_11897,N_6965,N_7453);
xnor U11898 (N_11898,N_7194,N_7140);
nor U11899 (N_11899,N_8892,N_7031);
or U11900 (N_11900,N_6442,N_7180);
and U11901 (N_11901,N_8546,N_7959);
xnor U11902 (N_11902,N_8651,N_7728);
xnor U11903 (N_11903,N_7048,N_9296);
and U11904 (N_11904,N_7357,N_6588);
or U11905 (N_11905,N_8771,N_7339);
nor U11906 (N_11906,N_7242,N_6840);
xor U11907 (N_11907,N_8983,N_9135);
and U11908 (N_11908,N_7740,N_7188);
nand U11909 (N_11909,N_6389,N_8877);
or U11910 (N_11910,N_6350,N_7783);
and U11911 (N_11911,N_8829,N_6941);
nor U11912 (N_11912,N_9068,N_6375);
or U11913 (N_11913,N_6346,N_8301);
nor U11914 (N_11914,N_8923,N_6797);
or U11915 (N_11915,N_7137,N_9242);
xnor U11916 (N_11916,N_8409,N_7543);
nand U11917 (N_11917,N_6955,N_8317);
xor U11918 (N_11918,N_7584,N_7144);
or U11919 (N_11919,N_7295,N_8280);
nor U11920 (N_11920,N_8907,N_7041);
and U11921 (N_11921,N_8600,N_8536);
nand U11922 (N_11922,N_7103,N_8733);
or U11923 (N_11923,N_6385,N_7714);
nor U11924 (N_11924,N_7076,N_8103);
and U11925 (N_11925,N_7220,N_7847);
nor U11926 (N_11926,N_7242,N_8689);
xor U11927 (N_11927,N_6974,N_7851);
nor U11928 (N_11928,N_8141,N_8258);
and U11929 (N_11929,N_7098,N_8148);
or U11930 (N_11930,N_7616,N_8761);
nand U11931 (N_11931,N_9304,N_6274);
or U11932 (N_11932,N_9115,N_6649);
xor U11933 (N_11933,N_9220,N_7504);
nor U11934 (N_11934,N_8522,N_8215);
nor U11935 (N_11935,N_8491,N_7839);
nand U11936 (N_11936,N_9301,N_7097);
nor U11937 (N_11937,N_9018,N_8002);
or U11938 (N_11938,N_6438,N_7031);
and U11939 (N_11939,N_8053,N_6895);
nand U11940 (N_11940,N_9308,N_7958);
and U11941 (N_11941,N_8207,N_6836);
and U11942 (N_11942,N_8469,N_9328);
or U11943 (N_11943,N_8714,N_7417);
nor U11944 (N_11944,N_9151,N_8573);
nand U11945 (N_11945,N_7230,N_7683);
nand U11946 (N_11946,N_7852,N_8256);
or U11947 (N_11947,N_7756,N_6527);
nand U11948 (N_11948,N_6359,N_7729);
nand U11949 (N_11949,N_6668,N_7166);
nor U11950 (N_11950,N_8506,N_7173);
nand U11951 (N_11951,N_6653,N_9326);
and U11952 (N_11952,N_6981,N_7749);
or U11953 (N_11953,N_8048,N_7296);
nor U11954 (N_11954,N_6856,N_8494);
and U11955 (N_11955,N_6579,N_8959);
nor U11956 (N_11956,N_7556,N_6345);
nor U11957 (N_11957,N_6658,N_6409);
or U11958 (N_11958,N_6469,N_7781);
and U11959 (N_11959,N_6768,N_8557);
nor U11960 (N_11960,N_7663,N_8478);
nor U11961 (N_11961,N_8824,N_7001);
nand U11962 (N_11962,N_9150,N_7862);
or U11963 (N_11963,N_7089,N_8005);
xor U11964 (N_11964,N_7121,N_6566);
nor U11965 (N_11965,N_8832,N_6906);
nor U11966 (N_11966,N_7361,N_7016);
xnor U11967 (N_11967,N_8333,N_9355);
nor U11968 (N_11968,N_7224,N_6657);
and U11969 (N_11969,N_8593,N_7236);
nand U11970 (N_11970,N_7984,N_8922);
nor U11971 (N_11971,N_7873,N_8319);
and U11972 (N_11972,N_8468,N_7355);
nand U11973 (N_11973,N_7547,N_8486);
or U11974 (N_11974,N_6659,N_8860);
xnor U11975 (N_11975,N_6281,N_7039);
and U11976 (N_11976,N_6897,N_9288);
nand U11977 (N_11977,N_8592,N_6715);
or U11978 (N_11978,N_7422,N_7199);
nor U11979 (N_11979,N_6998,N_8178);
nand U11980 (N_11980,N_8463,N_8180);
nand U11981 (N_11981,N_8296,N_7730);
nor U11982 (N_11982,N_8284,N_9222);
and U11983 (N_11983,N_8818,N_7174);
and U11984 (N_11984,N_6615,N_7151);
nor U11985 (N_11985,N_9262,N_7781);
and U11986 (N_11986,N_6643,N_8659);
nand U11987 (N_11987,N_8821,N_9366);
nor U11988 (N_11988,N_9180,N_9253);
nor U11989 (N_11989,N_7273,N_7510);
nand U11990 (N_11990,N_7973,N_8859);
nand U11991 (N_11991,N_6918,N_6495);
or U11992 (N_11992,N_8727,N_6424);
nand U11993 (N_11993,N_6660,N_9133);
nor U11994 (N_11994,N_8105,N_8391);
nor U11995 (N_11995,N_8665,N_8177);
and U11996 (N_11996,N_7879,N_7673);
and U11997 (N_11997,N_6570,N_6606);
nor U11998 (N_11998,N_8025,N_7351);
nor U11999 (N_11999,N_8064,N_8257);
or U12000 (N_12000,N_6846,N_7667);
nor U12001 (N_12001,N_7135,N_7786);
nor U12002 (N_12002,N_6934,N_8432);
nor U12003 (N_12003,N_8847,N_8136);
or U12004 (N_12004,N_7026,N_7118);
or U12005 (N_12005,N_7339,N_8908);
nand U12006 (N_12006,N_8254,N_7284);
or U12007 (N_12007,N_6691,N_6696);
xor U12008 (N_12008,N_6918,N_7812);
and U12009 (N_12009,N_8106,N_8371);
nor U12010 (N_12010,N_8450,N_8093);
and U12011 (N_12011,N_7742,N_7891);
nand U12012 (N_12012,N_6956,N_8717);
nor U12013 (N_12013,N_7317,N_7397);
or U12014 (N_12014,N_6747,N_9275);
or U12015 (N_12015,N_6335,N_7231);
and U12016 (N_12016,N_7661,N_8086);
or U12017 (N_12017,N_9183,N_7766);
nand U12018 (N_12018,N_8572,N_6717);
and U12019 (N_12019,N_6817,N_7993);
or U12020 (N_12020,N_7192,N_7515);
and U12021 (N_12021,N_8760,N_8191);
nor U12022 (N_12022,N_7753,N_7301);
xor U12023 (N_12023,N_8554,N_7608);
nor U12024 (N_12024,N_7282,N_7639);
or U12025 (N_12025,N_8047,N_6670);
xor U12026 (N_12026,N_6834,N_6903);
xor U12027 (N_12027,N_8210,N_8120);
nand U12028 (N_12028,N_8464,N_7521);
or U12029 (N_12029,N_9221,N_8254);
nor U12030 (N_12030,N_6786,N_6527);
and U12031 (N_12031,N_7111,N_7997);
or U12032 (N_12032,N_9256,N_9238);
and U12033 (N_12033,N_7446,N_8050);
or U12034 (N_12034,N_7554,N_9050);
and U12035 (N_12035,N_7595,N_7700);
or U12036 (N_12036,N_9287,N_6923);
nor U12037 (N_12037,N_8405,N_8799);
and U12038 (N_12038,N_7421,N_9245);
and U12039 (N_12039,N_6876,N_7217);
nand U12040 (N_12040,N_7943,N_8781);
xnor U12041 (N_12041,N_7801,N_8387);
and U12042 (N_12042,N_8644,N_6659);
or U12043 (N_12043,N_7047,N_7847);
nand U12044 (N_12044,N_7231,N_7549);
and U12045 (N_12045,N_6554,N_8614);
nor U12046 (N_12046,N_6651,N_8659);
xnor U12047 (N_12047,N_7443,N_7025);
xnor U12048 (N_12048,N_8974,N_9249);
nor U12049 (N_12049,N_9084,N_7161);
nor U12050 (N_12050,N_7143,N_6323);
nand U12051 (N_12051,N_6288,N_8356);
or U12052 (N_12052,N_9212,N_7592);
nor U12053 (N_12053,N_9191,N_7359);
xor U12054 (N_12054,N_8322,N_9343);
nand U12055 (N_12055,N_8783,N_7759);
nand U12056 (N_12056,N_8257,N_7174);
or U12057 (N_12057,N_7276,N_7128);
or U12058 (N_12058,N_7257,N_6890);
or U12059 (N_12059,N_7742,N_7065);
nor U12060 (N_12060,N_6845,N_8499);
and U12061 (N_12061,N_6535,N_8995);
nor U12062 (N_12062,N_7040,N_7816);
nand U12063 (N_12063,N_9011,N_8429);
or U12064 (N_12064,N_6881,N_7475);
and U12065 (N_12065,N_8885,N_8298);
nor U12066 (N_12066,N_6349,N_8917);
and U12067 (N_12067,N_7831,N_6798);
or U12068 (N_12068,N_7909,N_8069);
or U12069 (N_12069,N_8874,N_6782);
or U12070 (N_12070,N_8041,N_8661);
nand U12071 (N_12071,N_7690,N_7139);
nor U12072 (N_12072,N_8111,N_8698);
and U12073 (N_12073,N_8152,N_8083);
nand U12074 (N_12074,N_7183,N_9074);
nor U12075 (N_12075,N_7966,N_7057);
or U12076 (N_12076,N_7566,N_7740);
nor U12077 (N_12077,N_7485,N_6826);
and U12078 (N_12078,N_8639,N_8709);
and U12079 (N_12079,N_8098,N_7664);
nor U12080 (N_12080,N_6753,N_8009);
nand U12081 (N_12081,N_7103,N_9268);
or U12082 (N_12082,N_8422,N_7313);
or U12083 (N_12083,N_6301,N_8464);
nor U12084 (N_12084,N_6504,N_6399);
nand U12085 (N_12085,N_8321,N_6664);
or U12086 (N_12086,N_9119,N_8461);
or U12087 (N_12087,N_6344,N_8671);
or U12088 (N_12088,N_7191,N_7390);
and U12089 (N_12089,N_6959,N_8756);
or U12090 (N_12090,N_7698,N_7594);
xnor U12091 (N_12091,N_8192,N_7855);
or U12092 (N_12092,N_6411,N_7655);
nor U12093 (N_12093,N_6607,N_9263);
or U12094 (N_12094,N_7114,N_8032);
xnor U12095 (N_12095,N_7979,N_9286);
and U12096 (N_12096,N_7055,N_6499);
nor U12097 (N_12097,N_7603,N_7802);
nand U12098 (N_12098,N_6594,N_7322);
nand U12099 (N_12099,N_8451,N_6676);
or U12100 (N_12100,N_9253,N_7105);
nor U12101 (N_12101,N_6338,N_8393);
nor U12102 (N_12102,N_6454,N_6543);
nand U12103 (N_12103,N_7440,N_6716);
or U12104 (N_12104,N_6829,N_7359);
nand U12105 (N_12105,N_8789,N_6714);
nor U12106 (N_12106,N_8126,N_7269);
and U12107 (N_12107,N_8037,N_8704);
nor U12108 (N_12108,N_7628,N_9234);
and U12109 (N_12109,N_8841,N_7735);
nor U12110 (N_12110,N_8805,N_8484);
and U12111 (N_12111,N_9169,N_7617);
or U12112 (N_12112,N_8253,N_9256);
nand U12113 (N_12113,N_7928,N_8909);
nor U12114 (N_12114,N_6630,N_7674);
and U12115 (N_12115,N_6715,N_6724);
and U12116 (N_12116,N_6503,N_8428);
nor U12117 (N_12117,N_6581,N_8657);
xor U12118 (N_12118,N_9130,N_7062);
and U12119 (N_12119,N_8379,N_7766);
and U12120 (N_12120,N_7217,N_7317);
nand U12121 (N_12121,N_8616,N_8695);
xor U12122 (N_12122,N_6858,N_8739);
or U12123 (N_12123,N_9370,N_7611);
nor U12124 (N_12124,N_7107,N_8602);
or U12125 (N_12125,N_7356,N_6521);
or U12126 (N_12126,N_6365,N_9300);
nand U12127 (N_12127,N_8342,N_7694);
or U12128 (N_12128,N_6806,N_8901);
nor U12129 (N_12129,N_8194,N_6714);
and U12130 (N_12130,N_7784,N_6741);
nor U12131 (N_12131,N_8258,N_8388);
nor U12132 (N_12132,N_6309,N_7246);
and U12133 (N_12133,N_7207,N_7646);
nor U12134 (N_12134,N_7935,N_8877);
and U12135 (N_12135,N_8086,N_6705);
and U12136 (N_12136,N_6930,N_8270);
nor U12137 (N_12137,N_7293,N_6999);
and U12138 (N_12138,N_7375,N_6599);
nand U12139 (N_12139,N_8891,N_8065);
nand U12140 (N_12140,N_7167,N_6803);
nand U12141 (N_12141,N_8828,N_9007);
nor U12142 (N_12142,N_6921,N_7025);
nand U12143 (N_12143,N_7578,N_8150);
and U12144 (N_12144,N_8113,N_8795);
nor U12145 (N_12145,N_9340,N_6637);
or U12146 (N_12146,N_7876,N_6803);
nand U12147 (N_12147,N_9369,N_7654);
nand U12148 (N_12148,N_8439,N_7893);
and U12149 (N_12149,N_6530,N_9046);
nand U12150 (N_12150,N_6986,N_7804);
and U12151 (N_12151,N_8379,N_6375);
and U12152 (N_12152,N_9137,N_7065);
nor U12153 (N_12153,N_7259,N_9189);
and U12154 (N_12154,N_7783,N_9185);
and U12155 (N_12155,N_7627,N_8462);
xnor U12156 (N_12156,N_7365,N_9107);
nor U12157 (N_12157,N_8068,N_8458);
nand U12158 (N_12158,N_8073,N_8999);
or U12159 (N_12159,N_7109,N_7247);
or U12160 (N_12160,N_7883,N_6780);
or U12161 (N_12161,N_6855,N_6464);
or U12162 (N_12162,N_8683,N_8278);
or U12163 (N_12163,N_8155,N_8489);
and U12164 (N_12164,N_6644,N_8775);
or U12165 (N_12165,N_6337,N_7182);
nor U12166 (N_12166,N_9135,N_6505);
and U12167 (N_12167,N_6755,N_7044);
nand U12168 (N_12168,N_8558,N_6291);
nand U12169 (N_12169,N_9272,N_7923);
nor U12170 (N_12170,N_7779,N_7849);
and U12171 (N_12171,N_6750,N_7696);
and U12172 (N_12172,N_6995,N_7255);
and U12173 (N_12173,N_8831,N_9298);
or U12174 (N_12174,N_8660,N_7866);
and U12175 (N_12175,N_9103,N_8238);
nand U12176 (N_12176,N_6628,N_8323);
or U12177 (N_12177,N_8857,N_7013);
nand U12178 (N_12178,N_7671,N_7040);
and U12179 (N_12179,N_7535,N_7801);
xnor U12180 (N_12180,N_7358,N_8977);
nand U12181 (N_12181,N_9237,N_7576);
xor U12182 (N_12182,N_8163,N_7649);
or U12183 (N_12183,N_6821,N_6787);
nand U12184 (N_12184,N_6560,N_6810);
nor U12185 (N_12185,N_7884,N_6731);
or U12186 (N_12186,N_8023,N_6949);
nor U12187 (N_12187,N_6865,N_7291);
xor U12188 (N_12188,N_6269,N_6823);
or U12189 (N_12189,N_7253,N_8376);
or U12190 (N_12190,N_8761,N_7323);
xor U12191 (N_12191,N_6497,N_7311);
nand U12192 (N_12192,N_6411,N_6573);
nor U12193 (N_12193,N_8235,N_6296);
nor U12194 (N_12194,N_7306,N_7020);
nor U12195 (N_12195,N_8439,N_7458);
xnor U12196 (N_12196,N_6650,N_7052);
and U12197 (N_12197,N_8176,N_8331);
and U12198 (N_12198,N_7286,N_8298);
or U12199 (N_12199,N_9291,N_9282);
and U12200 (N_12200,N_8710,N_9166);
or U12201 (N_12201,N_6465,N_7479);
xnor U12202 (N_12202,N_8113,N_7419);
and U12203 (N_12203,N_7477,N_6717);
nand U12204 (N_12204,N_8436,N_7087);
nand U12205 (N_12205,N_9278,N_7245);
or U12206 (N_12206,N_9196,N_7847);
nand U12207 (N_12207,N_7479,N_8373);
nor U12208 (N_12208,N_8623,N_9358);
or U12209 (N_12209,N_8585,N_8201);
nand U12210 (N_12210,N_7429,N_7819);
nor U12211 (N_12211,N_8063,N_8576);
nand U12212 (N_12212,N_8340,N_7050);
or U12213 (N_12213,N_8430,N_7679);
or U12214 (N_12214,N_7034,N_7448);
nor U12215 (N_12215,N_8211,N_8079);
or U12216 (N_12216,N_6453,N_8398);
nor U12217 (N_12217,N_8920,N_7229);
xor U12218 (N_12218,N_7129,N_6501);
nor U12219 (N_12219,N_6582,N_6309);
xor U12220 (N_12220,N_8807,N_7238);
and U12221 (N_12221,N_7652,N_8659);
and U12222 (N_12222,N_8315,N_8828);
nand U12223 (N_12223,N_9346,N_7433);
nor U12224 (N_12224,N_8199,N_6263);
nand U12225 (N_12225,N_9322,N_8440);
nor U12226 (N_12226,N_8440,N_8610);
or U12227 (N_12227,N_8713,N_7415);
or U12228 (N_12228,N_8643,N_7282);
or U12229 (N_12229,N_7566,N_9049);
nor U12230 (N_12230,N_6415,N_7619);
nor U12231 (N_12231,N_8329,N_7475);
nand U12232 (N_12232,N_8716,N_7360);
nor U12233 (N_12233,N_6592,N_8876);
or U12234 (N_12234,N_8966,N_7371);
nor U12235 (N_12235,N_7382,N_6363);
xor U12236 (N_12236,N_7900,N_8870);
nor U12237 (N_12237,N_6342,N_8394);
nand U12238 (N_12238,N_9354,N_8129);
nor U12239 (N_12239,N_7469,N_7273);
nor U12240 (N_12240,N_6694,N_8490);
nor U12241 (N_12241,N_9341,N_6956);
and U12242 (N_12242,N_7687,N_9189);
and U12243 (N_12243,N_7036,N_9156);
and U12244 (N_12244,N_7320,N_8536);
xor U12245 (N_12245,N_8919,N_8766);
nor U12246 (N_12246,N_6530,N_7582);
nor U12247 (N_12247,N_6540,N_7110);
xnor U12248 (N_12248,N_6932,N_6943);
nand U12249 (N_12249,N_7041,N_7039);
or U12250 (N_12250,N_8634,N_6644);
and U12251 (N_12251,N_6541,N_7899);
or U12252 (N_12252,N_6814,N_8209);
nor U12253 (N_12253,N_7631,N_7577);
or U12254 (N_12254,N_6324,N_7097);
nor U12255 (N_12255,N_8372,N_7352);
and U12256 (N_12256,N_6832,N_9357);
and U12257 (N_12257,N_9106,N_6645);
and U12258 (N_12258,N_6255,N_8392);
and U12259 (N_12259,N_6983,N_8091);
or U12260 (N_12260,N_8337,N_6328);
nand U12261 (N_12261,N_9210,N_8585);
nand U12262 (N_12262,N_6402,N_6271);
xnor U12263 (N_12263,N_8116,N_8745);
nand U12264 (N_12264,N_8775,N_8407);
or U12265 (N_12265,N_9257,N_9107);
or U12266 (N_12266,N_7425,N_7424);
nand U12267 (N_12267,N_7927,N_8005);
or U12268 (N_12268,N_7103,N_7241);
nand U12269 (N_12269,N_6752,N_9260);
or U12270 (N_12270,N_6755,N_6973);
and U12271 (N_12271,N_8646,N_7367);
or U12272 (N_12272,N_8138,N_8404);
xor U12273 (N_12273,N_6782,N_7583);
or U12274 (N_12274,N_8444,N_8441);
or U12275 (N_12275,N_6389,N_8835);
or U12276 (N_12276,N_8313,N_8741);
nor U12277 (N_12277,N_7193,N_7659);
nor U12278 (N_12278,N_8904,N_6935);
or U12279 (N_12279,N_8925,N_6533);
nor U12280 (N_12280,N_8145,N_8989);
or U12281 (N_12281,N_7721,N_6988);
nand U12282 (N_12282,N_7529,N_6913);
nor U12283 (N_12283,N_8957,N_7100);
and U12284 (N_12284,N_8029,N_6286);
or U12285 (N_12285,N_7371,N_6563);
nand U12286 (N_12286,N_7503,N_8646);
nand U12287 (N_12287,N_7296,N_8858);
nand U12288 (N_12288,N_7901,N_7002);
nand U12289 (N_12289,N_9130,N_7478);
or U12290 (N_12290,N_7997,N_6977);
nand U12291 (N_12291,N_7245,N_6417);
nor U12292 (N_12292,N_9081,N_8321);
nand U12293 (N_12293,N_6981,N_6287);
xnor U12294 (N_12294,N_9149,N_7412);
xor U12295 (N_12295,N_7910,N_6984);
nor U12296 (N_12296,N_8232,N_9324);
nand U12297 (N_12297,N_8836,N_8084);
and U12298 (N_12298,N_8163,N_9058);
and U12299 (N_12299,N_8270,N_9371);
xor U12300 (N_12300,N_7038,N_8058);
or U12301 (N_12301,N_7744,N_6313);
nand U12302 (N_12302,N_6913,N_8908);
and U12303 (N_12303,N_6619,N_6674);
nor U12304 (N_12304,N_8704,N_9132);
or U12305 (N_12305,N_8055,N_8349);
and U12306 (N_12306,N_6666,N_7017);
nor U12307 (N_12307,N_8460,N_7849);
nand U12308 (N_12308,N_7639,N_8861);
nor U12309 (N_12309,N_6860,N_8274);
or U12310 (N_12310,N_8598,N_7957);
or U12311 (N_12311,N_6602,N_8620);
xnor U12312 (N_12312,N_9153,N_7990);
nand U12313 (N_12313,N_7105,N_8656);
xor U12314 (N_12314,N_7253,N_6439);
or U12315 (N_12315,N_8223,N_6501);
and U12316 (N_12316,N_7135,N_8595);
or U12317 (N_12317,N_8115,N_6493);
or U12318 (N_12318,N_8449,N_7802);
xnor U12319 (N_12319,N_7349,N_7939);
and U12320 (N_12320,N_9301,N_7398);
xnor U12321 (N_12321,N_7906,N_7255);
and U12322 (N_12322,N_7694,N_6404);
nand U12323 (N_12323,N_9353,N_7451);
nand U12324 (N_12324,N_8790,N_7431);
nand U12325 (N_12325,N_6428,N_7103);
xnor U12326 (N_12326,N_8593,N_6842);
xnor U12327 (N_12327,N_6694,N_8628);
nor U12328 (N_12328,N_7978,N_7549);
nor U12329 (N_12329,N_8201,N_6959);
nor U12330 (N_12330,N_6287,N_6898);
nor U12331 (N_12331,N_6548,N_9080);
nor U12332 (N_12332,N_8940,N_8524);
nor U12333 (N_12333,N_6446,N_8688);
nor U12334 (N_12334,N_8184,N_7942);
and U12335 (N_12335,N_8638,N_6984);
xor U12336 (N_12336,N_6915,N_8709);
or U12337 (N_12337,N_8994,N_7225);
and U12338 (N_12338,N_6836,N_9218);
nor U12339 (N_12339,N_7047,N_8676);
nor U12340 (N_12340,N_7872,N_9226);
nand U12341 (N_12341,N_9362,N_6482);
nand U12342 (N_12342,N_6949,N_8032);
nand U12343 (N_12343,N_8716,N_6615);
and U12344 (N_12344,N_7747,N_8592);
nand U12345 (N_12345,N_7229,N_8492);
and U12346 (N_12346,N_8146,N_6729);
or U12347 (N_12347,N_7427,N_6789);
nand U12348 (N_12348,N_8835,N_6771);
nand U12349 (N_12349,N_8047,N_7701);
and U12350 (N_12350,N_7414,N_6459);
xnor U12351 (N_12351,N_6483,N_8473);
or U12352 (N_12352,N_9373,N_7307);
and U12353 (N_12353,N_8688,N_8104);
nand U12354 (N_12354,N_6581,N_6327);
xor U12355 (N_12355,N_6265,N_8403);
and U12356 (N_12356,N_9111,N_9135);
nand U12357 (N_12357,N_7044,N_6311);
nor U12358 (N_12358,N_7396,N_9105);
or U12359 (N_12359,N_8121,N_8825);
nor U12360 (N_12360,N_6888,N_8018);
xnor U12361 (N_12361,N_7755,N_7981);
nor U12362 (N_12362,N_7369,N_7323);
or U12363 (N_12363,N_8768,N_9041);
nor U12364 (N_12364,N_8366,N_7843);
xnor U12365 (N_12365,N_6683,N_8170);
or U12366 (N_12366,N_7914,N_7246);
xnor U12367 (N_12367,N_7344,N_7463);
or U12368 (N_12368,N_8630,N_8769);
or U12369 (N_12369,N_8621,N_6408);
and U12370 (N_12370,N_8269,N_8200);
nand U12371 (N_12371,N_8003,N_7815);
xnor U12372 (N_12372,N_7971,N_7426);
nor U12373 (N_12373,N_9290,N_6668);
xor U12374 (N_12374,N_7248,N_7324);
nor U12375 (N_12375,N_7915,N_9125);
xor U12376 (N_12376,N_7618,N_7457);
or U12377 (N_12377,N_8597,N_8128);
and U12378 (N_12378,N_8512,N_8935);
nand U12379 (N_12379,N_9042,N_9259);
and U12380 (N_12380,N_8393,N_7110);
nand U12381 (N_12381,N_6819,N_8548);
nor U12382 (N_12382,N_8923,N_8962);
nor U12383 (N_12383,N_6760,N_6433);
or U12384 (N_12384,N_8745,N_6857);
nand U12385 (N_12385,N_7349,N_7326);
nand U12386 (N_12386,N_7522,N_7997);
nor U12387 (N_12387,N_7107,N_7567);
nand U12388 (N_12388,N_7404,N_8434);
or U12389 (N_12389,N_6548,N_9004);
xor U12390 (N_12390,N_8252,N_6783);
and U12391 (N_12391,N_7151,N_9328);
or U12392 (N_12392,N_8471,N_8113);
nor U12393 (N_12393,N_8783,N_8481);
nor U12394 (N_12394,N_8181,N_8345);
nand U12395 (N_12395,N_7350,N_6987);
nor U12396 (N_12396,N_7258,N_6740);
and U12397 (N_12397,N_7450,N_7983);
and U12398 (N_12398,N_9280,N_6459);
nor U12399 (N_12399,N_8406,N_9308);
and U12400 (N_12400,N_8928,N_9298);
xnor U12401 (N_12401,N_7064,N_6979);
or U12402 (N_12402,N_6525,N_7743);
and U12403 (N_12403,N_6589,N_8511);
nor U12404 (N_12404,N_7170,N_6857);
nand U12405 (N_12405,N_6492,N_7752);
and U12406 (N_12406,N_7999,N_8248);
nor U12407 (N_12407,N_8542,N_8039);
and U12408 (N_12408,N_9056,N_6397);
nand U12409 (N_12409,N_8855,N_7240);
xnor U12410 (N_12410,N_7943,N_9312);
nor U12411 (N_12411,N_8071,N_7116);
nand U12412 (N_12412,N_7785,N_8573);
nand U12413 (N_12413,N_7360,N_8389);
and U12414 (N_12414,N_7146,N_6914);
or U12415 (N_12415,N_8230,N_8590);
and U12416 (N_12416,N_9302,N_9291);
nand U12417 (N_12417,N_7265,N_8046);
and U12418 (N_12418,N_7408,N_9292);
or U12419 (N_12419,N_6997,N_8388);
nand U12420 (N_12420,N_8435,N_6888);
nor U12421 (N_12421,N_8270,N_6529);
or U12422 (N_12422,N_7360,N_8959);
nand U12423 (N_12423,N_7089,N_6743);
xnor U12424 (N_12424,N_8709,N_9001);
nand U12425 (N_12425,N_9266,N_6751);
or U12426 (N_12426,N_7300,N_8368);
and U12427 (N_12427,N_8221,N_8990);
xor U12428 (N_12428,N_6738,N_8980);
or U12429 (N_12429,N_7007,N_7814);
nand U12430 (N_12430,N_8347,N_6514);
nand U12431 (N_12431,N_8993,N_6713);
nand U12432 (N_12432,N_9246,N_8061);
or U12433 (N_12433,N_7955,N_6564);
and U12434 (N_12434,N_6494,N_8141);
and U12435 (N_12435,N_8131,N_9102);
xor U12436 (N_12436,N_7421,N_7248);
nor U12437 (N_12437,N_6453,N_8250);
and U12438 (N_12438,N_9157,N_6316);
and U12439 (N_12439,N_8068,N_8102);
xor U12440 (N_12440,N_8017,N_8916);
and U12441 (N_12441,N_8477,N_7363);
or U12442 (N_12442,N_7768,N_6399);
nand U12443 (N_12443,N_7344,N_6827);
nor U12444 (N_12444,N_7063,N_6654);
nand U12445 (N_12445,N_7029,N_8136);
and U12446 (N_12446,N_7903,N_6413);
nor U12447 (N_12447,N_7027,N_7564);
and U12448 (N_12448,N_7996,N_8016);
xor U12449 (N_12449,N_7584,N_7608);
nand U12450 (N_12450,N_9063,N_8849);
nor U12451 (N_12451,N_6433,N_8382);
or U12452 (N_12452,N_6604,N_7746);
or U12453 (N_12453,N_8232,N_8745);
nor U12454 (N_12454,N_6568,N_7970);
or U12455 (N_12455,N_8759,N_8848);
nand U12456 (N_12456,N_7955,N_7264);
or U12457 (N_12457,N_7966,N_6943);
nand U12458 (N_12458,N_7546,N_6922);
or U12459 (N_12459,N_8189,N_8334);
nor U12460 (N_12460,N_8532,N_6599);
and U12461 (N_12461,N_8407,N_8840);
nand U12462 (N_12462,N_7633,N_9237);
nor U12463 (N_12463,N_7448,N_7917);
nor U12464 (N_12464,N_8232,N_6701);
and U12465 (N_12465,N_6473,N_6648);
xor U12466 (N_12466,N_6751,N_8111);
and U12467 (N_12467,N_6981,N_7539);
nor U12468 (N_12468,N_8683,N_6712);
nor U12469 (N_12469,N_7846,N_6557);
xnor U12470 (N_12470,N_6765,N_8786);
nand U12471 (N_12471,N_6879,N_7776);
or U12472 (N_12472,N_9350,N_6992);
and U12473 (N_12473,N_8718,N_6457);
or U12474 (N_12474,N_7204,N_7405);
and U12475 (N_12475,N_6970,N_8271);
xnor U12476 (N_12476,N_6881,N_9229);
nand U12477 (N_12477,N_9333,N_7302);
or U12478 (N_12478,N_7724,N_7027);
xnor U12479 (N_12479,N_7154,N_7797);
nand U12480 (N_12480,N_6839,N_6588);
nand U12481 (N_12481,N_8758,N_8785);
and U12482 (N_12482,N_6710,N_6360);
nor U12483 (N_12483,N_8265,N_9184);
nand U12484 (N_12484,N_8784,N_7293);
xor U12485 (N_12485,N_9317,N_7426);
nand U12486 (N_12486,N_8976,N_7612);
and U12487 (N_12487,N_9296,N_7523);
nor U12488 (N_12488,N_8689,N_7198);
nand U12489 (N_12489,N_9079,N_6519);
nand U12490 (N_12490,N_8633,N_7012);
nor U12491 (N_12491,N_7293,N_7647);
nand U12492 (N_12492,N_6885,N_7045);
xor U12493 (N_12493,N_7533,N_9137);
nand U12494 (N_12494,N_8159,N_8771);
and U12495 (N_12495,N_8178,N_6763);
nand U12496 (N_12496,N_6564,N_8390);
or U12497 (N_12497,N_7876,N_8770);
nand U12498 (N_12498,N_6574,N_8349);
xnor U12499 (N_12499,N_6257,N_8174);
and U12500 (N_12500,N_12410,N_9868);
or U12501 (N_12501,N_11450,N_11001);
or U12502 (N_12502,N_10027,N_9597);
and U12503 (N_12503,N_9752,N_10203);
or U12504 (N_12504,N_10440,N_11232);
nand U12505 (N_12505,N_12344,N_10378);
xor U12506 (N_12506,N_10941,N_11841);
or U12507 (N_12507,N_10814,N_12231);
or U12508 (N_12508,N_11290,N_10508);
nor U12509 (N_12509,N_9781,N_9670);
nor U12510 (N_12510,N_12081,N_10765);
and U12511 (N_12511,N_9520,N_10822);
or U12512 (N_12512,N_11755,N_9620);
or U12513 (N_12513,N_9984,N_11452);
or U12514 (N_12514,N_9841,N_11224);
or U12515 (N_12515,N_12102,N_11368);
nor U12516 (N_12516,N_10148,N_11287);
nor U12517 (N_12517,N_9474,N_10946);
or U12518 (N_12518,N_12484,N_9462);
and U12519 (N_12519,N_12326,N_11939);
xor U12520 (N_12520,N_11797,N_12306);
nand U12521 (N_12521,N_10391,N_10471);
nand U12522 (N_12522,N_11218,N_10294);
nand U12523 (N_12523,N_12269,N_11093);
and U12524 (N_12524,N_10330,N_9491);
or U12525 (N_12525,N_11135,N_10301);
nor U12526 (N_12526,N_10468,N_10430);
and U12527 (N_12527,N_10190,N_10502);
or U12528 (N_12528,N_9917,N_10848);
nor U12529 (N_12529,N_11388,N_11745);
and U12530 (N_12530,N_11335,N_10965);
nand U12531 (N_12531,N_11882,N_10372);
or U12532 (N_12532,N_10002,N_9494);
nor U12533 (N_12533,N_10107,N_10449);
or U12534 (N_12534,N_11079,N_10083);
nand U12535 (N_12535,N_9649,N_9493);
and U12536 (N_12536,N_9519,N_12321);
nor U12537 (N_12537,N_11184,N_10269);
and U12538 (N_12538,N_11520,N_11554);
nor U12539 (N_12539,N_10927,N_11024);
nand U12540 (N_12540,N_11639,N_10735);
xnor U12541 (N_12541,N_10963,N_11676);
and U12542 (N_12542,N_9823,N_9742);
nand U12543 (N_12543,N_10284,N_12416);
nor U12544 (N_12544,N_12162,N_11713);
nand U12545 (N_12545,N_10337,N_9930);
nor U12546 (N_12546,N_10742,N_11375);
or U12547 (N_12547,N_12032,N_10703);
or U12548 (N_12548,N_10420,N_10135);
nand U12549 (N_12549,N_10004,N_10268);
xor U12550 (N_12550,N_10970,N_12130);
nor U12551 (N_12551,N_10078,N_11696);
xnor U12552 (N_12552,N_9825,N_11298);
nand U12553 (N_12553,N_10328,N_10580);
or U12554 (N_12554,N_9764,N_10839);
nand U12555 (N_12555,N_10369,N_11934);
nor U12556 (N_12556,N_9710,N_11245);
nor U12557 (N_12557,N_9961,N_9711);
and U12558 (N_12558,N_9587,N_12075);
nor U12559 (N_12559,N_9531,N_12006);
nand U12560 (N_12560,N_12235,N_11764);
nor U12561 (N_12561,N_9543,N_10241);
nor U12562 (N_12562,N_10724,N_10682);
nor U12563 (N_12563,N_9842,N_10071);
or U12564 (N_12564,N_11435,N_10650);
or U12565 (N_12565,N_12076,N_11010);
nand U12566 (N_12566,N_9640,N_10586);
or U12567 (N_12567,N_9403,N_11264);
nand U12568 (N_12568,N_10904,N_10755);
nor U12569 (N_12569,N_11201,N_9695);
and U12570 (N_12570,N_11162,N_10597);
or U12571 (N_12571,N_11836,N_12195);
nor U12572 (N_12572,N_9988,N_11629);
nand U12573 (N_12573,N_11947,N_9570);
xnor U12574 (N_12574,N_10496,N_10864);
nand U12575 (N_12575,N_10773,N_11609);
nor U12576 (N_12576,N_10697,N_11735);
xnor U12577 (N_12577,N_10286,N_11339);
and U12578 (N_12578,N_9458,N_11760);
nor U12579 (N_12579,N_10840,N_11805);
nor U12580 (N_12580,N_11969,N_9881);
or U12581 (N_12581,N_10295,N_9606);
nand U12582 (N_12582,N_10144,N_9685);
nand U12583 (N_12583,N_10776,N_9777);
nand U12584 (N_12584,N_10494,N_11033);
or U12585 (N_12585,N_12120,N_9870);
nor U12586 (N_12586,N_9614,N_11007);
or U12587 (N_12587,N_9628,N_11893);
nor U12588 (N_12588,N_11257,N_9435);
xnor U12589 (N_12589,N_9914,N_12337);
nand U12590 (N_12590,N_11381,N_10896);
nor U12591 (N_12591,N_11650,N_11559);
nand U12592 (N_12592,N_12180,N_9451);
and U12593 (N_12593,N_11046,N_12194);
nand U12594 (N_12594,N_9396,N_10416);
and U12595 (N_12595,N_10763,N_10110);
and U12596 (N_12596,N_9652,N_11250);
nor U12597 (N_12597,N_10595,N_11729);
or U12598 (N_12598,N_10231,N_9715);
nand U12599 (N_12599,N_12005,N_12174);
or U12600 (N_12600,N_11106,N_10237);
or U12601 (N_12601,N_10411,N_12428);
nor U12602 (N_12602,N_9768,N_11420);
and U12603 (N_12603,N_9753,N_9772);
nor U12604 (N_12604,N_9584,N_12134);
nand U12605 (N_12605,N_10234,N_11027);
and U12606 (N_12606,N_10618,N_10636);
nor U12607 (N_12607,N_11793,N_11921);
or U12608 (N_12608,N_10187,N_11100);
nor U12609 (N_12609,N_12425,N_11314);
nand U12610 (N_12610,N_9927,N_10335);
nor U12611 (N_12611,N_10945,N_10592);
and U12612 (N_12612,N_9774,N_10137);
and U12613 (N_12613,N_10455,N_10396);
and U12614 (N_12614,N_11295,N_10432);
or U12615 (N_12615,N_11321,N_9500);
and U12616 (N_12616,N_11794,N_10906);
nor U12617 (N_12617,N_10211,N_10583);
and U12618 (N_12618,N_12393,N_11053);
nor U12619 (N_12619,N_11225,N_11412);
and U12620 (N_12620,N_9588,N_11385);
nor U12621 (N_12621,N_10918,N_10731);
and U12622 (N_12622,N_11533,N_12118);
nor U12623 (N_12623,N_10092,N_11869);
or U12624 (N_12624,N_9903,N_10627);
xnor U12625 (N_12625,N_10448,N_11664);
nor U12626 (N_12626,N_12211,N_11081);
nand U12627 (N_12627,N_11874,N_11165);
xor U12628 (N_12628,N_10807,N_11564);
nor U12629 (N_12629,N_11401,N_11866);
and U12630 (N_12630,N_11700,N_9976);
nor U12631 (N_12631,N_11961,N_9720);
and U12632 (N_12632,N_9562,N_12127);
nor U12633 (N_12633,N_9566,N_9379);
nor U12634 (N_12634,N_10395,N_11179);
nand U12635 (N_12635,N_11424,N_10585);
or U12636 (N_12636,N_11627,N_11905);
nand U12637 (N_12637,N_9796,N_11671);
nand U12638 (N_12638,N_11394,N_10538);
nand U12639 (N_12639,N_11215,N_9585);
and U12640 (N_12640,N_10085,N_11431);
xor U12641 (N_12641,N_11367,N_11892);
nor U12642 (N_12642,N_11169,N_11510);
nor U12643 (N_12643,N_10133,N_10209);
nand U12644 (N_12644,N_11964,N_11606);
nand U12645 (N_12645,N_11739,N_12184);
nand U12646 (N_12646,N_11131,N_9873);
and U12647 (N_12647,N_11789,N_11877);
xor U12648 (N_12648,N_9946,N_11447);
or U12649 (N_12649,N_9681,N_11343);
xor U12650 (N_12650,N_12129,N_9957);
nand U12651 (N_12651,N_12288,N_10242);
xor U12652 (N_12652,N_10717,N_10521);
nand U12653 (N_12653,N_10457,N_10121);
xor U12654 (N_12654,N_10943,N_11369);
nor U12655 (N_12655,N_10908,N_10802);
xor U12656 (N_12656,N_11778,N_10379);
nor U12657 (N_12657,N_10748,N_10368);
and U12658 (N_12658,N_10619,N_10792);
or U12659 (N_12659,N_11115,N_11791);
nand U12660 (N_12660,N_12034,N_11453);
and U12661 (N_12661,N_10512,N_9632);
or U12662 (N_12662,N_12225,N_9838);
nor U12663 (N_12663,N_12398,N_9639);
and U12664 (N_12664,N_11055,N_9506);
xnor U12665 (N_12665,N_9446,N_10019);
nor U12666 (N_12666,N_12273,N_10949);
and U12667 (N_12667,N_9529,N_9673);
or U12668 (N_12668,N_10867,N_9763);
or U12669 (N_12669,N_10088,N_11479);
or U12670 (N_12670,N_11276,N_10948);
or U12671 (N_12671,N_11980,N_11175);
and U12672 (N_12672,N_12094,N_11732);
or U12673 (N_12673,N_11023,N_10947);
nand U12674 (N_12674,N_10020,N_10775);
and U12675 (N_12675,N_12031,N_10257);
nor U12676 (N_12676,N_10916,N_12254);
nand U12677 (N_12677,N_11396,N_11309);
or U12678 (N_12678,N_9511,N_10277);
and U12679 (N_12679,N_10493,N_10657);
nand U12680 (N_12680,N_10377,N_11800);
nor U12681 (N_12681,N_11665,N_9569);
or U12682 (N_12682,N_12475,N_11515);
and U12683 (N_12683,N_11300,N_10236);
or U12684 (N_12684,N_9682,N_12300);
xnor U12685 (N_12685,N_11084,N_11107);
nor U12686 (N_12686,N_10690,N_9440);
and U12687 (N_12687,N_9739,N_11407);
nand U12688 (N_12688,N_9641,N_11177);
nor U12689 (N_12689,N_9966,N_10439);
and U12690 (N_12690,N_9684,N_11119);
or U12691 (N_12691,N_11443,N_9980);
or U12692 (N_12692,N_11569,N_10159);
and U12693 (N_12693,N_11286,N_10045);
nand U12694 (N_12694,N_11283,N_10683);
xor U12695 (N_12695,N_11505,N_10550);
nand U12696 (N_12696,N_11281,N_9671);
xor U12697 (N_12697,N_11687,N_10143);
nand U12698 (N_12698,N_11563,N_9738);
nor U12699 (N_12699,N_9991,N_10499);
and U12700 (N_12700,N_10777,N_11472);
nand U12701 (N_12701,N_10291,N_11831);
nand U12702 (N_12702,N_11626,N_12001);
nand U12703 (N_12703,N_11152,N_9583);
nand U12704 (N_12704,N_9854,N_12210);
or U12705 (N_12705,N_10548,N_12304);
or U12706 (N_12706,N_10053,N_12479);
xnor U12707 (N_12707,N_10706,N_11054);
or U12708 (N_12708,N_12040,N_12320);
nor U12709 (N_12709,N_12041,N_11416);
nand U12710 (N_12710,N_10193,N_10033);
nand U12711 (N_12711,N_12328,N_12230);
nand U12712 (N_12712,N_10594,N_10172);
nand U12713 (N_12713,N_11073,N_12480);
nand U12714 (N_12714,N_11328,N_11379);
nand U12715 (N_12715,N_11460,N_9538);
or U12716 (N_12716,N_11973,N_10591);
nor U12717 (N_12717,N_10044,N_12299);
nand U12718 (N_12718,N_12250,N_11333);
nand U12719 (N_12719,N_12234,N_10977);
or U12720 (N_12720,N_9608,N_12445);
nand U12721 (N_12721,N_11349,N_10838);
nor U12722 (N_12722,N_11917,N_11589);
or U12723 (N_12723,N_11667,N_11903);
xor U12724 (N_12724,N_11875,N_11097);
nor U12725 (N_12725,N_11795,N_10264);
and U12726 (N_12726,N_11332,N_12116);
nand U12727 (N_12727,N_12206,N_9690);
or U12728 (N_12728,N_10425,N_9499);
nand U12729 (N_12729,N_12433,N_12310);
or U12730 (N_12730,N_12114,N_9848);
or U12731 (N_12731,N_11526,N_12429);
nor U12732 (N_12732,N_11701,N_10625);
nand U12733 (N_12733,N_9706,N_10076);
nor U12734 (N_12734,N_12220,N_12421);
and U12735 (N_12735,N_12448,N_9445);
or U12736 (N_12736,N_10727,N_10040);
and U12737 (N_12737,N_9634,N_11820);
xor U12738 (N_12738,N_11013,N_10983);
and U12739 (N_12739,N_12415,N_10542);
and U12740 (N_12740,N_11373,N_11551);
and U12741 (N_12741,N_11524,N_11421);
or U12742 (N_12742,N_10202,N_11262);
nor U12743 (N_12743,N_11469,N_12319);
nand U12744 (N_12744,N_11338,N_11012);
nand U12745 (N_12745,N_9655,N_12263);
nor U12746 (N_12746,N_9849,N_9895);
or U12747 (N_12747,N_9846,N_10556);
and U12748 (N_12748,N_10793,N_9479);
or U12749 (N_12749,N_10506,N_11751);
nor U12750 (N_12750,N_10737,N_10055);
nand U12751 (N_12751,N_11550,N_11132);
or U12752 (N_12752,N_11057,N_11694);
and U12753 (N_12753,N_9990,N_12322);
nor U12754 (N_12754,N_10113,N_10079);
xnor U12755 (N_12755,N_12271,N_10658);
or U12756 (N_12756,N_11906,N_10381);
nand U12757 (N_12757,N_9643,N_10060);
or U12758 (N_12758,N_12145,N_10794);
nand U12759 (N_12759,N_11766,N_12227);
nand U12760 (N_12760,N_11128,N_10582);
nand U12761 (N_12761,N_11014,N_11808);
nand U12762 (N_12762,N_9485,N_9782);
and U12763 (N_12763,N_10837,N_11914);
or U12764 (N_12764,N_11318,N_10451);
and U12765 (N_12765,N_11096,N_10680);
or U12766 (N_12766,N_10928,N_10723);
nor U12767 (N_12767,N_12143,N_11488);
nor U12768 (N_12768,N_9950,N_12488);
xnor U12769 (N_12769,N_10302,N_9567);
xnor U12770 (N_12770,N_9604,N_9830);
and U12771 (N_12771,N_10620,N_10100);
nor U12772 (N_12772,N_10520,N_9580);
or U12773 (N_12773,N_10632,N_9716);
nand U12774 (N_12774,N_10541,N_11835);
or U12775 (N_12775,N_11585,N_10890);
nor U12776 (N_12776,N_11355,N_9645);
nor U12777 (N_12777,N_10086,N_11608);
nor U12778 (N_12778,N_9871,N_11581);
nand U12779 (N_12779,N_11675,N_9644);
nand U12780 (N_12780,N_9769,N_9707);
xor U12781 (N_12781,N_9497,N_11943);
or U12782 (N_12782,N_11080,N_10528);
and U12783 (N_12783,N_11193,N_11727);
and U12784 (N_12784,N_11944,N_9415);
nand U12785 (N_12785,N_10146,N_11154);
nand U12786 (N_12786,N_11344,N_10299);
nand U12787 (N_12787,N_10487,N_10341);
nand U12788 (N_12788,N_12185,N_12060);
nor U12789 (N_12789,N_11704,N_12222);
and U12790 (N_12790,N_10179,N_10984);
nand U12791 (N_12791,N_11492,N_9664);
nor U12792 (N_12792,N_11932,N_10789);
nand U12793 (N_12793,N_9965,N_10177);
and U12794 (N_12794,N_11330,N_10705);
nand U12795 (N_12795,N_11830,N_12423);
or U12796 (N_12796,N_10996,N_12403);
nor U12797 (N_12797,N_10601,N_9481);
and U12798 (N_12798,N_10358,N_10589);
nor U12799 (N_12799,N_11736,N_11918);
nand U12800 (N_12800,N_10920,N_11026);
and U12801 (N_12801,N_10885,N_10570);
nand U12802 (N_12802,N_10571,N_10772);
nand U12803 (N_12803,N_11045,N_11315);
nand U12804 (N_12804,N_10424,N_11258);
nor U12805 (N_12805,N_10351,N_11904);
nor U12806 (N_12806,N_11773,N_9603);
and U12807 (N_12807,N_9425,N_11812);
nand U12808 (N_12808,N_12364,N_12178);
nand U12809 (N_12809,N_10898,N_11068);
nand U12810 (N_12810,N_10798,N_12440);
nor U12811 (N_12811,N_9509,N_11143);
and U12812 (N_12812,N_9648,N_9437);
nor U12813 (N_12813,N_11294,N_9721);
xnor U12814 (N_12814,N_11358,N_10648);
or U12815 (N_12815,N_11161,N_10799);
nor U12816 (N_12816,N_11485,N_11653);
nand U12817 (N_12817,N_10359,N_12142);
and U12818 (N_12818,N_11975,N_10955);
or U12819 (N_12819,N_9787,N_12157);
or U12820 (N_12820,N_10749,N_10509);
nand U12821 (N_12821,N_12019,N_10320);
nand U12822 (N_12822,N_10300,N_11908);
or U12823 (N_12823,N_9839,N_10954);
and U12824 (N_12824,N_10828,N_12239);
xor U12825 (N_12825,N_11644,N_12275);
nor U12826 (N_12826,N_9657,N_10347);
or U12827 (N_12827,N_9860,N_10901);
nor U12828 (N_12828,N_10819,N_9392);
nand U12829 (N_12829,N_11056,N_9941);
and U12830 (N_12830,N_10288,N_11928);
and U12831 (N_12831,N_9530,N_10791);
nand U12832 (N_12832,N_10293,N_12282);
and U12833 (N_12833,N_11669,N_10035);
nor U12834 (N_12834,N_9822,N_11242);
xor U12835 (N_12835,N_9422,N_10600);
or U12836 (N_12836,N_9916,N_10426);
and U12837 (N_12837,N_9388,N_11689);
xnor U12838 (N_12838,N_11968,N_11192);
nor U12839 (N_12839,N_9705,N_12384);
nand U12840 (N_12840,N_11094,N_10374);
or U12841 (N_12841,N_9843,N_11846);
or U12842 (N_12842,N_9663,N_11378);
nand U12843 (N_12843,N_10371,N_12377);
and U12844 (N_12844,N_10360,N_9890);
or U12845 (N_12845,N_10134,N_9426);
nand U12846 (N_12846,N_11804,N_11885);
nor U12847 (N_12847,N_9694,N_10080);
nor U12848 (N_12848,N_10373,N_10545);
nand U12849 (N_12849,N_10803,N_10830);
nand U12850 (N_12850,N_10221,N_11074);
nand U12851 (N_12851,N_10873,N_9886);
nand U12852 (N_12852,N_12066,N_11235);
and U12853 (N_12853,N_10292,N_11577);
nor U12854 (N_12854,N_9929,N_10176);
nand U12855 (N_12855,N_11004,N_10132);
nor U12856 (N_12856,N_12203,N_9488);
or U12857 (N_12857,N_11746,N_11386);
nor U12858 (N_12858,N_10871,N_9831);
nor U12859 (N_12859,N_12392,N_10997);
or U12860 (N_12860,N_12025,N_12069);
nand U12861 (N_12861,N_10279,N_10645);
nand U12862 (N_12862,N_11032,N_10101);
and U12863 (N_12863,N_11261,N_11734);
nand U12864 (N_12864,N_11611,N_10909);
nor U12865 (N_12865,N_9755,N_9453);
or U12866 (N_12866,N_11422,N_9476);
nand U12867 (N_12867,N_10480,N_10285);
nor U12868 (N_12868,N_12048,N_10549);
and U12869 (N_12869,N_9779,N_12097);
nor U12870 (N_12870,N_10326,N_12376);
nand U12871 (N_12871,N_10490,N_9611);
or U12872 (N_12872,N_10008,N_12389);
nand U12873 (N_12873,N_9869,N_11285);
nand U12874 (N_12874,N_9737,N_10750);
nor U12875 (N_12875,N_10223,N_10393);
xnor U12876 (N_12876,N_11855,N_11722);
nor U12877 (N_12877,N_11981,N_10778);
xnor U12878 (N_12878,N_11095,N_10801);
and U12879 (N_12879,N_9444,N_10246);
nand U12880 (N_12880,N_11002,N_10380);
nor U12881 (N_12881,N_10752,N_10046);
or U12882 (N_12882,N_9740,N_12061);
nor U12883 (N_12883,N_10445,N_10036);
xnor U12884 (N_12884,N_11677,N_9697);
nand U12885 (N_12885,N_10817,N_11540);
and U12886 (N_12886,N_11219,N_10175);
or U12887 (N_12887,N_12189,N_12274);
and U12888 (N_12888,N_11173,N_11486);
nor U12889 (N_12889,N_11353,N_10827);
or U12890 (N_12890,N_11036,N_10720);
and U12891 (N_12891,N_12303,N_10339);
nor U12892 (N_12892,N_11039,N_12305);
or U12893 (N_12893,N_12340,N_11529);
nand U12894 (N_12894,N_10478,N_10960);
nand U12895 (N_12895,N_11239,N_10059);
and U12896 (N_12896,N_11613,N_12113);
xnor U12897 (N_12897,N_12349,N_10385);
nor U12898 (N_12898,N_11887,N_10497);
and U12899 (N_12899,N_10721,N_10981);
nand U12900 (N_12900,N_11203,N_10766);
and U12901 (N_12901,N_10228,N_9610);
nand U12902 (N_12902,N_10857,N_9800);
and U12903 (N_12903,N_9743,N_9638);
and U12904 (N_12904,N_11635,N_10155);
nand U12905 (N_12905,N_11817,N_12351);
nor U12906 (N_12906,N_12387,N_10307);
and U12907 (N_12907,N_9999,N_11155);
nor U12908 (N_12908,N_11267,N_11845);
nand U12909 (N_12909,N_11718,N_11110);
and U12910 (N_12910,N_10441,N_11426);
nand U12911 (N_12911,N_10353,N_10786);
and U12912 (N_12912,N_9533,N_10122);
nor U12913 (N_12913,N_9963,N_9836);
nor U12914 (N_12914,N_10637,N_10073);
nor U12915 (N_12915,N_10780,N_12151);
or U12916 (N_12916,N_11979,N_11478);
nor U12917 (N_12917,N_9733,N_11832);
and U12918 (N_12918,N_11502,N_9808);
and U12919 (N_12919,N_12125,N_10310);
or U12920 (N_12920,N_11915,N_12408);
nor U12921 (N_12921,N_11138,N_11900);
nand U12922 (N_12922,N_11570,N_10082);
nand U12923 (N_12923,N_10452,N_9635);
nand U12924 (N_12924,N_11061,N_12456);
nor U12925 (N_12925,N_12270,N_9623);
and U12926 (N_12926,N_10068,N_10093);
and U12927 (N_12927,N_9933,N_11198);
nor U12928 (N_12928,N_10423,N_11465);
xor U12929 (N_12929,N_11482,N_11574);
xor U12930 (N_12930,N_11645,N_11436);
nand U12931 (N_12931,N_10875,N_11038);
nor U12932 (N_12932,N_10072,N_10476);
nand U12933 (N_12933,N_11157,N_9527);
and U12934 (N_12934,N_12447,N_10156);
or U12935 (N_12935,N_12316,N_9581);
nor U12936 (N_12936,N_9910,N_11935);
or U12937 (N_12937,N_10474,N_9773);
nor U12938 (N_12938,N_10563,N_10410);
or U12939 (N_12939,N_11433,N_9791);
nor U12940 (N_12940,N_11989,N_11767);
and U12941 (N_12941,N_11838,N_10039);
nand U12942 (N_12942,N_10930,N_12205);
nand U12943 (N_12943,N_10488,N_11252);
and U12944 (N_12944,N_11260,N_11933);
xor U12945 (N_12945,N_10034,N_11233);
and U12946 (N_12946,N_10089,N_12465);
or U12947 (N_12947,N_12087,N_9400);
and U12948 (N_12948,N_11658,N_10925);
and U12949 (N_12949,N_9879,N_10675);
and U12950 (N_12950,N_11890,N_9745);
or U12951 (N_12951,N_11592,N_10095);
nor U12952 (N_12952,N_11337,N_11307);
or U12953 (N_12953,N_11561,N_9922);
and U12954 (N_12954,N_9959,N_9680);
or U12955 (N_12955,N_11186,N_10051);
nor U12956 (N_12956,N_11197,N_10181);
xor U12957 (N_12957,N_11991,N_10511);
or U12958 (N_12958,N_10163,N_9935);
and U12959 (N_12959,N_10399,N_12251);
nor U12960 (N_12960,N_11047,N_11451);
nand U12961 (N_12961,N_10329,N_12407);
and U12962 (N_12962,N_10167,N_11000);
xor U12963 (N_12963,N_12082,N_12196);
nand U12964 (N_12964,N_10931,N_10868);
xor U12965 (N_12965,N_11384,N_11438);
nand U12966 (N_12966,N_10579,N_9821);
nor U12967 (N_12967,N_10016,N_10973);
or U12968 (N_12968,N_12495,N_9398);
nor U12969 (N_12969,N_12236,N_11850);
nand U12970 (N_12970,N_10312,N_9665);
nor U12971 (N_12971,N_11308,N_12276);
and U12972 (N_12972,N_9601,N_12202);
or U12973 (N_12973,N_11723,N_11527);
and U12974 (N_12974,N_11069,N_11610);
or U12975 (N_12975,N_10481,N_10783);
nand U12976 (N_12976,N_10774,N_10877);
and U12977 (N_12977,N_9911,N_11326);
nor U12978 (N_12978,N_10531,N_11126);
xor U12979 (N_12979,N_9947,N_11522);
nor U12980 (N_12980,N_9545,N_12167);
or U12981 (N_12981,N_12459,N_12381);
and U12982 (N_12982,N_9883,N_10205);
and U12983 (N_12983,N_10469,N_10306);
and U12984 (N_12984,N_11842,N_11634);
or U12985 (N_12985,N_9878,N_12168);
nand U12986 (N_12986,N_11387,N_9418);
nand U12987 (N_12987,N_11590,N_10180);
nor U12988 (N_12988,N_10647,N_11604);
or U12989 (N_12989,N_10050,N_10956);
nand U12990 (N_12990,N_9393,N_12046);
nand U12991 (N_12991,N_10689,N_11822);
or U12992 (N_12992,N_10421,N_9709);
nor U12993 (N_12993,N_9921,N_10437);
and U12994 (N_12994,N_11796,N_11573);
nor U12995 (N_12995,N_11752,N_11174);
nand U12996 (N_12996,N_9667,N_11114);
xnor U12997 (N_12997,N_12063,N_12311);
nor U12998 (N_12998,N_9377,N_10011);
nand U12999 (N_12999,N_9571,N_9487);
and U13000 (N_13000,N_10376,N_10355);
nand U13001 (N_13001,N_12119,N_11586);
nor U13002 (N_13002,N_10823,N_10845);
nand U13003 (N_13003,N_11166,N_11962);
nor U13004 (N_13004,N_10524,N_11471);
xor U13005 (N_13005,N_12244,N_11747);
nor U13006 (N_13006,N_9985,N_11316);
xnor U13007 (N_13007,N_10529,N_9411);
nand U13008 (N_13008,N_11603,N_9450);
nand U13009 (N_13009,N_9973,N_10751);
or U13010 (N_13010,N_10673,N_11702);
nand U13011 (N_13011,N_11030,N_9795);
or U13012 (N_13012,N_9750,N_10314);
or U13013 (N_13013,N_11448,N_10829);
and U13014 (N_13014,N_12062,N_10746);
or U13015 (N_13015,N_11619,N_10081);
or U13016 (N_13016,N_10250,N_12080);
xor U13017 (N_13017,N_10652,N_11632);
xor U13018 (N_13018,N_10206,N_10014);
or U13019 (N_13019,N_10869,N_10482);
and U13020 (N_13020,N_10405,N_12405);
nand U13021 (N_13021,N_9407,N_12138);
nor U13022 (N_13022,N_9590,N_10168);
and U13023 (N_13023,N_10387,N_10951);
nand U13024 (N_13024,N_10876,N_10934);
or U13025 (N_13025,N_10030,N_10674);
xnor U13026 (N_13026,N_12074,N_11116);
nor U13027 (N_13027,N_11580,N_11127);
nor U13028 (N_13028,N_11279,N_9932);
or U13029 (N_13029,N_12213,N_11019);
nor U13030 (N_13030,N_10781,N_12498);
nand U13031 (N_13031,N_10577,N_11521);
or U13032 (N_13032,N_10661,N_10362);
or U13033 (N_13033,N_9741,N_10240);
and U13034 (N_13034,N_9827,N_11924);
and U13035 (N_13035,N_10498,N_11409);
and U13036 (N_13036,N_10006,N_12295);
nor U13037 (N_13037,N_11693,N_9757);
nand U13038 (N_13038,N_11456,N_12382);
or U13039 (N_13039,N_11552,N_12132);
nand U13040 (N_13040,N_11506,N_12085);
and U13041 (N_13041,N_10893,N_11228);
nand U13042 (N_13042,N_11076,N_12240);
nand U13043 (N_13043,N_11303,N_11599);
and U13044 (N_13044,N_9789,N_10226);
or U13045 (N_13045,N_10733,N_10923);
and U13046 (N_13046,N_9565,N_11640);
nand U13047 (N_13047,N_10105,N_9853);
or U13048 (N_13048,N_10287,N_11357);
or U13049 (N_13049,N_11458,N_12432);
and U13050 (N_13050,N_11859,N_10989);
and U13051 (N_13051,N_10470,N_12248);
or U13052 (N_13052,N_12044,N_12033);
nor U13053 (N_13053,N_11414,N_11188);
nand U13054 (N_13054,N_12491,N_12362);
and U13055 (N_13055,N_10979,N_11136);
xor U13056 (N_13056,N_10345,N_10640);
nand U13057 (N_13057,N_11359,N_11238);
or U13058 (N_13058,N_10108,N_12233);
nand U13059 (N_13059,N_11516,N_10227);
or U13060 (N_13060,N_11756,N_10967);
and U13061 (N_13061,N_11549,N_10559);
nor U13062 (N_13062,N_12297,N_11299);
nor U13063 (N_13063,N_12221,N_9577);
and U13064 (N_13064,N_10711,N_10350);
xnor U13065 (N_13065,N_10835,N_11513);
nand U13066 (N_13066,N_12370,N_10450);
nand U13067 (N_13067,N_10598,N_11668);
xor U13068 (N_13068,N_9475,N_10075);
nor U13069 (N_13069,N_12226,N_11731);
or U13070 (N_13070,N_10136,N_10679);
nand U13071 (N_13071,N_9594,N_10160);
or U13072 (N_13072,N_11117,N_10599);
and U13073 (N_13073,N_12332,N_11710);
and U13074 (N_13074,N_10244,N_10260);
and U13075 (N_13075,N_9486,N_10037);
nand U13076 (N_13076,N_11191,N_12121);
nor U13077 (N_13077,N_11828,N_11364);
nand U13078 (N_13078,N_11077,N_10937);
nor U13079 (N_13079,N_10821,N_11725);
and U13080 (N_13080,N_11977,N_11404);
nand U13081 (N_13081,N_9595,N_12307);
or U13082 (N_13082,N_12173,N_12367);
nand U13083 (N_13083,N_10605,N_12397);
nor U13084 (N_13084,N_11158,N_9880);
and U13085 (N_13085,N_9882,N_10516);
nor U13086 (N_13086,N_9524,N_10692);
and U13087 (N_13087,N_11052,N_9460);
or U13088 (N_13088,N_10646,N_10003);
nand U13089 (N_13089,N_11098,N_9856);
and U13090 (N_13090,N_11967,N_10921);
or U13091 (N_13091,N_9887,N_11395);
nor U13092 (N_13092,N_11625,N_11528);
xnor U13093 (N_13093,N_9799,N_11113);
nand U13094 (N_13094,N_11199,N_10922);
and U13095 (N_13095,N_9771,N_9790);
or U13096 (N_13096,N_11123,N_11497);
nor U13097 (N_13097,N_12165,N_11868);
nor U13098 (N_13098,N_10500,N_9971);
nor U13099 (N_13099,N_10484,N_10334);
nand U13100 (N_13100,N_9642,N_11881);
and U13101 (N_13101,N_10744,N_12272);
and U13102 (N_13102,N_11200,N_10322);
and U13103 (N_13103,N_11814,N_9507);
nor U13104 (N_13104,N_10757,N_9420);
and U13105 (N_13105,N_11463,N_9688);
or U13106 (N_13106,N_11769,N_9812);
and U13107 (N_13107,N_9759,N_12375);
and U13108 (N_13108,N_11083,N_11772);
nor U13109 (N_13109,N_12458,N_9872);
xnor U13110 (N_13110,N_11945,N_10631);
or U13111 (N_13111,N_12329,N_11620);
nand U13112 (N_13112,N_12422,N_11878);
nor U13113 (N_13113,N_10539,N_9646);
or U13114 (N_13114,N_10165,N_11821);
or U13115 (N_13115,N_12318,N_11211);
and U13116 (N_13116,N_11867,N_12007);
xor U13117 (N_13117,N_12451,N_10384);
and U13118 (N_13118,N_9857,N_9723);
and U13119 (N_13119,N_10026,N_11495);
nand U13120 (N_13120,N_12036,N_9983);
nand U13121 (N_13121,N_11370,N_11405);
and U13122 (N_13122,N_10929,N_11699);
nand U13123 (N_13123,N_11317,N_9953);
xor U13124 (N_13124,N_9701,N_11206);
nand U13125 (N_13125,N_11737,N_10505);
nand U13126 (N_13126,N_9402,N_10198);
nand U13127 (N_13127,N_10590,N_10677);
nor U13128 (N_13128,N_11296,N_11415);
xnor U13129 (N_13129,N_10924,N_9861);
nand U13130 (N_13130,N_10564,N_10942);
or U13131 (N_13131,N_10966,N_10126);
nand U13132 (N_13132,N_10255,N_11125);
or U13133 (N_13133,N_11839,N_11523);
xor U13134 (N_13134,N_10884,N_11873);
nor U13135 (N_13135,N_10654,N_11329);
and U13136 (N_13136,N_10769,N_9482);
or U13137 (N_13137,N_10660,N_11066);
nor U13138 (N_13138,N_12345,N_10054);
or U13139 (N_13139,N_9852,N_10483);
and U13140 (N_13140,N_10321,N_10115);
or U13141 (N_13141,N_10874,N_12357);
nor U13142 (N_13142,N_12057,N_9693);
nand U13143 (N_13143,N_9589,N_12112);
or U13144 (N_13144,N_11342,N_11698);
nand U13145 (N_13145,N_12079,N_11009);
and U13146 (N_13146,N_12265,N_11771);
nor U13147 (N_13147,N_10811,N_11744);
nor U13148 (N_13148,N_11459,N_10104);
and U13149 (N_13149,N_11651,N_9465);
nand U13150 (N_13150,N_10324,N_12477);
nand U13151 (N_13151,N_10990,N_11636);
or U13152 (N_13152,N_11493,N_11040);
and U13153 (N_13153,N_11825,N_9702);
and U13154 (N_13154,N_11164,N_11750);
and U13155 (N_13155,N_10404,N_12022);
or U13156 (N_13156,N_10015,N_10681);
nor U13157 (N_13157,N_12473,N_11958);
nand U13158 (N_13158,N_12368,N_11065);
nor U13159 (N_13159,N_9677,N_9672);
xnor U13160 (N_13160,N_10861,N_12253);
or U13161 (N_13161,N_9780,N_11491);
nand U13162 (N_13162,N_10743,N_11615);
nor U13163 (N_13163,N_11195,N_11255);
or U13164 (N_13164,N_11146,N_10413);
nor U13165 (N_13165,N_11222,N_10005);
and U13166 (N_13166,N_10220,N_10894);
nor U13167 (N_13167,N_11168,N_12453);
xnor U13168 (N_13168,N_9972,N_9889);
nand U13169 (N_13169,N_9503,N_9837);
or U13170 (N_13170,N_12363,N_11788);
nand U13171 (N_13171,N_12045,N_10782);
nand U13172 (N_13172,N_10612,N_10912);
or U13173 (N_13173,N_12487,N_9455);
nand U13174 (N_13174,N_11854,N_9904);
and U13175 (N_13175,N_12043,N_11361);
nand U13176 (N_13176,N_12058,N_10447);
and U13177 (N_13177,N_9596,N_12216);
or U13178 (N_13178,N_10787,N_11861);
and U13179 (N_13179,N_11251,N_10573);
nor U13180 (N_13180,N_10406,N_10094);
or U13181 (N_13181,N_9429,N_11954);
nand U13182 (N_13182,N_11872,N_10961);
and U13183 (N_13183,N_11090,N_11966);
nor U13184 (N_13184,N_9586,N_10461);
nand U13185 (N_13185,N_11512,N_10913);
xor U13186 (N_13186,N_11247,N_9704);
nor U13187 (N_13187,N_12083,N_9598);
nand U13188 (N_13188,N_9654,N_9431);
xnor U13189 (N_13189,N_9386,N_9775);
nor U13190 (N_13190,N_12144,N_11560);
xor U13191 (N_13191,N_10854,N_11306);
nand U13192 (N_13192,N_11811,N_9384);
nand U13193 (N_13193,N_12490,N_10370);
nor U13194 (N_13194,N_9471,N_11362);
and U13195 (N_13195,N_12309,N_12027);
nor U13196 (N_13196,N_11473,N_10120);
and U13197 (N_13197,N_10125,N_9544);
nor U13198 (N_13198,N_9631,N_9528);
nor U13199 (N_13199,N_10976,N_12467);
and U13200 (N_13200,N_11578,N_9996);
or U13201 (N_13201,N_10653,N_11035);
nand U13202 (N_13202,N_12190,N_10809);
and U13203 (N_13203,N_11927,N_9484);
or U13204 (N_13204,N_12296,N_11272);
nor U13205 (N_13205,N_9502,N_10194);
xnor U13206 (N_13206,N_11774,N_9626);
or U13207 (N_13207,N_11142,N_12372);
nor U13208 (N_13208,N_12154,N_11331);
nor U13209 (N_13209,N_10888,N_10021);
nand U13210 (N_13210,N_10593,N_11950);
nand U13211 (N_13211,N_9809,N_9835);
or U13212 (N_13212,N_12373,N_9692);
nand U13213 (N_13213,N_11280,N_10555);
nand U13214 (N_13214,N_12466,N_12232);
or U13215 (N_13215,N_9760,N_10892);
nor U13216 (N_13216,N_10256,N_9826);
nor U13217 (N_13217,N_11496,N_9915);
and U13218 (N_13218,N_11716,N_9951);
and U13219 (N_13219,N_12077,N_12217);
nand U13220 (N_13220,N_9734,N_9477);
nand U13221 (N_13221,N_11942,N_11120);
and U13222 (N_13222,N_11579,N_12135);
and U13223 (N_13223,N_9483,N_10676);
and U13224 (N_13224,N_12176,N_12198);
xnor U13225 (N_13225,N_12149,N_11641);
and U13226 (N_13226,N_11685,N_10201);
xnor U13227 (N_13227,N_12155,N_9498);
or U13228 (N_13228,N_9810,N_11011);
and U13229 (N_13229,N_10131,N_11963);
nand U13230 (N_13230,N_12388,N_9718);
and U13231 (N_13231,N_10427,N_10964);
nor U13232 (N_13232,N_10454,N_9449);
and U13233 (N_13233,N_11034,N_12499);
xor U13234 (N_13234,N_12413,N_11282);
or U13235 (N_13235,N_11327,N_11277);
nand U13236 (N_13236,N_10238,N_12038);
or U13237 (N_13237,N_9452,N_12289);
and U13238 (N_13238,N_10278,N_11461);
nor U13239 (N_13239,N_10272,N_10588);
nor U13240 (N_13240,N_10214,N_10383);
nor U13241 (N_13241,N_11470,N_11647);
and U13242 (N_13242,N_11060,N_11457);
and U13243 (N_13243,N_10767,N_11230);
nor U13244 (N_13244,N_9703,N_12419);
or U13245 (N_13245,N_11946,N_11519);
nand U13246 (N_13246,N_10696,N_12186);
and U13247 (N_13247,N_12402,N_12298);
and U13248 (N_13248,N_10031,N_10608);
or U13249 (N_13249,N_12391,N_11530);
or U13250 (N_13250,N_11856,N_11508);
nor U13251 (N_13251,N_12104,N_11883);
nand U13252 (N_13252,N_12049,N_11088);
and U13253 (N_13253,N_9934,N_12424);
and U13254 (N_13254,N_11888,N_12172);
nand U13255 (N_13255,N_9463,N_11951);
or U13256 (N_13256,N_10386,N_12158);
nor U13257 (N_13257,N_11678,N_11227);
or U13258 (N_13258,N_11305,N_9439);
or U13259 (N_13259,N_10042,N_9540);
or U13260 (N_13260,N_11929,N_10210);
nand U13261 (N_13261,N_12286,N_10719);
xor U13262 (N_13262,N_11937,N_10806);
nor U13263 (N_13263,N_11572,N_11017);
xnor U13264 (N_13264,N_11638,N_12073);
xnor U13265 (N_13265,N_10340,N_11706);
or U13266 (N_13266,N_10161,N_11291);
nand U13267 (N_13267,N_10400,N_10764);
xor U13268 (N_13268,N_10154,N_9845);
nor U13269 (N_13269,N_9615,N_10048);
nor U13270 (N_13270,N_11244,N_10547);
or U13271 (N_13271,N_10962,N_9847);
or U13272 (N_13272,N_12207,N_12361);
and U13273 (N_13273,N_10953,N_10013);
and U13274 (N_13274,N_12052,N_9978);
nor U13275 (N_13275,N_10872,N_11899);
xnor U13276 (N_13276,N_10784,N_9728);
nand U13277 (N_13277,N_10842,N_12455);
xnor U13278 (N_13278,N_10736,N_11270);
or U13279 (N_13279,N_10218,N_11799);
or U13280 (N_13280,N_9952,N_12360);
nor U13281 (N_13281,N_9858,N_10818);
nand U13282 (N_13282,N_12278,N_10103);
and U13283 (N_13283,N_12463,N_10687);
xor U13284 (N_13284,N_11894,N_11724);
and U13285 (N_13285,N_11442,N_10662);
nand U13286 (N_13286,N_9442,N_11189);
or U13287 (N_13287,N_10858,N_12056);
xnor U13288 (N_13288,N_11539,N_11993);
or U13289 (N_13289,N_9945,N_9691);
or U13290 (N_13290,N_11784,N_10492);
or U13291 (N_13291,N_11754,N_11372);
nand U13292 (N_13292,N_12108,N_12099);
and U13293 (N_13293,N_11787,N_10392);
nand U13294 (N_13294,N_11759,N_12257);
xnor U13295 (N_13295,N_11434,N_11785);
and U13296 (N_13296,N_11417,N_12259);
and U13297 (N_13297,N_12212,N_12464);
nor U13298 (N_13298,N_11273,N_11949);
and U13299 (N_13299,N_10671,N_11432);
nand U13300 (N_13300,N_12444,N_10375);
and U13301 (N_13301,N_11205,N_11051);
and U13302 (N_13302,N_9748,N_11190);
and U13303 (N_13303,N_12140,N_11692);
or U13304 (N_13304,N_12371,N_10576);
nor U13305 (N_13305,N_11568,N_9964);
and U13306 (N_13306,N_9532,N_9801);
or U13307 (N_13307,N_10638,N_9512);
xnor U13308 (N_13308,N_10057,N_10422);
nor U13309 (N_13309,N_10366,N_11393);
nor U13310 (N_13310,N_10022,N_9783);
or U13311 (N_13311,N_9513,N_11596);
or U13312 (N_13312,N_10382,N_10917);
nand U13313 (N_13313,N_9441,N_11489);
nand U13314 (N_13314,N_10504,N_9918);
nor U13315 (N_13315,N_10865,N_9998);
and U13316 (N_13316,N_11490,N_11122);
or U13317 (N_13317,N_11231,N_11480);
nand U13318 (N_13318,N_11833,N_10153);
nand U13319 (N_13319,N_12312,N_10245);
or U13320 (N_13320,N_10064,N_9467);
nand U13321 (N_13321,N_11441,N_12039);
xnor U13322 (N_13322,N_12374,N_11809);
and U13323 (N_13323,N_10607,N_11714);
or U13324 (N_13324,N_9756,N_10536);
and U13325 (N_13325,N_10204,N_12133);
nor U13326 (N_13326,N_12159,N_11446);
and U13327 (N_13327,N_11236,N_11670);
nor U13328 (N_13328,N_9992,N_9785);
or U13329 (N_13329,N_10119,N_10007);
and U13330 (N_13330,N_11660,N_12192);
nand U13331 (N_13331,N_10394,N_10557);
xnor U13332 (N_13332,N_11071,N_12301);
nand U13333 (N_13333,N_11212,N_11323);
and U13334 (N_13334,N_11895,N_10308);
nand U13335 (N_13335,N_9574,N_12053);
nor U13336 (N_13336,N_11576,N_10415);
or U13337 (N_13337,N_9726,N_9979);
nor U13338 (N_13338,N_9659,N_11957);
xnor U13339 (N_13339,N_11376,N_10709);
xor U13340 (N_13340,N_9891,N_10233);
and U13341 (N_13341,N_11348,N_12246);
nor U13342 (N_13342,N_10208,N_9433);
and U13343 (N_13343,N_11208,N_11320);
nand U13344 (N_13344,N_9730,N_10253);
nor U13345 (N_13345,N_10639,N_9855);
or U13346 (N_13346,N_11425,N_11028);
or U13347 (N_13347,N_9390,N_11847);
and U13348 (N_13348,N_11707,N_10225);
nor U13349 (N_13349,N_10664,N_11265);
nor U13350 (N_13350,N_9807,N_12255);
nor U13351 (N_13351,N_10489,N_10017);
nand U13352 (N_13352,N_12065,N_9746);
nand U13353 (N_13353,N_9700,N_11085);
nand U13354 (N_13354,N_11891,N_9602);
nor U13355 (N_13355,N_11761,N_12485);
nand U13356 (N_13356,N_9937,N_9907);
nor U13357 (N_13357,N_11380,N_10063);
nor U13358 (N_13358,N_10919,N_11558);
nor U13359 (N_13359,N_11837,N_11567);
and U13360 (N_13360,N_11511,N_10911);
and U13361 (N_13361,N_9804,N_10718);
or U13362 (N_13362,N_11288,N_10635);
nor U13363 (N_13363,N_10695,N_9473);
nor U13364 (N_13364,N_11655,N_9784);
or U13365 (N_13365,N_9975,N_11477);
nand U13366 (N_13366,N_12342,N_11340);
nand U13367 (N_13367,N_10851,N_10980);
or U13368 (N_13368,N_10832,N_11948);
nand U13369 (N_13369,N_10024,N_12262);
nand U13370 (N_13370,N_10356,N_10271);
xnor U13371 (N_13371,N_11217,N_9770);
and U13372 (N_13372,N_11044,N_11449);
nand U13373 (N_13373,N_10863,N_10188);
or U13374 (N_13374,N_11301,N_10729);
xnor U13375 (N_13375,N_9522,N_9592);
and U13376 (N_13376,N_9811,N_10684);
nand U13377 (N_13377,N_10147,N_11753);
nand U13378 (N_13378,N_12059,N_10795);
nand U13379 (N_13379,N_11742,N_11413);
nor U13380 (N_13380,N_10098,N_11062);
nand U13381 (N_13381,N_11408,N_10762);
nor U13382 (N_13382,N_11160,N_11149);
and U13383 (N_13383,N_9521,N_11410);
nand U13384 (N_13384,N_9380,N_12200);
nor U13385 (N_13385,N_10621,N_9829);
xnor U13386 (N_13386,N_10971,N_9712);
and U13387 (N_13387,N_9541,N_10318);
or U13388 (N_13388,N_11015,N_10722);
and U13389 (N_13389,N_9609,N_10289);
nor U13390 (N_13390,N_11911,N_10141);
and U13391 (N_13391,N_9888,N_9679);
and U13392 (N_13392,N_9417,N_9573);
nor U13393 (N_13393,N_10077,N_9555);
or U13394 (N_13394,N_12169,N_11749);
or U13395 (N_13395,N_10672,N_9893);
or U13396 (N_13396,N_9876,N_10710);
xnor U13397 (N_13397,N_12214,N_9850);
nand U13398 (N_13398,N_12353,N_12404);
nor U13399 (N_13399,N_11118,N_10139);
nand U13400 (N_13400,N_12208,N_11940);
nor U13401 (N_13401,N_11719,N_9448);
nand U13402 (N_13402,N_10477,N_12401);
or U13403 (N_13403,N_11985,N_12379);
and U13404 (N_13404,N_12228,N_12050);
and U13405 (N_13405,N_10831,N_10230);
or U13406 (N_13406,N_10958,N_9568);
nor U13407 (N_13407,N_10708,N_11686);
nand U13408 (N_13408,N_10514,N_10443);
nor U13409 (N_13409,N_10409,N_11649);
and U13410 (N_13410,N_11181,N_12291);
and U13411 (N_13411,N_10609,N_9968);
nand U13412 (N_13412,N_11365,N_11622);
and U13413 (N_13413,N_12183,N_12249);
or U13414 (N_13414,N_11624,N_12111);
or U13415 (N_13415,N_9786,N_11140);
or U13416 (N_13416,N_11319,N_12385);
nor U13417 (N_13417,N_12193,N_11325);
or U13418 (N_13418,N_12237,N_11183);
nor U13419 (N_13419,N_12325,N_10467);
and U13420 (N_13420,N_9897,N_12330);
nor U13421 (N_13421,N_11269,N_11537);
and U13422 (N_13422,N_10124,N_12457);
nor U13423 (N_13423,N_11210,N_12283);
nor U13424 (N_13424,N_10617,N_9902);
nor U13425 (N_13425,N_12266,N_10535);
or U13426 (N_13426,N_12126,N_10634);
or U13427 (N_13427,N_10152,N_10900);
or U13428 (N_13428,N_10883,N_10938);
nor U13429 (N_13429,N_9546,N_10217);
and U13430 (N_13430,N_10754,N_11145);
nor U13431 (N_13431,N_9466,N_9536);
and U13432 (N_13432,N_10212,N_9698);
nand U13433 (N_13433,N_10354,N_11354);
xnor U13434 (N_13434,N_10694,N_10891);
nand U13435 (N_13435,N_11938,N_10297);
or U13436 (N_13436,N_9815,N_9468);
nor U13437 (N_13437,N_10173,N_10414);
nand U13438 (N_13438,N_9977,N_11016);
nor U13439 (N_13439,N_10084,N_11674);
and U13440 (N_13440,N_10568,N_12064);
nor U13441 (N_13441,N_12124,N_9803);
nor U13442 (N_13442,N_12261,N_10513);
or U13443 (N_13443,N_11428,N_11196);
or U13444 (N_13444,N_10847,N_12280);
or U13445 (N_13445,N_10316,N_11762);
and U13446 (N_13446,N_9647,N_10533);
and U13447 (N_13447,N_12204,N_9627);
and U13448 (N_13448,N_10558,N_9944);
and U13449 (N_13449,N_10523,N_10846);
nand U13450 (N_13450,N_12461,N_10074);
nor U13451 (N_13451,N_11690,N_10759);
or U13452 (N_13452,N_10606,N_9766);
nand U13453 (N_13453,N_10282,N_11187);
nand U13454 (N_13454,N_9813,N_11481);
and U13455 (N_13455,N_12241,N_10138);
nand U13456 (N_13456,N_9525,N_11876);
nand U13457 (N_13457,N_9725,N_12431);
nor U13458 (N_13458,N_9761,N_12023);
or U13459 (N_13459,N_10149,N_11992);
or U13460 (N_13460,N_9537,N_11843);
nand U13461 (N_13461,N_9579,N_9593);
nor U13462 (N_13462,N_11901,N_11688);
nand U13463 (N_13463,N_11633,N_12327);
nor U13464 (N_13464,N_11150,N_10349);
and U13465 (N_13465,N_10090,N_11476);
nand U13466 (N_13466,N_11860,N_10804);
and U13467 (N_13467,N_11246,N_9385);
nand U13468 (N_13468,N_9625,N_11816);
nand U13469 (N_13469,N_10991,N_12290);
nor U13470 (N_13470,N_11536,N_10761);
or U13471 (N_13471,N_9423,N_12086);
and U13472 (N_13472,N_10283,N_11249);
nand U13473 (N_13473,N_12029,N_9722);
and U13474 (N_13474,N_10649,N_12356);
xnor U13475 (N_13475,N_10102,N_10501);
and U13476 (N_13476,N_9401,N_10596);
nor U13477 (N_13477,N_9828,N_11263);
or U13478 (N_13478,N_11848,N_10889);
nand U13479 (N_13479,N_12400,N_11806);
or U13480 (N_13480,N_12331,N_11829);
nand U13481 (N_13481,N_10319,N_12469);
xor U13482 (N_13482,N_11105,N_11006);
nand U13483 (N_13483,N_11089,N_11602);
xor U13484 (N_13484,N_12348,N_12012);
and U13485 (N_13485,N_11091,N_10663);
or U13486 (N_13486,N_11363,N_11400);
nand U13487 (N_13487,N_10169,N_10902);
nor U13488 (N_13488,N_9794,N_10038);
xor U13489 (N_13489,N_9582,N_12323);
and U13490 (N_13490,N_10296,N_9605);
xor U13491 (N_13491,N_9956,N_10311);
and U13492 (N_13492,N_11628,N_12179);
and U13493 (N_13493,N_12110,N_12095);
nor U13494 (N_13494,N_11965,N_9909);
nand U13495 (N_13495,N_9719,N_11617);
or U13496 (N_13496,N_12078,N_9526);
and U13497 (N_13497,N_11941,N_11274);
nand U13498 (N_13498,N_10129,N_9713);
nor U13499 (N_13499,N_12439,N_12279);
and U13500 (N_13500,N_12137,N_11909);
and U13501 (N_13501,N_11614,N_9797);
nand U13502 (N_13502,N_12152,N_10261);
or U13503 (N_13503,N_9375,N_9687);
nand U13504 (N_13504,N_10615,N_11474);
xnor U13505 (N_13505,N_11583,N_11462);
nor U13506 (N_13506,N_10944,N_12474);
nand U13507 (N_13507,N_11936,N_10716);
nor U13508 (N_13508,N_9993,N_10895);
nand U13509 (N_13509,N_12359,N_10903);
nor U13510 (N_13510,N_10164,N_9469);
and U13511 (N_13511,N_10028,N_12191);
or U13512 (N_13512,N_9851,N_11982);
nand U13513 (N_13513,N_12308,N_10298);
nand U13514 (N_13514,N_10171,N_9931);
or U13515 (N_13515,N_9534,N_12004);
nand U13516 (N_13516,N_11852,N_10562);
or U13517 (N_13517,N_10974,N_12128);
nand U13518 (N_13518,N_12414,N_11503);
and U13519 (N_13519,N_11182,N_10348);
nand U13520 (N_13520,N_10325,N_9758);
xor U13521 (N_13521,N_9459,N_9496);
nand U13522 (N_13522,N_10191,N_10905);
and U13523 (N_13523,N_11109,N_12175);
nor U13524 (N_13524,N_10518,N_10841);
or U13525 (N_13525,N_11141,N_9970);
nor U13526 (N_13526,N_9653,N_12021);
or U13527 (N_13527,N_9940,N_12089);
xor U13528 (N_13528,N_10061,N_11827);
and U13529 (N_13529,N_11897,N_11663);
nand U13530 (N_13530,N_10670,N_12182);
nor U13531 (N_13531,N_11557,N_9378);
and U13532 (N_13532,N_11129,N_12171);
or U13533 (N_13533,N_11790,N_11289);
nand U13534 (N_13534,N_12091,N_10959);
or U13535 (N_13535,N_10760,N_9708);
xor U13536 (N_13536,N_12170,N_12072);
or U13537 (N_13537,N_9405,N_11185);
nand U13538 (N_13538,N_10843,N_11507);
nor U13539 (N_13539,N_9900,N_11798);
and U13540 (N_13540,N_10659,N_9412);
nor U13541 (N_13541,N_11292,N_10491);
or U13542 (N_13542,N_12000,N_11525);
and U13543 (N_13543,N_11419,N_9751);
nand U13544 (N_13544,N_10714,N_9816);
and U13545 (N_13545,N_10235,N_12471);
xnor U13546 (N_13546,N_9874,N_11757);
nand U13547 (N_13547,N_9724,N_11334);
nor U13548 (N_13548,N_11172,N_11324);
nor U13549 (N_13549,N_10826,N_10023);
nand U13550 (N_13550,N_9447,N_10408);
nand U13551 (N_13551,N_11803,N_11347);
nor U13552 (N_13552,N_10797,N_11072);
nor U13553 (N_13553,N_9557,N_12013);
and U13554 (N_13554,N_10957,N_11922);
and U13555 (N_13555,N_9958,N_11741);
nand U13556 (N_13556,N_9949,N_9986);
nor U13557 (N_13557,N_10247,N_12219);
nor U13558 (N_13558,N_11209,N_11468);
or U13559 (N_13559,N_10186,N_9905);
nor U13560 (N_13560,N_12302,N_10130);
nand U13561 (N_13561,N_11444,N_11666);
nand U13562 (N_13562,N_10886,N_11374);
nor U13563 (N_13563,N_12015,N_10280);
nand U13564 (N_13564,N_9814,N_9898);
and U13565 (N_13565,N_10142,N_12256);
and U13566 (N_13566,N_11758,N_11637);
nor U13567 (N_13567,N_11207,N_10118);
or U13568 (N_13568,N_11920,N_9517);
nand U13569 (N_13569,N_12339,N_11082);
or U13570 (N_13570,N_10336,N_10305);
nor U13571 (N_13571,N_12396,N_11826);
nand U13572 (N_13572,N_11466,N_10343);
or U13573 (N_13573,N_10525,N_10010);
nand U13574 (N_13574,N_11063,N_10850);
and U13575 (N_13575,N_10899,N_9404);
and U13576 (N_13576,N_11910,N_11819);
nor U13577 (N_13577,N_9419,N_11058);
and U13578 (N_13578,N_11930,N_12166);
nand U13579 (N_13579,N_10357,N_11851);
nor U13580 (N_13580,N_9607,N_11717);
nor U13581 (N_13581,N_10728,N_11711);
or U13582 (N_13582,N_9637,N_9490);
and U13583 (N_13583,N_11445,N_9865);
nand U13584 (N_13584,N_11499,N_9478);
xor U13585 (N_13585,N_10738,N_12483);
nand U13586 (N_13586,N_11733,N_11902);
nand U13587 (N_13587,N_9926,N_10982);
nor U13588 (N_13588,N_10434,N_10195);
nor U13589 (N_13589,N_11278,N_11313);
nand U13590 (N_13590,N_9877,N_10213);
and U13591 (N_13591,N_10691,N_12106);
nor U13592 (N_13592,N_11886,N_10734);
xor U13593 (N_13593,N_9383,N_10745);
nor U13594 (N_13594,N_11792,N_11673);
xnor U13595 (N_13595,N_11813,N_10860);
and U13596 (N_13596,N_11259,N_12355);
and U13597 (N_13597,N_9591,N_11176);
nand U13598 (N_13598,N_9859,N_10112);
nand U13599 (N_13599,N_9894,N_12084);
and U13600 (N_13600,N_10442,N_11531);
and U13601 (N_13601,N_12037,N_11912);
or U13602 (N_13602,N_11234,N_10418);
nor U13603 (N_13603,N_10753,N_10224);
and U13604 (N_13604,N_12478,N_12454);
or U13605 (N_13605,N_9749,N_9908);
or U13606 (N_13606,N_10702,N_11659);
nand U13607 (N_13607,N_12016,N_10614);
or U13608 (N_13608,N_11101,N_10726);
and U13609 (N_13609,N_11048,N_10047);
nand U13610 (N_13610,N_10707,N_10553);
and U13611 (N_13611,N_10581,N_11213);
or U13612 (N_13612,N_11870,N_10403);
or U13613 (N_13613,N_11454,N_10232);
and U13614 (N_13614,N_9428,N_10428);
nand U13615 (N_13615,N_10715,N_10933);
nor U13616 (N_13616,N_11587,N_9765);
xnor U13617 (N_13617,N_10192,N_11709);
and U13618 (N_13618,N_10276,N_9762);
nor U13619 (N_13619,N_12008,N_11455);
and U13620 (N_13620,N_9489,N_9818);
nand U13621 (N_13621,N_11159,N_11953);
or U13622 (N_13622,N_12482,N_10669);
and U13623 (N_13623,N_9793,N_11031);
nand U13624 (N_13624,N_11021,N_12277);
and U13625 (N_13625,N_10611,N_10785);
and U13626 (N_13626,N_12347,N_12260);
and U13627 (N_13627,N_10145,N_9923);
nand U13628 (N_13628,N_11059,N_10219);
and U13629 (N_13629,N_11546,N_12343);
or U13630 (N_13630,N_11341,N_9617);
or U13631 (N_13631,N_9523,N_10630);
and U13632 (N_13632,N_10222,N_11923);
nand U13633 (N_13633,N_11925,N_9427);
nand U13634 (N_13634,N_10097,N_10407);
xor U13635 (N_13635,N_12103,N_9995);
nor U13636 (N_13636,N_9862,N_11464);
nor U13637 (N_13637,N_11976,N_10364);
xnor U13638 (N_13638,N_11907,N_10507);
nor U13639 (N_13639,N_10578,N_10510);
nand U13640 (N_13640,N_9556,N_10546);
and U13641 (N_13641,N_12218,N_10978);
nand U13642 (N_13642,N_12434,N_10397);
nand U13643 (N_13643,N_11708,N_12201);
nor U13644 (N_13644,N_10936,N_11229);
nor U13645 (N_13645,N_11834,N_12109);
and U13646 (N_13646,N_12438,N_11984);
nand U13647 (N_13647,N_11726,N_10346);
nor U13648 (N_13648,N_11684,N_10887);
nand U13649 (N_13649,N_10070,N_9438);
and U13650 (N_13650,N_9559,N_10713);
nor U13651 (N_13651,N_10460,N_9678);
nand U13652 (N_13652,N_10000,N_10968);
nand U13653 (N_13653,N_12147,N_9955);
nand U13654 (N_13654,N_11221,N_10969);
nand U13655 (N_13655,N_9542,N_11104);
nand U13656 (N_13656,N_9805,N_10215);
nor U13657 (N_13657,N_10527,N_11399);
nor U13658 (N_13658,N_12460,N_10503);
nand U13659 (N_13659,N_9844,N_11439);
or U13660 (N_13660,N_10166,N_11959);
nor U13661 (N_13661,N_11167,N_11383);
nor U13662 (N_13662,N_10569,N_10067);
nor U13663 (N_13663,N_11297,N_10693);
nor U13664 (N_13664,N_10265,N_9387);
and U13665 (N_13665,N_11720,N_12493);
nand U13666 (N_13666,N_11423,N_12122);
nand U13667 (N_13667,N_10633,N_10747);
and U13668 (N_13668,N_11134,N_10836);
and U13669 (N_13669,N_10950,N_11075);
or U13670 (N_13670,N_11541,N_11043);
and U13671 (N_13671,N_10012,N_10446);
nand U13672 (N_13672,N_11345,N_9553);
or U13673 (N_13673,N_11712,N_9505);
and U13674 (N_13674,N_10910,N_12267);
and U13675 (N_13675,N_10058,N_11099);
and U13676 (N_13676,N_10431,N_10796);
nor U13677 (N_13677,N_12409,N_11102);
or U13678 (N_13678,N_11779,N_11241);
xor U13679 (N_13679,N_10032,N_10401);
and U13680 (N_13680,N_12136,N_10200);
nand U13681 (N_13681,N_10667,N_12394);
xor U13682 (N_13682,N_11997,N_11840);
or U13683 (N_13683,N_9560,N_11202);
nor U13684 (N_13684,N_11509,N_12350);
xnor U13685 (N_13685,N_10109,N_12026);
nand U13686 (N_13686,N_10532,N_10436);
nand U13687 (N_13687,N_10485,N_12494);
nand U13688 (N_13688,N_12358,N_10699);
nor U13689 (N_13689,N_12238,N_9549);
nand U13690 (N_13690,N_9391,N_9554);
nor U13691 (N_13691,N_12442,N_11137);
nor U13692 (N_13692,N_11391,N_10565);
and U13693 (N_13693,N_12496,N_9717);
nand U13694 (N_13694,N_10313,N_9802);
xor U13695 (N_13695,N_11064,N_12068);
nor U13696 (N_13696,N_10626,N_12024);
or U13697 (N_13697,N_12264,N_9397);
nor U13698 (N_13698,N_12245,N_9820);
nor U13699 (N_13699,N_10574,N_10655);
nand U13700 (N_13700,N_10281,N_12486);
or U13701 (N_13701,N_12187,N_10554);
or U13702 (N_13702,N_10174,N_10091);
or U13703 (N_13703,N_9928,N_11543);
nor U13704 (N_13704,N_12281,N_10515);
nand U13705 (N_13705,N_12412,N_11913);
or U13706 (N_13706,N_11029,N_10239);
nand U13707 (N_13707,N_11780,N_9621);
nand U13708 (N_13708,N_9863,N_10907);
and U13709 (N_13709,N_10106,N_9495);
nor U13710 (N_13710,N_11974,N_9651);
nand U13711 (N_13711,N_10438,N_9421);
and U13712 (N_13712,N_11597,N_10534);
or U13713 (N_13713,N_9599,N_11995);
nand U13714 (N_13714,N_12010,N_11680);
nand U13715 (N_13715,N_11411,N_12090);
nand U13716 (N_13716,N_11204,N_12181);
or U13717 (N_13717,N_9661,N_12420);
and U13718 (N_13718,N_12148,N_12268);
xnor U13719 (N_13719,N_11220,N_11547);
and U13720 (N_13720,N_12242,N_12028);
nand U13721 (N_13721,N_9994,N_12335);
nand U13722 (N_13722,N_12146,N_9936);
nor U13723 (N_13723,N_12105,N_10932);
nor U13724 (N_13724,N_10530,N_12177);
or U13725 (N_13725,N_10495,N_11336);
and U13726 (N_13726,N_9866,N_12247);
and U13727 (N_13727,N_11050,N_11657);
nand U13728 (N_13728,N_12003,N_9668);
nor U13729 (N_13729,N_9981,N_10116);
nand U13730 (N_13730,N_9727,N_11916);
nor U13731 (N_13731,N_12252,N_9747);
nor U13732 (N_13732,N_9938,N_10229);
nand U13733 (N_13733,N_10567,N_11738);
nand U13734 (N_13734,N_9699,N_11156);
xnor U13735 (N_13735,N_11858,N_9492);
nor U13736 (N_13736,N_9443,N_10417);
xor U13737 (N_13737,N_11588,N_11562);
or U13738 (N_13738,N_9516,N_11575);
or U13739 (N_13739,N_11170,N_11889);
and U13740 (N_13740,N_11926,N_10560);
nor U13741 (N_13741,N_9919,N_12437);
nand U13742 (N_13742,N_11544,N_9954);
nand U13743 (N_13743,N_11998,N_10644);
or U13744 (N_13744,N_11871,N_11037);
xnor U13745 (N_13745,N_12223,N_11631);
nand U13746 (N_13746,N_11275,N_10610);
nand U13747 (N_13747,N_11429,N_11987);
or U13748 (N_13748,N_10805,N_11801);
nand U13749 (N_13749,N_10361,N_11253);
xor U13750 (N_13750,N_10398,N_11402);
or U13751 (N_13751,N_9736,N_10704);
nand U13752 (N_13752,N_11654,N_10939);
or U13753 (N_13753,N_9669,N_11777);
nand U13754 (N_13754,N_11705,N_11392);
nand U13755 (N_13755,N_11823,N_10248);
or U13756 (N_13756,N_9613,N_12406);
and U13757 (N_13757,N_10249,N_11661);
and U13758 (N_13758,N_10433,N_9732);
and U13759 (N_13759,N_10975,N_11356);
xor U13760 (N_13760,N_9960,N_11648);
nand U13761 (N_13761,N_10458,N_11271);
nand U13762 (N_13762,N_12293,N_10665);
nor U13763 (N_13763,N_12163,N_10114);
and U13764 (N_13764,N_10056,N_11078);
and U13765 (N_13765,N_9432,N_12018);
nor U13766 (N_13766,N_11535,N_10678);
nor U13767 (N_13767,N_10389,N_9618);
nand U13768 (N_13768,N_10099,N_10813);
nor U13769 (N_13769,N_10111,N_10151);
nand U13770 (N_13770,N_11020,N_11139);
or U13771 (N_13771,N_11986,N_10184);
nor U13772 (N_13772,N_11240,N_11112);
and U13773 (N_13773,N_12450,N_10096);
nand U13774 (N_13774,N_12224,N_11679);
or U13775 (N_13775,N_9480,N_10332);
nor U13776 (N_13776,N_9806,N_9864);
or U13777 (N_13777,N_9675,N_9912);
or U13778 (N_13778,N_11740,N_11467);
nand U13779 (N_13779,N_12197,N_12417);
nand U13780 (N_13780,N_9461,N_11681);
nand U13781 (N_13781,N_11302,N_11815);
nor U13782 (N_13782,N_10365,N_10290);
and U13783 (N_13783,N_11691,N_10459);
nor U13784 (N_13784,N_11542,N_10881);
and U13785 (N_13785,N_10952,N_11147);
nand U13786 (N_13786,N_10926,N_11695);
nand U13787 (N_13787,N_10158,N_10189);
xnor U13788 (N_13788,N_10519,N_10856);
and U13789 (N_13789,N_10575,N_10275);
nand U13790 (N_13790,N_9636,N_12292);
nor U13791 (N_13791,N_10651,N_10259);
or U13792 (N_13792,N_10388,N_10540);
nand U13793 (N_13793,N_9399,N_11312);
nor U13794 (N_13794,N_11715,N_11896);
or U13795 (N_13795,N_11382,N_10183);
nor U13796 (N_13796,N_9434,N_10790);
nor U13797 (N_13797,N_9824,N_10486);
nand U13798 (N_13798,N_11133,N_11643);
and U13799 (N_13799,N_11594,N_11360);
or U13800 (N_13800,N_9616,N_10623);
xnor U13801 (N_13801,N_9899,N_9735);
nand U13802 (N_13802,N_10604,N_11124);
or U13803 (N_13803,N_12199,N_9658);
or U13804 (N_13804,N_11121,N_9656);
nand U13805 (N_13805,N_11697,N_10029);
xnor U13806 (N_13806,N_10435,N_9776);
nand U13807 (N_13807,N_10993,N_10456);
nand U13808 (N_13808,N_11545,N_12294);
and U13809 (N_13809,N_10254,N_12092);
or U13810 (N_13810,N_12047,N_9660);
xnor U13811 (N_13811,N_10741,N_11978);
nor U13812 (N_13812,N_11500,N_10363);
and U13813 (N_13813,N_11593,N_9622);
xor U13814 (N_13814,N_12035,N_11721);
nand U13815 (N_13815,N_10127,N_10182);
nand U13816 (N_13816,N_9906,N_11483);
and U13817 (N_13817,N_11008,N_11880);
or U13818 (N_13818,N_9457,N_12346);
nand U13819 (N_13819,N_12287,N_10820);
or U13820 (N_13820,N_9508,N_10331);
or U13821 (N_13821,N_10551,N_10317);
xnor U13822 (N_13822,N_12071,N_9676);
nor U13823 (N_13823,N_9884,N_10758);
or U13824 (N_13824,N_10196,N_11248);
and U13825 (N_13825,N_11807,N_12123);
or U13826 (N_13826,N_11612,N_12468);
nand U13827 (N_13827,N_10522,N_11086);
nor U13828 (N_13828,N_10866,N_9689);
nand U13829 (N_13829,N_11646,N_10859);
nand U13830 (N_13830,N_9612,N_9539);
nand U13831 (N_13831,N_10642,N_12160);
nand U13832 (N_13832,N_10808,N_9788);
and U13833 (N_13833,N_9901,N_11389);
xor U13834 (N_13834,N_11403,N_11350);
nand U13835 (N_13835,N_12164,N_9501);
or U13836 (N_13836,N_11514,N_10243);
and U13837 (N_13837,N_10641,N_10616);
nand U13838 (N_13838,N_11802,N_12443);
xnor U13839 (N_13839,N_10880,N_11605);
xnor U13840 (N_13840,N_10862,N_11621);
xor U13841 (N_13841,N_11600,N_11584);
nand U13842 (N_13842,N_12156,N_10267);
nor U13843 (N_13843,N_10561,N_10810);
and U13844 (N_13844,N_12315,N_12354);
nor U13845 (N_13845,N_11310,N_10049);
nand U13846 (N_13846,N_10262,N_10018);
nor U13847 (N_13847,N_12334,N_10465);
nor U13848 (N_13848,N_9662,N_12117);
xor U13849 (N_13849,N_9504,N_9600);
xnor U13850 (N_13850,N_9572,N_9925);
and U13851 (N_13851,N_12098,N_9406);
xor U13852 (N_13852,N_9547,N_9394);
and U13853 (N_13853,N_12131,N_9833);
or U13854 (N_13854,N_10685,N_10419);
xor U13855 (N_13855,N_9817,N_10087);
or U13856 (N_13856,N_11534,N_11775);
xor U13857 (N_13857,N_12014,N_10315);
and U13858 (N_13858,N_10025,N_11682);
or U13859 (N_13859,N_10812,N_10572);
or U13860 (N_13860,N_11862,N_10853);
xnor U13861 (N_13861,N_9650,N_9744);
and U13862 (N_13862,N_12462,N_10475);
or U13863 (N_13863,N_11351,N_9561);
nor U13864 (N_13864,N_12258,N_10628);
or U13865 (N_13865,N_9558,N_11810);
xor U13866 (N_13866,N_11430,N_12002);
or U13867 (N_13867,N_9408,N_10768);
or U13868 (N_13868,N_12441,N_11952);
nor U13869 (N_13869,N_11591,N_11864);
or U13870 (N_13870,N_11683,N_9518);
nor U13871 (N_13871,N_10517,N_11770);
nand U13872 (N_13872,N_10972,N_11163);
nor U13873 (N_13873,N_11130,N_10333);
or U13874 (N_13874,N_9424,N_10390);
and U13875 (N_13875,N_11884,N_10453);
or U13876 (N_13876,N_11556,N_11440);
and U13877 (N_13877,N_9389,N_11765);
or U13878 (N_13878,N_10128,N_9564);
or U13879 (N_13879,N_12051,N_11931);
and U13880 (N_13880,N_9939,N_9510);
and U13881 (N_13881,N_12009,N_11730);
nand U13882 (N_13882,N_11005,N_11565);
and U13883 (N_13883,N_12369,N_10879);
or U13884 (N_13884,N_9619,N_12115);
xor U13885 (N_13885,N_12229,N_11595);
nor U13886 (N_13886,N_10584,N_10412);
xor U13887 (N_13887,N_10844,N_10643);
xnor U13888 (N_13888,N_12093,N_9376);
or U13889 (N_13889,N_12352,N_9989);
nor U13890 (N_13890,N_11406,N_11566);
nand U13891 (N_13891,N_11748,N_10473);
xnor U13892 (N_13892,N_11879,N_11390);
and U13893 (N_13893,N_11582,N_11346);
or U13894 (N_13894,N_11652,N_11818);
nand U13895 (N_13895,N_10123,N_9896);
and U13896 (N_13896,N_12096,N_11553);
nand U13897 (N_13897,N_9624,N_12100);
and U13898 (N_13898,N_11254,N_11178);
nand U13899 (N_13899,N_11025,N_12426);
or U13900 (N_13900,N_10712,N_11366);
xnor U13901 (N_13901,N_12390,N_12435);
xor U13902 (N_13902,N_11266,N_12399);
nand U13903 (N_13903,N_11517,N_9674);
or U13904 (N_13904,N_10429,N_10740);
nand U13905 (N_13905,N_10344,N_11983);
or U13906 (N_13906,N_10603,N_9840);
or U13907 (N_13907,N_10273,N_10323);
and U13908 (N_13908,N_10698,N_10686);
nor U13909 (N_13909,N_9464,N_9942);
nor U13910 (N_13910,N_11662,N_9819);
or U13911 (N_13911,N_9714,N_10009);
or U13912 (N_13912,N_10770,N_11352);
and U13913 (N_13913,N_12067,N_10730);
nor U13914 (N_13914,N_11824,N_12209);
or U13915 (N_13915,N_11532,N_10207);
nor U13916 (N_13916,N_10800,N_10834);
xnor U13917 (N_13917,N_10526,N_11003);
or U13918 (N_13918,N_10252,N_11498);
and U13919 (N_13919,N_11865,N_10544);
nor U13920 (N_13920,N_10666,N_9629);
nor U13921 (N_13921,N_12386,N_12054);
or U13922 (N_13922,N_11999,N_11616);
nand U13923 (N_13923,N_9729,N_10629);
nor U13924 (N_13924,N_10987,N_12470);
xor U13925 (N_13925,N_11304,N_10566);
xnor U13926 (N_13926,N_12449,N_10062);
and U13927 (N_13927,N_9578,N_10771);
nand U13928 (N_13928,N_11018,N_9550);
nand U13929 (N_13929,N_11844,N_9867);
nand U13930 (N_13930,N_11223,N_12436);
nand U13931 (N_13931,N_11237,N_11786);
nand U13932 (N_13932,N_11598,N_12139);
or U13933 (N_13933,N_12333,N_11863);
nor U13934 (N_13934,N_11243,N_10066);
and U13935 (N_13935,N_11988,N_11504);
nand U13936 (N_13936,N_12395,N_10185);
nor U13937 (N_13937,N_10992,N_12472);
nor U13938 (N_13938,N_11216,N_9924);
nand U13939 (N_13939,N_9515,N_10303);
xor U13940 (N_13940,N_10998,N_9382);
xor U13941 (N_13941,N_10701,N_10444);
and U13942 (N_13942,N_9767,N_12383);
nand U13943 (N_13943,N_10739,N_9885);
xnor U13944 (N_13944,N_9552,N_9514);
or U13945 (N_13945,N_10258,N_11194);
or U13946 (N_13946,N_12338,N_10552);
or U13947 (N_13947,N_10543,N_12020);
xnor U13948 (N_13948,N_11518,N_11256);
nand U13949 (N_13949,N_11437,N_11776);
xnor U13950 (N_13950,N_9409,N_10995);
and U13951 (N_13951,N_10688,N_11656);
nand U13952 (N_13952,N_9666,N_9563);
or U13953 (N_13953,N_10852,N_9430);
and U13954 (N_13954,N_11151,N_11268);
nand U13955 (N_13955,N_10304,N_11703);
or U13956 (N_13956,N_12150,N_9982);
and U13957 (N_13957,N_10587,N_10725);
and U13958 (N_13958,N_9436,N_10935);
nor U13959 (N_13959,N_10352,N_9943);
or U13960 (N_13960,N_9875,N_9395);
xnor U13961 (N_13961,N_9551,N_11768);
nand U13962 (N_13962,N_11970,N_11782);
nor U13963 (N_13963,N_11487,N_11728);
and U13964 (N_13964,N_10216,N_11548);
xor U13965 (N_13965,N_10816,N_9630);
nand U13966 (N_13966,N_10266,N_12141);
or U13967 (N_13967,N_11571,N_10825);
nand U13968 (N_13968,N_11067,N_12055);
and U13969 (N_13969,N_12243,N_9778);
and U13970 (N_13970,N_11144,N_12411);
nor U13971 (N_13971,N_11311,N_11601);
nor U13972 (N_13972,N_12188,N_11041);
nand U13973 (N_13973,N_10668,N_9456);
and U13974 (N_13974,N_11956,N_10043);
nand U13975 (N_13975,N_10988,N_11153);
nor U13976 (N_13976,N_11630,N_11919);
nand U13977 (N_13977,N_11743,N_10622);
and U13978 (N_13978,N_12161,N_9454);
and U13979 (N_13979,N_10065,N_9832);
or U13980 (N_13980,N_10464,N_10756);
nor U13981 (N_13981,N_11763,N_10199);
nor U13982 (N_13982,N_10274,N_10613);
or U13983 (N_13983,N_9798,N_12497);
and U13984 (N_13984,N_11971,N_11501);
nor U13985 (N_13985,N_11398,N_11022);
or U13986 (N_13986,N_11994,N_9997);
and U13987 (N_13987,N_11148,N_10463);
nand U13988 (N_13988,N_11049,N_11618);
and U13989 (N_13989,N_10479,N_12446);
xnor U13990 (N_13990,N_10462,N_12378);
and U13991 (N_13991,N_9416,N_10162);
nor U13992 (N_13992,N_12452,N_11672);
nor U13993 (N_13993,N_11623,N_12489);
or U13994 (N_13994,N_10338,N_11996);
nand U13995 (N_13995,N_11418,N_12365);
or U13996 (N_13996,N_10197,N_10940);
or U13997 (N_13997,N_10140,N_11538);
nand U13998 (N_13998,N_10069,N_10985);
and U13999 (N_13999,N_11108,N_10263);
nand U14000 (N_14000,N_11111,N_11642);
or U14001 (N_14001,N_9754,N_10537);
and U14002 (N_14002,N_11171,N_10870);
nor U14003 (N_14003,N_11092,N_9410);
nor U14004 (N_14004,N_11070,N_12101);
or U14005 (N_14005,N_10915,N_9792);
xor U14006 (N_14006,N_10472,N_12017);
nand U14007 (N_14007,N_12314,N_9548);
and U14008 (N_14008,N_9576,N_11853);
or U14009 (N_14009,N_10878,N_10994);
nor U14010 (N_14010,N_11427,N_11484);
nor U14011 (N_14011,N_10342,N_11972);
nor U14012 (N_14012,N_10815,N_10882);
nand U14013 (N_14013,N_11103,N_12153);
or U14014 (N_14014,N_10270,N_10466);
and U14015 (N_14015,N_12380,N_11555);
or U14016 (N_14016,N_11377,N_9535);
xnor U14017 (N_14017,N_10833,N_9834);
or U14018 (N_14018,N_10170,N_11214);
and U14019 (N_14019,N_10001,N_12430);
nand U14020 (N_14020,N_12481,N_11180);
nor U14021 (N_14021,N_12313,N_9913);
and U14022 (N_14022,N_12427,N_10656);
and U14023 (N_14023,N_11087,N_10309);
and U14024 (N_14024,N_12317,N_9633);
nand U14025 (N_14025,N_10041,N_11042);
nor U14026 (N_14026,N_9974,N_12070);
nand U14027 (N_14027,N_12341,N_10849);
nor U14028 (N_14028,N_10788,N_11371);
and U14029 (N_14029,N_11284,N_11322);
and U14030 (N_14030,N_11781,N_10052);
nand U14031 (N_14031,N_9470,N_10367);
or U14032 (N_14032,N_9987,N_10732);
or U14033 (N_14033,N_9962,N_10824);
nand U14034 (N_14034,N_10157,N_12088);
nand U14035 (N_14035,N_11990,N_10986);
and U14036 (N_14036,N_10251,N_12011);
and U14037 (N_14037,N_9413,N_9892);
nand U14038 (N_14038,N_9381,N_10117);
xor U14039 (N_14039,N_9414,N_12324);
nor U14040 (N_14040,N_10150,N_11397);
and U14041 (N_14041,N_12042,N_10999);
nand U14042 (N_14042,N_12284,N_12336);
and U14043 (N_14043,N_11226,N_12492);
nor U14044 (N_14044,N_10914,N_9731);
nand U14045 (N_14045,N_9696,N_11494);
and U14046 (N_14046,N_11857,N_12030);
or U14047 (N_14047,N_10700,N_12476);
nor U14048 (N_14048,N_12366,N_12285);
and U14049 (N_14049,N_11849,N_11607);
nor U14050 (N_14050,N_11960,N_10855);
and U14051 (N_14051,N_10602,N_10402);
and U14052 (N_14052,N_9969,N_10624);
nand U14053 (N_14053,N_9967,N_12418);
or U14054 (N_14054,N_12215,N_9472);
nand U14055 (N_14055,N_11293,N_11898);
nand U14056 (N_14056,N_10327,N_10178);
nand U14057 (N_14057,N_10897,N_12107);
xnor U14058 (N_14058,N_9575,N_9948);
nor U14059 (N_14059,N_9683,N_11955);
xnor U14060 (N_14060,N_9920,N_9686);
nand U14061 (N_14061,N_11475,N_11783);
nor U14062 (N_14062,N_10779,N_10654);
or U14063 (N_14063,N_10711,N_10336);
nand U14064 (N_14064,N_11703,N_12007);
nor U14065 (N_14065,N_10267,N_12445);
nand U14066 (N_14066,N_12257,N_10509);
nor U14067 (N_14067,N_11489,N_11039);
nor U14068 (N_14068,N_11677,N_10200);
nand U14069 (N_14069,N_10310,N_10869);
nor U14070 (N_14070,N_10532,N_11332);
or U14071 (N_14071,N_11066,N_11263);
or U14072 (N_14072,N_11591,N_10901);
nor U14073 (N_14073,N_11510,N_9451);
and U14074 (N_14074,N_10421,N_9426);
or U14075 (N_14075,N_10559,N_11008);
nand U14076 (N_14076,N_9750,N_12132);
nand U14077 (N_14077,N_10477,N_11776);
and U14078 (N_14078,N_11820,N_10920);
or U14079 (N_14079,N_11970,N_9691);
or U14080 (N_14080,N_10784,N_10292);
nand U14081 (N_14081,N_11611,N_11229);
nand U14082 (N_14082,N_10395,N_11087);
nor U14083 (N_14083,N_9543,N_12454);
or U14084 (N_14084,N_12483,N_10758);
nor U14085 (N_14085,N_10921,N_11020);
or U14086 (N_14086,N_10980,N_12188);
xor U14087 (N_14087,N_10560,N_10734);
or U14088 (N_14088,N_10556,N_10160);
nand U14089 (N_14089,N_11140,N_10312);
or U14090 (N_14090,N_9607,N_10930);
nand U14091 (N_14091,N_10576,N_11436);
nor U14092 (N_14092,N_10956,N_12390);
xor U14093 (N_14093,N_11106,N_12369);
nand U14094 (N_14094,N_10237,N_10924);
and U14095 (N_14095,N_9818,N_9940);
nor U14096 (N_14096,N_11370,N_9620);
and U14097 (N_14097,N_12373,N_12250);
nor U14098 (N_14098,N_9538,N_11641);
nor U14099 (N_14099,N_10319,N_10164);
and U14100 (N_14100,N_12372,N_12238);
or U14101 (N_14101,N_12459,N_11359);
nand U14102 (N_14102,N_9679,N_9579);
and U14103 (N_14103,N_11419,N_10344);
nand U14104 (N_14104,N_10512,N_9674);
xor U14105 (N_14105,N_9818,N_11950);
and U14106 (N_14106,N_12342,N_10895);
or U14107 (N_14107,N_9996,N_12199);
xor U14108 (N_14108,N_10476,N_11725);
nor U14109 (N_14109,N_12216,N_9927);
nor U14110 (N_14110,N_11609,N_11988);
nand U14111 (N_14111,N_10331,N_10685);
nand U14112 (N_14112,N_11324,N_12135);
nor U14113 (N_14113,N_11840,N_11014);
nand U14114 (N_14114,N_10649,N_9451);
or U14115 (N_14115,N_11242,N_11138);
or U14116 (N_14116,N_10115,N_10130);
and U14117 (N_14117,N_10694,N_11653);
and U14118 (N_14118,N_11014,N_10130);
nand U14119 (N_14119,N_10930,N_11667);
and U14120 (N_14120,N_10161,N_10155);
or U14121 (N_14121,N_10118,N_11620);
xnor U14122 (N_14122,N_10550,N_9387);
nor U14123 (N_14123,N_9482,N_12336);
or U14124 (N_14124,N_9659,N_10967);
or U14125 (N_14125,N_10241,N_10757);
nand U14126 (N_14126,N_9454,N_11798);
or U14127 (N_14127,N_11295,N_11334);
nand U14128 (N_14128,N_10337,N_10825);
nor U14129 (N_14129,N_10468,N_11686);
nor U14130 (N_14130,N_12122,N_11641);
xnor U14131 (N_14131,N_10877,N_10467);
nor U14132 (N_14132,N_11989,N_10923);
and U14133 (N_14133,N_11348,N_10231);
and U14134 (N_14134,N_11045,N_12096);
nand U14135 (N_14135,N_12156,N_9923);
and U14136 (N_14136,N_10801,N_9800);
or U14137 (N_14137,N_10453,N_10005);
and U14138 (N_14138,N_12158,N_10899);
nand U14139 (N_14139,N_10304,N_9887);
or U14140 (N_14140,N_11951,N_11601);
xor U14141 (N_14141,N_10577,N_11887);
or U14142 (N_14142,N_10925,N_10228);
and U14143 (N_14143,N_9581,N_10907);
and U14144 (N_14144,N_11208,N_10529);
nand U14145 (N_14145,N_11275,N_10156);
and U14146 (N_14146,N_9912,N_11636);
or U14147 (N_14147,N_10760,N_11522);
and U14148 (N_14148,N_11351,N_9854);
nand U14149 (N_14149,N_9563,N_10392);
or U14150 (N_14150,N_9815,N_9576);
or U14151 (N_14151,N_10032,N_11863);
nand U14152 (N_14152,N_10902,N_10278);
nor U14153 (N_14153,N_12432,N_10607);
nor U14154 (N_14154,N_11902,N_11790);
nor U14155 (N_14155,N_10982,N_11705);
nand U14156 (N_14156,N_12035,N_10675);
nor U14157 (N_14157,N_9814,N_12104);
or U14158 (N_14158,N_10733,N_11716);
or U14159 (N_14159,N_12197,N_12471);
or U14160 (N_14160,N_10062,N_10225);
or U14161 (N_14161,N_11966,N_11010);
or U14162 (N_14162,N_11563,N_10248);
and U14163 (N_14163,N_9383,N_9553);
nor U14164 (N_14164,N_9618,N_11036);
or U14165 (N_14165,N_11730,N_9956);
nand U14166 (N_14166,N_10778,N_12321);
nor U14167 (N_14167,N_11930,N_12297);
or U14168 (N_14168,N_10937,N_9570);
xnor U14169 (N_14169,N_9918,N_10875);
and U14170 (N_14170,N_10956,N_12160);
nand U14171 (N_14171,N_10532,N_11629);
nand U14172 (N_14172,N_12181,N_11491);
nor U14173 (N_14173,N_11885,N_11041);
nand U14174 (N_14174,N_10102,N_11339);
or U14175 (N_14175,N_9458,N_9968);
nand U14176 (N_14176,N_11514,N_10026);
and U14177 (N_14177,N_9567,N_11855);
nor U14178 (N_14178,N_10934,N_9689);
nor U14179 (N_14179,N_11541,N_9385);
or U14180 (N_14180,N_12127,N_9577);
xor U14181 (N_14181,N_11307,N_10547);
xnor U14182 (N_14182,N_10151,N_11115);
nand U14183 (N_14183,N_10576,N_11079);
nand U14184 (N_14184,N_9865,N_10032);
and U14185 (N_14185,N_11631,N_11465);
nor U14186 (N_14186,N_12357,N_9420);
nor U14187 (N_14187,N_11989,N_10118);
nor U14188 (N_14188,N_10239,N_10785);
nor U14189 (N_14189,N_9709,N_12390);
and U14190 (N_14190,N_11825,N_12107);
nand U14191 (N_14191,N_10246,N_11957);
nand U14192 (N_14192,N_11911,N_9394);
nor U14193 (N_14193,N_9991,N_10495);
or U14194 (N_14194,N_10865,N_9468);
nand U14195 (N_14195,N_11443,N_11095);
or U14196 (N_14196,N_11494,N_9512);
or U14197 (N_14197,N_12487,N_11031);
xnor U14198 (N_14198,N_11327,N_11590);
or U14199 (N_14199,N_11097,N_11353);
and U14200 (N_14200,N_11036,N_12133);
or U14201 (N_14201,N_12094,N_11175);
and U14202 (N_14202,N_12066,N_10056);
nor U14203 (N_14203,N_9530,N_11306);
xor U14204 (N_14204,N_9929,N_11258);
nand U14205 (N_14205,N_10075,N_9714);
nor U14206 (N_14206,N_10299,N_11347);
nor U14207 (N_14207,N_11258,N_10825);
and U14208 (N_14208,N_10018,N_10404);
or U14209 (N_14209,N_10721,N_12226);
or U14210 (N_14210,N_11077,N_11586);
or U14211 (N_14211,N_11355,N_11526);
and U14212 (N_14212,N_10768,N_12228);
nand U14213 (N_14213,N_11679,N_9968);
or U14214 (N_14214,N_11184,N_11913);
nand U14215 (N_14215,N_11035,N_11736);
nand U14216 (N_14216,N_11422,N_12327);
nor U14217 (N_14217,N_11442,N_11573);
xnor U14218 (N_14218,N_12472,N_10339);
nor U14219 (N_14219,N_11151,N_11728);
and U14220 (N_14220,N_10496,N_11713);
nand U14221 (N_14221,N_11427,N_12463);
xor U14222 (N_14222,N_10798,N_12441);
nand U14223 (N_14223,N_9396,N_9872);
or U14224 (N_14224,N_12300,N_12062);
nor U14225 (N_14225,N_9772,N_12316);
and U14226 (N_14226,N_11147,N_10145);
and U14227 (N_14227,N_11941,N_9884);
and U14228 (N_14228,N_11630,N_10020);
nor U14229 (N_14229,N_10407,N_10674);
and U14230 (N_14230,N_9544,N_12483);
nor U14231 (N_14231,N_12233,N_10913);
nor U14232 (N_14232,N_10328,N_11509);
nand U14233 (N_14233,N_9448,N_10699);
nor U14234 (N_14234,N_10811,N_10477);
and U14235 (N_14235,N_9643,N_11457);
nor U14236 (N_14236,N_9762,N_10529);
nor U14237 (N_14237,N_11300,N_11872);
nor U14238 (N_14238,N_10253,N_11266);
or U14239 (N_14239,N_11772,N_9884);
nor U14240 (N_14240,N_11513,N_10610);
or U14241 (N_14241,N_10397,N_10380);
xor U14242 (N_14242,N_10515,N_10292);
and U14243 (N_14243,N_11004,N_12139);
nand U14244 (N_14244,N_10219,N_11318);
or U14245 (N_14245,N_12194,N_11451);
and U14246 (N_14246,N_11426,N_12242);
nor U14247 (N_14247,N_12402,N_11960);
xor U14248 (N_14248,N_11156,N_10269);
nor U14249 (N_14249,N_11494,N_9559);
nor U14250 (N_14250,N_12210,N_11967);
nand U14251 (N_14251,N_10232,N_12416);
and U14252 (N_14252,N_10343,N_11627);
xor U14253 (N_14253,N_10827,N_12332);
nor U14254 (N_14254,N_9469,N_10106);
or U14255 (N_14255,N_10576,N_11269);
nand U14256 (N_14256,N_12446,N_11688);
or U14257 (N_14257,N_11488,N_11609);
nor U14258 (N_14258,N_11632,N_11106);
and U14259 (N_14259,N_10197,N_9469);
and U14260 (N_14260,N_9901,N_11044);
xnor U14261 (N_14261,N_10555,N_10281);
nand U14262 (N_14262,N_10115,N_11537);
xnor U14263 (N_14263,N_10619,N_10066);
or U14264 (N_14264,N_9669,N_9908);
nand U14265 (N_14265,N_10005,N_10266);
xor U14266 (N_14266,N_10453,N_10067);
nand U14267 (N_14267,N_9862,N_10322);
or U14268 (N_14268,N_9412,N_11456);
nor U14269 (N_14269,N_12333,N_10781);
nor U14270 (N_14270,N_11786,N_10492);
nand U14271 (N_14271,N_11806,N_10975);
and U14272 (N_14272,N_10643,N_9665);
and U14273 (N_14273,N_10459,N_11828);
nor U14274 (N_14274,N_9403,N_9471);
nand U14275 (N_14275,N_12060,N_12477);
nand U14276 (N_14276,N_10414,N_11117);
nand U14277 (N_14277,N_10533,N_9388);
or U14278 (N_14278,N_12339,N_11776);
nor U14279 (N_14279,N_12348,N_12136);
xnor U14280 (N_14280,N_11666,N_10115);
or U14281 (N_14281,N_9989,N_10662);
or U14282 (N_14282,N_9938,N_12389);
nor U14283 (N_14283,N_10870,N_11115);
and U14284 (N_14284,N_11866,N_10992);
nand U14285 (N_14285,N_11117,N_10643);
or U14286 (N_14286,N_12407,N_11857);
nor U14287 (N_14287,N_10852,N_10813);
and U14288 (N_14288,N_11163,N_10120);
nand U14289 (N_14289,N_11060,N_11291);
xnor U14290 (N_14290,N_11315,N_11872);
xnor U14291 (N_14291,N_11999,N_10356);
nor U14292 (N_14292,N_11959,N_11132);
or U14293 (N_14293,N_11306,N_9509);
and U14294 (N_14294,N_12423,N_12498);
and U14295 (N_14295,N_9933,N_11902);
and U14296 (N_14296,N_10468,N_11541);
nor U14297 (N_14297,N_10268,N_10259);
or U14298 (N_14298,N_11700,N_12415);
nand U14299 (N_14299,N_11494,N_9926);
and U14300 (N_14300,N_11186,N_9690);
xnor U14301 (N_14301,N_10467,N_10517);
nand U14302 (N_14302,N_10053,N_10610);
and U14303 (N_14303,N_12347,N_10928);
nor U14304 (N_14304,N_11563,N_10270);
nand U14305 (N_14305,N_11830,N_10518);
nor U14306 (N_14306,N_10907,N_11597);
or U14307 (N_14307,N_10353,N_9821);
nand U14308 (N_14308,N_11877,N_9498);
and U14309 (N_14309,N_9466,N_11677);
xnor U14310 (N_14310,N_9930,N_11372);
nand U14311 (N_14311,N_11035,N_11000);
and U14312 (N_14312,N_12259,N_11522);
nand U14313 (N_14313,N_9727,N_12279);
nand U14314 (N_14314,N_10987,N_10535);
and U14315 (N_14315,N_12094,N_12336);
xor U14316 (N_14316,N_11968,N_10146);
nor U14317 (N_14317,N_11292,N_11331);
nand U14318 (N_14318,N_11044,N_9756);
nand U14319 (N_14319,N_11471,N_10556);
and U14320 (N_14320,N_9936,N_10847);
nand U14321 (N_14321,N_10485,N_11799);
or U14322 (N_14322,N_9678,N_10711);
nor U14323 (N_14323,N_10392,N_12020);
or U14324 (N_14324,N_12214,N_12125);
nand U14325 (N_14325,N_9929,N_10041);
nand U14326 (N_14326,N_10867,N_12312);
nor U14327 (N_14327,N_12245,N_12145);
xor U14328 (N_14328,N_10004,N_11890);
or U14329 (N_14329,N_10922,N_10587);
or U14330 (N_14330,N_10752,N_9552);
and U14331 (N_14331,N_9808,N_12271);
xor U14332 (N_14332,N_12436,N_11254);
nor U14333 (N_14333,N_9922,N_10934);
and U14334 (N_14334,N_11620,N_10394);
or U14335 (N_14335,N_12334,N_11668);
or U14336 (N_14336,N_11840,N_12301);
or U14337 (N_14337,N_12048,N_12154);
and U14338 (N_14338,N_10893,N_9660);
and U14339 (N_14339,N_11069,N_9988);
or U14340 (N_14340,N_9380,N_9918);
nand U14341 (N_14341,N_12461,N_10200);
nor U14342 (N_14342,N_12450,N_10016);
nor U14343 (N_14343,N_10944,N_11161);
nand U14344 (N_14344,N_12154,N_9492);
or U14345 (N_14345,N_10222,N_11738);
xnor U14346 (N_14346,N_11606,N_11168);
and U14347 (N_14347,N_10347,N_12477);
nor U14348 (N_14348,N_9605,N_12083);
or U14349 (N_14349,N_11662,N_12342);
and U14350 (N_14350,N_10667,N_12479);
nor U14351 (N_14351,N_9769,N_11200);
and U14352 (N_14352,N_9596,N_10835);
nor U14353 (N_14353,N_9863,N_12299);
or U14354 (N_14354,N_10194,N_10532);
or U14355 (N_14355,N_10092,N_9403);
xnor U14356 (N_14356,N_10964,N_10638);
and U14357 (N_14357,N_11085,N_10956);
and U14358 (N_14358,N_9475,N_9685);
or U14359 (N_14359,N_9839,N_10764);
xor U14360 (N_14360,N_10370,N_11688);
nor U14361 (N_14361,N_11711,N_12252);
nand U14362 (N_14362,N_10340,N_10508);
nand U14363 (N_14363,N_10290,N_10962);
nor U14364 (N_14364,N_12453,N_10968);
or U14365 (N_14365,N_9533,N_11534);
or U14366 (N_14366,N_11084,N_9676);
and U14367 (N_14367,N_10754,N_9705);
nand U14368 (N_14368,N_9598,N_11798);
or U14369 (N_14369,N_12225,N_10335);
or U14370 (N_14370,N_10171,N_10766);
or U14371 (N_14371,N_11132,N_9986);
and U14372 (N_14372,N_11389,N_9407);
and U14373 (N_14373,N_10206,N_10844);
and U14374 (N_14374,N_12231,N_10676);
or U14375 (N_14375,N_12233,N_10755);
or U14376 (N_14376,N_11430,N_10761);
nor U14377 (N_14377,N_12421,N_11412);
or U14378 (N_14378,N_9693,N_11983);
xnor U14379 (N_14379,N_11748,N_10534);
or U14380 (N_14380,N_11326,N_11178);
or U14381 (N_14381,N_11661,N_9841);
or U14382 (N_14382,N_11059,N_12263);
nor U14383 (N_14383,N_10658,N_10117);
or U14384 (N_14384,N_9728,N_9751);
and U14385 (N_14385,N_10512,N_10417);
nor U14386 (N_14386,N_9431,N_11924);
nor U14387 (N_14387,N_10655,N_11204);
nor U14388 (N_14388,N_11982,N_11878);
or U14389 (N_14389,N_10529,N_11639);
nand U14390 (N_14390,N_9957,N_9486);
nor U14391 (N_14391,N_10896,N_12393);
nand U14392 (N_14392,N_11600,N_10595);
nor U14393 (N_14393,N_11391,N_12230);
and U14394 (N_14394,N_9957,N_12491);
and U14395 (N_14395,N_10522,N_10422);
and U14396 (N_14396,N_11825,N_10867);
xnor U14397 (N_14397,N_10581,N_12460);
nor U14398 (N_14398,N_11367,N_10776);
or U14399 (N_14399,N_10610,N_10148);
nand U14400 (N_14400,N_11329,N_12370);
nand U14401 (N_14401,N_11416,N_11868);
nand U14402 (N_14402,N_11600,N_11217);
nand U14403 (N_14403,N_11510,N_9463);
and U14404 (N_14404,N_10835,N_10256);
or U14405 (N_14405,N_12134,N_9387);
or U14406 (N_14406,N_10423,N_9491);
and U14407 (N_14407,N_11450,N_9949);
nor U14408 (N_14408,N_11948,N_12194);
nand U14409 (N_14409,N_11310,N_11746);
and U14410 (N_14410,N_11007,N_10143);
or U14411 (N_14411,N_9590,N_9676);
and U14412 (N_14412,N_10438,N_10492);
nand U14413 (N_14413,N_10896,N_12198);
nand U14414 (N_14414,N_10426,N_11963);
nor U14415 (N_14415,N_11168,N_11239);
and U14416 (N_14416,N_11457,N_10635);
nand U14417 (N_14417,N_10457,N_11605);
nor U14418 (N_14418,N_11488,N_10388);
xnor U14419 (N_14419,N_10630,N_10542);
and U14420 (N_14420,N_11347,N_9597);
nor U14421 (N_14421,N_11364,N_10307);
and U14422 (N_14422,N_11867,N_11426);
and U14423 (N_14423,N_10616,N_12292);
nand U14424 (N_14424,N_9800,N_12268);
nor U14425 (N_14425,N_10006,N_11962);
xnor U14426 (N_14426,N_9880,N_9858);
and U14427 (N_14427,N_10496,N_12341);
or U14428 (N_14428,N_11016,N_10487);
and U14429 (N_14429,N_11123,N_12231);
nand U14430 (N_14430,N_9686,N_12027);
or U14431 (N_14431,N_9846,N_11303);
nand U14432 (N_14432,N_10078,N_10666);
nor U14433 (N_14433,N_10716,N_10996);
nor U14434 (N_14434,N_12499,N_11968);
xnor U14435 (N_14435,N_12411,N_11131);
and U14436 (N_14436,N_10051,N_11136);
nand U14437 (N_14437,N_11745,N_12209);
and U14438 (N_14438,N_11285,N_11528);
nand U14439 (N_14439,N_11653,N_9925);
or U14440 (N_14440,N_9928,N_10176);
nand U14441 (N_14441,N_11271,N_10673);
nor U14442 (N_14442,N_10263,N_11039);
and U14443 (N_14443,N_9468,N_11342);
or U14444 (N_14444,N_11964,N_10743);
or U14445 (N_14445,N_11170,N_11950);
nand U14446 (N_14446,N_10343,N_10266);
or U14447 (N_14447,N_11429,N_10901);
nor U14448 (N_14448,N_9522,N_9609);
and U14449 (N_14449,N_11904,N_10217);
or U14450 (N_14450,N_12148,N_9680);
or U14451 (N_14451,N_10007,N_9915);
and U14452 (N_14452,N_9493,N_11501);
nand U14453 (N_14453,N_11777,N_9471);
and U14454 (N_14454,N_11679,N_9869);
xor U14455 (N_14455,N_9951,N_11461);
nor U14456 (N_14456,N_12479,N_11594);
nor U14457 (N_14457,N_9654,N_10337);
xnor U14458 (N_14458,N_11159,N_12113);
nand U14459 (N_14459,N_12488,N_11362);
nand U14460 (N_14460,N_11124,N_12139);
and U14461 (N_14461,N_11217,N_11362);
and U14462 (N_14462,N_11919,N_11921);
or U14463 (N_14463,N_9513,N_11009);
nor U14464 (N_14464,N_11280,N_11435);
xor U14465 (N_14465,N_12048,N_11326);
and U14466 (N_14466,N_12184,N_11002);
nor U14467 (N_14467,N_10639,N_12248);
xnor U14468 (N_14468,N_10582,N_11312);
or U14469 (N_14469,N_9668,N_10672);
and U14470 (N_14470,N_10957,N_12348);
xnor U14471 (N_14471,N_12013,N_10734);
or U14472 (N_14472,N_10669,N_9884);
xor U14473 (N_14473,N_9376,N_11088);
or U14474 (N_14474,N_11316,N_11462);
or U14475 (N_14475,N_10399,N_10671);
and U14476 (N_14476,N_12236,N_10952);
nand U14477 (N_14477,N_11392,N_11473);
nand U14478 (N_14478,N_11186,N_11652);
xnor U14479 (N_14479,N_10485,N_11488);
nand U14480 (N_14480,N_11845,N_11537);
or U14481 (N_14481,N_9477,N_11437);
xnor U14482 (N_14482,N_12400,N_12296);
or U14483 (N_14483,N_9810,N_10146);
nor U14484 (N_14484,N_10504,N_10891);
nand U14485 (N_14485,N_10126,N_10614);
and U14486 (N_14486,N_11759,N_12379);
nor U14487 (N_14487,N_11137,N_12244);
nor U14488 (N_14488,N_10499,N_11719);
or U14489 (N_14489,N_12114,N_11722);
nand U14490 (N_14490,N_11929,N_9755);
nand U14491 (N_14491,N_12296,N_12317);
and U14492 (N_14492,N_11070,N_10928);
and U14493 (N_14493,N_11928,N_10634);
nand U14494 (N_14494,N_9393,N_9446);
xnor U14495 (N_14495,N_12487,N_10326);
and U14496 (N_14496,N_9853,N_9959);
or U14497 (N_14497,N_11567,N_12492);
nand U14498 (N_14498,N_10639,N_11335);
and U14499 (N_14499,N_11357,N_9875);
or U14500 (N_14500,N_12154,N_12316);
nand U14501 (N_14501,N_11259,N_12468);
nand U14502 (N_14502,N_10218,N_12011);
nor U14503 (N_14503,N_11559,N_11175);
or U14504 (N_14504,N_10076,N_10041);
and U14505 (N_14505,N_9903,N_10391);
or U14506 (N_14506,N_9701,N_11841);
nor U14507 (N_14507,N_12270,N_9738);
or U14508 (N_14508,N_9471,N_10520);
nand U14509 (N_14509,N_12029,N_10009);
nor U14510 (N_14510,N_11541,N_11808);
nor U14511 (N_14511,N_11777,N_12093);
nor U14512 (N_14512,N_11992,N_9450);
nor U14513 (N_14513,N_12196,N_10773);
nor U14514 (N_14514,N_11475,N_12323);
nand U14515 (N_14515,N_11536,N_10383);
nand U14516 (N_14516,N_9557,N_11436);
and U14517 (N_14517,N_10361,N_9505);
and U14518 (N_14518,N_12124,N_11755);
and U14519 (N_14519,N_9444,N_11746);
nand U14520 (N_14520,N_12454,N_11073);
or U14521 (N_14521,N_11791,N_12121);
or U14522 (N_14522,N_11659,N_12481);
and U14523 (N_14523,N_11860,N_11333);
nor U14524 (N_14524,N_11110,N_12383);
nand U14525 (N_14525,N_12185,N_11028);
nor U14526 (N_14526,N_10706,N_9541);
nand U14527 (N_14527,N_11711,N_9520);
and U14528 (N_14528,N_10283,N_10248);
xnor U14529 (N_14529,N_12031,N_9893);
and U14530 (N_14530,N_10858,N_12321);
nor U14531 (N_14531,N_9900,N_12376);
and U14532 (N_14532,N_11360,N_11236);
nor U14533 (N_14533,N_11073,N_12199);
and U14534 (N_14534,N_10176,N_11735);
nand U14535 (N_14535,N_10606,N_11091);
or U14536 (N_14536,N_10499,N_10439);
or U14537 (N_14537,N_12133,N_9564);
or U14538 (N_14538,N_12447,N_11961);
nand U14539 (N_14539,N_11644,N_10491);
or U14540 (N_14540,N_10762,N_9400);
nand U14541 (N_14541,N_9624,N_10284);
or U14542 (N_14542,N_10879,N_12499);
and U14543 (N_14543,N_9713,N_11281);
or U14544 (N_14544,N_12476,N_11887);
or U14545 (N_14545,N_11564,N_12231);
nand U14546 (N_14546,N_9581,N_10138);
or U14547 (N_14547,N_12375,N_10151);
and U14548 (N_14548,N_9750,N_10710);
and U14549 (N_14549,N_11335,N_10671);
and U14550 (N_14550,N_11681,N_10782);
nand U14551 (N_14551,N_12010,N_9726);
or U14552 (N_14552,N_9376,N_9533);
or U14553 (N_14553,N_10573,N_11095);
nand U14554 (N_14554,N_10696,N_10445);
xnor U14555 (N_14555,N_10937,N_10392);
or U14556 (N_14556,N_10645,N_12034);
nand U14557 (N_14557,N_10399,N_9671);
nor U14558 (N_14558,N_10794,N_11830);
and U14559 (N_14559,N_10408,N_11514);
xnor U14560 (N_14560,N_11312,N_11624);
or U14561 (N_14561,N_10513,N_10611);
xor U14562 (N_14562,N_12068,N_10966);
or U14563 (N_14563,N_9563,N_10587);
and U14564 (N_14564,N_10998,N_9526);
or U14565 (N_14565,N_10329,N_10642);
and U14566 (N_14566,N_10683,N_9622);
and U14567 (N_14567,N_11982,N_10081);
nor U14568 (N_14568,N_11661,N_10681);
and U14569 (N_14569,N_11863,N_10811);
nand U14570 (N_14570,N_9611,N_9727);
and U14571 (N_14571,N_9495,N_10498);
nor U14572 (N_14572,N_10089,N_10518);
nor U14573 (N_14573,N_10273,N_9391);
xnor U14574 (N_14574,N_11283,N_10087);
or U14575 (N_14575,N_9468,N_12088);
or U14576 (N_14576,N_11839,N_11483);
nand U14577 (N_14577,N_12039,N_11754);
xnor U14578 (N_14578,N_11923,N_12361);
nand U14579 (N_14579,N_11309,N_12374);
xor U14580 (N_14580,N_9497,N_10834);
or U14581 (N_14581,N_10147,N_9721);
and U14582 (N_14582,N_9464,N_9747);
nand U14583 (N_14583,N_11123,N_10990);
nand U14584 (N_14584,N_11753,N_9652);
or U14585 (N_14585,N_11836,N_11491);
and U14586 (N_14586,N_11796,N_11940);
nand U14587 (N_14587,N_10299,N_10000);
nor U14588 (N_14588,N_10464,N_9943);
or U14589 (N_14589,N_11143,N_10029);
nand U14590 (N_14590,N_11329,N_11795);
nand U14591 (N_14591,N_9912,N_9741);
or U14592 (N_14592,N_11692,N_12272);
nand U14593 (N_14593,N_11793,N_9767);
nor U14594 (N_14594,N_9813,N_9525);
nand U14595 (N_14595,N_10902,N_10385);
and U14596 (N_14596,N_10777,N_12330);
and U14597 (N_14597,N_9381,N_11655);
nand U14598 (N_14598,N_11898,N_10059);
or U14599 (N_14599,N_9971,N_10512);
and U14600 (N_14600,N_10366,N_11473);
and U14601 (N_14601,N_9569,N_12265);
nand U14602 (N_14602,N_9639,N_9921);
xnor U14603 (N_14603,N_10247,N_11726);
nor U14604 (N_14604,N_11183,N_10166);
nor U14605 (N_14605,N_10495,N_10144);
nand U14606 (N_14606,N_12014,N_11935);
or U14607 (N_14607,N_12043,N_10764);
nand U14608 (N_14608,N_9658,N_12376);
and U14609 (N_14609,N_10348,N_9790);
and U14610 (N_14610,N_12380,N_10435);
xor U14611 (N_14611,N_10944,N_12100);
nand U14612 (N_14612,N_11691,N_11323);
nand U14613 (N_14613,N_12175,N_11952);
nand U14614 (N_14614,N_11900,N_12052);
and U14615 (N_14615,N_12074,N_10540);
or U14616 (N_14616,N_10607,N_11752);
nor U14617 (N_14617,N_9408,N_11923);
nor U14618 (N_14618,N_12131,N_12158);
and U14619 (N_14619,N_10832,N_10181);
nor U14620 (N_14620,N_10357,N_9447);
nor U14621 (N_14621,N_10959,N_11179);
nor U14622 (N_14622,N_10358,N_9562);
nor U14623 (N_14623,N_12272,N_9975);
nand U14624 (N_14624,N_10675,N_10039);
or U14625 (N_14625,N_11564,N_11769);
or U14626 (N_14626,N_11028,N_10908);
nand U14627 (N_14627,N_10907,N_11468);
nand U14628 (N_14628,N_11603,N_9421);
nand U14629 (N_14629,N_11709,N_10098);
nand U14630 (N_14630,N_10954,N_11522);
nand U14631 (N_14631,N_10404,N_11559);
and U14632 (N_14632,N_10198,N_10834);
nand U14633 (N_14633,N_12122,N_12405);
nand U14634 (N_14634,N_10333,N_11717);
nand U14635 (N_14635,N_11513,N_9537);
nor U14636 (N_14636,N_11171,N_10677);
nand U14637 (N_14637,N_12362,N_10351);
and U14638 (N_14638,N_11829,N_11816);
or U14639 (N_14639,N_10918,N_11640);
and U14640 (N_14640,N_9934,N_10203);
or U14641 (N_14641,N_10734,N_10678);
nand U14642 (N_14642,N_12434,N_9451);
xor U14643 (N_14643,N_9909,N_10454);
nand U14644 (N_14644,N_11919,N_9875);
nand U14645 (N_14645,N_9493,N_9880);
nand U14646 (N_14646,N_11662,N_11376);
nand U14647 (N_14647,N_9675,N_11273);
or U14648 (N_14648,N_11270,N_11154);
and U14649 (N_14649,N_11509,N_9594);
and U14650 (N_14650,N_11749,N_9950);
nand U14651 (N_14651,N_11544,N_9530);
nand U14652 (N_14652,N_12176,N_11421);
and U14653 (N_14653,N_10437,N_12113);
xnor U14654 (N_14654,N_10516,N_9895);
or U14655 (N_14655,N_12464,N_9379);
and U14656 (N_14656,N_11290,N_11880);
and U14657 (N_14657,N_10411,N_11886);
nand U14658 (N_14658,N_11523,N_11049);
or U14659 (N_14659,N_11676,N_10622);
nand U14660 (N_14660,N_9925,N_12229);
or U14661 (N_14661,N_10160,N_11345);
and U14662 (N_14662,N_11053,N_11134);
xor U14663 (N_14663,N_10307,N_10428);
nand U14664 (N_14664,N_12210,N_12166);
nor U14665 (N_14665,N_12101,N_11040);
or U14666 (N_14666,N_10788,N_10542);
and U14667 (N_14667,N_11405,N_11597);
or U14668 (N_14668,N_11995,N_9531);
or U14669 (N_14669,N_11776,N_10857);
nor U14670 (N_14670,N_11411,N_9734);
nand U14671 (N_14671,N_10601,N_9427);
nand U14672 (N_14672,N_9853,N_10311);
nor U14673 (N_14673,N_10907,N_9890);
nor U14674 (N_14674,N_11105,N_10868);
nand U14675 (N_14675,N_12347,N_9502);
and U14676 (N_14676,N_11968,N_9740);
xnor U14677 (N_14677,N_11930,N_10268);
nand U14678 (N_14678,N_10724,N_9643);
or U14679 (N_14679,N_9498,N_10118);
nor U14680 (N_14680,N_10431,N_9764);
and U14681 (N_14681,N_11612,N_10773);
and U14682 (N_14682,N_10386,N_12494);
or U14683 (N_14683,N_10779,N_9825);
nand U14684 (N_14684,N_9648,N_11484);
nand U14685 (N_14685,N_10807,N_10308);
nor U14686 (N_14686,N_9698,N_9671);
and U14687 (N_14687,N_11112,N_10120);
nand U14688 (N_14688,N_11523,N_12062);
nand U14689 (N_14689,N_11770,N_9455);
and U14690 (N_14690,N_11333,N_9810);
or U14691 (N_14691,N_9457,N_11659);
nor U14692 (N_14692,N_10357,N_12217);
or U14693 (N_14693,N_9497,N_11398);
nor U14694 (N_14694,N_11142,N_9548);
xor U14695 (N_14695,N_12449,N_11295);
or U14696 (N_14696,N_9966,N_11201);
nor U14697 (N_14697,N_11888,N_10762);
and U14698 (N_14698,N_9695,N_11871);
or U14699 (N_14699,N_12037,N_11335);
and U14700 (N_14700,N_9976,N_11309);
nand U14701 (N_14701,N_11888,N_11066);
and U14702 (N_14702,N_9901,N_9501);
nor U14703 (N_14703,N_10920,N_9765);
nand U14704 (N_14704,N_11600,N_11590);
nor U14705 (N_14705,N_11129,N_11646);
or U14706 (N_14706,N_11180,N_9712);
and U14707 (N_14707,N_12191,N_9608);
and U14708 (N_14708,N_11555,N_10651);
or U14709 (N_14709,N_10922,N_9721);
nor U14710 (N_14710,N_12021,N_9457);
or U14711 (N_14711,N_11307,N_9833);
nand U14712 (N_14712,N_11166,N_9701);
or U14713 (N_14713,N_9948,N_12474);
and U14714 (N_14714,N_12248,N_11101);
and U14715 (N_14715,N_11621,N_11084);
and U14716 (N_14716,N_12255,N_11610);
and U14717 (N_14717,N_12108,N_10735);
xor U14718 (N_14718,N_11084,N_11278);
nand U14719 (N_14719,N_10926,N_10777);
nand U14720 (N_14720,N_10542,N_10408);
and U14721 (N_14721,N_9451,N_12361);
nand U14722 (N_14722,N_11991,N_12275);
nand U14723 (N_14723,N_12129,N_11878);
and U14724 (N_14724,N_10239,N_12207);
nor U14725 (N_14725,N_11713,N_11748);
and U14726 (N_14726,N_11560,N_11711);
or U14727 (N_14727,N_11310,N_11930);
nand U14728 (N_14728,N_12082,N_10708);
and U14729 (N_14729,N_11821,N_11517);
xnor U14730 (N_14730,N_12125,N_11651);
nand U14731 (N_14731,N_10711,N_10035);
nor U14732 (N_14732,N_9927,N_10927);
nor U14733 (N_14733,N_12269,N_12135);
or U14734 (N_14734,N_11199,N_10805);
nor U14735 (N_14735,N_10510,N_11619);
and U14736 (N_14736,N_10554,N_12424);
nor U14737 (N_14737,N_10309,N_10725);
and U14738 (N_14738,N_11348,N_9473);
and U14739 (N_14739,N_11791,N_9592);
and U14740 (N_14740,N_10607,N_12332);
and U14741 (N_14741,N_10533,N_11684);
nand U14742 (N_14742,N_11378,N_9920);
nor U14743 (N_14743,N_11046,N_11590);
or U14744 (N_14744,N_11029,N_10528);
nand U14745 (N_14745,N_10533,N_11360);
and U14746 (N_14746,N_10802,N_11828);
and U14747 (N_14747,N_10131,N_9778);
or U14748 (N_14748,N_11141,N_11145);
and U14749 (N_14749,N_12379,N_9693);
or U14750 (N_14750,N_10596,N_10047);
and U14751 (N_14751,N_10487,N_9891);
or U14752 (N_14752,N_11893,N_11724);
nor U14753 (N_14753,N_10292,N_10362);
nand U14754 (N_14754,N_11511,N_11541);
or U14755 (N_14755,N_10252,N_10477);
and U14756 (N_14756,N_10320,N_10008);
and U14757 (N_14757,N_9707,N_10811);
nor U14758 (N_14758,N_10908,N_11167);
and U14759 (N_14759,N_9947,N_11011);
nand U14760 (N_14760,N_9687,N_11431);
or U14761 (N_14761,N_12005,N_11647);
xor U14762 (N_14762,N_11580,N_10943);
or U14763 (N_14763,N_11845,N_12360);
xor U14764 (N_14764,N_10465,N_10742);
and U14765 (N_14765,N_12141,N_10958);
nor U14766 (N_14766,N_10051,N_11855);
or U14767 (N_14767,N_10647,N_10981);
xor U14768 (N_14768,N_12379,N_10162);
nor U14769 (N_14769,N_9974,N_10956);
nand U14770 (N_14770,N_11212,N_11234);
and U14771 (N_14771,N_10243,N_10214);
or U14772 (N_14772,N_12054,N_10238);
or U14773 (N_14773,N_10135,N_10922);
and U14774 (N_14774,N_12433,N_10810);
nor U14775 (N_14775,N_11599,N_9891);
nand U14776 (N_14776,N_9909,N_10590);
nor U14777 (N_14777,N_11142,N_10594);
nor U14778 (N_14778,N_10709,N_12337);
or U14779 (N_14779,N_10199,N_10009);
nand U14780 (N_14780,N_10353,N_11414);
and U14781 (N_14781,N_11536,N_11736);
and U14782 (N_14782,N_12100,N_12061);
nand U14783 (N_14783,N_12251,N_12356);
nor U14784 (N_14784,N_11988,N_10680);
nor U14785 (N_14785,N_9660,N_10398);
nor U14786 (N_14786,N_9900,N_11515);
or U14787 (N_14787,N_9791,N_12130);
nor U14788 (N_14788,N_12173,N_10812);
nor U14789 (N_14789,N_10162,N_9807);
xnor U14790 (N_14790,N_9999,N_11347);
nand U14791 (N_14791,N_10603,N_9635);
or U14792 (N_14792,N_9871,N_9865);
or U14793 (N_14793,N_11869,N_11691);
or U14794 (N_14794,N_11309,N_12273);
and U14795 (N_14795,N_9974,N_11491);
and U14796 (N_14796,N_10045,N_10441);
xor U14797 (N_14797,N_11585,N_11275);
and U14798 (N_14798,N_10060,N_10003);
nand U14799 (N_14799,N_11917,N_9853);
and U14800 (N_14800,N_11608,N_11577);
nand U14801 (N_14801,N_12296,N_10978);
and U14802 (N_14802,N_9976,N_12009);
nand U14803 (N_14803,N_10989,N_12082);
nor U14804 (N_14804,N_12192,N_10403);
nand U14805 (N_14805,N_10641,N_9802);
and U14806 (N_14806,N_9473,N_10518);
nand U14807 (N_14807,N_12184,N_9468);
and U14808 (N_14808,N_10107,N_9401);
nand U14809 (N_14809,N_10554,N_12193);
nor U14810 (N_14810,N_10924,N_9945);
nor U14811 (N_14811,N_11571,N_9478);
nand U14812 (N_14812,N_10035,N_11122);
and U14813 (N_14813,N_11443,N_10680);
and U14814 (N_14814,N_10876,N_12359);
and U14815 (N_14815,N_10148,N_12484);
and U14816 (N_14816,N_10463,N_12128);
and U14817 (N_14817,N_11466,N_12145);
nor U14818 (N_14818,N_9767,N_10688);
xor U14819 (N_14819,N_11817,N_11971);
nand U14820 (N_14820,N_11720,N_9657);
nand U14821 (N_14821,N_11460,N_11468);
nor U14822 (N_14822,N_9982,N_12159);
nand U14823 (N_14823,N_12465,N_10338);
or U14824 (N_14824,N_11177,N_10037);
xnor U14825 (N_14825,N_10396,N_11548);
xor U14826 (N_14826,N_12075,N_12341);
and U14827 (N_14827,N_11900,N_11156);
or U14828 (N_14828,N_11937,N_12489);
and U14829 (N_14829,N_12497,N_11834);
nor U14830 (N_14830,N_12314,N_12343);
xor U14831 (N_14831,N_10417,N_10649);
nor U14832 (N_14832,N_10891,N_12412);
xnor U14833 (N_14833,N_9564,N_10403);
and U14834 (N_14834,N_11427,N_10863);
xnor U14835 (N_14835,N_11924,N_9840);
or U14836 (N_14836,N_9520,N_12423);
and U14837 (N_14837,N_11137,N_9874);
nand U14838 (N_14838,N_10172,N_11553);
nand U14839 (N_14839,N_10413,N_10108);
nor U14840 (N_14840,N_11749,N_10837);
xnor U14841 (N_14841,N_10714,N_12459);
nor U14842 (N_14842,N_12371,N_11417);
nor U14843 (N_14843,N_11394,N_11769);
and U14844 (N_14844,N_11010,N_11518);
and U14845 (N_14845,N_11555,N_12270);
and U14846 (N_14846,N_9984,N_11400);
or U14847 (N_14847,N_11337,N_10213);
nor U14848 (N_14848,N_10401,N_10482);
nand U14849 (N_14849,N_11273,N_9796);
and U14850 (N_14850,N_11559,N_12201);
xnor U14851 (N_14851,N_10987,N_9829);
nand U14852 (N_14852,N_10630,N_9872);
nor U14853 (N_14853,N_12096,N_11150);
and U14854 (N_14854,N_10576,N_10208);
and U14855 (N_14855,N_9809,N_9427);
and U14856 (N_14856,N_11551,N_11175);
and U14857 (N_14857,N_10348,N_10340);
or U14858 (N_14858,N_10959,N_12083);
or U14859 (N_14859,N_12270,N_9468);
nand U14860 (N_14860,N_9789,N_11346);
or U14861 (N_14861,N_11448,N_10412);
nor U14862 (N_14862,N_12183,N_12108);
nor U14863 (N_14863,N_10980,N_10585);
nor U14864 (N_14864,N_12174,N_10501);
nand U14865 (N_14865,N_11454,N_11043);
nand U14866 (N_14866,N_10112,N_9768);
or U14867 (N_14867,N_11735,N_10020);
nor U14868 (N_14868,N_11981,N_10798);
and U14869 (N_14869,N_10288,N_9612);
nand U14870 (N_14870,N_10348,N_10528);
or U14871 (N_14871,N_10200,N_10002);
xor U14872 (N_14872,N_11593,N_11044);
or U14873 (N_14873,N_10774,N_9490);
nor U14874 (N_14874,N_12261,N_12231);
and U14875 (N_14875,N_10454,N_10711);
or U14876 (N_14876,N_11993,N_12229);
and U14877 (N_14877,N_10498,N_9393);
or U14878 (N_14878,N_11525,N_10604);
nand U14879 (N_14879,N_10451,N_11073);
and U14880 (N_14880,N_12181,N_11701);
nor U14881 (N_14881,N_11573,N_12418);
nand U14882 (N_14882,N_10422,N_11293);
and U14883 (N_14883,N_10328,N_10506);
nor U14884 (N_14884,N_9961,N_10181);
or U14885 (N_14885,N_12299,N_10721);
or U14886 (N_14886,N_10762,N_10715);
nand U14887 (N_14887,N_11919,N_10184);
nand U14888 (N_14888,N_10110,N_9612);
or U14889 (N_14889,N_11607,N_12122);
and U14890 (N_14890,N_11920,N_9567);
nor U14891 (N_14891,N_11149,N_10899);
nand U14892 (N_14892,N_10320,N_11634);
and U14893 (N_14893,N_9860,N_10845);
xnor U14894 (N_14894,N_11038,N_10435);
and U14895 (N_14895,N_10744,N_9667);
nor U14896 (N_14896,N_9382,N_10328);
or U14897 (N_14897,N_9704,N_9913);
nand U14898 (N_14898,N_12179,N_9678);
or U14899 (N_14899,N_9510,N_9732);
xor U14900 (N_14900,N_10369,N_11093);
nor U14901 (N_14901,N_9391,N_12041);
nor U14902 (N_14902,N_9440,N_12416);
nand U14903 (N_14903,N_10134,N_11227);
and U14904 (N_14904,N_10551,N_12373);
or U14905 (N_14905,N_9569,N_11351);
and U14906 (N_14906,N_10813,N_10374);
nand U14907 (N_14907,N_12349,N_11556);
and U14908 (N_14908,N_10595,N_9633);
and U14909 (N_14909,N_9390,N_12322);
nor U14910 (N_14910,N_11555,N_9590);
or U14911 (N_14911,N_9593,N_10549);
nand U14912 (N_14912,N_10255,N_12072);
or U14913 (N_14913,N_11165,N_10669);
nand U14914 (N_14914,N_10844,N_11356);
nor U14915 (N_14915,N_12056,N_11521);
nor U14916 (N_14916,N_9714,N_11986);
or U14917 (N_14917,N_9486,N_12383);
and U14918 (N_14918,N_10928,N_10749);
nor U14919 (N_14919,N_12313,N_9923);
or U14920 (N_14920,N_9650,N_10402);
nor U14921 (N_14921,N_9978,N_10176);
nor U14922 (N_14922,N_10552,N_10617);
nor U14923 (N_14923,N_11851,N_11123);
or U14924 (N_14924,N_9922,N_11467);
or U14925 (N_14925,N_10893,N_10314);
xor U14926 (N_14926,N_10502,N_10871);
nand U14927 (N_14927,N_10136,N_10863);
nor U14928 (N_14928,N_11479,N_12018);
nand U14929 (N_14929,N_10317,N_10349);
nand U14930 (N_14930,N_12069,N_10228);
or U14931 (N_14931,N_12105,N_11363);
or U14932 (N_14932,N_10157,N_11384);
nand U14933 (N_14933,N_11469,N_10497);
or U14934 (N_14934,N_10087,N_11376);
and U14935 (N_14935,N_10188,N_9682);
or U14936 (N_14936,N_12001,N_9502);
and U14937 (N_14937,N_9989,N_10110);
and U14938 (N_14938,N_12446,N_9684);
and U14939 (N_14939,N_9514,N_11541);
and U14940 (N_14940,N_11242,N_9837);
or U14941 (N_14941,N_12069,N_10817);
nor U14942 (N_14942,N_11267,N_10984);
and U14943 (N_14943,N_11928,N_12462);
or U14944 (N_14944,N_9416,N_11305);
nand U14945 (N_14945,N_10629,N_10393);
nor U14946 (N_14946,N_10162,N_10626);
and U14947 (N_14947,N_10393,N_9671);
nor U14948 (N_14948,N_9783,N_11695);
xnor U14949 (N_14949,N_10161,N_11818);
xnor U14950 (N_14950,N_9588,N_12242);
nand U14951 (N_14951,N_10380,N_10911);
nor U14952 (N_14952,N_10763,N_11303);
nand U14953 (N_14953,N_11970,N_12468);
and U14954 (N_14954,N_12385,N_10447);
or U14955 (N_14955,N_12009,N_12328);
nor U14956 (N_14956,N_9603,N_11799);
and U14957 (N_14957,N_10872,N_10942);
nor U14958 (N_14958,N_12023,N_9560);
and U14959 (N_14959,N_12291,N_10021);
nor U14960 (N_14960,N_10892,N_11401);
and U14961 (N_14961,N_10718,N_9809);
nand U14962 (N_14962,N_12388,N_11258);
nor U14963 (N_14963,N_11302,N_12326);
and U14964 (N_14964,N_11904,N_11103);
nand U14965 (N_14965,N_10020,N_10897);
nor U14966 (N_14966,N_10007,N_12466);
xnor U14967 (N_14967,N_12307,N_11690);
and U14968 (N_14968,N_10225,N_11128);
nand U14969 (N_14969,N_10015,N_9503);
nor U14970 (N_14970,N_11966,N_10474);
nand U14971 (N_14971,N_11946,N_9874);
and U14972 (N_14972,N_9859,N_12444);
nand U14973 (N_14973,N_10273,N_11959);
xnor U14974 (N_14974,N_10491,N_10220);
nand U14975 (N_14975,N_9550,N_10773);
nand U14976 (N_14976,N_11143,N_10306);
and U14977 (N_14977,N_11335,N_12156);
nor U14978 (N_14978,N_12021,N_11981);
and U14979 (N_14979,N_10829,N_12159);
xor U14980 (N_14980,N_11026,N_11266);
nand U14981 (N_14981,N_12365,N_11119);
and U14982 (N_14982,N_10033,N_10354);
and U14983 (N_14983,N_12386,N_10355);
nor U14984 (N_14984,N_11687,N_12160);
nand U14985 (N_14985,N_9971,N_11721);
and U14986 (N_14986,N_11709,N_11657);
nor U14987 (N_14987,N_11690,N_11891);
xor U14988 (N_14988,N_11933,N_10200);
nand U14989 (N_14989,N_9961,N_9677);
nand U14990 (N_14990,N_10956,N_12282);
nand U14991 (N_14991,N_12002,N_12090);
nor U14992 (N_14992,N_12143,N_10519);
nand U14993 (N_14993,N_10948,N_9987);
and U14994 (N_14994,N_11959,N_9847);
and U14995 (N_14995,N_12413,N_11847);
nand U14996 (N_14996,N_11182,N_11869);
or U14997 (N_14997,N_11023,N_10820);
nor U14998 (N_14998,N_11289,N_10402);
and U14999 (N_14999,N_9485,N_11677);
or U15000 (N_15000,N_11818,N_9820);
or U15001 (N_15001,N_10462,N_12063);
nand U15002 (N_15002,N_10932,N_9417);
and U15003 (N_15003,N_10599,N_9923);
nand U15004 (N_15004,N_11255,N_11969);
nand U15005 (N_15005,N_9424,N_11291);
and U15006 (N_15006,N_9523,N_9669);
and U15007 (N_15007,N_11246,N_11480);
xnor U15008 (N_15008,N_9512,N_11117);
and U15009 (N_15009,N_10285,N_11392);
xor U15010 (N_15010,N_11421,N_12360);
nand U15011 (N_15011,N_11013,N_12322);
and U15012 (N_15012,N_12402,N_10137);
nand U15013 (N_15013,N_12173,N_10112);
or U15014 (N_15014,N_10036,N_11491);
and U15015 (N_15015,N_11778,N_12157);
xor U15016 (N_15016,N_11272,N_10614);
or U15017 (N_15017,N_9978,N_11682);
or U15018 (N_15018,N_11130,N_10310);
or U15019 (N_15019,N_10261,N_10141);
nor U15020 (N_15020,N_11388,N_10885);
nand U15021 (N_15021,N_11693,N_9989);
nand U15022 (N_15022,N_10314,N_12001);
nand U15023 (N_15023,N_10909,N_11043);
and U15024 (N_15024,N_10874,N_12439);
nor U15025 (N_15025,N_11747,N_12388);
and U15026 (N_15026,N_10323,N_10412);
and U15027 (N_15027,N_9523,N_9812);
nand U15028 (N_15028,N_10759,N_11198);
and U15029 (N_15029,N_10886,N_11049);
nand U15030 (N_15030,N_9751,N_10671);
nor U15031 (N_15031,N_11946,N_9936);
or U15032 (N_15032,N_11921,N_10650);
or U15033 (N_15033,N_10924,N_12307);
nand U15034 (N_15034,N_11633,N_10476);
xnor U15035 (N_15035,N_10279,N_10352);
and U15036 (N_15036,N_9911,N_10604);
nor U15037 (N_15037,N_11407,N_9589);
nand U15038 (N_15038,N_12071,N_12393);
or U15039 (N_15039,N_9591,N_11161);
and U15040 (N_15040,N_12488,N_11944);
or U15041 (N_15041,N_10568,N_10479);
nand U15042 (N_15042,N_12098,N_12348);
nand U15043 (N_15043,N_11002,N_9765);
nor U15044 (N_15044,N_12237,N_11634);
nand U15045 (N_15045,N_11580,N_9734);
nor U15046 (N_15046,N_10475,N_10425);
or U15047 (N_15047,N_11715,N_12134);
nand U15048 (N_15048,N_10124,N_11105);
nand U15049 (N_15049,N_11790,N_9743);
nand U15050 (N_15050,N_11539,N_11968);
nor U15051 (N_15051,N_11895,N_11137);
nor U15052 (N_15052,N_9624,N_11420);
nor U15053 (N_15053,N_10439,N_11086);
or U15054 (N_15054,N_11303,N_10829);
and U15055 (N_15055,N_10856,N_9614);
and U15056 (N_15056,N_9809,N_11908);
nor U15057 (N_15057,N_10219,N_9647);
nor U15058 (N_15058,N_10142,N_9705);
nand U15059 (N_15059,N_9379,N_12254);
nand U15060 (N_15060,N_11246,N_10900);
or U15061 (N_15061,N_9835,N_12002);
nand U15062 (N_15062,N_9642,N_11126);
xnor U15063 (N_15063,N_12157,N_9412);
xor U15064 (N_15064,N_11688,N_11070);
nor U15065 (N_15065,N_10587,N_11819);
nor U15066 (N_15066,N_12023,N_9418);
and U15067 (N_15067,N_11785,N_12395);
nand U15068 (N_15068,N_12390,N_12458);
nor U15069 (N_15069,N_11279,N_11189);
nor U15070 (N_15070,N_11179,N_12065);
or U15071 (N_15071,N_11406,N_9890);
and U15072 (N_15072,N_12402,N_9591);
nand U15073 (N_15073,N_11232,N_12327);
xor U15074 (N_15074,N_12092,N_10057);
xor U15075 (N_15075,N_11827,N_11430);
nand U15076 (N_15076,N_10333,N_12172);
or U15077 (N_15077,N_9694,N_9496);
and U15078 (N_15078,N_10600,N_11416);
nand U15079 (N_15079,N_10056,N_11639);
nand U15080 (N_15080,N_12287,N_12307);
or U15081 (N_15081,N_10036,N_12172);
nor U15082 (N_15082,N_11892,N_12411);
nor U15083 (N_15083,N_11814,N_11140);
nand U15084 (N_15084,N_11628,N_10839);
nand U15085 (N_15085,N_10713,N_10172);
or U15086 (N_15086,N_11873,N_10553);
nand U15087 (N_15087,N_10073,N_11276);
nor U15088 (N_15088,N_12341,N_12463);
xnor U15089 (N_15089,N_9836,N_12025);
nand U15090 (N_15090,N_11430,N_11218);
or U15091 (N_15091,N_12206,N_12199);
nor U15092 (N_15092,N_10059,N_11493);
and U15093 (N_15093,N_11579,N_11157);
and U15094 (N_15094,N_10234,N_10289);
or U15095 (N_15095,N_10348,N_11097);
xnor U15096 (N_15096,N_10194,N_11720);
or U15097 (N_15097,N_11953,N_10677);
xnor U15098 (N_15098,N_10997,N_10785);
or U15099 (N_15099,N_12455,N_11360);
and U15100 (N_15100,N_9974,N_10742);
or U15101 (N_15101,N_10033,N_12392);
xnor U15102 (N_15102,N_10362,N_12260);
xnor U15103 (N_15103,N_10861,N_10675);
nand U15104 (N_15104,N_9568,N_10854);
xor U15105 (N_15105,N_10470,N_11525);
nand U15106 (N_15106,N_10851,N_11455);
nor U15107 (N_15107,N_11517,N_10563);
nor U15108 (N_15108,N_11639,N_11612);
nor U15109 (N_15109,N_11309,N_11088);
nor U15110 (N_15110,N_9948,N_9878);
or U15111 (N_15111,N_9971,N_11213);
nand U15112 (N_15112,N_9818,N_10580);
nor U15113 (N_15113,N_11050,N_11846);
xnor U15114 (N_15114,N_9781,N_10507);
nand U15115 (N_15115,N_10164,N_11444);
nor U15116 (N_15116,N_10319,N_10363);
nor U15117 (N_15117,N_11388,N_12326);
and U15118 (N_15118,N_10711,N_10611);
and U15119 (N_15119,N_12054,N_11136);
nor U15120 (N_15120,N_12478,N_12163);
nor U15121 (N_15121,N_11848,N_10414);
xnor U15122 (N_15122,N_9876,N_11958);
or U15123 (N_15123,N_9521,N_9990);
or U15124 (N_15124,N_11441,N_11823);
nor U15125 (N_15125,N_11556,N_10654);
or U15126 (N_15126,N_11222,N_12019);
nand U15127 (N_15127,N_12016,N_9620);
nor U15128 (N_15128,N_10801,N_10610);
xor U15129 (N_15129,N_9543,N_11863);
and U15130 (N_15130,N_9635,N_11529);
nor U15131 (N_15131,N_10123,N_9860);
xor U15132 (N_15132,N_10666,N_9608);
or U15133 (N_15133,N_10099,N_10439);
nor U15134 (N_15134,N_10860,N_11920);
or U15135 (N_15135,N_12135,N_9740);
nor U15136 (N_15136,N_10113,N_10007);
or U15137 (N_15137,N_11910,N_12362);
or U15138 (N_15138,N_12010,N_12159);
and U15139 (N_15139,N_10216,N_10631);
nor U15140 (N_15140,N_11797,N_11603);
nor U15141 (N_15141,N_10148,N_9525);
nor U15142 (N_15142,N_11002,N_11215);
and U15143 (N_15143,N_10979,N_9801);
and U15144 (N_15144,N_11977,N_11273);
or U15145 (N_15145,N_9843,N_11329);
nor U15146 (N_15146,N_9408,N_10244);
nor U15147 (N_15147,N_9939,N_9656);
nor U15148 (N_15148,N_11590,N_10005);
or U15149 (N_15149,N_9938,N_9737);
nand U15150 (N_15150,N_10322,N_10065);
and U15151 (N_15151,N_12318,N_12305);
or U15152 (N_15152,N_10364,N_11685);
nor U15153 (N_15153,N_11401,N_10877);
nor U15154 (N_15154,N_11428,N_11013);
xnor U15155 (N_15155,N_11669,N_12380);
nand U15156 (N_15156,N_9402,N_10285);
xnor U15157 (N_15157,N_10831,N_12341);
and U15158 (N_15158,N_10328,N_12347);
or U15159 (N_15159,N_12018,N_11899);
nand U15160 (N_15160,N_10054,N_10347);
nand U15161 (N_15161,N_12140,N_10891);
nand U15162 (N_15162,N_10574,N_12284);
nor U15163 (N_15163,N_9811,N_9860);
or U15164 (N_15164,N_9808,N_11896);
nor U15165 (N_15165,N_10434,N_10133);
nor U15166 (N_15166,N_10890,N_11298);
nor U15167 (N_15167,N_12053,N_11650);
nand U15168 (N_15168,N_12372,N_11699);
or U15169 (N_15169,N_11244,N_10959);
nor U15170 (N_15170,N_12324,N_11196);
nor U15171 (N_15171,N_9669,N_9453);
and U15172 (N_15172,N_10382,N_9653);
nor U15173 (N_15173,N_9658,N_9383);
nand U15174 (N_15174,N_10740,N_10203);
nor U15175 (N_15175,N_10561,N_11625);
and U15176 (N_15176,N_12054,N_11844);
or U15177 (N_15177,N_11288,N_10354);
nand U15178 (N_15178,N_11063,N_12005);
and U15179 (N_15179,N_10096,N_11255);
and U15180 (N_15180,N_9508,N_9858);
or U15181 (N_15181,N_12123,N_9965);
nand U15182 (N_15182,N_11690,N_12266);
or U15183 (N_15183,N_10769,N_10112);
or U15184 (N_15184,N_11219,N_12469);
and U15185 (N_15185,N_11127,N_10840);
or U15186 (N_15186,N_9705,N_11420);
and U15187 (N_15187,N_9644,N_9815);
nor U15188 (N_15188,N_10164,N_11979);
or U15189 (N_15189,N_11835,N_11803);
nand U15190 (N_15190,N_11436,N_9845);
nand U15191 (N_15191,N_10653,N_9638);
nor U15192 (N_15192,N_9456,N_11974);
nand U15193 (N_15193,N_12080,N_11616);
or U15194 (N_15194,N_11362,N_11836);
nor U15195 (N_15195,N_9839,N_10268);
nand U15196 (N_15196,N_11594,N_10814);
nor U15197 (N_15197,N_10481,N_10614);
nor U15198 (N_15198,N_11224,N_11873);
nor U15199 (N_15199,N_12163,N_10228);
xor U15200 (N_15200,N_9696,N_12390);
or U15201 (N_15201,N_10368,N_11839);
nand U15202 (N_15202,N_10245,N_11494);
nand U15203 (N_15203,N_11630,N_12459);
or U15204 (N_15204,N_11954,N_10873);
and U15205 (N_15205,N_10676,N_10021);
nor U15206 (N_15206,N_9772,N_9510);
xnor U15207 (N_15207,N_11997,N_12253);
and U15208 (N_15208,N_12489,N_11273);
nand U15209 (N_15209,N_10980,N_10074);
and U15210 (N_15210,N_12371,N_10249);
and U15211 (N_15211,N_10261,N_9710);
nand U15212 (N_15212,N_11510,N_11550);
or U15213 (N_15213,N_9823,N_12314);
and U15214 (N_15214,N_12253,N_11984);
nor U15215 (N_15215,N_12388,N_11661);
or U15216 (N_15216,N_11135,N_11922);
nor U15217 (N_15217,N_11658,N_10671);
or U15218 (N_15218,N_11100,N_10240);
nor U15219 (N_15219,N_10630,N_10464);
or U15220 (N_15220,N_11417,N_10214);
nand U15221 (N_15221,N_11906,N_9655);
and U15222 (N_15222,N_11484,N_12264);
or U15223 (N_15223,N_12380,N_11616);
nor U15224 (N_15224,N_12383,N_11980);
or U15225 (N_15225,N_9736,N_11909);
or U15226 (N_15226,N_11648,N_12351);
or U15227 (N_15227,N_11341,N_10269);
nand U15228 (N_15228,N_10453,N_10911);
nand U15229 (N_15229,N_12427,N_11879);
nor U15230 (N_15230,N_9942,N_11641);
nor U15231 (N_15231,N_10938,N_10138);
or U15232 (N_15232,N_11906,N_9583);
or U15233 (N_15233,N_9859,N_11439);
nor U15234 (N_15234,N_11503,N_11726);
nor U15235 (N_15235,N_10533,N_11659);
nand U15236 (N_15236,N_10072,N_9930);
nor U15237 (N_15237,N_9535,N_9569);
nand U15238 (N_15238,N_11579,N_11758);
nand U15239 (N_15239,N_11826,N_10955);
xor U15240 (N_15240,N_10399,N_12187);
and U15241 (N_15241,N_11982,N_10864);
xnor U15242 (N_15242,N_11554,N_10153);
or U15243 (N_15243,N_10990,N_11565);
nand U15244 (N_15244,N_10883,N_11348);
nand U15245 (N_15245,N_11192,N_9443);
and U15246 (N_15246,N_11401,N_10755);
nor U15247 (N_15247,N_12217,N_11874);
and U15248 (N_15248,N_10857,N_10614);
or U15249 (N_15249,N_9978,N_12481);
xnor U15250 (N_15250,N_9575,N_10568);
or U15251 (N_15251,N_11072,N_10358);
and U15252 (N_15252,N_11228,N_10346);
nand U15253 (N_15253,N_11255,N_10263);
xor U15254 (N_15254,N_9604,N_11311);
nor U15255 (N_15255,N_11406,N_9824);
or U15256 (N_15256,N_9785,N_12274);
and U15257 (N_15257,N_11484,N_11028);
and U15258 (N_15258,N_11437,N_9576);
xor U15259 (N_15259,N_11371,N_12383);
or U15260 (N_15260,N_10989,N_10058);
or U15261 (N_15261,N_12214,N_10513);
nand U15262 (N_15262,N_11823,N_11351);
and U15263 (N_15263,N_10703,N_9684);
and U15264 (N_15264,N_10349,N_10693);
nand U15265 (N_15265,N_10446,N_10526);
or U15266 (N_15266,N_10839,N_11696);
and U15267 (N_15267,N_9514,N_9877);
nand U15268 (N_15268,N_11864,N_11214);
nor U15269 (N_15269,N_11606,N_12094);
nand U15270 (N_15270,N_9375,N_11562);
nor U15271 (N_15271,N_11087,N_11525);
and U15272 (N_15272,N_10446,N_9552);
or U15273 (N_15273,N_11411,N_12370);
xor U15274 (N_15274,N_11279,N_10909);
nor U15275 (N_15275,N_11571,N_10475);
xnor U15276 (N_15276,N_11264,N_9573);
and U15277 (N_15277,N_10309,N_10106);
nand U15278 (N_15278,N_10434,N_10804);
xnor U15279 (N_15279,N_12032,N_11769);
or U15280 (N_15280,N_10740,N_10288);
xor U15281 (N_15281,N_10413,N_11332);
or U15282 (N_15282,N_10393,N_12487);
nor U15283 (N_15283,N_11388,N_10636);
and U15284 (N_15284,N_12069,N_11410);
nand U15285 (N_15285,N_10092,N_11701);
nand U15286 (N_15286,N_10291,N_9719);
nand U15287 (N_15287,N_10605,N_10379);
and U15288 (N_15288,N_10698,N_11536);
xor U15289 (N_15289,N_11283,N_9730);
and U15290 (N_15290,N_10838,N_10865);
and U15291 (N_15291,N_11124,N_10978);
nor U15292 (N_15292,N_10550,N_10761);
nand U15293 (N_15293,N_11248,N_11793);
and U15294 (N_15294,N_11649,N_12279);
nand U15295 (N_15295,N_11225,N_10818);
nand U15296 (N_15296,N_12134,N_11984);
and U15297 (N_15297,N_10187,N_11611);
and U15298 (N_15298,N_10986,N_12312);
and U15299 (N_15299,N_11235,N_11182);
nor U15300 (N_15300,N_9942,N_9877);
and U15301 (N_15301,N_10646,N_9920);
or U15302 (N_15302,N_11978,N_11916);
xnor U15303 (N_15303,N_11160,N_11260);
and U15304 (N_15304,N_11772,N_12490);
nor U15305 (N_15305,N_11142,N_10236);
nand U15306 (N_15306,N_9440,N_11612);
nand U15307 (N_15307,N_11677,N_10485);
nand U15308 (N_15308,N_11402,N_10021);
nand U15309 (N_15309,N_10251,N_10486);
and U15310 (N_15310,N_10649,N_12382);
nand U15311 (N_15311,N_9441,N_9774);
nor U15312 (N_15312,N_12370,N_10255);
nand U15313 (N_15313,N_11310,N_12266);
and U15314 (N_15314,N_9562,N_12088);
nand U15315 (N_15315,N_10035,N_10721);
and U15316 (N_15316,N_11418,N_12122);
nor U15317 (N_15317,N_9613,N_12105);
or U15318 (N_15318,N_10021,N_10313);
nand U15319 (N_15319,N_10714,N_11157);
or U15320 (N_15320,N_10244,N_11558);
and U15321 (N_15321,N_9804,N_10606);
nor U15322 (N_15322,N_11180,N_11429);
and U15323 (N_15323,N_12264,N_9602);
nand U15324 (N_15324,N_10327,N_9566);
and U15325 (N_15325,N_9780,N_9476);
nand U15326 (N_15326,N_12165,N_10288);
nor U15327 (N_15327,N_10535,N_10711);
nand U15328 (N_15328,N_11833,N_12461);
and U15329 (N_15329,N_11278,N_11784);
and U15330 (N_15330,N_10468,N_10356);
nor U15331 (N_15331,N_10358,N_11118);
nand U15332 (N_15332,N_10291,N_9950);
or U15333 (N_15333,N_10192,N_9585);
or U15334 (N_15334,N_9401,N_9752);
nand U15335 (N_15335,N_12181,N_12323);
nand U15336 (N_15336,N_12280,N_11970);
or U15337 (N_15337,N_11562,N_10126);
nand U15338 (N_15338,N_11075,N_11703);
and U15339 (N_15339,N_9841,N_11735);
nand U15340 (N_15340,N_12347,N_12147);
and U15341 (N_15341,N_10217,N_11127);
or U15342 (N_15342,N_11121,N_10648);
xor U15343 (N_15343,N_11462,N_9889);
and U15344 (N_15344,N_11271,N_12382);
or U15345 (N_15345,N_9726,N_9517);
nor U15346 (N_15346,N_12328,N_11264);
and U15347 (N_15347,N_10965,N_11958);
and U15348 (N_15348,N_12363,N_9796);
xor U15349 (N_15349,N_10634,N_10095);
and U15350 (N_15350,N_9802,N_10248);
xor U15351 (N_15351,N_10751,N_11284);
xnor U15352 (N_15352,N_9788,N_10585);
nor U15353 (N_15353,N_10337,N_10197);
xnor U15354 (N_15354,N_11889,N_11806);
and U15355 (N_15355,N_9503,N_11820);
nor U15356 (N_15356,N_10151,N_10327);
xor U15357 (N_15357,N_11893,N_11216);
nor U15358 (N_15358,N_10347,N_10030);
or U15359 (N_15359,N_11367,N_10435);
nor U15360 (N_15360,N_10769,N_11255);
xor U15361 (N_15361,N_10625,N_12114);
or U15362 (N_15362,N_11059,N_9851);
or U15363 (N_15363,N_12009,N_9833);
or U15364 (N_15364,N_10337,N_9763);
or U15365 (N_15365,N_11613,N_9716);
nor U15366 (N_15366,N_10368,N_11150);
and U15367 (N_15367,N_10873,N_10926);
nor U15368 (N_15368,N_10680,N_11957);
nand U15369 (N_15369,N_12334,N_10264);
or U15370 (N_15370,N_11677,N_11983);
and U15371 (N_15371,N_11465,N_9910);
and U15372 (N_15372,N_9561,N_11642);
nand U15373 (N_15373,N_9542,N_11410);
and U15374 (N_15374,N_11471,N_11474);
nand U15375 (N_15375,N_12489,N_9948);
and U15376 (N_15376,N_10318,N_10025);
nand U15377 (N_15377,N_9386,N_11149);
or U15378 (N_15378,N_9607,N_10403);
nor U15379 (N_15379,N_10170,N_11721);
nor U15380 (N_15380,N_9599,N_10145);
or U15381 (N_15381,N_10884,N_11179);
and U15382 (N_15382,N_12089,N_9424);
and U15383 (N_15383,N_12025,N_10140);
xnor U15384 (N_15384,N_12441,N_11824);
nor U15385 (N_15385,N_10390,N_12346);
and U15386 (N_15386,N_10315,N_10298);
nand U15387 (N_15387,N_11538,N_11890);
nor U15388 (N_15388,N_12446,N_10929);
or U15389 (N_15389,N_10045,N_10276);
and U15390 (N_15390,N_9704,N_12489);
and U15391 (N_15391,N_12196,N_11434);
nor U15392 (N_15392,N_10508,N_10991);
nor U15393 (N_15393,N_11605,N_10329);
or U15394 (N_15394,N_10880,N_11106);
nor U15395 (N_15395,N_9838,N_9775);
or U15396 (N_15396,N_12478,N_11248);
nor U15397 (N_15397,N_11328,N_11909);
xor U15398 (N_15398,N_12273,N_9929);
or U15399 (N_15399,N_11863,N_12051);
and U15400 (N_15400,N_10819,N_11315);
nor U15401 (N_15401,N_9821,N_11323);
and U15402 (N_15402,N_10670,N_9397);
or U15403 (N_15403,N_9799,N_9618);
or U15404 (N_15404,N_10268,N_11140);
nor U15405 (N_15405,N_12475,N_11683);
nor U15406 (N_15406,N_12164,N_12328);
nand U15407 (N_15407,N_10708,N_11323);
nor U15408 (N_15408,N_10401,N_9867);
nand U15409 (N_15409,N_11990,N_9429);
nand U15410 (N_15410,N_10101,N_12473);
nand U15411 (N_15411,N_11973,N_12432);
nor U15412 (N_15412,N_12160,N_11388);
xor U15413 (N_15413,N_11135,N_10737);
and U15414 (N_15414,N_11581,N_12133);
or U15415 (N_15415,N_10595,N_9406);
or U15416 (N_15416,N_11438,N_11714);
nand U15417 (N_15417,N_11505,N_11799);
or U15418 (N_15418,N_11169,N_10167);
nand U15419 (N_15419,N_11429,N_9729);
and U15420 (N_15420,N_10502,N_11819);
nor U15421 (N_15421,N_11554,N_12161);
and U15422 (N_15422,N_12183,N_12191);
nor U15423 (N_15423,N_12224,N_11584);
nor U15424 (N_15424,N_10360,N_12161);
xor U15425 (N_15425,N_12154,N_10768);
nand U15426 (N_15426,N_9427,N_10549);
and U15427 (N_15427,N_12443,N_10670);
and U15428 (N_15428,N_10520,N_12087);
nor U15429 (N_15429,N_11714,N_11589);
and U15430 (N_15430,N_11514,N_12453);
and U15431 (N_15431,N_10585,N_10013);
nor U15432 (N_15432,N_10800,N_10613);
or U15433 (N_15433,N_10473,N_10272);
and U15434 (N_15434,N_9963,N_12154);
or U15435 (N_15435,N_12232,N_10360);
nor U15436 (N_15436,N_11583,N_11063);
and U15437 (N_15437,N_10259,N_9554);
or U15438 (N_15438,N_9543,N_9822);
nor U15439 (N_15439,N_10649,N_11435);
or U15440 (N_15440,N_11849,N_10053);
or U15441 (N_15441,N_11785,N_12270);
nor U15442 (N_15442,N_10059,N_9531);
or U15443 (N_15443,N_12172,N_10985);
and U15444 (N_15444,N_11957,N_10882);
nand U15445 (N_15445,N_11038,N_9528);
and U15446 (N_15446,N_9400,N_9788);
and U15447 (N_15447,N_11405,N_9995);
and U15448 (N_15448,N_11154,N_9674);
and U15449 (N_15449,N_9452,N_9856);
nor U15450 (N_15450,N_10888,N_10084);
or U15451 (N_15451,N_10086,N_12423);
and U15452 (N_15452,N_11840,N_11443);
and U15453 (N_15453,N_11433,N_11025);
nand U15454 (N_15454,N_9409,N_12376);
nand U15455 (N_15455,N_12225,N_10879);
or U15456 (N_15456,N_9897,N_10989);
nand U15457 (N_15457,N_10350,N_11233);
nor U15458 (N_15458,N_9808,N_10171);
nor U15459 (N_15459,N_9818,N_9447);
and U15460 (N_15460,N_11562,N_10356);
nor U15461 (N_15461,N_10580,N_9742);
xor U15462 (N_15462,N_11447,N_11658);
nor U15463 (N_15463,N_12175,N_10607);
and U15464 (N_15464,N_10445,N_11720);
and U15465 (N_15465,N_10915,N_10557);
xor U15466 (N_15466,N_12235,N_10039);
nand U15467 (N_15467,N_10522,N_12423);
nand U15468 (N_15468,N_10219,N_10249);
and U15469 (N_15469,N_10767,N_9403);
or U15470 (N_15470,N_10498,N_10349);
nor U15471 (N_15471,N_10473,N_9976);
nand U15472 (N_15472,N_10267,N_11840);
and U15473 (N_15473,N_11912,N_11835);
or U15474 (N_15474,N_9708,N_12400);
nor U15475 (N_15475,N_12245,N_10491);
and U15476 (N_15476,N_11731,N_10206);
nor U15477 (N_15477,N_11987,N_11595);
nand U15478 (N_15478,N_11626,N_11833);
nor U15479 (N_15479,N_12031,N_12275);
nor U15480 (N_15480,N_10627,N_12496);
nor U15481 (N_15481,N_12007,N_9419);
nor U15482 (N_15482,N_10438,N_12458);
nand U15483 (N_15483,N_9645,N_11577);
and U15484 (N_15484,N_12032,N_12107);
nand U15485 (N_15485,N_10204,N_12488);
or U15486 (N_15486,N_11226,N_12017);
xor U15487 (N_15487,N_11785,N_9870);
nor U15488 (N_15488,N_10948,N_11823);
and U15489 (N_15489,N_9652,N_9736);
xnor U15490 (N_15490,N_11008,N_12419);
nor U15491 (N_15491,N_11358,N_11910);
nor U15492 (N_15492,N_9710,N_10279);
and U15493 (N_15493,N_9870,N_10772);
nand U15494 (N_15494,N_10941,N_9470);
xnor U15495 (N_15495,N_12105,N_9569);
and U15496 (N_15496,N_10923,N_10823);
and U15497 (N_15497,N_11493,N_10084);
nand U15498 (N_15498,N_11436,N_10120);
or U15499 (N_15499,N_9470,N_10226);
nand U15500 (N_15500,N_9643,N_9932);
and U15501 (N_15501,N_11678,N_9385);
nand U15502 (N_15502,N_11742,N_10788);
nand U15503 (N_15503,N_9418,N_10231);
nor U15504 (N_15504,N_12345,N_11121);
nor U15505 (N_15505,N_10472,N_9499);
or U15506 (N_15506,N_11616,N_11179);
xnor U15507 (N_15507,N_9631,N_11165);
nor U15508 (N_15508,N_12384,N_11063);
and U15509 (N_15509,N_9859,N_10965);
or U15510 (N_15510,N_9631,N_11817);
xnor U15511 (N_15511,N_9442,N_12309);
nand U15512 (N_15512,N_11048,N_11368);
nand U15513 (N_15513,N_10254,N_11336);
nor U15514 (N_15514,N_11668,N_10926);
nand U15515 (N_15515,N_9729,N_9426);
or U15516 (N_15516,N_9833,N_9487);
nor U15517 (N_15517,N_10766,N_11879);
nand U15518 (N_15518,N_11968,N_9929);
nor U15519 (N_15519,N_12037,N_10710);
xor U15520 (N_15520,N_10151,N_10968);
nand U15521 (N_15521,N_10961,N_12205);
nor U15522 (N_15522,N_12322,N_12219);
or U15523 (N_15523,N_10747,N_10942);
and U15524 (N_15524,N_12226,N_10299);
or U15525 (N_15525,N_9567,N_11900);
nand U15526 (N_15526,N_10170,N_11797);
nor U15527 (N_15527,N_12078,N_11952);
nand U15528 (N_15528,N_10916,N_12055);
and U15529 (N_15529,N_11562,N_11165);
or U15530 (N_15530,N_11150,N_12373);
or U15531 (N_15531,N_11752,N_9952);
nand U15532 (N_15532,N_10963,N_11648);
xor U15533 (N_15533,N_12044,N_11974);
or U15534 (N_15534,N_10350,N_9677);
or U15535 (N_15535,N_11603,N_10984);
nand U15536 (N_15536,N_10445,N_11674);
or U15537 (N_15537,N_10708,N_11067);
nand U15538 (N_15538,N_10612,N_11899);
nand U15539 (N_15539,N_12133,N_11208);
and U15540 (N_15540,N_11744,N_9860);
nor U15541 (N_15541,N_10177,N_9764);
nand U15542 (N_15542,N_9453,N_10901);
and U15543 (N_15543,N_9905,N_11766);
xor U15544 (N_15544,N_11175,N_10551);
nand U15545 (N_15545,N_10596,N_10143);
nor U15546 (N_15546,N_9607,N_12418);
or U15547 (N_15547,N_12010,N_9692);
nor U15548 (N_15548,N_9812,N_12330);
or U15549 (N_15549,N_10427,N_10989);
or U15550 (N_15550,N_9744,N_10299);
xnor U15551 (N_15551,N_11887,N_10321);
or U15552 (N_15552,N_11871,N_12087);
nor U15553 (N_15553,N_9626,N_11493);
nor U15554 (N_15554,N_11692,N_10929);
or U15555 (N_15555,N_9856,N_9594);
nand U15556 (N_15556,N_10068,N_11437);
xnor U15557 (N_15557,N_10864,N_11058);
nor U15558 (N_15558,N_11611,N_9487);
nand U15559 (N_15559,N_10653,N_12087);
nor U15560 (N_15560,N_11520,N_9721);
and U15561 (N_15561,N_11715,N_10439);
nor U15562 (N_15562,N_11189,N_11736);
or U15563 (N_15563,N_11380,N_9805);
and U15564 (N_15564,N_10964,N_11912);
xor U15565 (N_15565,N_12161,N_9383);
nand U15566 (N_15566,N_11821,N_10804);
nor U15567 (N_15567,N_11736,N_10712);
and U15568 (N_15568,N_11160,N_10549);
or U15569 (N_15569,N_11779,N_11900);
xor U15570 (N_15570,N_11230,N_11823);
or U15571 (N_15571,N_12066,N_11521);
nor U15572 (N_15572,N_11915,N_12024);
nand U15573 (N_15573,N_11699,N_10574);
nand U15574 (N_15574,N_11427,N_9924);
and U15575 (N_15575,N_12019,N_11350);
nand U15576 (N_15576,N_12386,N_11846);
nor U15577 (N_15577,N_9403,N_10645);
and U15578 (N_15578,N_9960,N_9932);
and U15579 (N_15579,N_11978,N_10886);
nor U15580 (N_15580,N_9701,N_11863);
and U15581 (N_15581,N_10623,N_10329);
or U15582 (N_15582,N_10398,N_12488);
or U15583 (N_15583,N_9876,N_12172);
or U15584 (N_15584,N_12328,N_9430);
or U15585 (N_15585,N_9689,N_10867);
nor U15586 (N_15586,N_11220,N_11139);
nor U15587 (N_15587,N_9555,N_9380);
xor U15588 (N_15588,N_11809,N_10707);
nor U15589 (N_15589,N_12153,N_10644);
nand U15590 (N_15590,N_9616,N_11318);
or U15591 (N_15591,N_9815,N_12370);
or U15592 (N_15592,N_10492,N_10027);
and U15593 (N_15593,N_11235,N_11671);
nand U15594 (N_15594,N_12065,N_9561);
nand U15595 (N_15595,N_11668,N_12453);
and U15596 (N_15596,N_10886,N_10637);
nor U15597 (N_15597,N_12433,N_11068);
and U15598 (N_15598,N_10333,N_12041);
xor U15599 (N_15599,N_10842,N_11221);
and U15600 (N_15600,N_11860,N_12332);
nand U15601 (N_15601,N_11898,N_11357);
nand U15602 (N_15602,N_11655,N_10132);
or U15603 (N_15603,N_9547,N_10949);
nand U15604 (N_15604,N_9533,N_9602);
nor U15605 (N_15605,N_11179,N_11129);
nand U15606 (N_15606,N_10320,N_11402);
nand U15607 (N_15607,N_12171,N_12477);
or U15608 (N_15608,N_9697,N_10968);
nand U15609 (N_15609,N_11116,N_10581);
and U15610 (N_15610,N_11498,N_12023);
nor U15611 (N_15611,N_10746,N_11433);
nand U15612 (N_15612,N_11800,N_12297);
nand U15613 (N_15613,N_10809,N_11314);
nand U15614 (N_15614,N_10209,N_11249);
and U15615 (N_15615,N_10383,N_12487);
and U15616 (N_15616,N_11017,N_10209);
nor U15617 (N_15617,N_11058,N_12238);
and U15618 (N_15618,N_10996,N_10783);
nor U15619 (N_15619,N_11422,N_11237);
nor U15620 (N_15620,N_12298,N_11215);
or U15621 (N_15621,N_10776,N_10875);
or U15622 (N_15622,N_9851,N_11676);
and U15623 (N_15623,N_10754,N_10064);
nand U15624 (N_15624,N_10950,N_9840);
or U15625 (N_15625,N_14910,N_12922);
or U15626 (N_15626,N_13338,N_15423);
and U15627 (N_15627,N_15401,N_14855);
nand U15628 (N_15628,N_15391,N_13277);
nand U15629 (N_15629,N_13599,N_13025);
nor U15630 (N_15630,N_12725,N_13127);
nand U15631 (N_15631,N_13763,N_14919);
xnor U15632 (N_15632,N_14276,N_12849);
xnor U15633 (N_15633,N_13583,N_13051);
nor U15634 (N_15634,N_15101,N_14453);
nor U15635 (N_15635,N_14601,N_13873);
and U15636 (N_15636,N_14637,N_13437);
nand U15637 (N_15637,N_14019,N_13436);
and U15638 (N_15638,N_14670,N_13145);
and U15639 (N_15639,N_15053,N_14828);
and U15640 (N_15640,N_13892,N_12748);
nand U15641 (N_15641,N_13645,N_14007);
nand U15642 (N_15642,N_13094,N_14722);
xor U15643 (N_15643,N_15441,N_14800);
or U15644 (N_15644,N_15308,N_12902);
or U15645 (N_15645,N_14398,N_14716);
nor U15646 (N_15646,N_13435,N_15597);
and U15647 (N_15647,N_12976,N_12925);
xnor U15648 (N_15648,N_13391,N_13691);
or U15649 (N_15649,N_13990,N_14255);
or U15650 (N_15650,N_14363,N_14020);
or U15651 (N_15651,N_13805,N_13114);
nand U15652 (N_15652,N_14188,N_12546);
nand U15653 (N_15653,N_14327,N_14149);
nand U15654 (N_15654,N_13273,N_14227);
nand U15655 (N_15655,N_12531,N_13309);
nor U15656 (N_15656,N_15220,N_15620);
nand U15657 (N_15657,N_14282,N_12993);
nand U15658 (N_15658,N_14901,N_15397);
or U15659 (N_15659,N_13631,N_14411);
nand U15660 (N_15660,N_15532,N_15099);
nor U15661 (N_15661,N_13900,N_13910);
nand U15662 (N_15662,N_13452,N_13070);
nand U15663 (N_15663,N_14711,N_13355);
nor U15664 (N_15664,N_15431,N_13296);
nor U15665 (N_15665,N_14139,N_14617);
nor U15666 (N_15666,N_15306,N_13684);
and U15667 (N_15667,N_15168,N_13155);
and U15668 (N_15668,N_15338,N_14425);
nor U15669 (N_15669,N_14444,N_12973);
and U15670 (N_15670,N_14339,N_14404);
or U15671 (N_15671,N_12550,N_15273);
nand U15672 (N_15672,N_12879,N_15572);
nand U15673 (N_15673,N_14459,N_13264);
or U15674 (N_15674,N_13586,N_15599);
nor U15675 (N_15675,N_13863,N_13383);
or U15676 (N_15676,N_12862,N_14392);
xor U15677 (N_15677,N_14563,N_13701);
or U15678 (N_15678,N_12569,N_13120);
and U15679 (N_15679,N_15267,N_15588);
and U15680 (N_15680,N_14538,N_12833);
nand U15681 (N_15681,N_15602,N_12788);
or U15682 (N_15682,N_13158,N_13405);
nor U15683 (N_15683,N_13749,N_14831);
nand U15684 (N_15684,N_14989,N_14541);
and U15685 (N_15685,N_14235,N_13058);
and U15686 (N_15686,N_14102,N_12974);
nand U15687 (N_15687,N_15547,N_15595);
nand U15688 (N_15688,N_13980,N_12617);
nand U15689 (N_15689,N_14301,N_15038);
xnor U15690 (N_15690,N_14456,N_15089);
nand U15691 (N_15691,N_13074,N_13425);
and U15692 (N_15692,N_14584,N_13585);
nor U15693 (N_15693,N_13231,N_12505);
and U15694 (N_15694,N_14706,N_13332);
nor U15695 (N_15695,N_12909,N_14835);
nand U15696 (N_15696,N_15440,N_14474);
and U15697 (N_15697,N_13546,N_15557);
nor U15698 (N_15698,N_14041,N_12824);
xor U15699 (N_15699,N_14480,N_14079);
and U15700 (N_15700,N_13780,N_15129);
nand U15701 (N_15701,N_13016,N_12627);
nor U15702 (N_15702,N_14649,N_12560);
and U15703 (N_15703,N_14166,N_14844);
nand U15704 (N_15704,N_14635,N_13642);
nand U15705 (N_15705,N_15248,N_15266);
or U15706 (N_15706,N_15536,N_13030);
and U15707 (N_15707,N_15203,N_15198);
and U15708 (N_15708,N_15132,N_13693);
or U15709 (N_15709,N_15243,N_14666);
xnor U15710 (N_15710,N_13854,N_15444);
nand U15711 (N_15711,N_15529,N_15057);
nand U15712 (N_15712,N_14168,N_13682);
nand U15713 (N_15713,N_13596,N_14135);
and U15714 (N_15714,N_12558,N_14894);
nor U15715 (N_15715,N_14050,N_13160);
or U15716 (N_15716,N_12948,N_15206);
nor U15717 (N_15717,N_13232,N_12591);
nor U15718 (N_15718,N_13036,N_12793);
xnor U15719 (N_15719,N_13233,N_15571);
nand U15720 (N_15720,N_12564,N_13415);
or U15721 (N_15721,N_13534,N_12562);
nand U15722 (N_15722,N_12723,N_14730);
nor U15723 (N_15723,N_13125,N_13397);
or U15724 (N_15724,N_14482,N_12586);
nand U15725 (N_15725,N_15347,N_15394);
nor U15726 (N_15726,N_14806,N_14984);
nand U15727 (N_15727,N_15584,N_13786);
and U15728 (N_15728,N_13241,N_13724);
and U15729 (N_15729,N_13941,N_14930);
and U15730 (N_15730,N_12878,N_13518);
or U15731 (N_15731,N_13150,N_14450);
and U15732 (N_15732,N_14509,N_14314);
nand U15733 (N_15733,N_12669,N_13300);
and U15734 (N_15734,N_14122,N_13837);
or U15735 (N_15735,N_12859,N_14898);
or U15736 (N_15736,N_13377,N_15174);
nand U15737 (N_15737,N_14228,N_12871);
nor U15738 (N_15738,N_13845,N_14423);
nor U15739 (N_15739,N_12556,N_13372);
and U15740 (N_15740,N_15442,N_12914);
nor U15741 (N_15741,N_15214,N_12540);
nand U15742 (N_15742,N_13455,N_12806);
nand U15743 (N_15743,N_13199,N_14513);
and U15744 (N_15744,N_13193,N_12514);
nand U15745 (N_15745,N_12903,N_12778);
or U15746 (N_15746,N_13390,N_15615);
and U15747 (N_15747,N_14794,N_14472);
and U15748 (N_15748,N_13832,N_14148);
or U15749 (N_15749,N_12657,N_14183);
and U15750 (N_15750,N_15066,N_13508);
and U15751 (N_15751,N_14832,N_15161);
and U15752 (N_15752,N_14194,N_14257);
nor U15753 (N_15753,N_14333,N_12855);
nand U15754 (N_15754,N_15356,N_13516);
nand U15755 (N_15755,N_15221,N_13381);
or U15756 (N_15756,N_14887,N_15288);
nand U15757 (N_15757,N_13686,N_15560);
or U15758 (N_15758,N_12729,N_14385);
nor U15759 (N_15759,N_14731,N_14893);
or U15760 (N_15760,N_13292,N_14746);
or U15761 (N_15761,N_13821,N_15353);
or U15762 (N_15762,N_14400,N_13625);
nand U15763 (N_15763,N_13023,N_13808);
or U15764 (N_15764,N_14605,N_15201);
or U15765 (N_15765,N_13608,N_14319);
or U15766 (N_15766,N_13616,N_12635);
or U15767 (N_15767,N_12544,N_13592);
nand U15768 (N_15768,N_14325,N_14117);
and U15769 (N_15769,N_12592,N_14749);
and U15770 (N_15770,N_15517,N_13773);
nor U15771 (N_15771,N_12938,N_14049);
and U15772 (N_15772,N_14214,N_13270);
or U15773 (N_15773,N_14738,N_14341);
nand U15774 (N_15774,N_15510,N_13271);
or U15775 (N_15775,N_14998,N_15514);
and U15776 (N_15776,N_13674,N_15540);
nand U15777 (N_15777,N_13593,N_14297);
xnor U15778 (N_15778,N_14209,N_13439);
or U15779 (N_15779,N_12685,N_15351);
and U15780 (N_15780,N_13812,N_15046);
nand U15781 (N_15781,N_12965,N_12554);
or U15782 (N_15782,N_12770,N_15199);
nand U15783 (N_15783,N_13028,N_15128);
xor U15784 (N_15784,N_13422,N_12579);
or U15785 (N_15785,N_13299,N_13267);
nand U15786 (N_15786,N_13429,N_12765);
xor U15787 (N_15787,N_12511,N_12646);
and U15788 (N_15788,N_13846,N_15462);
nor U15789 (N_15789,N_13416,N_15489);
nor U15790 (N_15790,N_14797,N_14084);
or U15791 (N_15791,N_13888,N_14163);
nand U15792 (N_15792,N_14728,N_13820);
or U15793 (N_15793,N_13419,N_14569);
xor U15794 (N_15794,N_14582,N_13612);
nand U15795 (N_15795,N_12769,N_14681);
and U15796 (N_15796,N_13803,N_15387);
nor U15797 (N_15797,N_13964,N_13302);
nor U15798 (N_15798,N_15458,N_15063);
or U15799 (N_15799,N_14184,N_13491);
and U15800 (N_15800,N_14526,N_12864);
nor U15801 (N_15801,N_13122,N_15017);
nand U15802 (N_15802,N_14743,N_13507);
nand U15803 (N_15803,N_13661,N_13263);
nand U15804 (N_15804,N_15265,N_15105);
nor U15805 (N_15805,N_12813,N_15549);
xnor U15806 (N_15806,N_12565,N_14345);
nand U15807 (N_15807,N_15177,N_14066);
or U15808 (N_15808,N_13144,N_15014);
and U15809 (N_15809,N_15190,N_13609);
and U15810 (N_15810,N_13056,N_12843);
or U15811 (N_15811,N_14395,N_15421);
and U15812 (N_15812,N_15433,N_14273);
and U15813 (N_15813,N_12994,N_13456);
nand U15814 (N_15814,N_14885,N_12566);
xor U15815 (N_15815,N_14171,N_15422);
and U15816 (N_15816,N_13359,N_14813);
or U15817 (N_15817,N_14552,N_13191);
nand U15818 (N_15818,N_12929,N_13665);
nand U15819 (N_15819,N_12536,N_15617);
xnor U15820 (N_15820,N_14144,N_12673);
nor U15821 (N_15821,N_15233,N_13620);
or U15822 (N_15822,N_13882,N_15405);
nor U15823 (N_15823,N_14631,N_15133);
or U15824 (N_15824,N_13929,N_13547);
nor U15825 (N_15825,N_13307,N_13444);
and U15826 (N_15826,N_14406,N_14954);
and U15827 (N_15827,N_12670,N_13205);
nor U15828 (N_15828,N_14976,N_12980);
and U15829 (N_15829,N_13240,N_13007);
nand U15830 (N_15830,N_15145,N_15372);
nand U15831 (N_15831,N_13458,N_15260);
nor U15832 (N_15832,N_13528,N_14751);
nor U15833 (N_15833,N_12817,N_15413);
and U15834 (N_15834,N_14527,N_13081);
nand U15835 (N_15835,N_14147,N_14372);
and U15836 (N_15836,N_13370,N_12743);
nor U15837 (N_15837,N_14197,N_13371);
or U15838 (N_15838,N_13079,N_13810);
or U15839 (N_15839,N_13552,N_15496);
and U15840 (N_15840,N_13047,N_14657);
xnor U15841 (N_15841,N_12555,N_14232);
nor U15842 (N_15842,N_15140,N_14119);
or U15843 (N_15843,N_15318,N_13417);
and U15844 (N_15844,N_14000,N_14767);
and U15845 (N_15845,N_13165,N_12692);
and U15846 (N_15846,N_13011,N_14890);
nor U15847 (N_15847,N_15159,N_14931);
nand U15848 (N_15848,N_14781,N_12777);
xnor U15849 (N_15849,N_13269,N_13935);
or U15850 (N_15850,N_14669,N_13113);
nand U15851 (N_15851,N_14988,N_13321);
nand U15852 (N_15852,N_14438,N_12709);
nor U15853 (N_15853,N_14698,N_14925);
nor U15854 (N_15854,N_14597,N_14857);
or U15855 (N_15855,N_14650,N_15217);
xor U15856 (N_15856,N_12798,N_15345);
nand U15857 (N_15857,N_14422,N_13958);
xor U15858 (N_15858,N_13375,N_12549);
or U15859 (N_15859,N_13146,N_14852);
nor U15860 (N_15860,N_14736,N_14229);
nor U15861 (N_15861,N_15426,N_13987);
nor U15862 (N_15862,N_14085,N_13989);
or U15863 (N_15863,N_15485,N_15360);
nor U15864 (N_15864,N_15621,N_14783);
and U15865 (N_15865,N_13636,N_15016);
or U15866 (N_15866,N_14495,N_13380);
nor U15867 (N_15867,N_13221,N_14758);
or U15868 (N_15868,N_13979,N_15279);
or U15869 (N_15869,N_13078,N_15488);
xor U15870 (N_15870,N_14934,N_12986);
nand U15871 (N_15871,N_12757,N_13176);
nand U15872 (N_15872,N_12895,N_13560);
or U15873 (N_15873,N_13339,N_12825);
and U15874 (N_15874,N_12866,N_14330);
and U15875 (N_15875,N_12571,N_15030);
or U15876 (N_15876,N_13274,N_12728);
and U15877 (N_15877,N_13067,N_14496);
nand U15878 (N_15878,N_13513,N_15131);
nand U15879 (N_15879,N_14030,N_13617);
nor U15880 (N_15880,N_15281,N_12889);
nor U15881 (N_15881,N_13450,N_13379);
or U15882 (N_15882,N_14981,N_15169);
or U15883 (N_15883,N_13001,N_15020);
nand U15884 (N_15884,N_14384,N_14487);
nor U15885 (N_15885,N_14130,N_13571);
and U15886 (N_15886,N_14664,N_12619);
xnor U15887 (N_15887,N_13602,N_14512);
and U15888 (N_15888,N_14708,N_15504);
or U15889 (N_15889,N_15611,N_13611);
and U15890 (N_15890,N_14172,N_14285);
nor U15891 (N_15891,N_14942,N_12991);
and U15892 (N_15892,N_13035,N_13476);
and U15893 (N_15893,N_13953,N_14556);
nor U15894 (N_15894,N_14982,N_13836);
xor U15895 (N_15895,N_15270,N_15027);
nor U15896 (N_15896,N_14274,N_14697);
and U15897 (N_15897,N_13503,N_14055);
nor U15898 (N_15898,N_14241,N_14573);
nand U15899 (N_15899,N_15227,N_15180);
and U15900 (N_15900,N_14864,N_13500);
or U15901 (N_15901,N_14607,N_12753);
nand U15902 (N_15902,N_12875,N_14927);
nand U15903 (N_15903,N_14338,N_13121);
nand U15904 (N_15904,N_14468,N_13077);
xnor U15905 (N_15905,N_15088,N_13000);
nor U15906 (N_15906,N_14958,N_12737);
or U15907 (N_15907,N_15494,N_14644);
or U15908 (N_15908,N_12663,N_15268);
nand U15909 (N_15909,N_13947,N_15034);
and U15910 (N_15910,N_15309,N_15204);
nand U15911 (N_15911,N_12921,N_14557);
nor U15912 (N_15912,N_13316,N_15127);
or U15913 (N_15913,N_13874,N_13795);
xnor U15914 (N_15914,N_15558,N_14225);
and U15915 (N_15915,N_13054,N_12677);
nand U15916 (N_15916,N_14719,N_15554);
and U15917 (N_15917,N_14275,N_15025);
nor U15918 (N_15918,N_13248,N_12578);
nand U15919 (N_15919,N_12885,N_14088);
and U15920 (N_15920,N_14303,N_13751);
and U15921 (N_15921,N_12744,N_14410);
or U15922 (N_15922,N_12810,N_14658);
or U15923 (N_15923,N_13209,N_14110);
or U15924 (N_15924,N_12664,N_13652);
or U15925 (N_15925,N_13533,N_13230);
or U15926 (N_15926,N_13069,N_15407);
and U15927 (N_15927,N_15104,N_12881);
xor U15928 (N_15928,N_14647,N_14280);
or U15929 (N_15929,N_12845,N_13341);
nor U15930 (N_15930,N_13920,N_13938);
xnor U15931 (N_15931,N_14865,N_14114);
and U15932 (N_15932,N_14814,N_13531);
and U15933 (N_15933,N_13511,N_15247);
nor U15934 (N_15934,N_13758,N_15241);
nor U15935 (N_15935,N_13861,N_14720);
xnor U15936 (N_15936,N_14881,N_15290);
nand U15937 (N_15937,N_12913,N_15098);
nand U15938 (N_15938,N_13673,N_14175);
nor U15939 (N_15939,N_12772,N_14244);
nand U15940 (N_15940,N_13747,N_13792);
nand U15941 (N_15941,N_13813,N_12874);
xnor U15942 (N_15942,N_13018,N_13662);
or U15943 (N_15943,N_15263,N_12880);
nand U15944 (N_15944,N_12856,N_15090);
nor U15945 (N_15945,N_13214,N_13817);
nor U15946 (N_15946,N_15417,N_13253);
nor U15947 (N_15947,N_15157,N_14393);
or U15948 (N_15948,N_14250,N_14922);
and U15949 (N_15949,N_14037,N_13502);
nor U15950 (N_15950,N_15464,N_13239);
and U15951 (N_15951,N_13843,N_14177);
or U15952 (N_15952,N_14186,N_14036);
nor U15953 (N_15953,N_14845,N_12694);
nor U15954 (N_15954,N_14291,N_14277);
nor U15955 (N_15955,N_13206,N_13746);
or U15956 (N_15956,N_14365,N_14320);
or U15957 (N_15957,N_13957,N_12911);
or U15958 (N_15958,N_14859,N_12930);
and U15959 (N_15959,N_15222,N_13789);
nor U15960 (N_15960,N_13830,N_15236);
or U15961 (N_15961,N_12726,N_13166);
and U15962 (N_15962,N_12924,N_13449);
and U15963 (N_15963,N_14141,N_14022);
nor U15964 (N_15964,N_14078,N_12771);
nand U15965 (N_15965,N_15003,N_14558);
xnor U15966 (N_15966,N_14326,N_13564);
nor U15967 (N_15967,N_14293,N_13988);
and U15968 (N_15968,N_15324,N_15522);
nor U15969 (N_15969,N_13734,N_14065);
and U15970 (N_15970,N_14413,N_12787);
nand U15971 (N_15971,N_12697,N_14245);
nand U15972 (N_15972,N_14642,N_14546);
xor U15973 (N_15973,N_13590,N_13086);
nand U15974 (N_15974,N_13772,N_13124);
or U15975 (N_15975,N_13613,N_14752);
nand U15976 (N_15976,N_14648,N_15479);
nand U15977 (N_15977,N_14471,N_13826);
xnor U15978 (N_15978,N_14010,N_14695);
and U15979 (N_15979,N_13978,N_13304);
nor U15980 (N_15980,N_13699,N_13290);
or U15981 (N_15981,N_13973,N_12671);
and U15982 (N_15982,N_15608,N_13418);
or U15983 (N_15983,N_15533,N_14217);
nand U15984 (N_15984,N_14869,N_13575);
xnor U15985 (N_15985,N_15610,N_13668);
nand U15986 (N_15986,N_14428,N_14279);
nor U15987 (N_15987,N_14021,N_15171);
or U15988 (N_15988,N_13912,N_12768);
and U15989 (N_15989,N_15100,N_13398);
nor U15990 (N_15990,N_14099,N_14770);
xor U15991 (N_15991,N_13965,N_13745);
xor U15992 (N_15992,N_14547,N_14315);
and U15993 (N_15993,N_13658,N_13291);
nor U15994 (N_15994,N_14440,N_12762);
and U15995 (N_15995,N_15587,N_12940);
and U15996 (N_15996,N_13128,N_13913);
or U15997 (N_15997,N_12686,N_14132);
nor U15998 (N_15998,N_14039,N_13393);
nand U15999 (N_15999,N_15342,N_14995);
and U16000 (N_16000,N_14003,N_15299);
or U16001 (N_16001,N_13265,N_13776);
xor U16002 (N_16002,N_13451,N_13557);
xor U16003 (N_16003,N_13457,N_12712);
nand U16004 (N_16004,N_14040,N_13570);
or U16005 (N_16005,N_15253,N_14374);
and U16006 (N_16006,N_13492,N_13565);
and U16007 (N_16007,N_13014,N_12504);
nand U16008 (N_16008,N_13619,N_13423);
nor U16009 (N_16009,N_12854,N_14073);
and U16010 (N_16010,N_12702,N_13713);
or U16011 (N_16011,N_14271,N_14189);
nand U16012 (N_16012,N_12972,N_12958);
or U16013 (N_16013,N_12501,N_15298);
nand U16014 (N_16014,N_13962,N_12735);
nand U16015 (N_16015,N_14957,N_13385);
xnor U16016 (N_16016,N_14801,N_15410);
or U16017 (N_16017,N_13387,N_15228);
nor U16018 (N_16018,N_15415,N_14692);
nor U16019 (N_16019,N_13465,N_12741);
or U16020 (N_16020,N_14101,N_15010);
nand U16021 (N_16021,N_13889,N_12525);
or U16022 (N_16022,N_12648,N_13768);
nand U16023 (N_16023,N_12872,N_14729);
nor U16024 (N_16024,N_13946,N_12513);
nor U16025 (N_16025,N_14784,N_12710);
nand U16026 (N_16026,N_13208,N_14053);
or U16027 (N_16027,N_12632,N_14691);
or U16028 (N_16028,N_13510,N_12755);
and U16029 (N_16029,N_14955,N_14762);
nand U16030 (N_16030,N_14246,N_13945);
xnor U16031 (N_16031,N_14790,N_13972);
nand U16032 (N_16032,N_13410,N_14609);
nor U16033 (N_16033,N_12818,N_13488);
or U16034 (N_16034,N_14242,N_13720);
or U16035 (N_16035,N_15466,N_15289);
or U16036 (N_16036,N_13303,N_14062);
nor U16037 (N_16037,N_13614,N_13196);
and U16038 (N_16038,N_13868,N_14427);
or U16039 (N_16039,N_13680,N_13757);
or U16040 (N_16040,N_12534,N_15028);
xor U16041 (N_16041,N_14771,N_15521);
nand U16042 (N_16042,N_13050,N_15400);
nand U16043 (N_16043,N_13345,N_15552);
or U16044 (N_16044,N_13403,N_14359);
nor U16045 (N_16045,N_15302,N_14048);
and U16046 (N_16046,N_15622,N_14252);
or U16047 (N_16047,N_13885,N_14264);
nand U16048 (N_16048,N_14873,N_14484);
or U16049 (N_16049,N_14505,N_15365);
or U16050 (N_16050,N_15402,N_14560);
or U16051 (N_16051,N_13532,N_13638);
or U16052 (N_16052,N_13936,N_12604);
xor U16053 (N_16053,N_12877,N_15175);
nor U16054 (N_16054,N_13840,N_13402);
nor U16055 (N_16055,N_13970,N_14348);
nand U16056 (N_16056,N_13698,N_12668);
xor U16057 (N_16057,N_13460,N_15370);
or U16058 (N_16058,N_15043,N_14863);
or U16059 (N_16059,N_14507,N_15144);
nand U16060 (N_16060,N_14551,N_15545);
nor U16061 (N_16061,N_12585,N_13222);
xor U16062 (N_16062,N_14778,N_12676);
nor U16063 (N_16063,N_12732,N_15501);
xnor U16064 (N_16064,N_13828,N_12779);
nand U16065 (N_16065,N_15179,N_14952);
and U16066 (N_16066,N_14151,N_15035);
nand U16067 (N_16067,N_15516,N_14860);
nand U16068 (N_16068,N_13259,N_14625);
and U16069 (N_16069,N_14997,N_14307);
nand U16070 (N_16070,N_12807,N_15114);
nor U16071 (N_16071,N_13897,N_14687);
and U16072 (N_16072,N_15600,N_15581);
and U16073 (N_16073,N_15429,N_12791);
or U16074 (N_16074,N_15383,N_12893);
nor U16075 (N_16075,N_14167,N_15395);
xor U16076 (N_16076,N_14023,N_13930);
xnor U16077 (N_16077,N_14170,N_13983);
nor U16078 (N_16078,N_14572,N_13750);
nor U16079 (N_16079,N_13783,N_13388);
and U16080 (N_16080,N_13931,N_13354);
and U16081 (N_16081,N_13759,N_12731);
and U16082 (N_16082,N_14856,N_13672);
nand U16083 (N_16083,N_13781,N_12738);
or U16084 (N_16084,N_14586,N_12522);
and U16085 (N_16085,N_13703,N_14671);
and U16086 (N_16086,N_13907,N_13842);
nor U16087 (N_16087,N_13234,N_15162);
or U16088 (N_16088,N_15254,N_12734);
or U16089 (N_16089,N_14621,N_13791);
nand U16090 (N_16090,N_15613,N_13186);
and U16091 (N_16091,N_12853,N_15346);
or U16092 (N_16092,N_15566,N_14334);
and U16093 (N_16093,N_12838,N_14185);
and U16094 (N_16094,N_14042,N_14858);
xnor U16095 (N_16095,N_12918,N_12713);
and U16096 (N_16096,N_14804,N_14915);
or U16097 (N_16097,N_14533,N_12666);
nand U16098 (N_16098,N_13597,N_15334);
and U16099 (N_16099,N_13347,N_14431);
or U16100 (N_16100,N_13095,N_15321);
nand U16101 (N_16101,N_14929,N_13862);
nor U16102 (N_16102,N_14713,N_14520);
nor U16103 (N_16103,N_13210,N_13389);
nor U16104 (N_16104,N_14435,N_12883);
xor U16105 (N_16105,N_15594,N_15379);
or U16106 (N_16106,N_14027,N_13580);
nor U16107 (N_16107,N_13778,N_14896);
or U16108 (N_16108,N_14260,N_13637);
nor U16109 (N_16109,N_12861,N_14972);
nor U16110 (N_16110,N_12827,N_14834);
or U16111 (N_16111,N_13092,N_12847);
xnor U16112 (N_16112,N_13089,N_13606);
nand U16113 (N_16113,N_12644,N_13715);
or U16114 (N_16114,N_15518,N_14861);
nor U16115 (N_16115,N_14539,N_15508);
or U16116 (N_16116,N_15238,N_13005);
and U16117 (N_16117,N_13649,N_13694);
nand U16118 (N_16118,N_15331,N_14416);
nand U16119 (N_16119,N_12959,N_14786);
nand U16120 (N_16120,N_13486,N_12588);
xor U16121 (N_16121,N_13323,N_13080);
xnor U16122 (N_16122,N_12814,N_13426);
nand U16123 (N_16123,N_13468,N_14061);
nand U16124 (N_16124,N_14205,N_13395);
or U16125 (N_16125,N_12943,N_13342);
nor U16126 (N_16126,N_14418,N_15001);
and U16127 (N_16127,N_14715,N_12634);
or U16128 (N_16128,N_13727,N_15492);
nor U16129 (N_16129,N_12722,N_13536);
or U16130 (N_16130,N_15339,N_14313);
nand U16131 (N_16131,N_13968,N_13112);
and U16132 (N_16132,N_13059,N_13087);
and U16133 (N_16133,N_12506,N_15330);
nor U16134 (N_16134,N_12840,N_12557);
or U16135 (N_16135,N_14689,N_15271);
and U16136 (N_16136,N_14802,N_14300);
nor U16137 (N_16137,N_15539,N_14535);
nor U16138 (N_16138,N_15355,N_13283);
or U16139 (N_16139,N_13107,N_14757);
xnor U16140 (N_16140,N_13003,N_13902);
nor U16141 (N_16141,N_14503,N_14100);
or U16142 (N_16142,N_14294,N_13358);
nor U16143 (N_16143,N_12543,N_15216);
and U16144 (N_16144,N_14408,N_14378);
and U16145 (N_16145,N_12981,N_13102);
nand U16146 (N_16146,N_13006,N_12652);
and U16147 (N_16147,N_15119,N_13040);
nor U16148 (N_16148,N_14529,N_15623);
or U16149 (N_16149,N_12870,N_14630);
and U16150 (N_16150,N_14939,N_14611);
or U16151 (N_16151,N_15392,N_14455);
or U16152 (N_16152,N_12915,N_12961);
or U16153 (N_16153,N_14531,N_13305);
nor U16154 (N_16154,N_14033,N_15231);
nand U16155 (N_16155,N_13519,N_14761);
or U16156 (N_16156,N_14121,N_12816);
nand U16157 (N_16157,N_14222,N_13601);
nand U16158 (N_16158,N_15574,N_15497);
and U16159 (N_16159,N_15320,N_12804);
and U16160 (N_16160,N_13903,N_14827);
or U16161 (N_16161,N_14707,N_13204);
nand U16162 (N_16162,N_14397,N_15437);
nor U16163 (N_16163,N_13041,N_15296);
or U16164 (N_16164,N_12615,N_14200);
or U16165 (N_16165,N_14819,N_14093);
or U16166 (N_16166,N_15548,N_14745);
nor U16167 (N_16167,N_15457,N_14986);
nor U16168 (N_16168,N_13870,N_13262);
or U16169 (N_16169,N_15195,N_14543);
xnor U16170 (N_16170,N_14867,N_14094);
nor U16171 (N_16171,N_14109,N_15576);
xnor U16172 (N_16172,N_15323,N_14795);
nor U16173 (N_16173,N_13085,N_13174);
xor U16174 (N_16174,N_14561,N_14879);
or U16175 (N_16175,N_14965,N_14268);
and U16176 (N_16176,N_14992,N_15065);
nor U16177 (N_16177,N_13841,N_14848);
or U16178 (N_16178,N_13877,N_15412);
xnor U16179 (N_16179,N_13117,N_15196);
nand U16180 (N_16180,N_13866,N_15167);
nand U16181 (N_16181,N_14299,N_14220);
or U16182 (N_16182,N_13245,N_15023);
nor U16183 (N_16183,N_14394,N_12637);
nor U16184 (N_16184,N_14096,N_13237);
and U16185 (N_16185,N_15122,N_13138);
nand U16186 (N_16186,N_14463,N_12581);
and U16187 (N_16187,N_15537,N_15008);
and U16188 (N_16188,N_13236,N_14152);
xnor U16189 (N_16189,N_15004,N_13850);
nand U16190 (N_16190,N_13105,N_15121);
nor U16191 (N_16191,N_13272,N_12721);
nor U16192 (N_16192,N_13581,N_13838);
or U16193 (N_16193,N_15050,N_15240);
nor U16194 (N_16194,N_14136,N_15586);
and U16195 (N_16195,N_13771,N_13522);
or U16196 (N_16196,N_12678,N_14705);
nor U16197 (N_16197,N_15303,N_13017);
or U16198 (N_16198,N_13297,N_14368);
nor U16199 (N_16199,N_15352,N_14026);
nor U16200 (N_16200,N_14936,N_13275);
and U16201 (N_16201,N_15341,N_13242);
nor U16202 (N_16202,N_13010,N_13899);
nand U16203 (N_16203,N_14581,N_12829);
and U16204 (N_16204,N_13676,N_14310);
or U16205 (N_16205,N_13667,N_15385);
nor U16206 (N_16206,N_14724,N_14914);
and U16207 (N_16207,N_13555,N_15278);
nor U16208 (N_16208,N_13223,N_15432);
and U16209 (N_16209,N_13632,N_13173);
nor U16210 (N_16210,N_13906,N_15310);
nor U16211 (N_16211,N_13554,N_13977);
xor U16212 (N_16212,N_12538,N_13481);
or U16213 (N_16213,N_13433,N_13100);
or U16214 (N_16214,N_14514,N_15060);
and U16215 (N_16215,N_12700,N_13670);
xor U16216 (N_16216,N_12628,N_14847);
nor U16217 (N_16217,N_13363,N_15287);
nor U16218 (N_16218,N_12541,N_15120);
nand U16219 (N_16219,N_14951,N_14306);
and U16220 (N_16220,N_15115,N_12898);
or U16221 (N_16221,N_14710,N_12587);
nor U16222 (N_16222,N_14116,N_13558);
nor U16223 (N_16223,N_12809,N_12799);
xor U16224 (N_16224,N_12933,N_13760);
xor U16225 (N_16225,N_14811,N_13368);
nor U16226 (N_16226,N_15388,N_12621);
nor U16227 (N_16227,N_14355,N_13443);
xor U16228 (N_16228,N_12764,N_14344);
or U16229 (N_16229,N_15482,N_13756);
nand U16230 (N_16230,N_14933,N_13950);
nand U16231 (N_16231,N_13995,N_13136);
or U16232 (N_16232,N_15062,N_12733);
nand U16233 (N_16233,N_14295,N_14842);
or U16234 (N_16234,N_12888,N_15565);
nor U16235 (N_16235,N_14755,N_13483);
or U16236 (N_16236,N_13579,N_15601);
and U16237 (N_16237,N_14994,N_15084);
or U16238 (N_16238,N_13951,N_15561);
and U16239 (N_16239,N_13689,N_13033);
nor U16240 (N_16240,N_14838,N_14401);
nor U16241 (N_16241,N_13521,N_14908);
and U16242 (N_16242,N_13349,N_13411);
nand U16243 (N_16243,N_15048,N_13331);
nor U16244 (N_16244,N_13217,N_14328);
and U16245 (N_16245,N_14287,N_15332);
nor U16246 (N_16246,N_12610,N_12518);
xor U16247 (N_16247,N_15439,N_14773);
nor U16248 (N_16248,N_13804,N_15246);
xor U16249 (N_16249,N_13220,N_14824);
or U16250 (N_16250,N_13847,N_14960);
nand U16251 (N_16251,N_12693,N_14791);
nor U16252 (N_16252,N_13523,N_12850);
xnor U16253 (N_16253,N_14764,N_14387);
or U16254 (N_16254,N_13190,N_13061);
nand U16255 (N_16255,N_14598,N_15262);
nand U16256 (N_16256,N_13711,N_15172);
and U16257 (N_16257,N_13099,N_13177);
nor U16258 (N_16258,N_14763,N_12599);
nor U16259 (N_16259,N_12561,N_14656);
nor U16260 (N_16260,N_14491,N_15230);
nand U16261 (N_16261,N_15052,N_13034);
nand U16262 (N_16262,N_12957,N_12756);
nor U16263 (N_16263,N_13905,N_13432);
or U16264 (N_16264,N_14946,N_12631);
or U16265 (N_16265,N_15007,N_14875);
nand U16266 (N_16266,N_14153,N_14466);
xor U16267 (N_16267,N_14343,N_14545);
or U16268 (N_16268,N_13741,N_13640);
nand U16269 (N_16269,N_13604,N_15209);
or U16270 (N_16270,N_15478,N_13811);
and U16271 (N_16271,N_15512,N_14074);
nor U16272 (N_16272,N_13430,N_14938);
nor U16273 (N_16273,N_14253,N_13188);
nand U16274 (N_16274,N_13256,N_13055);
nor U16275 (N_16275,N_15282,N_15139);
xor U16276 (N_16276,N_13948,N_15619);
nand U16277 (N_16277,N_13994,N_13201);
nor U16278 (N_16278,N_14045,N_13194);
or U16279 (N_16279,N_12608,N_14685);
nand U16280 (N_16280,N_15185,N_13911);
nand U16281 (N_16281,N_12629,N_15200);
xor U16282 (N_16282,N_14211,N_12519);
or U16283 (N_16283,N_13848,N_12868);
xnor U16284 (N_16284,N_12595,N_13104);
nor U16285 (N_16285,N_13921,N_13497);
or U16286 (N_16286,N_14447,N_13487);
nor U16287 (N_16287,N_13004,N_15445);
and U16288 (N_16288,N_15317,N_13603);
or U16289 (N_16289,N_14159,N_14377);
nand U16290 (N_16290,N_13677,N_14193);
nor U16291 (N_16291,N_12873,N_15456);
and U16292 (N_16292,N_13819,N_12790);
and U16293 (N_16293,N_12526,N_14473);
nand U16294 (N_16294,N_12695,N_15118);
nor U16295 (N_16295,N_13706,N_12969);
and U16296 (N_16296,N_12912,N_14308);
or U16297 (N_16297,N_14935,N_13301);
nor U16298 (N_16298,N_12907,N_14849);
nand U16299 (N_16299,N_15047,N_12999);
and U16300 (N_16300,N_14415,N_15403);
nand U16301 (N_16301,N_14850,N_13287);
nor U16302 (N_16302,N_14674,N_15555);
or U16303 (N_16303,N_13707,N_15258);
nor U16304 (N_16304,N_14445,N_12796);
nand U16305 (N_16305,N_14682,N_14361);
nand U16306 (N_16306,N_14980,N_15108);
or U16307 (N_16307,N_15390,N_14095);
nor U16308 (N_16308,N_13514,N_14288);
nand U16309 (N_16309,N_14080,N_12891);
nand U16310 (N_16310,N_15322,N_13482);
nand U16311 (N_16311,N_13740,N_14311);
or U16312 (N_16312,N_13688,N_13442);
and U16313 (N_16313,N_14479,N_12842);
or U16314 (N_16314,N_13876,N_15364);
nand U16315 (N_16315,N_15036,N_14382);
nor U16316 (N_16316,N_12763,N_14249);
and U16317 (N_16317,N_14360,N_14578);
nand U16318 (N_16318,N_15256,N_12786);
or U16319 (N_16319,N_12679,N_13624);
and U16320 (N_16320,N_15202,N_13446);
nor U16321 (N_16321,N_12899,N_15451);
nor U16322 (N_16322,N_14833,N_13728);
nor U16323 (N_16323,N_13883,N_14403);
or U16324 (N_16324,N_15019,N_12992);
nand U16325 (N_16325,N_12820,N_15575);
nand U16326 (N_16326,N_14588,N_15252);
and U16327 (N_16327,N_13551,N_15420);
nand U16328 (N_16328,N_14477,N_14086);
nor U16329 (N_16329,N_15283,N_12740);
nand U16330 (N_16330,N_15244,N_13044);
nor U16331 (N_16331,N_13156,N_13901);
or U16332 (N_16332,N_13284,N_14470);
nor U16333 (N_16333,N_13943,N_13101);
nor U16334 (N_16334,N_14038,N_12978);
or U16335 (N_16335,N_15404,N_12935);
nor U16336 (N_16336,N_15189,N_15436);
or U16337 (N_16337,N_15304,N_14964);
and U16338 (N_16338,N_14069,N_15211);
or U16339 (N_16339,N_13556,N_12714);
nor U16340 (N_16340,N_15480,N_13428);
and U16341 (N_16341,N_13879,N_13063);
or U16342 (N_16342,N_12523,N_13225);
and U16343 (N_16343,N_15312,N_14165);
and U16344 (N_16344,N_12782,N_15234);
xnor U16345 (N_16345,N_14478,N_13986);
nor U16346 (N_16346,N_15305,N_13961);
and U16347 (N_16347,N_13573,N_14131);
nor U16348 (N_16348,N_15146,N_13769);
and U16349 (N_16349,N_13710,N_14467);
nor U16350 (N_16350,N_14638,N_13037);
and U16351 (N_16351,N_12730,N_13373);
nand U16352 (N_16352,N_15344,N_13447);
nand U16353 (N_16353,N_13814,N_13400);
and U16354 (N_16354,N_13329,N_15335);
or U16355 (N_16355,N_14646,N_14145);
nor U16356 (N_16356,N_14882,N_12647);
or U16357 (N_16357,N_15011,N_14999);
or U16358 (N_16358,N_13312,N_15465);
xnor U16359 (N_16359,N_14349,N_14199);
or U16360 (N_16360,N_12984,N_14777);
nor U16361 (N_16361,N_15018,N_13227);
nor U16362 (N_16362,N_14375,N_14870);
nor U16363 (N_16363,N_15166,N_15382);
nand U16364 (N_16364,N_13927,N_14123);
xor U16365 (N_16365,N_13414,N_13412);
nand U16366 (N_16366,N_12720,N_13386);
and U16367 (N_16367,N_14178,N_13052);
and U16368 (N_16368,N_12509,N_14712);
nand U16369 (N_16369,N_13909,N_14923);
and U16370 (N_16370,N_14906,N_12836);
nor U16371 (N_16371,N_14693,N_15181);
and U16372 (N_16372,N_14688,N_13021);
or U16373 (N_16373,N_13438,N_13499);
and U16374 (N_16374,N_14125,N_14107);
or U16375 (N_16375,N_15580,N_14747);
nor U16376 (N_16376,N_13679,N_15039);
or U16377 (N_16377,N_13914,N_15068);
nor U16378 (N_16378,N_12917,N_15473);
or U16379 (N_16379,N_14880,N_13647);
or U16380 (N_16380,N_14971,N_15605);
nand U16381 (N_16381,N_13501,N_15430);
xor U16382 (N_16382,N_13115,N_14510);
nand U16383 (N_16383,N_13731,N_12659);
nand U16384 (N_16384,N_13408,N_15438);
or U16385 (N_16385,N_14155,N_13790);
nand U16386 (N_16386,N_14519,N_13923);
xor U16387 (N_16387,N_13175,N_14645);
or U16388 (N_16388,N_13134,N_14433);
nor U16389 (N_16389,N_15037,N_15551);
and U16390 (N_16390,N_14500,N_14146);
and U16391 (N_16391,N_12502,N_14718);
and U16392 (N_16392,N_14843,N_12937);
or U16393 (N_16393,N_14553,N_13932);
nand U16394 (N_16394,N_15092,N_14434);
or U16395 (N_16395,N_15081,N_14353);
nand U16396 (N_16396,N_13984,N_14632);
nand U16397 (N_16397,N_14296,N_13915);
xnor U16398 (N_16398,N_14158,N_14805);
or U16399 (N_16399,N_15328,N_14044);
nor U16400 (N_16400,N_13770,N_15472);
and U16401 (N_16401,N_14462,N_12609);
xor U16402 (N_16402,N_13477,N_15124);
or U16403 (N_16403,N_14540,N_14072);
nor U16404 (N_16404,N_14818,N_14821);
nand U16405 (N_16405,N_14665,N_13461);
nand U16406 (N_16406,N_12890,N_12985);
or U16407 (N_16407,N_14059,N_15374);
and U16408 (N_16408,N_14004,N_14017);
or U16409 (N_16409,N_14396,N_13974);
nand U16410 (N_16410,N_15326,N_12691);
and U16411 (N_16411,N_15543,N_14900);
or U16412 (N_16412,N_14945,N_14641);
nand U16413 (N_16413,N_13288,N_12801);
nor U16414 (N_16414,N_14201,N_12739);
nor U16415 (N_16415,N_14013,N_13954);
nor U16416 (N_16416,N_13512,N_14263);
or U16417 (N_16417,N_15515,N_13855);
xnor U16418 (N_16418,N_14134,N_15064);
nand U16419 (N_16419,N_12758,N_13473);
and U16420 (N_16420,N_15612,N_14124);
nor U16421 (N_16421,N_15087,N_14947);
or U16422 (N_16422,N_13306,N_13224);
or U16423 (N_16423,N_13111,N_13926);
and U16424 (N_16424,N_14494,N_12780);
nor U16425 (N_16425,N_12649,N_14236);
and U16426 (N_16426,N_13610,N_13195);
nand U16427 (N_16427,N_14810,N_12905);
or U16428 (N_16428,N_13925,N_14735);
nor U16429 (N_16429,N_14324,N_15005);
or U16430 (N_16430,N_15237,N_14057);
or U16431 (N_16431,N_15012,N_14699);
and U16432 (N_16432,N_14347,N_14595);
and U16433 (N_16433,N_14985,N_13949);
nand U16434 (N_16434,N_14179,N_15307);
nor U16435 (N_16435,N_12547,N_12711);
nand U16436 (N_16436,N_13966,N_13607);
nand U16437 (N_16437,N_14941,N_13761);
and U16438 (N_16438,N_15072,N_14663);
nand U16439 (N_16439,N_15021,N_13022);
xor U16440 (N_16440,N_15173,N_14991);
xnor U16441 (N_16441,N_15194,N_14481);
or U16442 (N_16442,N_12822,N_13801);
nor U16443 (N_16443,N_12812,N_13462);
nand U16444 (N_16444,N_13765,N_12696);
nand U16445 (N_16445,N_13895,N_13258);
and U16446 (N_16446,N_12987,N_12951);
xor U16447 (N_16447,N_14606,N_14518);
and U16448 (N_16448,N_12956,N_12655);
nor U16449 (N_16449,N_14161,N_15042);
nand U16450 (N_16450,N_15507,N_12953);
nor U16451 (N_16451,N_14304,N_14614);
or U16452 (N_16452,N_14610,N_12687);
nand U16453 (N_16453,N_15269,N_14732);
or U16454 (N_16454,N_15085,N_15205);
or U16455 (N_16455,N_13360,N_12602);
nand U16456 (N_16456,N_13969,N_12606);
or U16457 (N_16457,N_14812,N_13090);
and U16458 (N_16458,N_14542,N_12749);
and U16459 (N_16459,N_15376,N_12901);
nor U16460 (N_16460,N_14029,N_12594);
and U16461 (N_16461,N_15604,N_13330);
nand U16462 (N_16462,N_13027,N_12688);
or U16463 (N_16463,N_15276,N_14223);
or U16464 (N_16464,N_14600,N_12852);
and U16465 (N_16465,N_14202,N_14449);
nand U16466 (N_16466,N_13687,N_13441);
nand U16467 (N_16467,N_13281,N_14574);
nor U16468 (N_16468,N_13207,N_15232);
xor U16469 (N_16469,N_14460,N_13340);
nand U16470 (N_16470,N_15272,N_12783);
nand U16471 (N_16471,N_14231,N_12563);
and U16472 (N_16472,N_13197,N_15461);
or U16473 (N_16473,N_13181,N_14673);
or U16474 (N_16474,N_14809,N_15363);
xnor U16475 (N_16475,N_15490,N_12717);
nor U16476 (N_16476,N_12750,N_12989);
nand U16477 (N_16477,N_13695,N_12882);
and U16478 (N_16478,N_14622,N_12575);
nand U16479 (N_16479,N_13796,N_15300);
or U16480 (N_16480,N_14744,N_13189);
and U16481 (N_16481,N_14679,N_13285);
nand U16482 (N_16482,N_13542,N_12896);
nand U16483 (N_16483,N_14469,N_15075);
xnor U16484 (N_16484,N_13336,N_12596);
nand U16485 (N_16485,N_15154,N_14181);
and U16486 (N_16486,N_14369,N_14068);
and U16487 (N_16487,N_12623,N_13244);
nor U16488 (N_16488,N_14741,N_13179);
nand U16489 (N_16489,N_14937,N_15210);
nand U16490 (N_16490,N_14577,N_13666);
and U16491 (N_16491,N_13569,N_14846);
and U16492 (N_16492,N_14911,N_14417);
or U16493 (N_16493,N_13709,N_15583);
or U16494 (N_16494,N_15455,N_12539);
nand U16495 (N_16495,N_13043,N_13159);
nor U16496 (N_16496,N_13325,N_14677);
nand U16497 (N_16497,N_14702,N_15176);
nor U16498 (N_16498,N_15369,N_15449);
nor U16499 (N_16499,N_13993,N_14366);
nor U16500 (N_16500,N_15106,N_14789);
nor U16501 (N_16501,N_14009,N_13498);
or U16502 (N_16502,N_12797,N_14346);
nand U16503 (N_16503,N_13659,N_12802);
nand U16504 (N_16504,N_13739,N_14696);
or U16505 (N_16505,N_12900,N_14316);
and U16506 (N_16506,N_13294,N_15002);
or U16507 (N_16507,N_14515,N_14443);
or U16508 (N_16508,N_14091,N_14977);
nand U16509 (N_16509,N_14913,N_12927);
nor U16510 (N_16510,N_15524,N_15384);
and U16511 (N_16511,N_13849,N_15213);
nor U16512 (N_16512,N_15556,N_13149);
nand U16513 (N_16513,N_13143,N_12908);
and U16514 (N_16514,N_15418,N_14195);
or U16515 (N_16515,N_13568,N_14137);
nand U16516 (N_16516,N_15251,N_13816);
nor U16517 (N_16517,N_13183,N_14567);
nor U16518 (N_16518,N_15523,N_14337);
and U16519 (N_16519,N_12636,N_15377);
or U16520 (N_16520,N_15592,N_12574);
and U16521 (N_16521,N_14256,N_13545);
nand U16522 (N_16522,N_12897,N_13238);
nand U16523 (N_16523,N_12653,N_13337);
nor U16524 (N_16524,N_14426,N_14892);
nand U16525 (N_16525,N_14207,N_14379);
or U16526 (N_16526,N_14651,N_13584);
or U16527 (N_16527,N_12745,N_13748);
and U16528 (N_16528,N_12815,N_13937);
nor U16529 (N_16529,N_15411,N_14917);
or U16530 (N_16530,N_13348,N_14016);
nand U16531 (N_16531,N_13266,N_14424);
xnor U16532 (N_16532,N_14373,N_13320);
and U16533 (N_16533,N_14769,N_12520);
xor U16534 (N_16534,N_13917,N_12576);
nor U16535 (N_16535,N_15409,N_14815);
or U16536 (N_16536,N_13123,N_14653);
nand U16537 (N_16537,N_14414,N_12559);
nor U16538 (N_16538,N_14442,N_13716);
and U16539 (N_16539,N_12705,N_15152);
and U16540 (N_16540,N_15123,N_13916);
nor U16541 (N_16541,N_13737,N_13057);
and U16542 (N_16542,N_12704,N_14888);
or U16543 (N_16543,N_13406,N_14874);
or U16544 (N_16544,N_15563,N_13187);
nand U16545 (N_16545,N_14129,N_14364);
xnor U16546 (N_16546,N_14070,N_14949);
and U16547 (N_16547,N_13623,N_13243);
or U16548 (N_16548,N_15484,N_13356);
xor U16549 (N_16549,N_14570,N_14005);
nor U16550 (N_16550,N_12719,N_14792);
nand U16551 (N_16551,N_14523,N_13153);
and U16552 (N_16552,N_15280,N_15083);
nor U16553 (N_16553,N_15045,N_13683);
nand U16554 (N_16554,N_13072,N_13249);
xnor U16555 (N_16555,N_14549,N_13235);
nor U16556 (N_16556,N_13959,N_15223);
nor U16557 (N_16557,N_12766,N_14596);
or U16558 (N_16558,N_14192,N_15151);
nand U16559 (N_16559,N_14261,N_14221);
or U16560 (N_16560,N_13574,N_13777);
or U16561 (N_16561,N_12660,N_14680);
or U16562 (N_16562,N_13343,N_13960);
nor U16563 (N_16563,N_12633,N_13646);
xnor U16564 (N_16564,N_14258,N_14083);
nor U16565 (N_16565,N_13908,N_14475);
nand U16566 (N_16566,N_13470,N_13818);
or U16567 (N_16567,N_13009,N_13137);
xor U16568 (N_16568,N_14312,N_15264);
and U16569 (N_16569,N_12945,N_13129);
and U16570 (N_16570,N_13293,N_12583);
nand U16571 (N_16571,N_13543,N_15313);
or U16572 (N_16572,N_14562,N_13797);
or U16573 (N_16573,N_12781,N_14522);
or U16574 (N_16574,N_14226,N_14918);
or U16575 (N_16575,N_14613,N_12512);
and U16576 (N_16576,N_14592,N_14787);
and U16577 (N_16577,N_13282,N_15562);
or U16578 (N_16578,N_14340,N_14218);
or U16579 (N_16579,N_13815,N_14409);
nand U16580 (N_16580,N_12622,N_12952);
and U16581 (N_16581,N_13494,N_13762);
or U16582 (N_16582,N_13517,N_14975);
nand U16583 (N_16583,N_12593,N_14097);
and U16584 (N_16584,N_12742,N_14278);
nor U16585 (N_16585,N_15080,N_14499);
nand U16586 (N_16586,N_12651,N_13045);
nor U16587 (N_16587,N_13424,N_14461);
nand U16588 (N_16588,N_13226,N_12703);
or U16589 (N_16589,N_14269,N_14105);
nand U16590 (N_16590,N_12954,N_12851);
nand U16591 (N_16591,N_13335,N_14265);
or U16592 (N_16592,N_13871,N_14286);
and U16593 (N_16593,N_12776,N_14608);
and U16594 (N_16594,N_12998,N_15130);
nor U16595 (N_16595,N_13504,N_14615);
or U16596 (N_16596,N_14643,N_14517);
xor U16597 (N_16597,N_14302,N_13992);
nor U16598 (N_16598,N_12983,N_14357);
nand U16599 (N_16599,N_15559,N_12682);
nor U16600 (N_16600,N_14654,N_12532);
nor U16601 (N_16601,N_14871,N_15054);
or U16602 (N_16602,N_12654,N_13434);
or U16603 (N_16603,N_15568,N_15235);
or U16604 (N_16604,N_13520,N_14909);
nor U16605 (N_16605,N_13634,N_13807);
or U16606 (N_16606,N_15366,N_14904);
or U16607 (N_16607,N_14210,N_12630);
and U16608 (N_16608,N_14234,N_15567);
and U16609 (N_16609,N_13103,N_15301);
nand U16610 (N_16610,N_14979,N_14142);
and U16611 (N_16611,N_12548,N_14926);
nand U16612 (N_16612,N_12684,N_15325);
and U16613 (N_16613,N_13376,N_15109);
nand U16614 (N_16614,N_14554,N_15315);
and U16615 (N_16615,N_13696,N_14889);
nand U16616 (N_16616,N_13806,N_15474);
or U16617 (N_16617,N_12517,N_15358);
and U16618 (N_16618,N_14564,N_14962);
nor U16619 (N_16619,N_14247,N_14067);
nand U16620 (N_16620,N_12643,N_13038);
nand U16621 (N_16621,N_14281,N_12928);
or U16622 (N_16622,N_14162,N_13215);
and U16623 (N_16623,N_14133,N_12752);
xnor U16624 (N_16624,N_13878,N_12577);
nor U16625 (N_16625,N_13352,N_14948);
nor U16626 (N_16626,N_12774,N_14659);
or U16627 (N_16627,N_13148,N_12516);
and U16628 (N_16628,N_13735,N_14489);
xnor U16629 (N_16629,N_12761,N_12612);
nand U16630 (N_16630,N_12839,N_14089);
or U16631 (N_16631,N_12715,N_14448);
nand U16632 (N_16632,N_13702,N_13421);
nand U16633 (N_16633,N_14354,N_15135);
nor U16634 (N_16634,N_14943,N_15343);
nor U16635 (N_16635,N_12707,N_15094);
or U16636 (N_16636,N_15511,N_13644);
or U16637 (N_16637,N_13857,N_14701);
xor U16638 (N_16638,N_15593,N_14973);
or U16639 (N_16639,N_13648,N_14534);
and U16640 (N_16640,N_12841,N_15477);
nor U16641 (N_16641,N_13753,N_14950);
or U16642 (N_16642,N_13362,N_15375);
and U16643 (N_16643,N_13216,N_14239);
nand U16644 (N_16644,N_13279,N_13577);
or U16645 (N_16645,N_14604,N_14213);
nand U16646 (N_16646,N_14150,N_13685);
and U16647 (N_16647,N_13744,N_14905);
and U16648 (N_16648,N_14322,N_14511);
or U16649 (N_16649,N_14807,N_12865);
nor U16650 (N_16650,N_13132,N_14429);
nand U16651 (N_16651,N_14497,N_13280);
nor U16652 (N_16652,N_14868,N_12910);
or U16653 (N_16653,N_15354,N_13399);
and U16654 (N_16654,N_14779,N_14825);
xnor U16655 (N_16655,N_13084,N_14970);
nand U16656 (N_16656,N_13378,N_12625);
nor U16657 (N_16657,N_12528,N_14386);
nand U16658 (N_16658,N_14829,N_13971);
nand U16659 (N_16659,N_13322,N_14837);
and U16660 (N_16660,N_12831,N_14154);
nor U16661 (N_16661,N_15503,N_12916);
and U16662 (N_16662,N_13490,N_13328);
nor U16663 (N_16663,N_13012,N_12614);
or U16664 (N_16664,N_13708,N_15183);
nor U16665 (N_16665,N_13615,N_14580);
or U16666 (N_16666,N_14748,N_14987);
or U16667 (N_16667,N_15125,N_15525);
nor U16668 (N_16668,N_12582,N_13723);
and U16669 (N_16669,N_13448,N_12754);
and U16670 (N_16670,N_12527,N_15218);
nand U16671 (N_16671,N_12661,N_15491);
and U16672 (N_16672,N_14907,N_13867);
nand U16673 (N_16673,N_13904,N_15239);
and U16674 (N_16674,N_15015,N_14090);
or U16675 (N_16675,N_15542,N_15414);
nor U16676 (N_16676,N_14672,N_13982);
and U16677 (N_16677,N_14571,N_12701);
or U16678 (N_16678,N_13934,N_13212);
nor U16679 (N_16679,N_12886,N_13944);
and U16680 (N_16680,N_12674,N_13809);
or U16681 (N_16681,N_13890,N_15164);
nand U16682 (N_16682,N_14169,N_13141);
or U16683 (N_16683,N_14978,N_13939);
and U16684 (N_16684,N_12828,N_15073);
nor U16685 (N_16685,N_14897,N_13202);
and U16686 (N_16686,N_12795,N_13764);
or U16687 (N_16687,N_14884,N_13257);
xor U16688 (N_16688,N_13167,N_15591);
nor U16689 (N_16689,N_15535,N_13130);
or U16690 (N_16690,N_13655,N_14932);
and U16691 (N_16691,N_15408,N_14633);
or U16692 (N_16692,N_13639,N_15530);
and U16693 (N_16693,N_14187,N_14823);
nor U16694 (N_16694,N_15000,N_13663);
xnor U16695 (N_16695,N_15359,N_13382);
xor U16696 (N_16696,N_13109,N_13169);
and U16697 (N_16697,N_14270,N_13198);
nor U16698 (N_16698,N_14590,N_13839);
or U16699 (N_16699,N_12826,N_14230);
and U16700 (N_16700,N_15070,N_13471);
nand U16701 (N_16701,N_15013,N_15138);
nand U16702 (N_16702,N_13489,N_15097);
nor U16703 (N_16703,N_12699,N_13656);
and U16704 (N_16704,N_14996,N_12931);
nand U16705 (N_16705,N_13822,N_14902);
or U16706 (N_16706,N_12867,N_12667);
nor U16707 (N_16707,N_13042,N_15357);
nand U16708 (N_16708,N_13525,N_14830);
or U16709 (N_16709,N_13071,N_15495);
nand U16710 (N_16710,N_15368,N_14966);
nor U16711 (N_16711,N_14490,N_14331);
and U16712 (N_16712,N_15091,N_14714);
and U16713 (N_16713,N_13918,N_13324);
and U16714 (N_16714,N_13535,N_14628);
or U16715 (N_16715,N_12690,N_14536);
or U16716 (N_16716,N_14104,N_15624);
nand U16717 (N_16717,N_14483,N_15577);
nand U16718 (N_16718,N_15229,N_13785);
nor U16719 (N_16719,N_13697,N_12934);
or U16720 (N_16720,N_13725,N_15316);
and U16721 (N_16721,N_14391,N_15399);
nor U16722 (N_16722,N_14953,N_13999);
xor U16723 (N_16723,N_13743,N_14112);
or U16724 (N_16724,N_13184,N_13651);
xnor U16725 (N_16725,N_14421,N_13247);
xnor U16726 (N_16726,N_13108,N_15049);
and U16727 (N_16727,N_15606,N_13161);
and U16728 (N_16728,N_15163,N_14903);
or U16729 (N_16729,N_13131,N_14128);
nor U16730 (N_16730,N_14993,N_13333);
nor U16731 (N_16731,N_12680,N_13392);
nand U16732 (N_16732,N_14587,N_12767);
nand U16733 (N_16733,N_13566,N_15031);
and U16734 (N_16734,N_12638,N_15327);
xnor U16735 (N_16735,N_13013,N_14785);
and U16736 (N_16736,N_13046,N_14772);
nor U16737 (N_16737,N_13924,N_13200);
nand U16738 (N_16738,N_14052,N_14678);
and U16739 (N_16739,N_14766,N_13509);
nor U16740 (N_16740,N_13172,N_13480);
and U16741 (N_16741,N_14103,N_14028);
xor U16742 (N_16742,N_14001,N_13853);
and U16743 (N_16743,N_13261,N_12553);
nor U16744 (N_16744,N_15470,N_13752);
nor U16745 (N_16745,N_14899,N_13823);
nand U16746 (N_16746,N_15137,N_14756);
nand U16747 (N_16747,N_13367,N_13154);
or U16748 (N_16748,N_12535,N_14694);
nor U16749 (N_16749,N_15044,N_13633);
or U16750 (N_16750,N_14317,N_15427);
and U16751 (N_16751,N_15111,N_15476);
nand U16752 (N_16752,N_14524,N_14676);
nand U16753 (N_16753,N_15569,N_13872);
nand U16754 (N_16754,N_13048,N_13318);
nand U16755 (N_16755,N_15182,N_12611);
nor U16756 (N_16756,N_13774,N_14272);
and U16757 (N_16757,N_15607,N_15509);
and U16758 (N_16758,N_14782,N_14626);
or U16759 (N_16759,N_14332,N_13859);
nand U16760 (N_16760,N_15284,N_13278);
nand U16761 (N_16761,N_15531,N_13454);
or U16762 (N_16762,N_12946,N_15156);
and U16763 (N_16763,N_14959,N_14537);
and U16764 (N_16764,N_12641,N_15149);
or U16765 (N_16765,N_13928,N_15520);
or U16766 (N_16766,N_15443,N_12567);
nor U16767 (N_16767,N_13420,N_12573);
nand U16768 (N_16768,N_13286,N_13062);
xnor U16769 (N_16769,N_14668,N_13719);
nor U16770 (N_16770,N_14383,N_15459);
xor U16771 (N_16771,N_13825,N_13015);
nor U16772 (N_16772,N_14208,N_13985);
or U16773 (N_16773,N_15618,N_15396);
nand U16774 (N_16774,N_13991,N_15193);
nand U16775 (N_16775,N_14768,N_12971);
nor U16776 (N_16776,N_15032,N_14974);
nor U16777 (N_16777,N_12500,N_13587);
nor U16778 (N_16778,N_15147,N_14820);
and U16779 (N_16779,N_13162,N_13505);
nand U16780 (N_16780,N_13782,N_13692);
and U16781 (N_16781,N_13031,N_15033);
and U16782 (N_16782,N_13779,N_14636);
or U16783 (N_16783,N_13976,N_13567);
nand U16784 (N_16784,N_13967,N_14594);
nor U16785 (N_16785,N_13118,N_14111);
or U16786 (N_16786,N_13893,N_15250);
and U16787 (N_16787,N_13880,N_14655);
and U16788 (N_16788,N_13469,N_14963);
xor U16789 (N_16789,N_14182,N_15079);
and U16790 (N_16790,N_13250,N_14224);
nor U16791 (N_16791,N_12639,N_13493);
and U16792 (N_16792,N_15598,N_13135);
xnor U16793 (N_16793,N_13799,N_15471);
nor U16794 (N_16794,N_13260,N_15416);
and U16795 (N_16795,N_14486,N_14944);
nor U16796 (N_16796,N_14593,N_13598);
nand U16797 (N_16797,N_13091,N_12675);
xor U16798 (N_16798,N_14733,N_14075);
xor U16799 (N_16799,N_15603,N_13254);
and U16800 (N_16800,N_14575,N_13919);
nand U16801 (N_16801,N_13541,N_14530);
xor U16802 (N_16802,N_12848,N_15275);
nor U16803 (N_16803,N_14912,N_15528);
nand U16804 (N_16804,N_13766,N_13844);
nand U16805 (N_16805,N_13829,N_14464);
nand U16806 (N_16806,N_13704,N_13898);
and U16807 (N_16807,N_13478,N_12552);
or U16808 (N_16808,N_14662,N_12977);
and U16809 (N_16809,N_12932,N_14544);
or U16810 (N_16810,N_15286,N_15590);
nor U16811 (N_16811,N_14071,N_14196);
nor U16812 (N_16812,N_15460,N_15056);
and U16813 (N_16813,N_13858,N_12990);
nand U16814 (N_16814,N_15215,N_15112);
nor U16815 (N_16815,N_14836,N_15226);
nand U16816 (N_16816,N_14399,N_13549);
nor U16817 (N_16817,N_13981,N_14550);
nand U16818 (N_16818,N_14432,N_13787);
nand U16819 (N_16819,N_12966,N_12689);
nand U16820 (N_16820,N_15026,N_14390);
nand U16821 (N_16821,N_14799,N_15349);
and U16822 (N_16822,N_14683,N_13539);
nor U16823 (N_16823,N_14816,N_13365);
and U16824 (N_16824,N_14854,N_12794);
or U16825 (N_16825,N_12589,N_13346);
or U16826 (N_16826,N_15024,N_12894);
nand U16827 (N_16827,N_13942,N_14793);
and U16828 (N_16828,N_14156,N_15311);
or U16829 (N_16829,N_13627,N_13572);
nand U16830 (N_16830,N_13626,N_14335);
nand U16831 (N_16831,N_14243,N_14723);
or U16832 (N_16832,N_14639,N_13540);
xor U16833 (N_16833,N_13317,N_14011);
and U16834 (N_16834,N_15058,N_13002);
and U16835 (N_16835,N_15541,N_12844);
nor U16836 (N_16836,N_13163,N_14725);
and U16837 (N_16837,N_14336,N_13717);
nand U16838 (N_16838,N_13171,N_13168);
nand U16839 (N_16839,N_15277,N_12979);
or U16840 (N_16840,N_15178,N_12808);
nor U16841 (N_16841,N_14358,N_13589);
or U16842 (N_16842,N_13064,N_12607);
or U16843 (N_16843,N_14305,N_14419);
nand U16844 (N_16844,N_13147,N_13798);
xnor U16845 (N_16845,N_14381,N_13998);
nand U16846 (N_16846,N_12580,N_15336);
nor U16847 (N_16847,N_15134,N_14956);
nor U16848 (N_16848,N_15291,N_15255);
and U16849 (N_16849,N_15148,N_13445);
and U16850 (N_16850,N_14008,N_14528);
or U16851 (N_16851,N_14476,N_13019);
and U16852 (N_16852,N_14259,N_14839);
nor U16853 (N_16853,N_14452,N_14501);
nand U16854 (N_16854,N_13065,N_15294);
or U16855 (N_16855,N_13700,N_15446);
nand U16856 (N_16856,N_13327,N_13530);
or U16857 (N_16857,N_14412,N_14289);
xnor U16858 (N_16858,N_15245,N_14920);
nand U16859 (N_16859,N_13180,N_14006);
xor U16860 (N_16860,N_13083,N_15544);
xor U16861 (N_16861,N_14921,N_13211);
nand U16862 (N_16862,N_15208,N_14251);
nand U16863 (N_16863,N_14157,N_13831);
xnor U16864 (N_16864,N_15453,N_14619);
nor U16865 (N_16865,N_15450,N_15224);
nand U16866 (N_16866,N_12747,N_13213);
or U16867 (N_16867,N_13097,N_13246);
or U16868 (N_16868,N_12618,N_15487);
and U16869 (N_16869,N_13856,N_12923);
and U16870 (N_16870,N_14113,N_15040);
xor U16871 (N_16871,N_15519,N_15526);
and U16872 (N_16872,N_15191,N_13255);
or U16873 (N_16873,N_14290,N_14872);
or U16874 (N_16874,N_13788,N_13151);
nor U16875 (N_16875,N_14796,N_14284);
or U16876 (N_16876,N_15579,N_12751);
nand U16877 (N_16877,N_13170,N_12672);
nor U16878 (N_16878,N_13350,N_13334);
or U16879 (N_16879,N_13722,N_13896);
and U16880 (N_16880,N_12620,N_14441);
nand U16881 (N_16881,N_15116,N_15076);
nor U16882 (N_16882,N_12988,N_15573);
nand U16883 (N_16883,N_15212,N_14776);
and U16884 (N_16884,N_14488,N_12572);
xor U16885 (N_16885,N_13464,N_14063);
and U16886 (N_16886,N_15428,N_14565);
nand U16887 (N_16887,N_15505,N_13459);
nor U16888 (N_16888,N_13026,N_13139);
xnor U16889 (N_16889,N_14309,N_12650);
nor U16890 (N_16890,N_13495,N_14025);
nand U16891 (N_16891,N_13887,N_13394);
or U16892 (N_16892,N_13875,N_12759);
or U16893 (N_16893,N_13669,N_12584);
and U16894 (N_16894,N_13544,N_13671);
and U16895 (N_16895,N_14576,N_13053);
or U16896 (N_16896,N_14248,N_15329);
nor U16897 (N_16897,N_13319,N_12683);
or U16898 (N_16898,N_13550,N_14126);
or U16899 (N_16899,N_14485,N_14660);
nor U16900 (N_16900,N_13538,N_15454);
or U16901 (N_16901,N_14775,N_13622);
nand U16902 (N_16902,N_14454,N_14092);
and U16903 (N_16903,N_15103,N_14623);
and U16904 (N_16904,N_14173,N_13537);
nor U16905 (N_16905,N_14190,N_13315);
nand U16906 (N_16906,N_14579,N_13621);
and U16907 (N_16907,N_14620,N_13515);
nor U16908 (N_16908,N_12803,N_15386);
xor U16909 (N_16909,N_14098,N_14367);
and U16910 (N_16910,N_13073,N_13182);
or U16911 (N_16911,N_14624,N_13955);
or U16912 (N_16912,N_13933,N_13032);
nand U16913 (N_16913,N_15506,N_12533);
nor U16914 (N_16914,N_14342,N_12570);
and U16915 (N_16915,N_15406,N_14686);
nand U16916 (N_16916,N_14120,N_15564);
or U16917 (N_16917,N_13630,N_13526);
xnor U16918 (N_16918,N_13996,N_13653);
or U16919 (N_16919,N_13203,N_15113);
or U16920 (N_16920,N_14566,N_15550);
nand U16921 (N_16921,N_13738,N_15498);
and U16922 (N_16922,N_14652,N_13690);
and U16923 (N_16923,N_14389,N_12857);
and U16924 (N_16924,N_14940,N_13496);
xnor U16925 (N_16925,N_14046,N_13963);
nor U16926 (N_16926,N_13956,N_13314);
and U16927 (N_16927,N_15398,N_14204);
nor U16928 (N_16928,N_12785,N_13886);
nand U16929 (N_16929,N_13643,N_12887);
and U16930 (N_16930,N_14690,N_13218);
nand U16931 (N_16931,N_12537,N_14508);
nand U16932 (N_16932,N_15150,N_14446);
nor U16933 (N_16933,N_14143,N_14318);
nand U16934 (N_16934,N_13591,N_12542);
and U16935 (N_16935,N_14640,N_15293);
and U16936 (N_16936,N_13024,N_13884);
nand U16937 (N_16937,N_14127,N_13185);
or U16938 (N_16938,N_13364,N_14437);
nand U16939 (N_16939,N_14866,N_15082);
nand U16940 (N_16940,N_14262,N_13824);
nor U16941 (N_16941,N_14024,N_13576);
or U16942 (N_16942,N_12601,N_15468);
and U16943 (N_16943,N_13881,N_13096);
and U16944 (N_16944,N_14737,N_15585);
and U16945 (N_16945,N_15447,N_12568);
nor U16946 (N_16946,N_13467,N_13229);
nor U16947 (N_16947,N_13116,N_14851);
nand U16948 (N_16948,N_13730,N_13605);
nor U16949 (N_16949,N_12819,N_12524);
and U16950 (N_16950,N_13008,N_12736);
or U16951 (N_16951,N_13075,N_14983);
nor U16952 (N_16952,N_13548,N_13705);
and U16953 (N_16953,N_14742,N_14430);
nand U16954 (N_16954,N_15381,N_13407);
nand U16955 (N_16955,N_14822,N_12846);
and U16956 (N_16956,N_15467,N_15373);
or U16957 (N_16957,N_13152,N_15319);
and U16958 (N_16958,N_13440,N_14352);
nand U16959 (N_16959,N_15361,N_13192);
nor U16960 (N_16960,N_13068,N_14064);
or U16961 (N_16961,N_12947,N_13164);
nand U16962 (N_16962,N_12590,N_13066);
and U16963 (N_16963,N_15502,N_13326);
nand U16964 (N_16964,N_12681,N_15570);
nand U16965 (N_16965,N_14780,N_14629);
xor U16966 (N_16966,N_15197,N_13466);
or U16967 (N_16967,N_15126,N_13404);
nor U16968 (N_16968,N_14841,N_14176);
and U16969 (N_16969,N_15051,N_13366);
nor U16970 (N_16970,N_12507,N_15117);
nand U16971 (N_16971,N_15425,N_14961);
nand U16972 (N_16972,N_14140,N_14254);
nor U16973 (N_16973,N_14967,N_15389);
nand U16974 (N_16974,N_14700,N_14035);
and U16975 (N_16975,N_14684,N_15333);
and U16976 (N_16976,N_12995,N_14198);
and U16977 (N_16977,N_13827,N_15142);
nand U16978 (N_16978,N_13453,N_12662);
nand U16979 (N_16979,N_13228,N_13718);
nand U16980 (N_16980,N_13140,N_15069);
and U16981 (N_16981,N_14457,N_12789);
and U16982 (N_16982,N_12640,N_13110);
nand U16983 (N_16983,N_15463,N_13020);
nor U16984 (N_16984,N_15071,N_15143);
and U16985 (N_16985,N_12515,N_14138);
nor U16986 (N_16986,N_15061,N_14555);
nand U16987 (N_16987,N_14928,N_14853);
nand U16988 (N_16988,N_14916,N_14886);
nand U16989 (N_16989,N_15578,N_15582);
and U16990 (N_16990,N_14180,N_15170);
nand U16991 (N_16991,N_12926,N_15596);
xor U16992 (N_16992,N_12869,N_14759);
xor U16993 (N_16993,N_15475,N_15534);
nand U16994 (N_16994,N_12603,N_14323);
nand U16995 (N_16995,N_15337,N_13384);
nand U16996 (N_16996,N_13721,N_15187);
and U16997 (N_16997,N_13678,N_13276);
and U16998 (N_16998,N_14362,N_12996);
nor U16999 (N_16999,N_13754,N_14321);
and U17000 (N_17000,N_14525,N_13562);
nor U17001 (N_17001,N_12597,N_14568);
or U17002 (N_17002,N_13681,N_13413);
or U17003 (N_17003,N_15022,N_14504);
nand U17004 (N_17004,N_12521,N_12920);
xor U17005 (N_17005,N_13098,N_13479);
nor U17006 (N_17006,N_13344,N_14602);
nand U17007 (N_17007,N_13732,N_15188);
and U17008 (N_17008,N_13835,N_15469);
and U17009 (N_17009,N_13800,N_15483);
and U17010 (N_17010,N_13563,N_13865);
and U17011 (N_17011,N_14082,N_14599);
or U17012 (N_17012,N_15314,N_13157);
nand U17013 (N_17013,N_13852,N_15225);
nor U17014 (N_17014,N_14803,N_15285);
nor U17015 (N_17015,N_14817,N_14329);
nor U17016 (N_17016,N_15207,N_14585);
and U17017 (N_17017,N_14031,N_14726);
and U17018 (N_17018,N_13891,N_13635);
nand U17019 (N_17019,N_14283,N_14739);
or U17020 (N_17020,N_13374,N_13894);
or U17021 (N_17021,N_15486,N_14502);
and U17022 (N_17022,N_15393,N_13463);
or U17023 (N_17023,N_12775,N_12906);
or U17024 (N_17024,N_12624,N_15589);
and U17025 (N_17025,N_15499,N_13641);
xnor U17026 (N_17026,N_13736,N_12858);
xor U17027 (N_17027,N_12746,N_14118);
nor U17028 (N_17028,N_14405,N_13049);
nor U17029 (N_17029,N_14618,N_15192);
nor U17030 (N_17030,N_14388,N_14753);
nor U17031 (N_17031,N_15184,N_15096);
nand U17032 (N_17032,N_14675,N_13864);
nor U17033 (N_17033,N_12982,N_12939);
nand U17034 (N_17034,N_12811,N_13268);
and U17035 (N_17035,N_15362,N_13793);
nand U17036 (N_17036,N_14506,N_15078);
or U17037 (N_17037,N_15371,N_15055);
xnor U17038 (N_17038,N_14191,N_15435);
nor U17039 (N_17039,N_14521,N_12529);
nor U17040 (N_17040,N_12941,N_12950);
or U17041 (N_17041,N_12598,N_15350);
nor U17042 (N_17042,N_12503,N_14439);
and U17043 (N_17043,N_12510,N_15448);
nand U17044 (N_17044,N_12805,N_14969);
xnor U17045 (N_17045,N_13654,N_15513);
nand U17046 (N_17046,N_14548,N_14371);
nand U17047 (N_17047,N_15041,N_13093);
nor U17048 (N_17048,N_15186,N_15546);
nand U17049 (N_17049,N_15259,N_13289);
xnor U17050 (N_17050,N_15249,N_12784);
or U17051 (N_17051,N_13561,N_12773);
nor U17052 (N_17052,N_14233,N_14876);
and U17053 (N_17053,N_12944,N_13594);
nand U17054 (N_17054,N_12760,N_15609);
and U17055 (N_17055,N_14056,N_13219);
xor U17056 (N_17056,N_15295,N_15242);
nor U17057 (N_17057,N_13133,N_14034);
and U17058 (N_17058,N_14808,N_14420);
nand U17059 (N_17059,N_15006,N_12718);
and U17060 (N_17060,N_14402,N_14765);
and U17061 (N_17061,N_13527,N_13353);
nor U17062 (N_17062,N_13357,N_14115);
nor U17063 (N_17063,N_15095,N_12892);
and U17064 (N_17064,N_13409,N_14667);
nor U17065 (N_17065,N_14516,N_14493);
nor U17066 (N_17066,N_12884,N_12716);
or U17067 (N_17067,N_15107,N_13712);
or U17068 (N_17068,N_15093,N_12545);
nand U17069 (N_17069,N_15155,N_14164);
and U17070 (N_17070,N_13553,N_15340);
and U17071 (N_17071,N_15424,N_14877);
and U17072 (N_17072,N_13119,N_14014);
and U17073 (N_17073,N_14054,N_12860);
nor U17074 (N_17074,N_15059,N_13506);
nand U17075 (N_17075,N_12800,N_14267);
and U17076 (N_17076,N_14292,N_13975);
nand U17077 (N_17077,N_12876,N_13860);
or U17078 (N_17078,N_14216,N_14895);
or U17079 (N_17079,N_12960,N_14721);
or U17080 (N_17080,N_14616,N_13088);
nor U17081 (N_17081,N_13578,N_14212);
xor U17082 (N_17082,N_14002,N_13485);
or U17083 (N_17083,N_14583,N_12936);
nand U17084 (N_17084,N_13834,N_12613);
xor U17085 (N_17085,N_14750,N_13595);
nand U17086 (N_17086,N_14465,N_14589);
nor U17087 (N_17087,N_12955,N_13726);
and U17088 (N_17088,N_13997,N_14350);
or U17089 (N_17089,N_13784,N_13076);
or U17090 (N_17090,N_12904,N_13310);
xor U17091 (N_17091,N_14727,N_13650);
nor U17092 (N_17092,N_13952,N_14058);
nor U17093 (N_17093,N_13588,N_14108);
or U17094 (N_17094,N_15297,N_14087);
and U17095 (N_17095,N_14826,N_12832);
nor U17096 (N_17096,N_12919,N_13178);
and U17097 (N_17097,N_15378,N_13431);
or U17098 (N_17098,N_13559,N_12727);
or U17099 (N_17099,N_14298,N_13675);
and U17100 (N_17100,N_13755,N_15165);
or U17101 (N_17101,N_13940,N_14734);
xnor U17102 (N_17102,N_12834,N_14532);
nand U17103 (N_17103,N_14206,N_13714);
and U17104 (N_17104,N_13775,N_15348);
and U17105 (N_17105,N_14240,N_14492);
and U17106 (N_17106,N_14380,N_13351);
or U17107 (N_17107,N_14376,N_14703);
and U17108 (N_17108,N_14968,N_14498);
xnor U17109 (N_17109,N_13869,N_14356);
nand U17110 (N_17110,N_15553,N_14883);
nor U17111 (N_17111,N_12626,N_15141);
nor U17112 (N_17112,N_14238,N_12830);
nor U17113 (N_17113,N_14627,N_15160);
nor U17114 (N_17114,N_14774,N_12605);
xor U17115 (N_17115,N_12508,N_15274);
nor U17116 (N_17116,N_14436,N_12967);
and U17117 (N_17117,N_12642,N_14704);
and U17118 (N_17118,N_13082,N_13729);
and U17119 (N_17119,N_12821,N_12600);
xor U17120 (N_17120,N_15538,N_13664);
and U17121 (N_17121,N_12658,N_13126);
xor U17122 (N_17122,N_14603,N_14634);
or U17123 (N_17123,N_13618,N_12551);
xor U17124 (N_17124,N_15009,N_13142);
nand U17125 (N_17125,N_13833,N_14160);
and U17126 (N_17126,N_15153,N_13524);
nand U17127 (N_17127,N_13582,N_12963);
xor U17128 (N_17128,N_13657,N_14018);
nor U17129 (N_17129,N_13039,N_13851);
or U17130 (N_17130,N_13600,N_12837);
and U17131 (N_17131,N_15380,N_12863);
and U17132 (N_17132,N_15500,N_14990);
or U17133 (N_17133,N_14047,N_12792);
nand U17134 (N_17134,N_15527,N_12975);
nand U17135 (N_17135,N_12530,N_14174);
and U17136 (N_17136,N_12724,N_12708);
or U17137 (N_17137,N_13474,N_14709);
or U17138 (N_17138,N_13252,N_15029);
or U17139 (N_17139,N_13369,N_14924);
and U17140 (N_17140,N_13361,N_12656);
nand U17141 (N_17141,N_15452,N_14407);
or U17142 (N_17142,N_12962,N_15077);
nor U17143 (N_17143,N_14203,N_15292);
and U17144 (N_17144,N_14591,N_15257);
xnor U17145 (N_17145,N_14076,N_13029);
and U17146 (N_17146,N_12968,N_13660);
xnor U17147 (N_17147,N_14862,N_13733);
or U17148 (N_17148,N_13802,N_14717);
and U17149 (N_17149,N_15158,N_12698);
and U17150 (N_17150,N_15614,N_14788);
nand U17151 (N_17151,N_15367,N_14559);
or U17152 (N_17152,N_15086,N_14106);
nand U17153 (N_17153,N_15136,N_12706);
or U17154 (N_17154,N_13401,N_13298);
and U17155 (N_17155,N_12997,N_12964);
and U17156 (N_17156,N_15434,N_14219);
nor U17157 (N_17157,N_14661,N_13106);
nor U17158 (N_17158,N_13629,N_14878);
nand U17159 (N_17159,N_12949,N_15074);
xnor U17160 (N_17160,N_14266,N_14458);
and U17161 (N_17161,N_14077,N_14612);
and U17162 (N_17162,N_13742,N_13295);
nand U17163 (N_17163,N_14060,N_13396);
or U17164 (N_17164,N_15067,N_15493);
and U17165 (N_17165,N_12645,N_13427);
nand U17166 (N_17166,N_14760,N_12942);
or U17167 (N_17167,N_14043,N_14370);
xnor U17168 (N_17168,N_14451,N_15219);
nand U17169 (N_17169,N_14891,N_13529);
or U17170 (N_17170,N_13767,N_15481);
nor U17171 (N_17171,N_14351,N_13475);
xnor U17172 (N_17172,N_14051,N_13313);
or U17173 (N_17173,N_14215,N_15261);
nor U17174 (N_17174,N_13060,N_15102);
and U17175 (N_17175,N_12970,N_13311);
nor U17176 (N_17176,N_14798,N_14840);
nand U17177 (N_17177,N_12835,N_13251);
xnor U17178 (N_17178,N_13628,N_14740);
nor U17179 (N_17179,N_13308,N_12616);
nor U17180 (N_17180,N_15110,N_14012);
and U17181 (N_17181,N_14015,N_12823);
or U17182 (N_17182,N_15419,N_13922);
nand U17183 (N_17183,N_15616,N_14032);
xor U17184 (N_17184,N_12665,N_14237);
nor U17185 (N_17185,N_13794,N_13484);
nand U17186 (N_17186,N_13472,N_14754);
or U17187 (N_17187,N_14081,N_14792);
nand U17188 (N_17188,N_14126,N_14329);
or U17189 (N_17189,N_15440,N_13454);
and U17190 (N_17190,N_13137,N_15114);
and U17191 (N_17191,N_13071,N_13395);
or U17192 (N_17192,N_13543,N_13382);
nor U17193 (N_17193,N_14559,N_15449);
and U17194 (N_17194,N_15439,N_14457);
and U17195 (N_17195,N_14752,N_13010);
nand U17196 (N_17196,N_13133,N_13165);
nor U17197 (N_17197,N_14673,N_13127);
or U17198 (N_17198,N_14953,N_14955);
nand U17199 (N_17199,N_15181,N_14151);
nand U17200 (N_17200,N_14535,N_15226);
nor U17201 (N_17201,N_14351,N_12771);
and U17202 (N_17202,N_12793,N_13961);
nor U17203 (N_17203,N_14441,N_14868);
nor U17204 (N_17204,N_13340,N_14574);
nand U17205 (N_17205,N_12643,N_15493);
nor U17206 (N_17206,N_15271,N_13443);
nor U17207 (N_17207,N_14225,N_13182);
nor U17208 (N_17208,N_15140,N_13203);
nor U17209 (N_17209,N_13208,N_15212);
or U17210 (N_17210,N_13485,N_14011);
and U17211 (N_17211,N_12641,N_13767);
nand U17212 (N_17212,N_12526,N_13760);
nand U17213 (N_17213,N_14698,N_12681);
or U17214 (N_17214,N_14912,N_13921);
nand U17215 (N_17215,N_14052,N_15532);
and U17216 (N_17216,N_14113,N_15502);
nor U17217 (N_17217,N_13391,N_14913);
nand U17218 (N_17218,N_15085,N_14257);
or U17219 (N_17219,N_12967,N_14517);
nor U17220 (N_17220,N_13652,N_12809);
nor U17221 (N_17221,N_14126,N_13659);
xor U17222 (N_17222,N_14525,N_13283);
nor U17223 (N_17223,N_13468,N_15203);
and U17224 (N_17224,N_12851,N_13741);
nand U17225 (N_17225,N_15125,N_12700);
xor U17226 (N_17226,N_13733,N_12883);
nor U17227 (N_17227,N_13956,N_14569);
or U17228 (N_17228,N_13402,N_12851);
and U17229 (N_17229,N_14877,N_14785);
nand U17230 (N_17230,N_15447,N_14269);
xor U17231 (N_17231,N_12941,N_13132);
nor U17232 (N_17232,N_14200,N_12578);
and U17233 (N_17233,N_14757,N_15075);
nand U17234 (N_17234,N_14585,N_15265);
or U17235 (N_17235,N_14510,N_14426);
or U17236 (N_17236,N_14079,N_15302);
and U17237 (N_17237,N_12815,N_13002);
nor U17238 (N_17238,N_13334,N_13319);
or U17239 (N_17239,N_13039,N_14598);
nor U17240 (N_17240,N_14323,N_14967);
nor U17241 (N_17241,N_15157,N_14863);
or U17242 (N_17242,N_13204,N_13450);
nor U17243 (N_17243,N_14327,N_14184);
or U17244 (N_17244,N_13661,N_14969);
xnor U17245 (N_17245,N_14757,N_12863);
nor U17246 (N_17246,N_15045,N_12908);
nand U17247 (N_17247,N_12525,N_13203);
nor U17248 (N_17248,N_15611,N_13429);
or U17249 (N_17249,N_14308,N_13357);
and U17250 (N_17250,N_14371,N_15265);
nor U17251 (N_17251,N_15488,N_13274);
xnor U17252 (N_17252,N_12895,N_14958);
xnor U17253 (N_17253,N_13376,N_13610);
and U17254 (N_17254,N_14249,N_13337);
nor U17255 (N_17255,N_13620,N_12739);
and U17256 (N_17256,N_12751,N_13099);
xnor U17257 (N_17257,N_13277,N_12558);
nor U17258 (N_17258,N_12722,N_14345);
nand U17259 (N_17259,N_13489,N_15556);
or U17260 (N_17260,N_13253,N_14695);
or U17261 (N_17261,N_14705,N_14864);
xor U17262 (N_17262,N_12836,N_15049);
nor U17263 (N_17263,N_15182,N_15194);
nand U17264 (N_17264,N_14256,N_12793);
nor U17265 (N_17265,N_13587,N_12859);
nand U17266 (N_17266,N_15572,N_12657);
or U17267 (N_17267,N_14099,N_15143);
nor U17268 (N_17268,N_15243,N_13657);
nand U17269 (N_17269,N_13030,N_14647);
nor U17270 (N_17270,N_13973,N_13496);
or U17271 (N_17271,N_12755,N_13090);
nor U17272 (N_17272,N_12573,N_12652);
nand U17273 (N_17273,N_12785,N_13411);
and U17274 (N_17274,N_14900,N_14365);
nor U17275 (N_17275,N_14384,N_13607);
nand U17276 (N_17276,N_15167,N_12975);
xnor U17277 (N_17277,N_14487,N_15435);
and U17278 (N_17278,N_14169,N_13834);
and U17279 (N_17279,N_13195,N_15361);
and U17280 (N_17280,N_14773,N_14514);
nor U17281 (N_17281,N_13146,N_15316);
or U17282 (N_17282,N_15069,N_13766);
xor U17283 (N_17283,N_12755,N_12502);
or U17284 (N_17284,N_12919,N_15014);
xnor U17285 (N_17285,N_15389,N_13797);
nand U17286 (N_17286,N_14123,N_13286);
or U17287 (N_17287,N_14545,N_14486);
nor U17288 (N_17288,N_13736,N_15012);
nand U17289 (N_17289,N_12608,N_13672);
or U17290 (N_17290,N_15587,N_13973);
nor U17291 (N_17291,N_13513,N_13540);
xor U17292 (N_17292,N_15311,N_13518);
xnor U17293 (N_17293,N_12815,N_12998);
xnor U17294 (N_17294,N_13759,N_12851);
xnor U17295 (N_17295,N_13365,N_13051);
or U17296 (N_17296,N_13109,N_14800);
or U17297 (N_17297,N_13450,N_12938);
nor U17298 (N_17298,N_15235,N_12857);
and U17299 (N_17299,N_12616,N_14357);
or U17300 (N_17300,N_14539,N_13946);
nand U17301 (N_17301,N_13714,N_14025);
nand U17302 (N_17302,N_12978,N_14089);
or U17303 (N_17303,N_14477,N_15420);
nor U17304 (N_17304,N_13607,N_12771);
nor U17305 (N_17305,N_14957,N_14073);
nor U17306 (N_17306,N_14823,N_14789);
nand U17307 (N_17307,N_13860,N_14067);
xnor U17308 (N_17308,N_13051,N_14701);
and U17309 (N_17309,N_14216,N_12630);
xor U17310 (N_17310,N_14301,N_12726);
and U17311 (N_17311,N_13880,N_14931);
nor U17312 (N_17312,N_13020,N_15524);
and U17313 (N_17313,N_13202,N_12656);
xnor U17314 (N_17314,N_15525,N_12999);
or U17315 (N_17315,N_12623,N_13290);
nand U17316 (N_17316,N_12836,N_13324);
and U17317 (N_17317,N_13947,N_14733);
nor U17318 (N_17318,N_15353,N_14095);
or U17319 (N_17319,N_15621,N_14467);
nand U17320 (N_17320,N_14363,N_14408);
and U17321 (N_17321,N_14226,N_15067);
nor U17322 (N_17322,N_14421,N_14983);
nand U17323 (N_17323,N_13965,N_15465);
nor U17324 (N_17324,N_13409,N_12953);
and U17325 (N_17325,N_14000,N_12774);
and U17326 (N_17326,N_15305,N_15334);
and U17327 (N_17327,N_15620,N_14654);
nand U17328 (N_17328,N_15307,N_13576);
or U17329 (N_17329,N_13515,N_14544);
nand U17330 (N_17330,N_12503,N_14827);
nand U17331 (N_17331,N_15056,N_14216);
nor U17332 (N_17332,N_13429,N_12814);
and U17333 (N_17333,N_14368,N_13487);
nand U17334 (N_17334,N_14530,N_13830);
or U17335 (N_17335,N_12779,N_14469);
nand U17336 (N_17336,N_14889,N_13724);
nand U17337 (N_17337,N_14032,N_13201);
or U17338 (N_17338,N_14022,N_14044);
nand U17339 (N_17339,N_14845,N_13784);
nor U17340 (N_17340,N_13543,N_15188);
and U17341 (N_17341,N_15607,N_12576);
xnor U17342 (N_17342,N_13257,N_12748);
or U17343 (N_17343,N_14920,N_14667);
nor U17344 (N_17344,N_15340,N_14993);
xnor U17345 (N_17345,N_13217,N_14400);
xor U17346 (N_17346,N_14913,N_12738);
or U17347 (N_17347,N_15602,N_14230);
or U17348 (N_17348,N_14693,N_15018);
nor U17349 (N_17349,N_14333,N_15429);
xnor U17350 (N_17350,N_14643,N_12602);
nand U17351 (N_17351,N_14018,N_14508);
nor U17352 (N_17352,N_15388,N_12611);
nand U17353 (N_17353,N_12511,N_14384);
or U17354 (N_17354,N_14507,N_13451);
nand U17355 (N_17355,N_14745,N_12815);
nand U17356 (N_17356,N_14950,N_14012);
or U17357 (N_17357,N_14945,N_13715);
nor U17358 (N_17358,N_12538,N_15606);
and U17359 (N_17359,N_15536,N_14387);
nor U17360 (N_17360,N_14679,N_13284);
and U17361 (N_17361,N_14940,N_14225);
or U17362 (N_17362,N_13542,N_15133);
or U17363 (N_17363,N_14506,N_14436);
and U17364 (N_17364,N_14103,N_14374);
xnor U17365 (N_17365,N_14307,N_14872);
and U17366 (N_17366,N_13578,N_15456);
or U17367 (N_17367,N_13874,N_14126);
nor U17368 (N_17368,N_14948,N_15613);
and U17369 (N_17369,N_13226,N_14456);
and U17370 (N_17370,N_15118,N_14347);
nor U17371 (N_17371,N_15589,N_13465);
nand U17372 (N_17372,N_13244,N_14815);
xor U17373 (N_17373,N_14227,N_15010);
and U17374 (N_17374,N_13727,N_14487);
xor U17375 (N_17375,N_13418,N_13485);
nor U17376 (N_17376,N_13226,N_12608);
nor U17377 (N_17377,N_14094,N_13849);
xor U17378 (N_17378,N_14871,N_12836);
nor U17379 (N_17379,N_13709,N_14836);
nand U17380 (N_17380,N_14591,N_12548);
and U17381 (N_17381,N_13787,N_15613);
nor U17382 (N_17382,N_14440,N_13393);
xnor U17383 (N_17383,N_15487,N_13043);
nand U17384 (N_17384,N_14390,N_12645);
nor U17385 (N_17385,N_12799,N_12703);
nand U17386 (N_17386,N_14976,N_14880);
nor U17387 (N_17387,N_12708,N_14115);
or U17388 (N_17388,N_15283,N_14669);
and U17389 (N_17389,N_13591,N_14434);
xnor U17390 (N_17390,N_14693,N_12902);
or U17391 (N_17391,N_14536,N_14715);
nor U17392 (N_17392,N_13414,N_13087);
nand U17393 (N_17393,N_13622,N_12601);
or U17394 (N_17394,N_12567,N_13275);
or U17395 (N_17395,N_15224,N_14783);
nand U17396 (N_17396,N_12735,N_14412);
and U17397 (N_17397,N_14334,N_14622);
and U17398 (N_17398,N_13036,N_13553);
or U17399 (N_17399,N_13413,N_15391);
or U17400 (N_17400,N_12660,N_13552);
nor U17401 (N_17401,N_13415,N_14210);
or U17402 (N_17402,N_13702,N_13823);
or U17403 (N_17403,N_13862,N_15107);
nor U17404 (N_17404,N_14100,N_14378);
or U17405 (N_17405,N_13012,N_15428);
nand U17406 (N_17406,N_14186,N_15247);
nor U17407 (N_17407,N_13765,N_12984);
and U17408 (N_17408,N_15053,N_13909);
and U17409 (N_17409,N_14987,N_14373);
or U17410 (N_17410,N_15326,N_12652);
nor U17411 (N_17411,N_13354,N_15595);
or U17412 (N_17412,N_15466,N_15105);
nor U17413 (N_17413,N_12628,N_15561);
and U17414 (N_17414,N_14456,N_12680);
or U17415 (N_17415,N_15387,N_13713);
and U17416 (N_17416,N_13107,N_13075);
nor U17417 (N_17417,N_15406,N_12560);
nor U17418 (N_17418,N_15097,N_13191);
and U17419 (N_17419,N_15549,N_13836);
and U17420 (N_17420,N_12786,N_14371);
nor U17421 (N_17421,N_15543,N_15343);
nand U17422 (N_17422,N_15539,N_13057);
and U17423 (N_17423,N_12807,N_14559);
nand U17424 (N_17424,N_13057,N_12511);
or U17425 (N_17425,N_15093,N_14924);
or U17426 (N_17426,N_14198,N_15049);
nand U17427 (N_17427,N_13691,N_14497);
nor U17428 (N_17428,N_12563,N_13515);
and U17429 (N_17429,N_15226,N_14319);
nor U17430 (N_17430,N_13133,N_14617);
nor U17431 (N_17431,N_14136,N_13595);
nand U17432 (N_17432,N_13239,N_14172);
xnor U17433 (N_17433,N_13412,N_15022);
nand U17434 (N_17434,N_12978,N_14130);
and U17435 (N_17435,N_12941,N_15184);
and U17436 (N_17436,N_15527,N_13649);
or U17437 (N_17437,N_12901,N_13383);
and U17438 (N_17438,N_15581,N_13525);
nand U17439 (N_17439,N_12540,N_14308);
and U17440 (N_17440,N_12582,N_15570);
nor U17441 (N_17441,N_15263,N_15042);
nand U17442 (N_17442,N_14134,N_13590);
xor U17443 (N_17443,N_14296,N_13686);
nand U17444 (N_17444,N_13191,N_13891);
xor U17445 (N_17445,N_13351,N_14374);
and U17446 (N_17446,N_13206,N_13056);
nor U17447 (N_17447,N_14681,N_14359);
or U17448 (N_17448,N_12812,N_15120);
and U17449 (N_17449,N_12824,N_14991);
nand U17450 (N_17450,N_12576,N_14568);
nor U17451 (N_17451,N_12556,N_14935);
or U17452 (N_17452,N_13552,N_14969);
nand U17453 (N_17453,N_14706,N_14089);
or U17454 (N_17454,N_14759,N_15216);
nand U17455 (N_17455,N_13322,N_14271);
nand U17456 (N_17456,N_12728,N_14225);
and U17457 (N_17457,N_13475,N_12626);
nand U17458 (N_17458,N_14819,N_13534);
nand U17459 (N_17459,N_13831,N_14145);
nand U17460 (N_17460,N_14162,N_13524);
and U17461 (N_17461,N_14601,N_13353);
xnor U17462 (N_17462,N_13724,N_13734);
and U17463 (N_17463,N_14083,N_13002);
xor U17464 (N_17464,N_14173,N_15325);
nand U17465 (N_17465,N_13820,N_14895);
nor U17466 (N_17466,N_14794,N_14947);
and U17467 (N_17467,N_13820,N_13733);
nor U17468 (N_17468,N_13214,N_15320);
xnor U17469 (N_17469,N_15067,N_14134);
nor U17470 (N_17470,N_13846,N_14598);
nor U17471 (N_17471,N_15401,N_15087);
or U17472 (N_17472,N_14157,N_15346);
nor U17473 (N_17473,N_12537,N_13791);
or U17474 (N_17474,N_14596,N_14948);
or U17475 (N_17475,N_14914,N_15150);
nor U17476 (N_17476,N_15497,N_13331);
or U17477 (N_17477,N_15477,N_14372);
nor U17478 (N_17478,N_14022,N_14532);
nand U17479 (N_17479,N_13466,N_15539);
nand U17480 (N_17480,N_13071,N_13053);
and U17481 (N_17481,N_13967,N_13678);
or U17482 (N_17482,N_15233,N_13204);
nor U17483 (N_17483,N_13960,N_14546);
and U17484 (N_17484,N_15412,N_15512);
nand U17485 (N_17485,N_14182,N_14540);
nor U17486 (N_17486,N_13332,N_14738);
nand U17487 (N_17487,N_13990,N_15496);
nor U17488 (N_17488,N_15206,N_13920);
and U17489 (N_17489,N_13128,N_14300);
and U17490 (N_17490,N_14708,N_14039);
nor U17491 (N_17491,N_15164,N_14339);
nor U17492 (N_17492,N_14721,N_14420);
or U17493 (N_17493,N_14203,N_12815);
nand U17494 (N_17494,N_13272,N_14348);
nand U17495 (N_17495,N_14527,N_14332);
and U17496 (N_17496,N_15365,N_14928);
nor U17497 (N_17497,N_14208,N_15476);
nor U17498 (N_17498,N_13700,N_14801);
and U17499 (N_17499,N_13076,N_14271);
xor U17500 (N_17500,N_13755,N_15135);
or U17501 (N_17501,N_14636,N_12991);
nor U17502 (N_17502,N_13971,N_15249);
nor U17503 (N_17503,N_13546,N_13653);
nor U17504 (N_17504,N_13691,N_14618);
nand U17505 (N_17505,N_15085,N_15363);
nor U17506 (N_17506,N_12834,N_15028);
nand U17507 (N_17507,N_13893,N_15516);
and U17508 (N_17508,N_14693,N_13087);
or U17509 (N_17509,N_13366,N_15484);
and U17510 (N_17510,N_12954,N_13433);
or U17511 (N_17511,N_13161,N_12778);
nand U17512 (N_17512,N_14110,N_12657);
and U17513 (N_17513,N_13584,N_13676);
or U17514 (N_17514,N_15388,N_14850);
nand U17515 (N_17515,N_13424,N_15442);
nand U17516 (N_17516,N_12741,N_13267);
nor U17517 (N_17517,N_12905,N_12937);
and U17518 (N_17518,N_13146,N_12640);
xor U17519 (N_17519,N_14959,N_13661);
nor U17520 (N_17520,N_14064,N_14729);
nand U17521 (N_17521,N_14119,N_15329);
nand U17522 (N_17522,N_15306,N_13861);
xor U17523 (N_17523,N_14878,N_13650);
nor U17524 (N_17524,N_15517,N_12664);
xor U17525 (N_17525,N_13528,N_14726);
or U17526 (N_17526,N_15190,N_14352);
nor U17527 (N_17527,N_15283,N_13901);
or U17528 (N_17528,N_13002,N_12678);
nor U17529 (N_17529,N_15589,N_14886);
or U17530 (N_17530,N_14839,N_15138);
and U17531 (N_17531,N_13549,N_14767);
xnor U17532 (N_17532,N_14891,N_13324);
nand U17533 (N_17533,N_13464,N_12790);
nor U17534 (N_17534,N_15358,N_14152);
or U17535 (N_17535,N_15339,N_15525);
nor U17536 (N_17536,N_12847,N_12623);
xor U17537 (N_17537,N_15369,N_12845);
or U17538 (N_17538,N_14346,N_12525);
nand U17539 (N_17539,N_15552,N_13962);
or U17540 (N_17540,N_12737,N_13077);
nor U17541 (N_17541,N_14498,N_14899);
and U17542 (N_17542,N_12583,N_15546);
nand U17543 (N_17543,N_15249,N_15215);
nand U17544 (N_17544,N_13475,N_12795);
and U17545 (N_17545,N_14545,N_15428);
nor U17546 (N_17546,N_15291,N_14065);
xnor U17547 (N_17547,N_14918,N_13355);
and U17548 (N_17548,N_13360,N_15217);
or U17549 (N_17549,N_13701,N_13311);
xor U17550 (N_17550,N_14678,N_13961);
nand U17551 (N_17551,N_12722,N_14243);
nor U17552 (N_17552,N_14142,N_15114);
xor U17553 (N_17553,N_14414,N_15066);
nand U17554 (N_17554,N_15145,N_12738);
nor U17555 (N_17555,N_13974,N_13853);
or U17556 (N_17556,N_15324,N_14051);
and U17557 (N_17557,N_14976,N_13058);
and U17558 (N_17558,N_15553,N_15011);
nor U17559 (N_17559,N_14382,N_14908);
or U17560 (N_17560,N_12780,N_13911);
and U17561 (N_17561,N_12950,N_12972);
and U17562 (N_17562,N_14328,N_15045);
nand U17563 (N_17563,N_14930,N_13245);
or U17564 (N_17564,N_14257,N_13662);
nor U17565 (N_17565,N_14180,N_15482);
and U17566 (N_17566,N_12838,N_15388);
or U17567 (N_17567,N_13761,N_13668);
or U17568 (N_17568,N_13456,N_15388);
nor U17569 (N_17569,N_13549,N_14439);
or U17570 (N_17570,N_15442,N_15616);
or U17571 (N_17571,N_12909,N_14350);
and U17572 (N_17572,N_14138,N_12590);
or U17573 (N_17573,N_12801,N_14474);
nor U17574 (N_17574,N_12695,N_12558);
xor U17575 (N_17575,N_14893,N_14644);
and U17576 (N_17576,N_14311,N_13952);
or U17577 (N_17577,N_13975,N_13733);
nand U17578 (N_17578,N_15410,N_14853);
nand U17579 (N_17579,N_15327,N_15422);
or U17580 (N_17580,N_13789,N_14844);
or U17581 (N_17581,N_13242,N_15217);
nand U17582 (N_17582,N_13740,N_14594);
and U17583 (N_17583,N_12790,N_13688);
nor U17584 (N_17584,N_14061,N_12666);
nand U17585 (N_17585,N_15235,N_13496);
nor U17586 (N_17586,N_14584,N_13265);
and U17587 (N_17587,N_14066,N_15382);
or U17588 (N_17588,N_13953,N_14000);
and U17589 (N_17589,N_12737,N_12884);
nor U17590 (N_17590,N_14919,N_13024);
nand U17591 (N_17591,N_12693,N_13096);
nand U17592 (N_17592,N_13597,N_13639);
nor U17593 (N_17593,N_12716,N_15093);
nor U17594 (N_17594,N_13612,N_12898);
nand U17595 (N_17595,N_13256,N_13533);
or U17596 (N_17596,N_13224,N_13661);
nand U17597 (N_17597,N_14525,N_13019);
or U17598 (N_17598,N_13035,N_12939);
and U17599 (N_17599,N_15283,N_12793);
or U17600 (N_17600,N_15100,N_13310);
and U17601 (N_17601,N_13267,N_13288);
nand U17602 (N_17602,N_13931,N_14526);
nand U17603 (N_17603,N_13622,N_13528);
and U17604 (N_17604,N_14221,N_12638);
or U17605 (N_17605,N_13953,N_13840);
nor U17606 (N_17606,N_15210,N_12750);
or U17607 (N_17607,N_14713,N_14448);
nor U17608 (N_17608,N_14282,N_13871);
and U17609 (N_17609,N_14059,N_14136);
nor U17610 (N_17610,N_15220,N_14031);
nor U17611 (N_17611,N_14094,N_12990);
and U17612 (N_17612,N_13613,N_14089);
or U17613 (N_17613,N_13283,N_13521);
or U17614 (N_17614,N_12623,N_12737);
nor U17615 (N_17615,N_14768,N_13517);
nor U17616 (N_17616,N_15409,N_12595);
or U17617 (N_17617,N_12614,N_14460);
nor U17618 (N_17618,N_14827,N_14692);
or U17619 (N_17619,N_14666,N_13966);
xor U17620 (N_17620,N_14175,N_14478);
or U17621 (N_17621,N_14824,N_13945);
xnor U17622 (N_17622,N_15601,N_13898);
or U17623 (N_17623,N_14200,N_14512);
or U17624 (N_17624,N_13751,N_14006);
or U17625 (N_17625,N_13173,N_13635);
xnor U17626 (N_17626,N_13937,N_14013);
and U17627 (N_17627,N_13186,N_14205);
and U17628 (N_17628,N_13257,N_14949);
and U17629 (N_17629,N_13973,N_13676);
nor U17630 (N_17630,N_15019,N_13421);
and U17631 (N_17631,N_13818,N_14460);
and U17632 (N_17632,N_13080,N_15117);
or U17633 (N_17633,N_15246,N_14270);
nand U17634 (N_17634,N_13647,N_14261);
xnor U17635 (N_17635,N_12899,N_15431);
nand U17636 (N_17636,N_15362,N_15074);
nor U17637 (N_17637,N_13740,N_15372);
xor U17638 (N_17638,N_12814,N_12615);
or U17639 (N_17639,N_12768,N_15052);
xor U17640 (N_17640,N_14601,N_14306);
or U17641 (N_17641,N_12769,N_12682);
and U17642 (N_17642,N_14302,N_13659);
nand U17643 (N_17643,N_13389,N_15432);
nor U17644 (N_17644,N_14451,N_12570);
and U17645 (N_17645,N_14001,N_13237);
nand U17646 (N_17646,N_15070,N_12907);
or U17647 (N_17647,N_13216,N_14317);
nand U17648 (N_17648,N_12740,N_15526);
or U17649 (N_17649,N_14695,N_13812);
and U17650 (N_17650,N_14649,N_15336);
or U17651 (N_17651,N_14065,N_14007);
and U17652 (N_17652,N_13240,N_13302);
or U17653 (N_17653,N_12500,N_14851);
or U17654 (N_17654,N_13660,N_13668);
or U17655 (N_17655,N_14835,N_13544);
nand U17656 (N_17656,N_13806,N_14277);
and U17657 (N_17657,N_15595,N_12951);
nand U17658 (N_17658,N_13476,N_14199);
nand U17659 (N_17659,N_15476,N_14925);
xor U17660 (N_17660,N_13240,N_15565);
or U17661 (N_17661,N_14874,N_14296);
nor U17662 (N_17662,N_13465,N_15010);
or U17663 (N_17663,N_14980,N_14854);
or U17664 (N_17664,N_14563,N_13874);
nor U17665 (N_17665,N_14352,N_14200);
or U17666 (N_17666,N_14085,N_14718);
nor U17667 (N_17667,N_15338,N_14674);
nand U17668 (N_17668,N_14300,N_14625);
nor U17669 (N_17669,N_13921,N_15138);
nand U17670 (N_17670,N_13645,N_12705);
and U17671 (N_17671,N_12791,N_13082);
nand U17672 (N_17672,N_12991,N_12847);
xor U17673 (N_17673,N_12606,N_15522);
nand U17674 (N_17674,N_15527,N_12705);
or U17675 (N_17675,N_13087,N_14127);
or U17676 (N_17676,N_13274,N_15027);
nor U17677 (N_17677,N_14913,N_15228);
or U17678 (N_17678,N_15370,N_14140);
nor U17679 (N_17679,N_13266,N_12717);
and U17680 (N_17680,N_12928,N_14834);
or U17681 (N_17681,N_15311,N_13022);
nand U17682 (N_17682,N_12945,N_15276);
nor U17683 (N_17683,N_13083,N_13621);
nor U17684 (N_17684,N_12635,N_13113);
or U17685 (N_17685,N_15003,N_15153);
xnor U17686 (N_17686,N_13460,N_14686);
or U17687 (N_17687,N_14924,N_14986);
or U17688 (N_17688,N_12540,N_15542);
and U17689 (N_17689,N_14267,N_13222);
and U17690 (N_17690,N_14621,N_15120);
nand U17691 (N_17691,N_14569,N_15303);
nand U17692 (N_17692,N_15326,N_15029);
nor U17693 (N_17693,N_13279,N_14052);
or U17694 (N_17694,N_13926,N_13417);
or U17695 (N_17695,N_12757,N_13888);
nor U17696 (N_17696,N_14514,N_15550);
xor U17697 (N_17697,N_14404,N_14100);
or U17698 (N_17698,N_12882,N_14682);
and U17699 (N_17699,N_13584,N_13799);
or U17700 (N_17700,N_15077,N_12543);
nor U17701 (N_17701,N_13511,N_12918);
or U17702 (N_17702,N_13286,N_12816);
or U17703 (N_17703,N_15283,N_15450);
nand U17704 (N_17704,N_13716,N_13213);
nor U17705 (N_17705,N_15309,N_14421);
or U17706 (N_17706,N_13692,N_12872);
or U17707 (N_17707,N_14037,N_15360);
nand U17708 (N_17708,N_14096,N_12772);
nand U17709 (N_17709,N_12519,N_13129);
or U17710 (N_17710,N_12934,N_13326);
and U17711 (N_17711,N_14050,N_15222);
and U17712 (N_17712,N_13308,N_13491);
xor U17713 (N_17713,N_12705,N_14043);
and U17714 (N_17714,N_13360,N_12745);
nor U17715 (N_17715,N_13777,N_13234);
nor U17716 (N_17716,N_12821,N_13098);
xnor U17717 (N_17717,N_12883,N_13148);
or U17718 (N_17718,N_13425,N_15224);
or U17719 (N_17719,N_13578,N_15000);
and U17720 (N_17720,N_15308,N_13089);
or U17721 (N_17721,N_15240,N_14947);
nand U17722 (N_17722,N_14433,N_15512);
or U17723 (N_17723,N_14998,N_14377);
xor U17724 (N_17724,N_13035,N_15159);
and U17725 (N_17725,N_14686,N_13741);
nand U17726 (N_17726,N_14981,N_13214);
nand U17727 (N_17727,N_14957,N_15282);
or U17728 (N_17728,N_13570,N_14066);
nor U17729 (N_17729,N_13299,N_12820);
xnor U17730 (N_17730,N_13358,N_12995);
or U17731 (N_17731,N_14992,N_12577);
nor U17732 (N_17732,N_14683,N_12539);
nor U17733 (N_17733,N_13171,N_15030);
nor U17734 (N_17734,N_13859,N_12975);
nand U17735 (N_17735,N_14978,N_14991);
or U17736 (N_17736,N_15241,N_15322);
nand U17737 (N_17737,N_13625,N_13275);
nand U17738 (N_17738,N_14233,N_14785);
or U17739 (N_17739,N_14562,N_14306);
and U17740 (N_17740,N_13193,N_13153);
nand U17741 (N_17741,N_12511,N_14025);
or U17742 (N_17742,N_14845,N_13636);
xnor U17743 (N_17743,N_13875,N_13170);
and U17744 (N_17744,N_14356,N_12580);
or U17745 (N_17745,N_14498,N_15518);
nand U17746 (N_17746,N_14246,N_12950);
and U17747 (N_17747,N_13177,N_14113);
nor U17748 (N_17748,N_13655,N_15173);
nor U17749 (N_17749,N_13972,N_14423);
xor U17750 (N_17750,N_13863,N_12744);
and U17751 (N_17751,N_14279,N_12979);
nand U17752 (N_17752,N_14492,N_15541);
nor U17753 (N_17753,N_14548,N_14300);
and U17754 (N_17754,N_14580,N_15124);
and U17755 (N_17755,N_13705,N_13982);
xor U17756 (N_17756,N_14341,N_14951);
nor U17757 (N_17757,N_14572,N_12828);
or U17758 (N_17758,N_14936,N_14000);
and U17759 (N_17759,N_14858,N_13634);
nor U17760 (N_17760,N_12534,N_14220);
nand U17761 (N_17761,N_12744,N_13372);
nand U17762 (N_17762,N_14542,N_13868);
xor U17763 (N_17763,N_14109,N_14343);
or U17764 (N_17764,N_12825,N_13995);
nor U17765 (N_17765,N_13035,N_13574);
nand U17766 (N_17766,N_13545,N_12898);
or U17767 (N_17767,N_14230,N_14912);
nor U17768 (N_17768,N_15451,N_14902);
or U17769 (N_17769,N_15042,N_13676);
nand U17770 (N_17770,N_15237,N_13727);
and U17771 (N_17771,N_12565,N_14627);
and U17772 (N_17772,N_13199,N_14410);
nor U17773 (N_17773,N_14592,N_15620);
nand U17774 (N_17774,N_12554,N_12827);
nor U17775 (N_17775,N_15534,N_14181);
and U17776 (N_17776,N_14602,N_13706);
or U17777 (N_17777,N_13973,N_13182);
nor U17778 (N_17778,N_13650,N_12950);
and U17779 (N_17779,N_14412,N_13575);
or U17780 (N_17780,N_15334,N_13587);
or U17781 (N_17781,N_13318,N_15574);
nor U17782 (N_17782,N_15523,N_13851);
or U17783 (N_17783,N_15012,N_15391);
or U17784 (N_17784,N_13388,N_13635);
and U17785 (N_17785,N_13664,N_13220);
and U17786 (N_17786,N_13975,N_13159);
nor U17787 (N_17787,N_13302,N_12917);
nor U17788 (N_17788,N_15591,N_12580);
nor U17789 (N_17789,N_14678,N_12918);
nor U17790 (N_17790,N_13491,N_15523);
and U17791 (N_17791,N_13240,N_13198);
xor U17792 (N_17792,N_13320,N_14934);
nor U17793 (N_17793,N_12619,N_12949);
or U17794 (N_17794,N_14080,N_14307);
nand U17795 (N_17795,N_14487,N_14352);
and U17796 (N_17796,N_13045,N_13480);
nand U17797 (N_17797,N_15446,N_13410);
or U17798 (N_17798,N_13516,N_14366);
or U17799 (N_17799,N_15496,N_14194);
xor U17800 (N_17800,N_14300,N_14417);
nand U17801 (N_17801,N_14101,N_13120);
nor U17802 (N_17802,N_12882,N_15148);
or U17803 (N_17803,N_15135,N_15568);
and U17804 (N_17804,N_13654,N_13925);
and U17805 (N_17805,N_12975,N_13688);
nand U17806 (N_17806,N_15283,N_12692);
and U17807 (N_17807,N_14196,N_13082);
nor U17808 (N_17808,N_14231,N_12883);
nor U17809 (N_17809,N_14750,N_12789);
and U17810 (N_17810,N_15613,N_15321);
and U17811 (N_17811,N_13151,N_15198);
xnor U17812 (N_17812,N_14607,N_15162);
nor U17813 (N_17813,N_15025,N_15527);
nor U17814 (N_17814,N_12667,N_13794);
and U17815 (N_17815,N_14482,N_13861);
and U17816 (N_17816,N_14987,N_14016);
xor U17817 (N_17817,N_13391,N_13075);
nand U17818 (N_17818,N_13170,N_15059);
nor U17819 (N_17819,N_14840,N_14917);
xor U17820 (N_17820,N_13092,N_14674);
nor U17821 (N_17821,N_15414,N_12778);
and U17822 (N_17822,N_13653,N_13928);
nor U17823 (N_17823,N_12855,N_15456);
or U17824 (N_17824,N_14384,N_15196);
or U17825 (N_17825,N_14362,N_13698);
or U17826 (N_17826,N_12645,N_13539);
and U17827 (N_17827,N_12832,N_15284);
or U17828 (N_17828,N_13280,N_13495);
nand U17829 (N_17829,N_13101,N_13471);
nand U17830 (N_17830,N_13259,N_13751);
nand U17831 (N_17831,N_14682,N_12726);
and U17832 (N_17832,N_14571,N_14136);
and U17833 (N_17833,N_14447,N_14319);
nor U17834 (N_17834,N_14076,N_13439);
nand U17835 (N_17835,N_15012,N_14563);
or U17836 (N_17836,N_14409,N_12679);
nor U17837 (N_17837,N_12561,N_14914);
nor U17838 (N_17838,N_13781,N_14128);
nor U17839 (N_17839,N_14264,N_13567);
nand U17840 (N_17840,N_15619,N_14679);
xnor U17841 (N_17841,N_13766,N_15462);
or U17842 (N_17842,N_15564,N_13683);
nor U17843 (N_17843,N_13665,N_15430);
nand U17844 (N_17844,N_13263,N_14833);
nor U17845 (N_17845,N_13394,N_14557);
nor U17846 (N_17846,N_12506,N_12697);
nor U17847 (N_17847,N_13968,N_13576);
and U17848 (N_17848,N_14567,N_12715);
xnor U17849 (N_17849,N_13793,N_14332);
or U17850 (N_17850,N_12925,N_15414);
or U17851 (N_17851,N_13041,N_15610);
nand U17852 (N_17852,N_14942,N_14404);
nor U17853 (N_17853,N_13073,N_14206);
nand U17854 (N_17854,N_14361,N_15127);
and U17855 (N_17855,N_13597,N_14853);
nor U17856 (N_17856,N_12912,N_13230);
nand U17857 (N_17857,N_14853,N_13760);
nor U17858 (N_17858,N_14289,N_13962);
xnor U17859 (N_17859,N_14679,N_13565);
xnor U17860 (N_17860,N_15203,N_14876);
and U17861 (N_17861,N_13025,N_13079);
nand U17862 (N_17862,N_14552,N_14093);
or U17863 (N_17863,N_12678,N_15512);
or U17864 (N_17864,N_14315,N_14652);
xor U17865 (N_17865,N_14745,N_14675);
or U17866 (N_17866,N_12785,N_13499);
and U17867 (N_17867,N_14203,N_15070);
nor U17868 (N_17868,N_15614,N_13249);
or U17869 (N_17869,N_14170,N_14413);
or U17870 (N_17870,N_15463,N_15613);
nor U17871 (N_17871,N_15541,N_13900);
or U17872 (N_17872,N_15008,N_13115);
nor U17873 (N_17873,N_15609,N_15450);
xor U17874 (N_17874,N_13603,N_12595);
or U17875 (N_17875,N_12899,N_12806);
nand U17876 (N_17876,N_12851,N_13646);
nor U17877 (N_17877,N_12976,N_13520);
nor U17878 (N_17878,N_13847,N_14341);
and U17879 (N_17879,N_14856,N_14276);
nand U17880 (N_17880,N_13792,N_13230);
and U17881 (N_17881,N_13927,N_15117);
and U17882 (N_17882,N_13287,N_14289);
nor U17883 (N_17883,N_14651,N_14890);
or U17884 (N_17884,N_13523,N_15113);
and U17885 (N_17885,N_15017,N_15441);
or U17886 (N_17886,N_15374,N_14096);
nor U17887 (N_17887,N_15268,N_13220);
and U17888 (N_17888,N_15027,N_13752);
nand U17889 (N_17889,N_14554,N_14256);
nor U17890 (N_17890,N_12507,N_12769);
or U17891 (N_17891,N_12713,N_14332);
nand U17892 (N_17892,N_13229,N_13398);
or U17893 (N_17893,N_14062,N_15060);
nand U17894 (N_17894,N_15122,N_15369);
or U17895 (N_17895,N_14644,N_13197);
and U17896 (N_17896,N_14177,N_12797);
or U17897 (N_17897,N_12559,N_14317);
or U17898 (N_17898,N_15127,N_13789);
nand U17899 (N_17899,N_14625,N_12702);
nand U17900 (N_17900,N_15502,N_15605);
or U17901 (N_17901,N_14116,N_14917);
or U17902 (N_17902,N_14113,N_14458);
and U17903 (N_17903,N_13111,N_15488);
or U17904 (N_17904,N_13790,N_13985);
nor U17905 (N_17905,N_14938,N_14981);
or U17906 (N_17906,N_15175,N_12722);
and U17907 (N_17907,N_14899,N_13262);
nand U17908 (N_17908,N_14955,N_14576);
and U17909 (N_17909,N_14439,N_12673);
nand U17910 (N_17910,N_14506,N_14818);
nor U17911 (N_17911,N_14998,N_14162);
or U17912 (N_17912,N_15049,N_12637);
or U17913 (N_17913,N_15356,N_15433);
or U17914 (N_17914,N_14127,N_14021);
nor U17915 (N_17915,N_13229,N_13179);
xor U17916 (N_17916,N_12644,N_14590);
or U17917 (N_17917,N_13981,N_13480);
and U17918 (N_17918,N_13842,N_15210);
and U17919 (N_17919,N_13100,N_13336);
nor U17920 (N_17920,N_14125,N_12630);
nor U17921 (N_17921,N_15300,N_15427);
xor U17922 (N_17922,N_14237,N_14234);
or U17923 (N_17923,N_13448,N_13395);
xor U17924 (N_17924,N_13567,N_12783);
nand U17925 (N_17925,N_14124,N_13917);
and U17926 (N_17926,N_13017,N_13355);
nand U17927 (N_17927,N_13411,N_15237);
xor U17928 (N_17928,N_13955,N_15296);
or U17929 (N_17929,N_14677,N_13832);
and U17930 (N_17930,N_15139,N_12729);
and U17931 (N_17931,N_12832,N_12862);
or U17932 (N_17932,N_13568,N_13494);
nor U17933 (N_17933,N_15411,N_12764);
and U17934 (N_17934,N_13646,N_15184);
nor U17935 (N_17935,N_12746,N_14610);
nor U17936 (N_17936,N_14584,N_14759);
xor U17937 (N_17937,N_13743,N_15183);
nor U17938 (N_17938,N_13565,N_14299);
nand U17939 (N_17939,N_14295,N_12611);
nand U17940 (N_17940,N_14156,N_13920);
nor U17941 (N_17941,N_12599,N_13075);
or U17942 (N_17942,N_13876,N_13432);
nand U17943 (N_17943,N_15322,N_14395);
or U17944 (N_17944,N_15464,N_14774);
and U17945 (N_17945,N_15525,N_13536);
nand U17946 (N_17946,N_14265,N_15457);
xnor U17947 (N_17947,N_15296,N_15281);
nor U17948 (N_17948,N_14626,N_14056);
or U17949 (N_17949,N_14760,N_15489);
or U17950 (N_17950,N_14357,N_14711);
or U17951 (N_17951,N_14237,N_14191);
nor U17952 (N_17952,N_15048,N_14946);
xor U17953 (N_17953,N_13016,N_12635);
or U17954 (N_17954,N_14473,N_13055);
and U17955 (N_17955,N_13129,N_12549);
nand U17956 (N_17956,N_13724,N_14817);
xnor U17957 (N_17957,N_14386,N_13076);
nand U17958 (N_17958,N_12822,N_14391);
nor U17959 (N_17959,N_13854,N_13140);
nand U17960 (N_17960,N_14994,N_14401);
nand U17961 (N_17961,N_13302,N_15104);
xnor U17962 (N_17962,N_13877,N_13244);
or U17963 (N_17963,N_13023,N_12864);
or U17964 (N_17964,N_12567,N_14172);
nor U17965 (N_17965,N_14184,N_14186);
nand U17966 (N_17966,N_15489,N_13694);
nor U17967 (N_17967,N_15357,N_14120);
xor U17968 (N_17968,N_15495,N_15618);
or U17969 (N_17969,N_12701,N_13203);
nand U17970 (N_17970,N_12758,N_14540);
or U17971 (N_17971,N_14581,N_14862);
xor U17972 (N_17972,N_14643,N_14214);
and U17973 (N_17973,N_14359,N_15114);
nand U17974 (N_17974,N_14362,N_14998);
nor U17975 (N_17975,N_12923,N_15588);
or U17976 (N_17976,N_15102,N_12626);
nor U17977 (N_17977,N_14435,N_13616);
nand U17978 (N_17978,N_14766,N_15131);
or U17979 (N_17979,N_14933,N_14053);
nor U17980 (N_17980,N_13341,N_15327);
or U17981 (N_17981,N_14906,N_15149);
and U17982 (N_17982,N_13502,N_13923);
nor U17983 (N_17983,N_15619,N_12764);
and U17984 (N_17984,N_13250,N_13964);
and U17985 (N_17985,N_12549,N_13745);
xor U17986 (N_17986,N_14024,N_14326);
nor U17987 (N_17987,N_14619,N_13309);
nor U17988 (N_17988,N_14376,N_14383);
nand U17989 (N_17989,N_13521,N_15604);
or U17990 (N_17990,N_14564,N_13379);
or U17991 (N_17991,N_14283,N_15457);
and U17992 (N_17992,N_14264,N_13534);
and U17993 (N_17993,N_14684,N_13990);
or U17994 (N_17994,N_14851,N_13520);
nor U17995 (N_17995,N_15411,N_14570);
nand U17996 (N_17996,N_14719,N_13486);
nor U17997 (N_17997,N_13377,N_14198);
xnor U17998 (N_17998,N_14664,N_14015);
nand U17999 (N_17999,N_12757,N_14184);
or U18000 (N_18000,N_13177,N_14926);
nand U18001 (N_18001,N_15021,N_13470);
xnor U18002 (N_18002,N_15573,N_13544);
and U18003 (N_18003,N_13096,N_15614);
or U18004 (N_18004,N_15622,N_14942);
and U18005 (N_18005,N_14302,N_13393);
and U18006 (N_18006,N_14706,N_13740);
nand U18007 (N_18007,N_13078,N_14712);
nand U18008 (N_18008,N_13384,N_13908);
nand U18009 (N_18009,N_12564,N_13620);
and U18010 (N_18010,N_13737,N_15427);
and U18011 (N_18011,N_13982,N_14037);
nand U18012 (N_18012,N_14928,N_14252);
and U18013 (N_18013,N_14234,N_14206);
nor U18014 (N_18014,N_14221,N_15230);
nor U18015 (N_18015,N_15105,N_14306);
xor U18016 (N_18016,N_13498,N_12533);
nand U18017 (N_18017,N_14128,N_14508);
nand U18018 (N_18018,N_14361,N_14949);
nor U18019 (N_18019,N_12945,N_13497);
nor U18020 (N_18020,N_13853,N_14156);
or U18021 (N_18021,N_15457,N_15239);
nor U18022 (N_18022,N_13507,N_13914);
or U18023 (N_18023,N_13654,N_13450);
nand U18024 (N_18024,N_14181,N_14675);
nand U18025 (N_18025,N_14180,N_12720);
or U18026 (N_18026,N_14696,N_15396);
nor U18027 (N_18027,N_14013,N_14731);
nand U18028 (N_18028,N_13871,N_14015);
xnor U18029 (N_18029,N_14476,N_13478);
nor U18030 (N_18030,N_12951,N_12517);
nand U18031 (N_18031,N_14558,N_14724);
and U18032 (N_18032,N_15379,N_14501);
nor U18033 (N_18033,N_14659,N_14251);
or U18034 (N_18034,N_13475,N_15066);
and U18035 (N_18035,N_13917,N_14950);
nor U18036 (N_18036,N_14679,N_15155);
nand U18037 (N_18037,N_13560,N_14622);
nor U18038 (N_18038,N_15103,N_12571);
xnor U18039 (N_18039,N_12991,N_13298);
nor U18040 (N_18040,N_15542,N_13305);
nor U18041 (N_18041,N_13703,N_14572);
and U18042 (N_18042,N_12590,N_12598);
xnor U18043 (N_18043,N_12998,N_13699);
nand U18044 (N_18044,N_15303,N_14998);
and U18045 (N_18045,N_12514,N_13994);
and U18046 (N_18046,N_12503,N_13833);
nand U18047 (N_18047,N_15481,N_14748);
or U18048 (N_18048,N_13859,N_12510);
and U18049 (N_18049,N_14227,N_13275);
or U18050 (N_18050,N_12827,N_14094);
and U18051 (N_18051,N_13496,N_13697);
and U18052 (N_18052,N_14962,N_12937);
nor U18053 (N_18053,N_12623,N_14307);
or U18054 (N_18054,N_12938,N_12718);
nand U18055 (N_18055,N_14308,N_15492);
xnor U18056 (N_18056,N_13264,N_15513);
and U18057 (N_18057,N_15227,N_13971);
xor U18058 (N_18058,N_13814,N_15339);
and U18059 (N_18059,N_12835,N_15393);
nand U18060 (N_18060,N_14391,N_14008);
nor U18061 (N_18061,N_14981,N_14077);
and U18062 (N_18062,N_14896,N_14752);
and U18063 (N_18063,N_13959,N_13643);
and U18064 (N_18064,N_15624,N_13494);
xor U18065 (N_18065,N_15515,N_12848);
and U18066 (N_18066,N_15351,N_14960);
nor U18067 (N_18067,N_14319,N_14565);
nor U18068 (N_18068,N_12923,N_15243);
or U18069 (N_18069,N_14867,N_12510);
nand U18070 (N_18070,N_13257,N_12644);
nor U18071 (N_18071,N_14331,N_15326);
and U18072 (N_18072,N_12567,N_14224);
nor U18073 (N_18073,N_14320,N_12607);
nand U18074 (N_18074,N_14493,N_14040);
and U18075 (N_18075,N_14284,N_14002);
nand U18076 (N_18076,N_12751,N_15086);
and U18077 (N_18077,N_13206,N_12749);
and U18078 (N_18078,N_13497,N_13970);
nand U18079 (N_18079,N_13978,N_15079);
nand U18080 (N_18080,N_13804,N_15056);
and U18081 (N_18081,N_15301,N_14100);
or U18082 (N_18082,N_13319,N_13385);
nor U18083 (N_18083,N_13997,N_12568);
nor U18084 (N_18084,N_13398,N_14334);
nand U18085 (N_18085,N_14770,N_14296);
and U18086 (N_18086,N_14432,N_13449);
nor U18087 (N_18087,N_14599,N_13819);
and U18088 (N_18088,N_15193,N_12902);
nand U18089 (N_18089,N_12618,N_14199);
nor U18090 (N_18090,N_14453,N_15479);
and U18091 (N_18091,N_14983,N_12579);
and U18092 (N_18092,N_14595,N_13449);
nand U18093 (N_18093,N_13045,N_15596);
or U18094 (N_18094,N_12863,N_14156);
nand U18095 (N_18095,N_12574,N_13157);
or U18096 (N_18096,N_14716,N_12878);
or U18097 (N_18097,N_14550,N_12532);
and U18098 (N_18098,N_12752,N_12539);
and U18099 (N_18099,N_13991,N_12937);
and U18100 (N_18100,N_15016,N_13783);
and U18101 (N_18101,N_13278,N_13628);
xnor U18102 (N_18102,N_14726,N_14751);
and U18103 (N_18103,N_14233,N_12802);
xor U18104 (N_18104,N_14536,N_14727);
xor U18105 (N_18105,N_15242,N_14307);
and U18106 (N_18106,N_12726,N_15132);
nor U18107 (N_18107,N_14712,N_14219);
or U18108 (N_18108,N_15525,N_13453);
xnor U18109 (N_18109,N_14372,N_14143);
nor U18110 (N_18110,N_14669,N_13803);
and U18111 (N_18111,N_14818,N_13483);
and U18112 (N_18112,N_13953,N_13324);
xnor U18113 (N_18113,N_13141,N_12946);
nand U18114 (N_18114,N_12921,N_13095);
nand U18115 (N_18115,N_14471,N_14366);
and U18116 (N_18116,N_13079,N_13626);
or U18117 (N_18117,N_15559,N_13587);
and U18118 (N_18118,N_13545,N_13130);
or U18119 (N_18119,N_15017,N_14989);
xor U18120 (N_18120,N_15347,N_13029);
or U18121 (N_18121,N_14295,N_14620);
xnor U18122 (N_18122,N_14254,N_13968);
nor U18123 (N_18123,N_14424,N_12885);
or U18124 (N_18124,N_13211,N_12629);
nor U18125 (N_18125,N_13967,N_13522);
or U18126 (N_18126,N_13001,N_13992);
xnor U18127 (N_18127,N_13696,N_14439);
and U18128 (N_18128,N_12876,N_14737);
nor U18129 (N_18129,N_14595,N_13191);
and U18130 (N_18130,N_12739,N_15013);
nor U18131 (N_18131,N_15229,N_13710);
or U18132 (N_18132,N_12779,N_14383);
or U18133 (N_18133,N_14795,N_12802);
or U18134 (N_18134,N_13701,N_14724);
nor U18135 (N_18135,N_12582,N_15159);
or U18136 (N_18136,N_15277,N_13487);
or U18137 (N_18137,N_14661,N_13401);
nor U18138 (N_18138,N_13195,N_14584);
nor U18139 (N_18139,N_14331,N_14830);
nand U18140 (N_18140,N_13127,N_13772);
xor U18141 (N_18141,N_12665,N_14610);
nor U18142 (N_18142,N_14367,N_13945);
nand U18143 (N_18143,N_15261,N_13934);
or U18144 (N_18144,N_13747,N_15588);
or U18145 (N_18145,N_14998,N_15174);
nor U18146 (N_18146,N_13058,N_15388);
nor U18147 (N_18147,N_15081,N_14734);
and U18148 (N_18148,N_13850,N_14795);
or U18149 (N_18149,N_14755,N_14035);
nor U18150 (N_18150,N_15472,N_14789);
nor U18151 (N_18151,N_12758,N_13977);
xnor U18152 (N_18152,N_13934,N_15169);
or U18153 (N_18153,N_14052,N_15249);
nor U18154 (N_18154,N_15483,N_15037);
nand U18155 (N_18155,N_13189,N_14711);
nand U18156 (N_18156,N_14266,N_14478);
nand U18157 (N_18157,N_14918,N_14378);
nor U18158 (N_18158,N_12997,N_13668);
or U18159 (N_18159,N_13396,N_14049);
nor U18160 (N_18160,N_13849,N_13551);
or U18161 (N_18161,N_13837,N_14217);
and U18162 (N_18162,N_13106,N_13453);
or U18163 (N_18163,N_14625,N_15326);
or U18164 (N_18164,N_14668,N_13429);
or U18165 (N_18165,N_14335,N_14399);
nand U18166 (N_18166,N_15403,N_14277);
or U18167 (N_18167,N_14615,N_15072);
and U18168 (N_18168,N_13391,N_14113);
nand U18169 (N_18169,N_12907,N_14472);
nand U18170 (N_18170,N_14089,N_15484);
and U18171 (N_18171,N_14083,N_14035);
and U18172 (N_18172,N_14554,N_12745);
and U18173 (N_18173,N_14380,N_14804);
xor U18174 (N_18174,N_14954,N_14224);
and U18175 (N_18175,N_15561,N_13969);
xnor U18176 (N_18176,N_12881,N_14956);
nand U18177 (N_18177,N_13615,N_13425);
nand U18178 (N_18178,N_12727,N_14677);
and U18179 (N_18179,N_14566,N_14836);
nand U18180 (N_18180,N_13526,N_14647);
and U18181 (N_18181,N_14045,N_14549);
nor U18182 (N_18182,N_12843,N_13671);
nand U18183 (N_18183,N_13278,N_13403);
nand U18184 (N_18184,N_13133,N_15545);
or U18185 (N_18185,N_14360,N_12872);
nor U18186 (N_18186,N_13360,N_15342);
or U18187 (N_18187,N_14857,N_12582);
or U18188 (N_18188,N_12650,N_15564);
or U18189 (N_18189,N_12515,N_12942);
and U18190 (N_18190,N_15352,N_13255);
or U18191 (N_18191,N_15565,N_13498);
and U18192 (N_18192,N_13746,N_14698);
nor U18193 (N_18193,N_13879,N_14819);
or U18194 (N_18194,N_15165,N_13051);
nor U18195 (N_18195,N_14839,N_14632);
xnor U18196 (N_18196,N_13300,N_14649);
xor U18197 (N_18197,N_13210,N_13148);
and U18198 (N_18198,N_15032,N_13857);
nor U18199 (N_18199,N_15001,N_14237);
nand U18200 (N_18200,N_13788,N_13417);
or U18201 (N_18201,N_14170,N_13606);
nand U18202 (N_18202,N_13096,N_14234);
or U18203 (N_18203,N_14074,N_12937);
and U18204 (N_18204,N_14234,N_15116);
and U18205 (N_18205,N_13236,N_13873);
xor U18206 (N_18206,N_15085,N_13193);
nor U18207 (N_18207,N_12821,N_13457);
or U18208 (N_18208,N_12631,N_14372);
nand U18209 (N_18209,N_13274,N_14886);
or U18210 (N_18210,N_13024,N_13528);
nor U18211 (N_18211,N_15456,N_14914);
nand U18212 (N_18212,N_12660,N_14663);
nand U18213 (N_18213,N_12991,N_12906);
or U18214 (N_18214,N_13025,N_12787);
or U18215 (N_18215,N_13175,N_14000);
nor U18216 (N_18216,N_12883,N_14707);
nor U18217 (N_18217,N_14436,N_14429);
xnor U18218 (N_18218,N_13600,N_12500);
and U18219 (N_18219,N_15527,N_13884);
nor U18220 (N_18220,N_13100,N_14979);
and U18221 (N_18221,N_12964,N_14189);
and U18222 (N_18222,N_12529,N_12872);
xor U18223 (N_18223,N_13915,N_12661);
nor U18224 (N_18224,N_12783,N_14110);
or U18225 (N_18225,N_15597,N_13400);
or U18226 (N_18226,N_14072,N_13195);
or U18227 (N_18227,N_13474,N_13784);
nand U18228 (N_18228,N_14218,N_13786);
and U18229 (N_18229,N_15244,N_15072);
and U18230 (N_18230,N_14867,N_13971);
nand U18231 (N_18231,N_14670,N_15217);
nor U18232 (N_18232,N_12991,N_13335);
nor U18233 (N_18233,N_13221,N_13233);
xor U18234 (N_18234,N_13712,N_13772);
xnor U18235 (N_18235,N_13425,N_15612);
nand U18236 (N_18236,N_13967,N_15359);
nor U18237 (N_18237,N_12707,N_15290);
or U18238 (N_18238,N_12796,N_12799);
nand U18239 (N_18239,N_15280,N_13962);
or U18240 (N_18240,N_13598,N_13624);
and U18241 (N_18241,N_14920,N_13348);
and U18242 (N_18242,N_12509,N_14495);
nand U18243 (N_18243,N_15502,N_13281);
nor U18244 (N_18244,N_13206,N_15402);
and U18245 (N_18245,N_15268,N_15032);
nand U18246 (N_18246,N_14731,N_12852);
or U18247 (N_18247,N_14392,N_15570);
nor U18248 (N_18248,N_13257,N_15605);
and U18249 (N_18249,N_14959,N_14860);
nand U18250 (N_18250,N_13398,N_14106);
nor U18251 (N_18251,N_12933,N_12592);
and U18252 (N_18252,N_12761,N_13595);
or U18253 (N_18253,N_13587,N_15365);
nand U18254 (N_18254,N_15092,N_13716);
and U18255 (N_18255,N_12530,N_15269);
and U18256 (N_18256,N_15430,N_13779);
nand U18257 (N_18257,N_12984,N_13073);
or U18258 (N_18258,N_13859,N_13766);
nor U18259 (N_18259,N_13957,N_14643);
nand U18260 (N_18260,N_12891,N_14358);
or U18261 (N_18261,N_12831,N_12672);
nor U18262 (N_18262,N_13710,N_13911);
and U18263 (N_18263,N_14232,N_13892);
or U18264 (N_18264,N_15368,N_14236);
nor U18265 (N_18265,N_13740,N_15298);
nand U18266 (N_18266,N_14354,N_13048);
or U18267 (N_18267,N_13847,N_15089);
or U18268 (N_18268,N_14702,N_12690);
xor U18269 (N_18269,N_13635,N_13339);
and U18270 (N_18270,N_15522,N_15374);
and U18271 (N_18271,N_14856,N_12783);
xor U18272 (N_18272,N_13248,N_15311);
nor U18273 (N_18273,N_15132,N_13424);
nor U18274 (N_18274,N_14115,N_14469);
and U18275 (N_18275,N_13360,N_14893);
nor U18276 (N_18276,N_15447,N_14602);
or U18277 (N_18277,N_13650,N_14667);
xor U18278 (N_18278,N_14954,N_15455);
nand U18279 (N_18279,N_14007,N_15255);
or U18280 (N_18280,N_14753,N_15096);
nand U18281 (N_18281,N_13736,N_12545);
and U18282 (N_18282,N_15618,N_13602);
nand U18283 (N_18283,N_12915,N_12787);
nor U18284 (N_18284,N_14367,N_13287);
or U18285 (N_18285,N_15192,N_14356);
nand U18286 (N_18286,N_14581,N_15512);
and U18287 (N_18287,N_14479,N_14426);
nor U18288 (N_18288,N_14642,N_14064);
or U18289 (N_18289,N_15396,N_14363);
nand U18290 (N_18290,N_14606,N_14378);
nand U18291 (N_18291,N_15554,N_14589);
or U18292 (N_18292,N_14922,N_13625);
nand U18293 (N_18293,N_14583,N_12926);
and U18294 (N_18294,N_13605,N_14945);
nand U18295 (N_18295,N_12962,N_12689);
and U18296 (N_18296,N_13778,N_14270);
or U18297 (N_18297,N_14408,N_14391);
and U18298 (N_18298,N_14884,N_14051);
or U18299 (N_18299,N_12815,N_14316);
and U18300 (N_18300,N_15298,N_13896);
nor U18301 (N_18301,N_14814,N_14402);
nand U18302 (N_18302,N_13180,N_14221);
nand U18303 (N_18303,N_15390,N_13633);
or U18304 (N_18304,N_13668,N_13724);
and U18305 (N_18305,N_15056,N_13797);
and U18306 (N_18306,N_13116,N_14649);
and U18307 (N_18307,N_13609,N_15317);
nor U18308 (N_18308,N_14855,N_14673);
or U18309 (N_18309,N_15302,N_13995);
xnor U18310 (N_18310,N_14853,N_12564);
nor U18311 (N_18311,N_13143,N_12611);
nor U18312 (N_18312,N_14729,N_13112);
nor U18313 (N_18313,N_12581,N_13818);
and U18314 (N_18314,N_14215,N_13972);
nand U18315 (N_18315,N_14343,N_14420);
nand U18316 (N_18316,N_12550,N_13936);
nor U18317 (N_18317,N_14611,N_13276);
xor U18318 (N_18318,N_14703,N_13359);
and U18319 (N_18319,N_13730,N_12730);
and U18320 (N_18320,N_13444,N_15429);
nor U18321 (N_18321,N_13092,N_14317);
and U18322 (N_18322,N_14812,N_13485);
nand U18323 (N_18323,N_13591,N_15356);
and U18324 (N_18324,N_13269,N_13061);
xnor U18325 (N_18325,N_14698,N_13979);
nor U18326 (N_18326,N_14257,N_14923);
or U18327 (N_18327,N_13101,N_13394);
or U18328 (N_18328,N_14753,N_13521);
nor U18329 (N_18329,N_15074,N_14167);
and U18330 (N_18330,N_15025,N_13184);
nand U18331 (N_18331,N_12677,N_14071);
nand U18332 (N_18332,N_15559,N_13668);
nand U18333 (N_18333,N_13412,N_13163);
nand U18334 (N_18334,N_13546,N_14499);
or U18335 (N_18335,N_15015,N_13249);
nor U18336 (N_18336,N_13298,N_12661);
and U18337 (N_18337,N_13335,N_12917);
nand U18338 (N_18338,N_13638,N_15186);
or U18339 (N_18339,N_13845,N_15390);
nor U18340 (N_18340,N_12877,N_13537);
or U18341 (N_18341,N_13870,N_12785);
nor U18342 (N_18342,N_14356,N_13522);
and U18343 (N_18343,N_12726,N_14458);
or U18344 (N_18344,N_14744,N_13352);
and U18345 (N_18345,N_15528,N_13009);
nand U18346 (N_18346,N_15451,N_13541);
and U18347 (N_18347,N_12876,N_13558);
or U18348 (N_18348,N_15502,N_15558);
or U18349 (N_18349,N_15535,N_14086);
xnor U18350 (N_18350,N_15325,N_14342);
nand U18351 (N_18351,N_13583,N_13906);
nand U18352 (N_18352,N_14789,N_13540);
nor U18353 (N_18353,N_13457,N_13795);
and U18354 (N_18354,N_13061,N_13773);
nand U18355 (N_18355,N_15350,N_13170);
or U18356 (N_18356,N_14371,N_15167);
or U18357 (N_18357,N_13724,N_14055);
nor U18358 (N_18358,N_12515,N_14550);
or U18359 (N_18359,N_14978,N_12534);
nor U18360 (N_18360,N_14192,N_14893);
xor U18361 (N_18361,N_12733,N_15197);
nor U18362 (N_18362,N_14171,N_13463);
nand U18363 (N_18363,N_15350,N_14704);
or U18364 (N_18364,N_14315,N_15347);
or U18365 (N_18365,N_12644,N_13549);
or U18366 (N_18366,N_14213,N_13155);
and U18367 (N_18367,N_13889,N_14435);
and U18368 (N_18368,N_13380,N_12952);
or U18369 (N_18369,N_12881,N_15254);
or U18370 (N_18370,N_13118,N_13229);
xor U18371 (N_18371,N_13882,N_15551);
nor U18372 (N_18372,N_13187,N_13947);
nor U18373 (N_18373,N_14162,N_14450);
xor U18374 (N_18374,N_15314,N_14171);
nor U18375 (N_18375,N_14386,N_13631);
or U18376 (N_18376,N_15138,N_14927);
and U18377 (N_18377,N_15230,N_12970);
nor U18378 (N_18378,N_13855,N_13627);
and U18379 (N_18379,N_14523,N_15032);
nor U18380 (N_18380,N_15516,N_15620);
nor U18381 (N_18381,N_14584,N_13255);
and U18382 (N_18382,N_15048,N_15264);
and U18383 (N_18383,N_15223,N_15397);
and U18384 (N_18384,N_13280,N_13078);
nor U18385 (N_18385,N_13406,N_14562);
nor U18386 (N_18386,N_12694,N_13295);
or U18387 (N_18387,N_12917,N_15318);
nor U18388 (N_18388,N_13768,N_15406);
or U18389 (N_18389,N_15146,N_12751);
and U18390 (N_18390,N_13334,N_13775);
nor U18391 (N_18391,N_15402,N_13095);
nor U18392 (N_18392,N_13061,N_13284);
nor U18393 (N_18393,N_15496,N_14209);
or U18394 (N_18394,N_13037,N_13736);
or U18395 (N_18395,N_15281,N_12735);
xnor U18396 (N_18396,N_13144,N_14125);
nand U18397 (N_18397,N_13347,N_15097);
and U18398 (N_18398,N_15095,N_13354);
nor U18399 (N_18399,N_14680,N_15532);
and U18400 (N_18400,N_13466,N_13965);
xnor U18401 (N_18401,N_14542,N_13332);
or U18402 (N_18402,N_12575,N_15389);
and U18403 (N_18403,N_14524,N_13670);
nand U18404 (N_18404,N_13871,N_12952);
xnor U18405 (N_18405,N_13681,N_13572);
or U18406 (N_18406,N_14763,N_14739);
nor U18407 (N_18407,N_15002,N_12590);
and U18408 (N_18408,N_13171,N_13884);
xor U18409 (N_18409,N_13956,N_12951);
nand U18410 (N_18410,N_15329,N_13605);
xor U18411 (N_18411,N_13880,N_12877);
or U18412 (N_18412,N_12719,N_15520);
and U18413 (N_18413,N_15103,N_12716);
or U18414 (N_18414,N_14195,N_14560);
or U18415 (N_18415,N_14130,N_13698);
or U18416 (N_18416,N_13423,N_13884);
nand U18417 (N_18417,N_12718,N_15005);
nor U18418 (N_18418,N_13188,N_13581);
nand U18419 (N_18419,N_13593,N_13141);
nand U18420 (N_18420,N_13609,N_12624);
and U18421 (N_18421,N_14348,N_14272);
nor U18422 (N_18422,N_12553,N_13256);
or U18423 (N_18423,N_12770,N_14255);
or U18424 (N_18424,N_13837,N_12909);
xor U18425 (N_18425,N_12623,N_12665);
and U18426 (N_18426,N_13079,N_15316);
and U18427 (N_18427,N_13721,N_13181);
nand U18428 (N_18428,N_14596,N_12901);
nand U18429 (N_18429,N_15219,N_13507);
nor U18430 (N_18430,N_13451,N_14452);
nor U18431 (N_18431,N_13941,N_13623);
xor U18432 (N_18432,N_14652,N_12921);
or U18433 (N_18433,N_14456,N_12588);
nand U18434 (N_18434,N_13634,N_15369);
or U18435 (N_18435,N_13989,N_13128);
and U18436 (N_18436,N_15129,N_14086);
xor U18437 (N_18437,N_12546,N_14309);
or U18438 (N_18438,N_12943,N_13672);
nor U18439 (N_18439,N_13220,N_14388);
and U18440 (N_18440,N_14039,N_13541);
xnor U18441 (N_18441,N_12668,N_15182);
nand U18442 (N_18442,N_12887,N_15111);
nor U18443 (N_18443,N_13067,N_14227);
nand U18444 (N_18444,N_13450,N_13330);
and U18445 (N_18445,N_12658,N_13839);
and U18446 (N_18446,N_15230,N_14015);
nand U18447 (N_18447,N_14390,N_14862);
nand U18448 (N_18448,N_14991,N_12874);
or U18449 (N_18449,N_12817,N_15519);
nand U18450 (N_18450,N_14626,N_14700);
xor U18451 (N_18451,N_15411,N_12538);
and U18452 (N_18452,N_13443,N_13624);
nand U18453 (N_18453,N_14723,N_12961);
nand U18454 (N_18454,N_13901,N_13075);
or U18455 (N_18455,N_13719,N_14967);
nor U18456 (N_18456,N_12955,N_15576);
and U18457 (N_18457,N_15504,N_14534);
nor U18458 (N_18458,N_15109,N_14561);
xor U18459 (N_18459,N_14299,N_13731);
or U18460 (N_18460,N_15048,N_13864);
and U18461 (N_18461,N_13650,N_13085);
nor U18462 (N_18462,N_15116,N_14066);
nor U18463 (N_18463,N_14299,N_13204);
nand U18464 (N_18464,N_13424,N_12636);
or U18465 (N_18465,N_13817,N_12576);
and U18466 (N_18466,N_13417,N_15148);
xor U18467 (N_18467,N_14562,N_15169);
or U18468 (N_18468,N_12935,N_13758);
or U18469 (N_18469,N_14901,N_15244);
and U18470 (N_18470,N_14015,N_13961);
nor U18471 (N_18471,N_13424,N_12908);
and U18472 (N_18472,N_12843,N_12913);
or U18473 (N_18473,N_15448,N_14987);
and U18474 (N_18474,N_15148,N_15335);
xor U18475 (N_18475,N_14777,N_12952);
nand U18476 (N_18476,N_15340,N_15267);
or U18477 (N_18477,N_13696,N_13771);
and U18478 (N_18478,N_13301,N_12636);
nor U18479 (N_18479,N_15066,N_12858);
or U18480 (N_18480,N_12714,N_14601);
nand U18481 (N_18481,N_14193,N_13543);
or U18482 (N_18482,N_14633,N_14425);
or U18483 (N_18483,N_14486,N_14523);
nor U18484 (N_18484,N_14862,N_13457);
nand U18485 (N_18485,N_13830,N_13108);
nand U18486 (N_18486,N_14437,N_15535);
nor U18487 (N_18487,N_13494,N_14391);
or U18488 (N_18488,N_15351,N_14785);
and U18489 (N_18489,N_13851,N_13055);
xor U18490 (N_18490,N_15481,N_13197);
xnor U18491 (N_18491,N_12859,N_15393);
or U18492 (N_18492,N_15033,N_15325);
nor U18493 (N_18493,N_14308,N_14794);
nor U18494 (N_18494,N_15231,N_13424);
or U18495 (N_18495,N_14178,N_12627);
nor U18496 (N_18496,N_12964,N_14843);
nand U18497 (N_18497,N_12894,N_15591);
nor U18498 (N_18498,N_13816,N_14232);
nand U18499 (N_18499,N_15342,N_12600);
nor U18500 (N_18500,N_13216,N_14752);
nor U18501 (N_18501,N_15171,N_15176);
nor U18502 (N_18502,N_14521,N_15442);
nand U18503 (N_18503,N_13738,N_14956);
nand U18504 (N_18504,N_13013,N_15277);
and U18505 (N_18505,N_14517,N_14282);
xnor U18506 (N_18506,N_14217,N_14897);
nand U18507 (N_18507,N_13631,N_13275);
and U18508 (N_18508,N_13011,N_14432);
and U18509 (N_18509,N_14411,N_14488);
nand U18510 (N_18510,N_13042,N_13159);
xor U18511 (N_18511,N_15538,N_15618);
nand U18512 (N_18512,N_14165,N_13904);
xnor U18513 (N_18513,N_14124,N_15345);
and U18514 (N_18514,N_15383,N_15394);
and U18515 (N_18515,N_14552,N_15375);
or U18516 (N_18516,N_13815,N_14523);
or U18517 (N_18517,N_12698,N_13113);
nand U18518 (N_18518,N_13818,N_12552);
or U18519 (N_18519,N_13774,N_13094);
and U18520 (N_18520,N_13080,N_13381);
nor U18521 (N_18521,N_12755,N_12704);
or U18522 (N_18522,N_14603,N_12502);
nand U18523 (N_18523,N_15582,N_13525);
nand U18524 (N_18524,N_13068,N_15391);
nor U18525 (N_18525,N_15375,N_15607);
nand U18526 (N_18526,N_15159,N_14993);
nand U18527 (N_18527,N_13059,N_13749);
or U18528 (N_18528,N_12862,N_13418);
and U18529 (N_18529,N_13673,N_13901);
nor U18530 (N_18530,N_13462,N_14889);
nand U18531 (N_18531,N_14293,N_14480);
or U18532 (N_18532,N_13555,N_14221);
nand U18533 (N_18533,N_13435,N_14678);
nand U18534 (N_18534,N_13018,N_14784);
and U18535 (N_18535,N_13461,N_12578);
nand U18536 (N_18536,N_13225,N_14678);
nor U18537 (N_18537,N_13541,N_15498);
nand U18538 (N_18538,N_13526,N_15272);
nand U18539 (N_18539,N_13515,N_13065);
nand U18540 (N_18540,N_12923,N_14858);
and U18541 (N_18541,N_14141,N_14291);
nand U18542 (N_18542,N_12559,N_14224);
xor U18543 (N_18543,N_13508,N_14694);
and U18544 (N_18544,N_15170,N_15480);
and U18545 (N_18545,N_13704,N_14236);
xnor U18546 (N_18546,N_12545,N_14525);
nand U18547 (N_18547,N_14817,N_14528);
and U18548 (N_18548,N_14664,N_15254);
and U18549 (N_18549,N_14561,N_15438);
nor U18550 (N_18550,N_13492,N_14904);
or U18551 (N_18551,N_13885,N_14475);
nand U18552 (N_18552,N_14421,N_14222);
nor U18553 (N_18553,N_12679,N_15356);
or U18554 (N_18554,N_14553,N_13806);
nor U18555 (N_18555,N_15464,N_15528);
nor U18556 (N_18556,N_13266,N_14986);
or U18557 (N_18557,N_13411,N_13366);
and U18558 (N_18558,N_14860,N_13001);
and U18559 (N_18559,N_15055,N_15604);
or U18560 (N_18560,N_13119,N_13161);
and U18561 (N_18561,N_15397,N_14325);
or U18562 (N_18562,N_14172,N_13370);
nor U18563 (N_18563,N_14413,N_12788);
nand U18564 (N_18564,N_15480,N_14305);
and U18565 (N_18565,N_13823,N_15219);
nand U18566 (N_18566,N_12771,N_14540);
nor U18567 (N_18567,N_15054,N_12522);
nand U18568 (N_18568,N_15371,N_13475);
nand U18569 (N_18569,N_13514,N_12572);
and U18570 (N_18570,N_13302,N_14375);
nor U18571 (N_18571,N_15296,N_12860);
and U18572 (N_18572,N_13934,N_15077);
or U18573 (N_18573,N_14404,N_12510);
or U18574 (N_18574,N_13816,N_13248);
nor U18575 (N_18575,N_13428,N_15289);
xor U18576 (N_18576,N_14845,N_14684);
or U18577 (N_18577,N_12881,N_13667);
and U18578 (N_18578,N_13245,N_15598);
nand U18579 (N_18579,N_13671,N_14660);
nor U18580 (N_18580,N_13763,N_13162);
and U18581 (N_18581,N_12614,N_14112);
nand U18582 (N_18582,N_13284,N_15256);
or U18583 (N_18583,N_13995,N_13455);
or U18584 (N_18584,N_14312,N_14479);
and U18585 (N_18585,N_14642,N_13944);
and U18586 (N_18586,N_15514,N_12795);
and U18587 (N_18587,N_13557,N_13107);
and U18588 (N_18588,N_13636,N_14324);
nor U18589 (N_18589,N_15150,N_14214);
or U18590 (N_18590,N_12609,N_14864);
nor U18591 (N_18591,N_14107,N_15227);
and U18592 (N_18592,N_14261,N_14088);
or U18593 (N_18593,N_15211,N_14227);
nor U18594 (N_18594,N_14563,N_14266);
nand U18595 (N_18595,N_14645,N_15327);
or U18596 (N_18596,N_13421,N_13089);
nor U18597 (N_18597,N_15332,N_13303);
and U18598 (N_18598,N_13467,N_14846);
xor U18599 (N_18599,N_13195,N_15130);
nand U18600 (N_18600,N_13923,N_14774);
or U18601 (N_18601,N_15147,N_12726);
nor U18602 (N_18602,N_13598,N_13663);
nor U18603 (N_18603,N_15486,N_13308);
or U18604 (N_18604,N_15037,N_13338);
nand U18605 (N_18605,N_13893,N_15162);
nor U18606 (N_18606,N_15554,N_14230);
nand U18607 (N_18607,N_15201,N_15139);
or U18608 (N_18608,N_14651,N_13517);
and U18609 (N_18609,N_15178,N_15151);
nand U18610 (N_18610,N_14596,N_13808);
or U18611 (N_18611,N_14732,N_15054);
or U18612 (N_18612,N_13916,N_14527);
or U18613 (N_18613,N_15491,N_13297);
nor U18614 (N_18614,N_14607,N_13032);
nand U18615 (N_18615,N_15448,N_12772);
nor U18616 (N_18616,N_15602,N_14728);
nor U18617 (N_18617,N_13308,N_12961);
and U18618 (N_18618,N_15255,N_14725);
xor U18619 (N_18619,N_14963,N_13488);
xnor U18620 (N_18620,N_13247,N_13847);
xor U18621 (N_18621,N_13329,N_12594);
or U18622 (N_18622,N_15057,N_14344);
or U18623 (N_18623,N_12841,N_13685);
or U18624 (N_18624,N_14209,N_14128);
and U18625 (N_18625,N_13374,N_14572);
nor U18626 (N_18626,N_15613,N_12619);
nor U18627 (N_18627,N_13578,N_13027);
xnor U18628 (N_18628,N_14946,N_13041);
nand U18629 (N_18629,N_13733,N_14002);
and U18630 (N_18630,N_12727,N_13725);
nor U18631 (N_18631,N_14517,N_13601);
and U18632 (N_18632,N_15505,N_13669);
or U18633 (N_18633,N_14012,N_13255);
and U18634 (N_18634,N_14247,N_13555);
nor U18635 (N_18635,N_14063,N_13754);
nand U18636 (N_18636,N_13542,N_13530);
nand U18637 (N_18637,N_14289,N_14635);
nor U18638 (N_18638,N_13121,N_14379);
nand U18639 (N_18639,N_15586,N_12995);
and U18640 (N_18640,N_13485,N_14841);
nand U18641 (N_18641,N_12962,N_12759);
or U18642 (N_18642,N_13731,N_14348);
and U18643 (N_18643,N_13870,N_13142);
or U18644 (N_18644,N_14324,N_15615);
and U18645 (N_18645,N_13235,N_12974);
or U18646 (N_18646,N_12537,N_12719);
and U18647 (N_18647,N_14129,N_14101);
nand U18648 (N_18648,N_14686,N_14334);
nor U18649 (N_18649,N_12780,N_14723);
or U18650 (N_18650,N_13308,N_14870);
or U18651 (N_18651,N_14709,N_12674);
or U18652 (N_18652,N_15249,N_12782);
or U18653 (N_18653,N_15271,N_15041);
nor U18654 (N_18654,N_13939,N_14630);
nand U18655 (N_18655,N_13473,N_15299);
xor U18656 (N_18656,N_15197,N_14045);
nand U18657 (N_18657,N_12904,N_13598);
and U18658 (N_18658,N_13253,N_13748);
xor U18659 (N_18659,N_15105,N_14827);
or U18660 (N_18660,N_13304,N_14335);
nand U18661 (N_18661,N_12910,N_13036);
or U18662 (N_18662,N_13815,N_12916);
and U18663 (N_18663,N_14910,N_12762);
or U18664 (N_18664,N_12558,N_13510);
nor U18665 (N_18665,N_13245,N_15363);
xnor U18666 (N_18666,N_13982,N_12827);
nand U18667 (N_18667,N_13336,N_15163);
nor U18668 (N_18668,N_14714,N_12967);
nor U18669 (N_18669,N_12735,N_13629);
or U18670 (N_18670,N_15227,N_13112);
and U18671 (N_18671,N_13688,N_14875);
nand U18672 (N_18672,N_13025,N_14690);
or U18673 (N_18673,N_13758,N_14188);
xnor U18674 (N_18674,N_14517,N_15290);
nor U18675 (N_18675,N_13006,N_13255);
or U18676 (N_18676,N_14156,N_13420);
nand U18677 (N_18677,N_14600,N_14940);
nor U18678 (N_18678,N_14492,N_14194);
and U18679 (N_18679,N_12795,N_13156);
and U18680 (N_18680,N_14510,N_12969);
nand U18681 (N_18681,N_13220,N_15566);
xor U18682 (N_18682,N_14415,N_15424);
nor U18683 (N_18683,N_12921,N_15166);
nor U18684 (N_18684,N_13137,N_14603);
nor U18685 (N_18685,N_13971,N_15031);
nor U18686 (N_18686,N_13858,N_12549);
and U18687 (N_18687,N_15081,N_12655);
nand U18688 (N_18688,N_13903,N_13913);
and U18689 (N_18689,N_13692,N_15209);
or U18690 (N_18690,N_15018,N_15125);
nor U18691 (N_18691,N_14095,N_13909);
nor U18692 (N_18692,N_13417,N_13485);
and U18693 (N_18693,N_14683,N_12793);
nor U18694 (N_18694,N_13854,N_13016);
nor U18695 (N_18695,N_13521,N_14195);
xnor U18696 (N_18696,N_12708,N_12985);
or U18697 (N_18697,N_14447,N_13222);
nand U18698 (N_18698,N_14771,N_15321);
or U18699 (N_18699,N_15426,N_15566);
xnor U18700 (N_18700,N_13121,N_15165);
or U18701 (N_18701,N_13818,N_15561);
nand U18702 (N_18702,N_14577,N_13841);
xnor U18703 (N_18703,N_14126,N_14985);
and U18704 (N_18704,N_13438,N_14199);
nand U18705 (N_18705,N_13555,N_15140);
xor U18706 (N_18706,N_15214,N_12946);
or U18707 (N_18707,N_13357,N_14386);
and U18708 (N_18708,N_14060,N_14724);
nand U18709 (N_18709,N_12648,N_14645);
and U18710 (N_18710,N_15609,N_13267);
nand U18711 (N_18711,N_14016,N_13740);
or U18712 (N_18712,N_15435,N_13029);
nand U18713 (N_18713,N_13657,N_14022);
nand U18714 (N_18714,N_13135,N_14495);
xor U18715 (N_18715,N_14697,N_13896);
nand U18716 (N_18716,N_14647,N_12932);
nand U18717 (N_18717,N_12600,N_15158);
or U18718 (N_18718,N_12760,N_14207);
and U18719 (N_18719,N_15460,N_12519);
nand U18720 (N_18720,N_14393,N_13885);
and U18721 (N_18721,N_15554,N_14451);
nor U18722 (N_18722,N_14715,N_14061);
and U18723 (N_18723,N_14925,N_14120);
or U18724 (N_18724,N_13092,N_13982);
and U18725 (N_18725,N_14629,N_15449);
nor U18726 (N_18726,N_14075,N_15275);
nand U18727 (N_18727,N_15445,N_15089);
and U18728 (N_18728,N_12611,N_12896);
nor U18729 (N_18729,N_15261,N_14086);
xnor U18730 (N_18730,N_15446,N_12686);
nor U18731 (N_18731,N_13879,N_15355);
nand U18732 (N_18732,N_13171,N_15170);
and U18733 (N_18733,N_13670,N_13476);
and U18734 (N_18734,N_13489,N_12708);
or U18735 (N_18735,N_14270,N_15153);
nand U18736 (N_18736,N_15581,N_12776);
nand U18737 (N_18737,N_14959,N_13745);
nand U18738 (N_18738,N_14677,N_13838);
or U18739 (N_18739,N_14853,N_13957);
xor U18740 (N_18740,N_14271,N_13484);
nand U18741 (N_18741,N_14400,N_14407);
xor U18742 (N_18742,N_15397,N_13052);
or U18743 (N_18743,N_13484,N_15604);
and U18744 (N_18744,N_14656,N_15145);
or U18745 (N_18745,N_12671,N_13027);
xnor U18746 (N_18746,N_12732,N_15610);
or U18747 (N_18747,N_15365,N_14982);
nand U18748 (N_18748,N_15365,N_15062);
and U18749 (N_18749,N_12510,N_14373);
nor U18750 (N_18750,N_15806,N_17527);
or U18751 (N_18751,N_16949,N_18214);
nand U18752 (N_18752,N_18265,N_17442);
nor U18753 (N_18753,N_17202,N_18445);
or U18754 (N_18754,N_16625,N_17818);
and U18755 (N_18755,N_18558,N_18464);
or U18756 (N_18756,N_16697,N_18016);
nand U18757 (N_18757,N_17967,N_16872);
or U18758 (N_18758,N_18099,N_17238);
and U18759 (N_18759,N_18410,N_17324);
and U18760 (N_18760,N_18652,N_16168);
nand U18761 (N_18761,N_16636,N_17595);
nand U18762 (N_18762,N_17380,N_16790);
nand U18763 (N_18763,N_17878,N_16356);
or U18764 (N_18764,N_16808,N_18509);
xor U18765 (N_18765,N_17766,N_16875);
nand U18766 (N_18766,N_17980,N_15952);
nand U18767 (N_18767,N_18457,N_18698);
and U18768 (N_18768,N_16171,N_15734);
nor U18769 (N_18769,N_15626,N_15707);
nand U18770 (N_18770,N_17523,N_15930);
or U18771 (N_18771,N_17187,N_18158);
nor U18772 (N_18772,N_16129,N_18138);
nand U18773 (N_18773,N_16186,N_17506);
nor U18774 (N_18774,N_18363,N_15688);
or U18775 (N_18775,N_16983,N_17641);
or U18776 (N_18776,N_16229,N_16102);
and U18777 (N_18777,N_18080,N_17338);
nor U18778 (N_18778,N_17495,N_15931);
or U18779 (N_18779,N_15703,N_16624);
nand U18780 (N_18780,N_18173,N_16335);
and U18781 (N_18781,N_16459,N_16817);
nand U18782 (N_18782,N_15939,N_18317);
nand U18783 (N_18783,N_18338,N_16578);
nor U18784 (N_18784,N_18068,N_17140);
nor U18785 (N_18785,N_15935,N_16994);
and U18786 (N_18786,N_16517,N_18187);
nand U18787 (N_18787,N_15988,N_16009);
and U18788 (N_18788,N_15959,N_17814);
and U18789 (N_18789,N_17010,N_18682);
nor U18790 (N_18790,N_17018,N_16433);
nand U18791 (N_18791,N_17318,N_15788);
or U18792 (N_18792,N_15743,N_17756);
nor U18793 (N_18793,N_18147,N_15942);
nor U18794 (N_18794,N_18369,N_16680);
or U18795 (N_18795,N_16449,N_18216);
nand U18796 (N_18796,N_15632,N_18401);
xor U18797 (N_18797,N_18153,N_16669);
or U18798 (N_18798,N_17738,N_15675);
nand U18799 (N_18799,N_15728,N_17278);
nor U18800 (N_18800,N_18376,N_17131);
xor U18801 (N_18801,N_16791,N_16737);
and U18802 (N_18802,N_18228,N_17156);
and U18803 (N_18803,N_17886,N_15858);
and U18804 (N_18804,N_17037,N_18600);
or U18805 (N_18805,N_17768,N_16000);
nand U18806 (N_18806,N_16466,N_16405);
xor U18807 (N_18807,N_18518,N_17173);
nand U18808 (N_18808,N_17827,N_18143);
and U18809 (N_18809,N_17868,N_17731);
or U18810 (N_18810,N_16533,N_16868);
xnor U18811 (N_18811,N_17956,N_17463);
and U18812 (N_18812,N_15642,N_17168);
nand U18813 (N_18813,N_18045,N_17762);
nand U18814 (N_18814,N_16141,N_17460);
nor U18815 (N_18815,N_18358,N_17224);
nand U18816 (N_18816,N_18437,N_17352);
and U18817 (N_18817,N_16775,N_15779);
and U18818 (N_18818,N_16842,N_17057);
and U18819 (N_18819,N_16310,N_17340);
nand U18820 (N_18820,N_17082,N_16704);
nand U18821 (N_18821,N_16848,N_18106);
xor U18822 (N_18822,N_18390,N_16504);
or U18823 (N_18823,N_17081,N_16565);
nand U18824 (N_18824,N_18496,N_16178);
or U18825 (N_18825,N_17637,N_17013);
or U18826 (N_18826,N_16959,N_16022);
or U18827 (N_18827,N_16006,N_17543);
and U18828 (N_18828,N_15689,N_15872);
nor U18829 (N_18829,N_18641,N_17353);
or U18830 (N_18830,N_15831,N_17268);
nor U18831 (N_18831,N_16440,N_15915);
nand U18832 (N_18832,N_18744,N_16291);
or U18833 (N_18833,N_17555,N_17551);
or U18834 (N_18834,N_18672,N_16454);
or U18835 (N_18835,N_17369,N_16425);
nand U18836 (N_18836,N_17436,N_18010);
nor U18837 (N_18837,N_17488,N_18283);
xor U18838 (N_18838,N_17773,N_18510);
nor U18839 (N_18839,N_18667,N_16655);
or U18840 (N_18840,N_15681,N_18385);
or U18841 (N_18841,N_18485,N_17217);
nand U18842 (N_18842,N_16258,N_17011);
and U18843 (N_18843,N_16105,N_16410);
or U18844 (N_18844,N_17237,N_17476);
and U18845 (N_18845,N_17409,N_16396);
and U18846 (N_18846,N_17874,N_17405);
nand U18847 (N_18847,N_16308,N_18091);
or U18848 (N_18848,N_16314,N_16931);
and U18849 (N_18849,N_17751,N_18041);
nor U18850 (N_18850,N_15661,N_17284);
nor U18851 (N_18851,N_16593,N_17497);
nor U18852 (N_18852,N_18299,N_17663);
nand U18853 (N_18853,N_17758,N_18566);
or U18854 (N_18854,N_15916,N_17703);
or U18855 (N_18855,N_18629,N_15936);
nor U18856 (N_18856,N_17088,N_18524);
nand U18857 (N_18857,N_17402,N_15949);
or U18858 (N_18858,N_17556,N_16174);
and U18859 (N_18859,N_16820,N_17528);
nand U18860 (N_18860,N_17414,N_17293);
nor U18861 (N_18861,N_16999,N_15932);
nand U18862 (N_18862,N_17176,N_16555);
or U18863 (N_18863,N_17367,N_16892);
and U18864 (N_18864,N_18037,N_16830);
or U18865 (N_18865,N_15889,N_17931);
and U18866 (N_18866,N_17035,N_16123);
and U18867 (N_18867,N_18152,N_18590);
and U18868 (N_18868,N_17817,N_17458);
nor U18869 (N_18869,N_16929,N_17106);
and U18870 (N_18870,N_17295,N_18484);
nor U18871 (N_18871,N_17049,N_16420);
nand U18872 (N_18872,N_18271,N_18375);
xnor U18873 (N_18873,N_18666,N_17845);
and U18874 (N_18874,N_18017,N_18679);
or U18875 (N_18875,N_17784,N_16465);
or U18876 (N_18876,N_18393,N_16547);
or U18877 (N_18877,N_17421,N_15807);
and U18878 (N_18878,N_15818,N_17260);
nand U18879 (N_18879,N_16670,N_16380);
nor U18880 (N_18880,N_16423,N_17892);
nor U18881 (N_18881,N_16696,N_17547);
xnor U18882 (N_18882,N_17794,N_17733);
or U18883 (N_18883,N_18076,N_18710);
or U18884 (N_18884,N_17323,N_15857);
nand U18885 (N_18885,N_16430,N_18335);
nand U18886 (N_18886,N_17039,N_18218);
nor U18887 (N_18887,N_17152,N_15667);
nor U18888 (N_18888,N_17469,N_17916);
xor U18889 (N_18889,N_17507,N_18516);
nor U18890 (N_18890,N_18077,N_17234);
xnor U18891 (N_18891,N_16919,N_18210);
xor U18892 (N_18892,N_16523,N_17672);
nor U18893 (N_18893,N_16400,N_18399);
nand U18894 (N_18894,N_17554,N_18549);
xnor U18895 (N_18895,N_17433,N_16687);
and U18896 (N_18896,N_17658,N_16162);
nor U18897 (N_18897,N_16831,N_17939);
xor U18898 (N_18898,N_17000,N_17838);
nand U18899 (N_18899,N_18193,N_18126);
nor U18900 (N_18900,N_15762,N_18282);
xor U18901 (N_18901,N_18229,N_18243);
nand U18902 (N_18902,N_16752,N_16898);
or U18903 (N_18903,N_17913,N_16712);
nand U18904 (N_18904,N_16458,N_16520);
xor U18905 (N_18905,N_15683,N_18145);
and U18906 (N_18906,N_15691,N_16208);
or U18907 (N_18907,N_17091,N_17689);
nor U18908 (N_18908,N_17264,N_18064);
nor U18909 (N_18909,N_16341,N_16736);
or U18910 (N_18910,N_16126,N_15946);
nand U18911 (N_18911,N_17807,N_18511);
nand U18912 (N_18912,N_17483,N_18149);
nand U18913 (N_18913,N_17508,N_18256);
or U18914 (N_18914,N_16881,N_18148);
or U18915 (N_18915,N_16185,N_16716);
and U18916 (N_18916,N_15981,N_18150);
nand U18917 (N_18917,N_16793,N_17253);
or U18918 (N_18918,N_17372,N_17350);
or U18919 (N_18919,N_16197,N_16560);
and U18920 (N_18920,N_17148,N_17963);
and U18921 (N_18921,N_18088,N_17200);
and U18922 (N_18922,N_16726,N_17023);
and U18923 (N_18923,N_18571,N_15659);
nor U18924 (N_18924,N_16118,N_17851);
or U18925 (N_18925,N_17137,N_16821);
nor U18926 (N_18926,N_17865,N_17744);
nand U18927 (N_18927,N_16815,N_15989);
or U18928 (N_18928,N_17654,N_17928);
xor U18929 (N_18929,N_17968,N_18285);
nand U18930 (N_18930,N_16001,N_16557);
xnor U18931 (N_18931,N_18535,N_16537);
nand U18932 (N_18932,N_17438,N_18441);
nand U18933 (N_18933,N_16602,N_17855);
xor U18934 (N_18934,N_18300,N_17684);
or U18935 (N_18935,N_16033,N_17456);
and U18936 (N_18936,N_15972,N_18318);
and U18937 (N_18937,N_17999,N_18550);
xor U18938 (N_18938,N_16135,N_18264);
and U18939 (N_18939,N_18092,N_17019);
nand U18940 (N_18940,N_16407,N_16684);
and U18941 (N_18941,N_16442,N_16045);
or U18942 (N_18942,N_16613,N_18562);
nand U18943 (N_18943,N_16061,N_18542);
nor U18944 (N_18944,N_16021,N_17686);
and U18945 (N_18945,N_16605,N_18072);
nor U18946 (N_18946,N_16637,N_16414);
nor U18947 (N_18947,N_16247,N_17885);
and U18948 (N_18948,N_16481,N_16763);
and U18949 (N_18949,N_18279,N_15750);
and U18950 (N_18950,N_17782,N_16594);
nor U18951 (N_18951,N_15833,N_15870);
or U18952 (N_18952,N_16090,N_18043);
or U18953 (N_18953,N_15726,N_17820);
nor U18954 (N_18954,N_15684,N_16411);
nand U18955 (N_18955,N_17761,N_17186);
nand U18956 (N_18956,N_17804,N_18601);
nor U18957 (N_18957,N_18732,N_16603);
nor U18958 (N_18958,N_18697,N_16128);
and U18959 (N_18959,N_16453,N_18493);
nor U18960 (N_18960,N_17661,N_17989);
and U18961 (N_18961,N_16974,N_18684);
xnor U18962 (N_18962,N_16635,N_17447);
or U18963 (N_18963,N_18035,N_16644);
and U18964 (N_18964,N_17429,N_17104);
or U18965 (N_18965,N_16780,N_16270);
nor U18966 (N_18966,N_17065,N_18012);
or U18967 (N_18967,N_18166,N_17645);
nor U18968 (N_18968,N_17102,N_15682);
or U18969 (N_18969,N_15874,N_17258);
or U18970 (N_18970,N_15754,N_18458);
or U18971 (N_18971,N_17073,N_17946);
or U18972 (N_18972,N_18651,N_17009);
nor U18973 (N_18973,N_18224,N_18028);
or U18974 (N_18974,N_18361,N_15893);
nor U18975 (N_18975,N_16119,N_17164);
and U18976 (N_18976,N_17249,N_17671);
and U18977 (N_18977,N_18638,N_18523);
nor U18978 (N_18978,N_18132,N_16525);
nor U18979 (N_18979,N_16403,N_18545);
nand U18980 (N_18980,N_17191,N_17604);
nor U18981 (N_18981,N_18066,N_15848);
and U18982 (N_18982,N_18630,N_15881);
xor U18983 (N_18983,N_15634,N_18097);
or U18984 (N_18984,N_18482,N_15655);
nor U18985 (N_18985,N_17045,N_15644);
or U18986 (N_18986,N_16997,N_16721);
or U18987 (N_18987,N_17113,N_16012);
nand U18988 (N_18988,N_17064,N_18622);
and U18989 (N_18989,N_15671,N_18257);
nor U18990 (N_18990,N_16506,N_15747);
and U18991 (N_18991,N_18724,N_15637);
and U18992 (N_18992,N_17674,N_18422);
or U18993 (N_18993,N_18705,N_15853);
and U18994 (N_18994,N_15756,N_17247);
nand U18995 (N_18995,N_17815,N_16031);
or U18996 (N_18996,N_16535,N_16695);
or U18997 (N_18997,N_17917,N_18522);
and U18998 (N_18998,N_17386,N_17289);
and U18999 (N_18999,N_17403,N_17695);
or U19000 (N_19000,N_16779,N_16811);
or U19001 (N_19001,N_17477,N_16032);
or U19002 (N_19002,N_17841,N_17283);
and U19003 (N_19003,N_18397,N_16645);
and U19004 (N_19004,N_15776,N_17316);
nand U19005 (N_19005,N_18414,N_16773);
and U19006 (N_19006,N_18134,N_17683);
nand U19007 (N_19007,N_18480,N_17530);
and U19008 (N_19008,N_17538,N_17453);
nor U19009 (N_19009,N_16915,N_15654);
xor U19010 (N_19010,N_18115,N_16389);
and U19011 (N_19011,N_18525,N_18573);
and U19012 (N_19012,N_18089,N_15713);
xnor U19013 (N_19013,N_18661,N_15860);
nor U19014 (N_19014,N_17440,N_17591);
and U19015 (N_19015,N_17521,N_16142);
nor U19016 (N_19016,N_16127,N_17629);
nand U19017 (N_19017,N_17005,N_18624);
or U19018 (N_19018,N_16391,N_18577);
and U19019 (N_19019,N_18146,N_16293);
nor U19020 (N_19020,N_17948,N_18121);
or U19021 (N_19021,N_16026,N_18316);
and U19022 (N_19022,N_16798,N_16933);
nand U19023 (N_19023,N_18640,N_16436);
nor U19024 (N_19024,N_18122,N_16249);
xnor U19025 (N_19025,N_17618,N_16275);
nand U19026 (N_19026,N_16214,N_15794);
nand U19027 (N_19027,N_18280,N_18548);
nand U19028 (N_19028,N_15879,N_17145);
nand U19029 (N_19029,N_16524,N_16179);
nand U19030 (N_19030,N_16671,N_17896);
nand U19031 (N_19031,N_17667,N_18212);
nor U19032 (N_19032,N_18686,N_18704);
nand U19033 (N_19033,N_17408,N_18718);
xnor U19034 (N_19034,N_18230,N_17639);
or U19035 (N_19035,N_16538,N_17617);
nor U19036 (N_19036,N_17267,N_18534);
nand U19037 (N_19037,N_17589,N_16078);
nand U19038 (N_19038,N_18673,N_17392);
and U19039 (N_19039,N_16516,N_16722);
or U19040 (N_19040,N_16053,N_16058);
or U19041 (N_19041,N_16782,N_16110);
and U19042 (N_19042,N_17767,N_16512);
nand U19043 (N_19043,N_18253,N_15954);
and U19044 (N_19044,N_17001,N_17986);
nor U19045 (N_19045,N_17536,N_17864);
nor U19046 (N_19046,N_17741,N_15826);
nand U19047 (N_19047,N_16976,N_18060);
nor U19048 (N_19048,N_16859,N_18308);
nor U19049 (N_19049,N_17351,N_18565);
and U19050 (N_19050,N_17459,N_18270);
or U19051 (N_19051,N_15679,N_18483);
nor U19052 (N_19052,N_16357,N_17752);
nand U19053 (N_19053,N_17008,N_17016);
xor U19054 (N_19054,N_18498,N_17549);
or U19055 (N_19055,N_17921,N_16870);
or U19056 (N_19056,N_16472,N_17379);
xnor U19057 (N_19057,N_17336,N_17632);
or U19058 (N_19058,N_15962,N_17903);
or U19059 (N_19059,N_16418,N_16024);
or U19060 (N_19060,N_17895,N_17525);
and U19061 (N_19061,N_16665,N_17877);
or U19062 (N_19062,N_18274,N_18465);
and U19063 (N_19063,N_18082,N_18726);
and U19064 (N_19064,N_17537,N_15757);
and U19065 (N_19065,N_17753,N_16551);
nor U19066 (N_19066,N_16928,N_16324);
nand U19067 (N_19067,N_18249,N_18079);
nand U19068 (N_19068,N_18350,N_17711);
xnor U19069 (N_19069,N_18026,N_16794);
or U19070 (N_19070,N_15649,N_16920);
nand U19071 (N_19071,N_17032,N_18327);
and U19072 (N_19072,N_18286,N_18426);
or U19073 (N_19073,N_17613,N_17736);
and U19074 (N_19074,N_15639,N_18107);
and U19075 (N_19075,N_18380,N_17074);
or U19076 (N_19076,N_16772,N_16011);
nor U19077 (N_19077,N_16264,N_16166);
xnor U19078 (N_19078,N_17501,N_17155);
and U19079 (N_19079,N_17432,N_18367);
nor U19080 (N_19080,N_17068,N_18038);
nand U19081 (N_19081,N_18747,N_17242);
or U19082 (N_19082,N_18086,N_17116);
nor U19083 (N_19083,N_15862,N_16529);
and U19084 (N_19084,N_17211,N_15797);
nor U19085 (N_19085,N_16686,N_16239);
and U19086 (N_19086,N_15668,N_17244);
xor U19087 (N_19087,N_17180,N_17715);
and U19088 (N_19088,N_16640,N_16307);
nor U19089 (N_19089,N_17038,N_15868);
or U19090 (N_19090,N_16689,N_17254);
nand U19091 (N_19091,N_18746,N_18033);
or U19092 (N_19092,N_15838,N_18074);
nand U19093 (N_19093,N_16132,N_16664);
or U19094 (N_19094,N_18120,N_16663);
xnor U19095 (N_19095,N_16942,N_16151);
nor U19096 (N_19096,N_16413,N_17167);
nand U19097 (N_19097,N_17227,N_18172);
nand U19098 (N_19098,N_15852,N_17014);
nand U19099 (N_19099,N_18137,N_16246);
nand U19100 (N_19100,N_17363,N_17884);
nand U19101 (N_19101,N_16500,N_18749);
nand U19102 (N_19102,N_16130,N_17110);
nand U19103 (N_19103,N_18075,N_17232);
nand U19104 (N_19104,N_17089,N_16395);
xor U19105 (N_19105,N_16445,N_16518);
and U19106 (N_19106,N_18443,N_18289);
or U19107 (N_19107,N_18103,N_15929);
or U19108 (N_19108,N_18181,N_17566);
or U19109 (N_19109,N_18586,N_16702);
or U19110 (N_19110,N_16960,N_17216);
nor U19111 (N_19111,N_17976,N_18151);
nor U19112 (N_19112,N_17856,N_16956);
and U19113 (N_19113,N_17823,N_16294);
nor U19114 (N_19114,N_18027,N_16330);
nand U19115 (N_19115,N_17171,N_16879);
or U19116 (N_19116,N_18139,N_18301);
nand U19117 (N_19117,N_16302,N_16786);
or U19118 (N_19118,N_15774,N_16167);
or U19119 (N_19119,N_17912,N_17564);
nor U19120 (N_19120,N_15687,N_17748);
nand U19121 (N_19121,N_17170,N_18555);
nor U19122 (N_19122,N_15796,N_18052);
nor U19123 (N_19123,N_18078,N_16853);
nor U19124 (N_19124,N_16276,N_18462);
nor U19125 (N_19125,N_16987,N_15998);
and U19126 (N_19126,N_16550,N_16117);
nor U19127 (N_19127,N_18637,N_18556);
nor U19128 (N_19128,N_16804,N_16585);
nor U19129 (N_19129,N_16460,N_17286);
or U19130 (N_19130,N_16354,N_18610);
and U19131 (N_19131,N_18105,N_16347);
and U19132 (N_19132,N_16572,N_17947);
nor U19133 (N_19133,N_17522,N_16486);
and U19134 (N_19134,N_16498,N_15913);
or U19135 (N_19135,N_17612,N_15628);
nand U19136 (N_19136,N_17498,N_17520);
nand U19137 (N_19137,N_17754,N_15867);
and U19138 (N_19138,N_17450,N_16975);
or U19139 (N_19139,N_17359,N_16713);
or U19140 (N_19140,N_15710,N_18501);
nor U19141 (N_19141,N_15745,N_16296);
nand U19142 (N_19142,N_17151,N_18567);
or U19143 (N_19143,N_18602,N_17687);
and U19144 (N_19144,N_15740,N_17777);
xnor U19145 (N_19145,N_16406,N_16220);
and U19146 (N_19146,N_16703,N_17077);
and U19147 (N_19147,N_15702,N_15662);
and U19148 (N_19148,N_16388,N_18683);
or U19149 (N_19149,N_17586,N_17346);
nand U19150 (N_19150,N_17643,N_18715);
or U19151 (N_19151,N_18128,N_15795);
or U19152 (N_19152,N_15813,N_16649);
and U19153 (N_19153,N_15992,N_17378);
nand U19154 (N_19154,N_16828,N_15714);
nand U19155 (N_19155,N_17942,N_17337);
or U19156 (N_19156,N_18712,N_16352);
or U19157 (N_19157,N_18323,N_17142);
or U19158 (N_19158,N_15815,N_18305);
nor U19159 (N_19159,N_16200,N_17581);
or U19160 (N_19160,N_15722,N_16175);
and U19161 (N_19161,N_16378,N_16043);
or U19162 (N_19162,N_16741,N_17759);
or U19163 (N_19163,N_18728,N_17825);
nor U19164 (N_19164,N_18112,N_16944);
or U19165 (N_19165,N_15777,N_15887);
and U19166 (N_19166,N_15937,N_16172);
nor U19167 (N_19167,N_16143,N_18000);
nand U19168 (N_19168,N_17991,N_16195);
nand U19169 (N_19169,N_16943,N_17198);
nand U19170 (N_19170,N_18260,N_16646);
nor U19171 (N_19171,N_16099,N_17702);
or U19172 (N_19172,N_18540,N_18477);
nor U19173 (N_19173,N_16424,N_17422);
or U19174 (N_19174,N_17276,N_17446);
or U19175 (N_19175,N_16060,N_18636);
or U19176 (N_19176,N_16568,N_18722);
xnor U19177 (N_19177,N_16158,N_17412);
nand U19178 (N_19178,N_17382,N_17621);
nor U19179 (N_19179,N_18584,N_17925);
and U19180 (N_19180,N_16934,N_17983);
or U19181 (N_19181,N_17919,N_17785);
nand U19182 (N_19182,N_16202,N_17241);
nand U19183 (N_19183,N_18180,N_17568);
nor U19184 (N_19184,N_17574,N_17914);
nor U19185 (N_19185,N_18681,N_16274);
and U19186 (N_19186,N_17548,N_17389);
or U19187 (N_19187,N_16316,N_18160);
xor U19188 (N_19188,N_16470,N_18095);
or U19189 (N_19189,N_17630,N_15666);
nand U19190 (N_19190,N_16029,N_18634);
nor U19191 (N_19191,N_18188,N_17275);
nor U19192 (N_19192,N_18529,N_16865);
nor U19193 (N_19193,N_17926,N_15803);
and U19194 (N_19194,N_18170,N_15938);
xor U19195 (N_19195,N_18284,N_15866);
xnor U19196 (N_19196,N_15643,N_16211);
nand U19197 (N_19197,N_16907,N_16768);
or U19198 (N_19198,N_17087,N_16957);
nor U19199 (N_19199,N_17271,N_17584);
or U19200 (N_19200,N_17854,N_17857);
or U19201 (N_19201,N_18433,N_18592);
nor U19202 (N_19202,N_18278,N_18474);
nand U19203 (N_19203,N_15625,N_16309);
nor U19204 (N_19204,N_18406,N_17471);
or U19205 (N_19205,N_15890,N_17840);
and U19206 (N_19206,N_17210,N_16760);
and U19207 (N_19207,N_17570,N_16761);
and U19208 (N_19208,N_18475,N_16441);
nand U19209 (N_19209,N_15835,N_17132);
and U19210 (N_19210,N_18298,N_18687);
nand U19211 (N_19211,N_16322,N_18472);
nor U19212 (N_19212,N_15841,N_17890);
nor U19213 (N_19213,N_16085,N_17821);
nor U19214 (N_19214,N_16873,N_16511);
nor U19215 (N_19215,N_16776,N_18674);
xor U19216 (N_19216,N_15911,N_18677);
nor U19217 (N_19217,N_18449,N_17796);
nand U19218 (N_19218,N_16416,N_15708);
and U19219 (N_19219,N_15819,N_17331);
nand U19220 (N_19220,N_16724,N_16124);
nand U19221 (N_19221,N_18310,N_16361);
nor U19222 (N_19222,N_16279,N_16733);
xor U19223 (N_19223,N_17114,N_17345);
nand U19224 (N_19224,N_15814,N_16586);
and U19225 (N_19225,N_17594,N_18135);
and U19226 (N_19226,N_17682,N_17431);
nor U19227 (N_19227,N_17755,N_17256);
or U19228 (N_19228,N_16607,N_18597);
or U19229 (N_19229,N_17069,N_17099);
nor U19230 (N_19230,N_18574,N_18381);
or U19231 (N_19231,N_18727,N_16940);
and U19232 (N_19232,N_15995,N_17847);
nor U19233 (N_19233,N_16251,N_18307);
nor U19234 (N_19234,N_16982,N_16094);
nand U19235 (N_19235,N_16451,N_16005);
xor U19236 (N_19236,N_18500,N_16614);
or U19237 (N_19237,N_17084,N_17050);
and U19238 (N_19238,N_16355,N_17747);
or U19239 (N_19239,N_18093,N_18531);
nand U19240 (N_19240,N_18288,N_15696);
nor U19241 (N_19241,N_15771,N_16953);
and U19242 (N_19242,N_17529,N_17317);
and U19243 (N_19243,N_17396,N_15948);
xor U19244 (N_19244,N_16503,N_17326);
xnor U19245 (N_19245,N_16834,N_17296);
or U19246 (N_19246,N_17079,N_16332);
nor U19247 (N_19247,N_17954,N_16877);
xnor U19248 (N_19248,N_18039,N_17822);
nor U19249 (N_19249,N_16754,N_16850);
xor U19250 (N_19250,N_17012,N_16969);
or U19251 (N_19251,N_18100,N_16041);
or U19252 (N_19252,N_16304,N_16985);
and U19253 (N_19253,N_17519,N_17924);
nor U19254 (N_19254,N_17031,N_18290);
and U19255 (N_19255,N_17328,N_18312);
and U19256 (N_19256,N_17676,N_18502);
xnor U19257 (N_19257,N_16845,N_16660);
or U19258 (N_19258,N_17552,N_16629);
xnor U19259 (N_19259,N_17560,N_16209);
nand U19260 (N_19260,N_17384,N_17499);
nor U19261 (N_19261,N_16269,N_17615);
xor U19262 (N_19262,N_16924,N_18136);
or U19263 (N_19263,N_18415,N_16710);
and U19264 (N_19264,N_17370,N_16528);
or U19265 (N_19265,N_16014,N_16244);
nand U19266 (N_19266,N_17935,N_18258);
nand U19267 (N_19267,N_18678,N_17231);
xor U19268 (N_19268,N_17932,N_15720);
nor U19269 (N_19269,N_18067,N_17699);
nand U19270 (N_19270,N_16415,N_18463);
or U19271 (N_19271,N_18133,N_18319);
nor U19272 (N_19272,N_15731,N_16180);
or U19273 (N_19273,N_16764,N_16945);
or U19274 (N_19274,N_17022,N_17514);
nor U19275 (N_19275,N_18104,N_18362);
and U19276 (N_19276,N_17897,N_16905);
nand U19277 (N_19277,N_18167,N_16038);
nor U19278 (N_19278,N_18202,N_16390);
nand U19279 (N_19279,N_16428,N_15715);
and U19280 (N_19280,N_17559,N_17418);
and U19281 (N_19281,N_18733,N_16885);
or U19282 (N_19282,N_16328,N_17026);
nand U19283 (N_19283,N_16719,N_15724);
xor U19284 (N_19284,N_17648,N_18398);
nand U19285 (N_19285,N_17098,N_17881);
or U19286 (N_19286,N_17698,N_17420);
nand U19287 (N_19287,N_16243,N_16505);
nor U19288 (N_19288,N_16963,N_18419);
and U19289 (N_19289,N_15646,N_18175);
or U19290 (N_19290,N_17642,N_17719);
and U19291 (N_19291,N_17354,N_18619);
or U19292 (N_19292,N_17563,N_16984);
or U19293 (N_19293,N_18714,N_18025);
and U19294 (N_19294,N_17233,N_17934);
or U19295 (N_19295,N_17920,N_15997);
nand U19296 (N_19296,N_18685,N_17750);
and U19297 (N_19297,N_18015,N_16232);
xnor U19298 (N_19298,N_15749,N_18246);
and U19299 (N_19299,N_16096,N_16490);
or U19300 (N_19300,N_18425,N_17266);
nand U19301 (N_19301,N_17071,N_17330);
or U19302 (N_19302,N_17117,N_15744);
nand U19303 (N_19303,N_15760,N_16444);
and U19304 (N_19304,N_15837,N_15905);
and U19305 (N_19305,N_16371,N_16133);
nand U19306 (N_19306,N_17813,N_16751);
nand U19307 (N_19307,N_18250,N_17201);
or U19308 (N_19308,N_17334,N_16806);
or U19309 (N_19309,N_16131,N_16965);
nor U19310 (N_19310,N_18005,N_18528);
and U19311 (N_19311,N_15775,N_17974);
and U19312 (N_19312,N_16604,N_17806);
and U19313 (N_19313,N_17115,N_16954);
nand U19314 (N_19314,N_18455,N_17627);
nand U19315 (N_19315,N_15694,N_16338);
or U19316 (N_19316,N_17927,N_17837);
nor U19317 (N_19317,N_18623,N_17704);
nand U19318 (N_19318,N_18073,N_16497);
nor U19319 (N_19319,N_18254,N_17995);
nor U19320 (N_19320,N_18032,N_17473);
or U19321 (N_19321,N_16077,N_16679);
and U19322 (N_19322,N_17192,N_18626);
nand U19323 (N_19323,N_17670,N_16417);
nand U19324 (N_19324,N_18314,N_17047);
and U19325 (N_19325,N_16223,N_16619);
and U19326 (N_19326,N_18668,N_17871);
and U19327 (N_19327,N_16315,N_17491);
or U19328 (N_19328,N_17622,N_16588);
and U19329 (N_19329,N_16950,N_16295);
and U19330 (N_19330,N_18297,N_16730);
nand U19331 (N_19331,N_16777,N_17726);
nor U19332 (N_19332,N_16469,N_15907);
and U19333 (N_19333,N_18371,N_16502);
or U19334 (N_19334,N_17341,N_17571);
and U19335 (N_19335,N_16088,N_17938);
and U19336 (N_19336,N_16292,N_16977);
nor U19337 (N_19337,N_17130,N_15908);
and U19338 (N_19338,N_17395,N_15996);
xnor U19339 (N_19339,N_17580,N_17636);
nor U19340 (N_19340,N_16735,N_18551);
or U19341 (N_19341,N_16176,N_16321);
nand U19342 (N_19342,N_15823,N_16610);
nand U19343 (N_19343,N_18085,N_18084);
or U19344 (N_19344,N_15653,N_15676);
nor U19345 (N_19345,N_16228,N_16788);
nor U19346 (N_19346,N_16008,N_17787);
and U19347 (N_19347,N_16313,N_16583);
and U19348 (N_19348,N_15822,N_18315);
xor U19349 (N_19349,N_16899,N_17312);
and U19350 (N_19350,N_16918,N_15910);
nand U19351 (N_19351,N_17600,N_17902);
and U19352 (N_19352,N_18536,N_16025);
nand U19353 (N_19353,N_16037,N_16651);
nor U19354 (N_19354,N_18198,N_17859);
or U19355 (N_19355,N_16320,N_17095);
or U19356 (N_19356,N_16596,N_16711);
nand U19357 (N_19357,N_17561,N_18178);
xor U19358 (N_19358,N_15902,N_17608);
xnor U19359 (N_19359,N_17664,N_15864);
or U19360 (N_19360,N_18349,N_18707);
xor U19361 (N_19361,N_17185,N_15759);
xnor U19362 (N_19362,N_18447,N_18235);
nor U19363 (N_19363,N_18333,N_16926);
nor U19364 (N_19364,N_18420,N_16838);
or U19365 (N_19365,N_15909,N_16082);
or U19366 (N_19366,N_18580,N_16206);
xnor U19367 (N_19367,N_15976,N_16964);
or U19368 (N_19368,N_15993,N_16911);
and U19369 (N_19369,N_16962,N_16622);
or U19370 (N_19370,N_18430,N_16521);
nor U19371 (N_19371,N_15658,N_16839);
and U19372 (N_19372,N_15629,N_17329);
xor U19373 (N_19373,N_16204,N_16611);
nor U19374 (N_19374,N_18609,N_16348);
or U19375 (N_19375,N_15842,N_16946);
and U19376 (N_19376,N_16349,N_16137);
xnor U19377 (N_19377,N_16690,N_16157);
and U19378 (N_19378,N_18311,N_16114);
or U19379 (N_19379,N_16374,N_15674);
nor U19380 (N_19380,N_17846,N_18461);
nand U19381 (N_19381,N_18209,N_15631);
nand U19382 (N_19382,N_17588,N_17111);
or U19383 (N_19383,N_18199,N_17996);
nor U19384 (N_19384,N_17665,N_16219);
nor U19385 (N_19385,N_17517,N_18589);
xor U19386 (N_19386,N_15884,N_18019);
nand U19387 (N_19387,N_15914,N_16067);
xnor U19388 (N_19388,N_15650,N_17393);
or U19389 (N_19389,N_16844,N_15763);
nand U19390 (N_19390,N_16991,N_16851);
nand U19391 (N_19391,N_15920,N_17940);
and U19392 (N_19392,N_15978,N_17869);
nand U19393 (N_19393,N_16958,N_18632);
or U19394 (N_19394,N_16213,N_15966);
and U19395 (N_19395,N_17076,N_18388);
or U19396 (N_19396,N_18294,N_17647);
and U19397 (N_19397,N_18486,N_16615);
nand U19398 (N_19398,N_16729,N_17335);
nand U19399 (N_19399,N_16863,N_17486);
nor U19400 (N_19400,N_15651,N_18645);
or U19401 (N_19401,N_18723,N_16961);
nor U19402 (N_19402,N_18649,N_16173);
nor U19403 (N_19403,N_17223,N_17121);
nand U19404 (N_19404,N_18669,N_17062);
nand U19405 (N_19405,N_17655,N_16421);
nor U19406 (N_19406,N_18644,N_17366);
nor U19407 (N_19407,N_17998,N_17634);
nand U19408 (N_19408,N_17831,N_18125);
and U19409 (N_19409,N_15851,N_18647);
xor U19410 (N_19410,N_17789,N_16807);
or U19411 (N_19411,N_18538,N_18676);
or U19412 (N_19412,N_16570,N_17259);
nand U19413 (N_19413,N_16020,N_18409);
nand U19414 (N_19414,N_16039,N_18639);
and U19415 (N_19415,N_18141,N_18739);
or U19416 (N_19416,N_16177,N_16508);
nor U19417 (N_19417,N_18227,N_16641);
and U19418 (N_19418,N_18309,N_18047);
nand U19419 (N_19419,N_16862,N_16404);
nor U19420 (N_19420,N_16034,N_16160);
nand U19421 (N_19421,N_16080,N_17729);
nand U19422 (N_19422,N_18023,N_16193);
nand U19423 (N_19423,N_16682,N_15969);
or U19424 (N_19424,N_17860,N_16948);
or U19425 (N_19425,N_17322,N_16734);
or U19426 (N_19426,N_17593,N_18098);
or U19427 (N_19427,N_16639,N_15891);
nor U19428 (N_19428,N_18671,N_17475);
xor U19429 (N_19429,N_17515,N_16280);
nand U19430 (N_19430,N_17066,N_15956);
nand U19431 (N_19431,N_17652,N_17020);
nor U19432 (N_19432,N_17848,N_17572);
nand U19433 (N_19433,N_15832,N_16448);
nor U19434 (N_19434,N_17027,N_16819);
xor U19435 (N_19435,N_17090,N_17470);
nor U19436 (N_19436,N_17085,N_16483);
nand U19437 (N_19437,N_17697,N_17882);
nand U19438 (N_19438,N_16579,N_16097);
nor U19439 (N_19439,N_16561,N_18276);
and U19440 (N_19440,N_17302,N_15982);
nor U19441 (N_19441,N_15843,N_15958);
nor U19442 (N_19442,N_16473,N_15699);
nor U19443 (N_19443,N_16678,N_17133);
nor U19444 (N_19444,N_15999,N_18204);
xnor U19445 (N_19445,N_17828,N_17122);
nand U19446 (N_19446,N_17861,N_16706);
nor U19447 (N_19447,N_16801,N_18040);
and U19448 (N_19448,N_18508,N_18417);
or U19449 (N_19449,N_17710,N_16476);
nand U19450 (N_19450,N_16215,N_15711);
and U19451 (N_19451,N_18690,N_18743);
nand U19452 (N_19452,N_15965,N_15940);
nand U19453 (N_19453,N_16259,N_15753);
and U19454 (N_19454,N_18206,N_18203);
nor U19455 (N_19455,N_16050,N_17592);
and U19456 (N_19456,N_18142,N_18403);
xor U19457 (N_19457,N_17274,N_17108);
nand U19458 (N_19458,N_17222,N_16181);
and U19459 (N_19459,N_18337,N_18051);
and U19460 (N_19460,N_15855,N_18659);
nand U19461 (N_19461,N_16903,N_17096);
nor U19462 (N_19462,N_17725,N_17616);
or U19463 (N_19463,N_17377,N_15809);
and U19464 (N_19464,N_16238,N_15820);
nand U19465 (N_19465,N_15704,N_17272);
xor U19466 (N_19466,N_17355,N_17793);
nor U19467 (N_19467,N_16795,N_18334);
or U19468 (N_19468,N_18277,N_17732);
xnor U19469 (N_19469,N_16036,N_17006);
or U19470 (N_19470,N_18665,N_17512);
xnor U19471 (N_19471,N_18488,N_17836);
and U19472 (N_19472,N_16252,N_16890);
xnor U19473 (N_19473,N_17808,N_17763);
nor U19474 (N_19474,N_15840,N_16013);
or U19475 (N_19475,N_18438,N_16104);
nor U19476 (N_19476,N_18348,N_18706);
xor U19477 (N_19477,N_16519,N_17657);
and U19478 (N_19478,N_16283,N_17199);
nor U19479 (N_19479,N_18194,N_16951);
or U19480 (N_19480,N_17282,N_15638);
or U19481 (N_19481,N_16113,N_16569);
nand U19482 (N_19482,N_16471,N_17472);
or U19483 (N_19483,N_17614,N_17553);
xor U19484 (N_19484,N_16363,N_16393);
or U19485 (N_19485,N_16156,N_17757);
or U19486 (N_19486,N_18177,N_18386);
or U19487 (N_19487,N_18207,N_16125);
or U19488 (N_19488,N_16886,N_15793);
and U19489 (N_19489,N_16370,N_16002);
or U19490 (N_19490,N_17043,N_15786);
nand U19491 (N_19491,N_15636,N_15630);
and U19492 (N_19492,N_17666,N_18418);
xor U19493 (N_19493,N_16255,N_18526);
nor U19494 (N_19494,N_18110,N_17800);
and U19495 (N_19495,N_17333,N_17981);
and U19496 (N_19496,N_18576,N_17017);
nor U19497 (N_19497,N_18658,N_17364);
and U19498 (N_19498,N_17791,N_17205);
nor U19499 (N_19499,N_16358,N_18063);
nand U19500 (N_19500,N_17659,N_17292);
and U19501 (N_19501,N_18351,N_16144);
nand U19502 (N_19502,N_16727,N_16513);
or U19503 (N_19503,N_16564,N_16802);
or U19504 (N_19504,N_17374,N_17494);
nand U19505 (N_19505,N_15971,N_15784);
nand U19506 (N_19506,N_16643,N_16748);
or U19507 (N_19507,N_16774,N_16783);
or U19508 (N_19508,N_17716,N_18553);
xnor U19509 (N_19509,N_18313,N_15769);
and U19510 (N_19510,N_18220,N_16633);
and U19511 (N_19511,N_18579,N_18400);
nand U19512 (N_19512,N_16066,N_15967);
nand U19513 (N_19513,N_15925,N_18635);
nand U19514 (N_19514,N_17305,N_16120);
or U19515 (N_19515,N_16496,N_16311);
nor U19516 (N_19516,N_18268,N_15716);
nor U19517 (N_19517,N_15861,N_16480);
nor U19518 (N_19518,N_18740,N_15712);
nand U19519 (N_19519,N_18675,N_17609);
xnor U19520 (N_19520,N_18691,N_16545);
nor U19521 (N_19521,N_17417,N_17123);
xnor U19522 (N_19522,N_18164,N_18021);
or U19523 (N_19523,N_17906,N_15673);
nand U19524 (N_19524,N_16089,N_16281);
nor U19525 (N_19525,N_17953,N_15847);
nand U19526 (N_19526,N_15945,N_16688);
nand U19527 (N_19527,N_16343,N_17416);
nand U19528 (N_19528,N_15751,N_17631);
or U19529 (N_19529,N_17742,N_16621);
and U19530 (N_19530,N_16284,N_18321);
nand U19531 (N_19531,N_16152,N_17182);
xnor U19532 (N_19532,N_17597,N_16477);
nor U19533 (N_19533,N_16289,N_15839);
nand U19534 (N_19534,N_18185,N_15859);
xor U19535 (N_19535,N_17810,N_17034);
xor U19536 (N_19536,N_16326,N_16450);
nand U19537 (N_19537,N_18382,N_17582);
or U19538 (N_19538,N_16910,N_16253);
and U19539 (N_19539,N_17692,N_17315);
xor U19540 (N_19540,N_16359,N_18598);
and U19541 (N_19541,N_17679,N_16825);
nand U19542 (N_19542,N_16134,N_18293);
nor U19543 (N_19543,N_16499,N_16582);
and U19544 (N_19544,N_16256,N_15836);
or U19545 (N_19545,N_15770,N_17172);
and U19546 (N_19546,N_17531,N_16234);
or U19547 (N_19547,N_17261,N_18694);
nand U19548 (N_19548,N_16035,N_17730);
nand U19549 (N_19549,N_17401,N_16849);
and U19550 (N_19550,N_16803,N_16662);
nand U19551 (N_19551,N_18476,N_17721);
nand U19552 (N_19552,N_18320,N_17835);
and U19553 (N_19553,N_16809,N_16386);
nor U19554 (N_19554,N_16248,N_15799);
or U19555 (N_19555,N_15941,N_18604);
or U19556 (N_19556,N_16201,N_16447);
xor U19557 (N_19557,N_16589,N_15698);
or U19558 (N_19558,N_15727,N_17889);
nand U19559 (N_19559,N_18183,N_17194);
nand U19560 (N_19560,N_16191,N_16571);
nor U19561 (N_19561,N_17025,N_16146);
nand U19562 (N_19562,N_17562,N_18621);
nor U19563 (N_19563,N_16306,N_18266);
or U19564 (N_19564,N_16884,N_18007);
or U19565 (N_19565,N_18693,N_17576);
or U19566 (N_19566,N_17739,N_16789);
and U19567 (N_19567,N_18241,N_17228);
and U19568 (N_19568,N_15964,N_16676);
or U19569 (N_19569,N_15878,N_15693);
nand U19570 (N_19570,N_16981,N_17285);
and U19571 (N_19571,N_17072,N_18328);
nand U19572 (N_19572,N_16548,N_17143);
nand U19573 (N_19573,N_16541,N_17805);
and U19574 (N_19574,N_17373,N_18717);
or U19575 (N_19575,N_16377,N_17709);
and U19576 (N_19576,N_17966,N_15787);
or U19577 (N_19577,N_18154,N_16079);
and U19578 (N_19578,N_17635,N_15686);
and U19579 (N_19579,N_17399,N_17147);
and U19580 (N_19580,N_18618,N_17504);
nand U19581 (N_19581,N_17467,N_15718);
and U19582 (N_19582,N_17834,N_15994);
and U19583 (N_19583,N_16340,N_18346);
nor U19584 (N_19584,N_16916,N_17993);
or U19585 (N_19585,N_18720,N_18189);
nand U19586 (N_19586,N_16685,N_17875);
and U19587 (N_19587,N_18247,N_18520);
nand U19588 (N_19588,N_16861,N_18096);
nor U19589 (N_19589,N_17959,N_18130);
and U19590 (N_19590,N_17304,N_16154);
or U19591 (N_19591,N_15974,N_17381);
nand U19592 (N_19592,N_18664,N_16921);
and U19593 (N_19593,N_18552,N_16573);
xnor U19594 (N_19594,N_16367,N_18239);
and U19595 (N_19595,N_17650,N_17795);
xnor U19596 (N_19596,N_16303,N_17735);
and U19597 (N_19597,N_17545,N_17424);
xnor U19598 (N_19598,N_18054,N_18109);
nand U19599 (N_19599,N_17883,N_17368);
nand U19600 (N_19600,N_17585,N_16205);
nand U19601 (N_19601,N_16554,N_17307);
and U19602 (N_19602,N_16492,N_18653);
and U19603 (N_19603,N_16351,N_18231);
nand U19604 (N_19604,N_16056,N_18423);
nor U19605 (N_19605,N_16770,N_18124);
nor U19606 (N_19606,N_18631,N_17457);
or U19607 (N_19607,N_17029,N_17770);
or U19608 (N_19608,N_15790,N_16495);
and U19609 (N_19609,N_17159,N_17685);
nor U19610 (N_19610,N_15811,N_18357);
and U19611 (N_19611,N_15736,N_15781);
nor U19612 (N_19612,N_15664,N_18582);
and U19613 (N_19613,N_16431,N_17649);
nor U19614 (N_19614,N_18591,N_18497);
and U19615 (N_19615,N_17489,N_16659);
nand U19616 (N_19616,N_17623,N_18061);
xnor U19617 (N_19617,N_18387,N_17915);
xnor U19618 (N_19618,N_16267,N_16799);
nor U19619 (N_19619,N_16327,N_16530);
nor U19620 (N_19620,N_16217,N_15986);
xnor U19621 (N_19621,N_17105,N_18296);
or U19622 (N_19622,N_16979,N_17829);
and U19623 (N_19623,N_18379,N_16121);
or U19624 (N_19624,N_18656,N_17662);
xor U19625 (N_19625,N_16183,N_17466);
and U19626 (N_19626,N_17977,N_16732);
nor U19627 (N_19627,N_17092,N_17196);
nand U19628 (N_19628,N_17269,N_16221);
and U19629 (N_19629,N_17577,N_17792);
or U19630 (N_19630,N_17021,N_18123);
or U19631 (N_19631,N_17707,N_16108);
nand U19632 (N_19632,N_17833,N_16093);
and U19633 (N_19633,N_17534,N_17464);
nand U19634 (N_19634,N_15817,N_17443);
xnor U19635 (N_19635,N_17239,N_16048);
xor U19636 (N_19636,N_17979,N_17816);
or U19637 (N_19637,N_16922,N_18745);
xor U19638 (N_19638,N_17493,N_17961);
or U19639 (N_19639,N_18221,N_16235);
or U19640 (N_19640,N_16587,N_18737);
nand U19641 (N_19641,N_18287,N_16998);
xnor U19642 (N_19642,N_17251,N_16016);
or U19643 (N_19643,N_17188,N_15804);
nand U19644 (N_19644,N_17362,N_17949);
and U19645 (N_19645,N_15767,N_16913);
and U19646 (N_19646,N_16364,N_18049);
or U19647 (N_19647,N_17299,N_17061);
nor U19648 (N_19648,N_17542,N_18392);
nand U19649 (N_19649,N_16813,N_17779);
nand U19650 (N_19650,N_16297,N_18018);
and U19651 (N_19651,N_18395,N_18303);
xor U19652 (N_19652,N_15669,N_17426);
or U19653 (N_19653,N_16375,N_16816);
xor U19654 (N_19654,N_18663,N_16858);
nand U19655 (N_19655,N_15955,N_17899);
and U19656 (N_19656,N_17397,N_15865);
nand U19657 (N_19657,N_16744,N_16044);
nor U19658 (N_19658,N_18495,N_17936);
nand U19659 (N_19659,N_18354,N_15892);
and U19660 (N_19660,N_18599,N_18370);
nand U19661 (N_19661,N_17208,N_16653);
nand U19662 (N_19662,N_16973,N_18429);
nand U19663 (N_19663,N_16087,N_18176);
nand U19664 (N_19664,N_17843,N_15780);
nand U19665 (N_19665,N_16837,N_17680);
and U19666 (N_19666,N_17653,N_15828);
and U19667 (N_19667,N_16139,N_16489);
xnor U19668 (N_19668,N_16429,N_17051);
nand U19669 (N_19669,N_17383,N_17404);
xor U19670 (N_19670,N_17722,N_17126);
or U19671 (N_19671,N_16212,N_15979);
or U19672 (N_19672,N_18159,N_17911);
or U19673 (N_19673,N_16192,N_17918);
xor U19674 (N_19674,N_15752,N_16163);
nand U19675 (N_19675,N_18372,N_15729);
or U19676 (N_19676,N_16153,N_16866);
nand U19677 (N_19677,N_17135,N_16115);
nand U19678 (N_19678,N_17058,N_17826);
or U19679 (N_19679,N_16553,N_17605);
nor U19680 (N_19680,N_17197,N_16103);
nand U19681 (N_19681,N_16930,N_15738);
nand U19682 (N_19682,N_16576,N_16647);
nor U19683 (N_19683,N_16549,N_18006);
nand U19684 (N_19684,N_17500,N_16010);
and U19685 (N_19685,N_18168,N_16623);
nor U19686 (N_19686,N_18701,N_18251);
nor U19687 (N_19687,N_17080,N_17578);
or U19688 (N_19688,N_17717,N_15863);
and U19689 (N_19689,N_18660,N_16559);
or U19690 (N_19690,N_17681,N_18157);
and U19691 (N_19691,N_15741,N_16743);
nor U19692 (N_19692,N_16299,N_18440);
nor U19693 (N_19693,N_16278,N_16443);
nor U19694 (N_19694,N_16046,N_18412);
and U19695 (N_19695,N_16864,N_18487);
and U19696 (N_19696,N_15882,N_17160);
xnor U19697 (N_19697,N_18611,N_16437);
or U19698 (N_19698,N_15896,N_17872);
and U19699 (N_19699,N_18527,N_16996);
or U19700 (N_19700,N_18646,N_15886);
nor U19701 (N_19701,N_15773,N_16757);
nand U19702 (N_19702,N_18405,N_17298);
nand U19703 (N_19703,N_16222,N_15918);
nor U19704 (N_19704,N_16461,N_16581);
and U19705 (N_19705,N_16300,N_17046);
or U19706 (N_19706,N_16240,N_17503);
and U19707 (N_19707,N_16265,N_16017);
or U19708 (N_19708,N_15970,N_16231);
or U19709 (N_19709,N_15953,N_16546);
nand U19710 (N_19710,N_17907,N_17415);
nand U19711 (N_19711,N_17712,N_18201);
and U19712 (N_19712,N_18413,N_17790);
or U19713 (N_19713,N_15829,N_17449);
or U19714 (N_19714,N_17962,N_17052);
or U19715 (N_19715,N_16642,N_17250);
and U19716 (N_19716,N_15678,N_18161);
nand U19717 (N_19717,N_16542,N_18248);
xor U19718 (N_19718,N_18373,N_16882);
or U19719 (N_19719,N_17465,N_17599);
xnor U19720 (N_19720,N_18404,N_17675);
or U19721 (N_19721,N_16112,N_16630);
and U19722 (N_19722,N_18144,N_16739);
nor U19723 (N_19723,N_15748,N_18614);
xor U19724 (N_19724,N_16109,N_17206);
nor U19725 (N_19725,N_18191,N_16823);
nor U19726 (N_19726,N_16600,N_15758);
or U19727 (N_19727,N_18564,N_16758);
nand U19728 (N_19728,N_18517,N_15830);
and U19729 (N_19729,N_16740,N_17965);
or U19730 (N_19730,N_18344,N_18353);
nor U19731 (N_19731,N_16382,N_16147);
nor U19732 (N_19732,N_17252,N_17973);
nor U19733 (N_19733,N_18450,N_16365);
or U19734 (N_19734,N_16601,N_17007);
nand U19735 (N_19735,N_18368,N_17539);
nand U19736 (N_19736,N_17030,N_16230);
and U19737 (N_19737,N_16694,N_16658);
and U19738 (N_19738,N_16824,N_16194);
and U19739 (N_19739,N_18252,N_18237);
nand U19740 (N_19740,N_17060,N_16952);
or U19741 (N_19741,N_16236,N_15755);
or U19742 (N_19742,N_15917,N_18539);
nand U19743 (N_19743,N_18416,N_17590);
nand U19744 (N_19744,N_17134,N_18578);
nor U19745 (N_19745,N_16394,N_16475);
or U19746 (N_19746,N_15950,N_17706);
and U19747 (N_19747,N_18065,N_16971);
nand U19748 (N_19748,N_17437,N_18431);
or U19749 (N_19749,N_16874,N_18131);
and U19750 (N_19750,N_16992,N_15968);
nand U19751 (N_19751,N_15737,N_17905);
nor U19752 (N_19752,N_17688,N_15821);
nor U19753 (N_19753,N_18560,N_18512);
or U19754 (N_19754,N_18002,N_16876);
and U19755 (N_19755,N_17448,N_17950);
nand U19756 (N_19756,N_18689,N_18326);
nor U19757 (N_19757,N_16286,N_16891);
nor U19758 (N_19758,N_17644,N_17445);
nor U19759 (N_19759,N_16346,N_17189);
nand U19760 (N_19760,N_17700,N_16738);
or U19761 (N_19761,N_16707,N_16932);
or U19762 (N_19762,N_16342,N_15641);
nor U19763 (N_19763,N_17930,N_18340);
or U19764 (N_19764,N_16392,N_16438);
or U19765 (N_19765,N_17788,N_18059);
and U19766 (N_19766,N_15934,N_18118);
and U19767 (N_19767,N_15635,N_17541);
nor U19768 (N_19768,N_18515,N_17428);
nor U19769 (N_19769,N_15898,N_16812);
nand U19770 (N_19770,N_17427,N_17203);
nor U19771 (N_19771,N_16485,N_16970);
nor U19772 (N_19772,N_16860,N_18725);
nand U19773 (N_19773,N_18163,N_17347);
nand U19774 (N_19774,N_16069,N_18603);
and U19775 (N_19775,N_18347,N_16742);
xnor U19776 (N_19776,N_17696,N_18329);
or U19777 (N_19777,N_15798,N_18014);
and U19778 (N_19778,N_18471,N_15766);
and U19779 (N_19779,N_16620,N_16632);
nor U19780 (N_19780,N_16233,N_18011);
or U19781 (N_19781,N_17511,N_17054);
nand U19782 (N_19782,N_17876,N_17778);
xor U19783 (N_19783,N_16771,N_18568);
nor U19784 (N_19784,N_16301,N_17853);
nor U19785 (N_19785,N_16895,N_17398);
nand U19786 (N_19786,N_17195,N_17714);
nor U19787 (N_19787,N_17863,N_15944);
nor U19788 (N_19788,N_16978,N_17407);
nand U19789 (N_19789,N_18244,N_17485);
and U19790 (N_19790,N_16169,N_17811);
or U19791 (N_19791,N_18543,N_16990);
nor U19792 (N_19792,N_18225,N_16434);
or U19793 (N_19793,N_18473,N_17693);
and U19794 (N_19794,N_15991,N_16759);
nor U19795 (N_19795,N_17992,N_16241);
and U19796 (N_19796,N_15985,N_16136);
and U19797 (N_19797,N_16366,N_17669);
nand U19798 (N_19798,N_15922,N_15873);
and U19799 (N_19799,N_17957,N_17708);
or U19800 (N_19800,N_18069,N_17277);
and U19801 (N_19801,N_16709,N_16399);
nand U19802 (N_19802,N_17724,N_17139);
nand U19803 (N_19803,N_16925,N_17801);
and U19804 (N_19804,N_17028,N_17481);
or U19805 (N_19805,N_17390,N_18436);
nand U19806 (N_19806,N_17309,N_18343);
xnor U19807 (N_19807,N_17301,N_17033);
and U19808 (N_19808,N_16531,N_15695);
and U19809 (N_19809,N_16023,N_16030);
nor U19810 (N_19810,N_17602,N_16612);
nor U19811 (N_19811,N_16237,N_16908);
and U19812 (N_19812,N_16329,N_18605);
and U19813 (N_19813,N_17144,N_16691);
xnor U19814 (N_19814,N_16339,N_16203);
nor U19815 (N_19815,N_17994,N_16435);
or U19816 (N_19816,N_15791,N_17987);
nand U19817 (N_19817,N_17230,N_17225);
and U19818 (N_19818,N_16765,N_16784);
and U19819 (N_19819,N_17193,N_17349);
xor U19820 (N_19820,N_16869,N_18262);
nor U19821 (N_19821,N_17263,N_16698);
and U19822 (N_19822,N_18179,N_18394);
nand U19823 (N_19823,N_18554,N_17204);
nand U19824 (N_19824,N_16797,N_18261);
xnor U19825 (N_19825,N_16189,N_15903);
and U19826 (N_19826,N_17451,N_16076);
nand U19827 (N_19827,N_18478,N_16618);
xor U19828 (N_19828,N_18541,N_16226);
nor U19829 (N_19829,N_17727,N_16609);
and U19830 (N_19830,N_16841,N_17235);
or U19831 (N_19831,N_17975,N_16065);
nor U19832 (N_19832,N_16287,N_16262);
or U19833 (N_19833,N_16939,N_17297);
nand U19834 (N_19834,N_18140,N_16040);
nand U19835 (N_19835,N_17745,N_15800);
nand U19836 (N_19836,N_16446,N_16800);
and U19837 (N_19837,N_18378,N_15805);
nor U19838 (N_19838,N_15856,N_17893);
or U19839 (N_19839,N_16047,N_16319);
nand U19840 (N_19840,N_18596,N_17651);
nor U19841 (N_19841,N_17441,N_17533);
nor U19842 (N_19842,N_17557,N_16385);
nor U19843 (N_19843,N_15802,N_17056);
or U19844 (N_19844,N_17146,N_16369);
nand U19845 (N_19845,N_16867,N_16745);
or U19846 (N_19846,N_15984,N_17852);
xor U19847 (N_19847,N_16909,N_16165);
and U19848 (N_19848,N_16116,N_17625);
and U19849 (N_19849,N_15849,N_18408);
and U19850 (N_19850,N_16843,N_15746);
nor U19851 (N_19851,N_17439,N_16381);
or U19852 (N_19852,N_16083,N_18232);
nand U19853 (N_19853,N_16075,N_17190);
and U19854 (N_19854,N_18612,N_16616);
or U19855 (N_19855,N_16597,N_15816);
and U19856 (N_19856,N_17532,N_16263);
or U19857 (N_19857,N_16387,N_17774);
and U19858 (N_19858,N_15739,N_16897);
nand U19859 (N_19859,N_16753,N_16836);
or U19860 (N_19860,N_18642,N_18662);
nor U19861 (N_19861,N_18070,N_15850);
nor U19862 (N_19862,N_17601,N_18336);
nor U19863 (N_19863,N_18182,N_17569);
or U19864 (N_19864,N_15943,N_18585);
or U19865 (N_19865,N_18009,N_17078);
or U19866 (N_19866,N_16318,N_15960);
and U19867 (N_19867,N_18620,N_18192);
nor U19868 (N_19868,N_17219,N_18575);
nand U19869 (N_19869,N_18654,N_18608);
nor U19870 (N_19870,N_17348,N_18492);
nor U19871 (N_19871,N_15645,N_16101);
and U19872 (N_19872,N_16785,N_18519);
nand U19873 (N_19873,N_16781,N_16106);
or U19874 (N_19874,N_15846,N_16207);
nor U19875 (N_19875,N_18366,N_16507);
or U19876 (N_19876,N_16599,N_18730);
and U19877 (N_19877,N_17093,N_16271);
nand U19878 (N_19878,N_17136,N_17177);
or U19879 (N_19879,N_17468,N_17540);
or U19880 (N_19880,N_18703,N_16575);
nand U19881 (N_19881,N_15928,N_17988);
nand U19882 (N_19882,N_18374,N_17388);
nor U19883 (N_19883,N_16668,N_15845);
and U19884 (N_19884,N_17129,N_16462);
or U19885 (N_19885,N_16562,N_16778);
or U19886 (N_19886,N_18452,N_17118);
xor U19887 (N_19887,N_16254,N_16534);
nor U19888 (N_19888,N_18628,N_17786);
nor U19889 (N_19889,N_18466,N_18156);
nor U19890 (N_19890,N_15824,N_16540);
nand U19891 (N_19891,N_16457,N_15648);
nand U19892 (N_19892,N_18255,N_18238);
nand U19893 (N_19893,N_17243,N_18402);
nor U19894 (N_19894,N_18055,N_16648);
nor U19895 (N_19895,N_16723,N_16544);
or U19896 (N_19896,N_16468,N_18729);
and U19897 (N_19897,N_17809,N_16714);
and U19898 (N_19898,N_17737,N_16810);
and U19899 (N_19899,N_16474,N_16955);
and U19900 (N_19900,N_16019,N_18377);
and U19901 (N_19901,N_16049,N_15957);
nand U19902 (N_19902,N_17344,N_18186);
or U19903 (N_19903,N_18127,N_18384);
nor U19904 (N_19904,N_16847,N_16894);
nand U19905 (N_19905,N_17646,N_16906);
or U19906 (N_19906,N_17518,N_16282);
or U19907 (N_19907,N_18572,N_16700);
or U19908 (N_19908,N_15947,N_17303);
nor U19909 (N_19909,N_18442,N_16631);
or U19910 (N_19910,N_17358,N_16501);
nand U19911 (N_19911,N_18292,N_17127);
nand U19912 (N_19912,N_18205,N_18479);
or U19913 (N_19913,N_16972,N_18345);
or U19914 (N_19914,N_16705,N_18364);
and U19915 (N_19915,N_17042,N_17887);
or U19916 (N_19916,N_16325,N_16317);
nand U19917 (N_19917,N_18242,N_15633);
or U19918 (N_19918,N_17474,N_17596);
nand U19919 (N_19919,N_16675,N_17490);
and U19920 (N_19920,N_16580,N_15723);
and U19921 (N_19921,N_17313,N_16914);
and U19922 (N_19922,N_16362,N_16769);
nand U19923 (N_19923,N_16145,N_15975);
nor U19924 (N_19924,N_18291,N_17769);
or U19925 (N_19925,N_18053,N_16855);
or U19926 (N_19926,N_17454,N_15901);
and U19927 (N_19927,N_18533,N_16187);
nand U19928 (N_19928,N_16334,N_15670);
nand U19929 (N_19929,N_17888,N_18295);
and U19930 (N_19930,N_17740,N_18532);
and U19931 (N_19931,N_16268,N_17444);
xnor U19932 (N_19932,N_18360,N_18643);
or U19933 (N_19933,N_17112,N_15869);
and U19934 (N_19934,N_17971,N_17728);
nand U19935 (N_19935,N_16762,N_16479);
and U19936 (N_19936,N_18275,N_18116);
and U19937 (N_19937,N_18233,N_17677);
nand U19938 (N_19938,N_17094,N_16592);
xor U19939 (N_19939,N_17764,N_16336);
and U19940 (N_19940,N_16379,N_17356);
and U19941 (N_19941,N_17280,N_18169);
or U19942 (N_19942,N_16456,N_16539);
nor U19943 (N_19943,N_15983,N_18273);
or U19944 (N_19944,N_16833,N_16333);
or U19945 (N_19945,N_17990,N_18008);
or U19946 (N_19946,N_17900,N_16419);
and U19947 (N_19947,N_16617,N_17694);
nor U19948 (N_19948,N_16683,N_16856);
nor U19949 (N_19949,N_17413,N_16938);
nand U19950 (N_19950,N_18391,N_16989);
or U19951 (N_19951,N_18569,N_16360);
and U19952 (N_19952,N_15700,N_16590);
nand U19953 (N_19953,N_17771,N_17620);
nand U19954 (N_19954,N_17002,N_16988);
nand U19955 (N_19955,N_17273,N_18506);
or U19956 (N_19956,N_17749,N_16755);
nand U19957 (N_19957,N_16015,N_16257);
nor U19958 (N_19958,N_17387,N_16242);
and U19959 (N_19959,N_17839,N_17015);
nand U19960 (N_19960,N_17067,N_15640);
nand U19961 (N_19961,N_18234,N_16598);
nor U19962 (N_19962,N_17075,N_17482);
and U19963 (N_19963,N_17802,N_15951);
nor U19964 (N_19964,N_15761,N_18468);
or U19965 (N_19965,N_16923,N_17419);
xor U19966 (N_19966,N_17579,N_17898);
nor U19967 (N_19967,N_16652,N_16051);
nor U19968 (N_19968,N_18341,N_16893);
nor U19969 (N_19969,N_17213,N_15897);
nor U19970 (N_19970,N_17257,N_18020);
and U19971 (N_19971,N_17628,N_17929);
and U19972 (N_19972,N_16273,N_16628);
or U19973 (N_19973,N_16350,N_16227);
nand U19974 (N_19974,N_15732,N_16878);
nand U19975 (N_19975,N_17434,N_15927);
or U19976 (N_19976,N_16401,N_18171);
nand U19977 (N_19977,N_18226,N_16883);
nor U19978 (N_19978,N_18003,N_15660);
nor U19979 (N_19979,N_15883,N_18467);
nor U19980 (N_19980,N_18174,N_16650);
nand U19981 (N_19981,N_17166,N_16584);
or U19982 (N_19982,N_16967,N_18544);
or U19983 (N_19983,N_17162,N_16935);
xor U19984 (N_19984,N_16900,N_18046);
nand U19985 (N_19985,N_17978,N_17319);
nand U19986 (N_19986,N_17775,N_17343);
nand U19987 (N_19987,N_17803,N_17487);
nand U19988 (N_19988,N_17385,N_17997);
nor U19989 (N_19989,N_17430,N_18213);
nand U19990 (N_19990,N_16718,N_17435);
nor U19991 (N_19991,N_15733,N_18383);
nand U19992 (N_19992,N_18024,N_15665);
nor U19993 (N_19993,N_16514,N_15844);
nand U19994 (N_19994,N_16995,N_17360);
nor U19995 (N_19995,N_16827,N_16398);
nor U19996 (N_19996,N_17765,N_17107);
nor U19997 (N_19997,N_16059,N_16432);
and U19998 (N_19998,N_18721,N_17179);
nand U19999 (N_19999,N_15980,N_18269);
xor U20000 (N_20000,N_18503,N_18090);
nor U20001 (N_20001,N_17819,N_15785);
or U20002 (N_20002,N_18570,N_16566);
and U20003 (N_20003,N_17149,N_16111);
nand U20004 (N_20004,N_16250,N_17246);
nand U20005 (N_20005,N_18499,N_17452);
nor U20006 (N_20006,N_18469,N_16746);
nand U20007 (N_20007,N_17290,N_16427);
or U20008 (N_20008,N_18692,N_17908);
and U20009 (N_20009,N_17400,N_17776);
and U20010 (N_20010,N_16901,N_15987);
and U20011 (N_20011,N_16095,N_17945);
and U20012 (N_20012,N_17287,N_16552);
or U20013 (N_20013,N_18155,N_18306);
and U20014 (N_20014,N_15906,N_17455);
and U20015 (N_20015,N_16216,N_17103);
or U20016 (N_20016,N_17086,N_17964);
and U20017 (N_20017,N_17063,N_17640);
or U20018 (N_20018,N_16493,N_15899);
or U20019 (N_20019,N_17165,N_18735);
nor U20020 (N_20020,N_16993,N_16368);
or U20021 (N_20021,N_16889,N_16574);
nand U20022 (N_20022,N_17812,N_17513);
nor U20023 (N_20023,N_17425,N_17951);
and U20024 (N_20024,N_16452,N_17526);
or U20025 (N_20025,N_15990,N_17743);
nand U20026 (N_20026,N_18713,N_18050);
nor U20027 (N_20027,N_16947,N_16245);
and U20028 (N_20028,N_17505,N_18184);
and U20029 (N_20029,N_18583,N_18083);
nor U20030 (N_20030,N_16766,N_18259);
and U20031 (N_20031,N_16098,N_16100);
and U20032 (N_20032,N_16725,N_18245);
and U20033 (N_20033,N_16912,N_15961);
nand U20034 (N_20034,N_17873,N_17960);
nor U20035 (N_20035,N_16532,N_17391);
nor U20036 (N_20036,N_18196,N_17423);
and U20037 (N_20037,N_15663,N_17943);
nor U20038 (N_20038,N_17713,N_16656);
and U20039 (N_20039,N_18013,N_17097);
and U20040 (N_20040,N_17701,N_17327);
and U20041 (N_20041,N_16657,N_18615);
nor U20042 (N_20042,N_18494,N_15656);
nand U20043 (N_20043,N_16138,N_18489);
and U20044 (N_20044,N_17339,N_18627);
xnor U20045 (N_20045,N_18236,N_15977);
nor U20046 (N_20046,N_16210,N_16750);
nand U20047 (N_20047,N_18454,N_15717);
nor U20048 (N_20048,N_17365,N_15921);
or U20049 (N_20049,N_16312,N_17797);
nor U20050 (N_20050,N_17535,N_15919);
nor U20051 (N_20051,N_15854,N_18448);
and U20052 (N_20052,N_18434,N_18129);
xor U20053 (N_20053,N_18708,N_16677);
or U20054 (N_20054,N_17044,N_18324);
nor U20055 (N_20055,N_16887,N_16487);
or U20056 (N_20056,N_16062,N_17610);
nand U20057 (N_20057,N_18587,N_16693);
nor U20058 (N_20058,N_16543,N_16092);
nor U20059 (N_20059,N_15812,N_18304);
nand U20060 (N_20060,N_15701,N_17154);
nand U20061 (N_20061,N_17048,N_16455);
nor U20062 (N_20062,N_17832,N_16261);
nand U20063 (N_20063,N_15647,N_18537);
or U20064 (N_20064,N_18650,N_16701);
nor U20065 (N_20065,N_18670,N_18514);
and U20066 (N_20066,N_18240,N_18748);
nand U20067 (N_20067,N_15877,N_15768);
and U20068 (N_20068,N_18331,N_17174);
and U20069 (N_20069,N_15876,N_18048);
or U20070 (N_20070,N_17100,N_16383);
nor U20071 (N_20071,N_18741,N_16728);
or U20072 (N_20072,N_16591,N_16198);
or U20073 (N_20073,N_15827,N_15778);
or U20074 (N_20074,N_17781,N_16188);
or U20075 (N_20075,N_16422,N_17972);
or U20076 (N_20076,N_17583,N_17376);
nand U20077 (N_20077,N_18325,N_16556);
and U20078 (N_20078,N_16345,N_18655);
or U20079 (N_20079,N_17236,N_17314);
or U20080 (N_20080,N_18029,N_16170);
nand U20081 (N_20081,N_16510,N_17734);
and U20082 (N_20082,N_16814,N_18460);
nor U20083 (N_20083,N_15792,N_17624);
and U20084 (N_20084,N_17119,N_18561);
xor U20085 (N_20085,N_16627,N_16372);
and U20086 (N_20086,N_17321,N_16699);
xor U20087 (N_20087,N_17492,N_18352);
nand U20088 (N_20088,N_16904,N_17575);
xor U20089 (N_20089,N_15973,N_15706);
nor U20090 (N_20090,N_15895,N_18711);
xor U20091 (N_20091,N_17842,N_18459);
and U20092 (N_20092,N_16767,N_18062);
nand U20093 (N_20093,N_18365,N_18716);
and U20094 (N_20094,N_18389,N_16917);
or U20095 (N_20095,N_15685,N_16638);
xnor U20096 (N_20096,N_17958,N_16397);
or U20097 (N_20097,N_17633,N_18680);
and U20098 (N_20098,N_16412,N_17799);
nand U20099 (N_20099,N_18491,N_17070);
nor U20100 (N_20100,N_18594,N_15888);
or U20101 (N_20101,N_18081,N_18709);
or U20102 (N_20102,N_16681,N_16054);
and U20103 (N_20103,N_15697,N_16266);
nand U20104 (N_20104,N_17248,N_16224);
nand U20105 (N_20105,N_16936,N_16148);
nand U20106 (N_20106,N_17691,N_16463);
and U20107 (N_20107,N_18031,N_17746);
or U20108 (N_20108,N_17184,N_17375);
nor U20109 (N_20109,N_17040,N_17265);
nor U20110 (N_20110,N_16373,N_16285);
or U20111 (N_20111,N_16536,N_18359);
and U20112 (N_20112,N_16042,N_17984);
or U20113 (N_20113,N_18211,N_16084);
and U20114 (N_20114,N_16159,N_17830);
nor U20115 (N_20115,N_17320,N_18490);
and U20116 (N_20116,N_17516,N_16515);
nand U20117 (N_20117,N_17798,N_15894);
nand U20118 (N_20118,N_17281,N_16661);
xor U20119 (N_20119,N_18731,N_17300);
or U20120 (N_20120,N_16749,N_17255);
nor U20121 (N_20121,N_17509,N_16491);
nand U20122 (N_20122,N_17910,N_18267);
nor U20123 (N_20123,N_18339,N_17867);
nor U20124 (N_20124,N_17410,N_16464);
nor U20125 (N_20125,N_16880,N_16666);
nand U20126 (N_20126,N_16871,N_16826);
and U20127 (N_20127,N_17565,N_17603);
nor U20128 (N_20128,N_16966,N_17214);
or U20129 (N_20129,N_17394,N_17461);
or U20130 (N_20130,N_16941,N_17342);
or U20131 (N_20131,N_16595,N_15764);
and U20132 (N_20132,N_17985,N_18563);
and U20133 (N_20133,N_17550,N_15963);
nor U20134 (N_20134,N_16747,N_18263);
nand U20135 (N_20135,N_15801,N_17153);
or U20136 (N_20136,N_18702,N_16199);
nand U20137 (N_20137,N_18435,N_18004);
and U20138 (N_20138,N_18547,N_17270);
or U20139 (N_20139,N_16835,N_17862);
nor U20140 (N_20140,N_17638,N_18113);
nor U20141 (N_20141,N_16409,N_16353);
nand U20142 (N_20142,N_18087,N_17220);
nor U20143 (N_20143,N_17411,N_18719);
xnor U20144 (N_20144,N_18606,N_15765);
or U20145 (N_20145,N_16608,N_15904);
or U20146 (N_20146,N_16667,N_15735);
xor U20147 (N_20147,N_17923,N_16717);
nor U20148 (N_20148,N_15719,N_17024);
or U20149 (N_20149,N_16818,N_18456);
nand U20150 (N_20150,N_17866,N_18036);
nand U20151 (N_20151,N_18342,N_17357);
and U20152 (N_20152,N_17824,N_18504);
nor U20153 (N_20153,N_18613,N_16787);
nand U20154 (N_20154,N_17181,N_16164);
and U20155 (N_20155,N_17496,N_17484);
xnor U20156 (N_20156,N_16509,N_17544);
nor U20157 (N_20157,N_16057,N_18111);
xor U20158 (N_20158,N_18453,N_15627);
nand U20159 (N_20159,N_17844,N_15730);
or U20160 (N_20160,N_17660,N_18595);
xor U20161 (N_20161,N_16478,N_16408);
and U20162 (N_20162,N_16484,N_16337);
or U20163 (N_20163,N_17690,N_17510);
or U20164 (N_20164,N_16672,N_17626);
or U20165 (N_20165,N_16182,N_18030);
or U20166 (N_20166,N_18042,N_17101);
or U20167 (N_20167,N_18557,N_17870);
nor U20168 (N_20168,N_17969,N_15742);
nor U20169 (N_20169,N_16805,N_16150);
nor U20170 (N_20170,N_18332,N_17879);
and U20171 (N_20171,N_18688,N_18102);
nor U20172 (N_20172,N_17783,N_18022);
and U20173 (N_20173,N_17158,N_16149);
and U20174 (N_20174,N_16822,N_18424);
or U20175 (N_20175,N_17479,N_18421);
and U20176 (N_20176,N_16004,N_18505);
nand U20177 (N_20177,N_16720,N_18197);
nand U20178 (N_20178,N_16829,N_18588);
or U20179 (N_20179,N_15782,N_16606);
nand U20180 (N_20180,N_15721,N_16225);
or U20181 (N_20181,N_16068,N_16055);
xnor U20182 (N_20182,N_16155,N_17371);
and U20183 (N_20183,N_17294,N_18057);
nand U20184 (N_20184,N_17606,N_18444);
nand U20185 (N_20185,N_18736,N_16344);
xor U20186 (N_20186,N_18428,N_18648);
or U20187 (N_20187,N_16161,N_17567);
and U20188 (N_20188,N_17573,N_15871);
and U20189 (N_20189,N_16007,N_17944);
nor U20190 (N_20190,N_17937,N_18200);
or U20191 (N_20191,N_15912,N_17053);
or U20192 (N_20192,N_15725,N_16626);
xor U20193 (N_20193,N_16290,N_16840);
or U20194 (N_20194,N_17175,N_16190);
nand U20195 (N_20195,N_18633,N_16140);
or U20196 (N_20196,N_16854,N_16073);
nor U20197 (N_20197,N_17226,N_16323);
nor U20198 (N_20198,N_16692,N_17083);
nor U20199 (N_20199,N_15772,N_17308);
nand U20200 (N_20200,N_17128,N_18700);
xor U20201 (N_20201,N_18044,N_17891);
or U20202 (N_20202,N_17901,N_16577);
nand U20203 (N_20203,N_17209,N_18507);
nand U20204 (N_20204,N_15705,N_18058);
nor U20205 (N_20205,N_15692,N_16567);
nor U20206 (N_20206,N_18559,N_17524);
and U20207 (N_20207,N_16028,N_17607);
or U20208 (N_20208,N_15885,N_17141);
or U20209 (N_20209,N_16968,N_15789);
nor U20210 (N_20210,N_18593,N_17718);
xor U20211 (N_20211,N_18699,N_18530);
nor U20212 (N_20212,N_17922,N_18446);
nor U20213 (N_20213,N_16288,N_16196);
or U20214 (N_20214,N_15680,N_16488);
nor U20215 (N_20215,N_15926,N_17480);
nand U20216 (N_20216,N_17904,N_18217);
nand U20217 (N_20217,N_16063,N_18356);
and U20218 (N_20218,N_17858,N_18695);
and U20219 (N_20219,N_16218,N_18108);
nand U20220 (N_20220,N_17279,N_17245);
nor U20221 (N_20221,N_17157,N_16902);
nor U20222 (N_20222,N_17894,N_18521);
or U20223 (N_20223,N_16018,N_16937);
nor U20224 (N_20224,N_16298,N_17970);
nor U20225 (N_20225,N_16792,N_16708);
nor U20226 (N_20226,N_17941,N_16081);
xor U20227 (N_20227,N_17678,N_17546);
nor U20228 (N_20228,N_18738,N_17059);
nor U20229 (N_20229,N_16888,N_18190);
or U20230 (N_20230,N_17150,N_18411);
nand U20231 (N_20231,N_17361,N_15825);
and U20232 (N_20232,N_15690,N_16086);
nand U20233 (N_20233,N_16052,N_16071);
nand U20234 (N_20234,N_17218,N_16074);
and U20235 (N_20235,N_17673,N_16846);
nand U20236 (N_20236,N_18094,N_17041);
nor U20237 (N_20237,N_16122,N_18322);
or U20238 (N_20238,N_17109,N_18617);
nor U20239 (N_20239,N_17262,N_18657);
nor U20240 (N_20240,N_18581,N_16526);
nor U20241 (N_20241,N_18056,N_17462);
xnor U20242 (N_20242,N_17207,N_16091);
or U20243 (N_20243,N_18223,N_17656);
nand U20244 (N_20244,N_18396,N_18513);
or U20245 (N_20245,N_16426,N_17325);
and U20246 (N_20246,N_17933,N_17138);
and U20247 (N_20247,N_15808,N_15924);
or U20248 (N_20248,N_17772,N_17952);
nand U20249 (N_20249,N_17036,N_16563);
nor U20250 (N_20250,N_17478,N_18742);
nand U20251 (N_20251,N_17332,N_16064);
or U20252 (N_20252,N_16980,N_17161);
nor U20253 (N_20253,N_18330,N_18215);
and U20254 (N_20254,N_15880,N_18302);
and U20255 (N_20255,N_18734,N_17183);
and U20256 (N_20256,N_16654,N_17598);
nor U20257 (N_20257,N_18616,N_16072);
xor U20258 (N_20258,N_18696,N_18439);
nand U20259 (N_20259,N_15875,N_15677);
nand U20260 (N_20260,N_16482,N_16439);
nand U20261 (N_20261,N_16558,N_16027);
and U20262 (N_20262,N_16331,N_17288);
xor U20263 (N_20263,N_17221,N_16832);
and U20264 (N_20264,N_16673,N_17310);
and U20265 (N_20265,N_18407,N_17611);
nor U20266 (N_20266,N_18208,N_18114);
nand U20267 (N_20267,N_17502,N_16277);
nor U20268 (N_20268,N_17619,N_18119);
nand U20269 (N_20269,N_18281,N_15810);
nand U20270 (N_20270,N_16756,N_16305);
nand U20271 (N_20271,N_18101,N_18165);
nand U20272 (N_20272,N_17120,N_16402);
nand U20273 (N_20273,N_18272,N_15657);
xor U20274 (N_20274,N_18432,N_16184);
nand U20275 (N_20275,N_15672,N_16494);
and U20276 (N_20276,N_16527,N_16986);
nor U20277 (N_20277,N_17849,N_18470);
nor U20278 (N_20278,N_17880,N_17240);
nand U20279 (N_20279,N_17212,N_17163);
and U20280 (N_20280,N_16107,N_17306);
or U20281 (N_20281,N_16384,N_17558);
and U20282 (N_20282,N_18162,N_16674);
or U20283 (N_20283,N_16376,N_16715);
or U20284 (N_20284,N_16857,N_17215);
xor U20285 (N_20285,N_17004,N_18607);
xnor U20286 (N_20286,N_17124,N_18195);
nand U20287 (N_20287,N_18034,N_16852);
nand U20288 (N_20288,N_16272,N_16634);
nor U20289 (N_20289,N_18117,N_18546);
nand U20290 (N_20290,N_16927,N_15834);
and U20291 (N_20291,N_16896,N_17909);
nand U20292 (N_20292,N_17311,N_18427);
nand U20293 (N_20293,N_15900,N_17291);
nor U20294 (N_20294,N_15933,N_16731);
nor U20295 (N_20295,N_18355,N_17003);
and U20296 (N_20296,N_17760,N_17955);
and U20297 (N_20297,N_17668,N_17125);
or U20298 (N_20298,N_18071,N_17720);
nor U20299 (N_20299,N_15652,N_17850);
nor U20300 (N_20300,N_15783,N_16003);
nor U20301 (N_20301,N_16796,N_17723);
and U20302 (N_20302,N_17055,N_16467);
nand U20303 (N_20303,N_15923,N_18451);
nand U20304 (N_20304,N_17705,N_16070);
nand U20305 (N_20305,N_17178,N_15709);
and U20306 (N_20306,N_17780,N_17587);
and U20307 (N_20307,N_18625,N_16522);
nand U20308 (N_20308,N_17169,N_18222);
or U20309 (N_20309,N_18219,N_17406);
nor U20310 (N_20310,N_18001,N_17982);
nor U20311 (N_20311,N_18481,N_16260);
nand U20312 (N_20312,N_17229,N_18002);
nor U20313 (N_20313,N_18461,N_16650);
xor U20314 (N_20314,N_17057,N_18644);
nand U20315 (N_20315,N_17558,N_18397);
or U20316 (N_20316,N_17078,N_16216);
xnor U20317 (N_20317,N_18131,N_16133);
and U20318 (N_20318,N_16302,N_16752);
xor U20319 (N_20319,N_18209,N_16433);
or U20320 (N_20320,N_18581,N_15840);
nand U20321 (N_20321,N_17631,N_15745);
or U20322 (N_20322,N_16141,N_16756);
nand U20323 (N_20323,N_16816,N_16996);
and U20324 (N_20324,N_18286,N_17312);
and U20325 (N_20325,N_17762,N_16466);
and U20326 (N_20326,N_18361,N_18664);
and U20327 (N_20327,N_18471,N_18403);
or U20328 (N_20328,N_15627,N_17885);
nor U20329 (N_20329,N_16155,N_15691);
and U20330 (N_20330,N_15647,N_18386);
nand U20331 (N_20331,N_17836,N_16745);
or U20332 (N_20332,N_17713,N_17796);
or U20333 (N_20333,N_17581,N_17935);
nor U20334 (N_20334,N_17164,N_17332);
or U20335 (N_20335,N_16001,N_17190);
nand U20336 (N_20336,N_15932,N_18200);
or U20337 (N_20337,N_15839,N_16904);
xor U20338 (N_20338,N_17750,N_16113);
or U20339 (N_20339,N_17891,N_17725);
and U20340 (N_20340,N_17011,N_18344);
and U20341 (N_20341,N_15841,N_16920);
nor U20342 (N_20342,N_15811,N_17010);
nor U20343 (N_20343,N_16390,N_18453);
nor U20344 (N_20344,N_17683,N_17408);
or U20345 (N_20345,N_18422,N_16319);
and U20346 (N_20346,N_18576,N_16853);
nand U20347 (N_20347,N_18123,N_15714);
nor U20348 (N_20348,N_16130,N_16106);
or U20349 (N_20349,N_18615,N_16268);
nor U20350 (N_20350,N_17816,N_18248);
and U20351 (N_20351,N_18546,N_17565);
nand U20352 (N_20352,N_15955,N_16285);
and U20353 (N_20353,N_16056,N_17804);
nor U20354 (N_20354,N_15842,N_17030);
nor U20355 (N_20355,N_16887,N_17464);
or U20356 (N_20356,N_17421,N_18220);
nor U20357 (N_20357,N_17911,N_18341);
nand U20358 (N_20358,N_16983,N_17297);
and U20359 (N_20359,N_16645,N_17060);
or U20360 (N_20360,N_16798,N_16303);
and U20361 (N_20361,N_16254,N_18127);
nand U20362 (N_20362,N_16423,N_17340);
and U20363 (N_20363,N_18232,N_17924);
and U20364 (N_20364,N_16095,N_17974);
nor U20365 (N_20365,N_15684,N_17740);
and U20366 (N_20366,N_17555,N_16670);
and U20367 (N_20367,N_15917,N_17598);
nand U20368 (N_20368,N_17385,N_18549);
nor U20369 (N_20369,N_17102,N_16055);
or U20370 (N_20370,N_17860,N_18704);
and U20371 (N_20371,N_15774,N_18148);
and U20372 (N_20372,N_17987,N_17791);
nand U20373 (N_20373,N_17741,N_17379);
or U20374 (N_20374,N_16837,N_16292);
and U20375 (N_20375,N_18578,N_17465);
nand U20376 (N_20376,N_15929,N_16236);
or U20377 (N_20377,N_17876,N_16826);
nor U20378 (N_20378,N_16204,N_17117);
xor U20379 (N_20379,N_16395,N_16614);
nor U20380 (N_20380,N_16211,N_17615);
or U20381 (N_20381,N_17031,N_15658);
or U20382 (N_20382,N_16196,N_18523);
and U20383 (N_20383,N_15889,N_18617);
xnor U20384 (N_20384,N_17540,N_18117);
nand U20385 (N_20385,N_17861,N_18115);
nor U20386 (N_20386,N_15828,N_16611);
nand U20387 (N_20387,N_16334,N_16954);
and U20388 (N_20388,N_18265,N_16026);
and U20389 (N_20389,N_17250,N_16037);
and U20390 (N_20390,N_16746,N_18331);
nor U20391 (N_20391,N_15743,N_16255);
nand U20392 (N_20392,N_17766,N_16534);
nor U20393 (N_20393,N_18223,N_16530);
xnor U20394 (N_20394,N_18298,N_18620);
nor U20395 (N_20395,N_16453,N_17748);
xnor U20396 (N_20396,N_16117,N_18565);
nand U20397 (N_20397,N_16992,N_17094);
nor U20398 (N_20398,N_18093,N_16646);
nand U20399 (N_20399,N_16118,N_18327);
and U20400 (N_20400,N_16154,N_17952);
and U20401 (N_20401,N_18702,N_17957);
nand U20402 (N_20402,N_16278,N_17771);
and U20403 (N_20403,N_17917,N_17154);
nand U20404 (N_20404,N_16479,N_17735);
nand U20405 (N_20405,N_16559,N_16492);
or U20406 (N_20406,N_17589,N_18478);
nand U20407 (N_20407,N_17728,N_18058);
nand U20408 (N_20408,N_16089,N_16767);
and U20409 (N_20409,N_16607,N_16041);
nand U20410 (N_20410,N_16291,N_18519);
nand U20411 (N_20411,N_18296,N_18088);
or U20412 (N_20412,N_16214,N_17212);
nor U20413 (N_20413,N_16453,N_15988);
nand U20414 (N_20414,N_17777,N_17728);
and U20415 (N_20415,N_17554,N_17670);
xor U20416 (N_20416,N_17653,N_15738);
and U20417 (N_20417,N_18221,N_15920);
and U20418 (N_20418,N_15804,N_16053);
and U20419 (N_20419,N_16237,N_15966);
and U20420 (N_20420,N_16272,N_17711);
or U20421 (N_20421,N_17778,N_15851);
nand U20422 (N_20422,N_17248,N_17905);
and U20423 (N_20423,N_17985,N_16053);
nand U20424 (N_20424,N_16521,N_15970);
and U20425 (N_20425,N_17745,N_18338);
and U20426 (N_20426,N_16026,N_15672);
nand U20427 (N_20427,N_17507,N_16231);
or U20428 (N_20428,N_17487,N_16449);
nor U20429 (N_20429,N_17266,N_17533);
or U20430 (N_20430,N_17699,N_16784);
or U20431 (N_20431,N_16764,N_16677);
and U20432 (N_20432,N_15652,N_16254);
or U20433 (N_20433,N_17619,N_17726);
and U20434 (N_20434,N_16043,N_16354);
or U20435 (N_20435,N_16820,N_16445);
xor U20436 (N_20436,N_15691,N_15771);
and U20437 (N_20437,N_16911,N_17309);
nor U20438 (N_20438,N_16165,N_15632);
and U20439 (N_20439,N_16205,N_18630);
xor U20440 (N_20440,N_18580,N_16718);
nand U20441 (N_20441,N_17986,N_15960);
and U20442 (N_20442,N_16673,N_16039);
nor U20443 (N_20443,N_18552,N_15919);
nand U20444 (N_20444,N_17335,N_15641);
and U20445 (N_20445,N_17411,N_17123);
xnor U20446 (N_20446,N_18135,N_18614);
nand U20447 (N_20447,N_16040,N_18695);
and U20448 (N_20448,N_17335,N_16733);
nor U20449 (N_20449,N_17157,N_17135);
xnor U20450 (N_20450,N_16018,N_17912);
or U20451 (N_20451,N_17926,N_16538);
and U20452 (N_20452,N_16804,N_18191);
xnor U20453 (N_20453,N_17178,N_18330);
nor U20454 (N_20454,N_16062,N_17184);
and U20455 (N_20455,N_18252,N_15879);
and U20456 (N_20456,N_18002,N_17182);
nand U20457 (N_20457,N_16090,N_18090);
and U20458 (N_20458,N_15835,N_18485);
nand U20459 (N_20459,N_15674,N_17434);
and U20460 (N_20460,N_17081,N_16212);
or U20461 (N_20461,N_17464,N_16810);
and U20462 (N_20462,N_16328,N_18254);
and U20463 (N_20463,N_16573,N_17089);
or U20464 (N_20464,N_16051,N_16884);
nor U20465 (N_20465,N_17583,N_18570);
or U20466 (N_20466,N_18482,N_16901);
and U20467 (N_20467,N_16919,N_18499);
and U20468 (N_20468,N_16718,N_16600);
and U20469 (N_20469,N_18436,N_16232);
nor U20470 (N_20470,N_16429,N_17707);
nand U20471 (N_20471,N_17870,N_18548);
xnor U20472 (N_20472,N_18182,N_17741);
nor U20473 (N_20473,N_18416,N_15717);
and U20474 (N_20474,N_18551,N_17811);
nand U20475 (N_20475,N_16746,N_17335);
xor U20476 (N_20476,N_16628,N_17772);
nand U20477 (N_20477,N_15678,N_18502);
or U20478 (N_20478,N_16934,N_17475);
and U20479 (N_20479,N_17982,N_16317);
nor U20480 (N_20480,N_18737,N_15792);
and U20481 (N_20481,N_18434,N_15722);
or U20482 (N_20482,N_17169,N_15861);
xnor U20483 (N_20483,N_18098,N_17185);
or U20484 (N_20484,N_17552,N_15812);
or U20485 (N_20485,N_17750,N_18218);
nand U20486 (N_20486,N_17737,N_17098);
and U20487 (N_20487,N_16480,N_16139);
nand U20488 (N_20488,N_16192,N_17336);
nand U20489 (N_20489,N_18027,N_15930);
nand U20490 (N_20490,N_18187,N_18158);
and U20491 (N_20491,N_17173,N_18290);
nand U20492 (N_20492,N_16747,N_16404);
or U20493 (N_20493,N_17012,N_17317);
and U20494 (N_20494,N_16335,N_17363);
and U20495 (N_20495,N_17424,N_18311);
xnor U20496 (N_20496,N_18216,N_17316);
nand U20497 (N_20497,N_18315,N_16024);
or U20498 (N_20498,N_17762,N_16459);
nor U20499 (N_20499,N_16276,N_15853);
nand U20500 (N_20500,N_18432,N_17178);
nor U20501 (N_20501,N_18500,N_16510);
or U20502 (N_20502,N_15967,N_16178);
nor U20503 (N_20503,N_15879,N_17287);
nor U20504 (N_20504,N_17733,N_16638);
and U20505 (N_20505,N_16161,N_16417);
and U20506 (N_20506,N_16657,N_15782);
or U20507 (N_20507,N_18447,N_18516);
nand U20508 (N_20508,N_18580,N_15921);
nor U20509 (N_20509,N_15828,N_16735);
nor U20510 (N_20510,N_16436,N_16275);
and U20511 (N_20511,N_16790,N_18304);
xor U20512 (N_20512,N_17396,N_17613);
nor U20513 (N_20513,N_18490,N_16130);
nand U20514 (N_20514,N_16907,N_18317);
and U20515 (N_20515,N_17793,N_16660);
xor U20516 (N_20516,N_17118,N_18035);
nand U20517 (N_20517,N_16100,N_16562);
or U20518 (N_20518,N_15638,N_16459);
or U20519 (N_20519,N_16920,N_18586);
nor U20520 (N_20520,N_17035,N_18124);
nor U20521 (N_20521,N_17634,N_17474);
nand U20522 (N_20522,N_17896,N_16391);
nor U20523 (N_20523,N_17193,N_17574);
xor U20524 (N_20524,N_15692,N_15966);
nor U20525 (N_20525,N_15662,N_17043);
or U20526 (N_20526,N_16077,N_16423);
and U20527 (N_20527,N_16329,N_15880);
nand U20528 (N_20528,N_17033,N_16423);
and U20529 (N_20529,N_17985,N_17507);
and U20530 (N_20530,N_17138,N_17432);
and U20531 (N_20531,N_16753,N_18324);
xnor U20532 (N_20532,N_16569,N_15854);
or U20533 (N_20533,N_18442,N_16759);
and U20534 (N_20534,N_17170,N_15659);
and U20535 (N_20535,N_16522,N_18299);
nand U20536 (N_20536,N_18496,N_15803);
or U20537 (N_20537,N_17367,N_18654);
and U20538 (N_20538,N_16228,N_18464);
nand U20539 (N_20539,N_17700,N_17819);
nand U20540 (N_20540,N_17700,N_16144);
nand U20541 (N_20541,N_17910,N_16287);
nand U20542 (N_20542,N_17464,N_15691);
nor U20543 (N_20543,N_18130,N_18737);
or U20544 (N_20544,N_18000,N_17616);
nor U20545 (N_20545,N_17984,N_16767);
or U20546 (N_20546,N_15856,N_17744);
and U20547 (N_20547,N_17862,N_18454);
nand U20548 (N_20548,N_15644,N_18017);
and U20549 (N_20549,N_16389,N_15774);
xnor U20550 (N_20550,N_17910,N_18512);
or U20551 (N_20551,N_18740,N_18672);
or U20552 (N_20552,N_17984,N_18638);
and U20553 (N_20553,N_17815,N_16250);
and U20554 (N_20554,N_17565,N_17330);
nand U20555 (N_20555,N_15954,N_15994);
nor U20556 (N_20556,N_17463,N_15852);
or U20557 (N_20557,N_15853,N_15729);
xnor U20558 (N_20558,N_18620,N_16761);
nand U20559 (N_20559,N_15987,N_16553);
nor U20560 (N_20560,N_18298,N_17690);
and U20561 (N_20561,N_17251,N_17275);
and U20562 (N_20562,N_16535,N_18608);
or U20563 (N_20563,N_17129,N_17300);
or U20564 (N_20564,N_16396,N_17369);
or U20565 (N_20565,N_15909,N_16318);
xnor U20566 (N_20566,N_18568,N_18408);
nor U20567 (N_20567,N_17071,N_17898);
xor U20568 (N_20568,N_18457,N_18052);
nand U20569 (N_20569,N_18564,N_18215);
nand U20570 (N_20570,N_15816,N_15891);
nand U20571 (N_20571,N_18125,N_17114);
xnor U20572 (N_20572,N_17766,N_16884);
nor U20573 (N_20573,N_16274,N_17515);
nand U20574 (N_20574,N_17471,N_17238);
or U20575 (N_20575,N_18252,N_16306);
or U20576 (N_20576,N_18535,N_16394);
nor U20577 (N_20577,N_17908,N_17889);
xor U20578 (N_20578,N_17619,N_16577);
xnor U20579 (N_20579,N_17873,N_16797);
xnor U20580 (N_20580,N_18285,N_16585);
nor U20581 (N_20581,N_17304,N_16067);
and U20582 (N_20582,N_17113,N_18556);
or U20583 (N_20583,N_16743,N_16060);
nor U20584 (N_20584,N_17995,N_16425);
nor U20585 (N_20585,N_17060,N_18525);
nor U20586 (N_20586,N_18341,N_18266);
and U20587 (N_20587,N_18527,N_16114);
xor U20588 (N_20588,N_18473,N_17244);
nand U20589 (N_20589,N_17211,N_16529);
and U20590 (N_20590,N_17111,N_17680);
nand U20591 (N_20591,N_17414,N_18364);
nand U20592 (N_20592,N_17310,N_16367);
and U20593 (N_20593,N_17027,N_16146);
and U20594 (N_20594,N_15660,N_17444);
or U20595 (N_20595,N_18679,N_17180);
or U20596 (N_20596,N_18610,N_18351);
or U20597 (N_20597,N_18696,N_17059);
or U20598 (N_20598,N_18571,N_17417);
and U20599 (N_20599,N_18238,N_17407);
nand U20600 (N_20600,N_15775,N_17741);
nand U20601 (N_20601,N_15913,N_17484);
nor U20602 (N_20602,N_15796,N_15862);
nor U20603 (N_20603,N_16342,N_17180);
or U20604 (N_20604,N_15697,N_17601);
or U20605 (N_20605,N_18239,N_17823);
or U20606 (N_20606,N_17408,N_18599);
nor U20607 (N_20607,N_17966,N_16832);
nor U20608 (N_20608,N_15888,N_17373);
nand U20609 (N_20609,N_17178,N_17003);
xor U20610 (N_20610,N_16588,N_16557);
nor U20611 (N_20611,N_17068,N_16190);
nor U20612 (N_20612,N_16925,N_18630);
nor U20613 (N_20613,N_16160,N_18418);
nand U20614 (N_20614,N_17543,N_17903);
xor U20615 (N_20615,N_17633,N_17010);
or U20616 (N_20616,N_16546,N_15747);
and U20617 (N_20617,N_17652,N_16025);
nand U20618 (N_20618,N_17288,N_17953);
nand U20619 (N_20619,N_16989,N_16911);
or U20620 (N_20620,N_17016,N_17603);
or U20621 (N_20621,N_15822,N_18149);
nand U20622 (N_20622,N_17936,N_17393);
and U20623 (N_20623,N_16889,N_17469);
or U20624 (N_20624,N_15832,N_18400);
and U20625 (N_20625,N_17831,N_18681);
or U20626 (N_20626,N_18646,N_17184);
or U20627 (N_20627,N_17979,N_16415);
nor U20628 (N_20628,N_16714,N_17458);
nand U20629 (N_20629,N_17802,N_17411);
or U20630 (N_20630,N_16019,N_15704);
or U20631 (N_20631,N_17635,N_18076);
nand U20632 (N_20632,N_16064,N_16256);
or U20633 (N_20633,N_17206,N_16021);
or U20634 (N_20634,N_17824,N_15876);
or U20635 (N_20635,N_17253,N_16742);
xnor U20636 (N_20636,N_16936,N_17663);
xnor U20637 (N_20637,N_17841,N_17917);
nor U20638 (N_20638,N_17001,N_17676);
nor U20639 (N_20639,N_18532,N_17594);
nor U20640 (N_20640,N_16078,N_18059);
and U20641 (N_20641,N_18257,N_17635);
nand U20642 (N_20642,N_17055,N_16089);
and U20643 (N_20643,N_18321,N_16127);
nand U20644 (N_20644,N_15981,N_17770);
nand U20645 (N_20645,N_15952,N_15961);
xnor U20646 (N_20646,N_15938,N_18052);
nor U20647 (N_20647,N_16807,N_17710);
nor U20648 (N_20648,N_18093,N_18609);
nand U20649 (N_20649,N_17117,N_17513);
and U20650 (N_20650,N_16601,N_16690);
and U20651 (N_20651,N_18619,N_17745);
xor U20652 (N_20652,N_17448,N_15798);
nand U20653 (N_20653,N_17652,N_18450);
and U20654 (N_20654,N_16513,N_17693);
nor U20655 (N_20655,N_16886,N_18149);
nor U20656 (N_20656,N_17245,N_18484);
xor U20657 (N_20657,N_18209,N_16102);
and U20658 (N_20658,N_15927,N_18361);
nand U20659 (N_20659,N_18229,N_17315);
nor U20660 (N_20660,N_15958,N_17853);
or U20661 (N_20661,N_18432,N_17345);
or U20662 (N_20662,N_17022,N_17297);
or U20663 (N_20663,N_16467,N_17144);
xor U20664 (N_20664,N_16505,N_17694);
nand U20665 (N_20665,N_16187,N_16287);
xnor U20666 (N_20666,N_18411,N_17693);
and U20667 (N_20667,N_16164,N_15733);
nor U20668 (N_20668,N_16737,N_17425);
nor U20669 (N_20669,N_15859,N_16826);
nor U20670 (N_20670,N_18430,N_16522);
nor U20671 (N_20671,N_17025,N_18338);
and U20672 (N_20672,N_15845,N_16572);
nor U20673 (N_20673,N_18176,N_16339);
or U20674 (N_20674,N_16640,N_16955);
xor U20675 (N_20675,N_17156,N_17050);
or U20676 (N_20676,N_17757,N_17634);
nand U20677 (N_20677,N_18257,N_17562);
xnor U20678 (N_20678,N_17479,N_17527);
nor U20679 (N_20679,N_18345,N_17862);
nor U20680 (N_20680,N_17408,N_16752);
nor U20681 (N_20681,N_17398,N_16590);
nand U20682 (N_20682,N_15848,N_16012);
and U20683 (N_20683,N_18725,N_15882);
or U20684 (N_20684,N_16443,N_17686);
nand U20685 (N_20685,N_17906,N_18456);
and U20686 (N_20686,N_18360,N_18006);
or U20687 (N_20687,N_17662,N_16786);
xnor U20688 (N_20688,N_18715,N_16542);
nand U20689 (N_20689,N_16402,N_18060);
and U20690 (N_20690,N_18149,N_18155);
nand U20691 (N_20691,N_16047,N_16088);
nor U20692 (N_20692,N_17212,N_18028);
nor U20693 (N_20693,N_18076,N_16189);
and U20694 (N_20694,N_17974,N_17688);
nand U20695 (N_20695,N_18292,N_18012);
or U20696 (N_20696,N_16317,N_17786);
nor U20697 (N_20697,N_17965,N_17299);
nand U20698 (N_20698,N_17388,N_16240);
and U20699 (N_20699,N_18557,N_18417);
and U20700 (N_20700,N_15714,N_18683);
nor U20701 (N_20701,N_18733,N_15697);
nand U20702 (N_20702,N_18733,N_15898);
or U20703 (N_20703,N_18101,N_17236);
nand U20704 (N_20704,N_16512,N_16528);
xor U20705 (N_20705,N_16429,N_17422);
and U20706 (N_20706,N_16741,N_18721);
or U20707 (N_20707,N_16805,N_16874);
xnor U20708 (N_20708,N_17607,N_16185);
nand U20709 (N_20709,N_17492,N_16184);
or U20710 (N_20710,N_18075,N_16502);
nand U20711 (N_20711,N_16301,N_17500);
nor U20712 (N_20712,N_16255,N_17658);
nor U20713 (N_20713,N_16579,N_17204);
nor U20714 (N_20714,N_16343,N_17604);
or U20715 (N_20715,N_16118,N_18251);
nor U20716 (N_20716,N_17284,N_16893);
and U20717 (N_20717,N_16784,N_18506);
nor U20718 (N_20718,N_18423,N_18468);
nand U20719 (N_20719,N_17519,N_15883);
or U20720 (N_20720,N_18723,N_17801);
or U20721 (N_20721,N_17114,N_17656);
and U20722 (N_20722,N_16786,N_15936);
nand U20723 (N_20723,N_18492,N_18590);
xnor U20724 (N_20724,N_17645,N_18414);
or U20725 (N_20725,N_17410,N_15910);
or U20726 (N_20726,N_17674,N_18403);
and U20727 (N_20727,N_15946,N_16175);
nor U20728 (N_20728,N_18068,N_16733);
xor U20729 (N_20729,N_17849,N_18089);
and U20730 (N_20730,N_16953,N_17968);
xnor U20731 (N_20731,N_17126,N_15675);
nand U20732 (N_20732,N_17225,N_16085);
nand U20733 (N_20733,N_18534,N_17985);
nor U20734 (N_20734,N_18076,N_17869);
or U20735 (N_20735,N_17897,N_18113);
nor U20736 (N_20736,N_17585,N_17751);
nand U20737 (N_20737,N_16978,N_17730);
nor U20738 (N_20738,N_16000,N_16859);
and U20739 (N_20739,N_16077,N_18079);
nor U20740 (N_20740,N_17819,N_15812);
and U20741 (N_20741,N_18187,N_16887);
nand U20742 (N_20742,N_17156,N_16831);
and U20743 (N_20743,N_16446,N_18412);
nand U20744 (N_20744,N_16562,N_17756);
and U20745 (N_20745,N_17626,N_18227);
or U20746 (N_20746,N_18383,N_17583);
and U20747 (N_20747,N_18230,N_17497);
nand U20748 (N_20748,N_17888,N_18115);
or U20749 (N_20749,N_16706,N_16505);
or U20750 (N_20750,N_16812,N_17692);
nor U20751 (N_20751,N_16651,N_17972);
nor U20752 (N_20752,N_17181,N_17977);
nand U20753 (N_20753,N_17705,N_16215);
and U20754 (N_20754,N_15754,N_17486);
nand U20755 (N_20755,N_18245,N_17081);
or U20756 (N_20756,N_16156,N_17665);
nand U20757 (N_20757,N_16687,N_18258);
and U20758 (N_20758,N_18202,N_18240);
nor U20759 (N_20759,N_15868,N_17787);
xnor U20760 (N_20760,N_15727,N_16445);
and U20761 (N_20761,N_18595,N_17173);
nor U20762 (N_20762,N_18039,N_17039);
nand U20763 (N_20763,N_18565,N_16808);
and U20764 (N_20764,N_17799,N_17981);
and U20765 (N_20765,N_18080,N_17609);
or U20766 (N_20766,N_18151,N_16886);
and U20767 (N_20767,N_16505,N_16871);
nand U20768 (N_20768,N_16476,N_18403);
xor U20769 (N_20769,N_17337,N_16572);
or U20770 (N_20770,N_17046,N_18341);
nor U20771 (N_20771,N_17990,N_17306);
or U20772 (N_20772,N_17843,N_17556);
and U20773 (N_20773,N_17588,N_17140);
or U20774 (N_20774,N_18636,N_15711);
nor U20775 (N_20775,N_18203,N_16171);
and U20776 (N_20776,N_15712,N_16733);
nor U20777 (N_20777,N_18542,N_16016);
nor U20778 (N_20778,N_15771,N_15826);
nand U20779 (N_20779,N_18603,N_17845);
nand U20780 (N_20780,N_15761,N_16943);
or U20781 (N_20781,N_17510,N_15643);
nor U20782 (N_20782,N_16784,N_17838);
nor U20783 (N_20783,N_15968,N_16254);
xor U20784 (N_20784,N_18488,N_16232);
and U20785 (N_20785,N_16917,N_16779);
xnor U20786 (N_20786,N_18467,N_17778);
nand U20787 (N_20787,N_18274,N_18404);
nor U20788 (N_20788,N_16864,N_15949);
and U20789 (N_20789,N_17352,N_16899);
nand U20790 (N_20790,N_16932,N_18733);
xor U20791 (N_20791,N_18476,N_16971);
or U20792 (N_20792,N_18078,N_17764);
and U20793 (N_20793,N_17646,N_17537);
and U20794 (N_20794,N_17154,N_16081);
nand U20795 (N_20795,N_16948,N_18498);
xor U20796 (N_20796,N_17313,N_17708);
nand U20797 (N_20797,N_16946,N_17378);
nor U20798 (N_20798,N_17424,N_16075);
or U20799 (N_20799,N_17773,N_18491);
nor U20800 (N_20800,N_16866,N_17704);
nand U20801 (N_20801,N_16028,N_17889);
nor U20802 (N_20802,N_16952,N_15942);
and U20803 (N_20803,N_18219,N_17562);
nand U20804 (N_20804,N_17802,N_16912);
and U20805 (N_20805,N_15911,N_15802);
and U20806 (N_20806,N_17966,N_16795);
or U20807 (N_20807,N_15827,N_18327);
and U20808 (N_20808,N_18412,N_17626);
nor U20809 (N_20809,N_17007,N_16734);
nor U20810 (N_20810,N_15697,N_17061);
xnor U20811 (N_20811,N_18674,N_18460);
nor U20812 (N_20812,N_18519,N_17822);
nand U20813 (N_20813,N_18092,N_16284);
and U20814 (N_20814,N_16513,N_16794);
nand U20815 (N_20815,N_16616,N_17572);
nor U20816 (N_20816,N_17673,N_17886);
and U20817 (N_20817,N_18296,N_16128);
or U20818 (N_20818,N_16247,N_17858);
or U20819 (N_20819,N_15711,N_16217);
and U20820 (N_20820,N_17378,N_17849);
nand U20821 (N_20821,N_17243,N_15868);
or U20822 (N_20822,N_17887,N_16875);
nand U20823 (N_20823,N_16414,N_17721);
and U20824 (N_20824,N_16365,N_16829);
xnor U20825 (N_20825,N_17361,N_17069);
xor U20826 (N_20826,N_17988,N_17636);
and U20827 (N_20827,N_16838,N_16636);
xnor U20828 (N_20828,N_16642,N_17795);
or U20829 (N_20829,N_15716,N_16844);
or U20830 (N_20830,N_18000,N_16505);
or U20831 (N_20831,N_16198,N_17612);
nand U20832 (N_20832,N_18612,N_18400);
nor U20833 (N_20833,N_18588,N_18681);
xor U20834 (N_20834,N_16398,N_15685);
nand U20835 (N_20835,N_17386,N_15956);
xnor U20836 (N_20836,N_16739,N_18724);
or U20837 (N_20837,N_16754,N_16827);
nor U20838 (N_20838,N_18048,N_17102);
nand U20839 (N_20839,N_16869,N_18345);
nand U20840 (N_20840,N_18041,N_17464);
and U20841 (N_20841,N_17668,N_16003);
and U20842 (N_20842,N_17539,N_17552);
xor U20843 (N_20843,N_18282,N_16613);
nor U20844 (N_20844,N_18240,N_17807);
nand U20845 (N_20845,N_17882,N_16026);
and U20846 (N_20846,N_17056,N_16200);
and U20847 (N_20847,N_18336,N_17740);
nand U20848 (N_20848,N_16628,N_16265);
nor U20849 (N_20849,N_18540,N_16644);
nor U20850 (N_20850,N_17208,N_16003);
nor U20851 (N_20851,N_16328,N_16330);
nand U20852 (N_20852,N_16083,N_18555);
or U20853 (N_20853,N_17846,N_18217);
nor U20854 (N_20854,N_16081,N_17862);
and U20855 (N_20855,N_16058,N_17666);
or U20856 (N_20856,N_17215,N_18151);
and U20857 (N_20857,N_18563,N_16591);
nand U20858 (N_20858,N_18655,N_17047);
nor U20859 (N_20859,N_16537,N_17049);
nor U20860 (N_20860,N_18552,N_15883);
xor U20861 (N_20861,N_18304,N_16913);
and U20862 (N_20862,N_15669,N_15854);
nor U20863 (N_20863,N_17344,N_16840);
xnor U20864 (N_20864,N_16057,N_16375);
nor U20865 (N_20865,N_16948,N_18159);
nor U20866 (N_20866,N_15861,N_17042);
and U20867 (N_20867,N_18217,N_16498);
nor U20868 (N_20868,N_17800,N_15782);
xnor U20869 (N_20869,N_18718,N_17518);
or U20870 (N_20870,N_17114,N_17486);
and U20871 (N_20871,N_18571,N_17251);
nand U20872 (N_20872,N_16708,N_16319);
nor U20873 (N_20873,N_18000,N_16948);
and U20874 (N_20874,N_18257,N_17510);
nor U20875 (N_20875,N_18457,N_16618);
or U20876 (N_20876,N_16782,N_17073);
nor U20877 (N_20877,N_18035,N_16911);
or U20878 (N_20878,N_17362,N_18137);
xor U20879 (N_20879,N_16340,N_18109);
nor U20880 (N_20880,N_18168,N_18338);
or U20881 (N_20881,N_16352,N_17727);
nand U20882 (N_20882,N_17646,N_17164);
and U20883 (N_20883,N_17775,N_16119);
or U20884 (N_20884,N_17719,N_16482);
nand U20885 (N_20885,N_17073,N_15850);
and U20886 (N_20886,N_17132,N_16137);
and U20887 (N_20887,N_16482,N_16039);
nor U20888 (N_20888,N_16655,N_18596);
or U20889 (N_20889,N_16522,N_18171);
and U20890 (N_20890,N_17758,N_17309);
nor U20891 (N_20891,N_16676,N_16352);
nand U20892 (N_20892,N_15850,N_18092);
nand U20893 (N_20893,N_16355,N_16555);
nand U20894 (N_20894,N_16983,N_16592);
nor U20895 (N_20895,N_17012,N_17864);
nand U20896 (N_20896,N_18485,N_17468);
xor U20897 (N_20897,N_15760,N_15666);
and U20898 (N_20898,N_16433,N_18072);
or U20899 (N_20899,N_18693,N_16377);
nor U20900 (N_20900,N_18411,N_18748);
nand U20901 (N_20901,N_17823,N_17005);
or U20902 (N_20902,N_17017,N_17182);
xnor U20903 (N_20903,N_16236,N_16827);
nor U20904 (N_20904,N_18101,N_16792);
nand U20905 (N_20905,N_16120,N_17907);
or U20906 (N_20906,N_16808,N_15703);
xnor U20907 (N_20907,N_16529,N_16340);
or U20908 (N_20908,N_15707,N_15869);
or U20909 (N_20909,N_18264,N_18250);
and U20910 (N_20910,N_16956,N_17866);
and U20911 (N_20911,N_17212,N_16102);
nor U20912 (N_20912,N_17183,N_18714);
nand U20913 (N_20913,N_16737,N_16845);
or U20914 (N_20914,N_15910,N_18696);
or U20915 (N_20915,N_16243,N_18031);
xnor U20916 (N_20916,N_18402,N_16051);
or U20917 (N_20917,N_16196,N_16809);
and U20918 (N_20918,N_16330,N_15945);
and U20919 (N_20919,N_17096,N_16402);
or U20920 (N_20920,N_17222,N_17662);
nand U20921 (N_20921,N_18734,N_16713);
and U20922 (N_20922,N_17215,N_16744);
nand U20923 (N_20923,N_15996,N_18554);
or U20924 (N_20924,N_16244,N_17982);
xnor U20925 (N_20925,N_17440,N_18009);
and U20926 (N_20926,N_18699,N_17491);
xnor U20927 (N_20927,N_16521,N_18174);
nor U20928 (N_20928,N_16494,N_17061);
or U20929 (N_20929,N_17035,N_16904);
or U20930 (N_20930,N_17541,N_17523);
or U20931 (N_20931,N_16647,N_18281);
nor U20932 (N_20932,N_15875,N_17370);
nand U20933 (N_20933,N_17652,N_18396);
or U20934 (N_20934,N_16082,N_17404);
or U20935 (N_20935,N_17449,N_16506);
nand U20936 (N_20936,N_17090,N_16064);
and U20937 (N_20937,N_15854,N_17860);
xor U20938 (N_20938,N_16229,N_17121);
and U20939 (N_20939,N_18361,N_18735);
nand U20940 (N_20940,N_15904,N_16555);
or U20941 (N_20941,N_17428,N_17166);
nand U20942 (N_20942,N_17241,N_18337);
nor U20943 (N_20943,N_15829,N_16102);
nand U20944 (N_20944,N_17455,N_16652);
nand U20945 (N_20945,N_18730,N_15787);
nand U20946 (N_20946,N_16560,N_18673);
nor U20947 (N_20947,N_17955,N_15820);
and U20948 (N_20948,N_16383,N_16385);
nor U20949 (N_20949,N_17054,N_16290);
and U20950 (N_20950,N_18398,N_16862);
and U20951 (N_20951,N_16730,N_15714);
or U20952 (N_20952,N_16145,N_17921);
xor U20953 (N_20953,N_17701,N_17002);
nand U20954 (N_20954,N_18690,N_18536);
or U20955 (N_20955,N_16159,N_18705);
nand U20956 (N_20956,N_16293,N_17405);
nor U20957 (N_20957,N_18403,N_18274);
and U20958 (N_20958,N_15675,N_18657);
or U20959 (N_20959,N_15951,N_16725);
xnor U20960 (N_20960,N_16514,N_18599);
nand U20961 (N_20961,N_17411,N_16078);
or U20962 (N_20962,N_15884,N_17847);
nand U20963 (N_20963,N_17544,N_16999);
nor U20964 (N_20964,N_18214,N_16462);
and U20965 (N_20965,N_16274,N_16402);
nor U20966 (N_20966,N_17853,N_17052);
nand U20967 (N_20967,N_17513,N_18558);
nor U20968 (N_20968,N_16763,N_16413);
nand U20969 (N_20969,N_15753,N_15718);
or U20970 (N_20970,N_16516,N_17050);
or U20971 (N_20971,N_16881,N_16817);
or U20972 (N_20972,N_18304,N_17802);
nand U20973 (N_20973,N_18361,N_16216);
xor U20974 (N_20974,N_17958,N_16444);
nand U20975 (N_20975,N_16768,N_16623);
xor U20976 (N_20976,N_17488,N_18131);
and U20977 (N_20977,N_15739,N_18236);
or U20978 (N_20978,N_16142,N_17298);
and U20979 (N_20979,N_16171,N_15848);
and U20980 (N_20980,N_17472,N_16301);
nor U20981 (N_20981,N_16713,N_15732);
and U20982 (N_20982,N_17719,N_18074);
or U20983 (N_20983,N_18389,N_16248);
or U20984 (N_20984,N_16318,N_17932);
or U20985 (N_20985,N_17385,N_18048);
and U20986 (N_20986,N_17898,N_16738);
and U20987 (N_20987,N_17850,N_17358);
or U20988 (N_20988,N_16763,N_18621);
or U20989 (N_20989,N_18691,N_16653);
nand U20990 (N_20990,N_16453,N_18467);
nor U20991 (N_20991,N_16729,N_16596);
nand U20992 (N_20992,N_16746,N_17469);
nor U20993 (N_20993,N_18520,N_16503);
or U20994 (N_20994,N_18479,N_16535);
xor U20995 (N_20995,N_17829,N_17854);
nand U20996 (N_20996,N_16747,N_17345);
nor U20997 (N_20997,N_15651,N_16639);
nand U20998 (N_20998,N_16568,N_16130);
nand U20999 (N_20999,N_15944,N_17687);
nor U21000 (N_21000,N_17946,N_16156);
xnor U21001 (N_21001,N_18520,N_15677);
nand U21002 (N_21002,N_15982,N_18712);
nand U21003 (N_21003,N_15843,N_16004);
and U21004 (N_21004,N_17086,N_15971);
or U21005 (N_21005,N_16202,N_17355);
and U21006 (N_21006,N_16490,N_16789);
nand U21007 (N_21007,N_18303,N_16051);
nor U21008 (N_21008,N_17575,N_15897);
nor U21009 (N_21009,N_17329,N_18735);
and U21010 (N_21010,N_16544,N_16336);
nor U21011 (N_21011,N_18692,N_16900);
nor U21012 (N_21012,N_16031,N_18515);
or U21013 (N_21013,N_18006,N_17525);
nand U21014 (N_21014,N_18335,N_18704);
and U21015 (N_21015,N_18395,N_18412);
and U21016 (N_21016,N_17988,N_17904);
or U21017 (N_21017,N_18248,N_16686);
nor U21018 (N_21018,N_18571,N_16742);
and U21019 (N_21019,N_17017,N_15776);
or U21020 (N_21020,N_15752,N_18004);
and U21021 (N_21021,N_15942,N_16010);
xor U21022 (N_21022,N_17773,N_17854);
nor U21023 (N_21023,N_18435,N_18422);
nand U21024 (N_21024,N_16874,N_18492);
or U21025 (N_21025,N_16998,N_16715);
nor U21026 (N_21026,N_16338,N_17981);
nor U21027 (N_21027,N_17501,N_16149);
nor U21028 (N_21028,N_18420,N_15766);
nand U21029 (N_21029,N_16415,N_18103);
xnor U21030 (N_21030,N_17129,N_17426);
or U21031 (N_21031,N_15721,N_15895);
or U21032 (N_21032,N_16474,N_18297);
nand U21033 (N_21033,N_16251,N_17473);
nor U21034 (N_21034,N_17362,N_17157);
and U21035 (N_21035,N_18243,N_16300);
nand U21036 (N_21036,N_16506,N_16709);
nand U21037 (N_21037,N_17852,N_16812);
nand U21038 (N_21038,N_17769,N_17293);
xor U21039 (N_21039,N_18404,N_17381);
xnor U21040 (N_21040,N_18563,N_15703);
and U21041 (N_21041,N_15907,N_18305);
nand U21042 (N_21042,N_16428,N_16004);
nand U21043 (N_21043,N_15862,N_17051);
and U21044 (N_21044,N_17261,N_17610);
or U21045 (N_21045,N_17727,N_16007);
nor U21046 (N_21046,N_16939,N_16393);
and U21047 (N_21047,N_15886,N_16591);
and U21048 (N_21048,N_17566,N_18482);
nor U21049 (N_21049,N_17700,N_16100);
and U21050 (N_21050,N_17384,N_16898);
nor U21051 (N_21051,N_18434,N_17294);
and U21052 (N_21052,N_17282,N_16002);
nor U21053 (N_21053,N_16490,N_15864);
nand U21054 (N_21054,N_17397,N_18135);
nor U21055 (N_21055,N_18650,N_18246);
nor U21056 (N_21056,N_15758,N_18615);
and U21057 (N_21057,N_17048,N_16256);
and U21058 (N_21058,N_16785,N_15959);
and U21059 (N_21059,N_16558,N_16259);
xnor U21060 (N_21060,N_15745,N_18645);
and U21061 (N_21061,N_17986,N_15839);
xnor U21062 (N_21062,N_16098,N_17363);
or U21063 (N_21063,N_16793,N_17909);
or U21064 (N_21064,N_16911,N_18510);
nor U21065 (N_21065,N_17946,N_16230);
nand U21066 (N_21066,N_17500,N_15816);
or U21067 (N_21067,N_16874,N_16942);
nor U21068 (N_21068,N_15818,N_16957);
and U21069 (N_21069,N_17065,N_17759);
nor U21070 (N_21070,N_18688,N_15659);
or U21071 (N_21071,N_16868,N_15900);
and U21072 (N_21072,N_16130,N_16763);
nand U21073 (N_21073,N_17284,N_16469);
nor U21074 (N_21074,N_17803,N_17135);
nor U21075 (N_21075,N_16857,N_16722);
and U21076 (N_21076,N_18550,N_15963);
or U21077 (N_21077,N_16654,N_16272);
nor U21078 (N_21078,N_17722,N_18745);
xnor U21079 (N_21079,N_16636,N_18718);
nand U21080 (N_21080,N_16761,N_16426);
and U21081 (N_21081,N_16806,N_18392);
or U21082 (N_21082,N_18172,N_16649);
and U21083 (N_21083,N_17182,N_18008);
and U21084 (N_21084,N_16968,N_18434);
or U21085 (N_21085,N_17621,N_17844);
nand U21086 (N_21086,N_16164,N_17009);
nor U21087 (N_21087,N_16817,N_17946);
and U21088 (N_21088,N_16209,N_17546);
and U21089 (N_21089,N_18271,N_18238);
and U21090 (N_21090,N_16603,N_17588);
or U21091 (N_21091,N_16755,N_18392);
or U21092 (N_21092,N_17897,N_17704);
nor U21093 (N_21093,N_16826,N_16698);
and U21094 (N_21094,N_17812,N_15736);
xor U21095 (N_21095,N_17454,N_17731);
and U21096 (N_21096,N_18081,N_16063);
or U21097 (N_21097,N_17424,N_17569);
nor U21098 (N_21098,N_15718,N_17629);
or U21099 (N_21099,N_18457,N_15849);
nor U21100 (N_21100,N_18049,N_16828);
nand U21101 (N_21101,N_17563,N_17890);
or U21102 (N_21102,N_17214,N_18570);
and U21103 (N_21103,N_16200,N_16241);
and U21104 (N_21104,N_16649,N_16878);
nand U21105 (N_21105,N_15787,N_15941);
nor U21106 (N_21106,N_16445,N_17442);
nand U21107 (N_21107,N_15637,N_17119);
and U21108 (N_21108,N_15977,N_18656);
nand U21109 (N_21109,N_18640,N_16332);
nand U21110 (N_21110,N_16604,N_17943);
or U21111 (N_21111,N_15873,N_18043);
or U21112 (N_21112,N_17711,N_17919);
and U21113 (N_21113,N_15817,N_18022);
nand U21114 (N_21114,N_17874,N_18052);
nor U21115 (N_21115,N_15931,N_16105);
nor U21116 (N_21116,N_16532,N_15827);
nand U21117 (N_21117,N_17056,N_18672);
nor U21118 (N_21118,N_18028,N_17817);
or U21119 (N_21119,N_18011,N_17390);
xor U21120 (N_21120,N_16780,N_15629);
nand U21121 (N_21121,N_16264,N_16780);
and U21122 (N_21122,N_18172,N_18390);
or U21123 (N_21123,N_17677,N_15635);
nand U21124 (N_21124,N_18699,N_18576);
and U21125 (N_21125,N_17584,N_16605);
or U21126 (N_21126,N_18511,N_18403);
nor U21127 (N_21127,N_16336,N_15813);
and U21128 (N_21128,N_15800,N_16911);
nor U21129 (N_21129,N_18160,N_15972);
and U21130 (N_21130,N_18433,N_17168);
and U21131 (N_21131,N_15697,N_18618);
and U21132 (N_21132,N_18093,N_16057);
nand U21133 (N_21133,N_17021,N_16217);
nor U21134 (N_21134,N_17302,N_18074);
nand U21135 (N_21135,N_15944,N_18139);
and U21136 (N_21136,N_17081,N_16994);
xnor U21137 (N_21137,N_15659,N_18350);
nand U21138 (N_21138,N_17570,N_16755);
or U21139 (N_21139,N_16417,N_15862);
or U21140 (N_21140,N_17142,N_17050);
and U21141 (N_21141,N_16126,N_16224);
or U21142 (N_21142,N_16508,N_16133);
nand U21143 (N_21143,N_18121,N_18313);
nor U21144 (N_21144,N_18037,N_18697);
or U21145 (N_21145,N_18442,N_18121);
and U21146 (N_21146,N_16539,N_17203);
nor U21147 (N_21147,N_17947,N_18213);
xor U21148 (N_21148,N_16727,N_15639);
or U21149 (N_21149,N_15633,N_18554);
nor U21150 (N_21150,N_16193,N_16646);
nor U21151 (N_21151,N_16517,N_15933);
and U21152 (N_21152,N_16076,N_17160);
and U21153 (N_21153,N_15724,N_17446);
nand U21154 (N_21154,N_16776,N_17252);
or U21155 (N_21155,N_18649,N_16821);
or U21156 (N_21156,N_17687,N_17730);
or U21157 (N_21157,N_16179,N_16814);
nor U21158 (N_21158,N_17352,N_17879);
xnor U21159 (N_21159,N_15739,N_17882);
or U21160 (N_21160,N_17957,N_17885);
or U21161 (N_21161,N_17578,N_16614);
nand U21162 (N_21162,N_18273,N_18611);
and U21163 (N_21163,N_18628,N_17824);
or U21164 (N_21164,N_17432,N_18507);
nand U21165 (N_21165,N_16021,N_16119);
or U21166 (N_21166,N_16525,N_17923);
and U21167 (N_21167,N_18725,N_17708);
or U21168 (N_21168,N_17705,N_18248);
nand U21169 (N_21169,N_17773,N_17409);
nor U21170 (N_21170,N_16620,N_17598);
or U21171 (N_21171,N_17198,N_16252);
and U21172 (N_21172,N_18306,N_17498);
and U21173 (N_21173,N_16833,N_18188);
nor U21174 (N_21174,N_15741,N_18477);
nor U21175 (N_21175,N_16078,N_16698);
and U21176 (N_21176,N_18352,N_17717);
and U21177 (N_21177,N_15844,N_16537);
and U21178 (N_21178,N_17670,N_15734);
and U21179 (N_21179,N_17811,N_16882);
xnor U21180 (N_21180,N_18602,N_17407);
and U21181 (N_21181,N_15686,N_18537);
and U21182 (N_21182,N_17193,N_16291);
and U21183 (N_21183,N_18138,N_15911);
nor U21184 (N_21184,N_18624,N_18715);
nand U21185 (N_21185,N_16328,N_17600);
or U21186 (N_21186,N_16379,N_17429);
and U21187 (N_21187,N_15964,N_15776);
nand U21188 (N_21188,N_17079,N_16952);
or U21189 (N_21189,N_15677,N_18145);
or U21190 (N_21190,N_15928,N_18113);
nand U21191 (N_21191,N_16584,N_18661);
nor U21192 (N_21192,N_18663,N_16399);
xnor U21193 (N_21193,N_15814,N_17968);
or U21194 (N_21194,N_16648,N_16470);
and U21195 (N_21195,N_16139,N_15697);
or U21196 (N_21196,N_16419,N_17396);
and U21197 (N_21197,N_17002,N_18359);
or U21198 (N_21198,N_15880,N_17082);
or U21199 (N_21199,N_16549,N_18514);
and U21200 (N_21200,N_16239,N_16569);
and U21201 (N_21201,N_16017,N_16955);
nand U21202 (N_21202,N_18138,N_18672);
nand U21203 (N_21203,N_16783,N_16051);
and U21204 (N_21204,N_17994,N_17211);
nor U21205 (N_21205,N_16556,N_16735);
nor U21206 (N_21206,N_17373,N_16387);
or U21207 (N_21207,N_15898,N_17062);
nor U21208 (N_21208,N_16739,N_15702);
xor U21209 (N_21209,N_17694,N_16925);
or U21210 (N_21210,N_17748,N_16348);
xor U21211 (N_21211,N_16069,N_16698);
or U21212 (N_21212,N_16514,N_17159);
and U21213 (N_21213,N_17328,N_16656);
and U21214 (N_21214,N_17844,N_17847);
and U21215 (N_21215,N_16072,N_18034);
nand U21216 (N_21216,N_17119,N_16988);
or U21217 (N_21217,N_15890,N_17798);
nand U21218 (N_21218,N_17448,N_16564);
or U21219 (N_21219,N_16948,N_17739);
or U21220 (N_21220,N_18290,N_16382);
xor U21221 (N_21221,N_16123,N_16723);
or U21222 (N_21222,N_16849,N_17830);
nand U21223 (N_21223,N_18430,N_17756);
nand U21224 (N_21224,N_15654,N_17319);
nand U21225 (N_21225,N_16919,N_18656);
or U21226 (N_21226,N_18597,N_16894);
nand U21227 (N_21227,N_16705,N_17668);
and U21228 (N_21228,N_18651,N_17149);
or U21229 (N_21229,N_18736,N_18499);
and U21230 (N_21230,N_18685,N_15687);
and U21231 (N_21231,N_18646,N_16186);
and U21232 (N_21232,N_16549,N_17943);
nor U21233 (N_21233,N_17302,N_16970);
and U21234 (N_21234,N_16402,N_15705);
or U21235 (N_21235,N_18178,N_18598);
and U21236 (N_21236,N_15981,N_18129);
nand U21237 (N_21237,N_16429,N_17089);
and U21238 (N_21238,N_16056,N_17928);
and U21239 (N_21239,N_17911,N_18193);
nand U21240 (N_21240,N_17130,N_18062);
xnor U21241 (N_21241,N_18593,N_18258);
nand U21242 (N_21242,N_17855,N_16289);
or U21243 (N_21243,N_15763,N_17676);
and U21244 (N_21244,N_15914,N_17125);
xnor U21245 (N_21245,N_18658,N_16958);
or U21246 (N_21246,N_18266,N_15882);
nand U21247 (N_21247,N_17948,N_15748);
or U21248 (N_21248,N_16493,N_17475);
and U21249 (N_21249,N_18200,N_17298);
nor U21250 (N_21250,N_16797,N_17481);
xnor U21251 (N_21251,N_18056,N_18705);
nor U21252 (N_21252,N_16555,N_17525);
nand U21253 (N_21253,N_15876,N_15800);
xnor U21254 (N_21254,N_16746,N_17706);
nand U21255 (N_21255,N_17785,N_17062);
or U21256 (N_21256,N_16652,N_18381);
and U21257 (N_21257,N_16758,N_17825);
and U21258 (N_21258,N_17715,N_16782);
nor U21259 (N_21259,N_18213,N_16491);
nand U21260 (N_21260,N_18624,N_16238);
and U21261 (N_21261,N_17988,N_16684);
and U21262 (N_21262,N_18496,N_17933);
or U21263 (N_21263,N_18477,N_18661);
nor U21264 (N_21264,N_18237,N_17139);
nor U21265 (N_21265,N_17093,N_18323);
nor U21266 (N_21266,N_17310,N_17049);
nor U21267 (N_21267,N_18617,N_18561);
or U21268 (N_21268,N_16612,N_17268);
nand U21269 (N_21269,N_15912,N_16186);
nor U21270 (N_21270,N_15730,N_16819);
or U21271 (N_21271,N_15679,N_16849);
or U21272 (N_21272,N_15915,N_16039);
nand U21273 (N_21273,N_17011,N_18110);
and U21274 (N_21274,N_18101,N_16172);
and U21275 (N_21275,N_18681,N_18542);
or U21276 (N_21276,N_18629,N_17937);
nor U21277 (N_21277,N_17768,N_16746);
or U21278 (N_21278,N_17556,N_18300);
and U21279 (N_21279,N_16007,N_16437);
and U21280 (N_21280,N_17473,N_16824);
nor U21281 (N_21281,N_15944,N_18584);
nor U21282 (N_21282,N_16662,N_17354);
and U21283 (N_21283,N_18307,N_16818);
and U21284 (N_21284,N_17414,N_17908);
nand U21285 (N_21285,N_16275,N_16420);
and U21286 (N_21286,N_16797,N_17940);
or U21287 (N_21287,N_17168,N_16754);
nor U21288 (N_21288,N_17386,N_15831);
or U21289 (N_21289,N_15823,N_16534);
and U21290 (N_21290,N_17008,N_18279);
nand U21291 (N_21291,N_18726,N_18212);
nor U21292 (N_21292,N_17347,N_16817);
nor U21293 (N_21293,N_17344,N_17929);
and U21294 (N_21294,N_15731,N_18023);
nand U21295 (N_21295,N_18303,N_16489);
nand U21296 (N_21296,N_17015,N_15854);
or U21297 (N_21297,N_17717,N_18217);
and U21298 (N_21298,N_16713,N_17030);
nand U21299 (N_21299,N_17556,N_18503);
nor U21300 (N_21300,N_16603,N_15752);
and U21301 (N_21301,N_17655,N_18018);
and U21302 (N_21302,N_15652,N_17525);
nor U21303 (N_21303,N_18064,N_18475);
and U21304 (N_21304,N_18232,N_18289);
or U21305 (N_21305,N_17054,N_17324);
or U21306 (N_21306,N_18700,N_17593);
or U21307 (N_21307,N_16045,N_17644);
nand U21308 (N_21308,N_16662,N_17761);
nor U21309 (N_21309,N_16417,N_18701);
xnor U21310 (N_21310,N_16286,N_17959);
nor U21311 (N_21311,N_15699,N_18658);
and U21312 (N_21312,N_17726,N_15777);
nand U21313 (N_21313,N_15916,N_16144);
nor U21314 (N_21314,N_17267,N_16409);
and U21315 (N_21315,N_17576,N_16203);
and U21316 (N_21316,N_16600,N_18710);
and U21317 (N_21317,N_18305,N_18605);
nand U21318 (N_21318,N_17031,N_15701);
xor U21319 (N_21319,N_16473,N_17520);
xnor U21320 (N_21320,N_18346,N_18419);
or U21321 (N_21321,N_18425,N_16591);
and U21322 (N_21322,N_17627,N_16996);
xor U21323 (N_21323,N_16143,N_17634);
or U21324 (N_21324,N_16613,N_16384);
or U21325 (N_21325,N_18485,N_17656);
nand U21326 (N_21326,N_17375,N_18507);
and U21327 (N_21327,N_17985,N_15708);
or U21328 (N_21328,N_16507,N_18389);
xor U21329 (N_21329,N_18566,N_18454);
and U21330 (N_21330,N_17950,N_18373);
or U21331 (N_21331,N_16427,N_15893);
nand U21332 (N_21332,N_18143,N_16072);
nand U21333 (N_21333,N_16184,N_17603);
nor U21334 (N_21334,N_17723,N_16382);
nand U21335 (N_21335,N_17752,N_18411);
or U21336 (N_21336,N_18565,N_15937);
nor U21337 (N_21337,N_17478,N_16227);
nor U21338 (N_21338,N_17411,N_17274);
nand U21339 (N_21339,N_15754,N_17973);
nor U21340 (N_21340,N_15949,N_17950);
or U21341 (N_21341,N_16096,N_17750);
or U21342 (N_21342,N_17520,N_18096);
nor U21343 (N_21343,N_16761,N_18538);
or U21344 (N_21344,N_16015,N_17412);
nand U21345 (N_21345,N_17382,N_15896);
or U21346 (N_21346,N_17747,N_15751);
nor U21347 (N_21347,N_15936,N_17748);
or U21348 (N_21348,N_18003,N_17894);
nor U21349 (N_21349,N_15814,N_16072);
or U21350 (N_21350,N_16268,N_17393);
or U21351 (N_21351,N_16299,N_15916);
nor U21352 (N_21352,N_18064,N_15724);
nor U21353 (N_21353,N_16809,N_18510);
and U21354 (N_21354,N_17053,N_17609);
nand U21355 (N_21355,N_16091,N_16631);
or U21356 (N_21356,N_17363,N_15971);
or U21357 (N_21357,N_18671,N_16311);
nor U21358 (N_21358,N_18720,N_16510);
or U21359 (N_21359,N_16105,N_16048);
nand U21360 (N_21360,N_16166,N_16510);
nand U21361 (N_21361,N_16242,N_16498);
nand U21362 (N_21362,N_18633,N_16064);
nand U21363 (N_21363,N_18205,N_15712);
and U21364 (N_21364,N_17906,N_18013);
nand U21365 (N_21365,N_16161,N_16210);
or U21366 (N_21366,N_16972,N_18061);
or U21367 (N_21367,N_17121,N_16552);
nand U21368 (N_21368,N_16451,N_16420);
and U21369 (N_21369,N_18075,N_17042);
nand U21370 (N_21370,N_17002,N_16737);
and U21371 (N_21371,N_18735,N_15843);
or U21372 (N_21372,N_15950,N_17792);
or U21373 (N_21373,N_18259,N_16725);
nor U21374 (N_21374,N_17760,N_16331);
and U21375 (N_21375,N_16084,N_17486);
xor U21376 (N_21376,N_17834,N_16867);
xor U21377 (N_21377,N_17312,N_15928);
nand U21378 (N_21378,N_16448,N_18420);
or U21379 (N_21379,N_17755,N_17613);
nand U21380 (N_21380,N_16241,N_16613);
nand U21381 (N_21381,N_17262,N_18253);
xnor U21382 (N_21382,N_15705,N_18504);
nand U21383 (N_21383,N_16056,N_17670);
nor U21384 (N_21384,N_16876,N_17008);
and U21385 (N_21385,N_16980,N_16499);
nand U21386 (N_21386,N_17957,N_16957);
nand U21387 (N_21387,N_16538,N_16989);
or U21388 (N_21388,N_17954,N_16637);
or U21389 (N_21389,N_15773,N_17102);
and U21390 (N_21390,N_17549,N_16219);
xnor U21391 (N_21391,N_18341,N_18631);
nor U21392 (N_21392,N_16568,N_17078);
xor U21393 (N_21393,N_18350,N_16794);
and U21394 (N_21394,N_15927,N_18619);
nor U21395 (N_21395,N_15673,N_18038);
and U21396 (N_21396,N_16254,N_15875);
nand U21397 (N_21397,N_18612,N_15718);
xor U21398 (N_21398,N_18580,N_15972);
nand U21399 (N_21399,N_17317,N_18144);
or U21400 (N_21400,N_17410,N_16359);
or U21401 (N_21401,N_18293,N_16806);
nand U21402 (N_21402,N_15691,N_15827);
nand U21403 (N_21403,N_18654,N_16829);
or U21404 (N_21404,N_16879,N_16453);
nand U21405 (N_21405,N_18287,N_16300);
nor U21406 (N_21406,N_17099,N_16046);
and U21407 (N_21407,N_15856,N_18629);
nor U21408 (N_21408,N_16676,N_15960);
or U21409 (N_21409,N_17170,N_16909);
nand U21410 (N_21410,N_16640,N_17624);
or U21411 (N_21411,N_15781,N_18335);
nand U21412 (N_21412,N_16711,N_17385);
nand U21413 (N_21413,N_18381,N_18293);
and U21414 (N_21414,N_17113,N_17687);
nor U21415 (N_21415,N_18182,N_16829);
or U21416 (N_21416,N_17893,N_16302);
or U21417 (N_21417,N_16923,N_17369);
nand U21418 (N_21418,N_17992,N_18452);
and U21419 (N_21419,N_18553,N_17454);
or U21420 (N_21420,N_15968,N_16298);
nand U21421 (N_21421,N_16387,N_16991);
nor U21422 (N_21422,N_16621,N_15965);
xnor U21423 (N_21423,N_17014,N_16291);
and U21424 (N_21424,N_17717,N_18027);
and U21425 (N_21425,N_16821,N_15763);
xnor U21426 (N_21426,N_16328,N_17654);
or U21427 (N_21427,N_16725,N_16318);
nor U21428 (N_21428,N_17413,N_18238);
nor U21429 (N_21429,N_15743,N_17302);
nor U21430 (N_21430,N_17756,N_16214);
nand U21431 (N_21431,N_15643,N_16233);
and U21432 (N_21432,N_15717,N_17384);
nand U21433 (N_21433,N_18647,N_18078);
nand U21434 (N_21434,N_16955,N_16141);
nor U21435 (N_21435,N_16331,N_16719);
nand U21436 (N_21436,N_17141,N_17181);
xor U21437 (N_21437,N_18420,N_15635);
nor U21438 (N_21438,N_16698,N_17613);
or U21439 (N_21439,N_16817,N_16542);
nand U21440 (N_21440,N_16675,N_15898);
xnor U21441 (N_21441,N_16638,N_17867);
nand U21442 (N_21442,N_17530,N_16475);
and U21443 (N_21443,N_15700,N_16093);
and U21444 (N_21444,N_15697,N_18122);
nand U21445 (N_21445,N_15713,N_17848);
and U21446 (N_21446,N_16782,N_17160);
nand U21447 (N_21447,N_17506,N_16870);
nor U21448 (N_21448,N_18656,N_16106);
xnor U21449 (N_21449,N_17355,N_17014);
xor U21450 (N_21450,N_15906,N_18214);
and U21451 (N_21451,N_18547,N_17583);
nand U21452 (N_21452,N_17668,N_16416);
and U21453 (N_21453,N_17584,N_16252);
nor U21454 (N_21454,N_16903,N_17609);
or U21455 (N_21455,N_18307,N_16127);
or U21456 (N_21456,N_16842,N_17385);
nor U21457 (N_21457,N_18177,N_16049);
or U21458 (N_21458,N_15707,N_16694);
nand U21459 (N_21459,N_17088,N_15754);
nand U21460 (N_21460,N_15953,N_17381);
nand U21461 (N_21461,N_16099,N_17952);
or U21462 (N_21462,N_18663,N_17601);
nand U21463 (N_21463,N_17477,N_16548);
or U21464 (N_21464,N_18545,N_18058);
nand U21465 (N_21465,N_17013,N_18247);
or U21466 (N_21466,N_18572,N_16571);
nand U21467 (N_21467,N_17300,N_15861);
or U21468 (N_21468,N_18526,N_17577);
or U21469 (N_21469,N_17733,N_18452);
nand U21470 (N_21470,N_17528,N_17626);
nor U21471 (N_21471,N_18691,N_16736);
and U21472 (N_21472,N_17625,N_18562);
nor U21473 (N_21473,N_16898,N_17651);
nand U21474 (N_21474,N_15812,N_17012);
or U21475 (N_21475,N_17515,N_18621);
and U21476 (N_21476,N_17210,N_17805);
nand U21477 (N_21477,N_15911,N_18145);
or U21478 (N_21478,N_16094,N_16491);
xnor U21479 (N_21479,N_17845,N_17416);
nand U21480 (N_21480,N_18108,N_17219);
nand U21481 (N_21481,N_17661,N_16860);
nand U21482 (N_21482,N_15836,N_16068);
nand U21483 (N_21483,N_15820,N_17705);
nor U21484 (N_21484,N_16382,N_17924);
or U21485 (N_21485,N_17086,N_16863);
nor U21486 (N_21486,N_18698,N_17941);
xnor U21487 (N_21487,N_16209,N_17706);
or U21488 (N_21488,N_16649,N_18485);
nand U21489 (N_21489,N_16788,N_17242);
xnor U21490 (N_21490,N_15968,N_18270);
nand U21491 (N_21491,N_16203,N_18389);
nor U21492 (N_21492,N_17843,N_16723);
or U21493 (N_21493,N_16317,N_17037);
nor U21494 (N_21494,N_16314,N_18522);
xor U21495 (N_21495,N_16115,N_17444);
xnor U21496 (N_21496,N_18155,N_18043);
or U21497 (N_21497,N_18599,N_15911);
nand U21498 (N_21498,N_18495,N_16826);
and U21499 (N_21499,N_18109,N_16413);
nand U21500 (N_21500,N_16500,N_18337);
nand U21501 (N_21501,N_16270,N_18114);
nor U21502 (N_21502,N_18602,N_18689);
and U21503 (N_21503,N_17796,N_16018);
or U21504 (N_21504,N_15644,N_15871);
and U21505 (N_21505,N_17131,N_16571);
nor U21506 (N_21506,N_17971,N_18679);
nand U21507 (N_21507,N_16175,N_16650);
xnor U21508 (N_21508,N_17117,N_17371);
and U21509 (N_21509,N_15967,N_16615);
and U21510 (N_21510,N_15839,N_15952);
or U21511 (N_21511,N_18278,N_17181);
or U21512 (N_21512,N_15978,N_18564);
nand U21513 (N_21513,N_18548,N_18013);
or U21514 (N_21514,N_16167,N_17365);
nand U21515 (N_21515,N_16527,N_18589);
or U21516 (N_21516,N_16645,N_18573);
and U21517 (N_21517,N_17389,N_17380);
nand U21518 (N_21518,N_16558,N_18263);
nor U21519 (N_21519,N_15783,N_16958);
and U21520 (N_21520,N_18359,N_16362);
nor U21521 (N_21521,N_18158,N_16580);
or U21522 (N_21522,N_16057,N_18209);
nand U21523 (N_21523,N_16764,N_15944);
or U21524 (N_21524,N_17322,N_16246);
and U21525 (N_21525,N_17949,N_15960);
or U21526 (N_21526,N_18116,N_17122);
nor U21527 (N_21527,N_17116,N_16777);
xnor U21528 (N_21528,N_18255,N_17303);
nor U21529 (N_21529,N_15732,N_17954);
or U21530 (N_21530,N_17399,N_17182);
and U21531 (N_21531,N_17209,N_17596);
nor U21532 (N_21532,N_17814,N_16178);
nand U21533 (N_21533,N_18096,N_17029);
nand U21534 (N_21534,N_17828,N_16945);
or U21535 (N_21535,N_17375,N_15852);
nor U21536 (N_21536,N_16381,N_18057);
nor U21537 (N_21537,N_16469,N_18147);
nand U21538 (N_21538,N_18434,N_18000);
or U21539 (N_21539,N_16740,N_16206);
xor U21540 (N_21540,N_18103,N_16168);
xnor U21541 (N_21541,N_17984,N_16459);
nor U21542 (N_21542,N_17614,N_16315);
nor U21543 (N_21543,N_17990,N_17834);
nand U21544 (N_21544,N_17567,N_16864);
and U21545 (N_21545,N_16681,N_16232);
nand U21546 (N_21546,N_16879,N_16760);
nand U21547 (N_21547,N_15646,N_16972);
and U21548 (N_21548,N_18559,N_17031);
or U21549 (N_21549,N_15663,N_18603);
or U21550 (N_21550,N_17995,N_16874);
nor U21551 (N_21551,N_18610,N_18735);
nand U21552 (N_21552,N_17421,N_17072);
or U21553 (N_21553,N_17123,N_16343);
nor U21554 (N_21554,N_17025,N_15720);
xor U21555 (N_21555,N_15945,N_16945);
and U21556 (N_21556,N_18426,N_16451);
nand U21557 (N_21557,N_16774,N_18561);
and U21558 (N_21558,N_17648,N_17588);
xnor U21559 (N_21559,N_16018,N_16369);
or U21560 (N_21560,N_18604,N_16894);
and U21561 (N_21561,N_16467,N_18663);
nand U21562 (N_21562,N_15858,N_18089);
nand U21563 (N_21563,N_16815,N_16367);
nand U21564 (N_21564,N_17104,N_16677);
or U21565 (N_21565,N_17460,N_15828);
and U21566 (N_21566,N_17307,N_18649);
and U21567 (N_21567,N_17564,N_17732);
nand U21568 (N_21568,N_18473,N_15968);
xor U21569 (N_21569,N_15961,N_18099);
nor U21570 (N_21570,N_16975,N_18348);
nor U21571 (N_21571,N_17062,N_15714);
or U21572 (N_21572,N_16372,N_17034);
nor U21573 (N_21573,N_16878,N_17273);
nand U21574 (N_21574,N_18669,N_16540);
nor U21575 (N_21575,N_16707,N_15891);
and U21576 (N_21576,N_17076,N_18417);
xnor U21577 (N_21577,N_17473,N_18022);
nor U21578 (N_21578,N_17893,N_16596);
nor U21579 (N_21579,N_18678,N_15655);
and U21580 (N_21580,N_17561,N_17244);
or U21581 (N_21581,N_16912,N_16119);
and U21582 (N_21582,N_17745,N_18461);
and U21583 (N_21583,N_16096,N_17116);
nand U21584 (N_21584,N_16584,N_18014);
nand U21585 (N_21585,N_18269,N_16576);
nor U21586 (N_21586,N_17348,N_16791);
or U21587 (N_21587,N_16966,N_15773);
and U21588 (N_21588,N_18198,N_17745);
nand U21589 (N_21589,N_16341,N_18107);
or U21590 (N_21590,N_15728,N_16168);
nand U21591 (N_21591,N_16933,N_16350);
nor U21592 (N_21592,N_16525,N_17868);
xor U21593 (N_21593,N_17821,N_16486);
nand U21594 (N_21594,N_18062,N_18198);
or U21595 (N_21595,N_17909,N_18319);
or U21596 (N_21596,N_18164,N_17695);
nor U21597 (N_21597,N_16064,N_15782);
or U21598 (N_21598,N_18321,N_17728);
or U21599 (N_21599,N_15890,N_15813);
or U21600 (N_21600,N_15960,N_15650);
nand U21601 (N_21601,N_18701,N_16663);
xnor U21602 (N_21602,N_18320,N_16122);
nand U21603 (N_21603,N_15642,N_17078);
and U21604 (N_21604,N_16554,N_16431);
and U21605 (N_21605,N_17474,N_16113);
or U21606 (N_21606,N_16026,N_16945);
xnor U21607 (N_21607,N_17917,N_17117);
xor U21608 (N_21608,N_16054,N_18410);
or U21609 (N_21609,N_15937,N_18399);
nor U21610 (N_21610,N_16786,N_17158);
nand U21611 (N_21611,N_17488,N_18063);
nand U21612 (N_21612,N_17905,N_15906);
or U21613 (N_21613,N_16875,N_15848);
nor U21614 (N_21614,N_17654,N_16747);
xnor U21615 (N_21615,N_16280,N_17286);
xor U21616 (N_21616,N_16231,N_15773);
and U21617 (N_21617,N_15805,N_18747);
and U21618 (N_21618,N_15696,N_16911);
and U21619 (N_21619,N_17165,N_17711);
or U21620 (N_21620,N_17155,N_16007);
nor U21621 (N_21621,N_18544,N_17302);
xnor U21622 (N_21622,N_16247,N_16166);
nand U21623 (N_21623,N_17680,N_17493);
nor U21624 (N_21624,N_16599,N_17162);
nand U21625 (N_21625,N_18402,N_17654);
xor U21626 (N_21626,N_16117,N_18377);
and U21627 (N_21627,N_15673,N_17369);
nand U21628 (N_21628,N_16605,N_16013);
nor U21629 (N_21629,N_17509,N_15869);
nand U21630 (N_21630,N_17299,N_18517);
xor U21631 (N_21631,N_17127,N_18726);
nor U21632 (N_21632,N_17222,N_15754);
nand U21633 (N_21633,N_17806,N_18404);
and U21634 (N_21634,N_18491,N_17498);
and U21635 (N_21635,N_16499,N_15901);
xnor U21636 (N_21636,N_18322,N_18492);
or U21637 (N_21637,N_17467,N_17010);
nor U21638 (N_21638,N_18425,N_18595);
nand U21639 (N_21639,N_16841,N_17489);
nand U21640 (N_21640,N_17864,N_15853);
and U21641 (N_21641,N_15816,N_17826);
or U21642 (N_21642,N_15753,N_15877);
or U21643 (N_21643,N_18737,N_17074);
and U21644 (N_21644,N_16476,N_15792);
or U21645 (N_21645,N_18176,N_17721);
or U21646 (N_21646,N_17234,N_16053);
nor U21647 (N_21647,N_17105,N_17262);
nor U21648 (N_21648,N_17572,N_15634);
nand U21649 (N_21649,N_18559,N_16794);
nor U21650 (N_21650,N_16675,N_15841);
nand U21651 (N_21651,N_17437,N_18356);
nor U21652 (N_21652,N_17434,N_17255);
and U21653 (N_21653,N_18467,N_17609);
nor U21654 (N_21654,N_17963,N_17498);
and U21655 (N_21655,N_18263,N_17284);
and U21656 (N_21656,N_16487,N_17326);
or U21657 (N_21657,N_17682,N_17835);
nand U21658 (N_21658,N_18220,N_16919);
and U21659 (N_21659,N_16593,N_15625);
and U21660 (N_21660,N_18591,N_17316);
nor U21661 (N_21661,N_16655,N_17572);
or U21662 (N_21662,N_16402,N_16536);
nand U21663 (N_21663,N_18631,N_16504);
and U21664 (N_21664,N_18440,N_17307);
or U21665 (N_21665,N_17816,N_17140);
and U21666 (N_21666,N_15675,N_18073);
and U21667 (N_21667,N_17088,N_16862);
or U21668 (N_21668,N_17338,N_15693);
and U21669 (N_21669,N_16822,N_18253);
or U21670 (N_21670,N_17686,N_16421);
nor U21671 (N_21671,N_18667,N_18151);
nor U21672 (N_21672,N_16095,N_17844);
or U21673 (N_21673,N_17861,N_15802);
nand U21674 (N_21674,N_15954,N_16714);
xor U21675 (N_21675,N_18592,N_18687);
nand U21676 (N_21676,N_15822,N_17124);
and U21677 (N_21677,N_18159,N_17200);
nand U21678 (N_21678,N_17760,N_16507);
nand U21679 (N_21679,N_16272,N_15824);
and U21680 (N_21680,N_18005,N_18051);
nor U21681 (N_21681,N_17310,N_18296);
and U21682 (N_21682,N_15655,N_17777);
nand U21683 (N_21683,N_17878,N_15924);
xnor U21684 (N_21684,N_16623,N_16086);
and U21685 (N_21685,N_16322,N_16395);
and U21686 (N_21686,N_16556,N_17065);
xor U21687 (N_21687,N_17425,N_18007);
nand U21688 (N_21688,N_18609,N_17658);
nor U21689 (N_21689,N_17685,N_17534);
nand U21690 (N_21690,N_16030,N_15774);
xnor U21691 (N_21691,N_17362,N_16077);
or U21692 (N_21692,N_15791,N_17018);
or U21693 (N_21693,N_17736,N_18724);
or U21694 (N_21694,N_16834,N_18030);
nor U21695 (N_21695,N_18502,N_16051);
and U21696 (N_21696,N_17296,N_16188);
or U21697 (N_21697,N_18519,N_17631);
nor U21698 (N_21698,N_18289,N_15888);
nor U21699 (N_21699,N_17158,N_17916);
and U21700 (N_21700,N_16961,N_15682);
or U21701 (N_21701,N_17593,N_18707);
xnor U21702 (N_21702,N_18342,N_15987);
nand U21703 (N_21703,N_18633,N_17804);
and U21704 (N_21704,N_18184,N_18210);
or U21705 (N_21705,N_18055,N_17728);
and U21706 (N_21706,N_16516,N_15878);
or U21707 (N_21707,N_17083,N_16566);
nand U21708 (N_21708,N_18732,N_18094);
nand U21709 (N_21709,N_18356,N_15733);
or U21710 (N_21710,N_17850,N_18501);
nor U21711 (N_21711,N_17871,N_16547);
nor U21712 (N_21712,N_17570,N_18212);
nand U21713 (N_21713,N_15861,N_16272);
and U21714 (N_21714,N_18544,N_16753);
and U21715 (N_21715,N_17643,N_17849);
nand U21716 (N_21716,N_16701,N_18423);
and U21717 (N_21717,N_16917,N_17704);
nand U21718 (N_21718,N_18528,N_18610);
or U21719 (N_21719,N_18356,N_16699);
and U21720 (N_21720,N_17971,N_16339);
xnor U21721 (N_21721,N_16498,N_18523);
or U21722 (N_21722,N_18268,N_18401);
and U21723 (N_21723,N_16787,N_16474);
and U21724 (N_21724,N_18043,N_17976);
and U21725 (N_21725,N_16182,N_16210);
nand U21726 (N_21726,N_18401,N_16934);
nor U21727 (N_21727,N_18522,N_16542);
nor U21728 (N_21728,N_17870,N_18345);
nand U21729 (N_21729,N_17580,N_16228);
nor U21730 (N_21730,N_16797,N_15983);
nor U21731 (N_21731,N_15787,N_18615);
and U21732 (N_21732,N_17273,N_16845);
and U21733 (N_21733,N_16744,N_16182);
nand U21734 (N_21734,N_17946,N_17312);
or U21735 (N_21735,N_17665,N_17926);
nand U21736 (N_21736,N_15914,N_17576);
nand U21737 (N_21737,N_16587,N_18182);
nor U21738 (N_21738,N_15798,N_15683);
or U21739 (N_21739,N_15976,N_18455);
nand U21740 (N_21740,N_17409,N_16196);
and U21741 (N_21741,N_16873,N_16654);
and U21742 (N_21742,N_16275,N_18282);
and U21743 (N_21743,N_16821,N_16505);
nor U21744 (N_21744,N_17620,N_17574);
or U21745 (N_21745,N_18230,N_15705);
nor U21746 (N_21746,N_17589,N_15656);
nor U21747 (N_21747,N_17480,N_16147);
nand U21748 (N_21748,N_18068,N_16448);
nand U21749 (N_21749,N_17979,N_16543);
and U21750 (N_21750,N_17141,N_16044);
nor U21751 (N_21751,N_16342,N_16816);
nor U21752 (N_21752,N_17064,N_17948);
or U21753 (N_21753,N_17959,N_16788);
or U21754 (N_21754,N_18072,N_17173);
and U21755 (N_21755,N_16613,N_17946);
nand U21756 (N_21756,N_16067,N_17656);
nor U21757 (N_21757,N_16484,N_16551);
xor U21758 (N_21758,N_17046,N_17042);
nor U21759 (N_21759,N_18155,N_18702);
nand U21760 (N_21760,N_15910,N_17861);
and U21761 (N_21761,N_16850,N_18435);
nand U21762 (N_21762,N_15663,N_17595);
nand U21763 (N_21763,N_16860,N_17838);
and U21764 (N_21764,N_18609,N_15851);
and U21765 (N_21765,N_18632,N_18111);
nor U21766 (N_21766,N_17709,N_18220);
xnor U21767 (N_21767,N_18654,N_18197);
and U21768 (N_21768,N_16144,N_18622);
or U21769 (N_21769,N_17325,N_15687);
or U21770 (N_21770,N_16695,N_18735);
xnor U21771 (N_21771,N_18684,N_16733);
and U21772 (N_21772,N_17444,N_18247);
nor U21773 (N_21773,N_16745,N_17084);
nor U21774 (N_21774,N_17965,N_18527);
and U21775 (N_21775,N_16840,N_17721);
nor U21776 (N_21776,N_18552,N_16585);
or U21777 (N_21777,N_18330,N_18135);
or U21778 (N_21778,N_16467,N_15808);
or U21779 (N_21779,N_18445,N_17305);
xor U21780 (N_21780,N_17027,N_15687);
nand U21781 (N_21781,N_18404,N_16042);
and U21782 (N_21782,N_18680,N_17979);
or U21783 (N_21783,N_17323,N_18030);
or U21784 (N_21784,N_17733,N_17395);
nand U21785 (N_21785,N_15865,N_18201);
xor U21786 (N_21786,N_18537,N_16331);
or U21787 (N_21787,N_16871,N_18148);
nand U21788 (N_21788,N_18469,N_18518);
nor U21789 (N_21789,N_18600,N_18315);
nand U21790 (N_21790,N_17126,N_18185);
nand U21791 (N_21791,N_16090,N_17943);
and U21792 (N_21792,N_17216,N_18263);
or U21793 (N_21793,N_16579,N_18553);
and U21794 (N_21794,N_15748,N_17064);
and U21795 (N_21795,N_16033,N_17996);
and U21796 (N_21796,N_17148,N_18466);
nor U21797 (N_21797,N_17540,N_18118);
xnor U21798 (N_21798,N_18212,N_17069);
or U21799 (N_21799,N_16146,N_18472);
or U21800 (N_21800,N_17001,N_15985);
nor U21801 (N_21801,N_18634,N_17405);
xor U21802 (N_21802,N_15734,N_15825);
nand U21803 (N_21803,N_16129,N_16975);
or U21804 (N_21804,N_16254,N_16359);
nand U21805 (N_21805,N_15798,N_17065);
or U21806 (N_21806,N_15803,N_18565);
and U21807 (N_21807,N_18615,N_16651);
nor U21808 (N_21808,N_17148,N_16052);
or U21809 (N_21809,N_17413,N_15784);
xnor U21810 (N_21810,N_16676,N_17232);
nand U21811 (N_21811,N_18194,N_16118);
nand U21812 (N_21812,N_15732,N_16960);
nand U21813 (N_21813,N_16370,N_17971);
nand U21814 (N_21814,N_18237,N_18449);
nand U21815 (N_21815,N_17315,N_16525);
nand U21816 (N_21816,N_17722,N_16486);
or U21817 (N_21817,N_18224,N_17609);
xnor U21818 (N_21818,N_16442,N_16538);
and U21819 (N_21819,N_16196,N_15661);
xor U21820 (N_21820,N_17323,N_16565);
nand U21821 (N_21821,N_15970,N_16369);
or U21822 (N_21822,N_16593,N_17182);
nand U21823 (N_21823,N_15801,N_18056);
or U21824 (N_21824,N_15871,N_17511);
and U21825 (N_21825,N_18409,N_17213);
nand U21826 (N_21826,N_17372,N_16974);
nand U21827 (N_21827,N_17039,N_17651);
nand U21828 (N_21828,N_16537,N_18088);
and U21829 (N_21829,N_17772,N_17337);
nand U21830 (N_21830,N_18036,N_16672);
nand U21831 (N_21831,N_18086,N_17682);
and U21832 (N_21832,N_17195,N_16369);
or U21833 (N_21833,N_17937,N_17680);
nand U21834 (N_21834,N_18380,N_16499);
and U21835 (N_21835,N_15694,N_16105);
nor U21836 (N_21836,N_15847,N_15693);
or U21837 (N_21837,N_17330,N_18712);
nor U21838 (N_21838,N_16410,N_17198);
or U21839 (N_21839,N_16654,N_16227);
xor U21840 (N_21840,N_17299,N_17802);
and U21841 (N_21841,N_17857,N_15928);
nor U21842 (N_21842,N_18247,N_15886);
xnor U21843 (N_21843,N_16272,N_16612);
nand U21844 (N_21844,N_15844,N_18523);
xor U21845 (N_21845,N_17204,N_16387);
or U21846 (N_21846,N_18278,N_15886);
nor U21847 (N_21847,N_18023,N_16415);
or U21848 (N_21848,N_17047,N_18246);
nand U21849 (N_21849,N_16542,N_17037);
and U21850 (N_21850,N_16537,N_17289);
or U21851 (N_21851,N_16208,N_16576);
nor U21852 (N_21852,N_15950,N_17619);
xor U21853 (N_21853,N_18352,N_17073);
xor U21854 (N_21854,N_16293,N_16342);
and U21855 (N_21855,N_18069,N_17899);
nor U21856 (N_21856,N_18489,N_17980);
or U21857 (N_21857,N_16198,N_15982);
nand U21858 (N_21858,N_17478,N_17707);
nand U21859 (N_21859,N_17445,N_18706);
nand U21860 (N_21860,N_17506,N_18730);
nor U21861 (N_21861,N_17209,N_18677);
and U21862 (N_21862,N_18740,N_15749);
and U21863 (N_21863,N_17966,N_15916);
nor U21864 (N_21864,N_17688,N_18012);
or U21865 (N_21865,N_15656,N_16105);
and U21866 (N_21866,N_18194,N_16507);
nor U21867 (N_21867,N_16381,N_16587);
nand U21868 (N_21868,N_15993,N_16174);
nor U21869 (N_21869,N_18467,N_17360);
nand U21870 (N_21870,N_18064,N_17308);
nor U21871 (N_21871,N_16435,N_17732);
nor U21872 (N_21872,N_15787,N_18331);
nand U21873 (N_21873,N_15758,N_16985);
xnor U21874 (N_21874,N_18287,N_17561);
and U21875 (N_21875,N_21796,N_20305);
xor U21876 (N_21876,N_19581,N_20184);
nor U21877 (N_21877,N_21643,N_19456);
and U21878 (N_21878,N_20566,N_20897);
nand U21879 (N_21879,N_18818,N_19479);
and U21880 (N_21880,N_19691,N_19416);
nand U21881 (N_21881,N_19882,N_20269);
nor U21882 (N_21882,N_18973,N_21004);
nand U21883 (N_21883,N_21627,N_18763);
nand U21884 (N_21884,N_21854,N_21618);
or U21885 (N_21885,N_19465,N_21253);
nor U21886 (N_21886,N_19150,N_21164);
and U21887 (N_21887,N_20694,N_21441);
nand U21888 (N_21888,N_19334,N_19787);
or U21889 (N_21889,N_21523,N_21695);
nor U21890 (N_21890,N_19534,N_21148);
nand U21891 (N_21891,N_21280,N_19936);
and U21892 (N_21892,N_20020,N_20976);
nand U21893 (N_21893,N_18812,N_20090);
or U21894 (N_21894,N_21031,N_19547);
xor U21895 (N_21895,N_20428,N_21120);
nor U21896 (N_21896,N_19764,N_21783);
or U21897 (N_21897,N_20414,N_21760);
nand U21898 (N_21898,N_20087,N_20000);
and U21899 (N_21899,N_21642,N_19022);
and U21900 (N_21900,N_21577,N_20454);
and U21901 (N_21901,N_20960,N_18945);
nand U21902 (N_21902,N_21590,N_20293);
or U21903 (N_21903,N_20874,N_19056);
nor U21904 (N_21904,N_19475,N_21487);
nor U21905 (N_21905,N_20544,N_21873);
or U21906 (N_21906,N_20202,N_19193);
or U21907 (N_21907,N_18795,N_19784);
or U21908 (N_21908,N_20858,N_19810);
nor U21909 (N_21909,N_19621,N_20353);
and U21910 (N_21910,N_19363,N_20558);
and U21911 (N_21911,N_21299,N_19926);
nand U21912 (N_21912,N_20740,N_20675);
nand U21913 (N_21913,N_21073,N_18957);
or U21914 (N_21914,N_21451,N_19945);
and U21915 (N_21915,N_20218,N_21419);
xor U21916 (N_21916,N_20879,N_20713);
or U21917 (N_21917,N_19722,N_19954);
and U21918 (N_21918,N_20791,N_19113);
nor U21919 (N_21919,N_21728,N_21630);
or U21920 (N_21920,N_20160,N_18950);
or U21921 (N_21921,N_21176,N_19459);
and U21922 (N_21922,N_20528,N_21082);
and U21923 (N_21923,N_20001,N_20506);
and U21924 (N_21924,N_20751,N_19120);
or U21925 (N_21925,N_19136,N_19713);
xnor U21926 (N_21926,N_21220,N_19437);
or U21927 (N_21927,N_19156,N_19793);
xnor U21928 (N_21928,N_21600,N_19385);
nor U21929 (N_21929,N_20650,N_20527);
nand U21930 (N_21930,N_19745,N_19551);
nor U21931 (N_21931,N_21532,N_18808);
or U21932 (N_21932,N_21302,N_21175);
and U21933 (N_21933,N_21314,N_18780);
nor U21934 (N_21934,N_20907,N_18881);
nor U21935 (N_21935,N_21689,N_19932);
nand U21936 (N_21936,N_18983,N_20229);
or U21937 (N_21937,N_19349,N_21411);
nand U21938 (N_21938,N_19281,N_19019);
and U21939 (N_21939,N_18842,N_20339);
nand U21940 (N_21940,N_20590,N_20403);
xnor U21941 (N_21941,N_20749,N_21115);
nand U21942 (N_21942,N_19242,N_20790);
or U21943 (N_21943,N_20582,N_21713);
nor U21944 (N_21944,N_20298,N_21461);
nor U21945 (N_21945,N_20194,N_20760);
nand U21946 (N_21946,N_20977,N_21428);
or U21947 (N_21947,N_19159,N_21271);
or U21948 (N_21948,N_19244,N_21503);
nor U21949 (N_21949,N_19278,N_19122);
or U21950 (N_21950,N_20030,N_21071);
nand U21951 (N_21951,N_19170,N_18828);
nand U21952 (N_21952,N_20376,N_19739);
nand U21953 (N_21953,N_19606,N_21799);
and U21954 (N_21954,N_21711,N_21807);
or U21955 (N_21955,N_21602,N_18868);
nor U21956 (N_21956,N_20913,N_20810);
xor U21957 (N_21957,N_21749,N_19161);
and U21958 (N_21958,N_21746,N_21651);
nand U21959 (N_21959,N_18946,N_19627);
nor U21960 (N_21960,N_19243,N_21112);
nor U21961 (N_21961,N_19636,N_19994);
or U21962 (N_21962,N_20841,N_20754);
and U21963 (N_21963,N_21816,N_19004);
nor U21964 (N_21964,N_19608,N_19339);
and U21965 (N_21965,N_21397,N_21401);
and U21966 (N_21966,N_21632,N_21826);
xor U21967 (N_21967,N_19563,N_19322);
nand U21968 (N_21968,N_21544,N_20507);
and U21969 (N_21969,N_20833,N_20445);
or U21970 (N_21970,N_21505,N_18769);
xnor U21971 (N_21971,N_20663,N_19844);
nand U21972 (N_21972,N_19185,N_19637);
nand U21973 (N_21973,N_21391,N_21554);
and U21974 (N_21974,N_20965,N_20739);
and U21975 (N_21975,N_20662,N_20613);
nand U21976 (N_21976,N_20670,N_21156);
nor U21977 (N_21977,N_20473,N_21692);
or U21978 (N_21978,N_19286,N_19507);
nor U21979 (N_21979,N_20022,N_20925);
nand U21980 (N_21980,N_19643,N_19013);
nand U21981 (N_21981,N_19556,N_18887);
or U21982 (N_21982,N_20608,N_19696);
nand U21983 (N_21983,N_20538,N_18863);
nand U21984 (N_21984,N_20183,N_19881);
and U21985 (N_21985,N_19993,N_20526);
nor U21986 (N_21986,N_20917,N_21623);
xnor U21987 (N_21987,N_20993,N_20695);
and U21988 (N_21988,N_21693,N_20711);
or U21989 (N_21989,N_19069,N_21536);
and U21990 (N_21990,N_21768,N_20921);
nor U21991 (N_21991,N_20583,N_21238);
or U21992 (N_21992,N_21430,N_21133);
nor U21993 (N_21993,N_19460,N_19367);
nor U21994 (N_21994,N_21326,N_18858);
and U21995 (N_21995,N_21561,N_21181);
xnor U21996 (N_21996,N_18920,N_20618);
nor U21997 (N_21997,N_21438,N_19112);
or U21998 (N_21998,N_19721,N_20870);
xor U21999 (N_21999,N_20035,N_18952);
xor U22000 (N_22000,N_20824,N_19045);
nand U22001 (N_22001,N_20683,N_19918);
and U22002 (N_22002,N_20640,N_19491);
and U22003 (N_22003,N_19355,N_21404);
xor U22004 (N_22004,N_19231,N_20730);
or U22005 (N_22005,N_21315,N_20919);
nor U22006 (N_22006,N_20441,N_21677);
nor U22007 (N_22007,N_19222,N_19845);
nor U22008 (N_22008,N_18935,N_19094);
nor U22009 (N_22009,N_19296,N_21227);
nor U22010 (N_22010,N_19701,N_19423);
nor U22011 (N_22011,N_19749,N_21566);
nor U22012 (N_22012,N_20010,N_20591);
and U22013 (N_22013,N_20132,N_21568);
and U22014 (N_22014,N_18848,N_20867);
nor U22015 (N_22015,N_20788,N_21433);
or U22016 (N_22016,N_20005,N_18809);
nand U22017 (N_22017,N_19861,N_20188);
xnor U22018 (N_22018,N_19252,N_20575);
xor U22019 (N_22019,N_21736,N_21103);
or U22020 (N_22020,N_20532,N_21061);
and U22021 (N_22021,N_19843,N_20280);
or U22022 (N_22022,N_21712,N_20467);
and U22023 (N_22023,N_21174,N_20828);
or U22024 (N_22024,N_21370,N_21637);
or U22025 (N_22025,N_20058,N_21694);
or U22026 (N_22026,N_20343,N_20379);
and U22027 (N_22027,N_21207,N_20360);
nor U22028 (N_22028,N_21169,N_19111);
or U22029 (N_22029,N_21398,N_21560);
and U22030 (N_22030,N_19870,N_21131);
or U22031 (N_22031,N_19481,N_19664);
or U22032 (N_22032,N_19405,N_18777);
or U22033 (N_22033,N_19699,N_18792);
nor U22034 (N_22034,N_21237,N_19478);
or U22035 (N_22035,N_21747,N_21846);
and U22036 (N_22036,N_20103,N_19531);
nand U22037 (N_22037,N_20084,N_20500);
nor U22038 (N_22038,N_20761,N_20692);
or U22039 (N_22039,N_21501,N_18804);
xor U22040 (N_22040,N_19674,N_20073);
nand U22041 (N_22041,N_21466,N_20580);
or U22042 (N_22042,N_20419,N_20083);
nand U22043 (N_22043,N_18879,N_20632);
and U22044 (N_22044,N_21603,N_21795);
or U22045 (N_22045,N_20180,N_21596);
nor U22046 (N_22046,N_20674,N_21187);
nor U22047 (N_22047,N_19376,N_19440);
or U22048 (N_22048,N_20644,N_21425);
nor U22049 (N_22049,N_21841,N_19950);
or U22050 (N_22050,N_21321,N_21160);
and U22051 (N_22051,N_20914,N_20517);
nor U22052 (N_22052,N_21308,N_19922);
or U22053 (N_22053,N_20519,N_18930);
and U22054 (N_22054,N_18895,N_19390);
nor U22055 (N_22055,N_20394,N_19106);
nand U22056 (N_22056,N_20933,N_20451);
nand U22057 (N_22057,N_19435,N_21682);
nand U22058 (N_22058,N_21406,N_19154);
nand U22059 (N_22059,N_18872,N_21723);
and U22060 (N_22060,N_20823,N_20936);
nor U22061 (N_22061,N_20775,N_18932);
and U22062 (N_22062,N_19003,N_19285);
and U22063 (N_22063,N_19591,N_21234);
nor U22064 (N_22064,N_19153,N_19868);
nor U22065 (N_22065,N_19829,N_19450);
nor U22066 (N_22066,N_21099,N_18794);
nor U22067 (N_22067,N_21292,N_19017);
and U22068 (N_22068,N_19024,N_21773);
nand U22069 (N_22069,N_20915,N_21469);
or U22070 (N_22070,N_20186,N_19648);
or U22071 (N_22071,N_18773,N_20942);
xnor U22072 (N_22072,N_19358,N_20474);
nand U22073 (N_22073,N_19959,N_21146);
xnor U22074 (N_22074,N_19832,N_21110);
xor U22075 (N_22075,N_19370,N_21126);
and U22076 (N_22076,N_19657,N_21435);
or U22077 (N_22077,N_19653,N_21384);
nand U22078 (N_22078,N_19138,N_20258);
nor U22079 (N_22079,N_20271,N_20391);
and U22080 (N_22080,N_19714,N_21387);
nor U22081 (N_22081,N_21067,N_20901);
and U22082 (N_22082,N_21564,N_21222);
and U22083 (N_22083,N_19720,N_20863);
or U22084 (N_22084,N_18834,N_21400);
nor U22085 (N_22085,N_21094,N_19488);
nor U22086 (N_22086,N_20122,N_19028);
nand U22087 (N_22087,N_20570,N_19307);
nor U22088 (N_22088,N_20288,N_21049);
or U22089 (N_22089,N_21291,N_21765);
or U22090 (N_22090,N_20226,N_21814);
or U22091 (N_22091,N_20461,N_20254);
nor U22092 (N_22092,N_20105,N_21450);
or U22093 (N_22093,N_20520,N_20050);
nand U22094 (N_22094,N_19527,N_18953);
or U22095 (N_22095,N_21255,N_19082);
nor U22096 (N_22096,N_19357,N_19249);
nor U22097 (N_22097,N_19291,N_21454);
nand U22098 (N_22098,N_20211,N_19913);
or U22099 (N_22099,N_20829,N_19825);
or U22100 (N_22100,N_21836,N_20198);
nor U22101 (N_22101,N_20676,N_19140);
and U22102 (N_22102,N_19126,N_18978);
and U22103 (N_22103,N_20755,N_21277);
nand U22104 (N_22104,N_20869,N_20435);
nor U22105 (N_22105,N_19522,N_19444);
nor U22106 (N_22106,N_20889,N_20167);
or U22107 (N_22107,N_19215,N_21290);
and U22108 (N_22108,N_20911,N_19890);
or U22109 (N_22109,N_20368,N_20512);
and U22110 (N_22110,N_20827,N_19824);
or U22111 (N_22111,N_19638,N_20954);
nand U22112 (N_22112,N_19923,N_19631);
or U22113 (N_22113,N_20310,N_19279);
nand U22114 (N_22114,N_20373,N_20943);
nor U22115 (N_22115,N_21265,N_20701);
xnor U22116 (N_22116,N_19521,N_19345);
and U22117 (N_22117,N_21332,N_21123);
xor U22118 (N_22118,N_19403,N_20770);
or U22119 (N_22119,N_20492,N_19752);
xor U22120 (N_22120,N_21348,N_21236);
nand U22121 (N_22121,N_19395,N_21646);
or U22122 (N_22122,N_19333,N_19748);
xor U22123 (N_22123,N_19183,N_19842);
nor U22124 (N_22124,N_19678,N_21581);
nor U22125 (N_22125,N_19030,N_19441);
nand U22126 (N_22126,N_19175,N_19624);
or U22127 (N_22127,N_20546,N_21008);
nand U22128 (N_22128,N_21463,N_20706);
and U22129 (N_22129,N_20563,N_19509);
or U22130 (N_22130,N_19195,N_20436);
nand U22131 (N_22131,N_18940,N_18951);
xnor U22132 (N_22132,N_19869,N_21090);
or U22133 (N_22133,N_20496,N_19075);
and U22134 (N_22134,N_19535,N_19233);
or U22135 (N_22135,N_21871,N_21353);
and U22136 (N_22136,N_21076,N_20647);
nand U22137 (N_22137,N_21471,N_20329);
and U22138 (N_22138,N_19110,N_19240);
nand U22139 (N_22139,N_19559,N_21431);
nor U22140 (N_22140,N_19059,N_19434);
nor U22141 (N_22141,N_20205,N_20266);
and U22142 (N_22142,N_20127,N_19942);
or U22143 (N_22143,N_19010,N_20352);
nor U22144 (N_22144,N_18867,N_19568);
nand U22145 (N_22145,N_20830,N_19071);
and U22146 (N_22146,N_20876,N_20894);
nand U22147 (N_22147,N_21699,N_19301);
nor U22148 (N_22148,N_21859,N_20295);
and U22149 (N_22149,N_19805,N_20263);
or U22150 (N_22150,N_19482,N_18901);
nand U22151 (N_22151,N_20171,N_21831);
or U22152 (N_22152,N_20985,N_18924);
or U22153 (N_22153,N_18847,N_20299);
nand U22154 (N_22154,N_20072,N_20795);
and U22155 (N_22155,N_21645,N_19238);
and U22156 (N_22156,N_19241,N_19511);
nor U22157 (N_22157,N_19773,N_19862);
nand U22158 (N_22158,N_19054,N_20958);
or U22159 (N_22159,N_19590,N_21057);
or U22160 (N_22160,N_19576,N_21352);
or U22161 (N_22161,N_19600,N_19571);
and U22162 (N_22162,N_20729,N_21139);
nor U22163 (N_22163,N_20763,N_20465);
or U22164 (N_22164,N_21337,N_19109);
nor U22165 (N_22165,N_18779,N_19410);
nand U22166 (N_22166,N_21247,N_21531);
and U22167 (N_22167,N_19496,N_21200);
and U22168 (N_22168,N_19131,N_19001);
or U22169 (N_22169,N_21163,N_19319);
nand U22170 (N_22170,N_20148,N_19850);
nor U22171 (N_22171,N_19676,N_18996);
and U22172 (N_22172,N_18776,N_19523);
nand U22173 (N_22173,N_20844,N_19719);
xor U22174 (N_22174,N_20251,N_20471);
or U22175 (N_22175,N_20158,N_20117);
xor U22176 (N_22176,N_20571,N_20625);
nor U22177 (N_22177,N_19171,N_21781);
nor U22178 (N_22178,N_19809,N_20645);
nand U22179 (N_22179,N_21583,N_18866);
or U22180 (N_22180,N_18775,N_19048);
xor U22181 (N_22181,N_19618,N_19029);
nand U22182 (N_22182,N_21444,N_20115);
nand U22183 (N_22183,N_21874,N_21495);
nor U22184 (N_22184,N_20497,N_21415);
nor U22185 (N_22185,N_18984,N_21250);
nor U22186 (N_22186,N_19062,N_21734);
or U22187 (N_22187,N_21235,N_18928);
nand U22188 (N_22188,N_20185,N_21785);
nor U22189 (N_22189,N_19934,N_19340);
nand U22190 (N_22190,N_19542,N_20780);
or U22191 (N_22191,N_19461,N_19689);
or U22192 (N_22192,N_21525,N_19213);
nand U22193 (N_22193,N_19851,N_21818);
or U22194 (N_22194,N_20557,N_20243);
nor U22195 (N_22195,N_21500,N_21239);
or U22196 (N_22196,N_18825,N_20980);
or U22197 (N_22197,N_21449,N_21072);
nor U22198 (N_22198,N_20585,N_19529);
xor U22199 (N_22199,N_21180,N_19573);
xnor U22200 (N_22200,N_18990,N_18814);
and U22201 (N_22201,N_19985,N_19765);
nand U22202 (N_22202,N_20262,N_21312);
nand U22203 (N_22203,N_21533,N_20025);
nor U22204 (N_22204,N_20837,N_20388);
or U22205 (N_22205,N_18991,N_21231);
or U22206 (N_22206,N_19768,N_19378);
nand U22207 (N_22207,N_20076,N_21043);
xnor U22208 (N_22208,N_20899,N_20698);
and U22209 (N_22209,N_21607,N_20935);
xnor U22210 (N_22210,N_20438,N_19284);
nor U22211 (N_22211,N_19312,N_20479);
or U22212 (N_22212,N_19342,N_19178);
and U22213 (N_22213,N_20151,N_21104);
and U22214 (N_22214,N_21518,N_19409);
nor U22215 (N_22215,N_19858,N_19822);
nand U22216 (N_22216,N_19282,N_20283);
or U22217 (N_22217,N_21092,N_21625);
nand U22218 (N_22218,N_19124,N_21085);
nor U22219 (N_22219,N_20399,N_21153);
xor U22220 (N_22220,N_20460,N_19495);
or U22221 (N_22221,N_18832,N_19381);
and U22222 (N_22222,N_19451,N_19099);
nor U22223 (N_22223,N_19211,N_19063);
nor U22224 (N_22224,N_20957,N_19912);
or U22225 (N_22225,N_20865,N_20809);
nand U22226 (N_22226,N_21707,N_18903);
xor U22227 (N_22227,N_20717,N_19694);
nor U22228 (N_22228,N_20137,N_21744);
nor U22229 (N_22229,N_21171,N_21591);
xnor U22230 (N_22230,N_19100,N_19371);
nand U22231 (N_22231,N_20725,N_19086);
nor U22232 (N_22232,N_19204,N_20284);
and U22233 (N_22233,N_19426,N_21389);
nand U22234 (N_22234,N_21409,N_21722);
or U22235 (N_22235,N_19782,N_19073);
and U22236 (N_22236,N_18937,N_21548);
and U22237 (N_22237,N_20176,N_21702);
and U22238 (N_22238,N_21361,N_19514);
and U22239 (N_22239,N_19058,N_21296);
and U22240 (N_22240,N_20498,N_21266);
nand U22241 (N_22241,N_20236,N_19867);
or U22242 (N_22242,N_19207,N_19516);
nor U22243 (N_22243,N_21346,N_20478);
nor U22244 (N_22244,N_20055,N_20002);
and U22245 (N_22245,N_20099,N_21664);
and U22246 (N_22246,N_19192,N_21429);
or U22247 (N_22247,N_20365,N_19066);
nor U22248 (N_22248,N_21789,N_21371);
or U22249 (N_22249,N_21456,N_21655);
xor U22250 (N_22250,N_20562,N_19734);
xnor U22251 (N_22251,N_21184,N_19011);
xnor U22252 (N_22252,N_20118,N_20574);
nor U22253 (N_22253,N_19771,N_20313);
nand U22254 (N_22254,N_20318,N_19635);
nor U22255 (N_22255,N_19594,N_20777);
nor U22256 (N_22256,N_21243,N_19909);
xnor U22257 (N_22257,N_21520,N_19128);
nor U22258 (N_22258,N_21724,N_20104);
xor U22259 (N_22259,N_20979,N_20886);
nor U22260 (N_22260,N_21788,N_21041);
or U22261 (N_22261,N_18891,N_21065);
and U22262 (N_22262,N_20792,N_19148);
or U22263 (N_22263,N_20061,N_20691);
or U22264 (N_22264,N_21362,N_20753);
or U22265 (N_22265,N_21341,N_20709);
nor U22266 (N_22266,N_21135,N_20487);
nor U22267 (N_22267,N_19449,N_20733);
and U22268 (N_22268,N_21663,N_19228);
nor U22269 (N_22269,N_19807,N_19174);
or U22270 (N_22270,N_20346,N_19191);
and U22271 (N_22271,N_20668,N_19306);
nand U22272 (N_22272,N_20561,N_19798);
or U22273 (N_22273,N_18982,N_19610);
and U22274 (N_22274,N_20849,N_21660);
and U22275 (N_22275,N_21002,N_20069);
or U22276 (N_22276,N_18864,N_20011);
and U22277 (N_22277,N_18787,N_19373);
nand U22278 (N_22278,N_21268,N_21101);
or U22279 (N_22279,N_20439,N_19034);
nand U22280 (N_22280,N_21714,N_20534);
nor U22281 (N_22281,N_20366,N_19897);
nand U22282 (N_22282,N_21284,N_20195);
and U22283 (N_22283,N_20533,N_20896);
or U22284 (N_22284,N_19046,N_19997);
nor U22285 (N_22285,N_21576,N_19134);
nor U22286 (N_22286,N_19276,N_19504);
xnor U22287 (N_22287,N_19520,N_19593);
xor U22288 (N_22288,N_21051,N_20335);
and U22289 (N_22289,N_20155,N_21772);
nor U22290 (N_22290,N_19617,N_21629);
nor U22291 (N_22291,N_20665,N_19417);
or U22292 (N_22292,N_21829,N_20952);
or U22293 (N_22293,N_20509,N_19485);
or U22294 (N_22294,N_19025,N_20013);
or U22295 (N_22295,N_18791,N_21546);
and U22296 (N_22296,N_21249,N_19937);
and U22297 (N_22297,N_21739,N_21119);
and U22298 (N_22298,N_19014,N_21211);
nand U22299 (N_22299,N_20490,N_21611);
and U22300 (N_22300,N_19116,N_19583);
and U22301 (N_22301,N_19585,N_19431);
nand U22302 (N_22302,N_21124,N_20671);
or U22303 (N_22303,N_19038,N_19544);
nor U22304 (N_22304,N_19579,N_19991);
nand U22305 (N_22305,N_20859,N_20189);
nand U22306 (N_22306,N_19125,N_20276);
and U22307 (N_22307,N_21183,N_19633);
xor U22308 (N_22308,N_18939,N_19896);
and U22309 (N_22309,N_21155,N_20051);
and U22310 (N_22310,N_19566,N_20494);
nand U22311 (N_22311,N_21509,N_20455);
xor U22312 (N_22312,N_19295,N_19751);
or U22313 (N_22313,N_19698,N_21742);
nor U22314 (N_22314,N_21100,N_20719);
nand U22315 (N_22315,N_21423,N_19108);
nor U22316 (N_22316,N_21708,N_20610);
or U22317 (N_22317,N_20392,N_19210);
xor U22318 (N_22318,N_20934,N_21652);
or U22319 (N_22319,N_21628,N_21202);
nor U22320 (N_22320,N_21232,N_21759);
and U22321 (N_22321,N_21866,N_19558);
or U22322 (N_22322,N_18970,N_21798);
nor U22323 (N_22323,N_20997,N_19083);
or U22324 (N_22324,N_18772,N_21573);
xnor U22325 (N_22325,N_20992,N_19682);
nor U22326 (N_22326,N_21757,N_21309);
or U22327 (N_22327,N_20129,N_19040);
nand U22328 (N_22328,N_21482,N_21289);
or U22329 (N_22329,N_21805,N_20463);
nand U22330 (N_22330,N_21764,N_19671);
nor U22331 (N_22331,N_19708,N_18938);
and U22332 (N_22332,N_19761,N_21673);
and U22333 (N_22333,N_20415,N_20059);
xor U22334 (N_22334,N_19331,N_21510);
xnor U22335 (N_22335,N_20721,N_19865);
and U22336 (N_22336,N_21599,N_21021);
nand U22337 (N_22337,N_19401,N_19905);
nor U22338 (N_22338,N_19654,N_21074);
nor U22339 (N_22339,N_21730,N_19327);
nand U22340 (N_22340,N_21088,N_21706);
xnor U22341 (N_22341,N_19841,N_21011);
or U22342 (N_22342,N_21270,N_20967);
and U22343 (N_22343,N_19655,N_21125);
or U22344 (N_22344,N_20065,N_20611);
nor U22345 (N_22345,N_20842,N_21535);
and U22346 (N_22346,N_19533,N_19462);
or U22347 (N_22347,N_20397,N_19135);
xor U22348 (N_22348,N_21635,N_19639);
and U22349 (N_22349,N_21318,N_20248);
or U22350 (N_22350,N_21107,N_20955);
and U22351 (N_22351,N_21649,N_19960);
nor U22352 (N_22352,N_18761,N_19930);
xor U22353 (N_22353,N_20556,N_21242);
nand U22354 (N_22354,N_20742,N_21054);
or U22355 (N_22355,N_21549,N_21003);
nor U22356 (N_22356,N_18880,N_19219);
or U22357 (N_22357,N_21735,N_20409);
nand U22358 (N_22358,N_19601,N_18793);
nand U22359 (N_22359,N_20700,N_20705);
or U22360 (N_22360,N_19876,N_20172);
nor U22361 (N_22361,N_20696,N_19839);
nand U22362 (N_22362,N_18916,N_19854);
nand U22363 (N_22363,N_18788,N_19899);
or U22364 (N_22364,N_19194,N_18827);
or U22365 (N_22365,N_21776,N_19574);
or U22366 (N_22366,N_20756,N_20832);
or U22367 (N_22367,N_21530,N_19816);
or U22368 (N_22368,N_19543,N_21797);
xor U22369 (N_22369,N_19958,N_21279);
or U22370 (N_22370,N_19578,N_21497);
and U22371 (N_22371,N_19044,N_20200);
xor U22372 (N_22372,N_20861,N_18925);
or U22373 (N_22373,N_21203,N_20524);
or U22374 (N_22374,N_21354,N_21567);
nor U22375 (N_22375,N_19856,N_20722);
xnor U22376 (N_22376,N_19039,N_20996);
or U22377 (N_22377,N_20784,N_20146);
or U22378 (N_22378,N_20947,N_18765);
and U22379 (N_22379,N_20477,N_20208);
or U22380 (N_22380,N_19337,N_18826);
nor U22381 (N_22381,N_21096,N_19490);
or U22382 (N_22382,N_20250,N_21000);
nand U22383 (N_22383,N_20988,N_20355);
nor U22384 (N_22384,N_19834,N_18798);
nand U22385 (N_22385,N_19894,N_20530);
nor U22386 (N_22386,N_19928,N_21367);
nor U22387 (N_22387,N_19317,N_21381);
or U22388 (N_22388,N_19061,N_20245);
nor U22389 (N_22389,N_19589,N_20256);
and U22390 (N_22390,N_19127,N_20377);
nand U22391 (N_22391,N_20882,N_20937);
or U22392 (N_22392,N_20559,N_20905);
nand U22393 (N_22393,N_19952,N_19464);
or U22394 (N_22394,N_20426,N_20661);
or U22395 (N_22395,N_20892,N_18965);
nand U22396 (N_22396,N_21210,N_21813);
or U22397 (N_22397,N_21555,N_21335);
nand U22398 (N_22398,N_19394,N_20282);
nor U22399 (N_22399,N_20289,N_21138);
nand U22400 (N_22400,N_21364,N_20555);
or U22401 (N_22401,N_20910,N_20904);
nand U22402 (N_22402,N_19744,N_19467);
and U22403 (N_22403,N_19432,N_19087);
or U22404 (N_22404,N_18882,N_20982);
nor U22405 (N_22405,N_19293,N_19016);
nor U22406 (N_22406,N_20689,N_19321);
nor U22407 (N_22407,N_19402,N_20626);
or U22408 (N_22408,N_19452,N_21719);
or U22409 (N_22409,N_18875,N_21610);
or U22410 (N_22410,N_20015,N_19987);
nand U22411 (N_22411,N_21188,N_20893);
nand U22412 (N_22412,N_19107,N_21624);
nand U22413 (N_22413,N_19508,N_21486);
and U22414 (N_22414,N_20407,N_21079);
and U22415 (N_22415,N_20634,N_18986);
nor U22416 (N_22416,N_21824,N_19518);
nor U22417 (N_22417,N_20364,N_18908);
or U22418 (N_22418,N_20241,N_19634);
nand U22419 (N_22419,N_18754,N_20213);
nor U22420 (N_22420,N_19080,N_20606);
and U22421 (N_22421,N_20174,N_21662);
and U22422 (N_22422,N_19386,N_21661);
nor U22423 (N_22423,N_21276,N_21835);
and U22424 (N_22424,N_19000,N_19947);
nand U22425 (N_22425,N_19902,N_21393);
or U22426 (N_22426,N_20602,N_19454);
nand U22427 (N_22427,N_18941,N_21852);
or U22428 (N_22428,N_19962,N_19297);
and U22429 (N_22429,N_20273,N_20642);
or U22430 (N_22430,N_19077,N_20434);
and U22431 (N_22431,N_19209,N_20846);
or U22432 (N_22432,N_21044,N_21506);
and U22433 (N_22433,N_21062,N_19887);
xor U22434 (N_22434,N_21267,N_20680);
or U22435 (N_22435,N_19733,N_20096);
xor U22436 (N_22436,N_19666,N_21015);
nand U22437 (N_22437,N_19447,N_21578);
or U22438 (N_22438,N_19226,N_18797);
or U22439 (N_22439,N_19352,N_20932);
xor U22440 (N_22440,N_20086,N_19269);
nand U22441 (N_22441,N_20089,N_20963);
and U22442 (N_22442,N_21674,N_21275);
nand U22443 (N_22443,N_21027,N_19208);
nor U22444 (N_22444,N_21416,N_20765);
nor U22445 (N_22445,N_19256,N_20924);
nand U22446 (N_22446,N_19237,N_19515);
nor U22447 (N_22447,N_19780,N_21182);
and U22448 (N_22448,N_20314,N_21639);
nand U22449 (N_22449,N_20564,N_18989);
nor U22450 (N_22450,N_21331,N_20930);
or U22451 (N_22451,N_19860,N_21269);
and U22452 (N_22452,N_20504,N_19651);
or U22453 (N_22453,N_19348,N_19225);
nor U22454 (N_22454,N_18967,N_21521);
xor U22455 (N_22455,N_21844,N_21453);
xor U22456 (N_22456,N_21676,N_21861);
and U22457 (N_22457,N_20196,N_21737);
or U22458 (N_22458,N_19831,N_21667);
nand U22459 (N_22459,N_19383,N_19351);
or U22460 (N_22460,N_20396,N_19763);
or U22461 (N_22461,N_20877,N_21640);
and U22462 (N_22462,N_20502,N_21770);
or U22463 (N_22463,N_21111,N_21819);
and U22464 (N_22464,N_20684,N_20771);
and U22465 (N_22465,N_21856,N_20786);
nor U22466 (N_22466,N_21556,N_19347);
or U22467 (N_22467,N_20855,N_21066);
or U22468 (N_22468,N_21316,N_18942);
xnor U22469 (N_22469,N_21013,N_19955);
or U22470 (N_22470,N_19009,N_20277);
or U22471 (N_22471,N_19642,N_21395);
or U22472 (N_22472,N_20237,N_21390);
nand U22473 (N_22473,N_20781,N_20679);
and U22474 (N_22474,N_19102,N_19641);
nand U22475 (N_22475,N_21834,N_19826);
and U22476 (N_22476,N_19442,N_21761);
and U22477 (N_22477,N_20941,N_19203);
nand U22478 (N_22478,N_19626,N_19315);
nor U22479 (N_22479,N_20635,N_21686);
nand U22480 (N_22480,N_20003,N_19998);
xor U22481 (N_22481,N_21024,N_19888);
nand U22482 (N_22482,N_20095,N_20068);
and U22483 (N_22483,N_19605,N_20785);
or U22484 (N_22484,N_21621,N_21830);
and U22485 (N_22485,N_19448,N_19906);
nand U22486 (N_22486,N_19196,N_19255);
and U22487 (N_22487,N_20966,N_21310);
nor U22488 (N_22488,N_19302,N_19181);
and U22489 (N_22489,N_18889,N_21748);
and U22490 (N_22490,N_20845,N_21733);
and U22491 (N_22491,N_20384,N_20773);
xnor U22492 (N_22492,N_19530,N_21251);
xor U22493 (N_22493,N_19879,N_20449);
and U22494 (N_22494,N_20309,N_19463);
nand U22495 (N_22495,N_21178,N_19032);
and U22496 (N_22496,N_21372,N_19206);
nand U22497 (N_22497,N_19700,N_19772);
xnor U22498 (N_22498,N_19311,N_21173);
nand U22499 (N_22499,N_20333,N_21483);
nand U22500 (N_22500,N_19049,N_19663);
and U22501 (N_22501,N_18926,N_19387);
nor U22502 (N_22502,N_19157,N_21052);
or U22503 (N_22503,N_18892,N_20531);
or U22504 (N_22504,N_20412,N_20523);
nand U22505 (N_22505,N_20975,N_18948);
nand U22506 (N_22506,N_21191,N_20969);
and U22507 (N_22507,N_20539,N_19821);
nor U22508 (N_22508,N_20547,N_21281);
and U22509 (N_22509,N_19827,N_21817);
nand U22510 (N_22510,N_20600,N_20752);
or U22511 (N_22511,N_20049,N_19546);
nor U22512 (N_22512,N_20462,N_19480);
and U22513 (N_22513,N_21245,N_21644);
or U22514 (N_22514,N_19597,N_19716);
nand U22515 (N_22515,N_20116,N_19501);
nand U22516 (N_22516,N_18850,N_19972);
or U22517 (N_22517,N_21046,N_21669);
nor U22518 (N_22518,N_20092,N_21154);
or U22519 (N_22519,N_20727,N_20297);
nand U22520 (N_22520,N_18886,N_18750);
nor U22521 (N_22521,N_20983,N_21462);
and U22522 (N_22522,N_18988,N_20998);
and U22523 (N_22523,N_19817,N_19117);
nor U22524 (N_22524,N_21710,N_20831);
and U22525 (N_22525,N_21204,N_19725);
and U22526 (N_22526,N_19820,N_21023);
or U22527 (N_22527,N_20398,N_19536);
or U22528 (N_22528,N_19190,N_20287);
nand U22529 (N_22529,N_21828,N_20693);
and U22530 (N_22530,N_19470,N_21465);
and U22531 (N_22531,N_21687,N_19572);
xor U22532 (N_22532,N_19683,N_20815);
or U22533 (N_22533,N_20789,N_21215);
or U22534 (N_22534,N_21608,N_21418);
nand U22535 (N_22535,N_21803,N_20685);
and U22536 (N_22536,N_20316,N_19685);
nor U22537 (N_22537,N_19565,N_19884);
nor U22538 (N_22538,N_21006,N_18885);
nor U22539 (N_22539,N_21812,N_19272);
xor U22540 (N_22540,N_20080,N_18830);
nor U22541 (N_22541,N_21323,N_21185);
or U22542 (N_22542,N_20091,N_18768);
nor U22543 (N_22543,N_20431,N_19910);
nand U22544 (N_22544,N_20028,N_20769);
nand U22545 (N_22545,N_19259,N_21145);
or U22546 (N_22546,N_18870,N_19730);
and U22547 (N_22547,N_20703,N_20387);
or U22548 (N_22548,N_19853,N_19388);
xnor U22549 (N_22549,N_21399,N_19123);
nand U22550 (N_22550,N_21563,N_18824);
nand U22551 (N_22551,N_21009,N_21538);
and U22552 (N_22552,N_20622,N_20052);
or U22553 (N_22553,N_21262,N_21678);
xnor U22554 (N_22554,N_21165,N_19562);
nand U22555 (N_22555,N_21619,N_20801);
or U22556 (N_22556,N_21472,N_20170);
and U22557 (N_22557,N_19554,N_19130);
nand U22558 (N_22558,N_18964,N_21420);
nand U22559 (N_22559,N_20370,N_21675);
and U22560 (N_22560,N_19419,N_19260);
nor U22561 (N_22561,N_19155,N_20408);
nor U22562 (N_22562,N_21127,N_21448);
nor U22563 (N_22563,N_20926,N_21132);
nor U22564 (N_22564,N_19548,N_20652);
nor U22565 (N_22565,N_19224,N_20873);
and U22566 (N_22566,N_21575,N_19680);
and U22567 (N_22567,N_19672,N_21810);
nor U22568 (N_22568,N_19560,N_20970);
nand U22569 (N_22569,N_20973,N_19777);
nand U22570 (N_22570,N_20885,N_20162);
and U22571 (N_22571,N_19008,N_19891);
nand U22572 (N_22572,N_20321,N_20959);
xnor U22573 (N_22573,N_18962,N_21086);
and U22574 (N_22574,N_18944,N_21605);
and U22575 (N_22575,N_19473,N_19737);
and U22576 (N_22576,N_19645,N_21158);
xnor U22577 (N_22577,N_20888,N_20536);
and U22578 (N_22578,N_19197,N_19781);
and U22579 (N_22579,N_20677,N_20759);
and U22580 (N_22580,N_20878,N_19020);
or U22581 (N_22581,N_19555,N_19037);
xor U22582 (N_22582,N_21857,N_19863);
nand U22583 (N_22583,N_19497,N_20036);
xnor U22584 (N_22584,N_18865,N_19801);
or U22585 (N_22585,N_20840,N_20508);
and U22586 (N_22586,N_19330,N_20862);
or U22587 (N_22587,N_19659,N_19502);
nor U22588 (N_22588,N_19794,N_21380);
or U22589 (N_22589,N_20757,N_21545);
nor U22590 (N_22590,N_19969,N_21059);
and U22591 (N_22591,N_19979,N_21559);
or U22592 (N_22592,N_19489,N_19967);
nor U22593 (N_22593,N_21257,N_19422);
xnor U22594 (N_22594,N_18823,N_21014);
nor U22595 (N_22595,N_20552,N_19142);
and U22596 (N_22596,N_21007,N_21593);
nor U22597 (N_22597,N_21825,N_20193);
and U22598 (N_22598,N_18854,N_21282);
nand U22599 (N_22599,N_21439,N_19965);
or U22600 (N_22600,N_21870,N_19092);
or U22601 (N_22601,N_19726,N_18840);
nor U22602 (N_22602,N_18995,N_21839);
and U22603 (N_22603,N_20201,N_20075);
or U22604 (N_22604,N_21313,N_19673);
and U22605 (N_22605,N_20066,N_19961);
or U22606 (N_22606,N_18874,N_19369);
and U22607 (N_22607,N_21033,N_19944);
or U22608 (N_22608,N_19795,N_20067);
nor U22609 (N_22609,N_19776,N_18811);
and U22610 (N_22610,N_21791,N_19391);
and U22611 (N_22611,N_21141,N_21159);
and U22612 (N_22612,N_20820,N_19294);
nand U22613 (N_22613,N_21597,N_19915);
nand U22614 (N_22614,N_19679,N_19101);
nand U22615 (N_22615,N_21613,N_19248);
and U22616 (N_22616,N_20204,N_21128);
xor U22617 (N_22617,N_21565,N_21256);
and U22618 (N_22618,N_19420,N_19893);
nor U22619 (N_22619,N_21301,N_19974);
nand U22620 (N_22620,N_19081,N_20168);
and U22621 (N_22621,N_19021,N_20042);
or U22622 (N_22622,N_21726,N_20864);
nor U22623 (N_22623,N_21189,N_20163);
and U22624 (N_22624,N_21069,N_21572);
nor U22625 (N_22625,N_19778,N_20484);
nor U22626 (N_22626,N_21574,N_20741);
nand U22627 (N_22627,N_20902,N_21528);
xnor U22628 (N_22628,N_19684,N_19736);
nand U22629 (N_22629,N_20620,N_19229);
or U22630 (N_22630,N_19160,N_21725);
or U22631 (N_22631,N_18876,N_19318);
nor U22632 (N_22632,N_20553,N_19538);
or U22633 (N_22633,N_20159,N_20338);
and U22634 (N_22634,N_19356,N_18959);
nand U22635 (N_22635,N_20070,N_18949);
nor U22636 (N_22636,N_21762,N_21047);
and U22637 (N_22637,N_19172,N_20920);
and U22638 (N_22638,N_21507,N_20687);
nand U22639 (N_22639,N_19184,N_20944);
and U22640 (N_22640,N_20702,N_21840);
nand U22641 (N_22641,N_19287,N_19903);
nand U22642 (N_22642,N_21305,N_19917);
nor U22643 (N_22643,N_20274,N_21821);
xnor U22644 (N_22644,N_21832,N_20609);
and U22645 (N_22645,N_21190,N_19904);
xor U22646 (N_22646,N_20098,N_21755);
and U22647 (N_22647,N_18817,N_21327);
or U22648 (N_22648,N_20234,N_19625);
nor U22649 (N_22649,N_21218,N_18807);
and U22650 (N_22650,N_19785,N_20166);
nand U22651 (N_22651,N_20607,N_20678);
and U22652 (N_22652,N_21585,N_21478);
and U22653 (N_22653,N_19173,N_20233);
or U22654 (N_22654,N_20653,N_19943);
nand U22655 (N_22655,N_20133,N_20540);
or U22656 (N_22656,N_19596,N_21382);
nand U22657 (N_22657,N_20043,N_19760);
nand U22658 (N_22658,N_21786,N_18785);
or U22659 (N_22659,N_19837,N_20294);
nor U22660 (N_22660,N_19656,N_20342);
nand U22661 (N_22661,N_19090,N_20743);
or U22662 (N_22662,N_19951,N_21034);
and U22663 (N_22663,N_20150,N_21026);
or U22664 (N_22664,N_20257,N_19271);
and U22665 (N_22665,N_19283,N_21058);
and U22666 (N_22666,N_20386,N_19093);
xor U22667 (N_22667,N_19806,N_19541);
or U22668 (N_22668,N_20324,N_19788);
or U22669 (N_22669,N_21721,N_20636);
or U22670 (N_22670,N_18778,N_20802);
nor U22671 (N_22671,N_18987,N_21224);
nor U22672 (N_22672,N_20697,N_18915);
and U22673 (N_22673,N_20656,N_21515);
and U22674 (N_22674,N_20797,N_21068);
nor U22675 (N_22675,N_18767,N_20410);
and U22676 (N_22676,N_21688,N_20472);
nor U22677 (N_22677,N_20369,N_20097);
or U22678 (N_22678,N_21219,N_20078);
and U22679 (N_22679,N_19667,N_19740);
or U22680 (N_22680,N_20401,N_20779);
and U22681 (N_22681,N_21402,N_20594);
and U22682 (N_22682,N_19471,N_20682);
xnor U22683 (N_22683,N_20728,N_18917);
nand U22684 (N_22684,N_20102,N_21616);
nand U22685 (N_22685,N_20315,N_21490);
nor U22686 (N_22686,N_18816,N_19975);
or U22687 (N_22687,N_19525,N_20667);
nor U22688 (N_22688,N_19992,N_20071);
nand U22689 (N_22689,N_21845,N_19263);
xor U22690 (N_22690,N_19723,N_18933);
and U22691 (N_22691,N_19665,N_21018);
and U22692 (N_22692,N_21529,N_19060);
and U22693 (N_22693,N_19274,N_20940);
and U22694 (N_22694,N_21604,N_19067);
nor U22695 (N_22695,N_20220,N_20486);
nand U22696 (N_22696,N_19035,N_19786);
nor U22697 (N_22697,N_19907,N_20758);
and U22698 (N_22698,N_18852,N_21853);
nand U22699 (N_22699,N_19569,N_19115);
nor U22700 (N_22700,N_21102,N_21534);
or U22701 (N_22701,N_18836,N_20139);
or U22702 (N_22702,N_21095,N_18999);
nand U22703 (N_22703,N_21053,N_20079);
or U22704 (N_22704,N_18756,N_21569);
nor U22705 (N_22705,N_18789,N_19668);
and U22706 (N_22706,N_19586,N_20535);
xnor U22707 (N_22707,N_19836,N_18764);
nand U22708 (N_22708,N_19368,N_19324);
and U22709 (N_22709,N_20421,N_19098);
or U22710 (N_22710,N_19236,N_20746);
nand U22711 (N_22711,N_19517,N_20126);
or U22712 (N_22712,N_21087,N_18860);
nor U22713 (N_22713,N_19162,N_18923);
and U22714 (N_22714,N_21842,N_19078);
nor U22715 (N_22715,N_21386,N_19089);
nand U22716 (N_22716,N_19846,N_20125);
or U22717 (N_22717,N_20443,N_20259);
nand U22718 (N_22718,N_21498,N_19886);
xnor U22719 (N_22719,N_19553,N_19675);
and U22720 (N_22720,N_19189,N_19724);
nor U22721 (N_22721,N_20578,N_19731);
nor U22722 (N_22722,N_20515,N_21473);
nand U22723 (N_22723,N_19377,N_19418);
nor U22724 (N_22724,N_18929,N_20331);
nor U22725 (N_22725,N_18943,N_19644);
nand U22726 (N_22726,N_20628,N_21512);
xnor U22727 (N_22727,N_21240,N_19275);
or U22728 (N_22728,N_18900,N_20390);
nand U22729 (N_22729,N_20565,N_21363);
nor U22730 (N_22730,N_20576,N_20244);
nand U22731 (N_22731,N_19180,N_20215);
nor U22732 (N_22732,N_19096,N_20631);
or U22733 (N_22733,N_19996,N_20444);
nor U22734 (N_22734,N_21562,N_20745);
or U22735 (N_22735,N_20852,N_20411);
or U22736 (N_22736,N_21117,N_21622);
and U22737 (N_22737,N_19757,N_21769);
xnor U22738 (N_22738,N_20275,N_20776);
and U22739 (N_22739,N_20152,N_18781);
xnor U22740 (N_22740,N_19499,N_20114);
and U22741 (N_22741,N_20629,N_19277);
nand U22742 (N_22742,N_19220,N_20253);
xnor U22743 (N_22743,N_21837,N_19883);
and U22744 (N_22744,N_19920,N_19812);
nor U22745 (N_22745,N_20417,N_20584);
or U22746 (N_22746,N_20778,N_21648);
nand U22747 (N_22747,N_21142,N_20038);
nand U22748 (N_22748,N_21440,N_21077);
nor U22749 (N_22749,N_20747,N_20340);
nand U22750 (N_22750,N_21349,N_21300);
nor U22751 (N_22751,N_20605,N_20681);
and U22752 (N_22752,N_19702,N_19743);
or U22753 (N_22753,N_21376,N_19104);
nor U22754 (N_22754,N_20805,N_20927);
and U22755 (N_22755,N_19779,N_20308);
and U22756 (N_22756,N_21740,N_20587);
and U22757 (N_22757,N_21343,N_21860);
nand U22758 (N_22758,N_21149,N_18979);
nor U22759 (N_22759,N_19137,N_19429);
or U22760 (N_22760,N_19027,N_21001);
xnor U22761 (N_22761,N_21286,N_18800);
and U22762 (N_22762,N_19980,N_21863);
and U22763 (N_22763,N_18899,N_21480);
or U22764 (N_22764,N_20060,N_19603);
nand U22765 (N_22765,N_21540,N_19468);
nor U22766 (N_22766,N_20657,N_20476);
and U22767 (N_22767,N_19436,N_19649);
xnor U22768 (N_22768,N_19519,N_20483);
or U22769 (N_22769,N_19268,N_21230);
xor U22770 (N_22770,N_18906,N_18934);
or U22771 (N_22771,N_18931,N_20868);
and U22772 (N_22772,N_20599,N_19308);
or U22773 (N_22773,N_19595,N_19458);
or U22774 (N_22774,N_21365,N_20012);
xnor U22775 (N_22775,N_18977,N_19216);
nand U22776 (N_22776,N_19914,N_19505);
or U22777 (N_22777,N_20581,N_21684);
xnor U22778 (N_22778,N_20596,N_21484);
or U22779 (N_22779,N_21144,N_19949);
xnor U22780 (N_22780,N_20328,N_19898);
nand U22781 (N_22781,N_19852,N_21446);
or U22782 (N_22782,N_18752,N_19687);
or U22783 (N_22783,N_18783,N_21246);
and U22784 (N_22784,N_20811,N_18843);
nor U22785 (N_22785,N_20142,N_19033);
and U22786 (N_22786,N_19933,N_21194);
or U22787 (N_22787,N_20922,N_20714);
or U22788 (N_22788,N_19186,N_20224);
and U22789 (N_22789,N_18956,N_19407);
and U22790 (N_22790,N_19408,N_20130);
nand U22791 (N_22791,N_19759,N_18985);
or U22792 (N_22792,N_20192,N_20521);
nor U22793 (N_22793,N_19143,N_19164);
nand U22794 (N_22794,N_21502,N_20100);
nor U22795 (N_22795,N_21201,N_18919);
nor U22796 (N_22796,N_19221,N_21137);
nand U22797 (N_22797,N_21547,N_21715);
nand U22798 (N_22798,N_21850,N_19819);
nand U22799 (N_22799,N_20891,N_20615);
nand U22800 (N_22800,N_18904,N_18801);
and U22801 (N_22801,N_20264,N_20300);
nand U22802 (N_22802,N_20064,N_21340);
or U22803 (N_22803,N_20286,N_19791);
and U22804 (N_22804,N_19455,N_21615);
and U22805 (N_22805,N_18819,N_20951);
nor U22806 (N_22806,N_20281,N_21777);
xor U22807 (N_22807,N_21633,N_21815);
nor U22808 (N_22808,N_20179,N_21872);
xor U22809 (N_22809,N_20732,N_20999);
nor U22810 (N_22810,N_19074,N_20577);
or U22811 (N_22811,N_19895,N_20543);
and U22812 (N_22812,N_18910,N_19935);
or U22813 (N_22813,N_19908,N_20351);
or U22814 (N_22814,N_21248,N_21105);
and U22815 (N_22815,N_19669,N_19257);
or U22816 (N_22816,N_20413,N_19630);
and U22817 (N_22817,N_19006,N_19956);
and U22818 (N_22818,N_18803,N_21379);
nor U22819 (N_22819,N_18966,N_19697);
nor U22820 (N_22820,N_19177,N_20990);
nand U22821 (N_22821,N_18971,N_20354);
nor U22822 (N_22822,N_20207,N_21334);
or U22823 (N_22823,N_19804,N_21106);
or U22824 (N_22824,N_20210,N_18829);
nor U22825 (N_22825,N_21170,N_19838);
nand U22826 (N_22826,N_21168,N_21504);
and U22827 (N_22827,N_20279,N_20363);
nand U22828 (N_22828,N_20285,N_20601);
nor U22829 (N_22829,N_20489,N_19484);
or U22830 (N_22830,N_20738,N_19299);
nor U22831 (N_22831,N_19273,N_19424);
and U22832 (N_22832,N_20094,N_20589);
or U22833 (N_22833,N_21862,N_21325);
nand U22834 (N_22834,N_19261,N_20850);
nand U22835 (N_22835,N_20278,N_20173);
or U22836 (N_22836,N_19064,N_18838);
nor U22837 (N_22837,N_20715,N_21252);
nor U22838 (N_22838,N_20374,N_20107);
nor U22839 (N_22839,N_20045,N_20567);
or U22840 (N_22840,N_20212,N_21617);
nor U22841 (N_22841,N_19602,N_18796);
and U22842 (N_22842,N_19835,N_18954);
nand U22843 (N_22843,N_20307,N_19570);
or U22844 (N_22844,N_19379,N_20268);
nand U22845 (N_22845,N_19549,N_19346);
nand U22846 (N_22846,N_21208,N_20572);
nor U22847 (N_22847,N_19981,N_20804);
nand U22848 (N_22848,N_19265,N_21864);
nor U22849 (N_22849,N_21304,N_19341);
xor U22850 (N_22850,N_20866,N_21801);
nand U22851 (N_22851,N_19818,N_19990);
nand U22852 (N_22852,N_18845,N_20334);
nand U22853 (N_22853,N_19963,N_19717);
and U22854 (N_22854,N_21838,N_19103);
xnor U22855 (N_22855,N_21283,N_20044);
or U22856 (N_22856,N_20880,N_21295);
or U22857 (N_22857,N_21432,N_20736);
or U22858 (N_22858,N_21264,N_19532);
and U22859 (N_22859,N_21614,N_19382);
nor U22860 (N_22860,N_18961,N_21641);
or U22861 (N_22861,N_21671,N_20323);
and U22862 (N_22862,N_19580,N_19430);
nand U22863 (N_22863,N_20871,N_19957);
or U22864 (N_22864,N_20093,N_20787);
nor U22865 (N_22865,N_20029,N_18905);
and U22866 (N_22866,N_20551,N_20847);
and U22867 (N_22867,N_20056,N_19343);
nand U22868 (N_22868,N_19133,N_20032);
nand U22869 (N_22869,N_20974,N_19758);
and U22870 (N_22870,N_21221,N_20851);
nor U22871 (N_22871,N_20995,N_20641);
nor U22872 (N_22872,N_20624,N_21794);
and U22873 (N_22873,N_21550,N_20813);
or U22874 (N_22874,N_21445,N_20372);
xnor U22875 (N_22875,N_21311,N_20325);
or U22876 (N_22876,N_20448,N_21455);
nand U22877 (N_22877,N_20157,N_18751);
nand U22878 (N_22878,N_19076,N_20475);
nor U22879 (N_22879,N_19840,N_20453);
nor U22880 (N_22880,N_21691,N_20633);
nor U22881 (N_22881,N_20187,N_19176);
or U22882 (N_22882,N_18909,N_19792);
nand U22883 (N_22883,N_21612,N_19705);
nand U22884 (N_22884,N_21206,N_18969);
and U22885 (N_22885,N_21851,N_18810);
nor U22886 (N_22886,N_19984,N_20881);
and U22887 (N_22887,N_20782,N_21517);
nor U22888 (N_22888,N_20972,N_21727);
or U22889 (N_22889,N_19729,N_21492);
and U22890 (N_22890,N_19588,N_19650);
and U22891 (N_22891,N_19397,N_18762);
nor U22892 (N_22892,N_20994,N_20216);
nand U22893 (N_22893,N_19735,N_21039);
or U22894 (N_22894,N_21584,N_21690);
nor U22895 (N_22895,N_20336,N_20614);
or U22896 (N_22896,N_20406,N_20643);
nand U22897 (N_22897,N_19754,N_20549);
and U22898 (N_22898,N_18972,N_19769);
and U22899 (N_22899,N_18856,N_21849);
nor U22900 (N_22900,N_20347,N_20803);
or U22901 (N_22901,N_19715,N_19755);
nor U22902 (N_22902,N_20654,N_18980);
or U22903 (N_22903,N_20404,N_19057);
xor U22904 (N_22904,N_21338,N_21499);
nor U22905 (N_22905,N_19738,N_18820);
or U22906 (N_22906,N_21063,N_20219);
nor U22907 (N_22907,N_20385,N_21298);
and U22908 (N_22908,N_19483,N_18992);
nor U22909 (N_22909,N_19970,N_21143);
or U22910 (N_22910,N_19995,N_20040);
and U22911 (N_22911,N_19052,N_21035);
nor U22912 (N_22912,N_20240,N_18927);
or U22913 (N_22913,N_20875,N_21626);
nor U22914 (N_22914,N_18771,N_19258);
xnor U22915 (N_22915,N_20542,N_18936);
nor U22916 (N_22916,N_21359,N_20510);
nor U22917 (N_22917,N_20014,N_20814);
and U22918 (N_22918,N_20054,N_21775);
or U22919 (N_22919,N_20856,N_21778);
or U22920 (N_22920,N_19375,N_19750);
and U22921 (N_22921,N_19227,N_19537);
nand U22922 (N_22922,N_21129,N_20356);
nor U22923 (N_22923,N_21385,N_20659);
nand U22924 (N_22924,N_21508,N_20311);
nand U22925 (N_22925,N_20912,N_20664);
or U22926 (N_22926,N_19316,N_19332);
nor U22927 (N_22927,N_20041,N_18997);
or U22928 (N_22928,N_19230,N_18993);
and U22929 (N_22929,N_21464,N_19494);
xor U22930 (N_22930,N_21553,N_20322);
nand U22931 (N_22931,N_19811,N_19372);
nor U22932 (N_22932,N_20945,N_19187);
and U22933 (N_22933,N_21422,N_20707);
or U22934 (N_22934,N_19359,N_20371);
nand U22935 (N_22935,N_18805,N_21697);
nand U22936 (N_22936,N_20007,N_20793);
or U22937 (N_22937,N_19266,N_18855);
and U22938 (N_22938,N_20247,N_20121);
or U22939 (N_22939,N_18981,N_21192);
nand U22940 (N_22940,N_19149,N_20748);
nand U22941 (N_22941,N_20981,N_20383);
nand U22942 (N_22942,N_21017,N_21356);
and U22943 (N_22943,N_19335,N_19493);
nand U22944 (N_22944,N_21489,N_21016);
or U22945 (N_22945,N_19885,N_19072);
and U22946 (N_22946,N_18914,N_19746);
nand U22947 (N_22947,N_21743,N_21005);
and U22948 (N_22948,N_21447,N_18877);
or U22949 (N_22949,N_19362,N_19433);
or U22950 (N_22950,N_20481,N_19428);
and U22951 (N_22951,N_19799,N_18806);
and U22952 (N_22952,N_21317,N_21040);
nor U22953 (N_22953,N_19380,N_19050);
xnor U22954 (N_22954,N_21752,N_21598);
nand U22955 (N_22955,N_21700,N_19813);
nor U22956 (N_22956,N_19941,N_19977);
and U22957 (N_22957,N_19264,N_20724);
nor U22958 (N_22958,N_19438,N_21477);
or U22959 (N_22959,N_20303,N_21458);
and U22960 (N_22960,N_19728,N_21848);
nand U22961 (N_22961,N_19732,N_20514);
and U22962 (N_22962,N_20178,N_19756);
nand U22963 (N_22963,N_21665,N_19875);
nand U22964 (N_22964,N_20149,N_21330);
and U22965 (N_22965,N_20190,N_20304);
or U22966 (N_22966,N_21324,N_20718);
nand U22967 (N_22967,N_21179,N_20537);
nand U22968 (N_22968,N_21683,N_18960);
or U22969 (N_22969,N_20047,N_19292);
and U22970 (N_22970,N_21741,N_19767);
or U22971 (N_22971,N_19389,N_21205);
or U22972 (N_22972,N_19849,N_21685);
nor U22973 (N_22973,N_19647,N_21374);
nor U22974 (N_22974,N_19253,N_18912);
or U22975 (N_22975,N_18921,N_21656);
nand U22976 (N_22976,N_21360,N_20887);
or U22977 (N_22977,N_19540,N_20447);
and U22978 (N_22978,N_19978,N_20442);
xnor U22979 (N_22979,N_21260,N_19652);
nor U22980 (N_22980,N_20009,N_21285);
or U22981 (N_22981,N_21668,N_21527);
or U22982 (N_22982,N_19999,N_21254);
nand U22983 (N_22983,N_20991,N_20825);
and U22984 (N_22984,N_21060,N_19797);
or U22985 (N_22985,N_19762,N_20513);
nand U22986 (N_22986,N_18857,N_20260);
nand U22987 (N_22987,N_21514,N_19988);
or U22988 (N_22988,N_21036,N_21339);
and U22989 (N_22989,N_19313,N_20232);
nand U22990 (N_22990,N_20227,N_21056);
nor U22991 (N_22991,N_21526,N_21571);
or U22992 (N_22992,N_21522,N_18963);
or U22993 (N_22993,N_19513,N_21012);
and U22994 (N_22994,N_21496,N_20597);
or U22995 (N_22995,N_20433,N_20004);
and U22996 (N_22996,N_19848,N_18786);
nor U22997 (N_22997,N_20883,N_19068);
nor U22998 (N_22998,N_20772,N_21459);
nor U22999 (N_22999,N_20359,N_21537);
nor U23000 (N_23000,N_21010,N_19165);
nand U23001 (N_23001,N_21703,N_21443);
and U23002 (N_23002,N_21216,N_21320);
nand U23003 (N_23003,N_19823,N_21081);
or U23004 (N_23004,N_19427,N_19247);
nor U23005 (N_23005,N_21075,N_20550);
nand U23006 (N_23006,N_20712,N_19232);
and U23007 (N_23007,N_20783,N_21357);
nor U23008 (N_23008,N_19288,N_20182);
and U23009 (N_23009,N_21130,N_20560);
nor U23010 (N_23010,N_21855,N_21152);
or U23011 (N_23011,N_19880,N_21426);
and U23012 (N_23012,N_21787,N_19616);
or U23013 (N_23013,N_20948,N_20341);
or U23014 (N_23014,N_19023,N_20037);
nand U23015 (N_23015,N_19658,N_21050);
nand U23016 (N_23016,N_19393,N_19365);
nor U23017 (N_23017,N_19964,N_18853);
or U23018 (N_23018,N_20138,N_19718);
nor U23019 (N_23019,N_21716,N_21225);
xor U23020 (N_23020,N_21048,N_19280);
nand U23021 (N_23021,N_21322,N_20249);
and U23022 (N_23022,N_18790,N_20209);
nand U23023 (N_23023,N_19552,N_21580);
nor U23024 (N_23024,N_21091,N_21792);
xor U23025 (N_23025,N_20796,N_21579);
nor U23026 (N_23026,N_20836,N_21377);
nor U23027 (N_23027,N_20175,N_19802);
nand U23028 (N_23028,N_19587,N_18835);
or U23029 (N_23029,N_21541,N_19002);
nand U23030 (N_23030,N_19859,N_20423);
nor U23031 (N_23031,N_20147,N_20568);
and U23032 (N_23032,N_19202,N_20239);
and U23033 (N_23033,N_21732,N_20326);
or U23034 (N_23034,N_19132,N_19693);
xnor U23035 (N_23035,N_19234,N_18896);
xor U23036 (N_23036,N_21408,N_19144);
xnor U23037 (N_23037,N_21751,N_20437);
nor U23038 (N_23038,N_20598,N_19314);
nand U23039 (N_23039,N_20639,N_20918);
nor U23040 (N_23040,N_20222,N_20762);
and U23041 (N_23041,N_20939,N_21827);
xor U23042 (N_23042,N_21731,N_21193);
nor U23043 (N_23043,N_20135,N_20230);
nand U23044 (N_23044,N_20330,N_19400);
and U23045 (N_23045,N_21601,N_20242);
nor U23046 (N_23046,N_19304,N_21670);
and U23047 (N_23047,N_21121,N_19983);
or U23048 (N_23048,N_21650,N_21595);
or U23049 (N_23049,N_19599,N_20422);
nor U23050 (N_23050,N_20420,N_20393);
nor U23051 (N_23051,N_19492,N_19406);
and U23052 (N_23052,N_19613,N_20623);
nand U23053 (N_23053,N_19474,N_20818);
nand U23054 (N_23054,N_19619,N_19412);
nand U23055 (N_23055,N_18770,N_21022);
and U23056 (N_23056,N_20909,N_19201);
nor U23057 (N_23057,N_20424,N_20177);
nor U23058 (N_23058,N_21774,N_19015);
nor U23059 (N_23059,N_19550,N_20470);
nor U23060 (N_23060,N_19158,N_21793);
and U23061 (N_23061,N_19622,N_21278);
and U23062 (N_23062,N_19929,N_21720);
xnor U23063 (N_23063,N_21198,N_19878);
nor U23064 (N_23064,N_21373,N_20026);
and U23065 (N_23065,N_21226,N_21038);
nand U23066 (N_23066,N_20337,N_18918);
nand U23067 (N_23067,N_20113,N_19018);
and U23068 (N_23068,N_19384,N_20908);
and U23069 (N_23069,N_18841,N_18861);
and U23070 (N_23070,N_21136,N_20884);
nand U23071 (N_23071,N_21410,N_21434);
and U23072 (N_23072,N_20726,N_20456);
nand U23073 (N_23073,N_19510,N_20588);
or U23074 (N_23074,N_20081,N_20378);
nor U23075 (N_23075,N_20161,N_20181);
nor U23076 (N_23076,N_21516,N_20156);
or U23077 (N_23077,N_18994,N_18958);
nor U23078 (N_23078,N_21261,N_20088);
and U23079 (N_23079,N_19506,N_21551);
nand U23080 (N_23080,N_20332,N_20358);
and U23081 (N_23081,N_19163,N_20272);
or U23082 (N_23082,N_19704,N_20808);
or U23083 (N_23083,N_20485,N_19775);
nor U23084 (N_23084,N_20291,N_21098);
or U23085 (N_23085,N_19632,N_19053);
nand U23086 (N_23086,N_21823,N_19564);
or U23087 (N_23087,N_19710,N_21344);
nand U23088 (N_23088,N_21199,N_20111);
nand U23089 (N_23089,N_20843,N_20452);
and U23090 (N_23090,N_21738,N_18833);
and U23091 (N_23091,N_19105,N_21589);
and U23092 (N_23092,N_19085,N_21587);
and U23093 (N_23093,N_21594,N_19766);
nor U23094 (N_23094,N_21355,N_19199);
or U23095 (N_23095,N_20764,N_21476);
nand U23096 (N_23096,N_21437,N_18873);
nor U23097 (N_23097,N_20418,N_20950);
nand U23098 (N_23098,N_21294,N_19709);
xnor U23099 (N_23099,N_21020,N_20799);
or U23100 (N_23100,N_19790,N_20320);
and U23101 (N_23101,N_19808,N_21494);
or U23102 (N_23102,N_19703,N_18815);
nor U23103 (N_23103,N_21519,N_20019);
and U23104 (N_23104,N_20109,N_18782);
nor U23105 (N_23105,N_20024,N_19677);
or U23106 (N_23106,N_21479,N_20768);
nand U23107 (N_23107,N_20063,N_18831);
xor U23108 (N_23108,N_20817,N_21032);
nor U23109 (N_23109,N_21491,N_19289);
and U23110 (N_23110,N_21233,N_20164);
nor U23111 (N_23111,N_20821,N_20306);
nand U23112 (N_23112,N_18844,N_20731);
nand U23113 (N_23113,N_21167,N_20450);
xor U23114 (N_23114,N_18947,N_19707);
or U23115 (N_23115,N_20579,N_21753);
xnor U23116 (N_23116,N_19872,N_18862);
nor U23117 (N_23117,N_21064,N_21653);
or U23118 (N_23118,N_18890,N_19567);
and U23119 (N_23119,N_19976,N_19900);
or U23120 (N_23120,N_21347,N_18846);
or U23121 (N_23121,N_20459,N_20505);
nand U23122 (N_23122,N_19940,N_19374);
or U23123 (N_23123,N_21654,N_21293);
and U23124 (N_23124,N_21029,N_20429);
nor U23125 (N_23125,N_21750,N_20826);
nand U23126 (N_23126,N_20225,N_19857);
nand U23127 (N_23127,N_20357,N_20699);
nand U23128 (N_23128,N_19411,N_19609);
and U23129 (N_23129,N_21631,N_21195);
nor U23130 (N_23130,N_18898,N_21412);
and U23131 (N_23131,N_20430,N_21263);
or U23132 (N_23132,N_20928,N_19477);
and U23133 (N_23133,N_21333,N_21025);
nor U23134 (N_23134,N_19921,N_19354);
or U23135 (N_23135,N_19364,N_21414);
or U23136 (N_23136,N_19095,N_20946);
nand U23137 (N_23137,N_21582,N_21709);
xnor U23138 (N_23138,N_21151,N_19443);
xnor U23139 (N_23139,N_21166,N_21383);
and U23140 (N_23140,N_21638,N_20603);
xnor U23141 (N_23141,N_21452,N_19182);
or U23142 (N_23142,N_19404,N_18766);
nand U23143 (N_23143,N_20110,N_21319);
or U23144 (N_23144,N_19469,N_19692);
and U23145 (N_23145,N_21620,N_20964);
and U23146 (N_23146,N_21306,N_21229);
or U23147 (N_23147,N_21150,N_19303);
xnor U23148 (N_23148,N_20857,N_20903);
nand U23149 (N_23149,N_19871,N_20493);
or U23150 (N_23150,N_20468,N_20112);
nor U23151 (N_23151,N_20962,N_20349);
and U23152 (N_23152,N_20630,N_20627);
nor U23153 (N_23153,N_20191,N_19445);
xor U23154 (N_23154,N_20548,N_20141);
nand U23155 (N_23155,N_18968,N_19695);
nand U23156 (N_23156,N_20062,N_19966);
and U23157 (N_23157,N_19145,N_19686);
or U23158 (N_23158,N_20720,N_19300);
and U23159 (N_23159,N_19919,N_21228);
and U23160 (N_23160,N_19557,N_18757);
nand U23161 (N_23161,N_19007,N_19901);
xnor U23162 (N_23162,N_21767,N_19329);
xnor U23163 (N_23163,N_19047,N_20658);
or U23164 (N_23164,N_21396,N_21196);
or U23165 (N_23165,N_20734,N_20074);
nand U23166 (N_23166,N_20686,N_21118);
nand U23167 (N_23167,N_19250,N_20108);
or U23168 (N_23168,N_19660,N_19338);
xnor U23169 (N_23169,N_19305,N_20223);
nor U23170 (N_23170,N_19214,N_21696);
or U23171 (N_23171,N_20046,N_20529);
and U23172 (N_23172,N_21080,N_21394);
nand U23173 (N_23173,N_20806,N_20503);
and U23174 (N_23174,N_19681,N_21843);
or U23175 (N_23175,N_19939,N_20822);
nand U23176 (N_23176,N_21186,N_20134);
and U23177 (N_23177,N_21113,N_19097);
nor U23178 (N_23178,N_20120,N_20017);
nor U23179 (N_23179,N_19500,N_21288);
nor U23180 (N_23180,N_20301,N_20197);
and U23181 (N_23181,N_19309,N_21552);
nand U23182 (N_23182,N_20427,N_21609);
xnor U23183 (N_23183,N_19989,N_21328);
or U23184 (N_23184,N_20637,N_20416);
and U23185 (N_23185,N_19084,N_21809);
and U23186 (N_23186,N_21083,N_19789);
and U23187 (N_23187,N_20382,N_20522);
nor U23188 (N_23188,N_20361,N_21867);
and U23189 (N_23189,N_20495,N_21745);
nand U23190 (N_23190,N_20916,N_20949);
xnor U23191 (N_23191,N_18774,N_21672);
xor U23192 (N_23192,N_20710,N_20767);
nor U23193 (N_23193,N_19604,N_21718);
nand U23194 (N_23194,N_19361,N_19147);
and U23195 (N_23195,N_20501,N_19620);
nor U23196 (N_23196,N_21570,N_19360);
and U23197 (N_23197,N_20595,N_20140);
nand U23198 (N_23198,N_20938,N_20469);
nor U23199 (N_23199,N_21161,N_20077);
or U23200 (N_23200,N_19539,N_20735);
nand U23201 (N_23201,N_19741,N_19353);
nand U23202 (N_23202,N_21303,N_20604);
and U23203 (N_23203,N_19486,N_20389);
nand U23204 (N_23204,N_19398,N_19628);
nor U23205 (N_23205,N_19198,N_20270);
and U23206 (N_23206,N_20206,N_20612);
and U23207 (N_23207,N_19968,N_20039);
or U23208 (N_23208,N_20169,N_19245);
nand U23209 (N_23209,N_18976,N_19262);
or U23210 (N_23210,N_20153,N_19425);
nand U23211 (N_23211,N_19005,N_21543);
nand U23212 (N_23212,N_21704,N_20648);
nor U23213 (N_23213,N_20027,N_20021);
or U23214 (N_23214,N_19582,N_18784);
nand U23215 (N_23215,N_21771,N_18821);
and U23216 (N_23216,N_21847,N_21417);
nor U23217 (N_23217,N_20425,N_20953);
and U23218 (N_23218,N_21403,N_19344);
and U23219 (N_23219,N_20723,N_19200);
or U23220 (N_23220,N_20292,N_19026);
or U23221 (N_23221,N_19598,N_19042);
nand U23222 (N_23222,N_21055,N_18839);
nor U23223 (N_23223,N_19031,N_21806);
or U23224 (N_23224,N_19323,N_20491);
or U23225 (N_23225,N_19328,N_21258);
nand U23226 (N_23226,N_21679,N_18837);
or U23227 (N_23227,N_20199,N_19114);
nor U23228 (N_23228,N_21147,N_20774);
nand U23229 (N_23229,N_19267,N_20457);
xor U23230 (N_23230,N_19457,N_19727);
nand U23231 (N_23231,N_19828,N_20402);
nand U23232 (N_23232,N_19916,N_19415);
and U23233 (N_23233,N_19151,N_19223);
and U23234 (N_23234,N_19270,N_20906);
nor U23235 (N_23235,N_21822,N_21524);
nand U23236 (N_23236,N_20690,N_20480);
or U23237 (N_23237,N_19212,N_18955);
nand U23238 (N_23238,N_20344,N_19712);
nand U23239 (N_23239,N_19925,N_21758);
or U23240 (N_23240,N_21368,N_21470);
nor U23241 (N_23241,N_20154,N_20317);
or U23242 (N_23242,N_20673,N_20716);
or U23243 (N_23243,N_20458,N_19498);
nand U23244 (N_23244,N_19889,N_20312);
nor U23245 (N_23245,N_18753,N_21588);
nand U23246 (N_23246,N_20848,N_19139);
or U23247 (N_23247,N_20119,N_21259);
nand U23248 (N_23248,N_19629,N_21045);
nand U23249 (N_23249,N_20400,N_18878);
nor U23250 (N_23250,N_20807,N_19254);
nand U23251 (N_23251,N_20252,N_19152);
xor U23252 (N_23252,N_20638,N_20669);
and U23253 (N_23253,N_18802,N_20666);
nand U23254 (N_23254,N_19320,N_21375);
xnor U23255 (N_23255,N_20968,N_21392);
or U23256 (N_23256,N_20737,N_20145);
or U23257 (N_23257,N_20246,N_21868);
and U23258 (N_23258,N_19218,N_19088);
nor U23259 (N_23259,N_21865,N_20048);
or U23260 (N_23260,N_20290,N_21698);
and U23261 (N_23261,N_21140,N_18907);
or U23262 (N_23262,N_19188,N_20031);
and U23263 (N_23263,N_20238,N_21808);
nand U23264 (N_23264,N_19575,N_19833);
nand U23265 (N_23265,N_21019,N_19167);
and U23266 (N_23266,N_20482,N_18911);
nand U23267 (N_23267,N_18975,N_20367);
and U23268 (N_23268,N_21212,N_19091);
or U23269 (N_23269,N_19545,N_18760);
xor U23270 (N_23270,N_19246,N_20144);
nand U23271 (N_23271,N_20971,N_19971);
nand U23272 (N_23272,N_20987,N_20221);
xnor U23273 (N_23273,N_19070,N_20446);
and U23274 (N_23274,N_20265,N_20511);
nand U23275 (N_23275,N_20350,N_19526);
nand U23276 (N_23276,N_19336,N_21093);
xor U23277 (N_23277,N_19121,N_19662);
xnor U23278 (N_23278,N_20018,N_21369);
nand U23279 (N_23279,N_21421,N_20895);
and U23280 (N_23280,N_20800,N_20853);
xor U23281 (N_23281,N_21468,N_18822);
nand U23282 (N_23282,N_21351,N_21766);
nor U23283 (N_23283,N_21028,N_19041);
and U23284 (N_23284,N_21134,N_21366);
nand U23285 (N_23285,N_20085,N_20362);
nor U23286 (N_23286,N_21779,N_19413);
or U23287 (N_23287,N_18897,N_20525);
nor U23288 (N_23288,N_20672,N_20586);
nor U23289 (N_23289,N_21511,N_21442);
or U23290 (N_23290,N_20984,N_20348);
nor U23291 (N_23291,N_20432,N_19803);
nand U23292 (N_23292,N_18849,N_20616);
or U23293 (N_23293,N_21413,N_20798);
and U23294 (N_23294,N_20101,N_19770);
and U23295 (N_23295,N_18799,N_21307);
nand U23296 (N_23296,N_19711,N_21089);
and U23297 (N_23297,N_20123,N_18758);
nand U23298 (N_23298,N_21592,N_19065);
nor U23299 (N_23299,N_21209,N_21539);
or U23300 (N_23300,N_19043,N_21274);
and U23301 (N_23301,N_19169,N_18974);
nor U23302 (N_23302,N_19129,N_21214);
or U23303 (N_23303,N_20621,N_19036);
and U23304 (N_23304,N_21606,N_19607);
nor U23305 (N_23305,N_19118,N_19938);
nor U23306 (N_23306,N_20499,N_20569);
or U23307 (N_23307,N_21754,N_20516);
or U23308 (N_23308,N_21436,N_20898);
xor U23309 (N_23309,N_21467,N_21659);
nor U23310 (N_23310,N_19119,N_20165);
nand U23311 (N_23311,N_21457,N_19866);
nand U23312 (N_23312,N_18998,N_21475);
and U23313 (N_23313,N_20708,N_21342);
or U23314 (N_23314,N_20646,N_19614);
or U23315 (N_23315,N_19611,N_20860);
and U23316 (N_23316,N_19446,N_19051);
and U23317 (N_23317,N_19796,N_20267);
nand U23318 (N_23318,N_21217,N_21717);
or U23319 (N_23319,N_20053,N_18888);
or U23320 (N_23320,N_19800,N_20890);
nor U23321 (N_23321,N_19690,N_21782);
and U23322 (N_23322,N_21042,N_20136);
nor U23323 (N_23323,N_19453,N_19815);
or U23324 (N_23324,N_20345,N_21763);
and U23325 (N_23325,N_21666,N_21122);
and U23326 (N_23326,N_19584,N_21223);
or U23327 (N_23327,N_20956,N_19217);
nand U23328 (N_23328,N_21780,N_19830);
nand U23329 (N_23329,N_19615,N_20057);
or U23330 (N_23330,N_19877,N_20812);
and U23331 (N_23331,N_19623,N_18759);
xnor U23332 (N_23332,N_18922,N_21681);
and U23333 (N_23333,N_19753,N_21558);
or U23334 (N_23334,N_20816,N_21557);
or U23335 (N_23335,N_20617,N_19512);
nand U23336 (N_23336,N_19396,N_20655);
xor U23337 (N_23337,N_21078,N_20375);
or U23338 (N_23338,N_19982,N_21097);
nand U23339 (N_23339,N_19953,N_20978);
and U23340 (N_23340,N_21244,N_20016);
nor U23341 (N_23341,N_20006,N_19688);
nor U23342 (N_23342,N_21213,N_20834);
or U23343 (N_23343,N_21542,N_21157);
or U23344 (N_23344,N_21493,N_20573);
or U23345 (N_23345,N_21287,N_21488);
or U23346 (N_23346,N_19973,N_20900);
or U23347 (N_23347,N_21345,N_21474);
and U23348 (N_23348,N_21427,N_19946);
and U23349 (N_23349,N_20235,N_20214);
nor U23350 (N_23350,N_21802,N_20819);
nand U23351 (N_23351,N_20255,N_20106);
nor U23352 (N_23352,N_19646,N_21272);
and U23353 (N_23353,N_19747,N_20464);
or U23354 (N_23354,N_21336,N_19855);
or U23355 (N_23355,N_19141,N_19847);
nor U23356 (N_23356,N_21114,N_18883);
nor U23357 (N_23357,N_20380,N_20750);
and U23358 (N_23358,N_20986,N_21329);
and U23359 (N_23359,N_20541,N_19924);
nand U23360 (N_23360,N_19251,N_19392);
and U23361 (N_23361,N_21636,N_21197);
nand U23362 (N_23362,N_21273,N_19892);
and U23363 (N_23363,N_19239,N_19421);
nand U23364 (N_23364,N_20651,N_20319);
and U23365 (N_23365,N_21729,N_20688);
nand U23366 (N_23366,N_19350,N_19179);
or U23367 (N_23367,N_21680,N_20131);
nand U23368 (N_23368,N_19670,N_20261);
nor U23369 (N_23369,N_20231,N_20660);
or U23370 (N_23370,N_21586,N_18813);
nor U23371 (N_23371,N_19592,N_21378);
nand U23372 (N_23372,N_19487,N_19326);
and U23373 (N_23373,N_19235,N_21804);
nand U23374 (N_23374,N_20395,N_20128);
xor U23375 (N_23375,N_21513,N_21784);
nand U23376 (N_23376,N_18902,N_20082);
or U23377 (N_23377,N_20381,N_20619);
or U23378 (N_23378,N_21485,N_21790);
or U23379 (N_23379,N_20872,N_21756);
nand U23380 (N_23380,N_20023,N_20466);
and U23381 (N_23381,N_19612,N_20440);
or U23382 (N_23382,N_19661,N_21657);
nand U23383 (N_23383,N_19931,N_21647);
nor U23384 (N_23384,N_20649,N_18871);
and U23385 (N_23385,N_19561,N_20296);
and U23386 (N_23386,N_21869,N_19325);
nor U23387 (N_23387,N_19986,N_19466);
nor U23388 (N_23388,N_19864,N_21858);
nor U23389 (N_23389,N_21481,N_19528);
or U23390 (N_23390,N_20203,N_20488);
or U23391 (N_23391,N_20405,N_20143);
and U23392 (N_23392,N_21172,N_19055);
nand U23393 (N_23393,N_21820,N_18894);
nor U23394 (N_23394,N_21241,N_21800);
nor U23395 (N_23395,N_21705,N_20217);
nand U23396 (N_23396,N_18884,N_18851);
nand U23397 (N_23397,N_20327,N_20838);
or U23398 (N_23398,N_21030,N_20545);
and U23399 (N_23399,N_19911,N_19414);
nand U23400 (N_23400,N_21424,N_20744);
nand U23401 (N_23401,N_20008,N_21116);
or U23402 (N_23402,N_20124,N_20034);
and U23403 (N_23403,N_21297,N_21405);
or U23404 (N_23404,N_20518,N_19012);
nor U23405 (N_23405,N_21634,N_20794);
and U23406 (N_23406,N_19168,N_21388);
and U23407 (N_23407,N_20228,N_20302);
or U23408 (N_23408,N_20961,N_20593);
nor U23409 (N_23409,N_19205,N_21084);
nor U23410 (N_23410,N_19472,N_19774);
nand U23411 (N_23411,N_20592,N_20854);
or U23412 (N_23412,N_20704,N_21108);
or U23413 (N_23413,N_21162,N_21833);
or U23414 (N_23414,N_18869,N_21811);
and U23415 (N_23415,N_19503,N_20766);
or U23416 (N_23416,N_19399,N_19814);
nand U23417 (N_23417,N_19948,N_20929);
nor U23418 (N_23418,N_18913,N_19873);
and U23419 (N_23419,N_20923,N_19146);
nor U23420 (N_23420,N_19290,N_19927);
or U23421 (N_23421,N_19298,N_21358);
nor U23422 (N_23422,N_21070,N_20033);
and U23423 (N_23423,N_21460,N_19476);
nand U23424 (N_23424,N_19706,N_20554);
nor U23425 (N_23425,N_20839,N_21350);
and U23426 (N_23426,N_19640,N_20835);
and U23427 (N_23427,N_21037,N_19310);
or U23428 (N_23428,N_21109,N_19439);
nand U23429 (N_23429,N_19783,N_18859);
xor U23430 (N_23430,N_19166,N_19874);
or U23431 (N_23431,N_20931,N_18893);
or U23432 (N_23432,N_21177,N_21701);
xor U23433 (N_23433,N_18755,N_19079);
nor U23434 (N_23434,N_19366,N_19524);
nand U23435 (N_23435,N_21407,N_20989);
nor U23436 (N_23436,N_19742,N_21658);
nor U23437 (N_23437,N_19577,N_20900);
or U23438 (N_23438,N_21446,N_19984);
nor U23439 (N_23439,N_19892,N_19557);
nand U23440 (N_23440,N_21051,N_20951);
xor U23441 (N_23441,N_19000,N_19064);
nand U23442 (N_23442,N_19403,N_19635);
xnor U23443 (N_23443,N_19771,N_20602);
xnor U23444 (N_23444,N_20651,N_20836);
and U23445 (N_23445,N_20182,N_20073);
or U23446 (N_23446,N_19432,N_20871);
or U23447 (N_23447,N_20076,N_21654);
nand U23448 (N_23448,N_19660,N_20244);
or U23449 (N_23449,N_20912,N_21447);
nand U23450 (N_23450,N_21432,N_20579);
nor U23451 (N_23451,N_21646,N_20169);
nor U23452 (N_23452,N_18945,N_21705);
and U23453 (N_23453,N_21185,N_20128);
xor U23454 (N_23454,N_20328,N_21038);
or U23455 (N_23455,N_21078,N_20534);
nor U23456 (N_23456,N_21847,N_21619);
or U23457 (N_23457,N_21058,N_20290);
nand U23458 (N_23458,N_21147,N_19815);
or U23459 (N_23459,N_19762,N_19899);
nor U23460 (N_23460,N_21147,N_20807);
xor U23461 (N_23461,N_20523,N_21845);
nand U23462 (N_23462,N_20775,N_19144);
nor U23463 (N_23463,N_19152,N_21669);
nor U23464 (N_23464,N_20064,N_20903);
and U23465 (N_23465,N_18870,N_20797);
nor U23466 (N_23466,N_21629,N_19050);
or U23467 (N_23467,N_21045,N_20813);
nor U23468 (N_23468,N_20595,N_20670);
nor U23469 (N_23469,N_21067,N_20240);
and U23470 (N_23470,N_21342,N_21710);
and U23471 (N_23471,N_19845,N_19658);
or U23472 (N_23472,N_20660,N_20668);
nor U23473 (N_23473,N_19992,N_19090);
nand U23474 (N_23474,N_20965,N_21584);
nand U23475 (N_23475,N_18774,N_21348);
and U23476 (N_23476,N_20323,N_20745);
nand U23477 (N_23477,N_20103,N_19550);
and U23478 (N_23478,N_21819,N_19372);
nand U23479 (N_23479,N_20541,N_19219);
or U23480 (N_23480,N_20933,N_18848);
nor U23481 (N_23481,N_21833,N_21778);
or U23482 (N_23482,N_21838,N_20629);
nand U23483 (N_23483,N_20744,N_20602);
nor U23484 (N_23484,N_18941,N_19833);
or U23485 (N_23485,N_20047,N_20672);
or U23486 (N_23486,N_20051,N_19165);
nor U23487 (N_23487,N_20717,N_21161);
xnor U23488 (N_23488,N_19241,N_19520);
and U23489 (N_23489,N_19321,N_21186);
xor U23490 (N_23490,N_18777,N_19820);
and U23491 (N_23491,N_21052,N_19476);
nor U23492 (N_23492,N_21733,N_21020);
nand U23493 (N_23493,N_21244,N_19394);
nor U23494 (N_23494,N_20966,N_20822);
nor U23495 (N_23495,N_21421,N_21058);
or U23496 (N_23496,N_20930,N_19298);
xor U23497 (N_23497,N_19745,N_19349);
and U23498 (N_23498,N_19767,N_21130);
nand U23499 (N_23499,N_18988,N_20092);
or U23500 (N_23500,N_19901,N_20047);
nor U23501 (N_23501,N_19607,N_20631);
nand U23502 (N_23502,N_21353,N_21246);
xnor U23503 (N_23503,N_21170,N_19003);
and U23504 (N_23504,N_21723,N_20300);
or U23505 (N_23505,N_20785,N_20730);
or U23506 (N_23506,N_21263,N_20472);
and U23507 (N_23507,N_21310,N_19712);
nor U23508 (N_23508,N_21734,N_20938);
or U23509 (N_23509,N_21010,N_21140);
and U23510 (N_23510,N_19934,N_21759);
nand U23511 (N_23511,N_21758,N_20799);
nand U23512 (N_23512,N_19229,N_21076);
and U23513 (N_23513,N_20374,N_19007);
and U23514 (N_23514,N_19150,N_18947);
nor U23515 (N_23515,N_19632,N_21536);
nand U23516 (N_23516,N_21384,N_19845);
or U23517 (N_23517,N_20875,N_21697);
nand U23518 (N_23518,N_19909,N_20726);
and U23519 (N_23519,N_19514,N_19533);
xnor U23520 (N_23520,N_20061,N_19758);
and U23521 (N_23521,N_20793,N_19442);
and U23522 (N_23522,N_20962,N_20170);
nor U23523 (N_23523,N_18991,N_18920);
or U23524 (N_23524,N_20099,N_19527);
and U23525 (N_23525,N_19835,N_20224);
or U23526 (N_23526,N_21312,N_20440);
and U23527 (N_23527,N_19335,N_20823);
nand U23528 (N_23528,N_21506,N_19694);
xor U23529 (N_23529,N_21271,N_20071);
and U23530 (N_23530,N_19680,N_21651);
and U23531 (N_23531,N_21289,N_19055);
nand U23532 (N_23532,N_21239,N_18775);
or U23533 (N_23533,N_21285,N_19066);
nand U23534 (N_23534,N_21569,N_20507);
or U23535 (N_23535,N_19278,N_18966);
or U23536 (N_23536,N_18900,N_19155);
or U23537 (N_23537,N_19169,N_20630);
nor U23538 (N_23538,N_20053,N_21101);
nor U23539 (N_23539,N_21012,N_21511);
nor U23540 (N_23540,N_19849,N_19210);
or U23541 (N_23541,N_20508,N_20744);
or U23542 (N_23542,N_21547,N_19047);
nor U23543 (N_23543,N_20799,N_21620);
nand U23544 (N_23544,N_21644,N_21277);
xnor U23545 (N_23545,N_20036,N_20211);
xor U23546 (N_23546,N_21442,N_19944);
nand U23547 (N_23547,N_19543,N_19271);
or U23548 (N_23548,N_20974,N_21125);
and U23549 (N_23549,N_19943,N_20521);
nor U23550 (N_23550,N_20562,N_19413);
or U23551 (N_23551,N_19806,N_19830);
or U23552 (N_23552,N_20446,N_21668);
nor U23553 (N_23553,N_20855,N_20185);
xor U23554 (N_23554,N_19029,N_18927);
and U23555 (N_23555,N_20731,N_20911);
nor U23556 (N_23556,N_20398,N_21720);
nor U23557 (N_23557,N_21404,N_19507);
and U23558 (N_23558,N_20762,N_20688);
nand U23559 (N_23559,N_19754,N_19371);
nand U23560 (N_23560,N_20013,N_18834);
or U23561 (N_23561,N_19289,N_21516);
nand U23562 (N_23562,N_21541,N_21537);
or U23563 (N_23563,N_18839,N_21679);
and U23564 (N_23564,N_21386,N_19977);
nand U23565 (N_23565,N_21194,N_21298);
and U23566 (N_23566,N_21234,N_20365);
and U23567 (N_23567,N_20663,N_20367);
or U23568 (N_23568,N_21840,N_19833);
xor U23569 (N_23569,N_19526,N_20882);
xor U23570 (N_23570,N_19332,N_21611);
xnor U23571 (N_23571,N_20179,N_18984);
or U23572 (N_23572,N_20617,N_20965);
or U23573 (N_23573,N_21599,N_19904);
nor U23574 (N_23574,N_19709,N_21607);
or U23575 (N_23575,N_19385,N_20129);
and U23576 (N_23576,N_21804,N_19953);
or U23577 (N_23577,N_19405,N_19584);
nor U23578 (N_23578,N_20458,N_21243);
or U23579 (N_23579,N_20179,N_20227);
and U23580 (N_23580,N_19208,N_18816);
nand U23581 (N_23581,N_19505,N_19815);
nand U23582 (N_23582,N_19055,N_21525);
nor U23583 (N_23583,N_21346,N_19239);
and U23584 (N_23584,N_21482,N_19629);
and U23585 (N_23585,N_19404,N_20339);
nand U23586 (N_23586,N_20356,N_21113);
and U23587 (N_23587,N_19107,N_19986);
or U23588 (N_23588,N_18971,N_19700);
or U23589 (N_23589,N_19797,N_21673);
xnor U23590 (N_23590,N_21178,N_20240);
nor U23591 (N_23591,N_20401,N_21126);
xor U23592 (N_23592,N_20982,N_20823);
nor U23593 (N_23593,N_18940,N_21777);
and U23594 (N_23594,N_20838,N_18899);
and U23595 (N_23595,N_19047,N_19989);
nor U23596 (N_23596,N_19078,N_19732);
nand U23597 (N_23597,N_18833,N_21122);
or U23598 (N_23598,N_19507,N_20969);
nand U23599 (N_23599,N_19557,N_19440);
xor U23600 (N_23600,N_20459,N_18755);
nor U23601 (N_23601,N_18759,N_19555);
or U23602 (N_23602,N_21578,N_20529);
or U23603 (N_23603,N_20788,N_20168);
nor U23604 (N_23604,N_21656,N_21742);
nand U23605 (N_23605,N_21813,N_19181);
or U23606 (N_23606,N_19083,N_20349);
or U23607 (N_23607,N_21766,N_20102);
nor U23608 (N_23608,N_18790,N_19350);
xor U23609 (N_23609,N_20152,N_20840);
and U23610 (N_23610,N_21006,N_19738);
nand U23611 (N_23611,N_20718,N_21685);
nand U23612 (N_23612,N_19286,N_21392);
nor U23613 (N_23613,N_19592,N_20696);
nor U23614 (N_23614,N_20959,N_20834);
nor U23615 (N_23615,N_21357,N_21507);
and U23616 (N_23616,N_21418,N_21689);
nand U23617 (N_23617,N_19500,N_18984);
and U23618 (N_23618,N_19236,N_19991);
nor U23619 (N_23619,N_21238,N_19986);
or U23620 (N_23620,N_20002,N_21275);
and U23621 (N_23621,N_20636,N_19271);
and U23622 (N_23622,N_19251,N_21664);
nor U23623 (N_23623,N_20433,N_19416);
and U23624 (N_23624,N_19445,N_19461);
xnor U23625 (N_23625,N_19126,N_20994);
or U23626 (N_23626,N_19036,N_21710);
nor U23627 (N_23627,N_19066,N_20347);
or U23628 (N_23628,N_21801,N_19185);
or U23629 (N_23629,N_20871,N_19180);
nand U23630 (N_23630,N_19497,N_19449);
nor U23631 (N_23631,N_21783,N_20680);
nor U23632 (N_23632,N_20709,N_21471);
or U23633 (N_23633,N_19784,N_19159);
nor U23634 (N_23634,N_20567,N_21293);
nand U23635 (N_23635,N_21201,N_19757);
nand U23636 (N_23636,N_20228,N_21757);
xor U23637 (N_23637,N_19506,N_20510);
nor U23638 (N_23638,N_21787,N_21468);
or U23639 (N_23639,N_21592,N_20295);
and U23640 (N_23640,N_20940,N_21697);
and U23641 (N_23641,N_18985,N_21167);
nand U23642 (N_23642,N_20115,N_20743);
nor U23643 (N_23643,N_21754,N_19314);
or U23644 (N_23644,N_21696,N_20498);
and U23645 (N_23645,N_20266,N_18820);
nor U23646 (N_23646,N_21718,N_21776);
nand U23647 (N_23647,N_19671,N_19048);
or U23648 (N_23648,N_20243,N_20402);
xnor U23649 (N_23649,N_20805,N_21488);
xnor U23650 (N_23650,N_20274,N_20079);
and U23651 (N_23651,N_19020,N_21023);
or U23652 (N_23652,N_21345,N_20942);
and U23653 (N_23653,N_21738,N_18992);
nand U23654 (N_23654,N_20409,N_19019);
nor U23655 (N_23655,N_21731,N_20087);
xor U23656 (N_23656,N_20107,N_20565);
and U23657 (N_23657,N_21126,N_21818);
or U23658 (N_23658,N_20538,N_21652);
nand U23659 (N_23659,N_20629,N_21594);
and U23660 (N_23660,N_19416,N_20778);
and U23661 (N_23661,N_21692,N_21170);
nand U23662 (N_23662,N_21392,N_20412);
nand U23663 (N_23663,N_19556,N_20158);
nor U23664 (N_23664,N_21122,N_19683);
xor U23665 (N_23665,N_18842,N_20340);
nor U23666 (N_23666,N_21538,N_21305);
nand U23667 (N_23667,N_19363,N_19046);
xor U23668 (N_23668,N_21322,N_19727);
xnor U23669 (N_23669,N_21456,N_19518);
or U23670 (N_23670,N_20265,N_19144);
nor U23671 (N_23671,N_18871,N_19418);
nand U23672 (N_23672,N_19865,N_19487);
nor U23673 (N_23673,N_19258,N_19190);
or U23674 (N_23674,N_21696,N_21583);
nand U23675 (N_23675,N_19927,N_20004);
or U23676 (N_23676,N_18978,N_19051);
or U23677 (N_23677,N_18964,N_20795);
nand U23678 (N_23678,N_20688,N_20805);
or U23679 (N_23679,N_20026,N_19423);
nor U23680 (N_23680,N_20482,N_21740);
xnor U23681 (N_23681,N_18963,N_19227);
and U23682 (N_23682,N_21585,N_20907);
and U23683 (N_23683,N_20419,N_19731);
nand U23684 (N_23684,N_20306,N_21036);
nor U23685 (N_23685,N_20896,N_21140);
nor U23686 (N_23686,N_20536,N_21620);
nand U23687 (N_23687,N_21831,N_21307);
nor U23688 (N_23688,N_21252,N_21408);
xor U23689 (N_23689,N_21172,N_19333);
nor U23690 (N_23690,N_20987,N_18887);
and U23691 (N_23691,N_19348,N_19263);
xnor U23692 (N_23692,N_21369,N_21723);
xnor U23693 (N_23693,N_19885,N_20864);
nand U23694 (N_23694,N_21324,N_20807);
xnor U23695 (N_23695,N_20982,N_18945);
xor U23696 (N_23696,N_21218,N_20137);
or U23697 (N_23697,N_19068,N_19937);
nand U23698 (N_23698,N_19823,N_20950);
nor U23699 (N_23699,N_19901,N_19870);
nor U23700 (N_23700,N_21756,N_20798);
and U23701 (N_23701,N_19906,N_20700);
nand U23702 (N_23702,N_20525,N_20676);
nor U23703 (N_23703,N_21491,N_20099);
nand U23704 (N_23704,N_19285,N_19672);
and U23705 (N_23705,N_18830,N_20032);
and U23706 (N_23706,N_19748,N_21258);
nand U23707 (N_23707,N_21165,N_21728);
nor U23708 (N_23708,N_21145,N_21051);
and U23709 (N_23709,N_21352,N_19565);
and U23710 (N_23710,N_20142,N_19712);
nand U23711 (N_23711,N_19971,N_21378);
nand U23712 (N_23712,N_19673,N_19154);
and U23713 (N_23713,N_21160,N_20004);
nor U23714 (N_23714,N_20986,N_20152);
or U23715 (N_23715,N_20938,N_19138);
and U23716 (N_23716,N_20196,N_20775);
or U23717 (N_23717,N_18811,N_18840);
nor U23718 (N_23718,N_20484,N_21631);
and U23719 (N_23719,N_19021,N_20740);
and U23720 (N_23720,N_20832,N_20122);
and U23721 (N_23721,N_18897,N_21198);
nor U23722 (N_23722,N_20545,N_20458);
and U23723 (N_23723,N_20252,N_21234);
or U23724 (N_23724,N_21320,N_19371);
or U23725 (N_23725,N_21375,N_21658);
or U23726 (N_23726,N_18882,N_19981);
and U23727 (N_23727,N_20363,N_19222);
xor U23728 (N_23728,N_19775,N_19634);
and U23729 (N_23729,N_19679,N_18833);
or U23730 (N_23730,N_21648,N_19120);
or U23731 (N_23731,N_20686,N_20803);
and U23732 (N_23732,N_20135,N_19459);
or U23733 (N_23733,N_18961,N_20045);
nand U23734 (N_23734,N_20897,N_20977);
nor U23735 (N_23735,N_21578,N_19150);
or U23736 (N_23736,N_20964,N_20442);
nor U23737 (N_23737,N_19176,N_18988);
or U23738 (N_23738,N_20723,N_20390);
nor U23739 (N_23739,N_19604,N_21318);
and U23740 (N_23740,N_19245,N_21484);
or U23741 (N_23741,N_19100,N_21343);
and U23742 (N_23742,N_21493,N_20424);
nand U23743 (N_23743,N_21202,N_19946);
nor U23744 (N_23744,N_21035,N_18978);
or U23745 (N_23745,N_19725,N_21296);
or U23746 (N_23746,N_18829,N_19585);
or U23747 (N_23747,N_19109,N_19993);
and U23748 (N_23748,N_19679,N_19213);
and U23749 (N_23749,N_20949,N_18800);
nand U23750 (N_23750,N_19043,N_21487);
and U23751 (N_23751,N_20541,N_20109);
nor U23752 (N_23752,N_20479,N_19275);
xor U23753 (N_23753,N_21339,N_21790);
or U23754 (N_23754,N_21409,N_20585);
or U23755 (N_23755,N_20126,N_21393);
xnor U23756 (N_23756,N_20271,N_21825);
nor U23757 (N_23757,N_19338,N_21188);
xnor U23758 (N_23758,N_19885,N_20648);
or U23759 (N_23759,N_20514,N_19535);
xnor U23760 (N_23760,N_18917,N_20888);
nor U23761 (N_23761,N_20080,N_20690);
nor U23762 (N_23762,N_21553,N_20257);
nor U23763 (N_23763,N_19502,N_18825);
or U23764 (N_23764,N_20530,N_19039);
and U23765 (N_23765,N_18923,N_20047);
xnor U23766 (N_23766,N_19484,N_19714);
nor U23767 (N_23767,N_19616,N_19518);
nor U23768 (N_23768,N_21362,N_20894);
and U23769 (N_23769,N_21749,N_20970);
nand U23770 (N_23770,N_21864,N_20259);
nor U23771 (N_23771,N_21657,N_19698);
nor U23772 (N_23772,N_19536,N_19478);
and U23773 (N_23773,N_19767,N_21067);
nand U23774 (N_23774,N_18915,N_20979);
nor U23775 (N_23775,N_19291,N_21637);
and U23776 (N_23776,N_19671,N_19835);
nor U23777 (N_23777,N_20893,N_20853);
nand U23778 (N_23778,N_18845,N_21004);
nand U23779 (N_23779,N_20785,N_19745);
or U23780 (N_23780,N_20541,N_19406);
nor U23781 (N_23781,N_20743,N_20850);
or U23782 (N_23782,N_21109,N_21310);
nand U23783 (N_23783,N_19391,N_20332);
nor U23784 (N_23784,N_21614,N_21175);
or U23785 (N_23785,N_19314,N_21116);
and U23786 (N_23786,N_21432,N_19228);
nand U23787 (N_23787,N_19315,N_19518);
or U23788 (N_23788,N_19264,N_21422);
or U23789 (N_23789,N_18905,N_21062);
or U23790 (N_23790,N_19784,N_19788);
nand U23791 (N_23791,N_21357,N_20982);
or U23792 (N_23792,N_21667,N_21396);
nor U23793 (N_23793,N_19007,N_20375);
xnor U23794 (N_23794,N_19012,N_19168);
nor U23795 (N_23795,N_20385,N_19036);
xnor U23796 (N_23796,N_19263,N_21787);
nand U23797 (N_23797,N_19989,N_19720);
and U23798 (N_23798,N_20372,N_21058);
nand U23799 (N_23799,N_21142,N_20578);
or U23800 (N_23800,N_20839,N_19434);
nand U23801 (N_23801,N_19612,N_20355);
nand U23802 (N_23802,N_19827,N_19267);
nand U23803 (N_23803,N_19235,N_20383);
and U23804 (N_23804,N_19190,N_20267);
or U23805 (N_23805,N_20686,N_18754);
or U23806 (N_23806,N_18993,N_19629);
nand U23807 (N_23807,N_18848,N_19877);
and U23808 (N_23808,N_21777,N_21837);
or U23809 (N_23809,N_19718,N_20401);
and U23810 (N_23810,N_21158,N_19106);
and U23811 (N_23811,N_19903,N_19011);
xnor U23812 (N_23812,N_20400,N_20801);
nor U23813 (N_23813,N_21431,N_20662);
nor U23814 (N_23814,N_19867,N_21567);
nand U23815 (N_23815,N_21631,N_21500);
nor U23816 (N_23816,N_19087,N_21620);
nor U23817 (N_23817,N_21691,N_21344);
or U23818 (N_23818,N_19501,N_19645);
and U23819 (N_23819,N_20527,N_20034);
nor U23820 (N_23820,N_20686,N_19360);
nand U23821 (N_23821,N_20305,N_19408);
nand U23822 (N_23822,N_19895,N_18780);
and U23823 (N_23823,N_21870,N_21440);
or U23824 (N_23824,N_19381,N_21138);
nor U23825 (N_23825,N_18778,N_21855);
nor U23826 (N_23826,N_20386,N_19033);
and U23827 (N_23827,N_20308,N_21208);
and U23828 (N_23828,N_21833,N_21128);
nor U23829 (N_23829,N_21153,N_21084);
nand U23830 (N_23830,N_21125,N_19559);
and U23831 (N_23831,N_21143,N_21004);
and U23832 (N_23832,N_19920,N_20667);
or U23833 (N_23833,N_19480,N_19049);
nor U23834 (N_23834,N_20856,N_21219);
xnor U23835 (N_23835,N_21830,N_19319);
or U23836 (N_23836,N_21167,N_18792);
and U23837 (N_23837,N_19780,N_21642);
and U23838 (N_23838,N_20315,N_19720);
nand U23839 (N_23839,N_21128,N_20463);
or U23840 (N_23840,N_21261,N_21710);
or U23841 (N_23841,N_20827,N_21518);
nand U23842 (N_23842,N_20699,N_19521);
nand U23843 (N_23843,N_20165,N_19281);
or U23844 (N_23844,N_21739,N_19052);
and U23845 (N_23845,N_19722,N_20587);
xor U23846 (N_23846,N_19855,N_20441);
or U23847 (N_23847,N_20625,N_18909);
nand U23848 (N_23848,N_21489,N_19678);
or U23849 (N_23849,N_20004,N_21795);
xnor U23850 (N_23850,N_21125,N_21593);
xnor U23851 (N_23851,N_20928,N_21109);
nand U23852 (N_23852,N_19075,N_20900);
and U23853 (N_23853,N_21442,N_19662);
nand U23854 (N_23854,N_20551,N_21297);
and U23855 (N_23855,N_20653,N_20736);
and U23856 (N_23856,N_21313,N_20061);
nand U23857 (N_23857,N_19701,N_21047);
and U23858 (N_23858,N_21724,N_18891);
nand U23859 (N_23859,N_19115,N_21111);
and U23860 (N_23860,N_19146,N_20877);
xnor U23861 (N_23861,N_20254,N_19685);
or U23862 (N_23862,N_19096,N_19963);
and U23863 (N_23863,N_19943,N_19088);
and U23864 (N_23864,N_21565,N_21628);
or U23865 (N_23865,N_18916,N_18915);
and U23866 (N_23866,N_19007,N_21260);
nand U23867 (N_23867,N_20598,N_19286);
or U23868 (N_23868,N_19068,N_20753);
and U23869 (N_23869,N_20037,N_20528);
and U23870 (N_23870,N_19516,N_21823);
nand U23871 (N_23871,N_20781,N_19883);
nor U23872 (N_23872,N_21869,N_20267);
or U23873 (N_23873,N_19109,N_21092);
nand U23874 (N_23874,N_20629,N_19231);
nor U23875 (N_23875,N_19620,N_19330);
and U23876 (N_23876,N_19627,N_19596);
or U23877 (N_23877,N_21603,N_19942);
nor U23878 (N_23878,N_21256,N_18759);
or U23879 (N_23879,N_21292,N_21474);
or U23880 (N_23880,N_18992,N_20042);
nor U23881 (N_23881,N_21529,N_20474);
and U23882 (N_23882,N_18902,N_20462);
and U23883 (N_23883,N_21798,N_19155);
and U23884 (N_23884,N_21802,N_21055);
nor U23885 (N_23885,N_21056,N_20860);
nand U23886 (N_23886,N_20346,N_19633);
nor U23887 (N_23887,N_19096,N_21572);
and U23888 (N_23888,N_21068,N_20510);
and U23889 (N_23889,N_20668,N_21118);
nor U23890 (N_23890,N_21420,N_20825);
nor U23891 (N_23891,N_19287,N_21821);
nand U23892 (N_23892,N_19021,N_19307);
nand U23893 (N_23893,N_21742,N_21747);
nor U23894 (N_23894,N_19869,N_21536);
nor U23895 (N_23895,N_20831,N_19399);
nor U23896 (N_23896,N_20585,N_19684);
nor U23897 (N_23897,N_19445,N_19840);
and U23898 (N_23898,N_20963,N_19293);
nor U23899 (N_23899,N_21842,N_21678);
nor U23900 (N_23900,N_19856,N_21346);
or U23901 (N_23901,N_21575,N_20766);
nor U23902 (N_23902,N_21488,N_20743);
nand U23903 (N_23903,N_19570,N_20101);
nor U23904 (N_23904,N_20556,N_19742);
and U23905 (N_23905,N_21238,N_20343);
or U23906 (N_23906,N_20077,N_20045);
nor U23907 (N_23907,N_19712,N_19440);
nor U23908 (N_23908,N_21008,N_20708);
or U23909 (N_23909,N_20704,N_19637);
nor U23910 (N_23910,N_20227,N_19750);
xnor U23911 (N_23911,N_18843,N_21492);
nor U23912 (N_23912,N_21258,N_18781);
and U23913 (N_23913,N_19445,N_19320);
and U23914 (N_23914,N_20100,N_19407);
nand U23915 (N_23915,N_20794,N_20677);
nor U23916 (N_23916,N_19510,N_21700);
nand U23917 (N_23917,N_21143,N_20545);
nor U23918 (N_23918,N_21754,N_20953);
nand U23919 (N_23919,N_20412,N_19128);
or U23920 (N_23920,N_19810,N_21002);
nand U23921 (N_23921,N_21781,N_19842);
and U23922 (N_23922,N_21358,N_20010);
nand U23923 (N_23923,N_20597,N_19221);
nor U23924 (N_23924,N_20001,N_21790);
nor U23925 (N_23925,N_21313,N_21124);
or U23926 (N_23926,N_19454,N_19463);
and U23927 (N_23927,N_21299,N_21056);
xor U23928 (N_23928,N_21814,N_19579);
and U23929 (N_23929,N_19291,N_20673);
or U23930 (N_23930,N_20687,N_19463);
nand U23931 (N_23931,N_21507,N_19063);
nor U23932 (N_23932,N_20596,N_21002);
nor U23933 (N_23933,N_19069,N_21534);
nor U23934 (N_23934,N_19549,N_21792);
nand U23935 (N_23935,N_20446,N_19781);
or U23936 (N_23936,N_20322,N_20220);
nand U23937 (N_23937,N_20458,N_18778);
and U23938 (N_23938,N_20283,N_18939);
nor U23939 (N_23939,N_21749,N_20947);
or U23940 (N_23940,N_21828,N_21762);
nor U23941 (N_23941,N_20936,N_19604);
nor U23942 (N_23942,N_21342,N_21304);
xor U23943 (N_23943,N_18816,N_19123);
or U23944 (N_23944,N_19661,N_20046);
nand U23945 (N_23945,N_19723,N_21387);
and U23946 (N_23946,N_21671,N_19048);
or U23947 (N_23947,N_19903,N_21621);
or U23948 (N_23948,N_21655,N_19213);
nand U23949 (N_23949,N_20505,N_19110);
nor U23950 (N_23950,N_19416,N_20891);
or U23951 (N_23951,N_19703,N_20024);
nor U23952 (N_23952,N_21279,N_21183);
and U23953 (N_23953,N_20123,N_20461);
and U23954 (N_23954,N_21186,N_18782);
or U23955 (N_23955,N_21134,N_18983);
and U23956 (N_23956,N_19121,N_21468);
nor U23957 (N_23957,N_18981,N_21329);
or U23958 (N_23958,N_20560,N_20886);
nand U23959 (N_23959,N_20490,N_19482);
and U23960 (N_23960,N_20198,N_18954);
xor U23961 (N_23961,N_21029,N_19267);
xnor U23962 (N_23962,N_18840,N_21738);
and U23963 (N_23963,N_20284,N_20165);
nor U23964 (N_23964,N_19725,N_21048);
and U23965 (N_23965,N_19182,N_19290);
nand U23966 (N_23966,N_19364,N_18942);
nor U23967 (N_23967,N_20635,N_20537);
and U23968 (N_23968,N_20614,N_20727);
nor U23969 (N_23969,N_21201,N_19134);
nor U23970 (N_23970,N_21121,N_18828);
and U23971 (N_23971,N_20262,N_21663);
xor U23972 (N_23972,N_19800,N_19041);
or U23973 (N_23973,N_20083,N_20677);
and U23974 (N_23974,N_20248,N_19761);
and U23975 (N_23975,N_20952,N_19120);
xnor U23976 (N_23976,N_21318,N_20961);
nor U23977 (N_23977,N_20285,N_21125);
or U23978 (N_23978,N_19734,N_20091);
or U23979 (N_23979,N_20176,N_21555);
nor U23980 (N_23980,N_19037,N_20379);
nand U23981 (N_23981,N_21490,N_19199);
nand U23982 (N_23982,N_20088,N_21046);
and U23983 (N_23983,N_21351,N_19819);
or U23984 (N_23984,N_19480,N_19089);
or U23985 (N_23985,N_20208,N_21273);
nor U23986 (N_23986,N_19247,N_20415);
xor U23987 (N_23987,N_19424,N_21425);
or U23988 (N_23988,N_21061,N_20711);
and U23989 (N_23989,N_20449,N_20873);
nand U23990 (N_23990,N_20289,N_19468);
nor U23991 (N_23991,N_21610,N_21792);
nand U23992 (N_23992,N_21421,N_21413);
and U23993 (N_23993,N_19043,N_21587);
and U23994 (N_23994,N_19651,N_20238);
or U23995 (N_23995,N_21711,N_20116);
nand U23996 (N_23996,N_19577,N_19899);
or U23997 (N_23997,N_21826,N_21779);
and U23998 (N_23998,N_18867,N_21243);
and U23999 (N_23999,N_18919,N_19999);
and U24000 (N_24000,N_19154,N_21609);
nand U24001 (N_24001,N_18852,N_20774);
nor U24002 (N_24002,N_21337,N_19526);
nor U24003 (N_24003,N_19514,N_21136);
nor U24004 (N_24004,N_20945,N_19699);
nor U24005 (N_24005,N_19639,N_20180);
or U24006 (N_24006,N_19939,N_20558);
xor U24007 (N_24007,N_19499,N_21471);
xnor U24008 (N_24008,N_21466,N_20891);
or U24009 (N_24009,N_20926,N_21043);
nand U24010 (N_24010,N_21326,N_20895);
nor U24011 (N_24011,N_21260,N_20579);
nor U24012 (N_24012,N_20765,N_20047);
or U24013 (N_24013,N_20003,N_19140);
xnor U24014 (N_24014,N_19420,N_21747);
nor U24015 (N_24015,N_21392,N_20728);
nand U24016 (N_24016,N_21563,N_18993);
nor U24017 (N_24017,N_19056,N_20536);
and U24018 (N_24018,N_21851,N_20543);
nor U24019 (N_24019,N_20634,N_20035);
or U24020 (N_24020,N_21197,N_19576);
nand U24021 (N_24021,N_20831,N_21200);
nand U24022 (N_24022,N_21419,N_21065);
or U24023 (N_24023,N_18793,N_19460);
or U24024 (N_24024,N_20559,N_19312);
and U24025 (N_24025,N_18921,N_20397);
or U24026 (N_24026,N_21302,N_21703);
nor U24027 (N_24027,N_21400,N_19440);
and U24028 (N_24028,N_19337,N_19275);
nand U24029 (N_24029,N_19663,N_19123);
xnor U24030 (N_24030,N_19683,N_20303);
nand U24031 (N_24031,N_21749,N_21522);
xor U24032 (N_24032,N_21561,N_20452);
xor U24033 (N_24033,N_21299,N_19494);
nand U24034 (N_24034,N_21123,N_20221);
and U24035 (N_24035,N_19782,N_21066);
and U24036 (N_24036,N_19265,N_21267);
and U24037 (N_24037,N_21309,N_21017);
nand U24038 (N_24038,N_19516,N_20875);
nor U24039 (N_24039,N_20054,N_20893);
or U24040 (N_24040,N_19211,N_20602);
or U24041 (N_24041,N_18994,N_20097);
and U24042 (N_24042,N_19730,N_18795);
nor U24043 (N_24043,N_19067,N_20700);
nand U24044 (N_24044,N_21018,N_19699);
xnor U24045 (N_24045,N_19523,N_20255);
and U24046 (N_24046,N_21756,N_19803);
and U24047 (N_24047,N_20959,N_20659);
nor U24048 (N_24048,N_21092,N_20975);
and U24049 (N_24049,N_21130,N_21532);
and U24050 (N_24050,N_21588,N_20414);
and U24051 (N_24051,N_20232,N_20855);
nand U24052 (N_24052,N_20965,N_21256);
xor U24053 (N_24053,N_21824,N_20657);
nand U24054 (N_24054,N_19660,N_21561);
nand U24055 (N_24055,N_20944,N_20170);
and U24056 (N_24056,N_21450,N_21654);
nand U24057 (N_24057,N_18951,N_19973);
or U24058 (N_24058,N_21315,N_18805);
nand U24059 (N_24059,N_21428,N_21514);
nand U24060 (N_24060,N_21567,N_21578);
nor U24061 (N_24061,N_18797,N_19922);
nand U24062 (N_24062,N_21285,N_20576);
and U24063 (N_24063,N_19763,N_20073);
xnor U24064 (N_24064,N_20500,N_20285);
nor U24065 (N_24065,N_20681,N_21637);
or U24066 (N_24066,N_20944,N_20231);
and U24067 (N_24067,N_19872,N_21062);
and U24068 (N_24068,N_18822,N_20504);
nand U24069 (N_24069,N_20481,N_20478);
and U24070 (N_24070,N_18989,N_20953);
or U24071 (N_24071,N_20696,N_20866);
xnor U24072 (N_24072,N_21548,N_19707);
nor U24073 (N_24073,N_21396,N_20298);
nor U24074 (N_24074,N_21822,N_18969);
nand U24075 (N_24075,N_19088,N_19125);
or U24076 (N_24076,N_19266,N_20852);
or U24077 (N_24077,N_21287,N_21258);
nor U24078 (N_24078,N_19808,N_20792);
or U24079 (N_24079,N_20537,N_21031);
nor U24080 (N_24080,N_20581,N_19074);
and U24081 (N_24081,N_19946,N_21075);
xor U24082 (N_24082,N_19901,N_19776);
nor U24083 (N_24083,N_20811,N_21734);
xnor U24084 (N_24084,N_21428,N_19632);
nand U24085 (N_24085,N_20893,N_19590);
xnor U24086 (N_24086,N_19301,N_19049);
and U24087 (N_24087,N_21832,N_21471);
nor U24088 (N_24088,N_20427,N_19107);
nand U24089 (N_24089,N_21854,N_18818);
xnor U24090 (N_24090,N_19440,N_21100);
nor U24091 (N_24091,N_21635,N_19240);
and U24092 (N_24092,N_21094,N_20270);
xnor U24093 (N_24093,N_20427,N_21867);
and U24094 (N_24094,N_18756,N_20640);
nor U24095 (N_24095,N_19162,N_20222);
or U24096 (N_24096,N_21317,N_19289);
or U24097 (N_24097,N_19308,N_20290);
nand U24098 (N_24098,N_20751,N_21535);
xor U24099 (N_24099,N_19799,N_19045);
nor U24100 (N_24100,N_21106,N_21493);
xnor U24101 (N_24101,N_20636,N_19164);
nor U24102 (N_24102,N_21368,N_21779);
nor U24103 (N_24103,N_21121,N_20362);
nor U24104 (N_24104,N_21118,N_21494);
nor U24105 (N_24105,N_21306,N_20839);
nor U24106 (N_24106,N_21648,N_19773);
or U24107 (N_24107,N_20265,N_19086);
or U24108 (N_24108,N_19361,N_21450);
and U24109 (N_24109,N_19376,N_19284);
nor U24110 (N_24110,N_19815,N_18868);
and U24111 (N_24111,N_18870,N_21710);
nor U24112 (N_24112,N_20132,N_19227);
nor U24113 (N_24113,N_20369,N_21051);
xnor U24114 (N_24114,N_19863,N_19857);
nor U24115 (N_24115,N_21077,N_21697);
nand U24116 (N_24116,N_19535,N_21316);
nor U24117 (N_24117,N_19134,N_19853);
nor U24118 (N_24118,N_21105,N_21390);
nor U24119 (N_24119,N_19878,N_20337);
nor U24120 (N_24120,N_18850,N_19676);
nand U24121 (N_24121,N_20887,N_20724);
nor U24122 (N_24122,N_19175,N_18779);
nor U24123 (N_24123,N_19971,N_20801);
nand U24124 (N_24124,N_21562,N_19688);
nand U24125 (N_24125,N_20698,N_21802);
nor U24126 (N_24126,N_20462,N_19049);
nor U24127 (N_24127,N_19562,N_20456);
or U24128 (N_24128,N_20340,N_19618);
nand U24129 (N_24129,N_20607,N_20092);
nand U24130 (N_24130,N_21301,N_20437);
or U24131 (N_24131,N_21398,N_21034);
or U24132 (N_24132,N_21294,N_19766);
and U24133 (N_24133,N_18991,N_19638);
and U24134 (N_24134,N_20486,N_21329);
nand U24135 (N_24135,N_19904,N_19058);
and U24136 (N_24136,N_21704,N_20800);
nand U24137 (N_24137,N_20800,N_20434);
nand U24138 (N_24138,N_21356,N_19920);
nor U24139 (N_24139,N_19498,N_19613);
and U24140 (N_24140,N_21716,N_19400);
nor U24141 (N_24141,N_19744,N_20398);
xnor U24142 (N_24142,N_19660,N_19111);
and U24143 (N_24143,N_19380,N_19471);
nand U24144 (N_24144,N_19956,N_21693);
nand U24145 (N_24145,N_19570,N_21085);
and U24146 (N_24146,N_20969,N_19387);
or U24147 (N_24147,N_19552,N_20647);
or U24148 (N_24148,N_21367,N_21846);
nor U24149 (N_24149,N_20335,N_19963);
nand U24150 (N_24150,N_20307,N_21683);
nor U24151 (N_24151,N_20496,N_18947);
nand U24152 (N_24152,N_20496,N_21190);
and U24153 (N_24153,N_20891,N_20093);
nor U24154 (N_24154,N_20822,N_18792);
and U24155 (N_24155,N_18847,N_21590);
and U24156 (N_24156,N_19705,N_19744);
or U24157 (N_24157,N_20317,N_19424);
and U24158 (N_24158,N_21647,N_20995);
or U24159 (N_24159,N_20138,N_19627);
or U24160 (N_24160,N_19176,N_20894);
or U24161 (N_24161,N_21130,N_19933);
and U24162 (N_24162,N_20213,N_19315);
xor U24163 (N_24163,N_20474,N_20869);
xor U24164 (N_24164,N_21484,N_19454);
nor U24165 (N_24165,N_19653,N_18987);
and U24166 (N_24166,N_19686,N_20749);
nor U24167 (N_24167,N_19401,N_19465);
and U24168 (N_24168,N_21301,N_18923);
nand U24169 (N_24169,N_20661,N_18991);
nand U24170 (N_24170,N_19993,N_21485);
or U24171 (N_24171,N_21072,N_21493);
and U24172 (N_24172,N_19236,N_20304);
nor U24173 (N_24173,N_20747,N_21326);
nor U24174 (N_24174,N_19962,N_18802);
xnor U24175 (N_24175,N_20891,N_20665);
and U24176 (N_24176,N_19416,N_20327);
or U24177 (N_24177,N_18991,N_20962);
or U24178 (N_24178,N_19062,N_20728);
or U24179 (N_24179,N_20768,N_21082);
or U24180 (N_24180,N_20549,N_18922);
and U24181 (N_24181,N_18939,N_20666);
nor U24182 (N_24182,N_19151,N_21120);
or U24183 (N_24183,N_20492,N_18908);
or U24184 (N_24184,N_20462,N_19008);
and U24185 (N_24185,N_19020,N_19786);
and U24186 (N_24186,N_19992,N_20172);
nor U24187 (N_24187,N_20471,N_19372);
and U24188 (N_24188,N_19881,N_19337);
nor U24189 (N_24189,N_19301,N_21361);
nand U24190 (N_24190,N_18862,N_20666);
and U24191 (N_24191,N_20244,N_19449);
nand U24192 (N_24192,N_19558,N_20350);
nor U24193 (N_24193,N_20980,N_19365);
or U24194 (N_24194,N_20281,N_19783);
and U24195 (N_24195,N_18904,N_21865);
and U24196 (N_24196,N_21778,N_20859);
and U24197 (N_24197,N_19775,N_21415);
or U24198 (N_24198,N_18868,N_20845);
or U24199 (N_24199,N_20304,N_19154);
and U24200 (N_24200,N_19521,N_21146);
nand U24201 (N_24201,N_21863,N_19216);
nor U24202 (N_24202,N_20056,N_21254);
nand U24203 (N_24203,N_19757,N_19695);
nand U24204 (N_24204,N_21237,N_19423);
nand U24205 (N_24205,N_20810,N_19027);
nand U24206 (N_24206,N_21739,N_19739);
nor U24207 (N_24207,N_20750,N_21383);
or U24208 (N_24208,N_21742,N_19286);
xor U24209 (N_24209,N_18937,N_19548);
nand U24210 (N_24210,N_21491,N_20284);
nor U24211 (N_24211,N_19017,N_18885);
nor U24212 (N_24212,N_20095,N_20886);
nor U24213 (N_24213,N_19473,N_20820);
and U24214 (N_24214,N_19893,N_21578);
nor U24215 (N_24215,N_20274,N_19319);
nand U24216 (N_24216,N_20542,N_20692);
and U24217 (N_24217,N_20153,N_19991);
nor U24218 (N_24218,N_18875,N_20291);
xnor U24219 (N_24219,N_20210,N_20930);
and U24220 (N_24220,N_21867,N_20044);
and U24221 (N_24221,N_19476,N_19993);
or U24222 (N_24222,N_18904,N_18862);
nor U24223 (N_24223,N_21530,N_20112);
nand U24224 (N_24224,N_19398,N_19332);
nor U24225 (N_24225,N_21800,N_19622);
or U24226 (N_24226,N_19079,N_20406);
and U24227 (N_24227,N_20661,N_19613);
nand U24228 (N_24228,N_21498,N_21558);
nor U24229 (N_24229,N_20708,N_19853);
xor U24230 (N_24230,N_18760,N_19991);
and U24231 (N_24231,N_20269,N_21487);
nand U24232 (N_24232,N_20502,N_21836);
nand U24233 (N_24233,N_19643,N_19588);
or U24234 (N_24234,N_19126,N_19528);
or U24235 (N_24235,N_20089,N_21573);
nor U24236 (N_24236,N_20673,N_21631);
nor U24237 (N_24237,N_21125,N_20928);
and U24238 (N_24238,N_20056,N_21724);
or U24239 (N_24239,N_18999,N_19257);
and U24240 (N_24240,N_20658,N_21439);
and U24241 (N_24241,N_20601,N_19844);
nor U24242 (N_24242,N_20062,N_20302);
nand U24243 (N_24243,N_21664,N_18955);
nor U24244 (N_24244,N_21864,N_20766);
nand U24245 (N_24245,N_20590,N_21455);
nand U24246 (N_24246,N_21101,N_20008);
and U24247 (N_24247,N_21871,N_19690);
or U24248 (N_24248,N_18756,N_19627);
nand U24249 (N_24249,N_19772,N_19027);
and U24250 (N_24250,N_21220,N_19355);
or U24251 (N_24251,N_20522,N_19416);
or U24252 (N_24252,N_19227,N_21199);
nor U24253 (N_24253,N_21420,N_19222);
nand U24254 (N_24254,N_20947,N_19115);
nand U24255 (N_24255,N_20135,N_19630);
xor U24256 (N_24256,N_19514,N_20022);
and U24257 (N_24257,N_20721,N_21784);
nand U24258 (N_24258,N_20232,N_21108);
nor U24259 (N_24259,N_20156,N_21631);
nor U24260 (N_24260,N_19965,N_19079);
nand U24261 (N_24261,N_19399,N_21630);
and U24262 (N_24262,N_21072,N_21137);
nand U24263 (N_24263,N_20149,N_20667);
xor U24264 (N_24264,N_20958,N_21164);
xnor U24265 (N_24265,N_20197,N_19451);
nor U24266 (N_24266,N_20816,N_18993);
or U24267 (N_24267,N_20893,N_21415);
nand U24268 (N_24268,N_19344,N_19381);
nor U24269 (N_24269,N_19477,N_21264);
and U24270 (N_24270,N_21627,N_20327);
and U24271 (N_24271,N_20555,N_18940);
nand U24272 (N_24272,N_20698,N_19526);
nand U24273 (N_24273,N_19077,N_19689);
or U24274 (N_24274,N_19494,N_20407);
nand U24275 (N_24275,N_18984,N_20219);
and U24276 (N_24276,N_20530,N_18853);
nor U24277 (N_24277,N_21211,N_19957);
or U24278 (N_24278,N_19317,N_18893);
nor U24279 (N_24279,N_20901,N_21565);
nand U24280 (N_24280,N_21213,N_19902);
or U24281 (N_24281,N_19566,N_20215);
and U24282 (N_24282,N_21715,N_18849);
nand U24283 (N_24283,N_21872,N_18837);
and U24284 (N_24284,N_21812,N_19276);
or U24285 (N_24285,N_20628,N_20090);
nor U24286 (N_24286,N_18910,N_19565);
xnor U24287 (N_24287,N_21775,N_20833);
and U24288 (N_24288,N_21163,N_19817);
nand U24289 (N_24289,N_21858,N_18788);
nand U24290 (N_24290,N_20012,N_21070);
nor U24291 (N_24291,N_20637,N_21037);
and U24292 (N_24292,N_21085,N_20743);
nand U24293 (N_24293,N_20903,N_19583);
and U24294 (N_24294,N_19974,N_19012);
nand U24295 (N_24295,N_20320,N_19940);
nand U24296 (N_24296,N_19236,N_21020);
nand U24297 (N_24297,N_18793,N_19016);
and U24298 (N_24298,N_18937,N_20913);
nand U24299 (N_24299,N_20844,N_20785);
xor U24300 (N_24300,N_20392,N_21523);
nor U24301 (N_24301,N_19575,N_19400);
nand U24302 (N_24302,N_20246,N_21291);
and U24303 (N_24303,N_19501,N_19391);
nor U24304 (N_24304,N_18879,N_19387);
or U24305 (N_24305,N_19011,N_21249);
or U24306 (N_24306,N_20393,N_20477);
xnor U24307 (N_24307,N_20821,N_21490);
nor U24308 (N_24308,N_20606,N_19544);
or U24309 (N_24309,N_21635,N_20882);
xor U24310 (N_24310,N_21159,N_21582);
or U24311 (N_24311,N_19572,N_19866);
and U24312 (N_24312,N_19790,N_20121);
nor U24313 (N_24313,N_21809,N_21017);
nor U24314 (N_24314,N_20795,N_19164);
xor U24315 (N_24315,N_18778,N_20034);
nand U24316 (N_24316,N_20756,N_20671);
nor U24317 (N_24317,N_20191,N_19495);
or U24318 (N_24318,N_21045,N_21082);
and U24319 (N_24319,N_19528,N_19623);
nand U24320 (N_24320,N_20526,N_19606);
and U24321 (N_24321,N_21739,N_21602);
nor U24322 (N_24322,N_20074,N_21612);
nand U24323 (N_24323,N_19274,N_20509);
and U24324 (N_24324,N_19206,N_21239);
nor U24325 (N_24325,N_19842,N_21258);
and U24326 (N_24326,N_20981,N_21064);
and U24327 (N_24327,N_19326,N_21229);
nand U24328 (N_24328,N_21758,N_20458);
and U24329 (N_24329,N_20185,N_21707);
nor U24330 (N_24330,N_18996,N_21190);
nand U24331 (N_24331,N_21172,N_18804);
or U24332 (N_24332,N_19512,N_19081);
nor U24333 (N_24333,N_20700,N_21866);
nand U24334 (N_24334,N_19655,N_20370);
nor U24335 (N_24335,N_20080,N_19958);
and U24336 (N_24336,N_20076,N_18881);
xnor U24337 (N_24337,N_21552,N_18989);
xor U24338 (N_24338,N_20166,N_21127);
nor U24339 (N_24339,N_19731,N_21162);
nor U24340 (N_24340,N_21309,N_19766);
nand U24341 (N_24341,N_20075,N_19198);
and U24342 (N_24342,N_21689,N_21221);
nor U24343 (N_24343,N_20715,N_21612);
nor U24344 (N_24344,N_19391,N_20413);
or U24345 (N_24345,N_18989,N_20858);
nand U24346 (N_24346,N_18773,N_18898);
nor U24347 (N_24347,N_20506,N_18897);
nand U24348 (N_24348,N_19260,N_20163);
and U24349 (N_24349,N_19619,N_21447);
nand U24350 (N_24350,N_21289,N_18900);
nand U24351 (N_24351,N_19478,N_20782);
or U24352 (N_24352,N_19682,N_21824);
nand U24353 (N_24353,N_19483,N_21226);
nand U24354 (N_24354,N_20722,N_19989);
and U24355 (N_24355,N_18828,N_19585);
nand U24356 (N_24356,N_19004,N_18851);
nor U24357 (N_24357,N_21101,N_20218);
nand U24358 (N_24358,N_21780,N_21004);
nand U24359 (N_24359,N_20870,N_18835);
nand U24360 (N_24360,N_21744,N_21419);
and U24361 (N_24361,N_19636,N_20270);
and U24362 (N_24362,N_18832,N_18837);
nand U24363 (N_24363,N_20920,N_20036);
nor U24364 (N_24364,N_20761,N_21572);
and U24365 (N_24365,N_20350,N_21152);
nand U24366 (N_24366,N_19936,N_19092);
nand U24367 (N_24367,N_21443,N_20944);
and U24368 (N_24368,N_19846,N_20348);
nand U24369 (N_24369,N_19172,N_19163);
and U24370 (N_24370,N_20739,N_21396);
and U24371 (N_24371,N_19019,N_21376);
nand U24372 (N_24372,N_20427,N_21618);
nand U24373 (N_24373,N_20526,N_20974);
xnor U24374 (N_24374,N_20152,N_20061);
nand U24375 (N_24375,N_19372,N_19502);
xnor U24376 (N_24376,N_19095,N_18917);
nor U24377 (N_24377,N_20960,N_20430);
nor U24378 (N_24378,N_19277,N_19999);
nand U24379 (N_24379,N_19298,N_21386);
or U24380 (N_24380,N_20674,N_21429);
xnor U24381 (N_24381,N_20075,N_18981);
or U24382 (N_24382,N_19031,N_20128);
nor U24383 (N_24383,N_21854,N_20996);
or U24384 (N_24384,N_20866,N_21724);
nor U24385 (N_24385,N_19905,N_19060);
nor U24386 (N_24386,N_20333,N_20866);
nor U24387 (N_24387,N_19968,N_20476);
nand U24388 (N_24388,N_19084,N_21045);
nand U24389 (N_24389,N_19770,N_19629);
and U24390 (N_24390,N_20226,N_19743);
nor U24391 (N_24391,N_21387,N_18964);
or U24392 (N_24392,N_19461,N_20966);
xor U24393 (N_24393,N_18794,N_18945);
nor U24394 (N_24394,N_18780,N_21077);
nor U24395 (N_24395,N_19127,N_21356);
or U24396 (N_24396,N_19449,N_18955);
nor U24397 (N_24397,N_21264,N_21626);
or U24398 (N_24398,N_18931,N_19794);
xnor U24399 (N_24399,N_19549,N_20973);
or U24400 (N_24400,N_20344,N_19397);
and U24401 (N_24401,N_19206,N_21132);
nor U24402 (N_24402,N_20905,N_20637);
nand U24403 (N_24403,N_20064,N_21027);
nor U24404 (N_24404,N_20819,N_20098);
and U24405 (N_24405,N_20903,N_20683);
and U24406 (N_24406,N_21141,N_21808);
nand U24407 (N_24407,N_21107,N_19070);
nor U24408 (N_24408,N_19030,N_19813);
and U24409 (N_24409,N_19659,N_20884);
or U24410 (N_24410,N_20043,N_20390);
or U24411 (N_24411,N_21361,N_18851);
and U24412 (N_24412,N_19714,N_18763);
and U24413 (N_24413,N_21214,N_19941);
or U24414 (N_24414,N_18815,N_19096);
xor U24415 (N_24415,N_18807,N_18851);
or U24416 (N_24416,N_18807,N_21162);
nand U24417 (N_24417,N_19955,N_19433);
or U24418 (N_24418,N_20881,N_20665);
xor U24419 (N_24419,N_20710,N_19580);
nand U24420 (N_24420,N_19515,N_20621);
nand U24421 (N_24421,N_20478,N_20573);
or U24422 (N_24422,N_21141,N_21039);
or U24423 (N_24423,N_20371,N_19057);
or U24424 (N_24424,N_21027,N_21140);
nor U24425 (N_24425,N_19595,N_19108);
nand U24426 (N_24426,N_21337,N_19657);
nor U24427 (N_24427,N_19657,N_21066);
xnor U24428 (N_24428,N_19757,N_19242);
nand U24429 (N_24429,N_20498,N_21500);
or U24430 (N_24430,N_20709,N_19661);
nor U24431 (N_24431,N_20803,N_20123);
and U24432 (N_24432,N_20796,N_19780);
xor U24433 (N_24433,N_19214,N_19198);
and U24434 (N_24434,N_21601,N_19906);
and U24435 (N_24435,N_19255,N_21767);
xnor U24436 (N_24436,N_19662,N_21764);
and U24437 (N_24437,N_20260,N_20824);
or U24438 (N_24438,N_21363,N_20754);
or U24439 (N_24439,N_21470,N_21600);
nand U24440 (N_24440,N_20424,N_19754);
or U24441 (N_24441,N_19582,N_20824);
and U24442 (N_24442,N_20809,N_19328);
or U24443 (N_24443,N_21225,N_21091);
and U24444 (N_24444,N_19204,N_20463);
nor U24445 (N_24445,N_19213,N_19496);
nand U24446 (N_24446,N_19507,N_19013);
and U24447 (N_24447,N_19558,N_19150);
nor U24448 (N_24448,N_19890,N_19818);
nand U24449 (N_24449,N_19914,N_18889);
nand U24450 (N_24450,N_19223,N_18962);
nand U24451 (N_24451,N_19201,N_21651);
and U24452 (N_24452,N_21234,N_20145);
nand U24453 (N_24453,N_19812,N_20876);
nor U24454 (N_24454,N_21873,N_20388);
and U24455 (N_24455,N_19136,N_21838);
nor U24456 (N_24456,N_19516,N_20152);
or U24457 (N_24457,N_19394,N_21377);
or U24458 (N_24458,N_20066,N_21283);
nor U24459 (N_24459,N_19726,N_20064);
nand U24460 (N_24460,N_21265,N_20692);
and U24461 (N_24461,N_19273,N_21833);
nor U24462 (N_24462,N_21154,N_21568);
xor U24463 (N_24463,N_21042,N_19903);
or U24464 (N_24464,N_21480,N_20166);
xor U24465 (N_24465,N_20390,N_20935);
or U24466 (N_24466,N_21393,N_19777);
nand U24467 (N_24467,N_21001,N_21136);
or U24468 (N_24468,N_19910,N_20388);
nor U24469 (N_24469,N_21341,N_19078);
or U24470 (N_24470,N_19370,N_21764);
nand U24471 (N_24471,N_20763,N_19988);
or U24472 (N_24472,N_19685,N_21479);
and U24473 (N_24473,N_21079,N_18787);
or U24474 (N_24474,N_20532,N_21138);
or U24475 (N_24475,N_19820,N_21584);
and U24476 (N_24476,N_19523,N_19948);
or U24477 (N_24477,N_21242,N_20520);
or U24478 (N_24478,N_21368,N_21833);
nor U24479 (N_24479,N_21579,N_18903);
and U24480 (N_24480,N_21648,N_20100);
nor U24481 (N_24481,N_19028,N_20923);
nand U24482 (N_24482,N_19209,N_20804);
or U24483 (N_24483,N_19588,N_19734);
nor U24484 (N_24484,N_20771,N_20539);
nor U24485 (N_24485,N_20554,N_21668);
or U24486 (N_24486,N_21348,N_20461);
nor U24487 (N_24487,N_19662,N_21254);
nor U24488 (N_24488,N_21582,N_20318);
or U24489 (N_24489,N_19430,N_20230);
xor U24490 (N_24490,N_21709,N_19761);
nor U24491 (N_24491,N_21452,N_19128);
or U24492 (N_24492,N_20392,N_20379);
nand U24493 (N_24493,N_20193,N_19126);
nand U24494 (N_24494,N_21424,N_20418);
or U24495 (N_24495,N_21514,N_19640);
nand U24496 (N_24496,N_19040,N_19146);
and U24497 (N_24497,N_21398,N_19948);
or U24498 (N_24498,N_19455,N_20959);
nand U24499 (N_24499,N_20243,N_18992);
nor U24500 (N_24500,N_19429,N_19676);
or U24501 (N_24501,N_21074,N_19313);
and U24502 (N_24502,N_19611,N_20387);
or U24503 (N_24503,N_19601,N_20193);
nor U24504 (N_24504,N_19372,N_21468);
or U24505 (N_24505,N_19558,N_19174);
nor U24506 (N_24506,N_19063,N_18854);
nor U24507 (N_24507,N_20190,N_21059);
xor U24508 (N_24508,N_21339,N_20806);
or U24509 (N_24509,N_19849,N_21366);
and U24510 (N_24510,N_20193,N_18786);
nand U24511 (N_24511,N_20079,N_19595);
and U24512 (N_24512,N_20139,N_19479);
and U24513 (N_24513,N_20023,N_20803);
or U24514 (N_24514,N_20295,N_19653);
nand U24515 (N_24515,N_20784,N_20779);
nand U24516 (N_24516,N_19836,N_19321);
nand U24517 (N_24517,N_21659,N_21313);
xnor U24518 (N_24518,N_18883,N_21624);
nand U24519 (N_24519,N_19291,N_21628);
and U24520 (N_24520,N_19712,N_19321);
and U24521 (N_24521,N_19423,N_19551);
nand U24522 (N_24522,N_19563,N_19358);
and U24523 (N_24523,N_20737,N_20270);
or U24524 (N_24524,N_21042,N_19908);
nor U24525 (N_24525,N_21608,N_20195);
nor U24526 (N_24526,N_20456,N_20236);
xnor U24527 (N_24527,N_19028,N_21661);
nand U24528 (N_24528,N_19941,N_18750);
or U24529 (N_24529,N_21760,N_19753);
nand U24530 (N_24530,N_20294,N_21807);
or U24531 (N_24531,N_21373,N_20357);
or U24532 (N_24532,N_19678,N_18871);
nand U24533 (N_24533,N_21564,N_20347);
or U24534 (N_24534,N_20640,N_19365);
nor U24535 (N_24535,N_20995,N_19995);
nor U24536 (N_24536,N_21712,N_19043);
and U24537 (N_24537,N_20582,N_21233);
nand U24538 (N_24538,N_18977,N_20285);
nand U24539 (N_24539,N_20860,N_19435);
and U24540 (N_24540,N_18915,N_19870);
nor U24541 (N_24541,N_19480,N_20751);
nor U24542 (N_24542,N_20547,N_21060);
and U24543 (N_24543,N_19777,N_21260);
nand U24544 (N_24544,N_21287,N_20453);
nor U24545 (N_24545,N_21377,N_19692);
nand U24546 (N_24546,N_18970,N_21774);
nor U24547 (N_24547,N_19308,N_20802);
nand U24548 (N_24548,N_20289,N_20185);
nor U24549 (N_24549,N_21643,N_19683);
or U24550 (N_24550,N_21417,N_19311);
nand U24551 (N_24551,N_21329,N_19542);
xnor U24552 (N_24552,N_19743,N_21091);
nor U24553 (N_24553,N_21177,N_18957);
and U24554 (N_24554,N_19422,N_21616);
nand U24555 (N_24555,N_20925,N_20187);
xnor U24556 (N_24556,N_21412,N_21738);
nor U24557 (N_24557,N_20584,N_21431);
or U24558 (N_24558,N_19989,N_19726);
or U24559 (N_24559,N_20886,N_18824);
and U24560 (N_24560,N_19267,N_20740);
nand U24561 (N_24561,N_20015,N_21045);
xor U24562 (N_24562,N_18850,N_19415);
nand U24563 (N_24563,N_20175,N_20776);
nand U24564 (N_24564,N_20620,N_20214);
xnor U24565 (N_24565,N_20414,N_20289);
nor U24566 (N_24566,N_20163,N_21187);
and U24567 (N_24567,N_19913,N_19401);
nand U24568 (N_24568,N_20410,N_20833);
nor U24569 (N_24569,N_20345,N_19597);
nor U24570 (N_24570,N_21583,N_21152);
nor U24571 (N_24571,N_20654,N_21019);
xnor U24572 (N_24572,N_20061,N_19146);
xnor U24573 (N_24573,N_21713,N_20877);
or U24574 (N_24574,N_19319,N_21506);
and U24575 (N_24575,N_19243,N_20881);
and U24576 (N_24576,N_19299,N_21735);
or U24577 (N_24577,N_21000,N_21541);
or U24578 (N_24578,N_20218,N_21053);
xnor U24579 (N_24579,N_21038,N_19969);
and U24580 (N_24580,N_20457,N_20960);
xor U24581 (N_24581,N_20943,N_21466);
nor U24582 (N_24582,N_20425,N_18907);
xnor U24583 (N_24583,N_21185,N_19165);
and U24584 (N_24584,N_20959,N_21671);
and U24585 (N_24585,N_19063,N_19685);
and U24586 (N_24586,N_20581,N_20679);
or U24587 (N_24587,N_21201,N_19614);
or U24588 (N_24588,N_20304,N_19314);
nand U24589 (N_24589,N_19216,N_21763);
nor U24590 (N_24590,N_18794,N_21601);
nand U24591 (N_24591,N_19227,N_20662);
or U24592 (N_24592,N_18906,N_21839);
or U24593 (N_24593,N_20300,N_20826);
and U24594 (N_24594,N_21557,N_18969);
nand U24595 (N_24595,N_20136,N_21204);
or U24596 (N_24596,N_20230,N_19125);
or U24597 (N_24597,N_21276,N_20655);
xor U24598 (N_24598,N_20832,N_19234);
or U24599 (N_24599,N_19605,N_18830);
or U24600 (N_24600,N_19796,N_20223);
or U24601 (N_24601,N_20605,N_18814);
or U24602 (N_24602,N_20549,N_21013);
and U24603 (N_24603,N_21702,N_21832);
nor U24604 (N_24604,N_19655,N_21208);
or U24605 (N_24605,N_21707,N_20007);
nand U24606 (N_24606,N_21714,N_19982);
nor U24607 (N_24607,N_20895,N_20477);
nor U24608 (N_24608,N_20521,N_19082);
nand U24609 (N_24609,N_19413,N_21052);
or U24610 (N_24610,N_21065,N_20849);
xnor U24611 (N_24611,N_19404,N_19611);
nor U24612 (N_24612,N_20269,N_20483);
nor U24613 (N_24613,N_18790,N_19970);
nor U24614 (N_24614,N_21708,N_21364);
and U24615 (N_24615,N_20761,N_21709);
and U24616 (N_24616,N_18902,N_20298);
xor U24617 (N_24617,N_20788,N_20542);
nor U24618 (N_24618,N_21018,N_18821);
nor U24619 (N_24619,N_19800,N_19013);
xnor U24620 (N_24620,N_21775,N_19858);
or U24621 (N_24621,N_20734,N_19005);
nor U24622 (N_24622,N_20354,N_21364);
nand U24623 (N_24623,N_21119,N_20772);
nor U24624 (N_24624,N_21436,N_20261);
or U24625 (N_24625,N_21313,N_19066);
xnor U24626 (N_24626,N_20989,N_21635);
and U24627 (N_24627,N_19492,N_19842);
and U24628 (N_24628,N_21331,N_21666);
or U24629 (N_24629,N_20794,N_20139);
or U24630 (N_24630,N_18771,N_19263);
or U24631 (N_24631,N_19160,N_20043);
or U24632 (N_24632,N_21429,N_20356);
or U24633 (N_24633,N_21649,N_20571);
or U24634 (N_24634,N_21831,N_19466);
and U24635 (N_24635,N_20085,N_20293);
or U24636 (N_24636,N_20459,N_20769);
and U24637 (N_24637,N_20625,N_20347);
and U24638 (N_24638,N_20393,N_21495);
nand U24639 (N_24639,N_21062,N_19547);
or U24640 (N_24640,N_21584,N_21801);
xnor U24641 (N_24641,N_19208,N_21669);
or U24642 (N_24642,N_20631,N_21768);
nand U24643 (N_24643,N_21814,N_20441);
and U24644 (N_24644,N_20744,N_21261);
xnor U24645 (N_24645,N_20594,N_21747);
nand U24646 (N_24646,N_19986,N_21622);
or U24647 (N_24647,N_20321,N_19049);
or U24648 (N_24648,N_18967,N_20216);
nor U24649 (N_24649,N_18841,N_21866);
and U24650 (N_24650,N_20349,N_18757);
or U24651 (N_24651,N_21288,N_20204);
xnor U24652 (N_24652,N_19526,N_21580);
xnor U24653 (N_24653,N_19539,N_21646);
xnor U24654 (N_24654,N_20497,N_20363);
xor U24655 (N_24655,N_20970,N_19637);
xor U24656 (N_24656,N_21249,N_20253);
nor U24657 (N_24657,N_19998,N_21718);
nand U24658 (N_24658,N_21732,N_20466);
and U24659 (N_24659,N_21258,N_19031);
and U24660 (N_24660,N_21856,N_20401);
xnor U24661 (N_24661,N_21522,N_18761);
nor U24662 (N_24662,N_19751,N_19462);
and U24663 (N_24663,N_20445,N_20053);
nand U24664 (N_24664,N_19934,N_19744);
nor U24665 (N_24665,N_21035,N_18874);
nor U24666 (N_24666,N_20510,N_20045);
and U24667 (N_24667,N_21167,N_21178);
nor U24668 (N_24668,N_21140,N_20185);
nor U24669 (N_24669,N_20407,N_18958);
nor U24670 (N_24670,N_20490,N_20046);
and U24671 (N_24671,N_21382,N_20628);
and U24672 (N_24672,N_19762,N_20747);
nand U24673 (N_24673,N_18775,N_20327);
and U24674 (N_24674,N_21201,N_20738);
nor U24675 (N_24675,N_19849,N_19361);
nand U24676 (N_24676,N_19059,N_21210);
xor U24677 (N_24677,N_21187,N_19361);
nand U24678 (N_24678,N_20657,N_21651);
and U24679 (N_24679,N_19548,N_19148);
nor U24680 (N_24680,N_19527,N_18952);
or U24681 (N_24681,N_18818,N_20492);
nor U24682 (N_24682,N_21464,N_18779);
or U24683 (N_24683,N_21248,N_21249);
nor U24684 (N_24684,N_19751,N_20807);
nor U24685 (N_24685,N_21812,N_21355);
nor U24686 (N_24686,N_20584,N_20992);
nand U24687 (N_24687,N_19901,N_20516);
and U24688 (N_24688,N_21299,N_20120);
nor U24689 (N_24689,N_20634,N_21547);
and U24690 (N_24690,N_21640,N_21575);
nor U24691 (N_24691,N_20498,N_19941);
or U24692 (N_24692,N_20580,N_19722);
and U24693 (N_24693,N_20708,N_19865);
nor U24694 (N_24694,N_19237,N_20889);
and U24695 (N_24695,N_20383,N_20389);
or U24696 (N_24696,N_20632,N_20152);
or U24697 (N_24697,N_19523,N_21568);
nand U24698 (N_24698,N_19281,N_19825);
or U24699 (N_24699,N_20518,N_20630);
and U24700 (N_24700,N_21013,N_19507);
nand U24701 (N_24701,N_20940,N_21071);
nor U24702 (N_24702,N_19044,N_19747);
nand U24703 (N_24703,N_19297,N_19084);
nor U24704 (N_24704,N_20783,N_19980);
or U24705 (N_24705,N_18761,N_21365);
or U24706 (N_24706,N_19084,N_19456);
and U24707 (N_24707,N_21610,N_21343);
or U24708 (N_24708,N_20442,N_21043);
nand U24709 (N_24709,N_21419,N_18996);
or U24710 (N_24710,N_19951,N_20636);
and U24711 (N_24711,N_20522,N_20416);
and U24712 (N_24712,N_19733,N_20109);
nor U24713 (N_24713,N_20428,N_20782);
nor U24714 (N_24714,N_18943,N_20113);
xor U24715 (N_24715,N_20556,N_19211);
or U24716 (N_24716,N_21489,N_20402);
and U24717 (N_24717,N_20944,N_19599);
and U24718 (N_24718,N_20678,N_19931);
or U24719 (N_24719,N_19788,N_21866);
xor U24720 (N_24720,N_20951,N_19500);
xor U24721 (N_24721,N_21743,N_21491);
and U24722 (N_24722,N_19689,N_20217);
and U24723 (N_24723,N_21318,N_19820);
and U24724 (N_24724,N_20741,N_21481);
nor U24725 (N_24725,N_21792,N_20151);
or U24726 (N_24726,N_21164,N_20685);
nor U24727 (N_24727,N_18872,N_19551);
xor U24728 (N_24728,N_20737,N_18789);
and U24729 (N_24729,N_20606,N_18920);
nand U24730 (N_24730,N_21596,N_20395);
nand U24731 (N_24731,N_20716,N_19576);
and U24732 (N_24732,N_19866,N_19475);
or U24733 (N_24733,N_20018,N_20779);
and U24734 (N_24734,N_20931,N_18978);
or U24735 (N_24735,N_20125,N_19321);
or U24736 (N_24736,N_21868,N_19036);
or U24737 (N_24737,N_19362,N_19344);
and U24738 (N_24738,N_19513,N_21826);
nand U24739 (N_24739,N_21873,N_20852);
nor U24740 (N_24740,N_19644,N_21844);
and U24741 (N_24741,N_21776,N_20992);
nor U24742 (N_24742,N_19281,N_20840);
or U24743 (N_24743,N_20061,N_20787);
and U24744 (N_24744,N_20616,N_21628);
and U24745 (N_24745,N_20797,N_21256);
nor U24746 (N_24746,N_18916,N_20196);
nand U24747 (N_24747,N_20337,N_19554);
nand U24748 (N_24748,N_21231,N_20913);
nand U24749 (N_24749,N_20561,N_20910);
and U24750 (N_24750,N_19370,N_21199);
nand U24751 (N_24751,N_19036,N_21387);
nand U24752 (N_24752,N_20861,N_19568);
or U24753 (N_24753,N_20890,N_21373);
or U24754 (N_24754,N_20771,N_20407);
xor U24755 (N_24755,N_19698,N_19427);
or U24756 (N_24756,N_21842,N_19707);
nand U24757 (N_24757,N_19861,N_21627);
and U24758 (N_24758,N_19692,N_18849);
nor U24759 (N_24759,N_20636,N_19975);
nand U24760 (N_24760,N_18764,N_19608);
nand U24761 (N_24761,N_21551,N_19654);
and U24762 (N_24762,N_19703,N_21678);
nand U24763 (N_24763,N_19154,N_19543);
and U24764 (N_24764,N_20032,N_21187);
xor U24765 (N_24765,N_21007,N_21778);
nor U24766 (N_24766,N_19141,N_19416);
and U24767 (N_24767,N_19410,N_20604);
nand U24768 (N_24768,N_20440,N_20705);
nor U24769 (N_24769,N_18919,N_19560);
and U24770 (N_24770,N_20407,N_20976);
nand U24771 (N_24771,N_19492,N_20284);
nor U24772 (N_24772,N_20930,N_20222);
nand U24773 (N_24773,N_20930,N_18963);
and U24774 (N_24774,N_19258,N_18919);
nand U24775 (N_24775,N_21043,N_20986);
and U24776 (N_24776,N_20738,N_20210);
or U24777 (N_24777,N_21393,N_19243);
xor U24778 (N_24778,N_20378,N_19271);
nand U24779 (N_24779,N_18901,N_20604);
and U24780 (N_24780,N_21667,N_20811);
xnor U24781 (N_24781,N_20431,N_20856);
and U24782 (N_24782,N_21597,N_19646);
nand U24783 (N_24783,N_20040,N_20878);
nor U24784 (N_24784,N_20623,N_18826);
and U24785 (N_24785,N_21643,N_19036);
or U24786 (N_24786,N_21385,N_21605);
xor U24787 (N_24787,N_19790,N_19062);
and U24788 (N_24788,N_20363,N_21308);
nor U24789 (N_24789,N_20635,N_19162);
or U24790 (N_24790,N_20992,N_18810);
nor U24791 (N_24791,N_20804,N_19417);
nor U24792 (N_24792,N_20522,N_21753);
and U24793 (N_24793,N_21166,N_19583);
nor U24794 (N_24794,N_20550,N_21828);
and U24795 (N_24795,N_20760,N_20230);
nand U24796 (N_24796,N_19511,N_19443);
and U24797 (N_24797,N_18783,N_20297);
and U24798 (N_24798,N_20855,N_20092);
or U24799 (N_24799,N_19348,N_19702);
nor U24800 (N_24800,N_20660,N_19546);
nand U24801 (N_24801,N_19767,N_19144);
nor U24802 (N_24802,N_20448,N_20801);
nor U24803 (N_24803,N_19719,N_20064);
xor U24804 (N_24804,N_19053,N_21790);
nand U24805 (N_24805,N_21153,N_18914);
or U24806 (N_24806,N_21401,N_21662);
nor U24807 (N_24807,N_21307,N_21548);
and U24808 (N_24808,N_19950,N_19812);
nand U24809 (N_24809,N_19730,N_20271);
nand U24810 (N_24810,N_20287,N_20088);
or U24811 (N_24811,N_19029,N_21196);
nor U24812 (N_24812,N_20181,N_20428);
nand U24813 (N_24813,N_19976,N_19962);
nand U24814 (N_24814,N_19336,N_21519);
xor U24815 (N_24815,N_21784,N_19903);
and U24816 (N_24816,N_19240,N_19884);
nor U24817 (N_24817,N_20686,N_20002);
and U24818 (N_24818,N_20836,N_19503);
nor U24819 (N_24819,N_19946,N_21179);
or U24820 (N_24820,N_21804,N_19402);
nand U24821 (N_24821,N_20302,N_19173);
nand U24822 (N_24822,N_21551,N_20744);
and U24823 (N_24823,N_19942,N_19153);
nor U24824 (N_24824,N_20516,N_19408);
nor U24825 (N_24825,N_21462,N_19769);
or U24826 (N_24826,N_19603,N_19065);
nand U24827 (N_24827,N_20828,N_19354);
and U24828 (N_24828,N_21643,N_20701);
and U24829 (N_24829,N_20294,N_19194);
or U24830 (N_24830,N_19671,N_20725);
nand U24831 (N_24831,N_20464,N_20434);
or U24832 (N_24832,N_20077,N_20537);
nor U24833 (N_24833,N_19779,N_19455);
or U24834 (N_24834,N_21731,N_19752);
and U24835 (N_24835,N_19862,N_20180);
nand U24836 (N_24836,N_19537,N_20042);
and U24837 (N_24837,N_19869,N_19295);
or U24838 (N_24838,N_20942,N_19548);
nand U24839 (N_24839,N_19521,N_21268);
and U24840 (N_24840,N_18999,N_21378);
or U24841 (N_24841,N_21631,N_20868);
xor U24842 (N_24842,N_19665,N_21442);
nor U24843 (N_24843,N_20670,N_19989);
nor U24844 (N_24844,N_19247,N_19003);
or U24845 (N_24845,N_21700,N_20657);
or U24846 (N_24846,N_19792,N_21003);
nand U24847 (N_24847,N_18756,N_19432);
nand U24848 (N_24848,N_20218,N_19277);
nand U24849 (N_24849,N_20126,N_21824);
or U24850 (N_24850,N_20590,N_20258);
nand U24851 (N_24851,N_21299,N_21475);
nand U24852 (N_24852,N_19108,N_20978);
nor U24853 (N_24853,N_20285,N_20873);
xor U24854 (N_24854,N_20089,N_18785);
nor U24855 (N_24855,N_19190,N_19951);
and U24856 (N_24856,N_20734,N_19825);
and U24857 (N_24857,N_21427,N_19061);
nand U24858 (N_24858,N_18959,N_21170);
nor U24859 (N_24859,N_20000,N_19803);
or U24860 (N_24860,N_21431,N_21472);
or U24861 (N_24861,N_19970,N_19547);
or U24862 (N_24862,N_19199,N_21112);
or U24863 (N_24863,N_19147,N_20338);
nand U24864 (N_24864,N_18923,N_19232);
or U24865 (N_24865,N_19583,N_20034);
nand U24866 (N_24866,N_21628,N_21249);
or U24867 (N_24867,N_21552,N_19296);
xor U24868 (N_24868,N_20995,N_20964);
nor U24869 (N_24869,N_20963,N_20631);
nand U24870 (N_24870,N_21073,N_20337);
and U24871 (N_24871,N_19973,N_19971);
and U24872 (N_24872,N_19081,N_19375);
and U24873 (N_24873,N_19155,N_19937);
and U24874 (N_24874,N_20395,N_18969);
nor U24875 (N_24875,N_21720,N_19489);
or U24876 (N_24876,N_18971,N_21613);
nand U24877 (N_24877,N_20274,N_21300);
or U24878 (N_24878,N_19921,N_21427);
xor U24879 (N_24879,N_20268,N_20308);
and U24880 (N_24880,N_19670,N_19701);
and U24881 (N_24881,N_21451,N_20397);
nand U24882 (N_24882,N_18833,N_21001);
or U24883 (N_24883,N_19305,N_19449);
nand U24884 (N_24884,N_19938,N_18769);
nand U24885 (N_24885,N_20071,N_21790);
nor U24886 (N_24886,N_19434,N_19378);
nand U24887 (N_24887,N_19158,N_19833);
and U24888 (N_24888,N_21833,N_21238);
nor U24889 (N_24889,N_21768,N_19751);
nand U24890 (N_24890,N_20311,N_18861);
and U24891 (N_24891,N_20828,N_21769);
or U24892 (N_24892,N_21072,N_21684);
and U24893 (N_24893,N_20118,N_19004);
or U24894 (N_24894,N_21264,N_19706);
nor U24895 (N_24895,N_20406,N_20010);
nand U24896 (N_24896,N_18902,N_19909);
and U24897 (N_24897,N_21445,N_20818);
xor U24898 (N_24898,N_20535,N_21132);
nor U24899 (N_24899,N_19929,N_20403);
xor U24900 (N_24900,N_21104,N_18804);
or U24901 (N_24901,N_21757,N_19747);
nor U24902 (N_24902,N_21674,N_19537);
xnor U24903 (N_24903,N_19072,N_20199);
or U24904 (N_24904,N_19177,N_20366);
and U24905 (N_24905,N_20051,N_19371);
nand U24906 (N_24906,N_21735,N_21090);
and U24907 (N_24907,N_21256,N_20236);
nand U24908 (N_24908,N_19324,N_21567);
and U24909 (N_24909,N_19255,N_19233);
nand U24910 (N_24910,N_20213,N_21635);
nor U24911 (N_24911,N_20953,N_20365);
and U24912 (N_24912,N_21359,N_20334);
or U24913 (N_24913,N_21378,N_21847);
nor U24914 (N_24914,N_21487,N_20481);
nand U24915 (N_24915,N_21564,N_19078);
or U24916 (N_24916,N_18776,N_19634);
and U24917 (N_24917,N_21787,N_20337);
and U24918 (N_24918,N_19805,N_20871);
or U24919 (N_24919,N_19519,N_18881);
nand U24920 (N_24920,N_20622,N_21014);
and U24921 (N_24921,N_20692,N_21316);
or U24922 (N_24922,N_20071,N_21421);
nor U24923 (N_24923,N_19128,N_19103);
and U24924 (N_24924,N_20986,N_18842);
nand U24925 (N_24925,N_20992,N_20579);
nand U24926 (N_24926,N_20970,N_20575);
xor U24927 (N_24927,N_21498,N_21094);
nor U24928 (N_24928,N_20026,N_21211);
nor U24929 (N_24929,N_21031,N_19922);
or U24930 (N_24930,N_21626,N_21644);
nor U24931 (N_24931,N_21865,N_19656);
nor U24932 (N_24932,N_19977,N_20458);
and U24933 (N_24933,N_20357,N_21285);
nand U24934 (N_24934,N_19270,N_21282);
and U24935 (N_24935,N_19771,N_21555);
nor U24936 (N_24936,N_20246,N_20780);
nor U24937 (N_24937,N_19524,N_20406);
and U24938 (N_24938,N_19021,N_20732);
nand U24939 (N_24939,N_20550,N_21192);
and U24940 (N_24940,N_19525,N_20909);
nand U24941 (N_24941,N_19980,N_20761);
xor U24942 (N_24942,N_21491,N_21410);
and U24943 (N_24943,N_19882,N_21005);
nor U24944 (N_24944,N_20288,N_19257);
nand U24945 (N_24945,N_21438,N_20733);
or U24946 (N_24946,N_19047,N_19799);
and U24947 (N_24947,N_21710,N_18828);
nor U24948 (N_24948,N_20155,N_20066);
nor U24949 (N_24949,N_21115,N_21765);
and U24950 (N_24950,N_21873,N_19796);
or U24951 (N_24951,N_20396,N_21438);
or U24952 (N_24952,N_21212,N_19251);
and U24953 (N_24953,N_18965,N_21377);
nand U24954 (N_24954,N_21096,N_19154);
nand U24955 (N_24955,N_19552,N_21436);
nand U24956 (N_24956,N_21289,N_20795);
nand U24957 (N_24957,N_20125,N_21270);
nor U24958 (N_24958,N_19341,N_20439);
nor U24959 (N_24959,N_18945,N_20664);
nand U24960 (N_24960,N_19500,N_18819);
nor U24961 (N_24961,N_19163,N_19022);
nand U24962 (N_24962,N_18956,N_19910);
and U24963 (N_24963,N_19868,N_21870);
xor U24964 (N_24964,N_20451,N_19452);
nor U24965 (N_24965,N_18758,N_20035);
nand U24966 (N_24966,N_20667,N_19947);
and U24967 (N_24967,N_18841,N_21400);
or U24968 (N_24968,N_18872,N_20549);
or U24969 (N_24969,N_19192,N_19304);
or U24970 (N_24970,N_20950,N_20481);
nand U24971 (N_24971,N_21569,N_21798);
nand U24972 (N_24972,N_20893,N_20624);
nor U24973 (N_24973,N_21179,N_19647);
nand U24974 (N_24974,N_19361,N_21371);
nor U24975 (N_24975,N_18814,N_18800);
nor U24976 (N_24976,N_20178,N_20784);
or U24977 (N_24977,N_19566,N_19335);
and U24978 (N_24978,N_20796,N_21627);
nand U24979 (N_24979,N_19204,N_21281);
or U24980 (N_24980,N_20346,N_19231);
or U24981 (N_24981,N_20806,N_19684);
and U24982 (N_24982,N_19552,N_20779);
nor U24983 (N_24983,N_19990,N_21387);
nor U24984 (N_24984,N_19192,N_20588);
and U24985 (N_24985,N_20377,N_20275);
nor U24986 (N_24986,N_20060,N_20030);
or U24987 (N_24987,N_19421,N_20787);
nor U24988 (N_24988,N_20128,N_20489);
or U24989 (N_24989,N_19108,N_19858);
nand U24990 (N_24990,N_20884,N_19089);
and U24991 (N_24991,N_20008,N_19234);
or U24992 (N_24992,N_20735,N_21586);
nand U24993 (N_24993,N_20163,N_20368);
nor U24994 (N_24994,N_19903,N_21279);
and U24995 (N_24995,N_19441,N_19723);
nor U24996 (N_24996,N_21813,N_19158);
xor U24997 (N_24997,N_18837,N_20371);
or U24998 (N_24998,N_21827,N_20868);
or U24999 (N_24999,N_20946,N_20352);
xnor UO_0 (O_0,N_23914,N_23355);
nor UO_1 (O_1,N_22372,N_24164);
or UO_2 (O_2,N_22409,N_23558);
nand UO_3 (O_3,N_23305,N_24022);
nor UO_4 (O_4,N_23237,N_24797);
nand UO_5 (O_5,N_22319,N_24477);
and UO_6 (O_6,N_22887,N_22877);
or UO_7 (O_7,N_24306,N_24557);
and UO_8 (O_8,N_23662,N_24648);
nor UO_9 (O_9,N_23204,N_24357);
nand UO_10 (O_10,N_23924,N_23654);
and UO_11 (O_11,N_24624,N_22453);
nor UO_12 (O_12,N_23025,N_23438);
and UO_13 (O_13,N_24345,N_22296);
xnor UO_14 (O_14,N_24805,N_24770);
nor UO_15 (O_15,N_22027,N_24969);
xor UO_16 (O_16,N_23306,N_22418);
or UO_17 (O_17,N_22661,N_23968);
or UO_18 (O_18,N_23883,N_22899);
nand UO_19 (O_19,N_23314,N_22175);
nor UO_20 (O_20,N_24577,N_22898);
nand UO_21 (O_21,N_22591,N_22184);
nand UO_22 (O_22,N_23313,N_23343);
nor UO_23 (O_23,N_23118,N_23207);
nand UO_24 (O_24,N_22406,N_24752);
or UO_25 (O_25,N_24379,N_22224);
and UO_26 (O_26,N_22645,N_23031);
and UO_27 (O_27,N_23960,N_22426);
and UO_28 (O_28,N_21956,N_22618);
xor UO_29 (O_29,N_24513,N_22068);
and UO_30 (O_30,N_22365,N_22780);
or UO_31 (O_31,N_22346,N_24524);
or UO_32 (O_32,N_24413,N_22366);
nand UO_33 (O_33,N_24330,N_24963);
nor UO_34 (O_34,N_24548,N_22929);
and UO_35 (O_35,N_24251,N_24849);
xnor UO_36 (O_36,N_22496,N_24394);
nor UO_37 (O_37,N_22157,N_22022);
nand UO_38 (O_38,N_23178,N_24706);
nand UO_39 (O_39,N_22716,N_22676);
or UO_40 (O_40,N_24593,N_22480);
and UO_41 (O_41,N_23901,N_22606);
or UO_42 (O_42,N_21944,N_23231);
or UO_43 (O_43,N_22949,N_22578);
and UO_44 (O_44,N_23564,N_22544);
and UO_45 (O_45,N_22803,N_22468);
or UO_46 (O_46,N_24917,N_24173);
or UO_47 (O_47,N_24886,N_24728);
nor UO_48 (O_48,N_24778,N_24180);
nand UO_49 (O_49,N_24630,N_23711);
nand UO_50 (O_50,N_22793,N_24780);
nor UO_51 (O_51,N_22718,N_24262);
and UO_52 (O_52,N_22145,N_23021);
and UO_53 (O_53,N_22056,N_24584);
and UO_54 (O_54,N_23106,N_23568);
xnor UO_55 (O_55,N_24182,N_24922);
or UO_56 (O_56,N_23104,N_23296);
or UO_57 (O_57,N_23257,N_22118);
nor UO_58 (O_58,N_22125,N_22099);
nor UO_59 (O_59,N_23605,N_22592);
nor UO_60 (O_60,N_22279,N_22080);
or UO_61 (O_61,N_24415,N_21903);
or UO_62 (O_62,N_22684,N_22045);
or UO_63 (O_63,N_23395,N_22124);
nand UO_64 (O_64,N_24505,N_22412);
nor UO_65 (O_65,N_24263,N_23202);
or UO_66 (O_66,N_24581,N_24384);
nor UO_67 (O_67,N_22422,N_24564);
and UO_68 (O_68,N_23818,N_22802);
or UO_69 (O_69,N_22156,N_23548);
or UO_70 (O_70,N_23693,N_24868);
and UO_71 (O_71,N_24785,N_24095);
and UO_72 (O_72,N_24240,N_22892);
nor UO_73 (O_73,N_21963,N_22138);
xor UO_74 (O_74,N_23732,N_22910);
nand UO_75 (O_75,N_22518,N_24021);
or UO_76 (O_76,N_23199,N_24081);
nor UO_77 (O_77,N_22262,N_23612);
nand UO_78 (O_78,N_23926,N_22729);
nand UO_79 (O_79,N_23132,N_22546);
and UO_80 (O_80,N_22069,N_22536);
nor UO_81 (O_81,N_22404,N_22007);
nand UO_82 (O_82,N_23990,N_22025);
or UO_83 (O_83,N_24586,N_21886);
or UO_84 (O_84,N_24450,N_22074);
and UO_85 (O_85,N_24799,N_22355);
and UO_86 (O_86,N_22927,N_23386);
nor UO_87 (O_87,N_24439,N_23403);
nand UO_88 (O_88,N_22013,N_24016);
nor UO_89 (O_89,N_22547,N_24430);
nor UO_90 (O_90,N_24762,N_23004);
nor UO_91 (O_91,N_24209,N_24870);
nand UO_92 (O_92,N_22221,N_24665);
or UO_93 (O_93,N_24709,N_24918);
nor UO_94 (O_94,N_23093,N_22416);
nor UO_95 (O_95,N_24984,N_22255);
or UO_96 (O_96,N_23371,N_22072);
nor UO_97 (O_97,N_23534,N_23201);
xnor UO_98 (O_98,N_22754,N_21922);
and UO_99 (O_99,N_24539,N_23253);
nand UO_100 (O_100,N_23051,N_23293);
and UO_101 (O_101,N_23978,N_23298);
nor UO_102 (O_102,N_22467,N_23733);
nor UO_103 (O_103,N_24769,N_22227);
nand UO_104 (O_104,N_23047,N_24526);
nor UO_105 (O_105,N_22897,N_23740);
nand UO_106 (O_106,N_23946,N_23414);
and UO_107 (O_107,N_22644,N_23663);
nand UO_108 (O_108,N_24832,N_24606);
or UO_109 (O_109,N_22024,N_24879);
and UO_110 (O_110,N_23328,N_22539);
nand UO_111 (O_111,N_23085,N_24236);
nor UO_112 (O_112,N_23811,N_24775);
or UO_113 (O_113,N_24342,N_24928);
and UO_114 (O_114,N_22843,N_24206);
and UO_115 (O_115,N_24341,N_22607);
nand UO_116 (O_116,N_23760,N_23768);
or UO_117 (O_117,N_23060,N_22253);
and UO_118 (O_118,N_22408,N_21964);
nand UO_119 (O_119,N_24566,N_22169);
and UO_120 (O_120,N_23727,N_21883);
nand UO_121 (O_121,N_22706,N_23723);
or UO_122 (O_122,N_23420,N_22581);
xor UO_123 (O_123,N_22593,N_23588);
nand UO_124 (O_124,N_22839,N_24226);
and UO_125 (O_125,N_22755,N_22904);
and UO_126 (O_126,N_24090,N_23792);
nand UO_127 (O_127,N_23890,N_24239);
and UO_128 (O_128,N_22267,N_24625);
or UO_129 (O_129,N_23412,N_22776);
or UO_130 (O_130,N_22957,N_23376);
or UO_131 (O_131,N_22598,N_24714);
nor UO_132 (O_132,N_23073,N_22541);
nor UO_133 (O_133,N_23399,N_24175);
nand UO_134 (O_134,N_23142,N_22719);
or UO_135 (O_135,N_24827,N_22482);
nor UO_136 (O_136,N_22713,N_23533);
nand UO_137 (O_137,N_23868,N_24145);
and UO_138 (O_138,N_23056,N_21986);
xnor UO_139 (O_139,N_24733,N_23308);
xnor UO_140 (O_140,N_23489,N_24196);
and UO_141 (O_141,N_24616,N_22924);
nor UO_142 (O_142,N_24372,N_23666);
nand UO_143 (O_143,N_24587,N_23200);
and UO_144 (O_144,N_23180,N_22316);
nand UO_145 (O_145,N_24949,N_21904);
and UO_146 (O_146,N_22911,N_23170);
nand UO_147 (O_147,N_21995,N_23432);
and UO_148 (O_148,N_22251,N_24700);
or UO_149 (O_149,N_22167,N_22178);
nand UO_150 (O_150,N_24461,N_22309);
nand UO_151 (O_151,N_24633,N_23444);
nor UO_152 (O_152,N_22801,N_24193);
nor UO_153 (O_153,N_23808,N_22234);
and UO_154 (O_154,N_22306,N_22509);
and UO_155 (O_155,N_23235,N_24109);
and UO_156 (O_156,N_22739,N_22465);
and UO_157 (O_157,N_24781,N_24426);
nor UO_158 (O_158,N_24754,N_22762);
nand UO_159 (O_159,N_23518,N_22486);
and UO_160 (O_160,N_23363,N_24722);
and UO_161 (O_161,N_22525,N_22474);
or UO_162 (O_162,N_23501,N_22935);
or UO_163 (O_163,N_23135,N_24594);
xor UO_164 (O_164,N_23687,N_21941);
or UO_165 (O_165,N_24340,N_23148);
or UO_166 (O_166,N_22636,N_23222);
or UO_167 (O_167,N_23155,N_22471);
or UO_168 (O_168,N_23684,N_24598);
and UO_169 (O_169,N_22726,N_23380);
nand UO_170 (O_170,N_23767,N_23105);
and UO_171 (O_171,N_22140,N_23023);
xor UO_172 (O_172,N_22494,N_22413);
or UO_173 (O_173,N_24067,N_23160);
nand UO_174 (O_174,N_22315,N_24100);
nand UO_175 (O_175,N_24739,N_23973);
nand UO_176 (O_176,N_22747,N_23712);
nor UO_177 (O_177,N_24491,N_23166);
nor UO_178 (O_178,N_22815,N_21960);
or UO_179 (O_179,N_24831,N_22604);
and UO_180 (O_180,N_22102,N_21950);
and UO_181 (O_181,N_24147,N_22048);
nor UO_182 (O_182,N_22545,N_24271);
nor UO_183 (O_183,N_22003,N_23778);
xnor UO_184 (O_184,N_23907,N_24128);
nand UO_185 (O_185,N_24623,N_24891);
nand UO_186 (O_186,N_22625,N_23941);
nor UO_187 (O_187,N_24853,N_24774);
xor UO_188 (O_188,N_23967,N_24794);
nor UO_189 (O_189,N_22236,N_23485);
nor UO_190 (O_190,N_24458,N_22724);
or UO_191 (O_191,N_24688,N_22039);
xnor UO_192 (O_192,N_23702,N_22415);
or UO_193 (O_193,N_22216,N_22520);
nor UO_194 (O_194,N_24446,N_24899);
or UO_195 (O_195,N_22475,N_21939);
nand UO_196 (O_196,N_24315,N_23992);
nand UO_197 (O_197,N_22497,N_22466);
nand UO_198 (O_198,N_22531,N_24523);
or UO_199 (O_199,N_23350,N_22344);
or UO_200 (O_200,N_22798,N_22026);
nor UO_201 (O_201,N_22381,N_24936);
nor UO_202 (O_202,N_23841,N_22063);
xnor UO_203 (O_203,N_23545,N_24708);
xnor UO_204 (O_204,N_24117,N_23896);
or UO_205 (O_205,N_24179,N_22004);
or UO_206 (O_206,N_23365,N_23109);
nand UO_207 (O_207,N_23950,N_23310);
and UO_208 (O_208,N_24821,N_24144);
or UO_209 (O_209,N_22860,N_23301);
nand UO_210 (O_210,N_23359,N_22387);
and UO_211 (O_211,N_23826,N_24773);
and UO_212 (O_212,N_23205,N_24452);
nor UO_213 (O_213,N_24332,N_21881);
and UO_214 (O_214,N_22222,N_22638);
nand UO_215 (O_215,N_23194,N_22385);
or UO_216 (O_216,N_24008,N_23391);
and UO_217 (O_217,N_24914,N_21970);
nand UO_218 (O_218,N_23873,N_22955);
nor UO_219 (O_219,N_23110,N_24977);
or UO_220 (O_220,N_22001,N_22340);
nor UO_221 (O_221,N_23161,N_23303);
and UO_222 (O_222,N_23824,N_24822);
or UO_223 (O_223,N_23481,N_23172);
or UO_224 (O_224,N_21893,N_23103);
nor UO_225 (O_225,N_24646,N_22945);
and UO_226 (O_226,N_22808,N_23796);
nor UO_227 (O_227,N_24863,N_24388);
or UO_228 (O_228,N_22677,N_22608);
or UO_229 (O_229,N_23835,N_22299);
or UO_230 (O_230,N_23435,N_24540);
nor UO_231 (O_231,N_23427,N_23278);
nand UO_232 (O_232,N_24242,N_24046);
or UO_233 (O_233,N_23260,N_23806);
nor UO_234 (O_234,N_23117,N_22235);
xor UO_235 (O_235,N_22014,N_24790);
xnor UO_236 (O_236,N_23368,N_22177);
nand UO_237 (O_237,N_22799,N_23216);
nand UO_238 (O_238,N_24208,N_23229);
and UO_239 (O_239,N_24416,N_24801);
nor UO_240 (O_240,N_22720,N_24360);
xor UO_241 (O_241,N_23863,N_24682);
nand UO_242 (O_242,N_21932,N_23440);
or UO_243 (O_243,N_22841,N_22654);
and UO_244 (O_244,N_23746,N_24083);
or UO_245 (O_245,N_22771,N_24750);
or UO_246 (O_246,N_23254,N_24932);
or UO_247 (O_247,N_23516,N_21996);
or UO_248 (O_248,N_23398,N_24314);
nand UO_249 (O_249,N_23979,N_23624);
nand UO_250 (O_250,N_22553,N_22884);
or UO_251 (O_251,N_24149,N_24847);
nor UO_252 (O_252,N_24010,N_23459);
nor UO_253 (O_253,N_23602,N_23816);
or UO_254 (O_254,N_24268,N_23163);
nand UO_255 (O_255,N_24634,N_24293);
xnor UO_256 (O_256,N_23921,N_24380);
nor UO_257 (O_257,N_22737,N_24954);
or UO_258 (O_258,N_22139,N_24560);
nor UO_259 (O_259,N_22923,N_24280);
nor UO_260 (O_260,N_24712,N_22212);
nor UO_261 (O_261,N_24002,N_21914);
nand UO_262 (O_262,N_24609,N_22452);
and UO_263 (O_263,N_24228,N_24194);
nor UO_264 (O_264,N_23638,N_22953);
nor UO_265 (O_265,N_23880,N_23095);
nand UO_266 (O_266,N_24789,N_23127);
nor UO_267 (O_267,N_22864,N_23652);
nor UO_268 (O_268,N_21889,N_22688);
and UO_269 (O_269,N_23698,N_23214);
and UO_270 (O_270,N_22079,N_24448);
nor UO_271 (O_271,N_24290,N_24343);
nor UO_272 (O_272,N_24213,N_24627);
or UO_273 (O_273,N_24215,N_22161);
xor UO_274 (O_274,N_24892,N_24019);
or UO_275 (O_275,N_22031,N_23582);
nand UO_276 (O_276,N_22217,N_24747);
nor UO_277 (O_277,N_24382,N_24684);
nand UO_278 (O_278,N_24864,N_22882);
nand UO_279 (O_279,N_21984,N_23614);
or UO_280 (O_280,N_22894,N_24088);
or UO_281 (O_281,N_24359,N_22116);
and UO_282 (O_282,N_23504,N_21901);
nand UO_283 (O_283,N_24070,N_22988);
or UO_284 (O_284,N_24044,N_23657);
nor UO_285 (O_285,N_22601,N_23251);
nor UO_286 (O_286,N_24979,N_24060);
nor UO_287 (O_287,N_22809,N_24571);
and UO_288 (O_288,N_22557,N_22272);
nor UO_289 (O_289,N_24504,N_22917);
or UO_290 (O_290,N_24432,N_23859);
and UO_291 (O_291,N_22368,N_23265);
or UO_292 (O_292,N_24231,N_22081);
and UO_293 (O_293,N_22370,N_24107);
nand UO_294 (O_294,N_22332,N_22663);
nor UO_295 (O_295,N_23780,N_23949);
nand UO_296 (O_296,N_22390,N_24947);
or UO_297 (O_297,N_22800,N_22238);
nand UO_298 (O_298,N_24668,N_21968);
nand UO_299 (O_299,N_21877,N_24862);
and UO_300 (O_300,N_23938,N_23832);
xor UO_301 (O_301,N_22653,N_21913);
and UO_302 (O_302,N_23488,N_24738);
xor UO_303 (O_303,N_23299,N_22784);
and UO_304 (O_304,N_24035,N_22743);
nor UO_305 (O_305,N_24056,N_22979);
nor UO_306 (O_306,N_24387,N_22363);
and UO_307 (O_307,N_22854,N_23182);
or UO_308 (O_308,N_23243,N_24026);
or UO_309 (O_309,N_23130,N_23895);
and UO_310 (O_310,N_22219,N_23893);
nand UO_311 (O_311,N_24576,N_23367);
nor UO_312 (O_312,N_22303,N_24256);
or UO_313 (O_313,N_23219,N_23665);
and UO_314 (O_314,N_24985,N_22264);
or UO_315 (O_315,N_23012,N_24732);
nand UO_316 (O_316,N_22660,N_24172);
xnor UO_317 (O_317,N_21938,N_23678);
nor UO_318 (O_318,N_24945,N_23410);
or UO_319 (O_319,N_23951,N_23874);
or UO_320 (O_320,N_23286,N_23577);
and UO_321 (O_321,N_24080,N_23206);
nor UO_322 (O_322,N_23053,N_23011);
or UO_323 (O_323,N_23351,N_22195);
nor UO_324 (O_324,N_22727,N_23667);
nand UO_325 (O_325,N_21954,N_23225);
nand UO_326 (O_326,N_23016,N_23976);
and UO_327 (O_327,N_23675,N_22098);
nor UO_328 (O_328,N_24933,N_24906);
nor UO_329 (O_329,N_22556,N_24214);
nor UO_330 (O_330,N_23961,N_22640);
or UO_331 (O_331,N_24096,N_22840);
nor UO_332 (O_332,N_23294,N_23943);
and UO_333 (O_333,N_24381,N_23987);
xnor UO_334 (O_334,N_22115,N_22912);
nor UO_335 (O_335,N_24846,N_23423);
and UO_336 (O_336,N_23636,N_24850);
nor UO_337 (O_337,N_23404,N_23454);
nand UO_338 (O_338,N_23779,N_22326);
nand UO_339 (O_339,N_24270,N_22517);
and UO_340 (O_340,N_22964,N_22974);
nor UO_341 (O_341,N_24065,N_24097);
and UO_342 (O_342,N_22246,N_23035);
nor UO_343 (O_343,N_24744,N_24592);
nor UO_344 (O_344,N_24480,N_24195);
or UO_345 (O_345,N_23542,N_23252);
nor UO_346 (O_346,N_23326,N_23944);
and UO_347 (O_347,N_22394,N_23385);
and UO_348 (O_348,N_23147,N_23584);
or UO_349 (O_349,N_24303,N_22772);
nand UO_350 (O_350,N_23370,N_23458);
nor UO_351 (O_351,N_23587,N_23933);
and UO_352 (O_352,N_22906,N_23608);
nor UO_353 (O_353,N_24077,N_24111);
nor UO_354 (O_354,N_22313,N_23217);
nor UO_355 (O_355,N_22659,N_23094);
nand UO_356 (O_356,N_23168,N_23664);
nand UO_357 (O_357,N_23366,N_24465);
nand UO_358 (O_358,N_22276,N_23619);
or UO_359 (O_359,N_22745,N_24261);
nand UO_360 (O_360,N_23471,N_23998);
or UO_361 (O_361,N_23099,N_24237);
nor UO_362 (O_362,N_23932,N_24205);
or UO_363 (O_363,N_24723,N_22532);
nor UO_364 (O_364,N_24437,N_24007);
and UO_365 (O_365,N_23898,N_24444);
nor UO_366 (O_366,N_23424,N_22970);
nand UO_367 (O_367,N_22392,N_23633);
and UO_368 (O_368,N_24143,N_24575);
or UO_369 (O_369,N_24645,N_23394);
and UO_370 (O_370,N_24113,N_24973);
xnor UO_371 (O_371,N_23270,N_24024);
and UO_372 (O_372,N_23994,N_22519);
nand UO_373 (O_373,N_24835,N_24074);
and UO_374 (O_374,N_24061,N_22628);
nor UO_375 (O_375,N_22484,N_22511);
and UO_376 (O_376,N_22844,N_23342);
or UO_377 (O_377,N_22571,N_24377);
nand UO_378 (O_378,N_22041,N_23646);
xnor UO_379 (O_379,N_24786,N_24460);
and UO_380 (O_380,N_23390,N_24441);
xor UO_381 (O_381,N_22992,N_21884);
nand UO_382 (O_382,N_24588,N_22209);
and UO_383 (O_383,N_24844,N_23115);
nor UO_384 (O_384,N_24788,N_23030);
and UO_385 (O_385,N_22549,N_23793);
nor UO_386 (O_386,N_23795,N_22835);
nor UO_387 (O_387,N_23809,N_22277);
nor UO_388 (O_388,N_23750,N_24400);
and UO_389 (O_389,N_24493,N_24897);
xor UO_390 (O_390,N_23112,N_24644);
xor UO_391 (O_391,N_24654,N_23197);
or UO_392 (O_392,N_22521,N_23829);
and UO_393 (O_393,N_22086,N_24680);
and UO_394 (O_394,N_24503,N_23869);
nand UO_395 (O_395,N_24285,N_22164);
nor UO_396 (O_396,N_22837,N_23397);
or UO_397 (O_397,N_24494,N_23354);
or UO_398 (O_398,N_24392,N_24102);
nor UO_399 (O_399,N_23451,N_24475);
nand UO_400 (O_400,N_22971,N_24287);
nor UO_401 (O_401,N_24294,N_22916);
nand UO_402 (O_402,N_22621,N_23295);
or UO_403 (O_403,N_24866,N_22562);
or UO_404 (O_404,N_24442,N_24601);
or UO_405 (O_405,N_22528,N_23919);
nor UO_406 (O_406,N_24058,N_23009);
and UO_407 (O_407,N_22275,N_22588);
xor UO_408 (O_408,N_24227,N_22627);
nor UO_409 (O_409,N_24885,N_22490);
or UO_410 (O_410,N_22694,N_22749);
xnor UO_411 (O_411,N_22523,N_24150);
and UO_412 (O_412,N_24968,N_23965);
or UO_413 (O_413,N_22443,N_22637);
or UO_414 (O_414,N_22347,N_22967);
or UO_415 (O_415,N_24676,N_22172);
or UO_416 (O_416,N_22704,N_22855);
or UO_417 (O_417,N_22903,N_24146);
nor UO_418 (O_418,N_24185,N_22119);
nand UO_419 (O_419,N_22789,N_23971);
nand UO_420 (O_420,N_22165,N_23259);
nor UO_421 (O_421,N_22895,N_24707);
or UO_422 (O_422,N_24273,N_23126);
xor UO_423 (O_423,N_24856,N_24495);
and UO_424 (O_424,N_24838,N_22351);
or UO_425 (O_425,N_22260,N_23589);
and UO_426 (O_426,N_24408,N_23770);
or UO_427 (O_427,N_24905,N_22058);
and UO_428 (O_428,N_23381,N_23617);
nor UO_429 (O_429,N_23570,N_24803);
or UO_430 (O_430,N_23039,N_21962);
or UO_431 (O_431,N_23606,N_24254);
nor UO_432 (O_432,N_23524,N_24089);
nand UO_433 (O_433,N_22020,N_24986);
or UO_434 (O_434,N_23574,N_24716);
nand UO_435 (O_435,N_24124,N_22575);
and UO_436 (O_436,N_22938,N_24551);
and UO_437 (O_437,N_22846,N_24565);
or UO_438 (O_438,N_21933,N_23282);
nand UO_439 (O_439,N_23755,N_22462);
and UO_440 (O_440,N_24265,N_24030);
and UO_441 (O_441,N_23709,N_24942);
and UO_442 (O_442,N_24923,N_23555);
or UO_443 (O_443,N_24148,N_24583);
or UO_444 (O_444,N_23121,N_23659);
nand UO_445 (O_445,N_23042,N_22008);
nor UO_446 (O_446,N_22134,N_23289);
nor UO_447 (O_447,N_22649,N_21898);
or UO_448 (O_448,N_22769,N_22869);
or UO_449 (O_449,N_22990,N_23374);
or UO_450 (O_450,N_23484,N_23773);
nand UO_451 (O_451,N_22652,N_24235);
or UO_452 (O_452,N_22770,N_23529);
and UO_453 (O_453,N_24597,N_22642);
nor UO_454 (O_454,N_24715,N_22176);
nand UO_455 (O_455,N_24316,N_24243);
or UO_456 (O_456,N_22962,N_21955);
and UO_457 (O_457,N_24292,N_24915);
or UO_458 (O_458,N_23757,N_23552);
or UO_459 (O_459,N_22088,N_23615);
nand UO_460 (O_460,N_23375,N_23569);
nand UO_461 (O_461,N_24223,N_24286);
nand UO_462 (O_462,N_23854,N_23651);
and UO_463 (O_463,N_22513,N_24741);
nand UO_464 (O_464,N_24980,N_22695);
nand UO_465 (O_465,N_23406,N_22858);
xor UO_466 (O_466,N_23911,N_22215);
nor UO_467 (O_467,N_24375,N_23362);
nor UO_468 (O_468,N_22282,N_21953);
nand UO_469 (O_469,N_24943,N_23910);
nand UO_470 (O_470,N_22261,N_24283);
or UO_471 (O_471,N_22325,N_24927);
nor UO_472 (O_472,N_22428,N_22483);
or UO_473 (O_473,N_24166,N_23464);
nand UO_474 (O_474,N_22237,N_24536);
xnor UO_475 (O_475,N_22090,N_24031);
nand UO_476 (O_476,N_23597,N_23974);
nor UO_477 (O_477,N_24397,N_24826);
and UO_478 (O_478,N_23437,N_23500);
or UO_479 (O_479,N_22985,N_24649);
or UO_480 (O_480,N_22091,N_23771);
xnor UO_481 (O_481,N_22503,N_23877);
and UO_482 (O_482,N_23450,N_22009);
or UO_483 (O_483,N_23553,N_22722);
or UO_484 (O_484,N_22459,N_22850);
and UO_485 (O_485,N_24554,N_24502);
or UO_486 (O_486,N_24371,N_22900);
and UO_487 (O_487,N_22147,N_21948);
nor UO_488 (O_488,N_24804,N_24659);
nor UO_489 (O_489,N_24361,N_24546);
or UO_490 (O_490,N_23331,N_23108);
nor UO_491 (O_491,N_24244,N_23575);
nor UO_492 (O_492,N_23493,N_24912);
or UO_493 (O_493,N_22456,N_21879);
and UO_494 (O_494,N_23507,N_24084);
or UO_495 (O_495,N_23729,N_23226);
nor UO_496 (O_496,N_22812,N_24757);
and UO_497 (O_497,N_22092,N_23748);
or UO_498 (O_498,N_23520,N_23672);
or UO_499 (O_499,N_23645,N_22450);
nor UO_500 (O_500,N_22201,N_24241);
nand UO_501 (O_501,N_23157,N_23329);
nor UO_502 (O_502,N_23761,N_21966);
nand UO_503 (O_503,N_24042,N_24643);
and UO_504 (O_504,N_24313,N_22470);
xor UO_505 (O_505,N_23983,N_24764);
or UO_506 (O_506,N_24550,N_21892);
xnor UO_507 (O_507,N_23514,N_24855);
nand UO_508 (O_508,N_23563,N_22302);
or UO_509 (O_509,N_22391,N_24989);
xor UO_510 (O_510,N_24673,N_24935);
and UO_511 (O_511,N_22248,N_22508);
and UO_512 (O_512,N_23187,N_24086);
xor UO_513 (O_513,N_22300,N_24013);
and UO_514 (O_514,N_22181,N_23899);
or UO_515 (O_515,N_23133,N_23947);
nand UO_516 (O_516,N_23443,N_24165);
or UO_517 (O_517,N_23878,N_24473);
nor UO_518 (O_518,N_23113,N_24177);
xnor UO_519 (O_519,N_22744,N_23521);
and UO_520 (O_520,N_23167,N_23862);
and UO_521 (O_521,N_24131,N_23906);
or UO_522 (O_522,N_23373,N_23154);
or UO_523 (O_523,N_23071,N_22263);
nor UO_524 (O_524,N_24881,N_23777);
nor UO_525 (O_525,N_23699,N_21975);
or UO_526 (O_526,N_22613,N_23218);
nand UO_527 (O_527,N_22421,N_23063);
and UO_528 (O_528,N_22414,N_24946);
xnor UO_529 (O_529,N_24798,N_22752);
nand UO_530 (O_530,N_21973,N_21896);
nand UO_531 (O_531,N_22499,N_23323);
or UO_532 (O_532,N_23630,N_23688);
and UO_533 (O_533,N_21977,N_24559);
nand UO_534 (O_534,N_21979,N_22397);
nand UO_535 (O_535,N_24040,N_24266);
nor UO_536 (O_536,N_24574,N_22786);
nor UO_537 (O_537,N_22689,N_24167);
xnor UO_538 (O_538,N_23988,N_23230);
nand UO_539 (O_539,N_24647,N_22671);
nor UO_540 (O_540,N_22582,N_22611);
nand UO_541 (O_541,N_23057,N_23731);
nor UO_542 (O_542,N_23361,N_23211);
nand UO_543 (O_543,N_23676,N_23312);
nor UO_544 (O_544,N_22298,N_24689);
nor UO_545 (O_545,N_24319,N_23752);
nand UO_546 (O_546,N_22631,N_23647);
nor UO_547 (O_547,N_22535,N_23124);
or UO_548 (O_548,N_23003,N_23146);
or UO_549 (O_549,N_24347,N_24776);
and UO_550 (O_550,N_23872,N_22889);
xnor UO_551 (O_551,N_24721,N_23642);
xor UO_552 (O_552,N_24880,N_23122);
nand UO_553 (O_553,N_24390,N_22386);
xnor UO_554 (O_554,N_24211,N_23819);
nand UO_555 (O_555,N_23143,N_24795);
and UO_556 (O_556,N_23635,N_22909);
and UO_557 (O_557,N_22329,N_23052);
xnor UO_558 (O_558,N_24669,N_24735);
nand UO_559 (O_559,N_22740,N_23894);
xnor UO_560 (O_560,N_24763,N_23957);
or UO_561 (O_561,N_23245,N_22614);
and UO_562 (O_562,N_23046,N_24514);
nand UO_563 (O_563,N_23291,N_24806);
nand UO_564 (O_564,N_24824,N_24398);
and UO_565 (O_565,N_24053,N_24204);
nor UO_566 (O_566,N_22651,N_23421);
nand UO_567 (O_567,N_23220,N_24697);
nor UO_568 (O_568,N_23482,N_22266);
xor UO_569 (O_569,N_22965,N_23707);
and UO_570 (O_570,N_23685,N_22920);
or UO_571 (O_571,N_23153,N_23156);
or UO_572 (O_572,N_23930,N_22597);
nor UO_573 (O_573,N_23865,N_22952);
or UO_574 (O_574,N_22083,N_23904);
nand UO_575 (O_575,N_23928,N_23991);
and UO_576 (O_576,N_24636,N_24499);
and UO_577 (O_577,N_24055,N_24105);
or UO_578 (O_578,N_22596,N_23812);
nor UO_579 (O_579,N_23677,N_21997);
and UO_580 (O_580,N_24889,N_23072);
nand UO_581 (O_581,N_23141,N_23517);
xor UO_582 (O_582,N_22759,N_22551);
and UO_583 (O_583,N_22702,N_21969);
nand UO_584 (O_584,N_24274,N_22057);
nand UO_585 (O_585,N_22791,N_23223);
and UO_586 (O_586,N_23544,N_23720);
nand UO_587 (O_587,N_23333,N_23766);
and UO_588 (O_588,N_22586,N_23798);
or UO_589 (O_589,N_24663,N_24894);
xnor UO_590 (O_590,N_24957,N_23628);
or UO_591 (O_591,N_22021,N_24229);
nand UO_592 (O_592,N_24489,N_23581);
and UO_593 (O_593,N_22875,N_24521);
nand UO_594 (O_594,N_21958,N_23839);
nand UO_595 (O_595,N_22986,N_23149);
nand UO_596 (O_596,N_23319,N_23954);
nor UO_597 (O_597,N_22336,N_24027);
nor UO_598 (O_598,N_23886,N_22773);
or UO_599 (O_599,N_24034,N_22190);
xor UO_600 (O_600,N_23722,N_22382);
nand UO_601 (O_601,N_24501,N_23683);
nand UO_602 (O_602,N_22991,N_22220);
nand UO_603 (O_603,N_22454,N_24159);
or UO_604 (O_604,N_22297,N_23753);
nor UO_605 (O_605,N_24520,N_21924);
xor UO_606 (O_606,N_22295,N_23853);
xnor UO_607 (O_607,N_24525,N_24834);
nand UO_608 (O_608,N_22552,N_24253);
nor UO_609 (O_609,N_22244,N_24157);
nor UO_610 (O_610,N_24186,N_23340);
xnor UO_611 (O_611,N_21882,N_24568);
and UO_612 (O_612,N_23392,N_22448);
and UO_613 (O_613,N_22384,N_23080);
and UO_614 (O_614,N_23005,N_22978);
nor UO_615 (O_615,N_24796,N_22493);
nand UO_616 (O_616,N_22818,N_24079);
nand UO_617 (O_617,N_24538,N_24192);
nor UO_618 (O_618,N_22968,N_24518);
or UO_619 (O_619,N_22851,N_24155);
or UO_620 (O_620,N_23595,N_24637);
and UO_621 (O_621,N_22573,N_23820);
and UO_622 (O_622,N_22427,N_23639);
xnor UO_623 (O_623,N_24217,N_22533);
nor UO_624 (O_624,N_24828,N_23879);
and UO_625 (O_625,N_22097,N_21982);
or UO_626 (O_626,N_23915,N_22650);
xnor UO_627 (O_627,N_24865,N_24940);
or UO_628 (O_628,N_24825,N_22871);
nand UO_629 (O_629,N_22269,N_23913);
and UO_630 (O_630,N_24991,N_24385);
nand UO_631 (O_631,N_24093,N_23396);
nand UO_632 (O_632,N_22491,N_24861);
nand UO_633 (O_633,N_23179,N_24043);
nand UO_634 (O_634,N_23283,N_23559);
or UO_635 (O_635,N_24188,N_22830);
nor UO_636 (O_636,N_23528,N_23592);
nor UO_637 (O_637,N_24807,N_22543);
nor UO_638 (O_638,N_22566,N_24569);
or UO_639 (O_639,N_22699,N_23369);
and UO_640 (O_640,N_24809,N_22580);
and UO_641 (O_641,N_23613,N_24820);
or UO_642 (O_642,N_24170,N_24662);
and UO_643 (O_643,N_22205,N_23448);
nand UO_644 (O_644,N_24367,N_24958);
and UO_645 (O_645,N_22192,N_24001);
nand UO_646 (O_646,N_24317,N_22078);
or UO_647 (O_647,N_24199,N_22766);
and UO_648 (O_648,N_22228,N_23185);
nor UO_649 (O_649,N_24118,N_23271);
xnor UO_650 (O_650,N_22128,N_24032);
nand UO_651 (O_651,N_23334,N_24875);
nand UO_652 (O_652,N_24370,N_23706);
nor UO_653 (O_653,N_24547,N_24104);
nor UO_654 (O_654,N_24249,N_24068);
nand UO_655 (O_655,N_23674,N_23357);
or UO_656 (O_656,N_23840,N_24189);
or UO_657 (O_657,N_24903,N_22230);
nand UO_658 (O_658,N_23281,N_24900);
or UO_659 (O_659,N_22018,N_24289);
nor UO_660 (O_660,N_22960,N_23040);
xor UO_661 (O_661,N_22507,N_21952);
or UO_662 (O_662,N_22746,N_22357);
xnor UO_663 (O_663,N_24033,N_23660);
nand UO_664 (O_664,N_22885,N_23316);
or UO_665 (O_665,N_22589,N_22918);
xor UO_666 (O_666,N_24063,N_24607);
nor UO_667 (O_667,N_23781,N_24054);
or UO_668 (O_668,N_22180,N_24777);
nand UO_669 (O_669,N_24877,N_24528);
or UO_670 (O_670,N_22257,N_24471);
and UO_671 (O_671,N_23134,N_22646);
nor UO_672 (O_672,N_22498,N_24421);
or UO_673 (O_673,N_21985,N_24742);
xnor UO_674 (O_674,N_22526,N_24216);
nor UO_675 (O_675,N_22207,N_23543);
or UO_676 (O_676,N_23601,N_21878);
or UO_677 (O_677,N_22066,N_21974);
or UO_678 (O_678,N_24036,N_23138);
nand UO_679 (O_679,N_22856,N_22795);
nand UO_680 (O_680,N_24591,N_21959);
nor UO_681 (O_681,N_23114,N_23327);
and UO_682 (O_682,N_22461,N_23567);
or UO_683 (O_683,N_22210,N_23338);
and UO_684 (O_684,N_22204,N_23430);
nor UO_685 (O_685,N_23629,N_22914);
nor UO_686 (O_686,N_23083,N_22250);
nand UO_687 (O_687,N_22240,N_22405);
or UO_688 (O_688,N_23304,N_23803);
and UO_689 (O_689,N_23515,N_23942);
and UO_690 (O_690,N_24057,N_24041);
nand UO_691 (O_691,N_24555,N_23922);
nand UO_692 (O_692,N_24472,N_23579);
nand UO_693 (O_693,N_22813,N_24685);
and UO_694 (O_694,N_22630,N_23980);
xor UO_695 (O_695,N_23360,N_22880);
or UO_696 (O_696,N_24507,N_24896);
nand UO_697 (O_697,N_23549,N_23018);
nand UO_698 (O_698,N_23782,N_24690);
and UO_699 (O_699,N_22534,N_24466);
and UO_700 (O_700,N_22687,N_23769);
nor UO_701 (O_701,N_23461,N_24248);
and UO_702 (O_702,N_23843,N_23875);
or UO_703 (O_703,N_23737,N_22350);
xnor UO_704 (O_704,N_24882,N_24848);
nor UO_705 (O_705,N_22043,N_24655);
or UO_706 (O_706,N_22669,N_24218);
xnor UO_707 (O_707,N_24171,N_23775);
or UO_708 (O_708,N_24755,N_23330);
nor UO_709 (O_709,N_23572,N_23344);
and UO_710 (O_710,N_22886,N_22112);
xnor UO_711 (O_711,N_24039,N_24871);
nor UO_712 (O_712,N_23152,N_24966);
xor UO_713 (O_713,N_23513,N_23815);
or UO_714 (O_714,N_22691,N_22656);
or UO_715 (O_715,N_22155,N_22442);
and UO_716 (O_716,N_23656,N_22681);
nand UO_717 (O_717,N_23348,N_21943);
xnor UO_718 (O_718,N_24403,N_23007);
and UO_719 (O_719,N_24011,N_22038);
nand UO_720 (O_720,N_22283,N_23277);
or UO_721 (O_721,N_24071,N_24561);
nand UO_722 (O_722,N_23210,N_22289);
and UO_723 (O_723,N_22281,N_22106);
nor UO_724 (O_724,N_22311,N_23475);
or UO_725 (O_725,N_24926,N_21947);
nand UO_726 (O_726,N_24629,N_22788);
nor UO_727 (O_727,N_23681,N_23492);
and UO_728 (O_728,N_23765,N_23641);
and UO_729 (O_729,N_22584,N_24378);
nor UO_730 (O_730,N_22223,N_22756);
and UO_731 (O_731,N_24904,N_24913);
nand UO_732 (O_732,N_22943,N_24014);
or UO_733 (O_733,N_24959,N_23159);
nand UO_734 (O_734,N_22379,N_22131);
nand UO_735 (O_735,N_24717,N_24758);
and UO_736 (O_736,N_23002,N_23028);
nand UO_737 (O_737,N_23184,N_22989);
and UO_738 (O_738,N_22017,N_23655);
or UO_739 (O_739,N_23062,N_24511);
or UO_740 (O_740,N_23786,N_23714);
and UO_741 (O_741,N_23276,N_22976);
nor UO_742 (O_742,N_22328,N_24457);
xnor UO_743 (O_743,N_24727,N_22199);
and UO_744 (O_744,N_23925,N_24406);
nor UO_745 (O_745,N_23140,N_21907);
nand UO_746 (O_746,N_24486,N_21918);
or UO_747 (O_747,N_23325,N_24693);
and UO_748 (O_748,N_24134,N_22065);
nand UO_749 (O_749,N_23297,N_22129);
and UO_750 (O_750,N_23241,N_24258);
or UO_751 (O_751,N_24817,N_23596);
and UO_752 (O_752,N_24529,N_23934);
nand UO_753 (O_753,N_23409,N_22348);
and UO_754 (O_754,N_23591,N_22093);
or UO_755 (O_755,N_21880,N_22323);
nor UO_756 (O_756,N_21919,N_23195);
and UO_757 (O_757,N_24614,N_24373);
and UO_758 (O_758,N_24278,N_23997);
nor UO_759 (O_759,N_22015,N_24572);
nand UO_760 (O_760,N_23466,N_23959);
and UO_761 (O_761,N_23648,N_24103);
or UO_762 (O_762,N_23789,N_22120);
or UO_763 (O_763,N_22292,N_23322);
xor UO_764 (O_764,N_23996,N_24048);
nor UO_765 (O_765,N_21920,N_22460);
and UO_766 (O_766,N_24496,N_24478);
nor UO_767 (O_767,N_23181,N_23856);
or UO_768 (O_768,N_23759,N_23300);
nor UO_769 (O_769,N_22194,N_23849);
nor UO_770 (O_770,N_24020,N_23213);
and UO_771 (O_771,N_22554,N_23238);
xnor UO_772 (O_772,N_22542,N_22942);
nor UO_773 (O_773,N_22055,N_24544);
and UO_774 (O_774,N_22337,N_22407);
nand UO_775 (O_775,N_22371,N_24638);
xnor UO_776 (O_776,N_24396,N_22763);
nor UO_777 (O_777,N_23209,N_22327);
nor UO_778 (O_778,N_23097,N_22954);
or UO_779 (O_779,N_22265,N_23311);
or UO_780 (O_780,N_24414,N_23058);
or UO_781 (O_781,N_24296,N_24766);
and UO_782 (O_782,N_22996,N_23525);
xor UO_783 (O_783,N_24409,N_23240);
nor UO_784 (O_784,N_24418,N_24508);
or UO_785 (O_785,N_22108,N_24288);
nor UO_786 (O_786,N_24431,N_22469);
nand UO_787 (O_787,N_23452,N_22583);
nand UO_788 (O_788,N_23790,N_24429);
nor UO_789 (O_789,N_24687,N_22934);
nand UO_790 (O_790,N_22089,N_22023);
and UO_791 (O_791,N_22130,N_24600);
or UO_792 (O_792,N_24672,N_23096);
and UO_793 (O_793,N_24995,N_24012);
nand UO_794 (O_794,N_22288,N_23164);
and UO_795 (O_795,N_24901,N_23710);
and UO_796 (O_796,N_24652,N_24481);
nand UO_797 (O_797,N_22389,N_22451);
nand UO_798 (O_798,N_22305,N_23070);
or UO_799 (O_799,N_24300,N_22940);
nand UO_800 (O_800,N_22247,N_24941);
nor UO_801 (O_801,N_23033,N_22890);
xor UO_802 (O_802,N_23477,N_24299);
or UO_803 (O_803,N_24309,N_24468);
nor UO_804 (O_804,N_21971,N_22930);
and UO_805 (O_805,N_24407,N_24028);
nor UO_806 (O_806,N_22019,N_24327);
nand UO_807 (O_807,N_21894,N_22783);
nand UO_808 (O_808,N_22358,N_22868);
and UO_809 (O_809,N_22734,N_22861);
or UO_810 (O_810,N_22434,N_23017);
and UO_811 (O_811,N_23449,N_22975);
nor UO_812 (O_812,N_22785,N_23337);
nor UO_813 (O_813,N_23176,N_22150);
nand UO_814 (O_814,N_24883,N_22479);
nor UO_815 (O_815,N_22548,N_24389);
and UO_816 (O_816,N_23627,N_22665);
nor UO_817 (O_817,N_24944,N_23643);
xor UO_818 (O_818,N_22304,N_22524);
and UO_819 (O_819,N_22286,N_22438);
xnor UO_820 (O_820,N_23964,N_24664);
or UO_821 (O_821,N_23536,N_24515);
nand UO_822 (O_822,N_23479,N_24363);
nand UO_823 (O_823,N_22042,N_24500);
and UO_824 (O_824,N_22603,N_23347);
nand UO_825 (O_825,N_22362,N_22411);
xor UO_826 (O_826,N_24840,N_23125);
or UO_827 (O_827,N_23273,N_21876);
nor UO_828 (O_828,N_24842,N_22050);
or UO_829 (O_829,N_24761,N_22403);
nand UO_830 (O_830,N_24867,N_24651);
and UO_831 (O_831,N_23799,N_23669);
nand UO_832 (O_832,N_23855,N_24729);
nand UO_833 (O_833,N_24395,N_23049);
and UO_834 (O_834,N_24939,N_23456);
xor UO_835 (O_835,N_22594,N_23177);
nand UO_836 (O_836,N_22142,N_22728);
nand UO_837 (O_837,N_23224,N_24321);
or UO_838 (O_838,N_23650,N_22805);
nand UO_839 (O_839,N_22820,N_24355);
and UO_840 (O_840,N_23701,N_23339);
or UO_841 (O_841,N_24066,N_22958);
xnor UO_842 (O_842,N_23668,N_24420);
or UO_843 (O_843,N_22576,N_23417);
or UO_844 (O_844,N_23136,N_23442);
and UO_845 (O_845,N_24006,N_23952);
nor UO_846 (O_846,N_24474,N_22429);
and UO_847 (O_847,N_22214,N_22290);
nand UO_848 (O_848,N_23349,N_22133);
nand UO_849 (O_849,N_23302,N_22258);
or UO_850 (O_850,N_22565,N_23151);
nor UO_851 (O_851,N_24318,N_24003);
nand UO_852 (O_852,N_22619,N_22635);
and UO_853 (O_853,N_23993,N_23384);
nand UO_854 (O_854,N_24666,N_24073);
nor UO_855 (O_855,N_24916,N_24990);
nand UO_856 (O_856,N_24930,N_23745);
and UO_857 (O_857,N_23741,N_24233);
and UO_858 (O_858,N_23173,N_23001);
and UO_859 (O_859,N_23228,N_22076);
or UO_860 (O_860,N_22040,N_23499);
nor UO_861 (O_861,N_24391,N_22711);
and UO_862 (O_862,N_22946,N_24924);
nand UO_863 (O_863,N_23268,N_23480);
and UO_864 (O_864,N_22312,N_24818);
or UO_865 (O_865,N_23174,N_22136);
nand UO_866 (O_866,N_24141,N_21906);
and UO_867 (O_867,N_22595,N_23963);
nor UO_868 (O_868,N_24281,N_24671);
nand UO_869 (O_869,N_24004,N_22824);
xnor UO_870 (O_870,N_23335,N_22399);
nor UO_871 (O_871,N_24338,N_23196);
nand UO_872 (O_872,N_24632,N_22873);
xor UO_873 (O_873,N_21983,N_24449);
nand UO_874 (O_874,N_23119,N_24698);
xor UO_875 (O_875,N_24626,N_23264);
and UO_876 (O_876,N_23772,N_23604);
or UO_877 (O_877,N_23422,N_22028);
and UO_878 (O_878,N_23445,N_23034);
and UO_879 (O_879,N_23754,N_24247);
or UO_880 (O_880,N_24686,N_24470);
or UO_881 (O_881,N_23465,N_22959);
xor UO_882 (O_882,N_24759,N_21917);
nand UO_883 (O_883,N_22832,N_23026);
nor UO_884 (O_884,N_22135,N_24812);
nor UO_885 (O_885,N_21992,N_23503);
nand UO_886 (O_886,N_24934,N_23813);
nand UO_887 (O_887,N_23532,N_22198);
nand UO_888 (O_888,N_23455,N_24767);
and UO_889 (O_889,N_23900,N_23876);
or UO_890 (O_890,N_23931,N_24425);
or UO_891 (O_891,N_23089,N_22060);
nor UO_892 (O_892,N_24642,N_24410);
and UO_893 (O_893,N_24353,N_22559);
xor UO_894 (O_894,N_22231,N_22622);
or UO_895 (O_895,N_24641,N_22550);
or UO_896 (O_896,N_22944,N_22342);
nor UO_897 (O_897,N_22599,N_23460);
nor UO_898 (O_898,N_23692,N_22431);
or UO_899 (O_899,N_22229,N_24650);
nor UO_900 (O_900,N_24312,N_23321);
or UO_901 (O_901,N_23747,N_22182);
nor UO_902 (O_902,N_22819,N_24025);
or UO_903 (O_903,N_21936,N_23429);
and UO_904 (O_904,N_21967,N_23927);
and UO_905 (O_905,N_24993,N_24836);
nand UO_906 (O_906,N_23019,N_24130);
nor UO_907 (O_907,N_24615,N_23434);
and UO_908 (O_908,N_22568,N_23690);
nor UO_909 (O_909,N_22564,N_24537);
xor UO_910 (O_910,N_24417,N_22373);
nor UO_911 (O_911,N_22879,N_22123);
xnor UO_912 (O_912,N_23857,N_21885);
and UO_913 (O_913,N_23866,N_23621);
or UO_914 (O_914,N_22941,N_23345);
or UO_915 (O_915,N_22685,N_22712);
and UO_916 (O_916,N_22101,N_24631);
nor UO_917 (O_917,N_22569,N_24888);
or UO_918 (O_918,N_22883,N_22143);
nor UO_919 (O_919,N_24988,N_23020);
or UO_920 (O_920,N_22902,N_24611);
xnor UO_921 (O_921,N_22032,N_22848);
nand UO_922 (O_922,N_23065,N_22765);
xor UO_923 (O_923,N_24931,N_22705);
or UO_924 (O_924,N_24219,N_22171);
xor UO_925 (O_925,N_23905,N_23607);
or UO_926 (O_926,N_23721,N_23519);
xor UO_927 (O_927,N_23888,N_23137);
and UO_928 (O_928,N_24260,N_23742);
nand UO_929 (O_929,N_24596,N_22878);
nand UO_930 (O_930,N_22396,N_22162);
xor UO_931 (O_931,N_22693,N_23618);
nor UO_932 (O_932,N_24760,N_23726);
nand UO_933 (O_933,N_22951,N_23848);
or UO_934 (O_934,N_22639,N_23082);
or UO_935 (O_935,N_24257,N_22672);
or UO_936 (O_936,N_23887,N_24152);
and UO_937 (O_937,N_24116,N_22270);
nand UO_938 (O_938,N_23560,N_22464);
nand UO_939 (O_939,N_24779,N_24740);
nand UO_940 (O_940,N_23100,N_22322);
nand UO_941 (O_941,N_24451,N_22433);
and UO_942 (O_942,N_23661,N_24350);
nand UO_943 (O_943,N_24369,N_22686);
xor UO_944 (O_944,N_23852,N_22356);
nor UO_945 (O_945,N_24782,N_22208);
and UO_946 (O_946,N_24787,N_22146);
or UO_947 (O_947,N_22527,N_22838);
nand UO_948 (O_948,N_23263,N_21940);
and UO_949 (O_949,N_22318,N_23008);
nand UO_950 (O_950,N_22777,N_24743);
and UO_951 (O_951,N_23565,N_23912);
and UO_952 (O_952,N_23836,N_24677);
nand UO_953 (O_953,N_24308,N_22792);
nor UO_954 (O_954,N_24628,N_24580);
nor UO_955 (O_955,N_24884,N_24112);
nand UO_956 (O_956,N_22683,N_22067);
or UO_957 (O_957,N_24232,N_24037);
or UO_958 (O_958,N_22273,N_22402);
nand UO_959 (O_959,N_24553,N_23837);
or UO_960 (O_960,N_23736,N_22420);
xor UO_961 (O_961,N_23794,N_24252);
nand UO_962 (O_962,N_22388,N_24509);
or UO_963 (O_963,N_24691,N_23415);
nand UO_964 (O_964,N_23972,N_22540);
or UO_965 (O_965,N_24635,N_21909);
or UO_966 (O_966,N_23956,N_24519);
nand UO_967 (O_967,N_24200,N_23735);
xnor UO_968 (O_968,N_23496,N_22796);
nor UO_969 (O_969,N_22061,N_23823);
nor UO_970 (O_970,N_24181,N_23576);
nand UO_971 (O_971,N_22617,N_22094);
or UO_972 (O_972,N_22335,N_22280);
nor UO_973 (O_973,N_23116,N_24908);
nand UO_974 (O_974,N_22148,N_22966);
xor UO_975 (O_975,N_24366,N_22790);
xnor UO_976 (O_976,N_23700,N_23077);
xor UO_977 (O_977,N_22703,N_23469);
or UO_978 (O_978,N_24535,N_24603);
nand UO_979 (O_979,N_23955,N_22213);
and UO_980 (O_980,N_24187,N_23787);
and UO_981 (O_981,N_23724,N_23215);
nand UO_982 (O_982,N_23165,N_22842);
and UO_983 (O_983,N_22767,N_24710);
and UO_984 (O_984,N_22913,N_22439);
and UO_985 (O_985,N_24830,N_23540);
nand UO_986 (O_986,N_23236,N_22932);
xor UO_987 (O_987,N_22376,N_24953);
nand UO_988 (O_988,N_24772,N_23756);
and UO_989 (O_989,N_24983,N_24874);
nand UO_990 (O_990,N_22425,N_22338);
or UO_991 (O_991,N_24562,N_24487);
or UO_992 (O_992,N_23834,N_24333);
and UO_993 (O_993,N_23708,N_21931);
or UO_994 (O_994,N_24678,N_24955);
nor UO_995 (O_995,N_22698,N_24981);
or UO_996 (O_996,N_23457,N_23494);
xor UO_997 (O_997,N_22680,N_22852);
nor UO_998 (O_998,N_22561,N_24595);
nand UO_999 (O_999,N_22441,N_23962);
xor UO_1000 (O_1000,N_23111,N_24907);
xnor UO_1001 (O_1001,N_24009,N_23352);
or UO_1002 (O_1002,N_23188,N_24210);
or UO_1003 (O_1003,N_22051,N_23064);
and UO_1004 (O_1004,N_24049,N_23881);
nand UO_1005 (O_1005,N_24302,N_22249);
nor UO_1006 (O_1006,N_21990,N_24064);
nor UO_1007 (O_1007,N_22424,N_22817);
or UO_1008 (O_1008,N_22126,N_23632);
and UO_1009 (O_1009,N_23419,N_23242);
nand UO_1010 (O_1010,N_22095,N_23918);
and UO_1011 (O_1011,N_24910,N_23599);
or UO_1012 (O_1012,N_23920,N_23716);
nand UO_1013 (O_1013,N_22037,N_24810);
or UO_1014 (O_1014,N_22781,N_24704);
and UO_1015 (O_1015,N_23844,N_24833);
nand UO_1016 (O_1016,N_24573,N_24142);
nand UO_1017 (O_1017,N_23084,N_23232);
and UO_1018 (O_1018,N_23372,N_22915);
or UO_1019 (O_1019,N_22005,N_24506);
xnor UO_1020 (O_1020,N_24909,N_23076);
nor UO_1021 (O_1021,N_24695,N_22537);
nand UO_1022 (O_1022,N_24419,N_23284);
nand UO_1023 (O_1023,N_23145,N_22369);
nand UO_1024 (O_1024,N_23749,N_22600);
nor UO_1025 (O_1025,N_23418,N_23966);
xor UO_1026 (O_1026,N_24701,N_23696);
and UO_1027 (O_1027,N_23400,N_24582);
nand UO_1028 (O_1028,N_23622,N_22398);
and UO_1029 (O_1029,N_24469,N_22084);
nor UO_1030 (O_1030,N_21927,N_23092);
nand UO_1031 (O_1031,N_23262,N_23838);
xor UO_1032 (O_1032,N_24522,N_24921);
or UO_1033 (O_1033,N_23889,N_22410);
nand UO_1034 (O_1034,N_21916,N_24276);
nor UO_1035 (O_1035,N_22036,N_22950);
nand UO_1036 (O_1036,N_23066,N_24492);
and UO_1037 (O_1037,N_22487,N_22064);
or UO_1038 (O_1038,N_23892,N_22657);
and UO_1039 (O_1039,N_21925,N_22062);
nand UO_1040 (O_1040,N_24622,N_23871);
and UO_1041 (O_1041,N_22696,N_24222);
nor UO_1042 (O_1042,N_24151,N_24975);
or UO_1043 (O_1043,N_24099,N_22000);
nor UO_1044 (O_1044,N_21998,N_23550);
or UO_1045 (O_1045,N_22476,N_23945);
nor UO_1046 (O_1046,N_24119,N_22104);
or UO_1047 (O_1047,N_23649,N_24436);
nor UO_1048 (O_1048,N_22570,N_23074);
or UO_1049 (O_1049,N_23686,N_23817);
or UO_1050 (O_1050,N_24005,N_24362);
and UO_1051 (O_1051,N_23858,N_24246);
or UO_1052 (O_1052,N_21942,N_22200);
xnor UO_1053 (O_1053,N_22623,N_24567);
nor UO_1054 (O_1054,N_22107,N_22972);
nor UO_1055 (O_1055,N_23860,N_22983);
and UO_1056 (O_1056,N_24784,N_22359);
nor UO_1057 (O_1057,N_24335,N_23509);
nand UO_1058 (O_1058,N_24532,N_23102);
nand UO_1059 (O_1059,N_24517,N_24110);
nand UO_1060 (O_1060,N_22154,N_23044);
nor UO_1061 (O_1061,N_23940,N_22998);
nor UO_1062 (O_1062,N_24344,N_23006);
and UO_1063 (O_1063,N_22211,N_23916);
or UO_1064 (O_1064,N_24658,N_23833);
nand UO_1065 (O_1065,N_22969,N_24545);
or UO_1066 (O_1066,N_23530,N_22748);
or UO_1067 (O_1067,N_24987,N_24621);
nor UO_1068 (O_1068,N_24198,N_22105);
or UO_1069 (O_1069,N_22936,N_23758);
or UO_1070 (O_1070,N_22477,N_23498);
or UO_1071 (O_1071,N_23387,N_22113);
or UO_1072 (O_1072,N_21946,N_24476);
or UO_1073 (O_1073,N_24510,N_21987);
nor UO_1074 (O_1074,N_23267,N_22052);
nand UO_1075 (O_1075,N_22339,N_23718);
and UO_1076 (O_1076,N_24878,N_23439);
and UO_1077 (O_1077,N_23013,N_22697);
nor UO_1078 (O_1078,N_24996,N_23431);
nor UO_1079 (O_1079,N_22241,N_22485);
nor UO_1080 (O_1080,N_24029,N_24837);
and UO_1081 (O_1081,N_23929,N_24952);
nand UO_1082 (O_1082,N_23239,N_21980);
nand UO_1083 (O_1083,N_22605,N_24793);
nand UO_1084 (O_1084,N_24950,N_23827);
nand UO_1085 (O_1085,N_22378,N_21905);
nand UO_1086 (O_1086,N_22049,N_23221);
nand UO_1087 (O_1087,N_23131,N_24291);
xor UO_1088 (O_1088,N_24018,N_24734);
and UO_1089 (O_1089,N_24072,N_22764);
or UO_1090 (O_1090,N_22197,N_23556);
or UO_1091 (O_1091,N_23290,N_22173);
and UO_1092 (O_1092,N_23538,N_24816);
and UO_1093 (O_1093,N_24138,N_24534);
nand UO_1094 (O_1094,N_22343,N_22753);
nand UO_1095 (O_1095,N_22806,N_22862);
and UO_1096 (O_1096,N_24351,N_24543);
and UO_1097 (O_1097,N_24284,N_23609);
nor UO_1098 (O_1098,N_24311,N_23436);
nand UO_1099 (O_1099,N_22925,N_22002);
or UO_1100 (O_1100,N_24749,N_23244);
or UO_1101 (O_1101,N_22110,N_24570);
nor UO_1102 (O_1102,N_22341,N_24563);
or UO_1103 (O_1103,N_23658,N_24530);
or UO_1104 (O_1104,N_24220,N_22847);
nor UO_1105 (O_1105,N_22831,N_24696);
nor UO_1106 (O_1106,N_23640,N_23495);
nand UO_1107 (O_1107,N_24911,N_22310);
or UO_1108 (O_1108,N_24125,N_22602);
and UO_1109 (O_1109,N_22186,N_24305);
nand UO_1110 (O_1110,N_23939,N_22512);
and UO_1111 (O_1111,N_22073,N_22896);
nor UO_1112 (O_1112,N_22907,N_23247);
nor UO_1113 (O_1113,N_22430,N_22811);
nand UO_1114 (O_1114,N_24106,N_22881);
and UO_1115 (O_1115,N_24094,N_23842);
and UO_1116 (O_1116,N_24212,N_23433);
nor UO_1117 (O_1117,N_24541,N_22679);
and UO_1118 (O_1118,N_23090,N_23531);
and UO_1119 (O_1119,N_21965,N_22187);
or UO_1120 (O_1120,N_23075,N_24608);
nor UO_1121 (O_1121,N_24301,N_23580);
or UO_1122 (O_1122,N_24814,N_24971);
nand UO_1123 (O_1123,N_22432,N_24887);
and UO_1124 (O_1124,N_22845,N_24736);
and UO_1125 (O_1125,N_23791,N_22481);
and UO_1126 (O_1126,N_24435,N_21911);
and UO_1127 (O_1127,N_22445,N_23703);
or UO_1128 (O_1128,N_24768,N_24737);
and UO_1129 (O_1129,N_24579,N_24640);
and UO_1130 (O_1130,N_24670,N_22271);
and UO_1131 (O_1131,N_24295,N_24895);
nand UO_1132 (O_1132,N_24994,N_22046);
and UO_1133 (O_1133,N_24620,N_24498);
nand UO_1134 (O_1134,N_23388,N_23478);
and UO_1135 (O_1135,N_24092,N_24602);
or UO_1136 (O_1136,N_23186,N_24412);
and UO_1137 (O_1137,N_24589,N_24705);
nand UO_1138 (O_1138,N_24322,N_23474);
nand UO_1139 (O_1139,N_22629,N_22560);
or UO_1140 (O_1140,N_24771,N_24792);
xor UO_1141 (O_1141,N_23193,N_23250);
nand UO_1142 (O_1142,N_24890,N_22867);
nor UO_1143 (O_1143,N_24713,N_21934);
nand UO_1144 (O_1144,N_22203,N_23069);
nand UO_1145 (O_1145,N_24140,N_23150);
nor UO_1146 (O_1146,N_24617,N_24203);
xor UO_1147 (O_1147,N_23670,N_24599);
and UO_1148 (O_1148,N_24605,N_24531);
nand UO_1149 (O_1149,N_23999,N_22011);
and UO_1150 (O_1150,N_24590,N_22624);
nand UO_1151 (O_1151,N_24578,N_24765);
or UO_1152 (O_1152,N_24269,N_22361);
and UO_1153 (O_1153,N_22191,N_22152);
nand UO_1154 (O_1154,N_24337,N_22577);
nor UO_1155 (O_1155,N_24998,N_23037);
and UO_1156 (O_1156,N_24352,N_24527);
nor UO_1157 (O_1157,N_24813,N_24860);
nor UO_1158 (O_1158,N_24358,N_23162);
nor UO_1159 (O_1159,N_23585,N_22075);
nor UO_1160 (O_1160,N_22647,N_24191);
nand UO_1161 (O_1161,N_22933,N_23320);
and UO_1162 (O_1162,N_24422,N_24962);
nand UO_1163 (O_1163,N_24730,N_23266);
and UO_1164 (O_1164,N_23625,N_22268);
and UO_1165 (O_1165,N_22810,N_21895);
or UO_1166 (O_1166,N_22779,N_23845);
and UO_1167 (O_1167,N_23129,N_23208);
nand UO_1168 (O_1168,N_24753,N_23603);
and UO_1169 (O_1169,N_24453,N_23719);
nand UO_1170 (O_1170,N_24135,N_22463);
nand UO_1171 (O_1171,N_22853,N_23679);
nand UO_1172 (O_1172,N_23523,N_24154);
and UO_1173 (O_1173,N_22664,N_23382);
nor UO_1174 (O_1174,N_24873,N_23441);
and UO_1175 (O_1175,N_23784,N_23800);
nor UO_1176 (O_1176,N_23969,N_24681);
nand UO_1177 (O_1177,N_23537,N_22193);
or UO_1178 (O_1178,N_22324,N_23882);
and UO_1179 (O_1179,N_23586,N_23505);
and UO_1180 (O_1180,N_24516,N_23870);
and UO_1181 (O_1181,N_22670,N_24153);
nor UO_1182 (O_1182,N_24920,N_24972);
or UO_1183 (O_1183,N_24585,N_22908);
nor UO_1184 (O_1184,N_22242,N_24168);
or UO_1185 (O_1185,N_22662,N_22741);
nor UO_1186 (O_1186,N_24331,N_24434);
and UO_1187 (O_1187,N_22395,N_23902);
nand UO_1188 (O_1188,N_22054,N_24612);
or UO_1189 (O_1189,N_24349,N_23261);
and UO_1190 (O_1190,N_24556,N_22849);
nor UO_1191 (O_1191,N_22768,N_23975);
nor UO_1192 (O_1192,N_24085,N_22436);
nor UO_1193 (O_1193,N_23081,N_22928);
xnor UO_1194 (O_1194,N_22758,N_24169);
or UO_1195 (O_1195,N_22821,N_24201);
xnor UO_1196 (O_1196,N_22274,N_22708);
and UO_1197 (O_1197,N_21928,N_23198);
nor UO_1198 (O_1198,N_22400,N_22232);
nor UO_1199 (O_1199,N_22179,N_24960);
or UO_1200 (O_1200,N_22993,N_24657);
or UO_1201 (O_1201,N_23705,N_24062);
or UO_1202 (O_1202,N_23831,N_24718);
xor UO_1203 (O_1203,N_24961,N_24951);
or UO_1204 (O_1204,N_24137,N_23600);
and UO_1205 (O_1205,N_23982,N_22334);
or UO_1206 (O_1206,N_24619,N_22939);
or UO_1207 (O_1207,N_23948,N_21991);
or UO_1208 (O_1208,N_23408,N_24115);
and UO_1209 (O_1209,N_22291,N_21875);
nor UO_1210 (O_1210,N_23426,N_24699);
nand UO_1211 (O_1211,N_22567,N_23411);
or UO_1212 (O_1212,N_23923,N_24184);
and UO_1213 (O_1213,N_22174,N_23958);
and UO_1214 (O_1214,N_24978,N_22721);
or UO_1215 (O_1215,N_24956,N_24937);
or UO_1216 (O_1216,N_23098,N_22354);
or UO_1217 (O_1217,N_22674,N_23107);
and UO_1218 (O_1218,N_24965,N_21957);
or UO_1219 (O_1219,N_24433,N_22678);
nor UO_1220 (O_1220,N_23189,N_24121);
or UO_1221 (O_1221,N_24919,N_23128);
nand UO_1222 (O_1222,N_24161,N_22367);
or UO_1223 (O_1223,N_22574,N_23547);
nor UO_1224 (O_1224,N_22804,N_21999);
xor UO_1225 (O_1225,N_22980,N_22774);
nand UO_1226 (O_1226,N_24158,N_23734);
or UO_1227 (O_1227,N_22829,N_24156);
nor UO_1228 (O_1228,N_22572,N_22137);
or UO_1229 (O_1229,N_23984,N_22506);
nor UO_1230 (O_1230,N_22828,N_24823);
nor UO_1231 (O_1231,N_23541,N_22029);
nor UO_1232 (O_1232,N_23249,N_23346);
nor UO_1233 (O_1233,N_23139,N_23680);
and UO_1234 (O_1234,N_23086,N_23903);
and UO_1235 (O_1235,N_24323,N_22609);
nand UO_1236 (O_1236,N_23682,N_23341);
or UO_1237 (O_1237,N_22059,N_21993);
and UO_1238 (O_1238,N_23038,N_22836);
nand UO_1239 (O_1239,N_23088,N_24854);
or UO_1240 (O_1240,N_24872,N_23287);
nor UO_1241 (O_1241,N_24839,N_24282);
nor UO_1242 (O_1242,N_24497,N_22196);
and UO_1243 (O_1243,N_23377,N_22301);
xnor UO_1244 (O_1244,N_23054,N_23691);
nand UO_1245 (O_1245,N_24462,N_24230);
xor UO_1246 (O_1246,N_24132,N_23797);
or UO_1247 (O_1247,N_23425,N_22293);
and UO_1248 (O_1248,N_22620,N_24310);
and UO_1249 (O_1249,N_23594,N_22891);
or UO_1250 (O_1250,N_22701,N_23447);
and UO_1251 (O_1251,N_22492,N_22717);
and UO_1252 (O_1252,N_22888,N_22202);
or UO_1253 (O_1253,N_24122,N_23407);
nor UO_1254 (O_1254,N_22901,N_24334);
nor UO_1255 (O_1255,N_24133,N_22675);
and UO_1256 (O_1256,N_22100,N_22530);
xnor UO_1257 (O_1257,N_22320,N_23061);
nand UO_1258 (O_1258,N_24401,N_22984);
nor UO_1259 (O_1259,N_23233,N_23059);
or UO_1260 (O_1260,N_21949,N_24967);
and UO_1261 (O_1261,N_23487,N_22127);
and UO_1262 (O_1262,N_23356,N_22866);
xor UO_1263 (O_1263,N_23032,N_23644);
nand UO_1264 (O_1264,N_24120,N_24087);
and UO_1265 (O_1265,N_22307,N_22963);
and UO_1266 (O_1266,N_23805,N_23762);
nor UO_1267 (O_1267,N_22349,N_22666);
and UO_1268 (O_1268,N_24259,N_23041);
nor UO_1269 (O_1269,N_22668,N_23783);
or UO_1270 (O_1270,N_23158,N_22563);
nor UO_1271 (O_1271,N_22794,N_24304);
and UO_1272 (O_1272,N_22006,N_23191);
and UO_1273 (O_1273,N_23307,N_24843);
nand UO_1274 (O_1274,N_23269,N_22189);
and UO_1275 (O_1275,N_24255,N_23467);
and UO_1276 (O_1276,N_24745,N_23353);
and UO_1277 (O_1277,N_22700,N_23087);
and UO_1278 (O_1278,N_22612,N_22782);
nand UO_1279 (O_1279,N_22034,N_23318);
or UO_1280 (O_1280,N_23078,N_22226);
nor UO_1281 (O_1281,N_22632,N_24999);
or UO_1282 (O_1282,N_23275,N_24829);
or UO_1283 (O_1283,N_22473,N_21887);
xor UO_1284 (O_1284,N_23554,N_23067);
nand UO_1285 (O_1285,N_23288,N_23024);
and UO_1286 (O_1286,N_24859,N_23486);
and UO_1287 (O_1287,N_22997,N_22044);
nand UO_1288 (O_1288,N_23416,N_23981);
and UO_1289 (O_1289,N_24976,N_23413);
or UO_1290 (O_1290,N_22529,N_22254);
xor UO_1291 (O_1291,N_24272,N_22188);
nor UO_1292 (O_1292,N_24402,N_23144);
nor UO_1293 (O_1293,N_24970,N_22440);
or UO_1294 (O_1294,N_21915,N_24679);
or UO_1295 (O_1295,N_24692,N_24069);
or UO_1296 (O_1296,N_24225,N_24123);
and UO_1297 (O_1297,N_23897,N_22206);
nand UO_1298 (O_1298,N_24207,N_22826);
and UO_1299 (O_1299,N_24558,N_23203);
or UO_1300 (O_1300,N_23497,N_22510);
and UO_1301 (O_1301,N_24483,N_22233);
and UO_1302 (O_1302,N_24245,N_23402);
nand UO_1303 (O_1303,N_24320,N_22423);
or UO_1304 (O_1304,N_22419,N_23728);
or UO_1305 (O_1305,N_23557,N_23830);
and UO_1306 (O_1306,N_21921,N_22905);
and UO_1307 (O_1307,N_24250,N_23743);
and UO_1308 (O_1308,N_22360,N_22585);
nor UO_1309 (O_1309,N_22961,N_24456);
or UO_1310 (O_1310,N_22383,N_23562);
nand UO_1311 (O_1311,N_24542,N_22030);
or UO_1312 (O_1312,N_23539,N_24512);
xnor UO_1313 (O_1313,N_23043,N_24052);
or UO_1314 (O_1314,N_24667,N_23694);
and UO_1315 (O_1315,N_23985,N_24423);
nor UO_1316 (O_1316,N_23631,N_24405);
and UO_1317 (O_1317,N_22243,N_22995);
and UO_1318 (O_1318,N_23739,N_22330);
nor UO_1319 (O_1319,N_22579,N_21972);
or UO_1320 (O_1320,N_23891,N_24463);
and UO_1321 (O_1321,N_21902,N_23937);
and UO_1322 (O_1322,N_23814,N_22956);
nor UO_1323 (O_1323,N_23029,N_23620);
and UO_1324 (O_1324,N_22515,N_22333);
and UO_1325 (O_1325,N_24267,N_22709);
nor UO_1326 (O_1326,N_22016,N_24045);
xnor UO_1327 (O_1327,N_22814,N_21945);
nand UO_1328 (O_1328,N_21912,N_24238);
nor UO_1329 (O_1329,N_24190,N_24326);
nor UO_1330 (O_1330,N_22218,N_22947);
nand UO_1331 (O_1331,N_23055,N_24162);
nor UO_1332 (O_1332,N_22446,N_22153);
or UO_1333 (O_1333,N_23358,N_24411);
or UO_1334 (O_1334,N_22757,N_24221);
nand UO_1335 (O_1335,N_23774,N_22735);
and UO_1336 (O_1336,N_23510,N_23590);
nand UO_1337 (O_1337,N_23593,N_23571);
nand UO_1338 (O_1338,N_24059,N_22715);
nor UO_1339 (O_1339,N_23256,N_24440);
or UO_1340 (O_1340,N_23807,N_24000);
xnor UO_1341 (O_1341,N_24938,N_22750);
xnor UO_1342 (O_1342,N_24339,N_23192);
or UO_1343 (O_1343,N_24447,N_24091);
or UO_1344 (O_1344,N_23274,N_21888);
nor UO_1345 (O_1345,N_21929,N_22331);
nor UO_1346 (O_1346,N_24869,N_22284);
or UO_1347 (O_1347,N_24791,N_22033);
and UO_1348 (O_1348,N_24841,N_22141);
nor UO_1349 (O_1349,N_22314,N_22457);
and UO_1350 (O_1350,N_22807,N_24703);
or UO_1351 (O_1351,N_23738,N_22981);
and UO_1352 (O_1352,N_22096,N_22375);
and UO_1353 (O_1353,N_24325,N_22047);
or UO_1354 (O_1354,N_24845,N_24174);
or UO_1355 (O_1355,N_24808,N_24746);
nor UO_1356 (O_1356,N_24459,N_24108);
or UO_1357 (O_1357,N_22994,N_23573);
nand UO_1358 (O_1358,N_24898,N_23704);
or UO_1359 (O_1359,N_24050,N_24346);
xor UO_1360 (O_1360,N_23512,N_23014);
xnor UO_1361 (O_1361,N_23473,N_24484);
nor UO_1362 (O_1362,N_24948,N_22641);
nand UO_1363 (O_1363,N_24126,N_23610);
or UO_1364 (O_1364,N_22633,N_23935);
or UO_1365 (O_1365,N_23522,N_21951);
nand UO_1366 (O_1366,N_23483,N_24618);
nor UO_1367 (O_1367,N_24354,N_23190);
nor UO_1368 (O_1368,N_23611,N_23785);
or UO_1369 (O_1369,N_23234,N_24702);
and UO_1370 (O_1370,N_24139,N_22922);
nand UO_1371 (O_1371,N_24076,N_21989);
nor UO_1372 (O_1372,N_24675,N_22321);
and UO_1373 (O_1373,N_21930,N_22377);
and UO_1374 (O_1374,N_24455,N_22259);
or UO_1375 (O_1375,N_22827,N_22160);
or UO_1376 (O_1376,N_22982,N_24925);
or UO_1377 (O_1377,N_23175,N_24393);
and UO_1378 (O_1378,N_24163,N_23506);
or UO_1379 (O_1379,N_23183,N_22121);
nor UO_1380 (O_1380,N_23953,N_22071);
nand UO_1381 (O_1381,N_22393,N_23010);
nand UO_1382 (O_1382,N_22287,N_22797);
or UO_1383 (O_1383,N_24017,N_22308);
and UO_1384 (O_1384,N_23861,N_22667);
or UO_1385 (O_1385,N_22505,N_22731);
and UO_1386 (O_1386,N_22502,N_24178);
and UO_1387 (O_1387,N_22682,N_22103);
nand UO_1388 (O_1388,N_22070,N_23000);
or UO_1389 (O_1389,N_24533,N_24376);
or UO_1390 (O_1390,N_23428,N_24129);
nand UO_1391 (O_1391,N_22863,N_21910);
nor UO_1392 (O_1392,N_24098,N_23171);
and UO_1393 (O_1393,N_23637,N_22999);
nor UO_1394 (O_1394,N_21890,N_22876);
or UO_1395 (O_1395,N_22053,N_23535);
or UO_1396 (O_1396,N_22558,N_23810);
or UO_1397 (O_1397,N_24136,N_22893);
nand UO_1398 (O_1398,N_22648,N_23764);
nand UO_1399 (O_1399,N_22610,N_22489);
and UO_1400 (O_1400,N_23598,N_24467);
nor UO_1401 (O_1401,N_24275,N_22775);
nand UO_1402 (O_1402,N_23788,N_23626);
nor UO_1403 (O_1403,N_23917,N_24482);
nand UO_1404 (O_1404,N_24893,N_23048);
and UO_1405 (O_1405,N_22417,N_23405);
and UO_1406 (O_1406,N_24399,N_22655);
nor UO_1407 (O_1407,N_23364,N_23050);
nor UO_1408 (O_1408,N_22626,N_24552);
nor UO_1409 (O_1409,N_23015,N_24490);
xnor UO_1410 (O_1410,N_22751,N_22285);
and UO_1411 (O_1411,N_23309,N_24997);
nand UO_1412 (O_1412,N_23689,N_23279);
or UO_1413 (O_1413,N_23378,N_22615);
or UO_1414 (O_1414,N_22730,N_24445);
nor UO_1415 (O_1415,N_22380,N_22714);
nand UO_1416 (O_1416,N_23255,N_23970);
nor UO_1417 (O_1417,N_24051,N_22345);
nor UO_1418 (O_1418,N_23476,N_23526);
or UO_1419 (O_1419,N_23583,N_22159);
or UO_1420 (O_1420,N_22872,N_23091);
xnor UO_1421 (O_1421,N_24613,N_22163);
xnor UO_1422 (O_1422,N_24815,N_24811);
nand UO_1423 (O_1423,N_22183,N_23393);
nand UO_1424 (O_1424,N_22449,N_23821);
nand UO_1425 (O_1425,N_21988,N_24549);
nand UO_1426 (O_1426,N_22733,N_22948);
and UO_1427 (O_1427,N_22673,N_23285);
nor UO_1428 (O_1428,N_22012,N_24297);
nand UO_1429 (O_1429,N_24719,N_23995);
nand UO_1430 (O_1430,N_24307,N_21908);
and UO_1431 (O_1431,N_21978,N_23977);
nand UO_1432 (O_1432,N_24454,N_24176);
and UO_1433 (O_1433,N_22931,N_22364);
and UO_1434 (O_1434,N_24720,N_23079);
nor UO_1435 (O_1435,N_23258,N_23730);
or UO_1436 (O_1436,N_23324,N_21935);
or UO_1437 (O_1437,N_24726,N_23623);
nor UO_1438 (O_1438,N_22977,N_22353);
nand UO_1439 (O_1439,N_22692,N_22401);
nand UO_1440 (O_1440,N_23453,N_23713);
or UO_1441 (O_1441,N_24802,N_22437);
nor UO_1442 (O_1442,N_23336,N_24078);
nor UO_1443 (O_1443,N_24047,N_23986);
nand UO_1444 (O_1444,N_23490,N_23884);
or UO_1445 (O_1445,N_22256,N_22761);
nand UO_1446 (O_1446,N_23246,N_24183);
and UO_1447 (O_1447,N_23864,N_24329);
and UO_1448 (O_1448,N_22870,N_24800);
nand UO_1449 (O_1449,N_24202,N_23546);
and UO_1450 (O_1450,N_22170,N_22919);
nand UO_1451 (O_1451,N_22500,N_24364);
and UO_1452 (O_1452,N_22825,N_22117);
xnor UO_1453 (O_1453,N_22077,N_24639);
and UO_1454 (O_1454,N_24661,N_24756);
nand UO_1455 (O_1455,N_23989,N_23101);
xor UO_1456 (O_1456,N_23491,N_23511);
xnor UO_1457 (O_1457,N_21900,N_24876);
and UO_1458 (O_1458,N_24683,N_24075);
or UO_1459 (O_1459,N_24160,N_23715);
nor UO_1460 (O_1460,N_23292,N_24428);
and UO_1461 (O_1461,N_24197,N_23502);
or UO_1462 (O_1462,N_23825,N_23673);
and UO_1463 (O_1463,N_23272,N_22738);
or UO_1464 (O_1464,N_22736,N_23379);
nor UO_1465 (O_1465,N_21981,N_24038);
nand UO_1466 (O_1466,N_24857,N_22225);
nor UO_1467 (O_1467,N_23801,N_23763);
and UO_1468 (O_1468,N_22278,N_22495);
or UO_1469 (O_1469,N_22158,N_23027);
or UO_1470 (O_1470,N_24851,N_22504);
xnor UO_1471 (O_1471,N_22114,N_24404);
and UO_1472 (O_1472,N_23847,N_24336);
nor UO_1473 (O_1473,N_23248,N_24610);
or UO_1474 (O_1474,N_23697,N_22778);
nor UO_1475 (O_1475,N_24674,N_24234);
xor UO_1476 (O_1476,N_24751,N_22973);
or UO_1477 (O_1477,N_22874,N_24101);
nand UO_1478 (O_1478,N_23383,N_22501);
nand UO_1479 (O_1479,N_23169,N_22760);
and UO_1480 (O_1480,N_23851,N_22857);
xor UO_1481 (O_1481,N_23462,N_22590);
xnor UO_1482 (O_1482,N_23744,N_23909);
nor UO_1483 (O_1483,N_21961,N_22132);
and UO_1484 (O_1484,N_22294,N_24443);
and UO_1485 (O_1485,N_22616,N_23036);
or UO_1486 (O_1486,N_22447,N_24488);
nand UO_1487 (O_1487,N_23776,N_23804);
or UO_1488 (O_1488,N_24277,N_22444);
and UO_1489 (O_1489,N_24365,N_22514);
nand UO_1490 (O_1490,N_22937,N_24324);
nor UO_1491 (O_1491,N_24479,N_21994);
nand UO_1492 (O_1492,N_22634,N_21897);
nor UO_1493 (O_1493,N_21899,N_23828);
xnor UO_1494 (O_1494,N_22317,N_22149);
and UO_1495 (O_1495,N_22435,N_22643);
or UO_1496 (O_1496,N_24298,N_23332);
or UO_1497 (O_1497,N_24023,N_22239);
or UO_1498 (O_1498,N_23578,N_23867);
nor UO_1499 (O_1499,N_21891,N_22488);
or UO_1500 (O_1500,N_22010,N_23472);
or UO_1501 (O_1501,N_23227,N_22082);
or UO_1502 (O_1502,N_22352,N_22455);
nor UO_1503 (O_1503,N_24653,N_22834);
and UO_1504 (O_1504,N_22823,N_22252);
or UO_1505 (O_1505,N_23463,N_21937);
nand UO_1506 (O_1506,N_22168,N_24368);
nor UO_1507 (O_1507,N_23317,N_22087);
nand UO_1508 (O_1508,N_22587,N_24464);
and UO_1509 (O_1509,N_22109,N_23846);
nor UO_1510 (O_1510,N_22859,N_24438);
or UO_1511 (O_1511,N_22538,N_22725);
xnor UO_1512 (O_1512,N_24974,N_22122);
nand UO_1513 (O_1513,N_23822,N_24485);
nor UO_1514 (O_1514,N_22707,N_23123);
or UO_1515 (O_1515,N_23389,N_23885);
or UO_1516 (O_1516,N_22723,N_22144);
and UO_1517 (O_1517,N_22822,N_22151);
and UO_1518 (O_1518,N_24374,N_23802);
and UO_1519 (O_1519,N_22472,N_24127);
or UO_1520 (O_1520,N_24604,N_23401);
or UO_1521 (O_1521,N_24731,N_24264);
xnor UO_1522 (O_1522,N_22111,N_22926);
nand UO_1523 (O_1523,N_24082,N_24279);
nand UO_1524 (O_1524,N_23671,N_23634);
and UO_1525 (O_1525,N_24982,N_22921);
or UO_1526 (O_1526,N_24114,N_23315);
and UO_1527 (O_1527,N_22710,N_23468);
and UO_1528 (O_1528,N_24711,N_23120);
and UO_1529 (O_1529,N_22522,N_23212);
and UO_1530 (O_1530,N_23470,N_23280);
nand UO_1531 (O_1531,N_23908,N_22690);
or UO_1532 (O_1532,N_24992,N_22816);
and UO_1533 (O_1533,N_22987,N_24748);
or UO_1534 (O_1534,N_23022,N_22555);
or UO_1535 (O_1535,N_22478,N_23527);
or UO_1536 (O_1536,N_24424,N_24386);
nand UO_1537 (O_1537,N_22245,N_24725);
nor UO_1538 (O_1538,N_23725,N_23653);
nand UO_1539 (O_1539,N_24783,N_23561);
or UO_1540 (O_1540,N_24356,N_22732);
xor UO_1541 (O_1541,N_22035,N_24819);
or UO_1542 (O_1542,N_23751,N_23717);
or UO_1543 (O_1543,N_22865,N_24015);
nand UO_1544 (O_1544,N_24902,N_24224);
nor UO_1545 (O_1545,N_23936,N_23551);
or UO_1546 (O_1546,N_22085,N_22166);
nand UO_1547 (O_1547,N_23850,N_24660);
nor UO_1548 (O_1548,N_22516,N_24383);
and UO_1549 (O_1549,N_21976,N_24929);
and UO_1550 (O_1550,N_24427,N_23566);
nand UO_1551 (O_1551,N_23508,N_24328);
and UO_1552 (O_1552,N_23695,N_22374);
or UO_1553 (O_1553,N_24694,N_21926);
or UO_1554 (O_1554,N_22833,N_24348);
nand UO_1555 (O_1555,N_23045,N_22185);
and UO_1556 (O_1556,N_23068,N_24858);
or UO_1557 (O_1557,N_24852,N_22787);
or UO_1558 (O_1558,N_23446,N_24724);
and UO_1559 (O_1559,N_24964,N_24656);
nor UO_1560 (O_1560,N_21923,N_23616);
or UO_1561 (O_1561,N_22458,N_22658);
nor UO_1562 (O_1562,N_22742,N_24111);
nand UO_1563 (O_1563,N_24887,N_24954);
xor UO_1564 (O_1564,N_24977,N_23558);
xnor UO_1565 (O_1565,N_22350,N_23846);
nor UO_1566 (O_1566,N_22853,N_24698);
nand UO_1567 (O_1567,N_24354,N_23346);
and UO_1568 (O_1568,N_24693,N_23553);
xnor UO_1569 (O_1569,N_22536,N_24674);
or UO_1570 (O_1570,N_24173,N_24972);
nand UO_1571 (O_1571,N_24824,N_22397);
and UO_1572 (O_1572,N_24449,N_22220);
nor UO_1573 (O_1573,N_22063,N_24228);
xnor UO_1574 (O_1574,N_22892,N_22883);
nor UO_1575 (O_1575,N_22995,N_22552);
nand UO_1576 (O_1576,N_22293,N_24272);
or UO_1577 (O_1577,N_24339,N_24552);
or UO_1578 (O_1578,N_23258,N_22766);
nand UO_1579 (O_1579,N_23677,N_24079);
and UO_1580 (O_1580,N_23769,N_23949);
nor UO_1581 (O_1581,N_24766,N_24819);
nand UO_1582 (O_1582,N_22234,N_24892);
and UO_1583 (O_1583,N_23736,N_24573);
and UO_1584 (O_1584,N_23318,N_23836);
nand UO_1585 (O_1585,N_24037,N_23914);
and UO_1586 (O_1586,N_23670,N_22994);
nand UO_1587 (O_1587,N_24677,N_24917);
or UO_1588 (O_1588,N_22281,N_23465);
and UO_1589 (O_1589,N_23581,N_22809);
or UO_1590 (O_1590,N_22564,N_23383);
nand UO_1591 (O_1591,N_22113,N_22492);
nand UO_1592 (O_1592,N_23254,N_22335);
nand UO_1593 (O_1593,N_24819,N_24400);
and UO_1594 (O_1594,N_22812,N_24062);
and UO_1595 (O_1595,N_22490,N_21920);
and UO_1596 (O_1596,N_24297,N_22105);
xor UO_1597 (O_1597,N_24506,N_22293);
and UO_1598 (O_1598,N_23936,N_23950);
or UO_1599 (O_1599,N_23181,N_22862);
or UO_1600 (O_1600,N_22787,N_23202);
or UO_1601 (O_1601,N_23200,N_22289);
nand UO_1602 (O_1602,N_24009,N_23775);
or UO_1603 (O_1603,N_24415,N_22285);
nand UO_1604 (O_1604,N_23628,N_22052);
or UO_1605 (O_1605,N_24975,N_23978);
and UO_1606 (O_1606,N_21916,N_22259);
nor UO_1607 (O_1607,N_24161,N_24392);
and UO_1608 (O_1608,N_22722,N_22048);
nor UO_1609 (O_1609,N_23535,N_24999);
or UO_1610 (O_1610,N_24709,N_24286);
and UO_1611 (O_1611,N_23540,N_22312);
and UO_1612 (O_1612,N_23380,N_21983);
or UO_1613 (O_1613,N_24557,N_22035);
or UO_1614 (O_1614,N_23450,N_23680);
and UO_1615 (O_1615,N_24461,N_23684);
nand UO_1616 (O_1616,N_22591,N_22903);
nor UO_1617 (O_1617,N_23443,N_24668);
and UO_1618 (O_1618,N_24014,N_22108);
xnor UO_1619 (O_1619,N_22021,N_24682);
or UO_1620 (O_1620,N_24622,N_23574);
and UO_1621 (O_1621,N_22894,N_23445);
nor UO_1622 (O_1622,N_23886,N_23264);
nand UO_1623 (O_1623,N_23112,N_22550);
nand UO_1624 (O_1624,N_24583,N_24966);
nand UO_1625 (O_1625,N_21914,N_22427);
nor UO_1626 (O_1626,N_23384,N_22150);
nand UO_1627 (O_1627,N_22726,N_24731);
and UO_1628 (O_1628,N_24360,N_24178);
and UO_1629 (O_1629,N_22744,N_24705);
or UO_1630 (O_1630,N_23965,N_23555);
nand UO_1631 (O_1631,N_24763,N_24222);
and UO_1632 (O_1632,N_23928,N_23236);
and UO_1633 (O_1633,N_23279,N_21980);
or UO_1634 (O_1634,N_23868,N_22063);
or UO_1635 (O_1635,N_22205,N_23599);
or UO_1636 (O_1636,N_22645,N_22682);
nand UO_1637 (O_1637,N_24143,N_22042);
nand UO_1638 (O_1638,N_23292,N_22104);
xnor UO_1639 (O_1639,N_22771,N_22955);
or UO_1640 (O_1640,N_23587,N_23110);
nor UO_1641 (O_1641,N_22424,N_23292);
xor UO_1642 (O_1642,N_24536,N_24547);
nand UO_1643 (O_1643,N_21941,N_23634);
and UO_1644 (O_1644,N_21892,N_22267);
and UO_1645 (O_1645,N_23574,N_22474);
or UO_1646 (O_1646,N_22546,N_22388);
and UO_1647 (O_1647,N_24161,N_24641);
nand UO_1648 (O_1648,N_24075,N_22818);
or UO_1649 (O_1649,N_22759,N_22682);
nor UO_1650 (O_1650,N_21924,N_22675);
nand UO_1651 (O_1651,N_22384,N_23666);
and UO_1652 (O_1652,N_23954,N_23002);
nor UO_1653 (O_1653,N_22432,N_24536);
nor UO_1654 (O_1654,N_22503,N_24381);
and UO_1655 (O_1655,N_24894,N_23456);
nand UO_1656 (O_1656,N_24800,N_23694);
or UO_1657 (O_1657,N_24573,N_24499);
or UO_1658 (O_1658,N_24884,N_24584);
nand UO_1659 (O_1659,N_23729,N_24743);
and UO_1660 (O_1660,N_24336,N_24977);
or UO_1661 (O_1661,N_24995,N_23106);
nor UO_1662 (O_1662,N_22260,N_23173);
or UO_1663 (O_1663,N_22310,N_22697);
or UO_1664 (O_1664,N_22433,N_24542);
and UO_1665 (O_1665,N_23471,N_22686);
and UO_1666 (O_1666,N_23364,N_23292);
and UO_1667 (O_1667,N_22508,N_23682);
nand UO_1668 (O_1668,N_22006,N_24577);
nand UO_1669 (O_1669,N_23228,N_23203);
nor UO_1670 (O_1670,N_23803,N_24005);
xor UO_1671 (O_1671,N_22530,N_24034);
and UO_1672 (O_1672,N_24285,N_22016);
nand UO_1673 (O_1673,N_22175,N_24359);
nand UO_1674 (O_1674,N_23917,N_24652);
nor UO_1675 (O_1675,N_24301,N_24565);
nand UO_1676 (O_1676,N_22228,N_22611);
nand UO_1677 (O_1677,N_24297,N_23486);
and UO_1678 (O_1678,N_22390,N_24188);
or UO_1679 (O_1679,N_24151,N_24218);
and UO_1680 (O_1680,N_24672,N_22012);
nor UO_1681 (O_1681,N_22408,N_23151);
nor UO_1682 (O_1682,N_22538,N_23552);
or UO_1683 (O_1683,N_22517,N_22008);
nand UO_1684 (O_1684,N_23338,N_22140);
nor UO_1685 (O_1685,N_22957,N_23337);
or UO_1686 (O_1686,N_23232,N_22651);
nand UO_1687 (O_1687,N_24409,N_24480);
nand UO_1688 (O_1688,N_23925,N_24344);
nor UO_1689 (O_1689,N_24563,N_23272);
or UO_1690 (O_1690,N_24009,N_24702);
and UO_1691 (O_1691,N_24591,N_24885);
nor UO_1692 (O_1692,N_24375,N_23011);
and UO_1693 (O_1693,N_21883,N_23306);
nor UO_1694 (O_1694,N_23887,N_23015);
nand UO_1695 (O_1695,N_24586,N_22446);
xnor UO_1696 (O_1696,N_24088,N_24754);
xnor UO_1697 (O_1697,N_21993,N_24942);
and UO_1698 (O_1698,N_24623,N_23894);
or UO_1699 (O_1699,N_23461,N_23266);
or UO_1700 (O_1700,N_23642,N_23695);
nor UO_1701 (O_1701,N_23098,N_24811);
and UO_1702 (O_1702,N_22808,N_24821);
nand UO_1703 (O_1703,N_23323,N_23015);
or UO_1704 (O_1704,N_22639,N_24888);
or UO_1705 (O_1705,N_22278,N_22842);
nor UO_1706 (O_1706,N_23178,N_23130);
or UO_1707 (O_1707,N_24810,N_24648);
and UO_1708 (O_1708,N_23038,N_24499);
xor UO_1709 (O_1709,N_22559,N_23456);
nor UO_1710 (O_1710,N_22263,N_22271);
nor UO_1711 (O_1711,N_24146,N_24577);
and UO_1712 (O_1712,N_24957,N_24475);
nand UO_1713 (O_1713,N_24489,N_22742);
or UO_1714 (O_1714,N_22567,N_22408);
or UO_1715 (O_1715,N_22712,N_23090);
or UO_1716 (O_1716,N_24747,N_23666);
or UO_1717 (O_1717,N_23333,N_21901);
xor UO_1718 (O_1718,N_24265,N_24972);
or UO_1719 (O_1719,N_22215,N_23235);
xor UO_1720 (O_1720,N_23809,N_24123);
and UO_1721 (O_1721,N_23371,N_22061);
or UO_1722 (O_1722,N_22748,N_24189);
or UO_1723 (O_1723,N_23215,N_23995);
or UO_1724 (O_1724,N_23357,N_24089);
nand UO_1725 (O_1725,N_24010,N_23083);
nand UO_1726 (O_1726,N_23754,N_21911);
nand UO_1727 (O_1727,N_24737,N_23483);
xnor UO_1728 (O_1728,N_22696,N_24983);
and UO_1729 (O_1729,N_22975,N_24349);
nand UO_1730 (O_1730,N_23807,N_24642);
and UO_1731 (O_1731,N_22349,N_24040);
nand UO_1732 (O_1732,N_23997,N_24166);
or UO_1733 (O_1733,N_22884,N_24140);
nand UO_1734 (O_1734,N_24748,N_24727);
or UO_1735 (O_1735,N_22142,N_23162);
nand UO_1736 (O_1736,N_23136,N_24849);
nor UO_1737 (O_1737,N_23189,N_22090);
and UO_1738 (O_1738,N_24203,N_22439);
nor UO_1739 (O_1739,N_23150,N_22019);
nor UO_1740 (O_1740,N_24232,N_22009);
xor UO_1741 (O_1741,N_24823,N_24705);
nor UO_1742 (O_1742,N_23273,N_23827);
or UO_1743 (O_1743,N_23325,N_24670);
xor UO_1744 (O_1744,N_21976,N_23531);
and UO_1745 (O_1745,N_24815,N_22184);
xor UO_1746 (O_1746,N_24760,N_23968);
nor UO_1747 (O_1747,N_23805,N_23440);
nand UO_1748 (O_1748,N_21918,N_24506);
and UO_1749 (O_1749,N_22645,N_24956);
nand UO_1750 (O_1750,N_23298,N_24656);
or UO_1751 (O_1751,N_24798,N_24510);
and UO_1752 (O_1752,N_23517,N_22839);
nand UO_1753 (O_1753,N_21921,N_23331);
or UO_1754 (O_1754,N_24444,N_22557);
nand UO_1755 (O_1755,N_22624,N_22339);
nand UO_1756 (O_1756,N_24854,N_24030);
xor UO_1757 (O_1757,N_22795,N_24359);
nor UO_1758 (O_1758,N_24462,N_24290);
nand UO_1759 (O_1759,N_24733,N_23443);
or UO_1760 (O_1760,N_22587,N_21991);
xnor UO_1761 (O_1761,N_21877,N_24431);
nor UO_1762 (O_1762,N_24586,N_24073);
or UO_1763 (O_1763,N_23627,N_24499);
or UO_1764 (O_1764,N_22870,N_22485);
and UO_1765 (O_1765,N_23152,N_22126);
and UO_1766 (O_1766,N_23464,N_23526);
or UO_1767 (O_1767,N_22864,N_23540);
nand UO_1768 (O_1768,N_24304,N_22711);
nand UO_1769 (O_1769,N_23379,N_24258);
and UO_1770 (O_1770,N_23403,N_22176);
or UO_1771 (O_1771,N_22046,N_24834);
or UO_1772 (O_1772,N_24307,N_24731);
or UO_1773 (O_1773,N_23855,N_22557);
xor UO_1774 (O_1774,N_23508,N_22194);
xor UO_1775 (O_1775,N_24755,N_22129);
and UO_1776 (O_1776,N_22280,N_22362);
or UO_1777 (O_1777,N_22572,N_22750);
xor UO_1778 (O_1778,N_24142,N_22007);
nand UO_1779 (O_1779,N_24014,N_22668);
and UO_1780 (O_1780,N_22975,N_22749);
nor UO_1781 (O_1781,N_22090,N_22047);
and UO_1782 (O_1782,N_23738,N_23650);
nand UO_1783 (O_1783,N_22474,N_24485);
xnor UO_1784 (O_1784,N_24348,N_22530);
nand UO_1785 (O_1785,N_23864,N_22981);
xor UO_1786 (O_1786,N_22632,N_23738);
or UO_1787 (O_1787,N_22664,N_22966);
nor UO_1788 (O_1788,N_23346,N_22718);
nand UO_1789 (O_1789,N_24179,N_24648);
nor UO_1790 (O_1790,N_21970,N_22843);
nand UO_1791 (O_1791,N_24807,N_22237);
nor UO_1792 (O_1792,N_24026,N_22955);
nand UO_1793 (O_1793,N_22717,N_23345);
nor UO_1794 (O_1794,N_24935,N_23032);
nor UO_1795 (O_1795,N_23657,N_22470);
and UO_1796 (O_1796,N_22015,N_22555);
nor UO_1797 (O_1797,N_24259,N_24362);
nor UO_1798 (O_1798,N_24069,N_22280);
and UO_1799 (O_1799,N_23264,N_23929);
and UO_1800 (O_1800,N_23219,N_22162);
nand UO_1801 (O_1801,N_23849,N_22149);
nor UO_1802 (O_1802,N_23603,N_24340);
nor UO_1803 (O_1803,N_23916,N_24046);
nand UO_1804 (O_1804,N_24190,N_23455);
nor UO_1805 (O_1805,N_23420,N_23851);
nand UO_1806 (O_1806,N_24707,N_24199);
xnor UO_1807 (O_1807,N_22002,N_24495);
nand UO_1808 (O_1808,N_23325,N_21966);
xor UO_1809 (O_1809,N_24816,N_22160);
or UO_1810 (O_1810,N_22753,N_22249);
or UO_1811 (O_1811,N_22198,N_24051);
or UO_1812 (O_1812,N_23869,N_23467);
and UO_1813 (O_1813,N_23311,N_22340);
or UO_1814 (O_1814,N_23171,N_22293);
nor UO_1815 (O_1815,N_23879,N_22573);
nand UO_1816 (O_1816,N_23593,N_22754);
and UO_1817 (O_1817,N_22403,N_24528);
and UO_1818 (O_1818,N_23793,N_24294);
xor UO_1819 (O_1819,N_24177,N_24133);
xnor UO_1820 (O_1820,N_23755,N_22185);
and UO_1821 (O_1821,N_23036,N_22568);
xor UO_1822 (O_1822,N_22935,N_22623);
xor UO_1823 (O_1823,N_23204,N_23623);
nor UO_1824 (O_1824,N_23570,N_23462);
nor UO_1825 (O_1825,N_24956,N_22677);
xor UO_1826 (O_1826,N_24563,N_22260);
nor UO_1827 (O_1827,N_22710,N_22025);
and UO_1828 (O_1828,N_24717,N_22838);
nor UO_1829 (O_1829,N_24967,N_24018);
nor UO_1830 (O_1830,N_22106,N_24285);
nor UO_1831 (O_1831,N_24517,N_23818);
and UO_1832 (O_1832,N_24311,N_24569);
and UO_1833 (O_1833,N_24168,N_23672);
nand UO_1834 (O_1834,N_24540,N_22780);
or UO_1835 (O_1835,N_23095,N_22845);
and UO_1836 (O_1836,N_22884,N_23128);
nand UO_1837 (O_1837,N_24932,N_23569);
and UO_1838 (O_1838,N_22790,N_24531);
nor UO_1839 (O_1839,N_23858,N_22542);
nor UO_1840 (O_1840,N_24966,N_22690);
and UO_1841 (O_1841,N_24384,N_24304);
nor UO_1842 (O_1842,N_24386,N_24691);
xor UO_1843 (O_1843,N_22149,N_22761);
and UO_1844 (O_1844,N_24657,N_24359);
nand UO_1845 (O_1845,N_22302,N_23821);
nand UO_1846 (O_1846,N_22678,N_23097);
nand UO_1847 (O_1847,N_23251,N_23439);
or UO_1848 (O_1848,N_24487,N_23357);
nor UO_1849 (O_1849,N_24091,N_24281);
nor UO_1850 (O_1850,N_23969,N_24655);
nand UO_1851 (O_1851,N_22407,N_21921);
or UO_1852 (O_1852,N_22959,N_23300);
xor UO_1853 (O_1853,N_24820,N_23583);
and UO_1854 (O_1854,N_22697,N_22194);
xor UO_1855 (O_1855,N_23774,N_23289);
and UO_1856 (O_1856,N_22739,N_22496);
nor UO_1857 (O_1857,N_24969,N_23234);
nand UO_1858 (O_1858,N_22665,N_24535);
and UO_1859 (O_1859,N_22780,N_22449);
and UO_1860 (O_1860,N_24570,N_23517);
or UO_1861 (O_1861,N_22071,N_22197);
nand UO_1862 (O_1862,N_23669,N_23181);
xnor UO_1863 (O_1863,N_22647,N_22203);
or UO_1864 (O_1864,N_23066,N_24884);
or UO_1865 (O_1865,N_24156,N_22123);
or UO_1866 (O_1866,N_22657,N_24969);
or UO_1867 (O_1867,N_23975,N_23384);
xor UO_1868 (O_1868,N_23687,N_24296);
or UO_1869 (O_1869,N_23359,N_23994);
and UO_1870 (O_1870,N_22725,N_22695);
xnor UO_1871 (O_1871,N_22933,N_22807);
or UO_1872 (O_1872,N_24357,N_23602);
xor UO_1873 (O_1873,N_24245,N_23737);
and UO_1874 (O_1874,N_22423,N_23265);
nand UO_1875 (O_1875,N_22912,N_24704);
and UO_1876 (O_1876,N_23455,N_22906);
and UO_1877 (O_1877,N_23096,N_22823);
nand UO_1878 (O_1878,N_23657,N_22850);
nor UO_1879 (O_1879,N_22697,N_22665);
nand UO_1880 (O_1880,N_21962,N_24846);
or UO_1881 (O_1881,N_21959,N_24974);
nand UO_1882 (O_1882,N_22621,N_24246);
or UO_1883 (O_1883,N_23646,N_23492);
or UO_1884 (O_1884,N_22378,N_22318);
nor UO_1885 (O_1885,N_21939,N_23553);
nand UO_1886 (O_1886,N_24510,N_22441);
xor UO_1887 (O_1887,N_22901,N_22643);
nand UO_1888 (O_1888,N_22047,N_24414);
nor UO_1889 (O_1889,N_21937,N_24320);
nand UO_1890 (O_1890,N_22305,N_22700);
and UO_1891 (O_1891,N_24371,N_24971);
xor UO_1892 (O_1892,N_24573,N_24779);
and UO_1893 (O_1893,N_24654,N_23701);
or UO_1894 (O_1894,N_24611,N_24792);
or UO_1895 (O_1895,N_22343,N_24582);
nor UO_1896 (O_1896,N_23732,N_22468);
or UO_1897 (O_1897,N_22397,N_22957);
and UO_1898 (O_1898,N_22967,N_24658);
xnor UO_1899 (O_1899,N_24935,N_22817);
and UO_1900 (O_1900,N_22051,N_24982);
nor UO_1901 (O_1901,N_23119,N_24656);
xnor UO_1902 (O_1902,N_23901,N_23417);
nor UO_1903 (O_1903,N_24890,N_23635);
nor UO_1904 (O_1904,N_24795,N_22268);
nand UO_1905 (O_1905,N_24186,N_24443);
nand UO_1906 (O_1906,N_24869,N_24642);
nand UO_1907 (O_1907,N_24409,N_22064);
nor UO_1908 (O_1908,N_23288,N_23586);
or UO_1909 (O_1909,N_23105,N_22944);
nor UO_1910 (O_1910,N_21983,N_24395);
xor UO_1911 (O_1911,N_21909,N_21960);
and UO_1912 (O_1912,N_24000,N_23501);
or UO_1913 (O_1913,N_24835,N_24654);
nor UO_1914 (O_1914,N_22595,N_24437);
nand UO_1915 (O_1915,N_22839,N_23996);
and UO_1916 (O_1916,N_22652,N_23744);
and UO_1917 (O_1917,N_24092,N_23944);
xor UO_1918 (O_1918,N_24582,N_22866);
nand UO_1919 (O_1919,N_22788,N_24950);
nor UO_1920 (O_1920,N_22319,N_22764);
and UO_1921 (O_1921,N_24133,N_23738);
and UO_1922 (O_1922,N_22812,N_22229);
nand UO_1923 (O_1923,N_23156,N_24723);
and UO_1924 (O_1924,N_24043,N_23155);
nor UO_1925 (O_1925,N_22349,N_24558);
or UO_1926 (O_1926,N_23979,N_23429);
or UO_1927 (O_1927,N_23547,N_22143);
and UO_1928 (O_1928,N_23329,N_22705);
and UO_1929 (O_1929,N_24992,N_22217);
nor UO_1930 (O_1930,N_23658,N_22344);
nand UO_1931 (O_1931,N_23993,N_23657);
and UO_1932 (O_1932,N_24137,N_22751);
nor UO_1933 (O_1933,N_23670,N_22274);
and UO_1934 (O_1934,N_24891,N_22615);
xor UO_1935 (O_1935,N_24501,N_23423);
nand UO_1936 (O_1936,N_22197,N_24331);
nor UO_1937 (O_1937,N_22653,N_24060);
or UO_1938 (O_1938,N_22170,N_22241);
or UO_1939 (O_1939,N_22489,N_24981);
nor UO_1940 (O_1940,N_23925,N_24919);
nand UO_1941 (O_1941,N_22717,N_23097);
nor UO_1942 (O_1942,N_23876,N_23453);
and UO_1943 (O_1943,N_24198,N_24853);
nor UO_1944 (O_1944,N_22666,N_22881);
nand UO_1945 (O_1945,N_22304,N_24428);
xnor UO_1946 (O_1946,N_23658,N_24439);
or UO_1947 (O_1947,N_22278,N_22357);
and UO_1948 (O_1948,N_23187,N_22874);
nand UO_1949 (O_1949,N_22966,N_23603);
nor UO_1950 (O_1950,N_22268,N_23651);
xor UO_1951 (O_1951,N_23252,N_24682);
nand UO_1952 (O_1952,N_24742,N_23817);
and UO_1953 (O_1953,N_22620,N_23790);
nand UO_1954 (O_1954,N_23441,N_24383);
and UO_1955 (O_1955,N_21984,N_22300);
and UO_1956 (O_1956,N_24475,N_22128);
or UO_1957 (O_1957,N_24440,N_22713);
and UO_1958 (O_1958,N_22603,N_21887);
nor UO_1959 (O_1959,N_24545,N_24900);
or UO_1960 (O_1960,N_23429,N_23875);
nand UO_1961 (O_1961,N_24446,N_24863);
or UO_1962 (O_1962,N_24457,N_22954);
nand UO_1963 (O_1963,N_24032,N_22482);
and UO_1964 (O_1964,N_22417,N_24924);
or UO_1965 (O_1965,N_23967,N_24744);
nor UO_1966 (O_1966,N_22187,N_21974);
nand UO_1967 (O_1967,N_24040,N_24108);
nor UO_1968 (O_1968,N_24489,N_24980);
and UO_1969 (O_1969,N_22777,N_22940);
or UO_1970 (O_1970,N_23313,N_24113);
nand UO_1971 (O_1971,N_21963,N_22358);
nor UO_1972 (O_1972,N_24387,N_21888);
or UO_1973 (O_1973,N_23924,N_24624);
nor UO_1974 (O_1974,N_24913,N_24266);
and UO_1975 (O_1975,N_22954,N_23911);
nor UO_1976 (O_1976,N_22454,N_23223);
nor UO_1977 (O_1977,N_24050,N_22045);
nand UO_1978 (O_1978,N_23299,N_23594);
nand UO_1979 (O_1979,N_22401,N_23923);
nor UO_1980 (O_1980,N_23947,N_24195);
nand UO_1981 (O_1981,N_23966,N_22305);
or UO_1982 (O_1982,N_23770,N_23277);
xor UO_1983 (O_1983,N_22368,N_24366);
nor UO_1984 (O_1984,N_24788,N_21880);
nor UO_1985 (O_1985,N_23868,N_22648);
and UO_1986 (O_1986,N_23352,N_24939);
nor UO_1987 (O_1987,N_24702,N_22164);
or UO_1988 (O_1988,N_23418,N_24450);
and UO_1989 (O_1989,N_22964,N_22839);
nand UO_1990 (O_1990,N_22893,N_24149);
nand UO_1991 (O_1991,N_23481,N_24209);
or UO_1992 (O_1992,N_22045,N_22264);
nand UO_1993 (O_1993,N_23025,N_22209);
nor UO_1994 (O_1994,N_22821,N_24581);
and UO_1995 (O_1995,N_23141,N_23034);
nor UO_1996 (O_1996,N_22370,N_21881);
nand UO_1997 (O_1997,N_22392,N_22198);
and UO_1998 (O_1998,N_23011,N_23671);
xnor UO_1999 (O_1999,N_22182,N_23973);
xor UO_2000 (O_2000,N_23848,N_23558);
nand UO_2001 (O_2001,N_23611,N_21875);
xnor UO_2002 (O_2002,N_24226,N_24512);
nand UO_2003 (O_2003,N_24370,N_23391);
nand UO_2004 (O_2004,N_22417,N_24213);
or UO_2005 (O_2005,N_24674,N_24783);
nand UO_2006 (O_2006,N_23728,N_22450);
and UO_2007 (O_2007,N_22746,N_22031);
or UO_2008 (O_2008,N_23330,N_22173);
or UO_2009 (O_2009,N_24527,N_23820);
or UO_2010 (O_2010,N_22278,N_23019);
and UO_2011 (O_2011,N_22079,N_24816);
xnor UO_2012 (O_2012,N_22388,N_23113);
nand UO_2013 (O_2013,N_23846,N_22850);
and UO_2014 (O_2014,N_22437,N_24975);
nand UO_2015 (O_2015,N_23357,N_24578);
xor UO_2016 (O_2016,N_24335,N_21981);
or UO_2017 (O_2017,N_24570,N_24704);
nand UO_2018 (O_2018,N_22669,N_24312);
or UO_2019 (O_2019,N_23589,N_22983);
and UO_2020 (O_2020,N_24040,N_23841);
nand UO_2021 (O_2021,N_24587,N_24902);
and UO_2022 (O_2022,N_24053,N_22345);
and UO_2023 (O_2023,N_22937,N_22296);
xnor UO_2024 (O_2024,N_24720,N_22151);
or UO_2025 (O_2025,N_24401,N_22109);
nand UO_2026 (O_2026,N_23461,N_24467);
nand UO_2027 (O_2027,N_24127,N_23583);
nand UO_2028 (O_2028,N_24183,N_23504);
or UO_2029 (O_2029,N_22566,N_24578);
xnor UO_2030 (O_2030,N_22926,N_24067);
nand UO_2031 (O_2031,N_24953,N_24070);
or UO_2032 (O_2032,N_22708,N_22246);
and UO_2033 (O_2033,N_23896,N_23037);
nand UO_2034 (O_2034,N_24627,N_23391);
nor UO_2035 (O_2035,N_24858,N_23943);
and UO_2036 (O_2036,N_22169,N_24789);
nor UO_2037 (O_2037,N_23381,N_23297);
nand UO_2038 (O_2038,N_23495,N_24558);
nand UO_2039 (O_2039,N_22745,N_23230);
or UO_2040 (O_2040,N_23402,N_23916);
or UO_2041 (O_2041,N_24606,N_24129);
or UO_2042 (O_2042,N_24501,N_22611);
xnor UO_2043 (O_2043,N_22018,N_24337);
and UO_2044 (O_2044,N_23040,N_23402);
or UO_2045 (O_2045,N_24742,N_22948);
or UO_2046 (O_2046,N_23074,N_22589);
or UO_2047 (O_2047,N_23468,N_24978);
nand UO_2048 (O_2048,N_24961,N_21961);
and UO_2049 (O_2049,N_23130,N_23612);
or UO_2050 (O_2050,N_24378,N_24133);
and UO_2051 (O_2051,N_22176,N_22846);
or UO_2052 (O_2052,N_24522,N_24051);
nor UO_2053 (O_2053,N_22730,N_22075);
or UO_2054 (O_2054,N_22346,N_23598);
nor UO_2055 (O_2055,N_24139,N_24991);
nor UO_2056 (O_2056,N_24408,N_24055);
nor UO_2057 (O_2057,N_22800,N_23653);
or UO_2058 (O_2058,N_23532,N_22534);
and UO_2059 (O_2059,N_23028,N_23228);
nor UO_2060 (O_2060,N_23143,N_24250);
nand UO_2061 (O_2061,N_23343,N_22793);
and UO_2062 (O_2062,N_24587,N_24870);
nand UO_2063 (O_2063,N_24230,N_24254);
and UO_2064 (O_2064,N_22948,N_24584);
and UO_2065 (O_2065,N_24271,N_24934);
or UO_2066 (O_2066,N_23891,N_23955);
and UO_2067 (O_2067,N_23763,N_23049);
nor UO_2068 (O_2068,N_24246,N_23150);
nand UO_2069 (O_2069,N_24661,N_22354);
or UO_2070 (O_2070,N_24393,N_23850);
nand UO_2071 (O_2071,N_24334,N_22076);
nor UO_2072 (O_2072,N_22444,N_24954);
and UO_2073 (O_2073,N_23114,N_23492);
and UO_2074 (O_2074,N_24446,N_22858);
nor UO_2075 (O_2075,N_22094,N_24455);
nor UO_2076 (O_2076,N_22554,N_22244);
nor UO_2077 (O_2077,N_23013,N_22732);
nand UO_2078 (O_2078,N_23454,N_22221);
nor UO_2079 (O_2079,N_24202,N_24833);
nand UO_2080 (O_2080,N_22233,N_23987);
or UO_2081 (O_2081,N_21894,N_23381);
and UO_2082 (O_2082,N_23249,N_24779);
and UO_2083 (O_2083,N_22811,N_21914);
nor UO_2084 (O_2084,N_24869,N_24817);
and UO_2085 (O_2085,N_24903,N_23007);
xor UO_2086 (O_2086,N_24580,N_24004);
nand UO_2087 (O_2087,N_22040,N_23948);
nand UO_2088 (O_2088,N_24833,N_21878);
xnor UO_2089 (O_2089,N_24916,N_23778);
and UO_2090 (O_2090,N_23247,N_21919);
and UO_2091 (O_2091,N_23050,N_22642);
nor UO_2092 (O_2092,N_23798,N_22821);
and UO_2093 (O_2093,N_24255,N_22000);
nand UO_2094 (O_2094,N_23688,N_24555);
or UO_2095 (O_2095,N_24109,N_22545);
nor UO_2096 (O_2096,N_22649,N_23704);
xnor UO_2097 (O_2097,N_24683,N_24602);
and UO_2098 (O_2098,N_22971,N_23012);
nor UO_2099 (O_2099,N_24318,N_24616);
and UO_2100 (O_2100,N_23720,N_23903);
or UO_2101 (O_2101,N_24489,N_24427);
and UO_2102 (O_2102,N_23468,N_23850);
and UO_2103 (O_2103,N_22821,N_24702);
nor UO_2104 (O_2104,N_22282,N_23904);
nor UO_2105 (O_2105,N_21961,N_22099);
and UO_2106 (O_2106,N_24327,N_21964);
nor UO_2107 (O_2107,N_24139,N_22247);
and UO_2108 (O_2108,N_24711,N_22961);
nor UO_2109 (O_2109,N_22087,N_24365);
xnor UO_2110 (O_2110,N_23870,N_21989);
nor UO_2111 (O_2111,N_22283,N_22829);
or UO_2112 (O_2112,N_24581,N_23410);
or UO_2113 (O_2113,N_23948,N_22017);
nand UO_2114 (O_2114,N_22026,N_23439);
or UO_2115 (O_2115,N_24883,N_23975);
nor UO_2116 (O_2116,N_22895,N_23845);
and UO_2117 (O_2117,N_22871,N_22127);
or UO_2118 (O_2118,N_24953,N_23989);
and UO_2119 (O_2119,N_22176,N_23534);
xnor UO_2120 (O_2120,N_22814,N_23278);
xor UO_2121 (O_2121,N_24741,N_22397);
or UO_2122 (O_2122,N_22169,N_22281);
or UO_2123 (O_2123,N_23066,N_24743);
and UO_2124 (O_2124,N_23633,N_22842);
xor UO_2125 (O_2125,N_24452,N_22661);
or UO_2126 (O_2126,N_23667,N_22460);
nor UO_2127 (O_2127,N_22246,N_21990);
nand UO_2128 (O_2128,N_23290,N_23440);
or UO_2129 (O_2129,N_22100,N_22073);
nor UO_2130 (O_2130,N_22957,N_24003);
nor UO_2131 (O_2131,N_23706,N_23443);
and UO_2132 (O_2132,N_22475,N_24196);
or UO_2133 (O_2133,N_24709,N_23638);
and UO_2134 (O_2134,N_24988,N_22532);
and UO_2135 (O_2135,N_22775,N_22705);
and UO_2136 (O_2136,N_22513,N_24060);
xnor UO_2137 (O_2137,N_22522,N_23893);
nand UO_2138 (O_2138,N_23063,N_23709);
nand UO_2139 (O_2139,N_24031,N_23861);
nand UO_2140 (O_2140,N_22641,N_24779);
or UO_2141 (O_2141,N_23864,N_24378);
and UO_2142 (O_2142,N_23043,N_24676);
or UO_2143 (O_2143,N_22591,N_23625);
or UO_2144 (O_2144,N_22790,N_23425);
and UO_2145 (O_2145,N_22466,N_22801);
xnor UO_2146 (O_2146,N_22444,N_24870);
and UO_2147 (O_2147,N_24138,N_23511);
nor UO_2148 (O_2148,N_23237,N_24784);
xnor UO_2149 (O_2149,N_22406,N_24845);
and UO_2150 (O_2150,N_23752,N_22645);
nand UO_2151 (O_2151,N_22614,N_23606);
nand UO_2152 (O_2152,N_23563,N_22807);
nand UO_2153 (O_2153,N_23919,N_24013);
xor UO_2154 (O_2154,N_24229,N_23535);
nor UO_2155 (O_2155,N_23915,N_22071);
xor UO_2156 (O_2156,N_24408,N_24474);
nor UO_2157 (O_2157,N_24028,N_22285);
nor UO_2158 (O_2158,N_24367,N_24157);
nand UO_2159 (O_2159,N_24806,N_23963);
and UO_2160 (O_2160,N_23517,N_24581);
nor UO_2161 (O_2161,N_23332,N_22022);
and UO_2162 (O_2162,N_22940,N_24547);
nor UO_2163 (O_2163,N_23625,N_24190);
xnor UO_2164 (O_2164,N_24808,N_24627);
nor UO_2165 (O_2165,N_24928,N_22311);
or UO_2166 (O_2166,N_24763,N_23066);
nand UO_2167 (O_2167,N_22277,N_22571);
or UO_2168 (O_2168,N_24758,N_23221);
nor UO_2169 (O_2169,N_22738,N_23866);
xor UO_2170 (O_2170,N_22096,N_22166);
or UO_2171 (O_2171,N_22905,N_22107);
and UO_2172 (O_2172,N_22876,N_23753);
nand UO_2173 (O_2173,N_24494,N_23030);
or UO_2174 (O_2174,N_24047,N_22528);
and UO_2175 (O_2175,N_22593,N_23980);
nand UO_2176 (O_2176,N_24716,N_23866);
or UO_2177 (O_2177,N_22689,N_22017);
and UO_2178 (O_2178,N_24609,N_23614);
xnor UO_2179 (O_2179,N_24665,N_23445);
or UO_2180 (O_2180,N_24509,N_24263);
nor UO_2181 (O_2181,N_24281,N_23844);
nand UO_2182 (O_2182,N_23677,N_22136);
nand UO_2183 (O_2183,N_23866,N_24495);
nor UO_2184 (O_2184,N_22341,N_21907);
or UO_2185 (O_2185,N_22601,N_23536);
nand UO_2186 (O_2186,N_22731,N_24463);
and UO_2187 (O_2187,N_24092,N_22104);
or UO_2188 (O_2188,N_24605,N_22523);
nor UO_2189 (O_2189,N_23127,N_22128);
nand UO_2190 (O_2190,N_23210,N_24020);
or UO_2191 (O_2191,N_21975,N_22434);
or UO_2192 (O_2192,N_23821,N_24625);
or UO_2193 (O_2193,N_22551,N_23108);
nand UO_2194 (O_2194,N_23575,N_24143);
nand UO_2195 (O_2195,N_24221,N_23928);
xnor UO_2196 (O_2196,N_22611,N_23413);
nand UO_2197 (O_2197,N_22051,N_24611);
and UO_2198 (O_2198,N_23936,N_24433);
xnor UO_2199 (O_2199,N_24862,N_23101);
nand UO_2200 (O_2200,N_23360,N_22882);
nand UO_2201 (O_2201,N_23907,N_22552);
and UO_2202 (O_2202,N_24296,N_22536);
and UO_2203 (O_2203,N_23770,N_24493);
and UO_2204 (O_2204,N_24446,N_23795);
nor UO_2205 (O_2205,N_22685,N_23364);
nand UO_2206 (O_2206,N_22440,N_22656);
nand UO_2207 (O_2207,N_23635,N_23856);
nor UO_2208 (O_2208,N_22892,N_24839);
or UO_2209 (O_2209,N_24586,N_22094);
or UO_2210 (O_2210,N_24495,N_23528);
nor UO_2211 (O_2211,N_21939,N_24270);
and UO_2212 (O_2212,N_24153,N_24826);
or UO_2213 (O_2213,N_22923,N_23984);
or UO_2214 (O_2214,N_24960,N_22198);
and UO_2215 (O_2215,N_23190,N_22275);
nand UO_2216 (O_2216,N_23291,N_22227);
nor UO_2217 (O_2217,N_21930,N_22083);
or UO_2218 (O_2218,N_22172,N_24443);
nor UO_2219 (O_2219,N_22668,N_23359);
xnor UO_2220 (O_2220,N_23336,N_22640);
xor UO_2221 (O_2221,N_22871,N_22152);
nand UO_2222 (O_2222,N_24257,N_22992);
nor UO_2223 (O_2223,N_21984,N_24835);
or UO_2224 (O_2224,N_22799,N_23834);
nand UO_2225 (O_2225,N_24106,N_22640);
or UO_2226 (O_2226,N_22008,N_24751);
or UO_2227 (O_2227,N_24879,N_23294);
nor UO_2228 (O_2228,N_22889,N_23299);
xor UO_2229 (O_2229,N_24202,N_23929);
nand UO_2230 (O_2230,N_22670,N_23460);
nand UO_2231 (O_2231,N_24069,N_24344);
or UO_2232 (O_2232,N_21914,N_24769);
and UO_2233 (O_2233,N_21913,N_23770);
or UO_2234 (O_2234,N_22785,N_22327);
or UO_2235 (O_2235,N_22800,N_22055);
nor UO_2236 (O_2236,N_23130,N_23440);
nor UO_2237 (O_2237,N_24046,N_24538);
or UO_2238 (O_2238,N_22656,N_24048);
xor UO_2239 (O_2239,N_24432,N_22049);
and UO_2240 (O_2240,N_24443,N_22532);
or UO_2241 (O_2241,N_23067,N_22472);
nor UO_2242 (O_2242,N_22868,N_23713);
and UO_2243 (O_2243,N_24826,N_23736);
nor UO_2244 (O_2244,N_22422,N_24920);
nand UO_2245 (O_2245,N_22758,N_22105);
and UO_2246 (O_2246,N_22808,N_24221);
or UO_2247 (O_2247,N_24030,N_23257);
nand UO_2248 (O_2248,N_24519,N_24069);
or UO_2249 (O_2249,N_22825,N_22183);
nand UO_2250 (O_2250,N_23782,N_24794);
and UO_2251 (O_2251,N_24966,N_22773);
xor UO_2252 (O_2252,N_22521,N_23566);
nand UO_2253 (O_2253,N_24206,N_23827);
nand UO_2254 (O_2254,N_23342,N_24196);
and UO_2255 (O_2255,N_24207,N_22192);
and UO_2256 (O_2256,N_23739,N_24408);
nand UO_2257 (O_2257,N_24925,N_24367);
and UO_2258 (O_2258,N_24628,N_22431);
or UO_2259 (O_2259,N_24415,N_22914);
or UO_2260 (O_2260,N_21997,N_24022);
nand UO_2261 (O_2261,N_24688,N_22888);
nand UO_2262 (O_2262,N_23491,N_22686);
nor UO_2263 (O_2263,N_22874,N_24660);
or UO_2264 (O_2264,N_24322,N_22007);
or UO_2265 (O_2265,N_23846,N_22835);
and UO_2266 (O_2266,N_24578,N_23016);
nand UO_2267 (O_2267,N_22706,N_23734);
or UO_2268 (O_2268,N_22169,N_22929);
and UO_2269 (O_2269,N_22209,N_22268);
nand UO_2270 (O_2270,N_24795,N_23508);
nand UO_2271 (O_2271,N_24769,N_23167);
or UO_2272 (O_2272,N_22341,N_22600);
or UO_2273 (O_2273,N_23590,N_23379);
or UO_2274 (O_2274,N_24161,N_21900);
or UO_2275 (O_2275,N_23703,N_23449);
nor UO_2276 (O_2276,N_24118,N_23824);
nor UO_2277 (O_2277,N_22348,N_22693);
nor UO_2278 (O_2278,N_24279,N_22550);
or UO_2279 (O_2279,N_23492,N_23230);
nand UO_2280 (O_2280,N_24929,N_24336);
or UO_2281 (O_2281,N_22198,N_22219);
nand UO_2282 (O_2282,N_24481,N_22007);
and UO_2283 (O_2283,N_22746,N_22903);
nand UO_2284 (O_2284,N_24763,N_23996);
or UO_2285 (O_2285,N_22185,N_24736);
nor UO_2286 (O_2286,N_22600,N_21943);
nor UO_2287 (O_2287,N_23471,N_22738);
nand UO_2288 (O_2288,N_24723,N_23438);
or UO_2289 (O_2289,N_22441,N_22737);
nand UO_2290 (O_2290,N_24495,N_23651);
nor UO_2291 (O_2291,N_23179,N_23552);
nor UO_2292 (O_2292,N_22235,N_22386);
nand UO_2293 (O_2293,N_22264,N_24778);
nor UO_2294 (O_2294,N_24546,N_22663);
or UO_2295 (O_2295,N_21934,N_24777);
and UO_2296 (O_2296,N_24805,N_24746);
nor UO_2297 (O_2297,N_22470,N_22960);
nand UO_2298 (O_2298,N_23574,N_23193);
xor UO_2299 (O_2299,N_23569,N_24769);
or UO_2300 (O_2300,N_22072,N_23436);
nand UO_2301 (O_2301,N_24269,N_24934);
nand UO_2302 (O_2302,N_23627,N_24175);
nand UO_2303 (O_2303,N_24703,N_22936);
and UO_2304 (O_2304,N_22675,N_23633);
nand UO_2305 (O_2305,N_24778,N_22902);
or UO_2306 (O_2306,N_24437,N_24215);
nand UO_2307 (O_2307,N_24687,N_23065);
nand UO_2308 (O_2308,N_22117,N_24755);
and UO_2309 (O_2309,N_22570,N_22178);
or UO_2310 (O_2310,N_23832,N_22953);
xnor UO_2311 (O_2311,N_24575,N_24337);
nand UO_2312 (O_2312,N_23725,N_23068);
or UO_2313 (O_2313,N_23879,N_24306);
and UO_2314 (O_2314,N_23013,N_22234);
nor UO_2315 (O_2315,N_22257,N_23782);
or UO_2316 (O_2316,N_22031,N_22099);
or UO_2317 (O_2317,N_22959,N_23494);
and UO_2318 (O_2318,N_24975,N_23765);
or UO_2319 (O_2319,N_24465,N_24128);
nor UO_2320 (O_2320,N_22770,N_24362);
nor UO_2321 (O_2321,N_24765,N_22492);
nor UO_2322 (O_2322,N_23589,N_22978);
and UO_2323 (O_2323,N_23101,N_22000);
nor UO_2324 (O_2324,N_23034,N_22938);
nor UO_2325 (O_2325,N_23516,N_23411);
and UO_2326 (O_2326,N_24010,N_22560);
or UO_2327 (O_2327,N_22130,N_22600);
and UO_2328 (O_2328,N_24088,N_23931);
nor UO_2329 (O_2329,N_22892,N_22189);
and UO_2330 (O_2330,N_22317,N_21943);
and UO_2331 (O_2331,N_22651,N_23997);
or UO_2332 (O_2332,N_24260,N_24683);
and UO_2333 (O_2333,N_22559,N_23752);
nand UO_2334 (O_2334,N_22056,N_23438);
nor UO_2335 (O_2335,N_24289,N_24966);
nor UO_2336 (O_2336,N_22120,N_23568);
or UO_2337 (O_2337,N_23542,N_23165);
nor UO_2338 (O_2338,N_22931,N_22129);
nor UO_2339 (O_2339,N_22795,N_22878);
or UO_2340 (O_2340,N_22921,N_24792);
and UO_2341 (O_2341,N_23091,N_24365);
and UO_2342 (O_2342,N_23553,N_24854);
or UO_2343 (O_2343,N_24901,N_24133);
and UO_2344 (O_2344,N_24323,N_24843);
nor UO_2345 (O_2345,N_24879,N_23652);
nand UO_2346 (O_2346,N_23030,N_24652);
nor UO_2347 (O_2347,N_22718,N_22671);
xnor UO_2348 (O_2348,N_24265,N_22355);
nor UO_2349 (O_2349,N_22019,N_24165);
nor UO_2350 (O_2350,N_22115,N_22255);
and UO_2351 (O_2351,N_24945,N_23585);
xor UO_2352 (O_2352,N_22560,N_24826);
xor UO_2353 (O_2353,N_23870,N_24039);
and UO_2354 (O_2354,N_22553,N_24398);
or UO_2355 (O_2355,N_23853,N_23199);
and UO_2356 (O_2356,N_22087,N_22531);
nand UO_2357 (O_2357,N_23125,N_24797);
or UO_2358 (O_2358,N_24765,N_23077);
nand UO_2359 (O_2359,N_24662,N_23177);
nor UO_2360 (O_2360,N_24500,N_24049);
nand UO_2361 (O_2361,N_23799,N_24663);
nand UO_2362 (O_2362,N_24572,N_22982);
nand UO_2363 (O_2363,N_22965,N_22916);
or UO_2364 (O_2364,N_24677,N_24900);
nand UO_2365 (O_2365,N_24049,N_21904);
nor UO_2366 (O_2366,N_23779,N_22232);
nor UO_2367 (O_2367,N_22155,N_23300);
and UO_2368 (O_2368,N_23595,N_24659);
xor UO_2369 (O_2369,N_24030,N_24256);
xor UO_2370 (O_2370,N_24252,N_22557);
nand UO_2371 (O_2371,N_24458,N_22968);
xnor UO_2372 (O_2372,N_23846,N_24671);
and UO_2373 (O_2373,N_23477,N_23670);
and UO_2374 (O_2374,N_23481,N_24430);
nor UO_2375 (O_2375,N_22163,N_22177);
and UO_2376 (O_2376,N_22970,N_24198);
and UO_2377 (O_2377,N_24229,N_23524);
nor UO_2378 (O_2378,N_22893,N_22706);
and UO_2379 (O_2379,N_24044,N_24024);
nand UO_2380 (O_2380,N_22008,N_24816);
nor UO_2381 (O_2381,N_22698,N_22243);
and UO_2382 (O_2382,N_22170,N_24909);
or UO_2383 (O_2383,N_23032,N_21896);
or UO_2384 (O_2384,N_22327,N_24056);
xnor UO_2385 (O_2385,N_22929,N_24697);
nand UO_2386 (O_2386,N_24672,N_23519);
nand UO_2387 (O_2387,N_23458,N_22200);
nand UO_2388 (O_2388,N_23293,N_24748);
nor UO_2389 (O_2389,N_24051,N_22147);
or UO_2390 (O_2390,N_22148,N_24258);
and UO_2391 (O_2391,N_22825,N_24008);
nor UO_2392 (O_2392,N_21890,N_22893);
and UO_2393 (O_2393,N_22965,N_22730);
or UO_2394 (O_2394,N_22933,N_23175);
and UO_2395 (O_2395,N_23544,N_23795);
nor UO_2396 (O_2396,N_22097,N_24230);
and UO_2397 (O_2397,N_23356,N_24130);
nand UO_2398 (O_2398,N_22375,N_23319);
nor UO_2399 (O_2399,N_24746,N_23242);
and UO_2400 (O_2400,N_22567,N_23295);
or UO_2401 (O_2401,N_23619,N_22722);
nand UO_2402 (O_2402,N_23576,N_22297);
xor UO_2403 (O_2403,N_23579,N_23412);
and UO_2404 (O_2404,N_24901,N_24985);
xor UO_2405 (O_2405,N_24639,N_22096);
nor UO_2406 (O_2406,N_24842,N_22433);
or UO_2407 (O_2407,N_24047,N_24454);
nand UO_2408 (O_2408,N_23684,N_24375);
or UO_2409 (O_2409,N_22815,N_24812);
or UO_2410 (O_2410,N_22049,N_22042);
and UO_2411 (O_2411,N_23838,N_21922);
and UO_2412 (O_2412,N_24655,N_23471);
and UO_2413 (O_2413,N_22769,N_24241);
nor UO_2414 (O_2414,N_23882,N_24611);
nor UO_2415 (O_2415,N_21908,N_23900);
xnor UO_2416 (O_2416,N_24088,N_24710);
xor UO_2417 (O_2417,N_24337,N_22628);
and UO_2418 (O_2418,N_24663,N_22732);
xnor UO_2419 (O_2419,N_23757,N_23554);
and UO_2420 (O_2420,N_24264,N_24737);
nor UO_2421 (O_2421,N_23245,N_24989);
nand UO_2422 (O_2422,N_24529,N_22795);
or UO_2423 (O_2423,N_24946,N_22578);
and UO_2424 (O_2424,N_24386,N_21976);
nor UO_2425 (O_2425,N_22755,N_22095);
nand UO_2426 (O_2426,N_24831,N_22553);
or UO_2427 (O_2427,N_23648,N_23375);
xnor UO_2428 (O_2428,N_23230,N_22692);
nand UO_2429 (O_2429,N_24635,N_24993);
xnor UO_2430 (O_2430,N_24729,N_24636);
xor UO_2431 (O_2431,N_22541,N_24401);
nor UO_2432 (O_2432,N_22534,N_22459);
and UO_2433 (O_2433,N_24967,N_23988);
or UO_2434 (O_2434,N_23102,N_23468);
nor UO_2435 (O_2435,N_23687,N_22477);
xor UO_2436 (O_2436,N_24349,N_24314);
nand UO_2437 (O_2437,N_24982,N_22029);
or UO_2438 (O_2438,N_22726,N_24280);
or UO_2439 (O_2439,N_22418,N_22859);
nand UO_2440 (O_2440,N_22270,N_24989);
and UO_2441 (O_2441,N_24454,N_23404);
or UO_2442 (O_2442,N_22394,N_22211);
nor UO_2443 (O_2443,N_24571,N_22724);
nand UO_2444 (O_2444,N_23847,N_23695);
and UO_2445 (O_2445,N_23136,N_23853);
or UO_2446 (O_2446,N_22703,N_22184);
nand UO_2447 (O_2447,N_24919,N_23381);
nor UO_2448 (O_2448,N_22292,N_23914);
or UO_2449 (O_2449,N_22379,N_24470);
and UO_2450 (O_2450,N_22960,N_22600);
or UO_2451 (O_2451,N_23428,N_23673);
xnor UO_2452 (O_2452,N_23063,N_23611);
xor UO_2453 (O_2453,N_23656,N_24564);
or UO_2454 (O_2454,N_23558,N_22988);
xor UO_2455 (O_2455,N_22920,N_23245);
or UO_2456 (O_2456,N_24624,N_21903);
and UO_2457 (O_2457,N_23652,N_23824);
and UO_2458 (O_2458,N_23857,N_22311);
xor UO_2459 (O_2459,N_24592,N_23267);
nor UO_2460 (O_2460,N_22736,N_22734);
nor UO_2461 (O_2461,N_24021,N_22786);
nand UO_2462 (O_2462,N_24967,N_24101);
or UO_2463 (O_2463,N_23875,N_22839);
nor UO_2464 (O_2464,N_24359,N_23508);
nor UO_2465 (O_2465,N_23539,N_22988);
and UO_2466 (O_2466,N_24882,N_22175);
or UO_2467 (O_2467,N_22916,N_22544);
and UO_2468 (O_2468,N_24068,N_23698);
nand UO_2469 (O_2469,N_24888,N_23455);
nor UO_2470 (O_2470,N_24238,N_21887);
xnor UO_2471 (O_2471,N_22210,N_24427);
or UO_2472 (O_2472,N_23746,N_23389);
and UO_2473 (O_2473,N_24198,N_22628);
xor UO_2474 (O_2474,N_24088,N_22619);
nand UO_2475 (O_2475,N_22788,N_24537);
nand UO_2476 (O_2476,N_24429,N_24230);
and UO_2477 (O_2477,N_22336,N_24238);
and UO_2478 (O_2478,N_24248,N_23119);
nand UO_2479 (O_2479,N_23477,N_23656);
nand UO_2480 (O_2480,N_24738,N_23376);
nor UO_2481 (O_2481,N_23422,N_24110);
and UO_2482 (O_2482,N_22244,N_24395);
nand UO_2483 (O_2483,N_22108,N_24659);
nor UO_2484 (O_2484,N_22318,N_24881);
and UO_2485 (O_2485,N_24273,N_24793);
nand UO_2486 (O_2486,N_23196,N_24546);
nor UO_2487 (O_2487,N_21984,N_22860);
and UO_2488 (O_2488,N_23492,N_22111);
xnor UO_2489 (O_2489,N_24657,N_23013);
or UO_2490 (O_2490,N_21876,N_22489);
and UO_2491 (O_2491,N_24103,N_23432);
nand UO_2492 (O_2492,N_23552,N_23523);
or UO_2493 (O_2493,N_22313,N_22114);
nor UO_2494 (O_2494,N_24971,N_24021);
and UO_2495 (O_2495,N_22261,N_24369);
xnor UO_2496 (O_2496,N_23892,N_23725);
nand UO_2497 (O_2497,N_24075,N_22277);
nor UO_2498 (O_2498,N_24281,N_24430);
xnor UO_2499 (O_2499,N_22998,N_23337);
nor UO_2500 (O_2500,N_23215,N_23514);
nor UO_2501 (O_2501,N_23978,N_22000);
or UO_2502 (O_2502,N_23581,N_24064);
or UO_2503 (O_2503,N_22824,N_22390);
and UO_2504 (O_2504,N_24449,N_24060);
or UO_2505 (O_2505,N_24386,N_22718);
nor UO_2506 (O_2506,N_24869,N_22859);
and UO_2507 (O_2507,N_24366,N_24149);
nor UO_2508 (O_2508,N_24775,N_23064);
nand UO_2509 (O_2509,N_24161,N_22550);
and UO_2510 (O_2510,N_23569,N_22702);
and UO_2511 (O_2511,N_22862,N_22680);
nand UO_2512 (O_2512,N_24529,N_22255);
nand UO_2513 (O_2513,N_23637,N_23026);
nand UO_2514 (O_2514,N_22467,N_24050);
or UO_2515 (O_2515,N_24525,N_23467);
nor UO_2516 (O_2516,N_24315,N_23257);
and UO_2517 (O_2517,N_23575,N_22932);
nand UO_2518 (O_2518,N_23279,N_24002);
nand UO_2519 (O_2519,N_23158,N_24227);
or UO_2520 (O_2520,N_23072,N_24314);
or UO_2521 (O_2521,N_22040,N_23898);
and UO_2522 (O_2522,N_22082,N_22114);
or UO_2523 (O_2523,N_22295,N_24355);
and UO_2524 (O_2524,N_24260,N_23232);
or UO_2525 (O_2525,N_24097,N_22617);
nor UO_2526 (O_2526,N_22785,N_24193);
nor UO_2527 (O_2527,N_21918,N_22945);
xor UO_2528 (O_2528,N_23503,N_24054);
nor UO_2529 (O_2529,N_22962,N_23254);
and UO_2530 (O_2530,N_23652,N_24832);
nor UO_2531 (O_2531,N_23173,N_24844);
or UO_2532 (O_2532,N_24616,N_22178);
nor UO_2533 (O_2533,N_24833,N_24258);
and UO_2534 (O_2534,N_22413,N_22927);
nor UO_2535 (O_2535,N_24387,N_23906);
nor UO_2536 (O_2536,N_23822,N_21885);
nor UO_2537 (O_2537,N_24606,N_24304);
xor UO_2538 (O_2538,N_23447,N_23311);
nand UO_2539 (O_2539,N_24237,N_24185);
nand UO_2540 (O_2540,N_24963,N_23861);
nor UO_2541 (O_2541,N_22029,N_24436);
nor UO_2542 (O_2542,N_22987,N_24951);
and UO_2543 (O_2543,N_23909,N_22370);
or UO_2544 (O_2544,N_22238,N_22260);
xnor UO_2545 (O_2545,N_23669,N_23871);
nand UO_2546 (O_2546,N_24430,N_22093);
nand UO_2547 (O_2547,N_24892,N_24429);
and UO_2548 (O_2548,N_24600,N_23688);
or UO_2549 (O_2549,N_21975,N_22645);
or UO_2550 (O_2550,N_21909,N_24036);
nor UO_2551 (O_2551,N_24971,N_23557);
and UO_2552 (O_2552,N_22247,N_24924);
xnor UO_2553 (O_2553,N_22511,N_22960);
nand UO_2554 (O_2554,N_22856,N_24488);
nor UO_2555 (O_2555,N_22695,N_23605);
nor UO_2556 (O_2556,N_24098,N_23773);
and UO_2557 (O_2557,N_22781,N_23531);
or UO_2558 (O_2558,N_22520,N_22885);
nor UO_2559 (O_2559,N_22929,N_24031);
nor UO_2560 (O_2560,N_24254,N_23649);
nor UO_2561 (O_2561,N_21908,N_22731);
or UO_2562 (O_2562,N_22141,N_23011);
or UO_2563 (O_2563,N_24051,N_23110);
or UO_2564 (O_2564,N_24608,N_22718);
or UO_2565 (O_2565,N_23786,N_22833);
nor UO_2566 (O_2566,N_23996,N_23162);
or UO_2567 (O_2567,N_24480,N_23908);
nand UO_2568 (O_2568,N_24426,N_22891);
and UO_2569 (O_2569,N_23386,N_23857);
xor UO_2570 (O_2570,N_23000,N_21956);
and UO_2571 (O_2571,N_23343,N_23037);
or UO_2572 (O_2572,N_22693,N_22248);
xnor UO_2573 (O_2573,N_24718,N_23497);
or UO_2574 (O_2574,N_24725,N_23281);
nand UO_2575 (O_2575,N_22262,N_22103);
or UO_2576 (O_2576,N_23877,N_24189);
nor UO_2577 (O_2577,N_24308,N_22968);
and UO_2578 (O_2578,N_24321,N_22046);
nand UO_2579 (O_2579,N_23204,N_24562);
or UO_2580 (O_2580,N_22966,N_22250);
nand UO_2581 (O_2581,N_22169,N_24606);
or UO_2582 (O_2582,N_23814,N_24286);
nor UO_2583 (O_2583,N_22005,N_24344);
and UO_2584 (O_2584,N_24136,N_23032);
nor UO_2585 (O_2585,N_22242,N_22756);
nand UO_2586 (O_2586,N_24481,N_21926);
and UO_2587 (O_2587,N_23565,N_23189);
and UO_2588 (O_2588,N_23944,N_22223);
or UO_2589 (O_2589,N_24097,N_22735);
nor UO_2590 (O_2590,N_22895,N_22209);
nand UO_2591 (O_2591,N_22476,N_23029);
nor UO_2592 (O_2592,N_24722,N_21937);
nor UO_2593 (O_2593,N_23859,N_24185);
nor UO_2594 (O_2594,N_23339,N_22909);
nor UO_2595 (O_2595,N_23719,N_22934);
and UO_2596 (O_2596,N_22657,N_22302);
or UO_2597 (O_2597,N_23093,N_22373);
and UO_2598 (O_2598,N_23313,N_22898);
or UO_2599 (O_2599,N_24039,N_22262);
or UO_2600 (O_2600,N_24970,N_23795);
and UO_2601 (O_2601,N_22323,N_24057);
or UO_2602 (O_2602,N_23852,N_24676);
nor UO_2603 (O_2603,N_24755,N_24154);
nor UO_2604 (O_2604,N_22513,N_24986);
and UO_2605 (O_2605,N_24198,N_24272);
or UO_2606 (O_2606,N_22229,N_24066);
or UO_2607 (O_2607,N_22337,N_24536);
and UO_2608 (O_2608,N_24766,N_23367);
nand UO_2609 (O_2609,N_24491,N_22943);
nand UO_2610 (O_2610,N_24827,N_24791);
and UO_2611 (O_2611,N_23989,N_23653);
xnor UO_2612 (O_2612,N_23748,N_23186);
nor UO_2613 (O_2613,N_24999,N_21889);
nor UO_2614 (O_2614,N_22518,N_22055);
or UO_2615 (O_2615,N_23623,N_24987);
nor UO_2616 (O_2616,N_24726,N_22411);
nand UO_2617 (O_2617,N_23521,N_23674);
nor UO_2618 (O_2618,N_24012,N_22767);
nand UO_2619 (O_2619,N_23847,N_22312);
nor UO_2620 (O_2620,N_22232,N_24781);
and UO_2621 (O_2621,N_23065,N_22695);
or UO_2622 (O_2622,N_22827,N_22435);
nand UO_2623 (O_2623,N_23563,N_24925);
and UO_2624 (O_2624,N_22899,N_24555);
nor UO_2625 (O_2625,N_24730,N_22664);
nand UO_2626 (O_2626,N_23502,N_24858);
nor UO_2627 (O_2627,N_22958,N_23959);
and UO_2628 (O_2628,N_23879,N_22366);
or UO_2629 (O_2629,N_24149,N_22850);
nand UO_2630 (O_2630,N_23823,N_24177);
nand UO_2631 (O_2631,N_21906,N_22157);
or UO_2632 (O_2632,N_23873,N_23369);
and UO_2633 (O_2633,N_24431,N_23043);
and UO_2634 (O_2634,N_24686,N_24543);
nor UO_2635 (O_2635,N_22098,N_22687);
and UO_2636 (O_2636,N_24201,N_22455);
and UO_2637 (O_2637,N_22493,N_24844);
or UO_2638 (O_2638,N_22582,N_22475);
or UO_2639 (O_2639,N_22843,N_23608);
and UO_2640 (O_2640,N_24492,N_22395);
or UO_2641 (O_2641,N_23673,N_22611);
nand UO_2642 (O_2642,N_22172,N_23515);
and UO_2643 (O_2643,N_22715,N_23421);
nor UO_2644 (O_2644,N_23665,N_24618);
and UO_2645 (O_2645,N_23947,N_24505);
or UO_2646 (O_2646,N_23404,N_21922);
and UO_2647 (O_2647,N_24602,N_24735);
nand UO_2648 (O_2648,N_24106,N_23535);
or UO_2649 (O_2649,N_23786,N_24486);
or UO_2650 (O_2650,N_22191,N_22415);
or UO_2651 (O_2651,N_23109,N_22128);
nand UO_2652 (O_2652,N_22391,N_23094);
or UO_2653 (O_2653,N_22787,N_22607);
nand UO_2654 (O_2654,N_21951,N_23694);
xnor UO_2655 (O_2655,N_24198,N_23104);
nor UO_2656 (O_2656,N_21961,N_24919);
and UO_2657 (O_2657,N_23760,N_22635);
or UO_2658 (O_2658,N_24793,N_23379);
nand UO_2659 (O_2659,N_24888,N_21902);
and UO_2660 (O_2660,N_24749,N_22469);
nor UO_2661 (O_2661,N_23659,N_22374);
nor UO_2662 (O_2662,N_24214,N_23291);
nor UO_2663 (O_2663,N_23123,N_24588);
or UO_2664 (O_2664,N_22829,N_23381);
nor UO_2665 (O_2665,N_24718,N_22921);
and UO_2666 (O_2666,N_23790,N_22220);
or UO_2667 (O_2667,N_24898,N_22239);
nand UO_2668 (O_2668,N_24889,N_24055);
or UO_2669 (O_2669,N_23666,N_24859);
nand UO_2670 (O_2670,N_23009,N_23168);
nor UO_2671 (O_2671,N_24587,N_22245);
and UO_2672 (O_2672,N_22407,N_23947);
nor UO_2673 (O_2673,N_23011,N_22337);
nand UO_2674 (O_2674,N_23609,N_23198);
nor UO_2675 (O_2675,N_24033,N_22388);
and UO_2676 (O_2676,N_24974,N_24734);
and UO_2677 (O_2677,N_24271,N_22341);
xnor UO_2678 (O_2678,N_24684,N_23400);
or UO_2679 (O_2679,N_22230,N_24305);
nor UO_2680 (O_2680,N_24148,N_24520);
nor UO_2681 (O_2681,N_23313,N_24455);
nand UO_2682 (O_2682,N_23917,N_21878);
and UO_2683 (O_2683,N_23956,N_22337);
or UO_2684 (O_2684,N_23658,N_23907);
xnor UO_2685 (O_2685,N_22481,N_23653);
nand UO_2686 (O_2686,N_23644,N_22193);
nand UO_2687 (O_2687,N_24732,N_21982);
and UO_2688 (O_2688,N_23824,N_23655);
and UO_2689 (O_2689,N_22311,N_22974);
nor UO_2690 (O_2690,N_23852,N_22901);
and UO_2691 (O_2691,N_22656,N_23576);
nor UO_2692 (O_2692,N_22447,N_22786);
xor UO_2693 (O_2693,N_22583,N_21902);
and UO_2694 (O_2694,N_22725,N_24869);
xnor UO_2695 (O_2695,N_24799,N_23150);
nor UO_2696 (O_2696,N_22232,N_22558);
and UO_2697 (O_2697,N_23202,N_23432);
nand UO_2698 (O_2698,N_24599,N_23587);
nand UO_2699 (O_2699,N_22615,N_23696);
or UO_2700 (O_2700,N_24583,N_24733);
and UO_2701 (O_2701,N_22544,N_24533);
nand UO_2702 (O_2702,N_22927,N_23070);
nor UO_2703 (O_2703,N_24175,N_22466);
nor UO_2704 (O_2704,N_24193,N_24997);
and UO_2705 (O_2705,N_22818,N_23026);
nor UO_2706 (O_2706,N_23442,N_23107);
and UO_2707 (O_2707,N_22105,N_24751);
nor UO_2708 (O_2708,N_23727,N_23877);
nand UO_2709 (O_2709,N_23461,N_22305);
nor UO_2710 (O_2710,N_23321,N_22862);
and UO_2711 (O_2711,N_22732,N_23128);
or UO_2712 (O_2712,N_24853,N_24280);
and UO_2713 (O_2713,N_23809,N_24075);
nand UO_2714 (O_2714,N_24558,N_23307);
or UO_2715 (O_2715,N_24840,N_23253);
nor UO_2716 (O_2716,N_24556,N_22266);
or UO_2717 (O_2717,N_23456,N_23473);
or UO_2718 (O_2718,N_22287,N_22555);
nand UO_2719 (O_2719,N_22432,N_24802);
nor UO_2720 (O_2720,N_23053,N_22379);
nor UO_2721 (O_2721,N_23292,N_22550);
and UO_2722 (O_2722,N_23226,N_21943);
nand UO_2723 (O_2723,N_23848,N_23530);
or UO_2724 (O_2724,N_22575,N_22639);
nand UO_2725 (O_2725,N_24046,N_23169);
and UO_2726 (O_2726,N_24356,N_24930);
and UO_2727 (O_2727,N_23070,N_23308);
nand UO_2728 (O_2728,N_24125,N_24075);
or UO_2729 (O_2729,N_21917,N_24983);
nand UO_2730 (O_2730,N_23853,N_24653);
or UO_2731 (O_2731,N_23795,N_23752);
or UO_2732 (O_2732,N_22499,N_23223);
xnor UO_2733 (O_2733,N_24446,N_24675);
nand UO_2734 (O_2734,N_21964,N_22844);
xnor UO_2735 (O_2735,N_22423,N_24408);
nand UO_2736 (O_2736,N_23021,N_22039);
xnor UO_2737 (O_2737,N_23543,N_24904);
nand UO_2738 (O_2738,N_24530,N_22324);
nand UO_2739 (O_2739,N_23484,N_23122);
nand UO_2740 (O_2740,N_24717,N_22107);
or UO_2741 (O_2741,N_23723,N_24501);
or UO_2742 (O_2742,N_22556,N_24856);
nor UO_2743 (O_2743,N_24117,N_22574);
or UO_2744 (O_2744,N_22888,N_22654);
nand UO_2745 (O_2745,N_23816,N_24387);
and UO_2746 (O_2746,N_24580,N_22245);
nand UO_2747 (O_2747,N_23696,N_24241);
nor UO_2748 (O_2748,N_24990,N_22323);
or UO_2749 (O_2749,N_24246,N_23588);
nand UO_2750 (O_2750,N_22090,N_24863);
or UO_2751 (O_2751,N_23589,N_22876);
nand UO_2752 (O_2752,N_22876,N_22532);
or UO_2753 (O_2753,N_23965,N_23336);
or UO_2754 (O_2754,N_24746,N_22901);
nand UO_2755 (O_2755,N_21971,N_22444);
and UO_2756 (O_2756,N_22351,N_22625);
nor UO_2757 (O_2757,N_24256,N_22581);
xnor UO_2758 (O_2758,N_24043,N_22404);
or UO_2759 (O_2759,N_23315,N_23314);
nor UO_2760 (O_2760,N_23711,N_24538);
and UO_2761 (O_2761,N_22761,N_22287);
nand UO_2762 (O_2762,N_22712,N_21997);
and UO_2763 (O_2763,N_24145,N_24060);
nor UO_2764 (O_2764,N_22890,N_24125);
or UO_2765 (O_2765,N_22850,N_24848);
nor UO_2766 (O_2766,N_23219,N_22749);
xor UO_2767 (O_2767,N_23526,N_24166);
and UO_2768 (O_2768,N_22795,N_24805);
nor UO_2769 (O_2769,N_23699,N_24546);
nand UO_2770 (O_2770,N_22758,N_22331);
or UO_2771 (O_2771,N_24681,N_22363);
nor UO_2772 (O_2772,N_24485,N_23109);
xor UO_2773 (O_2773,N_22180,N_23620);
and UO_2774 (O_2774,N_24663,N_24912);
and UO_2775 (O_2775,N_24946,N_24837);
or UO_2776 (O_2776,N_23168,N_24853);
and UO_2777 (O_2777,N_24119,N_22011);
or UO_2778 (O_2778,N_22695,N_24518);
nor UO_2779 (O_2779,N_21901,N_23830);
nor UO_2780 (O_2780,N_22415,N_24733);
and UO_2781 (O_2781,N_23699,N_22442);
and UO_2782 (O_2782,N_23702,N_22065);
or UO_2783 (O_2783,N_22238,N_24902);
or UO_2784 (O_2784,N_22657,N_22315);
or UO_2785 (O_2785,N_22999,N_23029);
nor UO_2786 (O_2786,N_24010,N_24368);
nor UO_2787 (O_2787,N_24355,N_23014);
nor UO_2788 (O_2788,N_23052,N_23619);
nand UO_2789 (O_2789,N_24351,N_23024);
nor UO_2790 (O_2790,N_24603,N_24839);
nand UO_2791 (O_2791,N_23747,N_22731);
and UO_2792 (O_2792,N_23123,N_23171);
xnor UO_2793 (O_2793,N_22419,N_23660);
or UO_2794 (O_2794,N_22322,N_23101);
and UO_2795 (O_2795,N_24303,N_22098);
nor UO_2796 (O_2796,N_24602,N_22668);
nand UO_2797 (O_2797,N_22058,N_23828);
xnor UO_2798 (O_2798,N_24831,N_23165);
and UO_2799 (O_2799,N_21977,N_22910);
nand UO_2800 (O_2800,N_23407,N_23516);
nand UO_2801 (O_2801,N_22796,N_23621);
or UO_2802 (O_2802,N_24735,N_23041);
and UO_2803 (O_2803,N_22661,N_23560);
nor UO_2804 (O_2804,N_24113,N_23746);
and UO_2805 (O_2805,N_23201,N_24747);
nand UO_2806 (O_2806,N_23209,N_22274);
nand UO_2807 (O_2807,N_22755,N_24403);
nand UO_2808 (O_2808,N_24420,N_22820);
xnor UO_2809 (O_2809,N_24326,N_22109);
or UO_2810 (O_2810,N_24891,N_22505);
or UO_2811 (O_2811,N_22824,N_23185);
and UO_2812 (O_2812,N_22406,N_24718);
and UO_2813 (O_2813,N_23977,N_22057);
or UO_2814 (O_2814,N_24768,N_23405);
nor UO_2815 (O_2815,N_22491,N_23022);
nor UO_2816 (O_2816,N_24719,N_23052);
nand UO_2817 (O_2817,N_24342,N_22317);
and UO_2818 (O_2818,N_24962,N_21937);
xnor UO_2819 (O_2819,N_24481,N_22271);
or UO_2820 (O_2820,N_23023,N_23822);
and UO_2821 (O_2821,N_22726,N_24703);
nor UO_2822 (O_2822,N_22514,N_24513);
nor UO_2823 (O_2823,N_24109,N_24339);
nand UO_2824 (O_2824,N_23632,N_23743);
nor UO_2825 (O_2825,N_24215,N_23612);
xor UO_2826 (O_2826,N_23852,N_23053);
or UO_2827 (O_2827,N_24292,N_24763);
nand UO_2828 (O_2828,N_23151,N_23321);
and UO_2829 (O_2829,N_22172,N_24476);
or UO_2830 (O_2830,N_22371,N_22127);
nor UO_2831 (O_2831,N_22897,N_24515);
or UO_2832 (O_2832,N_22384,N_23921);
and UO_2833 (O_2833,N_23032,N_23543);
or UO_2834 (O_2834,N_23320,N_22487);
nand UO_2835 (O_2835,N_22766,N_22758);
nand UO_2836 (O_2836,N_23671,N_24042);
nand UO_2837 (O_2837,N_24507,N_23057);
nor UO_2838 (O_2838,N_22420,N_24479);
nand UO_2839 (O_2839,N_24061,N_23452);
xnor UO_2840 (O_2840,N_23339,N_23485);
nor UO_2841 (O_2841,N_22081,N_22154);
nor UO_2842 (O_2842,N_23173,N_24944);
nand UO_2843 (O_2843,N_21922,N_23895);
or UO_2844 (O_2844,N_23862,N_24218);
xor UO_2845 (O_2845,N_23035,N_24785);
and UO_2846 (O_2846,N_22133,N_23335);
nand UO_2847 (O_2847,N_23804,N_24133);
and UO_2848 (O_2848,N_23179,N_24154);
or UO_2849 (O_2849,N_22238,N_24142);
or UO_2850 (O_2850,N_24303,N_21986);
xnor UO_2851 (O_2851,N_22870,N_22851);
and UO_2852 (O_2852,N_23014,N_24930);
or UO_2853 (O_2853,N_24067,N_24579);
xor UO_2854 (O_2854,N_23631,N_24106);
and UO_2855 (O_2855,N_24479,N_23881);
and UO_2856 (O_2856,N_24675,N_23614);
nand UO_2857 (O_2857,N_24033,N_23875);
nor UO_2858 (O_2858,N_21902,N_24451);
or UO_2859 (O_2859,N_24652,N_23834);
xor UO_2860 (O_2860,N_24138,N_24721);
and UO_2861 (O_2861,N_23553,N_24244);
nor UO_2862 (O_2862,N_22145,N_22322);
nand UO_2863 (O_2863,N_23151,N_22767);
and UO_2864 (O_2864,N_22588,N_23595);
xnor UO_2865 (O_2865,N_23879,N_24317);
nand UO_2866 (O_2866,N_24366,N_24732);
and UO_2867 (O_2867,N_24109,N_22313);
xor UO_2868 (O_2868,N_22767,N_23959);
nor UO_2869 (O_2869,N_24340,N_24558);
or UO_2870 (O_2870,N_24030,N_23741);
nor UO_2871 (O_2871,N_22160,N_22340);
and UO_2872 (O_2872,N_22236,N_22695);
nor UO_2873 (O_2873,N_23004,N_22888);
or UO_2874 (O_2874,N_24234,N_23310);
and UO_2875 (O_2875,N_24417,N_22139);
and UO_2876 (O_2876,N_23534,N_22369);
or UO_2877 (O_2877,N_23309,N_24831);
nor UO_2878 (O_2878,N_23441,N_23565);
nand UO_2879 (O_2879,N_22932,N_23347);
or UO_2880 (O_2880,N_23356,N_24749);
or UO_2881 (O_2881,N_24149,N_24846);
xor UO_2882 (O_2882,N_24816,N_23078);
xnor UO_2883 (O_2883,N_23773,N_22100);
nor UO_2884 (O_2884,N_22722,N_24522);
or UO_2885 (O_2885,N_22960,N_21988);
xor UO_2886 (O_2886,N_22839,N_22834);
xnor UO_2887 (O_2887,N_23502,N_24372);
nand UO_2888 (O_2888,N_24924,N_22288);
nand UO_2889 (O_2889,N_23560,N_23523);
and UO_2890 (O_2890,N_22087,N_23659);
nor UO_2891 (O_2891,N_22647,N_23643);
nor UO_2892 (O_2892,N_22113,N_21922);
and UO_2893 (O_2893,N_23679,N_24457);
nor UO_2894 (O_2894,N_23808,N_22878);
nor UO_2895 (O_2895,N_22121,N_24882);
xor UO_2896 (O_2896,N_23949,N_22238);
or UO_2897 (O_2897,N_22438,N_24508);
nand UO_2898 (O_2898,N_22756,N_22291);
and UO_2899 (O_2899,N_22811,N_22969);
nand UO_2900 (O_2900,N_23590,N_23016);
and UO_2901 (O_2901,N_24719,N_22736);
nor UO_2902 (O_2902,N_22738,N_21895);
nand UO_2903 (O_2903,N_23536,N_22091);
xnor UO_2904 (O_2904,N_23590,N_22953);
or UO_2905 (O_2905,N_23952,N_21882);
or UO_2906 (O_2906,N_24042,N_21897);
nor UO_2907 (O_2907,N_24018,N_24643);
and UO_2908 (O_2908,N_22439,N_22448);
or UO_2909 (O_2909,N_24294,N_24959);
and UO_2910 (O_2910,N_23289,N_24713);
nand UO_2911 (O_2911,N_22453,N_24798);
nand UO_2912 (O_2912,N_23043,N_22033);
nor UO_2913 (O_2913,N_23924,N_24520);
nor UO_2914 (O_2914,N_22473,N_22639);
or UO_2915 (O_2915,N_23630,N_22980);
xor UO_2916 (O_2916,N_21899,N_22257);
xor UO_2917 (O_2917,N_22740,N_21966);
and UO_2918 (O_2918,N_24417,N_23363);
or UO_2919 (O_2919,N_24708,N_24094);
and UO_2920 (O_2920,N_24351,N_22961);
xnor UO_2921 (O_2921,N_22611,N_23172);
nand UO_2922 (O_2922,N_23416,N_22431);
nor UO_2923 (O_2923,N_23109,N_24601);
nand UO_2924 (O_2924,N_23944,N_24173);
or UO_2925 (O_2925,N_22319,N_22717);
and UO_2926 (O_2926,N_24117,N_23453);
xor UO_2927 (O_2927,N_21938,N_23742);
nor UO_2928 (O_2928,N_22811,N_22693);
and UO_2929 (O_2929,N_24616,N_23558);
nor UO_2930 (O_2930,N_23636,N_24514);
and UO_2931 (O_2931,N_22619,N_24272);
xor UO_2932 (O_2932,N_24161,N_22361);
nand UO_2933 (O_2933,N_24762,N_23818);
and UO_2934 (O_2934,N_22880,N_22573);
and UO_2935 (O_2935,N_23263,N_23577);
xor UO_2936 (O_2936,N_23957,N_23922);
nor UO_2937 (O_2937,N_22188,N_23637);
nand UO_2938 (O_2938,N_23263,N_22693);
or UO_2939 (O_2939,N_24433,N_24015);
or UO_2940 (O_2940,N_22521,N_24153);
nand UO_2941 (O_2941,N_23950,N_22291);
and UO_2942 (O_2942,N_21990,N_23703);
xnor UO_2943 (O_2943,N_22618,N_24138);
and UO_2944 (O_2944,N_23677,N_23427);
and UO_2945 (O_2945,N_22854,N_24296);
nand UO_2946 (O_2946,N_24262,N_23099);
nor UO_2947 (O_2947,N_24407,N_24867);
and UO_2948 (O_2948,N_24424,N_22307);
or UO_2949 (O_2949,N_22442,N_23621);
or UO_2950 (O_2950,N_23375,N_22634);
and UO_2951 (O_2951,N_24447,N_23216);
nand UO_2952 (O_2952,N_22295,N_23098);
nor UO_2953 (O_2953,N_23424,N_24330);
nand UO_2954 (O_2954,N_23880,N_22763);
nor UO_2955 (O_2955,N_22500,N_24211);
or UO_2956 (O_2956,N_23412,N_22706);
nand UO_2957 (O_2957,N_22396,N_22263);
and UO_2958 (O_2958,N_22226,N_23897);
or UO_2959 (O_2959,N_24684,N_23411);
nor UO_2960 (O_2960,N_23480,N_23497);
nor UO_2961 (O_2961,N_24004,N_24239);
or UO_2962 (O_2962,N_23467,N_23760);
or UO_2963 (O_2963,N_23794,N_23454);
or UO_2964 (O_2964,N_23185,N_22064);
nand UO_2965 (O_2965,N_24241,N_23056);
nor UO_2966 (O_2966,N_23259,N_24471);
or UO_2967 (O_2967,N_24606,N_22823);
nand UO_2968 (O_2968,N_23472,N_22889);
and UO_2969 (O_2969,N_22523,N_22798);
and UO_2970 (O_2970,N_22171,N_21977);
and UO_2971 (O_2971,N_21898,N_24179);
and UO_2972 (O_2972,N_22624,N_21945);
nor UO_2973 (O_2973,N_22745,N_23657);
nor UO_2974 (O_2974,N_23866,N_23822);
or UO_2975 (O_2975,N_24888,N_24980);
xor UO_2976 (O_2976,N_23008,N_21929);
nand UO_2977 (O_2977,N_23474,N_24738);
xor UO_2978 (O_2978,N_21953,N_23236);
nand UO_2979 (O_2979,N_23858,N_24091);
or UO_2980 (O_2980,N_24611,N_23413);
or UO_2981 (O_2981,N_24200,N_23915);
and UO_2982 (O_2982,N_24166,N_22131);
and UO_2983 (O_2983,N_24080,N_23763);
nor UO_2984 (O_2984,N_22646,N_22725);
or UO_2985 (O_2985,N_23912,N_23004);
nor UO_2986 (O_2986,N_23530,N_24425);
xnor UO_2987 (O_2987,N_23697,N_22589);
or UO_2988 (O_2988,N_23287,N_23726);
xnor UO_2989 (O_2989,N_23533,N_22417);
nand UO_2990 (O_2990,N_22506,N_23707);
xor UO_2991 (O_2991,N_22024,N_24604);
nor UO_2992 (O_2992,N_24374,N_22148);
nor UO_2993 (O_2993,N_24612,N_22480);
and UO_2994 (O_2994,N_23844,N_23370);
xor UO_2995 (O_2995,N_23651,N_22042);
xnor UO_2996 (O_2996,N_22664,N_23638);
xor UO_2997 (O_2997,N_21943,N_22257);
and UO_2998 (O_2998,N_24111,N_22935);
or UO_2999 (O_2999,N_24555,N_24030);
endmodule