module basic_500_3000_500_5_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_176,In_435);
nor U1 (N_1,In_392,In_372);
or U2 (N_2,In_113,In_79);
and U3 (N_3,In_404,In_41);
nand U4 (N_4,In_199,In_377);
and U5 (N_5,In_452,In_354);
or U6 (N_6,In_8,In_105);
or U7 (N_7,In_429,In_461);
xnor U8 (N_8,In_60,In_92);
or U9 (N_9,In_385,In_38);
nor U10 (N_10,In_467,In_151);
and U11 (N_11,In_69,In_171);
nor U12 (N_12,In_177,In_244);
nand U13 (N_13,In_325,In_450);
nor U14 (N_14,In_490,In_247);
and U15 (N_15,In_342,In_389);
nand U16 (N_16,In_123,In_102);
and U17 (N_17,In_403,In_219);
and U18 (N_18,In_388,In_178);
or U19 (N_19,In_266,In_409);
and U20 (N_20,In_390,In_246);
or U21 (N_21,In_417,In_65);
or U22 (N_22,In_71,In_98);
and U23 (N_23,In_215,In_464);
nand U24 (N_24,In_424,In_360);
nor U25 (N_25,In_327,In_411);
and U26 (N_26,In_191,In_357);
nor U27 (N_27,In_498,In_434);
nand U28 (N_28,In_96,In_276);
or U29 (N_29,In_27,In_189);
nand U30 (N_30,In_363,In_295);
nor U31 (N_31,In_317,In_449);
nor U32 (N_32,In_154,In_144);
or U33 (N_33,In_400,In_164);
nand U34 (N_34,In_155,In_413);
nand U35 (N_35,In_208,In_355);
nor U36 (N_36,In_93,In_15);
nand U37 (N_37,In_402,In_484);
nand U38 (N_38,In_456,In_274);
nor U39 (N_39,In_222,In_420);
nand U40 (N_40,In_486,In_476);
nor U41 (N_41,In_73,In_153);
and U42 (N_42,In_200,In_234);
and U43 (N_43,In_462,In_39);
or U44 (N_44,In_135,In_380);
or U45 (N_45,In_255,In_346);
nor U46 (N_46,In_235,In_344);
nand U47 (N_47,In_386,In_336);
nor U48 (N_48,In_109,In_348);
and U49 (N_49,In_114,In_283);
nor U50 (N_50,In_211,In_112);
nand U51 (N_51,In_125,In_87);
and U52 (N_52,In_333,In_243);
nand U53 (N_53,In_481,In_425);
nand U54 (N_54,In_157,In_458);
nor U55 (N_55,In_373,In_488);
or U56 (N_56,In_119,In_227);
xor U57 (N_57,In_459,In_339);
and U58 (N_58,In_395,In_312);
or U59 (N_59,In_127,In_492);
nor U60 (N_60,In_24,In_401);
or U61 (N_61,In_122,In_58);
or U62 (N_62,In_307,In_453);
and U63 (N_63,In_1,In_361);
nand U64 (N_64,In_22,In_381);
and U65 (N_65,In_32,In_260);
or U66 (N_66,In_131,In_173);
nand U67 (N_67,In_95,In_257);
and U68 (N_68,In_397,In_382);
nor U69 (N_69,In_341,In_188);
or U70 (N_70,In_40,In_9);
nand U71 (N_71,In_223,In_310);
and U72 (N_72,In_440,In_72);
nand U73 (N_73,In_258,In_54);
and U74 (N_74,In_265,In_427);
and U75 (N_75,In_76,In_80);
and U76 (N_76,In_207,In_5);
nand U77 (N_77,In_47,In_451);
nor U78 (N_78,In_419,In_11);
nand U79 (N_79,In_110,In_124);
or U80 (N_80,In_31,In_68);
nor U81 (N_81,In_170,In_82);
xor U82 (N_82,In_286,In_81);
nand U83 (N_83,In_431,In_268);
or U84 (N_84,In_328,In_428);
and U85 (N_85,In_469,In_35);
or U86 (N_86,In_314,In_245);
or U87 (N_87,In_85,In_349);
nand U88 (N_88,In_140,In_470);
or U89 (N_89,In_479,In_220);
or U90 (N_90,In_120,In_248);
or U91 (N_91,In_229,In_213);
nor U92 (N_92,In_167,In_489);
nand U93 (N_93,In_443,In_446);
nand U94 (N_94,In_26,In_273);
or U95 (N_95,In_480,In_2);
nor U96 (N_96,In_291,In_193);
and U97 (N_97,In_426,In_90);
nor U98 (N_98,In_437,In_324);
or U99 (N_99,In_237,In_137);
nor U100 (N_100,In_201,In_30);
or U101 (N_101,In_297,In_279);
and U102 (N_102,In_74,In_23);
and U103 (N_103,In_10,In_146);
or U104 (N_104,In_66,In_3);
or U105 (N_105,In_107,In_353);
and U106 (N_106,In_351,In_298);
nor U107 (N_107,In_77,In_168);
nand U108 (N_108,In_442,In_166);
xnor U109 (N_109,In_371,In_309);
or U110 (N_110,In_315,In_362);
nand U111 (N_111,In_145,In_44);
and U112 (N_112,In_366,In_350);
or U113 (N_113,In_115,In_196);
nor U114 (N_114,In_141,In_230);
and U115 (N_115,In_267,In_455);
nor U116 (N_116,In_318,In_147);
nor U117 (N_117,In_59,In_422);
nor U118 (N_118,In_218,In_457);
or U119 (N_119,In_280,In_423);
nand U120 (N_120,In_6,In_226);
or U121 (N_121,In_97,In_225);
nand U122 (N_122,In_214,In_473);
and U123 (N_123,In_421,In_84);
nor U124 (N_124,In_477,In_187);
and U125 (N_125,In_104,In_180);
and U126 (N_126,In_364,In_332);
and U127 (N_127,In_83,In_275);
nor U128 (N_128,In_195,In_101);
xor U129 (N_129,In_204,In_4);
and U130 (N_130,In_485,In_17);
nand U131 (N_131,In_209,In_272);
and U132 (N_132,In_496,In_182);
or U133 (N_133,In_439,In_284);
or U134 (N_134,In_345,In_499);
or U135 (N_135,In_259,In_185);
and U136 (N_136,In_210,In_67);
and U137 (N_137,In_475,In_399);
and U138 (N_138,In_378,In_368);
nand U139 (N_139,In_48,In_251);
or U140 (N_140,In_50,In_337);
nor U141 (N_141,In_43,In_138);
or U142 (N_142,In_282,In_483);
and U143 (N_143,In_281,In_487);
nand U144 (N_144,In_376,In_448);
nor U145 (N_145,In_57,In_190);
or U146 (N_146,In_88,In_306);
or U147 (N_147,In_416,In_51);
and U148 (N_148,In_472,In_197);
or U149 (N_149,In_296,In_302);
nor U150 (N_150,In_148,In_288);
nand U151 (N_151,In_42,In_497);
nand U152 (N_152,In_316,In_165);
nor U153 (N_153,In_19,In_78);
nor U154 (N_154,In_28,In_216);
and U155 (N_155,In_0,In_61);
or U156 (N_156,In_264,In_183);
or U157 (N_157,In_46,In_460);
or U158 (N_158,In_444,In_319);
and U159 (N_159,In_285,In_174);
nand U160 (N_160,In_13,In_163);
or U161 (N_161,In_12,In_393);
nor U162 (N_162,In_430,In_128);
nor U163 (N_163,In_300,In_94);
xnor U164 (N_164,In_118,In_21);
or U165 (N_165,In_116,In_313);
or U166 (N_166,In_228,In_320);
nand U167 (N_167,In_491,In_249);
nand U168 (N_168,In_108,In_25);
and U169 (N_169,In_175,In_261);
nand U170 (N_170,In_294,In_181);
and U171 (N_171,In_311,In_143);
or U172 (N_172,In_256,In_29);
nand U173 (N_173,In_495,In_263);
nor U174 (N_174,In_156,In_406);
and U175 (N_175,In_270,In_160);
nand U176 (N_176,In_494,In_408);
nor U177 (N_177,In_179,In_55);
nor U178 (N_178,In_172,In_184);
and U179 (N_179,In_252,In_347);
or U180 (N_180,In_384,In_438);
xnor U181 (N_181,In_236,In_387);
xor U182 (N_182,In_482,In_356);
or U183 (N_183,In_326,In_445);
or U184 (N_184,In_329,In_89);
and U185 (N_185,In_52,In_340);
or U186 (N_186,In_262,In_202);
and U187 (N_187,In_405,In_198);
and U188 (N_188,In_308,In_142);
or U189 (N_189,In_396,In_292);
and U190 (N_190,In_303,In_159);
and U191 (N_191,In_86,In_130);
or U192 (N_192,In_322,In_343);
and U193 (N_193,In_139,In_394);
nor U194 (N_194,In_91,In_335);
or U195 (N_195,In_33,In_233);
or U196 (N_196,In_18,In_100);
nand U197 (N_197,In_415,In_454);
nor U198 (N_198,In_134,In_231);
nor U199 (N_199,In_441,In_287);
or U200 (N_200,In_301,In_203);
nor U201 (N_201,In_242,In_103);
or U202 (N_202,In_205,In_224);
and U203 (N_203,In_466,In_239);
nand U204 (N_204,In_99,In_414);
nand U205 (N_205,In_241,In_53);
and U206 (N_206,In_117,In_254);
and U207 (N_207,In_278,In_358);
xnor U208 (N_208,In_289,In_290);
and U209 (N_209,In_238,In_240);
nand U210 (N_210,In_62,In_158);
nand U211 (N_211,In_121,In_493);
or U212 (N_212,In_474,In_304);
and U213 (N_213,In_34,In_149);
nand U214 (N_214,In_169,In_111);
or U215 (N_215,In_129,In_271);
nand U216 (N_216,In_436,In_407);
nand U217 (N_217,In_63,In_162);
nor U218 (N_218,In_468,In_253);
or U219 (N_219,In_432,In_16);
nand U220 (N_220,In_20,In_161);
and U221 (N_221,In_56,In_338);
and U222 (N_222,In_277,In_367);
nand U223 (N_223,In_232,In_305);
nor U224 (N_224,In_410,In_150);
or U225 (N_225,In_217,In_132);
xor U226 (N_226,In_70,In_49);
or U227 (N_227,In_152,In_370);
nor U228 (N_228,In_375,In_64);
nor U229 (N_229,In_37,In_192);
nand U230 (N_230,In_299,In_45);
or U231 (N_231,In_186,In_331);
or U232 (N_232,In_379,In_250);
nand U233 (N_233,In_418,In_206);
nor U234 (N_234,In_194,In_374);
or U235 (N_235,In_478,In_133);
and U236 (N_236,In_7,In_398);
nand U237 (N_237,In_75,In_126);
nand U238 (N_238,In_269,In_330);
nor U239 (N_239,In_106,In_293);
nand U240 (N_240,In_334,In_447);
nand U241 (N_241,In_463,In_383);
and U242 (N_242,In_212,In_352);
nand U243 (N_243,In_391,In_321);
and U244 (N_244,In_14,In_221);
nand U245 (N_245,In_433,In_36);
xnor U246 (N_246,In_412,In_323);
and U247 (N_247,In_465,In_365);
or U248 (N_248,In_369,In_471);
and U249 (N_249,In_359,In_136);
nor U250 (N_250,In_321,In_195);
nand U251 (N_251,In_158,In_394);
and U252 (N_252,In_105,In_482);
or U253 (N_253,In_214,In_253);
nor U254 (N_254,In_248,In_139);
and U255 (N_255,In_444,In_249);
nand U256 (N_256,In_432,In_82);
nor U257 (N_257,In_247,In_448);
nor U258 (N_258,In_462,In_418);
and U259 (N_259,In_463,In_72);
or U260 (N_260,In_348,In_278);
and U261 (N_261,In_367,In_267);
or U262 (N_262,In_258,In_438);
nand U263 (N_263,In_238,In_56);
nand U264 (N_264,In_50,In_57);
and U265 (N_265,In_276,In_236);
nand U266 (N_266,In_96,In_159);
and U267 (N_267,In_97,In_131);
and U268 (N_268,In_450,In_125);
and U269 (N_269,In_323,In_222);
nand U270 (N_270,In_467,In_346);
or U271 (N_271,In_142,In_71);
nor U272 (N_272,In_410,In_385);
and U273 (N_273,In_476,In_469);
or U274 (N_274,In_354,In_210);
and U275 (N_275,In_154,In_29);
xor U276 (N_276,In_272,In_387);
nand U277 (N_277,In_408,In_240);
and U278 (N_278,In_274,In_317);
nand U279 (N_279,In_57,In_328);
or U280 (N_280,In_392,In_272);
and U281 (N_281,In_293,In_370);
or U282 (N_282,In_55,In_363);
nor U283 (N_283,In_356,In_208);
or U284 (N_284,In_249,In_228);
and U285 (N_285,In_485,In_313);
nor U286 (N_286,In_212,In_92);
or U287 (N_287,In_286,In_348);
and U288 (N_288,In_59,In_19);
nand U289 (N_289,In_104,In_332);
nand U290 (N_290,In_48,In_226);
nor U291 (N_291,In_413,In_408);
and U292 (N_292,In_409,In_323);
and U293 (N_293,In_457,In_470);
or U294 (N_294,In_8,In_225);
nor U295 (N_295,In_365,In_167);
and U296 (N_296,In_269,In_411);
or U297 (N_297,In_105,In_489);
and U298 (N_298,In_154,In_279);
nand U299 (N_299,In_90,In_127);
or U300 (N_300,In_278,In_461);
nor U301 (N_301,In_327,In_485);
nand U302 (N_302,In_435,In_198);
nor U303 (N_303,In_422,In_20);
nand U304 (N_304,In_363,In_218);
nor U305 (N_305,In_312,In_293);
and U306 (N_306,In_415,In_284);
nor U307 (N_307,In_181,In_232);
nor U308 (N_308,In_412,In_455);
nand U309 (N_309,In_188,In_389);
and U310 (N_310,In_177,In_292);
nor U311 (N_311,In_235,In_409);
and U312 (N_312,In_172,In_10);
or U313 (N_313,In_152,In_23);
nor U314 (N_314,In_360,In_486);
nor U315 (N_315,In_306,In_169);
or U316 (N_316,In_13,In_404);
nor U317 (N_317,In_390,In_236);
and U318 (N_318,In_253,In_243);
and U319 (N_319,In_20,In_277);
nor U320 (N_320,In_106,In_363);
nand U321 (N_321,In_495,In_219);
and U322 (N_322,In_402,In_235);
nand U323 (N_323,In_391,In_300);
nand U324 (N_324,In_135,In_122);
nand U325 (N_325,In_421,In_114);
nor U326 (N_326,In_490,In_463);
nor U327 (N_327,In_183,In_208);
and U328 (N_328,In_279,In_44);
nor U329 (N_329,In_7,In_456);
or U330 (N_330,In_266,In_301);
nand U331 (N_331,In_109,In_392);
and U332 (N_332,In_395,In_450);
nand U333 (N_333,In_356,In_108);
and U334 (N_334,In_233,In_215);
nor U335 (N_335,In_299,In_97);
and U336 (N_336,In_324,In_110);
nand U337 (N_337,In_217,In_48);
nand U338 (N_338,In_356,In_264);
and U339 (N_339,In_266,In_352);
and U340 (N_340,In_45,In_240);
nor U341 (N_341,In_299,In_200);
or U342 (N_342,In_319,In_183);
and U343 (N_343,In_388,In_300);
and U344 (N_344,In_136,In_56);
and U345 (N_345,In_243,In_420);
and U346 (N_346,In_473,In_114);
nand U347 (N_347,In_102,In_42);
and U348 (N_348,In_172,In_312);
nor U349 (N_349,In_433,In_46);
and U350 (N_350,In_358,In_156);
or U351 (N_351,In_271,In_312);
or U352 (N_352,In_222,In_439);
nand U353 (N_353,In_215,In_445);
nor U354 (N_354,In_91,In_28);
or U355 (N_355,In_168,In_345);
nor U356 (N_356,In_445,In_479);
or U357 (N_357,In_265,In_74);
nand U358 (N_358,In_278,In_338);
nor U359 (N_359,In_230,In_329);
and U360 (N_360,In_93,In_165);
nand U361 (N_361,In_351,In_188);
and U362 (N_362,In_30,In_52);
or U363 (N_363,In_74,In_83);
nor U364 (N_364,In_93,In_273);
nor U365 (N_365,In_241,In_398);
nor U366 (N_366,In_119,In_213);
nor U367 (N_367,In_3,In_372);
nor U368 (N_368,In_254,In_491);
or U369 (N_369,In_289,In_482);
nor U370 (N_370,In_389,In_299);
nand U371 (N_371,In_55,In_57);
or U372 (N_372,In_393,In_30);
nand U373 (N_373,In_105,In_461);
nand U374 (N_374,In_13,In_80);
and U375 (N_375,In_433,In_113);
nor U376 (N_376,In_202,In_356);
nor U377 (N_377,In_37,In_339);
xnor U378 (N_378,In_143,In_134);
and U379 (N_379,In_394,In_284);
nor U380 (N_380,In_331,In_145);
and U381 (N_381,In_287,In_127);
nand U382 (N_382,In_149,In_389);
and U383 (N_383,In_24,In_261);
nor U384 (N_384,In_260,In_336);
nor U385 (N_385,In_41,In_77);
or U386 (N_386,In_401,In_436);
nor U387 (N_387,In_194,In_135);
and U388 (N_388,In_35,In_57);
nor U389 (N_389,In_25,In_265);
nand U390 (N_390,In_210,In_1);
or U391 (N_391,In_21,In_79);
or U392 (N_392,In_4,In_135);
nor U393 (N_393,In_272,In_225);
nand U394 (N_394,In_462,In_29);
nand U395 (N_395,In_478,In_430);
nand U396 (N_396,In_392,In_145);
nand U397 (N_397,In_249,In_448);
and U398 (N_398,In_496,In_74);
nand U399 (N_399,In_289,In_411);
nand U400 (N_400,In_238,In_64);
or U401 (N_401,In_378,In_257);
and U402 (N_402,In_71,In_118);
or U403 (N_403,In_193,In_220);
and U404 (N_404,In_279,In_95);
and U405 (N_405,In_410,In_297);
nor U406 (N_406,In_60,In_159);
or U407 (N_407,In_137,In_485);
nor U408 (N_408,In_232,In_470);
nand U409 (N_409,In_322,In_0);
and U410 (N_410,In_61,In_86);
nor U411 (N_411,In_134,In_145);
or U412 (N_412,In_237,In_27);
or U413 (N_413,In_419,In_57);
or U414 (N_414,In_59,In_17);
nand U415 (N_415,In_53,In_410);
nand U416 (N_416,In_213,In_468);
or U417 (N_417,In_264,In_122);
or U418 (N_418,In_240,In_140);
and U419 (N_419,In_410,In_473);
nor U420 (N_420,In_99,In_67);
nand U421 (N_421,In_134,In_275);
xor U422 (N_422,In_212,In_154);
and U423 (N_423,In_209,In_86);
nor U424 (N_424,In_120,In_398);
and U425 (N_425,In_381,In_250);
nor U426 (N_426,In_246,In_72);
nand U427 (N_427,In_494,In_391);
or U428 (N_428,In_137,In_37);
nor U429 (N_429,In_309,In_330);
and U430 (N_430,In_420,In_488);
or U431 (N_431,In_99,In_200);
or U432 (N_432,In_31,In_48);
or U433 (N_433,In_393,In_29);
nand U434 (N_434,In_22,In_333);
nor U435 (N_435,In_41,In_394);
nand U436 (N_436,In_125,In_324);
or U437 (N_437,In_445,In_206);
and U438 (N_438,In_343,In_290);
and U439 (N_439,In_144,In_160);
nor U440 (N_440,In_102,In_380);
nor U441 (N_441,In_152,In_399);
nand U442 (N_442,In_241,In_465);
and U443 (N_443,In_34,In_422);
or U444 (N_444,In_406,In_231);
or U445 (N_445,In_459,In_93);
or U446 (N_446,In_122,In_67);
nand U447 (N_447,In_495,In_467);
and U448 (N_448,In_320,In_342);
nand U449 (N_449,In_245,In_53);
nand U450 (N_450,In_9,In_264);
and U451 (N_451,In_55,In_33);
nor U452 (N_452,In_446,In_394);
nand U453 (N_453,In_103,In_191);
or U454 (N_454,In_316,In_242);
or U455 (N_455,In_103,In_251);
nor U456 (N_456,In_198,In_411);
nor U457 (N_457,In_481,In_256);
nor U458 (N_458,In_40,In_215);
and U459 (N_459,In_300,In_30);
nand U460 (N_460,In_444,In_202);
nor U461 (N_461,In_68,In_170);
or U462 (N_462,In_155,In_275);
nor U463 (N_463,In_29,In_100);
or U464 (N_464,In_202,In_458);
nor U465 (N_465,In_86,In_370);
nor U466 (N_466,In_490,In_343);
or U467 (N_467,In_416,In_104);
and U468 (N_468,In_140,In_211);
nand U469 (N_469,In_156,In_220);
nor U470 (N_470,In_219,In_473);
or U471 (N_471,In_421,In_272);
nand U472 (N_472,In_276,In_63);
nand U473 (N_473,In_416,In_162);
or U474 (N_474,In_242,In_147);
and U475 (N_475,In_418,In_374);
or U476 (N_476,In_130,In_305);
nand U477 (N_477,In_227,In_29);
nand U478 (N_478,In_121,In_414);
nor U479 (N_479,In_33,In_106);
and U480 (N_480,In_226,In_96);
or U481 (N_481,In_165,In_260);
nand U482 (N_482,In_220,In_99);
or U483 (N_483,In_312,In_154);
nand U484 (N_484,In_33,In_60);
nand U485 (N_485,In_195,In_155);
and U486 (N_486,In_439,In_272);
and U487 (N_487,In_371,In_246);
and U488 (N_488,In_423,In_275);
nand U489 (N_489,In_319,In_255);
nor U490 (N_490,In_32,In_365);
and U491 (N_491,In_103,In_353);
nor U492 (N_492,In_391,In_56);
or U493 (N_493,In_211,In_297);
nor U494 (N_494,In_249,In_487);
nand U495 (N_495,In_333,In_417);
nand U496 (N_496,In_167,In_135);
or U497 (N_497,In_492,In_283);
and U498 (N_498,In_138,In_131);
nor U499 (N_499,In_345,In_489);
or U500 (N_500,In_390,In_381);
nor U501 (N_501,In_106,In_422);
nor U502 (N_502,In_229,In_60);
nor U503 (N_503,In_222,In_477);
or U504 (N_504,In_260,In_289);
or U505 (N_505,In_324,In_405);
nand U506 (N_506,In_254,In_235);
or U507 (N_507,In_439,In_480);
or U508 (N_508,In_420,In_438);
nand U509 (N_509,In_459,In_179);
and U510 (N_510,In_27,In_423);
or U511 (N_511,In_29,In_345);
nand U512 (N_512,In_265,In_309);
nand U513 (N_513,In_133,In_333);
or U514 (N_514,In_442,In_259);
and U515 (N_515,In_432,In_358);
nand U516 (N_516,In_275,In_240);
xor U517 (N_517,In_196,In_34);
or U518 (N_518,In_4,In_235);
nand U519 (N_519,In_21,In_30);
or U520 (N_520,In_47,In_82);
nand U521 (N_521,In_351,In_60);
nor U522 (N_522,In_349,In_201);
nor U523 (N_523,In_250,In_64);
nand U524 (N_524,In_332,In_70);
or U525 (N_525,In_326,In_264);
nand U526 (N_526,In_355,In_78);
nor U527 (N_527,In_190,In_23);
and U528 (N_528,In_33,In_91);
and U529 (N_529,In_491,In_218);
or U530 (N_530,In_210,In_458);
nor U531 (N_531,In_418,In_78);
nor U532 (N_532,In_37,In_173);
or U533 (N_533,In_183,In_344);
nor U534 (N_534,In_488,In_115);
nor U535 (N_535,In_219,In_438);
nand U536 (N_536,In_306,In_150);
nor U537 (N_537,In_296,In_58);
nand U538 (N_538,In_51,In_91);
nor U539 (N_539,In_329,In_284);
nand U540 (N_540,In_168,In_340);
xnor U541 (N_541,In_484,In_380);
and U542 (N_542,In_334,In_275);
or U543 (N_543,In_113,In_124);
and U544 (N_544,In_28,In_80);
nor U545 (N_545,In_16,In_227);
or U546 (N_546,In_42,In_417);
nor U547 (N_547,In_452,In_22);
nor U548 (N_548,In_16,In_318);
nor U549 (N_549,In_449,In_316);
nand U550 (N_550,In_161,In_118);
nor U551 (N_551,In_19,In_272);
nor U552 (N_552,In_168,In_104);
xnor U553 (N_553,In_182,In_318);
nor U554 (N_554,In_326,In_87);
and U555 (N_555,In_167,In_433);
and U556 (N_556,In_307,In_277);
or U557 (N_557,In_494,In_33);
or U558 (N_558,In_395,In_65);
and U559 (N_559,In_57,In_302);
or U560 (N_560,In_441,In_362);
or U561 (N_561,In_494,In_142);
nand U562 (N_562,In_125,In_194);
nand U563 (N_563,In_361,In_492);
nand U564 (N_564,In_467,In_458);
nand U565 (N_565,In_41,In_30);
or U566 (N_566,In_271,In_138);
nor U567 (N_567,In_262,In_216);
nor U568 (N_568,In_344,In_455);
and U569 (N_569,In_66,In_78);
nand U570 (N_570,In_83,In_319);
nor U571 (N_571,In_51,In_79);
and U572 (N_572,In_93,In_364);
or U573 (N_573,In_35,In_152);
nor U574 (N_574,In_62,In_273);
or U575 (N_575,In_25,In_137);
or U576 (N_576,In_265,In_487);
or U577 (N_577,In_63,In_403);
nand U578 (N_578,In_284,In_56);
or U579 (N_579,In_449,In_216);
or U580 (N_580,In_302,In_456);
or U581 (N_581,In_435,In_175);
nand U582 (N_582,In_113,In_373);
xor U583 (N_583,In_262,In_40);
nor U584 (N_584,In_139,In_374);
or U585 (N_585,In_388,In_136);
nand U586 (N_586,In_316,In_117);
or U587 (N_587,In_65,In_4);
and U588 (N_588,In_52,In_369);
nor U589 (N_589,In_352,In_193);
nand U590 (N_590,In_374,In_185);
xnor U591 (N_591,In_97,In_70);
and U592 (N_592,In_201,In_223);
and U593 (N_593,In_248,In_204);
nand U594 (N_594,In_439,In_333);
and U595 (N_595,In_74,In_213);
nor U596 (N_596,In_468,In_30);
and U597 (N_597,In_229,In_75);
nand U598 (N_598,In_336,In_193);
or U599 (N_599,In_113,In_200);
and U600 (N_600,N_558,N_570);
nor U601 (N_601,N_54,N_374);
xor U602 (N_602,N_457,N_201);
and U603 (N_603,N_64,N_135);
nand U604 (N_604,N_398,N_517);
nor U605 (N_605,N_399,N_118);
or U606 (N_606,N_475,N_252);
nor U607 (N_607,N_486,N_230);
nor U608 (N_608,N_577,N_199);
and U609 (N_609,N_358,N_341);
and U610 (N_610,N_216,N_43);
nor U611 (N_611,N_593,N_169);
nor U612 (N_612,N_172,N_537);
nor U613 (N_613,N_328,N_61);
nand U614 (N_614,N_109,N_559);
nand U615 (N_615,N_207,N_287);
or U616 (N_616,N_412,N_275);
nand U617 (N_617,N_149,N_366);
or U618 (N_618,N_117,N_292);
or U619 (N_619,N_270,N_178);
xnor U620 (N_620,N_533,N_331);
nand U621 (N_621,N_464,N_567);
nand U622 (N_622,N_102,N_566);
nor U623 (N_623,N_493,N_211);
nor U624 (N_624,N_373,N_29);
and U625 (N_625,N_309,N_186);
nand U626 (N_626,N_532,N_385);
or U627 (N_627,N_53,N_599);
or U628 (N_628,N_195,N_91);
nand U629 (N_629,N_62,N_98);
and U630 (N_630,N_500,N_498);
nor U631 (N_631,N_286,N_254);
and U632 (N_632,N_454,N_145);
and U633 (N_633,N_370,N_89);
xnor U634 (N_634,N_393,N_356);
and U635 (N_635,N_143,N_585);
and U636 (N_636,N_239,N_535);
nand U637 (N_637,N_438,N_364);
nor U638 (N_638,N_227,N_88);
nor U639 (N_639,N_137,N_241);
nor U640 (N_640,N_168,N_305);
nor U641 (N_641,N_487,N_437);
nand U642 (N_642,N_588,N_442);
nor U643 (N_643,N_506,N_565);
xor U644 (N_644,N_446,N_189);
nor U645 (N_645,N_104,N_416);
and U646 (N_646,N_428,N_329);
nand U647 (N_647,N_233,N_285);
nor U648 (N_648,N_108,N_190);
or U649 (N_649,N_41,N_209);
or U650 (N_650,N_379,N_539);
xnor U651 (N_651,N_140,N_403);
or U652 (N_652,N_449,N_543);
nor U653 (N_653,N_161,N_293);
or U654 (N_654,N_184,N_150);
or U655 (N_655,N_170,N_520);
xnor U656 (N_656,N_455,N_4);
nand U657 (N_657,N_522,N_492);
or U658 (N_658,N_353,N_116);
or U659 (N_659,N_74,N_278);
or U660 (N_660,N_362,N_39);
nand U661 (N_661,N_431,N_361);
and U662 (N_662,N_544,N_295);
nand U663 (N_663,N_37,N_282);
or U664 (N_664,N_504,N_294);
or U665 (N_665,N_246,N_365);
nand U666 (N_666,N_488,N_156);
nand U667 (N_667,N_47,N_525);
or U668 (N_668,N_501,N_268);
or U669 (N_669,N_269,N_237);
and U670 (N_670,N_210,N_404);
and U671 (N_671,N_551,N_23);
and U672 (N_672,N_218,N_141);
or U673 (N_673,N_56,N_472);
or U674 (N_674,N_394,N_99);
nor U675 (N_675,N_524,N_306);
nand U676 (N_676,N_144,N_598);
nor U677 (N_677,N_65,N_477);
and U678 (N_678,N_253,N_129);
and U679 (N_679,N_244,N_107);
or U680 (N_680,N_193,N_166);
nand U681 (N_681,N_380,N_279);
and U682 (N_682,N_511,N_489);
or U683 (N_683,N_10,N_273);
and U684 (N_684,N_38,N_461);
nor U685 (N_685,N_490,N_213);
or U686 (N_686,N_342,N_127);
or U687 (N_687,N_304,N_513);
or U688 (N_688,N_214,N_155);
nand U689 (N_689,N_72,N_20);
nand U690 (N_690,N_238,N_519);
or U691 (N_691,N_540,N_34);
and U692 (N_692,N_68,N_435);
and U693 (N_693,N_443,N_436);
or U694 (N_694,N_13,N_27);
or U695 (N_695,N_527,N_222);
and U696 (N_696,N_575,N_298);
or U697 (N_697,N_71,N_384);
nand U698 (N_698,N_348,N_45);
or U699 (N_699,N_174,N_499);
nor U700 (N_700,N_354,N_367);
or U701 (N_701,N_159,N_330);
or U702 (N_702,N_447,N_549);
nor U703 (N_703,N_202,N_235);
or U704 (N_704,N_456,N_473);
nand U705 (N_705,N_30,N_547);
and U706 (N_706,N_564,N_265);
nand U707 (N_707,N_314,N_458);
or U708 (N_708,N_267,N_103);
and U709 (N_709,N_471,N_263);
or U710 (N_710,N_121,N_70);
or U711 (N_711,N_204,N_125);
nor U712 (N_712,N_459,N_16);
xor U713 (N_713,N_548,N_576);
nand U714 (N_714,N_360,N_171);
and U715 (N_715,N_440,N_100);
nor U716 (N_716,N_14,N_280);
or U717 (N_717,N_531,N_448);
and U718 (N_718,N_6,N_590);
or U719 (N_719,N_90,N_261);
or U720 (N_720,N_553,N_200);
nor U721 (N_721,N_28,N_9);
nor U722 (N_722,N_153,N_523);
and U723 (N_723,N_297,N_220);
nand U724 (N_724,N_321,N_332);
or U725 (N_725,N_48,N_79);
nor U726 (N_726,N_378,N_248);
nand U727 (N_727,N_391,N_568);
nor U728 (N_728,N_439,N_26);
nor U729 (N_729,N_73,N_232);
nor U730 (N_730,N_77,N_78);
or U731 (N_731,N_180,N_101);
nand U732 (N_732,N_441,N_465);
or U733 (N_733,N_333,N_162);
nand U734 (N_734,N_327,N_479);
or U735 (N_735,N_18,N_390);
and U736 (N_736,N_318,N_433);
or U737 (N_737,N_343,N_434);
nor U738 (N_738,N_518,N_132);
and U739 (N_739,N_120,N_468);
or U740 (N_740,N_388,N_242);
nand U741 (N_741,N_7,N_445);
or U742 (N_742,N_80,N_592);
and U743 (N_743,N_346,N_396);
and U744 (N_744,N_369,N_50);
nand U745 (N_745,N_290,N_19);
nor U746 (N_746,N_301,N_260);
nor U747 (N_747,N_582,N_320);
and U748 (N_748,N_452,N_427);
and U749 (N_749,N_389,N_316);
nand U750 (N_750,N_583,N_347);
nor U751 (N_751,N_281,N_325);
or U752 (N_752,N_587,N_160);
or U753 (N_753,N_276,N_485);
and U754 (N_754,N_417,N_251);
or U755 (N_755,N_429,N_49);
nor U756 (N_756,N_175,N_315);
and U757 (N_757,N_187,N_382);
nand U758 (N_758,N_467,N_421);
nand U759 (N_759,N_406,N_383);
and U760 (N_760,N_115,N_188);
nand U761 (N_761,N_40,N_550);
xnor U762 (N_762,N_336,N_0);
or U763 (N_763,N_397,N_418);
or U764 (N_764,N_63,N_512);
nand U765 (N_765,N_257,N_51);
or U766 (N_766,N_212,N_158);
nand U767 (N_767,N_494,N_334);
and U768 (N_768,N_596,N_432);
and U769 (N_769,N_584,N_528);
nor U770 (N_770,N_515,N_131);
and U771 (N_771,N_338,N_480);
or U772 (N_772,N_67,N_572);
nor U773 (N_773,N_484,N_60);
and U774 (N_774,N_476,N_84);
nor U775 (N_775,N_381,N_546);
nor U776 (N_776,N_81,N_142);
and U777 (N_777,N_194,N_478);
and U778 (N_778,N_224,N_296);
or U779 (N_779,N_368,N_250);
nand U780 (N_780,N_372,N_249);
xor U781 (N_781,N_217,N_482);
nor U782 (N_782,N_495,N_196);
nor U783 (N_783,N_387,N_264);
xor U784 (N_784,N_277,N_355);
or U785 (N_785,N_123,N_205);
nor U786 (N_786,N_262,N_469);
and U787 (N_787,N_554,N_221);
nor U788 (N_788,N_339,N_119);
or U789 (N_789,N_597,N_136);
nand U790 (N_790,N_534,N_271);
and U791 (N_791,N_502,N_148);
nor U792 (N_792,N_594,N_173);
or U793 (N_793,N_573,N_110);
and U794 (N_794,N_185,N_312);
nor U795 (N_795,N_530,N_113);
and U796 (N_796,N_133,N_283);
and U797 (N_797,N_176,N_307);
and U798 (N_798,N_344,N_538);
and U799 (N_799,N_337,N_351);
nor U800 (N_800,N_401,N_579);
and U801 (N_801,N_272,N_291);
xnor U802 (N_802,N_557,N_560);
and U803 (N_803,N_243,N_408);
and U804 (N_804,N_76,N_508);
and U805 (N_805,N_411,N_430);
and U806 (N_806,N_52,N_147);
nand U807 (N_807,N_496,N_55);
and U808 (N_808,N_44,N_154);
nand U809 (N_809,N_580,N_376);
or U810 (N_810,N_208,N_300);
nor U811 (N_811,N_335,N_12);
or U812 (N_812,N_92,N_424);
and U813 (N_813,N_491,N_96);
nor U814 (N_814,N_521,N_31);
or U815 (N_815,N_138,N_42);
or U816 (N_816,N_24,N_310);
or U817 (N_817,N_58,N_359);
and U818 (N_818,N_386,N_470);
nand U819 (N_819,N_563,N_395);
nand U820 (N_820,N_66,N_400);
or U821 (N_821,N_453,N_22);
nor U822 (N_822,N_181,N_545);
or U823 (N_823,N_444,N_503);
or U824 (N_824,N_419,N_422);
nand U825 (N_825,N_128,N_152);
nand U826 (N_826,N_274,N_352);
and U827 (N_827,N_326,N_122);
or U828 (N_828,N_203,N_555);
nand U829 (N_829,N_223,N_32);
or U830 (N_830,N_569,N_466);
and U831 (N_831,N_266,N_595);
nor U832 (N_832,N_191,N_288);
nor U833 (N_833,N_556,N_192);
nand U834 (N_834,N_284,N_256);
nand U835 (N_835,N_198,N_231);
and U836 (N_836,N_371,N_112);
nor U837 (N_837,N_59,N_2);
or U838 (N_838,N_299,N_345);
and U839 (N_839,N_83,N_322);
and U840 (N_840,N_11,N_111);
nor U841 (N_841,N_402,N_124);
or U842 (N_842,N_151,N_197);
nor U843 (N_843,N_134,N_349);
nor U844 (N_844,N_57,N_97);
or U845 (N_845,N_33,N_323);
or U846 (N_846,N_126,N_36);
nor U847 (N_847,N_516,N_561);
nand U848 (N_848,N_1,N_423);
or U849 (N_849,N_225,N_303);
and U850 (N_850,N_497,N_226);
or U851 (N_851,N_481,N_392);
or U852 (N_852,N_462,N_308);
and U853 (N_853,N_589,N_591);
xor U854 (N_854,N_165,N_552);
or U855 (N_855,N_258,N_106);
nor U856 (N_856,N_94,N_93);
nand U857 (N_857,N_311,N_460);
and U858 (N_858,N_215,N_229);
nand U859 (N_859,N_426,N_164);
nand U860 (N_860,N_450,N_415);
xnor U861 (N_861,N_409,N_240);
nand U862 (N_862,N_571,N_167);
and U863 (N_863,N_377,N_245);
and U864 (N_864,N_317,N_146);
nor U865 (N_865,N_114,N_228);
nand U866 (N_866,N_206,N_259);
xor U867 (N_867,N_578,N_69);
or U868 (N_868,N_529,N_340);
and U869 (N_869,N_541,N_25);
or U870 (N_870,N_247,N_483);
or U871 (N_871,N_86,N_82);
nand U872 (N_872,N_3,N_375);
and U873 (N_873,N_219,N_324);
nor U874 (N_874,N_363,N_179);
and U875 (N_875,N_350,N_586);
nor U876 (N_876,N_95,N_21);
xnor U877 (N_877,N_15,N_536);
nor U878 (N_878,N_562,N_420);
and U879 (N_879,N_5,N_85);
nand U880 (N_880,N_463,N_46);
or U881 (N_881,N_302,N_182);
nor U882 (N_882,N_509,N_581);
nand U883 (N_883,N_130,N_157);
nor U884 (N_884,N_510,N_183);
or U885 (N_885,N_425,N_255);
nor U886 (N_886,N_87,N_526);
nor U887 (N_887,N_35,N_474);
and U888 (N_888,N_313,N_574);
or U889 (N_889,N_177,N_405);
nor U890 (N_890,N_451,N_413);
and U891 (N_891,N_17,N_75);
and U892 (N_892,N_139,N_542);
or U893 (N_893,N_410,N_8);
nand U894 (N_894,N_514,N_505);
or U895 (N_895,N_507,N_407);
nor U896 (N_896,N_319,N_414);
nand U897 (N_897,N_163,N_357);
and U898 (N_898,N_105,N_234);
nor U899 (N_899,N_289,N_236);
nand U900 (N_900,N_318,N_99);
or U901 (N_901,N_268,N_110);
nor U902 (N_902,N_37,N_166);
and U903 (N_903,N_581,N_531);
nand U904 (N_904,N_280,N_21);
nor U905 (N_905,N_279,N_63);
nor U906 (N_906,N_324,N_182);
and U907 (N_907,N_260,N_1);
and U908 (N_908,N_151,N_287);
or U909 (N_909,N_376,N_141);
nand U910 (N_910,N_296,N_457);
and U911 (N_911,N_25,N_17);
nand U912 (N_912,N_267,N_205);
nor U913 (N_913,N_289,N_472);
nor U914 (N_914,N_255,N_422);
nand U915 (N_915,N_238,N_359);
and U916 (N_916,N_113,N_177);
nor U917 (N_917,N_561,N_206);
nor U918 (N_918,N_471,N_313);
and U919 (N_919,N_512,N_27);
and U920 (N_920,N_578,N_202);
nand U921 (N_921,N_397,N_562);
and U922 (N_922,N_346,N_399);
nand U923 (N_923,N_311,N_227);
or U924 (N_924,N_581,N_535);
or U925 (N_925,N_457,N_374);
nor U926 (N_926,N_593,N_566);
or U927 (N_927,N_550,N_1);
or U928 (N_928,N_219,N_122);
and U929 (N_929,N_396,N_270);
nand U930 (N_930,N_198,N_72);
or U931 (N_931,N_262,N_308);
nor U932 (N_932,N_290,N_480);
nand U933 (N_933,N_508,N_57);
nor U934 (N_934,N_548,N_47);
nand U935 (N_935,N_416,N_213);
nor U936 (N_936,N_340,N_523);
and U937 (N_937,N_188,N_523);
or U938 (N_938,N_360,N_267);
nor U939 (N_939,N_113,N_423);
nand U940 (N_940,N_478,N_422);
nor U941 (N_941,N_408,N_226);
nor U942 (N_942,N_413,N_394);
or U943 (N_943,N_207,N_534);
nor U944 (N_944,N_198,N_286);
and U945 (N_945,N_537,N_187);
or U946 (N_946,N_404,N_74);
or U947 (N_947,N_145,N_72);
nor U948 (N_948,N_566,N_290);
and U949 (N_949,N_437,N_419);
nor U950 (N_950,N_203,N_197);
and U951 (N_951,N_14,N_510);
or U952 (N_952,N_383,N_434);
nand U953 (N_953,N_381,N_533);
or U954 (N_954,N_21,N_304);
nor U955 (N_955,N_126,N_435);
nor U956 (N_956,N_216,N_377);
and U957 (N_957,N_464,N_508);
nand U958 (N_958,N_351,N_590);
nor U959 (N_959,N_474,N_403);
and U960 (N_960,N_179,N_36);
and U961 (N_961,N_181,N_159);
or U962 (N_962,N_51,N_78);
and U963 (N_963,N_552,N_253);
nor U964 (N_964,N_176,N_221);
and U965 (N_965,N_179,N_34);
and U966 (N_966,N_258,N_264);
nand U967 (N_967,N_226,N_413);
nor U968 (N_968,N_522,N_178);
or U969 (N_969,N_276,N_216);
and U970 (N_970,N_480,N_39);
nor U971 (N_971,N_138,N_569);
and U972 (N_972,N_99,N_240);
nand U973 (N_973,N_422,N_69);
and U974 (N_974,N_429,N_241);
nand U975 (N_975,N_248,N_537);
nor U976 (N_976,N_304,N_577);
nor U977 (N_977,N_126,N_446);
nor U978 (N_978,N_159,N_116);
and U979 (N_979,N_574,N_520);
nand U980 (N_980,N_86,N_268);
or U981 (N_981,N_479,N_101);
and U982 (N_982,N_284,N_60);
nand U983 (N_983,N_367,N_239);
nand U984 (N_984,N_289,N_492);
nor U985 (N_985,N_188,N_372);
and U986 (N_986,N_197,N_344);
nand U987 (N_987,N_36,N_533);
nor U988 (N_988,N_346,N_199);
and U989 (N_989,N_212,N_442);
or U990 (N_990,N_181,N_171);
nor U991 (N_991,N_412,N_519);
and U992 (N_992,N_261,N_128);
nand U993 (N_993,N_364,N_587);
nor U994 (N_994,N_28,N_475);
and U995 (N_995,N_126,N_503);
nor U996 (N_996,N_185,N_246);
nor U997 (N_997,N_102,N_460);
nand U998 (N_998,N_376,N_527);
nor U999 (N_999,N_7,N_381);
xnor U1000 (N_1000,N_241,N_393);
and U1001 (N_1001,N_155,N_395);
and U1002 (N_1002,N_486,N_211);
nor U1003 (N_1003,N_517,N_42);
nor U1004 (N_1004,N_156,N_344);
nand U1005 (N_1005,N_29,N_293);
and U1006 (N_1006,N_67,N_274);
nand U1007 (N_1007,N_163,N_455);
or U1008 (N_1008,N_424,N_454);
nor U1009 (N_1009,N_146,N_437);
nand U1010 (N_1010,N_586,N_258);
nand U1011 (N_1011,N_490,N_209);
nand U1012 (N_1012,N_492,N_265);
and U1013 (N_1013,N_152,N_234);
xnor U1014 (N_1014,N_413,N_580);
or U1015 (N_1015,N_496,N_568);
or U1016 (N_1016,N_352,N_103);
nor U1017 (N_1017,N_514,N_166);
or U1018 (N_1018,N_426,N_220);
nor U1019 (N_1019,N_182,N_382);
nand U1020 (N_1020,N_288,N_149);
nor U1021 (N_1021,N_250,N_475);
nand U1022 (N_1022,N_284,N_294);
and U1023 (N_1023,N_86,N_139);
or U1024 (N_1024,N_79,N_269);
nand U1025 (N_1025,N_513,N_599);
or U1026 (N_1026,N_551,N_593);
and U1027 (N_1027,N_505,N_456);
or U1028 (N_1028,N_432,N_49);
or U1029 (N_1029,N_419,N_193);
nor U1030 (N_1030,N_207,N_525);
nor U1031 (N_1031,N_160,N_106);
or U1032 (N_1032,N_408,N_64);
nor U1033 (N_1033,N_52,N_111);
nand U1034 (N_1034,N_519,N_371);
nor U1035 (N_1035,N_504,N_546);
nand U1036 (N_1036,N_461,N_125);
xor U1037 (N_1037,N_329,N_190);
nand U1038 (N_1038,N_545,N_470);
nand U1039 (N_1039,N_539,N_447);
nor U1040 (N_1040,N_15,N_218);
xor U1041 (N_1041,N_380,N_195);
or U1042 (N_1042,N_162,N_157);
and U1043 (N_1043,N_146,N_66);
xor U1044 (N_1044,N_420,N_513);
or U1045 (N_1045,N_266,N_567);
and U1046 (N_1046,N_401,N_39);
nor U1047 (N_1047,N_87,N_507);
nor U1048 (N_1048,N_152,N_441);
and U1049 (N_1049,N_231,N_208);
nor U1050 (N_1050,N_9,N_217);
and U1051 (N_1051,N_591,N_236);
nand U1052 (N_1052,N_271,N_464);
xnor U1053 (N_1053,N_267,N_552);
nand U1054 (N_1054,N_412,N_153);
or U1055 (N_1055,N_313,N_399);
or U1056 (N_1056,N_188,N_579);
nand U1057 (N_1057,N_268,N_513);
and U1058 (N_1058,N_251,N_327);
xnor U1059 (N_1059,N_16,N_235);
nand U1060 (N_1060,N_415,N_367);
and U1061 (N_1061,N_158,N_400);
or U1062 (N_1062,N_80,N_33);
or U1063 (N_1063,N_273,N_379);
or U1064 (N_1064,N_369,N_465);
nor U1065 (N_1065,N_100,N_83);
nor U1066 (N_1066,N_212,N_293);
or U1067 (N_1067,N_345,N_385);
nor U1068 (N_1068,N_81,N_524);
and U1069 (N_1069,N_406,N_248);
nand U1070 (N_1070,N_313,N_596);
nor U1071 (N_1071,N_212,N_167);
nand U1072 (N_1072,N_131,N_328);
nand U1073 (N_1073,N_59,N_176);
or U1074 (N_1074,N_574,N_207);
or U1075 (N_1075,N_513,N_108);
nor U1076 (N_1076,N_331,N_350);
nor U1077 (N_1077,N_159,N_435);
nor U1078 (N_1078,N_134,N_541);
or U1079 (N_1079,N_242,N_496);
nand U1080 (N_1080,N_367,N_385);
nand U1081 (N_1081,N_497,N_566);
nand U1082 (N_1082,N_52,N_226);
or U1083 (N_1083,N_112,N_282);
nand U1084 (N_1084,N_449,N_211);
nor U1085 (N_1085,N_330,N_371);
nor U1086 (N_1086,N_311,N_247);
nor U1087 (N_1087,N_224,N_112);
or U1088 (N_1088,N_343,N_456);
or U1089 (N_1089,N_523,N_144);
or U1090 (N_1090,N_500,N_297);
or U1091 (N_1091,N_480,N_220);
nor U1092 (N_1092,N_554,N_477);
nand U1093 (N_1093,N_514,N_139);
nor U1094 (N_1094,N_301,N_397);
nor U1095 (N_1095,N_405,N_229);
or U1096 (N_1096,N_472,N_538);
nand U1097 (N_1097,N_256,N_211);
nand U1098 (N_1098,N_327,N_222);
nand U1099 (N_1099,N_86,N_394);
and U1100 (N_1100,N_284,N_435);
nor U1101 (N_1101,N_275,N_374);
nor U1102 (N_1102,N_30,N_88);
nor U1103 (N_1103,N_450,N_384);
nand U1104 (N_1104,N_541,N_428);
nand U1105 (N_1105,N_80,N_557);
xnor U1106 (N_1106,N_83,N_488);
and U1107 (N_1107,N_498,N_481);
and U1108 (N_1108,N_330,N_61);
or U1109 (N_1109,N_115,N_13);
nor U1110 (N_1110,N_400,N_362);
nand U1111 (N_1111,N_3,N_211);
nor U1112 (N_1112,N_59,N_34);
nor U1113 (N_1113,N_412,N_179);
or U1114 (N_1114,N_300,N_324);
xor U1115 (N_1115,N_298,N_246);
nor U1116 (N_1116,N_84,N_511);
nand U1117 (N_1117,N_328,N_575);
nand U1118 (N_1118,N_246,N_200);
and U1119 (N_1119,N_586,N_432);
and U1120 (N_1120,N_77,N_135);
and U1121 (N_1121,N_246,N_531);
nor U1122 (N_1122,N_28,N_263);
or U1123 (N_1123,N_463,N_438);
nor U1124 (N_1124,N_569,N_477);
or U1125 (N_1125,N_469,N_6);
nor U1126 (N_1126,N_550,N_365);
and U1127 (N_1127,N_503,N_404);
nand U1128 (N_1128,N_205,N_583);
nor U1129 (N_1129,N_556,N_212);
nor U1130 (N_1130,N_190,N_191);
and U1131 (N_1131,N_312,N_411);
nand U1132 (N_1132,N_18,N_135);
and U1133 (N_1133,N_415,N_59);
nor U1134 (N_1134,N_13,N_107);
nor U1135 (N_1135,N_44,N_100);
nor U1136 (N_1136,N_5,N_500);
nor U1137 (N_1137,N_454,N_68);
nand U1138 (N_1138,N_117,N_344);
nor U1139 (N_1139,N_140,N_158);
xor U1140 (N_1140,N_468,N_274);
nor U1141 (N_1141,N_379,N_550);
or U1142 (N_1142,N_404,N_255);
and U1143 (N_1143,N_485,N_79);
xor U1144 (N_1144,N_491,N_152);
or U1145 (N_1145,N_83,N_135);
or U1146 (N_1146,N_10,N_204);
or U1147 (N_1147,N_529,N_375);
nand U1148 (N_1148,N_598,N_208);
nand U1149 (N_1149,N_310,N_585);
nor U1150 (N_1150,N_421,N_141);
nor U1151 (N_1151,N_84,N_385);
and U1152 (N_1152,N_69,N_376);
or U1153 (N_1153,N_139,N_464);
nor U1154 (N_1154,N_410,N_65);
nor U1155 (N_1155,N_553,N_503);
nor U1156 (N_1156,N_102,N_74);
and U1157 (N_1157,N_84,N_434);
nand U1158 (N_1158,N_299,N_119);
or U1159 (N_1159,N_256,N_238);
nor U1160 (N_1160,N_481,N_115);
nor U1161 (N_1161,N_154,N_231);
and U1162 (N_1162,N_326,N_102);
and U1163 (N_1163,N_361,N_323);
and U1164 (N_1164,N_267,N_28);
and U1165 (N_1165,N_473,N_10);
xnor U1166 (N_1166,N_278,N_510);
nor U1167 (N_1167,N_512,N_551);
nand U1168 (N_1168,N_8,N_197);
nor U1169 (N_1169,N_399,N_121);
or U1170 (N_1170,N_148,N_87);
nand U1171 (N_1171,N_46,N_132);
and U1172 (N_1172,N_341,N_531);
and U1173 (N_1173,N_538,N_505);
or U1174 (N_1174,N_325,N_51);
nor U1175 (N_1175,N_134,N_465);
or U1176 (N_1176,N_12,N_522);
and U1177 (N_1177,N_597,N_367);
nor U1178 (N_1178,N_486,N_48);
nor U1179 (N_1179,N_298,N_407);
and U1180 (N_1180,N_347,N_273);
or U1181 (N_1181,N_140,N_38);
or U1182 (N_1182,N_375,N_101);
nor U1183 (N_1183,N_305,N_594);
nand U1184 (N_1184,N_419,N_90);
nor U1185 (N_1185,N_402,N_174);
or U1186 (N_1186,N_305,N_377);
nor U1187 (N_1187,N_131,N_183);
or U1188 (N_1188,N_571,N_48);
nor U1189 (N_1189,N_277,N_144);
or U1190 (N_1190,N_568,N_488);
nor U1191 (N_1191,N_321,N_38);
nor U1192 (N_1192,N_593,N_131);
nand U1193 (N_1193,N_97,N_338);
nor U1194 (N_1194,N_511,N_45);
and U1195 (N_1195,N_463,N_472);
nand U1196 (N_1196,N_588,N_150);
xnor U1197 (N_1197,N_270,N_300);
or U1198 (N_1198,N_331,N_94);
nand U1199 (N_1199,N_570,N_488);
and U1200 (N_1200,N_691,N_1054);
nand U1201 (N_1201,N_1077,N_1190);
nand U1202 (N_1202,N_910,N_640);
nand U1203 (N_1203,N_925,N_763);
or U1204 (N_1204,N_736,N_972);
nor U1205 (N_1205,N_883,N_1008);
and U1206 (N_1206,N_1127,N_998);
or U1207 (N_1207,N_1068,N_817);
nand U1208 (N_1208,N_710,N_1081);
nand U1209 (N_1209,N_1197,N_909);
and U1210 (N_1210,N_951,N_1089);
or U1211 (N_1211,N_1142,N_865);
nor U1212 (N_1212,N_665,N_666);
and U1213 (N_1213,N_862,N_1122);
nand U1214 (N_1214,N_931,N_784);
and U1215 (N_1215,N_1112,N_1066);
and U1216 (N_1216,N_687,N_1168);
nand U1217 (N_1217,N_908,N_995);
nor U1218 (N_1218,N_1123,N_1098);
and U1219 (N_1219,N_932,N_730);
nor U1220 (N_1220,N_839,N_647);
nand U1221 (N_1221,N_1136,N_844);
nor U1222 (N_1222,N_644,N_786);
or U1223 (N_1223,N_809,N_988);
nand U1224 (N_1224,N_1144,N_620);
nand U1225 (N_1225,N_621,N_626);
nor U1226 (N_1226,N_1117,N_966);
or U1227 (N_1227,N_1103,N_820);
nand U1228 (N_1228,N_846,N_713);
or U1229 (N_1229,N_994,N_828);
nand U1230 (N_1230,N_772,N_1088);
nand U1231 (N_1231,N_624,N_794);
nor U1232 (N_1232,N_717,N_670);
nor U1233 (N_1233,N_878,N_777);
and U1234 (N_1234,N_723,N_943);
and U1235 (N_1235,N_1003,N_1034);
or U1236 (N_1236,N_824,N_742);
xnor U1237 (N_1237,N_1185,N_711);
nand U1238 (N_1238,N_712,N_635);
or U1239 (N_1239,N_975,N_950);
nor U1240 (N_1240,N_1056,N_1111);
nor U1241 (N_1241,N_858,N_1099);
nand U1242 (N_1242,N_1035,N_1134);
nor U1243 (N_1243,N_1194,N_811);
and U1244 (N_1244,N_1082,N_997);
or U1245 (N_1245,N_871,N_1093);
or U1246 (N_1246,N_1120,N_807);
and U1247 (N_1247,N_655,N_1073);
nor U1248 (N_1248,N_1118,N_1029);
or U1249 (N_1249,N_942,N_706);
nor U1250 (N_1250,N_896,N_659);
or U1251 (N_1251,N_1163,N_840);
or U1252 (N_1252,N_979,N_607);
nor U1253 (N_1253,N_753,N_1137);
nand U1254 (N_1254,N_613,N_696);
nand U1255 (N_1255,N_1133,N_926);
nand U1256 (N_1256,N_701,N_922);
or U1257 (N_1257,N_881,N_845);
nor U1258 (N_1258,N_984,N_1047);
or U1259 (N_1259,N_1031,N_917);
and U1260 (N_1260,N_1052,N_882);
nand U1261 (N_1261,N_1028,N_646);
and U1262 (N_1262,N_754,N_652);
or U1263 (N_1263,N_729,N_894);
or U1264 (N_1264,N_747,N_782);
nor U1265 (N_1265,N_808,N_1092);
nand U1266 (N_1266,N_1170,N_802);
nor U1267 (N_1267,N_1044,N_664);
and U1268 (N_1268,N_1062,N_986);
or U1269 (N_1269,N_1116,N_870);
nand U1270 (N_1270,N_1014,N_737);
and U1271 (N_1271,N_1187,N_1143);
nor U1272 (N_1272,N_695,N_1160);
or U1273 (N_1273,N_798,N_916);
and U1274 (N_1274,N_780,N_693);
and U1275 (N_1275,N_958,N_761);
and U1276 (N_1276,N_999,N_911);
nand U1277 (N_1277,N_1076,N_1189);
nand U1278 (N_1278,N_961,N_728);
and U1279 (N_1279,N_1059,N_785);
and U1280 (N_1280,N_604,N_921);
and U1281 (N_1281,N_638,N_676);
or U1282 (N_1282,N_918,N_619);
or U1283 (N_1283,N_980,N_907);
and U1284 (N_1284,N_969,N_949);
or U1285 (N_1285,N_965,N_1017);
and U1286 (N_1286,N_981,N_609);
nand U1287 (N_1287,N_1007,N_775);
or U1288 (N_1288,N_603,N_993);
nor U1289 (N_1289,N_1013,N_987);
nand U1290 (N_1290,N_1004,N_903);
nand U1291 (N_1291,N_978,N_861);
or U1292 (N_1292,N_792,N_684);
nor U1293 (N_1293,N_1039,N_976);
nand U1294 (N_1294,N_797,N_738);
or U1295 (N_1295,N_1074,N_816);
nor U1296 (N_1296,N_1131,N_1049);
nand U1297 (N_1297,N_731,N_641);
and U1298 (N_1298,N_852,N_629);
nor U1299 (N_1299,N_799,N_1001);
and U1300 (N_1300,N_860,N_721);
and U1301 (N_1301,N_1006,N_1141);
nor U1302 (N_1302,N_1179,N_741);
or U1303 (N_1303,N_956,N_1171);
or U1304 (N_1304,N_1057,N_1005);
or U1305 (N_1305,N_1115,N_1140);
nand U1306 (N_1306,N_924,N_855);
nor U1307 (N_1307,N_778,N_1174);
nand U1308 (N_1308,N_834,N_727);
xnor U1309 (N_1309,N_1186,N_899);
nor U1310 (N_1310,N_1095,N_1151);
or U1311 (N_1311,N_822,N_789);
and U1312 (N_1312,N_600,N_906);
nor U1313 (N_1313,N_774,N_851);
nand U1314 (N_1314,N_937,N_623);
and U1315 (N_1315,N_1169,N_1102);
or U1316 (N_1316,N_773,N_915);
nand U1317 (N_1317,N_793,N_1018);
nand U1318 (N_1318,N_838,N_756);
nand U1319 (N_1319,N_867,N_1072);
xor U1320 (N_1320,N_954,N_663);
nor U1321 (N_1321,N_806,N_748);
nand U1322 (N_1322,N_1178,N_1161);
nand U1323 (N_1323,N_847,N_1037);
nand U1324 (N_1324,N_1097,N_971);
nand U1325 (N_1325,N_680,N_1058);
and U1326 (N_1326,N_758,N_933);
and U1327 (N_1327,N_1135,N_708);
and U1328 (N_1328,N_983,N_1158);
and U1329 (N_1329,N_982,N_890);
nor U1330 (N_1330,N_1022,N_694);
nand U1331 (N_1331,N_1070,N_857);
nand U1332 (N_1332,N_945,N_1159);
nand U1333 (N_1333,N_1191,N_1096);
xnor U1334 (N_1334,N_989,N_601);
nor U1335 (N_1335,N_977,N_927);
and U1336 (N_1336,N_892,N_866);
nor U1337 (N_1337,N_1033,N_627);
or U1338 (N_1338,N_726,N_869);
and U1339 (N_1339,N_682,N_1011);
nor U1340 (N_1340,N_1156,N_991);
or U1341 (N_1341,N_749,N_946);
and U1342 (N_1342,N_936,N_920);
or U1343 (N_1343,N_672,N_944);
or U1344 (N_1344,N_656,N_854);
nor U1345 (N_1345,N_677,N_1084);
and U1346 (N_1346,N_678,N_1104);
or U1347 (N_1347,N_760,N_996);
nand U1348 (N_1348,N_853,N_681);
and U1349 (N_1349,N_1038,N_849);
nor U1350 (N_1350,N_889,N_1154);
and U1351 (N_1351,N_650,N_649);
nand U1352 (N_1352,N_764,N_1042);
nand U1353 (N_1353,N_832,N_1045);
nand U1354 (N_1354,N_960,N_795);
nand U1355 (N_1355,N_1162,N_631);
nor U1356 (N_1356,N_1175,N_690);
nand U1357 (N_1357,N_617,N_671);
nor U1358 (N_1358,N_1065,N_990);
or U1359 (N_1359,N_614,N_823);
nor U1360 (N_1360,N_843,N_875);
nand U1361 (N_1361,N_692,N_1105);
nand U1362 (N_1362,N_1138,N_616);
and U1363 (N_1363,N_1119,N_874);
nand U1364 (N_1364,N_891,N_1172);
or U1365 (N_1365,N_715,N_940);
xor U1366 (N_1366,N_1015,N_622);
nor U1367 (N_1367,N_725,N_648);
and U1368 (N_1368,N_645,N_1090);
nor U1369 (N_1369,N_683,N_859);
nand U1370 (N_1370,N_673,N_1150);
nor U1371 (N_1371,N_1046,N_992);
nand U1372 (N_1372,N_643,N_1021);
and U1373 (N_1373,N_697,N_880);
xor U1374 (N_1374,N_699,N_755);
nor U1375 (N_1375,N_939,N_947);
and U1376 (N_1376,N_1173,N_876);
nor U1377 (N_1377,N_1061,N_1107);
nand U1378 (N_1378,N_732,N_733);
and U1379 (N_1379,N_974,N_653);
and U1380 (N_1380,N_759,N_1083);
and U1381 (N_1381,N_1176,N_704);
or U1382 (N_1382,N_743,N_842);
and U1383 (N_1383,N_1026,N_675);
or U1384 (N_1384,N_985,N_897);
and U1385 (N_1385,N_781,N_744);
or U1386 (N_1386,N_800,N_660);
and U1387 (N_1387,N_810,N_928);
and U1388 (N_1388,N_801,N_1146);
nor U1389 (N_1389,N_1063,N_739);
and U1390 (N_1390,N_1041,N_1125);
nand U1391 (N_1391,N_1165,N_1153);
and U1392 (N_1392,N_905,N_1055);
and U1393 (N_1393,N_1094,N_804);
nor U1394 (N_1394,N_606,N_662);
nor U1395 (N_1395,N_790,N_724);
and U1396 (N_1396,N_1101,N_796);
or U1397 (N_1397,N_833,N_767);
or U1398 (N_1398,N_746,N_1180);
or U1399 (N_1399,N_679,N_904);
and U1400 (N_1400,N_1196,N_815);
nor U1401 (N_1401,N_895,N_1183);
and U1402 (N_1402,N_783,N_615);
and U1403 (N_1403,N_955,N_1114);
nand U1404 (N_1404,N_667,N_873);
nor U1405 (N_1405,N_967,N_923);
nand U1406 (N_1406,N_1025,N_669);
or U1407 (N_1407,N_618,N_605);
nand U1408 (N_1408,N_850,N_769);
nor U1409 (N_1409,N_1149,N_1030);
or U1410 (N_1410,N_1091,N_1121);
and U1411 (N_1411,N_1195,N_685);
and U1412 (N_1412,N_1177,N_689);
nor U1413 (N_1413,N_1106,N_1043);
nand U1414 (N_1414,N_632,N_829);
and U1415 (N_1415,N_1113,N_929);
and U1416 (N_1416,N_1124,N_1139);
nor U1417 (N_1417,N_634,N_900);
and U1418 (N_1418,N_818,N_1036);
nor U1419 (N_1419,N_1199,N_1128);
nand U1420 (N_1420,N_1020,N_1009);
nand U1421 (N_1421,N_938,N_1071);
nor U1422 (N_1422,N_803,N_657);
or U1423 (N_1423,N_1100,N_722);
nor U1424 (N_1424,N_1000,N_779);
and U1425 (N_1425,N_821,N_830);
or U1426 (N_1426,N_825,N_718);
or U1427 (N_1427,N_1192,N_1109);
nand U1428 (N_1428,N_668,N_768);
xor U1429 (N_1429,N_957,N_887);
or U1430 (N_1430,N_831,N_1182);
or U1431 (N_1431,N_1147,N_770);
or U1432 (N_1432,N_1198,N_841);
nand U1433 (N_1433,N_1016,N_970);
or U1434 (N_1434,N_856,N_973);
nor U1435 (N_1435,N_1188,N_639);
nor U1436 (N_1436,N_661,N_819);
or U1437 (N_1437,N_863,N_602);
or U1438 (N_1438,N_884,N_805);
nor U1439 (N_1439,N_707,N_864);
or U1440 (N_1440,N_962,N_1126);
nand U1441 (N_1441,N_952,N_953);
xor U1442 (N_1442,N_752,N_1010);
or U1443 (N_1443,N_877,N_714);
or U1444 (N_1444,N_827,N_885);
nand U1445 (N_1445,N_893,N_1019);
and U1446 (N_1446,N_757,N_745);
nor U1447 (N_1447,N_835,N_935);
nand U1448 (N_1448,N_703,N_686);
or U1449 (N_1449,N_888,N_610);
and U1450 (N_1450,N_1067,N_1108);
nor U1451 (N_1451,N_1080,N_709);
nand U1452 (N_1452,N_963,N_1048);
nor U1453 (N_1453,N_654,N_902);
nor U1454 (N_1454,N_1060,N_914);
and U1455 (N_1455,N_1164,N_1130);
and U1456 (N_1456,N_740,N_1193);
nor U1457 (N_1457,N_1012,N_1002);
or U1458 (N_1458,N_766,N_813);
and U1459 (N_1459,N_826,N_1040);
nor U1460 (N_1460,N_913,N_1079);
nor U1461 (N_1461,N_1132,N_1064);
nor U1462 (N_1462,N_1181,N_751);
nand U1463 (N_1463,N_611,N_868);
nor U1464 (N_1464,N_912,N_812);
or U1465 (N_1465,N_628,N_898);
nor U1466 (N_1466,N_1166,N_633);
nor U1467 (N_1467,N_959,N_700);
nand U1468 (N_1468,N_1167,N_1155);
nand U1469 (N_1469,N_688,N_720);
or U1470 (N_1470,N_948,N_814);
or U1471 (N_1471,N_1086,N_636);
nand U1472 (N_1472,N_750,N_787);
and U1473 (N_1473,N_886,N_1085);
or U1474 (N_1474,N_608,N_1110);
and U1475 (N_1475,N_1145,N_934);
and U1476 (N_1476,N_941,N_716);
nor U1477 (N_1477,N_919,N_788);
or U1478 (N_1478,N_1024,N_1027);
or U1479 (N_1479,N_1152,N_1053);
and U1480 (N_1480,N_1078,N_719);
nand U1481 (N_1481,N_1050,N_836);
and U1482 (N_1482,N_930,N_901);
nand U1483 (N_1483,N_734,N_791);
nor U1484 (N_1484,N_848,N_765);
nand U1485 (N_1485,N_1129,N_1051);
xor U1486 (N_1486,N_612,N_651);
or U1487 (N_1487,N_1023,N_642);
nand U1488 (N_1488,N_702,N_637);
or U1489 (N_1489,N_735,N_1032);
nor U1490 (N_1490,N_762,N_658);
nand U1491 (N_1491,N_964,N_1075);
or U1492 (N_1492,N_771,N_776);
and U1493 (N_1493,N_837,N_1184);
nand U1494 (N_1494,N_1148,N_879);
nor U1495 (N_1495,N_625,N_705);
and U1496 (N_1496,N_1069,N_1087);
nor U1497 (N_1497,N_1157,N_674);
nor U1498 (N_1498,N_872,N_968);
or U1499 (N_1499,N_630,N_698);
nand U1500 (N_1500,N_1170,N_1172);
and U1501 (N_1501,N_817,N_1129);
and U1502 (N_1502,N_1040,N_620);
nor U1503 (N_1503,N_879,N_974);
and U1504 (N_1504,N_1064,N_875);
nand U1505 (N_1505,N_614,N_882);
nand U1506 (N_1506,N_1174,N_1078);
or U1507 (N_1507,N_842,N_826);
nor U1508 (N_1508,N_1023,N_672);
and U1509 (N_1509,N_728,N_611);
or U1510 (N_1510,N_734,N_1096);
or U1511 (N_1511,N_958,N_713);
nor U1512 (N_1512,N_1136,N_911);
nor U1513 (N_1513,N_812,N_664);
nor U1514 (N_1514,N_930,N_728);
nand U1515 (N_1515,N_1021,N_922);
or U1516 (N_1516,N_1193,N_949);
xor U1517 (N_1517,N_1150,N_941);
nand U1518 (N_1518,N_966,N_1096);
or U1519 (N_1519,N_1178,N_613);
or U1520 (N_1520,N_847,N_1105);
and U1521 (N_1521,N_699,N_998);
and U1522 (N_1522,N_1147,N_1133);
nand U1523 (N_1523,N_1028,N_874);
and U1524 (N_1524,N_801,N_1182);
or U1525 (N_1525,N_1156,N_842);
nor U1526 (N_1526,N_695,N_818);
or U1527 (N_1527,N_632,N_783);
or U1528 (N_1528,N_952,N_1025);
and U1529 (N_1529,N_747,N_1040);
nor U1530 (N_1530,N_991,N_1151);
nand U1531 (N_1531,N_630,N_1130);
and U1532 (N_1532,N_1051,N_928);
or U1533 (N_1533,N_881,N_1186);
nand U1534 (N_1534,N_1175,N_625);
nand U1535 (N_1535,N_1143,N_717);
or U1536 (N_1536,N_716,N_907);
or U1537 (N_1537,N_813,N_965);
and U1538 (N_1538,N_856,N_711);
nor U1539 (N_1539,N_820,N_991);
or U1540 (N_1540,N_653,N_654);
nand U1541 (N_1541,N_639,N_931);
nor U1542 (N_1542,N_1017,N_832);
nand U1543 (N_1543,N_1172,N_1069);
nor U1544 (N_1544,N_782,N_867);
and U1545 (N_1545,N_744,N_1006);
nand U1546 (N_1546,N_615,N_778);
nor U1547 (N_1547,N_939,N_963);
nand U1548 (N_1548,N_1069,N_845);
and U1549 (N_1549,N_719,N_754);
and U1550 (N_1550,N_1101,N_667);
and U1551 (N_1551,N_1046,N_811);
nand U1552 (N_1552,N_1114,N_966);
nor U1553 (N_1553,N_1020,N_1136);
or U1554 (N_1554,N_968,N_890);
and U1555 (N_1555,N_884,N_1069);
or U1556 (N_1556,N_989,N_1022);
xnor U1557 (N_1557,N_1151,N_833);
or U1558 (N_1558,N_1121,N_1076);
nand U1559 (N_1559,N_1039,N_1032);
or U1560 (N_1560,N_1152,N_1110);
nor U1561 (N_1561,N_1068,N_1181);
and U1562 (N_1562,N_685,N_667);
or U1563 (N_1563,N_838,N_1155);
and U1564 (N_1564,N_1187,N_1063);
and U1565 (N_1565,N_1130,N_734);
or U1566 (N_1566,N_1154,N_913);
nand U1567 (N_1567,N_820,N_846);
nand U1568 (N_1568,N_859,N_862);
nand U1569 (N_1569,N_807,N_682);
nor U1570 (N_1570,N_974,N_707);
or U1571 (N_1571,N_959,N_621);
and U1572 (N_1572,N_1142,N_985);
or U1573 (N_1573,N_861,N_1109);
and U1574 (N_1574,N_926,N_692);
and U1575 (N_1575,N_901,N_684);
nor U1576 (N_1576,N_900,N_888);
or U1577 (N_1577,N_634,N_1060);
or U1578 (N_1578,N_834,N_946);
or U1579 (N_1579,N_888,N_603);
nor U1580 (N_1580,N_1119,N_987);
and U1581 (N_1581,N_850,N_602);
nor U1582 (N_1582,N_825,N_672);
nor U1583 (N_1583,N_665,N_985);
or U1584 (N_1584,N_1035,N_758);
or U1585 (N_1585,N_768,N_624);
nor U1586 (N_1586,N_948,N_1045);
or U1587 (N_1587,N_827,N_751);
nor U1588 (N_1588,N_940,N_751);
xor U1589 (N_1589,N_812,N_618);
nand U1590 (N_1590,N_838,N_1157);
or U1591 (N_1591,N_1114,N_732);
or U1592 (N_1592,N_943,N_1077);
or U1593 (N_1593,N_1155,N_1133);
nand U1594 (N_1594,N_1059,N_738);
and U1595 (N_1595,N_811,N_961);
nor U1596 (N_1596,N_1115,N_973);
nand U1597 (N_1597,N_932,N_764);
or U1598 (N_1598,N_628,N_672);
xnor U1599 (N_1599,N_1121,N_926);
and U1600 (N_1600,N_864,N_744);
and U1601 (N_1601,N_921,N_1027);
nand U1602 (N_1602,N_1033,N_649);
nand U1603 (N_1603,N_966,N_724);
nand U1604 (N_1604,N_834,N_704);
and U1605 (N_1605,N_761,N_1173);
or U1606 (N_1606,N_716,N_1134);
nor U1607 (N_1607,N_640,N_953);
and U1608 (N_1608,N_697,N_734);
nor U1609 (N_1609,N_977,N_965);
or U1610 (N_1610,N_774,N_625);
nand U1611 (N_1611,N_930,N_892);
nor U1612 (N_1612,N_1053,N_653);
xor U1613 (N_1613,N_635,N_920);
or U1614 (N_1614,N_856,N_629);
nor U1615 (N_1615,N_688,N_1006);
nand U1616 (N_1616,N_618,N_749);
and U1617 (N_1617,N_1049,N_1101);
or U1618 (N_1618,N_837,N_1173);
nand U1619 (N_1619,N_961,N_1190);
and U1620 (N_1620,N_759,N_1122);
nor U1621 (N_1621,N_1106,N_677);
nor U1622 (N_1622,N_655,N_708);
and U1623 (N_1623,N_1019,N_1171);
nand U1624 (N_1624,N_989,N_935);
and U1625 (N_1625,N_1107,N_835);
or U1626 (N_1626,N_1051,N_1130);
nor U1627 (N_1627,N_655,N_637);
and U1628 (N_1628,N_969,N_918);
or U1629 (N_1629,N_912,N_756);
nor U1630 (N_1630,N_910,N_614);
and U1631 (N_1631,N_727,N_1117);
or U1632 (N_1632,N_981,N_775);
and U1633 (N_1633,N_1027,N_1134);
and U1634 (N_1634,N_622,N_1078);
nand U1635 (N_1635,N_939,N_1182);
nand U1636 (N_1636,N_1184,N_1003);
or U1637 (N_1637,N_1007,N_976);
nand U1638 (N_1638,N_1090,N_1097);
and U1639 (N_1639,N_893,N_1109);
and U1640 (N_1640,N_780,N_877);
nand U1641 (N_1641,N_944,N_716);
nor U1642 (N_1642,N_790,N_627);
nor U1643 (N_1643,N_817,N_726);
and U1644 (N_1644,N_929,N_977);
and U1645 (N_1645,N_940,N_965);
nand U1646 (N_1646,N_1006,N_935);
and U1647 (N_1647,N_1099,N_1166);
xnor U1648 (N_1648,N_1166,N_1071);
nor U1649 (N_1649,N_926,N_1183);
nand U1650 (N_1650,N_984,N_722);
or U1651 (N_1651,N_1119,N_853);
nand U1652 (N_1652,N_813,N_726);
xor U1653 (N_1653,N_628,N_1080);
or U1654 (N_1654,N_1101,N_656);
and U1655 (N_1655,N_616,N_893);
and U1656 (N_1656,N_1197,N_814);
or U1657 (N_1657,N_666,N_663);
and U1658 (N_1658,N_926,N_1061);
nand U1659 (N_1659,N_897,N_901);
nor U1660 (N_1660,N_789,N_929);
or U1661 (N_1661,N_1010,N_623);
nand U1662 (N_1662,N_1160,N_629);
nand U1663 (N_1663,N_749,N_760);
and U1664 (N_1664,N_1082,N_1132);
nor U1665 (N_1665,N_870,N_880);
and U1666 (N_1666,N_620,N_879);
nand U1667 (N_1667,N_855,N_844);
or U1668 (N_1668,N_1051,N_1012);
nor U1669 (N_1669,N_971,N_685);
nand U1670 (N_1670,N_693,N_869);
nand U1671 (N_1671,N_1043,N_1022);
and U1672 (N_1672,N_853,N_800);
and U1673 (N_1673,N_935,N_995);
and U1674 (N_1674,N_703,N_625);
nand U1675 (N_1675,N_861,N_1068);
nand U1676 (N_1676,N_1104,N_705);
and U1677 (N_1677,N_969,N_972);
nand U1678 (N_1678,N_983,N_645);
and U1679 (N_1679,N_1150,N_840);
or U1680 (N_1680,N_854,N_978);
nor U1681 (N_1681,N_720,N_618);
and U1682 (N_1682,N_1051,N_946);
and U1683 (N_1683,N_820,N_799);
nor U1684 (N_1684,N_761,N_1174);
nor U1685 (N_1685,N_1042,N_1166);
or U1686 (N_1686,N_1101,N_801);
and U1687 (N_1687,N_853,N_609);
nor U1688 (N_1688,N_1118,N_1021);
xor U1689 (N_1689,N_827,N_794);
nor U1690 (N_1690,N_1030,N_709);
nand U1691 (N_1691,N_958,N_1106);
nand U1692 (N_1692,N_823,N_1187);
nor U1693 (N_1693,N_1056,N_1019);
and U1694 (N_1694,N_1048,N_977);
nor U1695 (N_1695,N_728,N_1080);
nor U1696 (N_1696,N_1019,N_1132);
and U1697 (N_1697,N_893,N_1000);
nor U1698 (N_1698,N_948,N_874);
and U1699 (N_1699,N_740,N_649);
nand U1700 (N_1700,N_684,N_616);
and U1701 (N_1701,N_653,N_951);
or U1702 (N_1702,N_760,N_926);
nor U1703 (N_1703,N_847,N_721);
nand U1704 (N_1704,N_1178,N_941);
xor U1705 (N_1705,N_846,N_747);
nand U1706 (N_1706,N_999,N_914);
nand U1707 (N_1707,N_666,N_1089);
nand U1708 (N_1708,N_1071,N_680);
nor U1709 (N_1709,N_1066,N_916);
nor U1710 (N_1710,N_1153,N_1145);
nor U1711 (N_1711,N_880,N_1079);
nand U1712 (N_1712,N_959,N_672);
and U1713 (N_1713,N_911,N_963);
and U1714 (N_1714,N_1134,N_927);
and U1715 (N_1715,N_1040,N_867);
xor U1716 (N_1716,N_758,N_1158);
or U1717 (N_1717,N_843,N_1063);
or U1718 (N_1718,N_1174,N_1074);
nor U1719 (N_1719,N_1027,N_608);
nand U1720 (N_1720,N_665,N_1080);
nand U1721 (N_1721,N_659,N_702);
xnor U1722 (N_1722,N_954,N_757);
nand U1723 (N_1723,N_804,N_1051);
or U1724 (N_1724,N_770,N_1037);
nand U1725 (N_1725,N_854,N_1079);
nor U1726 (N_1726,N_867,N_956);
and U1727 (N_1727,N_763,N_780);
and U1728 (N_1728,N_933,N_720);
nand U1729 (N_1729,N_1173,N_1130);
and U1730 (N_1730,N_815,N_1148);
nor U1731 (N_1731,N_641,N_674);
nand U1732 (N_1732,N_1021,N_984);
nand U1733 (N_1733,N_957,N_982);
nand U1734 (N_1734,N_1153,N_920);
or U1735 (N_1735,N_731,N_913);
or U1736 (N_1736,N_921,N_850);
and U1737 (N_1737,N_1052,N_667);
nand U1738 (N_1738,N_937,N_1130);
and U1739 (N_1739,N_615,N_967);
or U1740 (N_1740,N_864,N_1179);
nand U1741 (N_1741,N_721,N_809);
and U1742 (N_1742,N_1094,N_623);
nor U1743 (N_1743,N_870,N_625);
nand U1744 (N_1744,N_881,N_673);
or U1745 (N_1745,N_864,N_1180);
nor U1746 (N_1746,N_740,N_828);
and U1747 (N_1747,N_642,N_968);
nor U1748 (N_1748,N_1050,N_696);
and U1749 (N_1749,N_1086,N_972);
nand U1750 (N_1750,N_1004,N_961);
and U1751 (N_1751,N_1150,N_647);
or U1752 (N_1752,N_1084,N_703);
nand U1753 (N_1753,N_1050,N_959);
nor U1754 (N_1754,N_958,N_913);
nor U1755 (N_1755,N_827,N_1173);
nand U1756 (N_1756,N_1092,N_1112);
or U1757 (N_1757,N_683,N_1001);
nand U1758 (N_1758,N_1102,N_945);
and U1759 (N_1759,N_1008,N_1116);
or U1760 (N_1760,N_792,N_869);
and U1761 (N_1761,N_1114,N_634);
nor U1762 (N_1762,N_831,N_1114);
or U1763 (N_1763,N_878,N_1100);
nand U1764 (N_1764,N_672,N_1182);
nor U1765 (N_1765,N_1076,N_883);
and U1766 (N_1766,N_1114,N_909);
nor U1767 (N_1767,N_899,N_907);
nand U1768 (N_1768,N_705,N_1050);
nand U1769 (N_1769,N_928,N_988);
and U1770 (N_1770,N_863,N_1198);
or U1771 (N_1771,N_810,N_673);
and U1772 (N_1772,N_1007,N_1154);
and U1773 (N_1773,N_749,N_815);
and U1774 (N_1774,N_604,N_937);
nand U1775 (N_1775,N_883,N_622);
or U1776 (N_1776,N_877,N_680);
and U1777 (N_1777,N_1090,N_1168);
or U1778 (N_1778,N_833,N_956);
xnor U1779 (N_1779,N_681,N_627);
and U1780 (N_1780,N_637,N_1181);
nand U1781 (N_1781,N_932,N_953);
xnor U1782 (N_1782,N_1009,N_1021);
nor U1783 (N_1783,N_1180,N_1086);
and U1784 (N_1784,N_1052,N_957);
nor U1785 (N_1785,N_793,N_1149);
nor U1786 (N_1786,N_1174,N_967);
nor U1787 (N_1787,N_1125,N_1184);
nand U1788 (N_1788,N_1142,N_744);
or U1789 (N_1789,N_992,N_706);
nor U1790 (N_1790,N_1111,N_1028);
nor U1791 (N_1791,N_688,N_759);
nand U1792 (N_1792,N_907,N_806);
nor U1793 (N_1793,N_1104,N_966);
and U1794 (N_1794,N_659,N_716);
or U1795 (N_1795,N_675,N_639);
nor U1796 (N_1796,N_762,N_1127);
nor U1797 (N_1797,N_761,N_1109);
or U1798 (N_1798,N_712,N_1176);
and U1799 (N_1799,N_661,N_1065);
nand U1800 (N_1800,N_1725,N_1733);
nand U1801 (N_1801,N_1221,N_1430);
or U1802 (N_1802,N_1347,N_1653);
nand U1803 (N_1803,N_1525,N_1554);
and U1804 (N_1804,N_1514,N_1569);
or U1805 (N_1805,N_1238,N_1438);
nand U1806 (N_1806,N_1707,N_1295);
and U1807 (N_1807,N_1278,N_1714);
and U1808 (N_1808,N_1216,N_1476);
nor U1809 (N_1809,N_1768,N_1406);
xor U1810 (N_1810,N_1542,N_1510);
and U1811 (N_1811,N_1746,N_1567);
nor U1812 (N_1812,N_1630,N_1582);
nor U1813 (N_1813,N_1572,N_1676);
nand U1814 (N_1814,N_1469,N_1297);
or U1815 (N_1815,N_1645,N_1709);
and U1816 (N_1816,N_1499,N_1609);
or U1817 (N_1817,N_1698,N_1329);
nand U1818 (N_1818,N_1423,N_1454);
or U1819 (N_1819,N_1259,N_1775);
nand U1820 (N_1820,N_1316,N_1282);
nor U1821 (N_1821,N_1710,N_1334);
nor U1822 (N_1822,N_1446,N_1792);
or U1823 (N_1823,N_1659,N_1531);
nand U1824 (N_1824,N_1363,N_1380);
or U1825 (N_1825,N_1234,N_1479);
and U1826 (N_1826,N_1563,N_1581);
and U1827 (N_1827,N_1694,N_1570);
and U1828 (N_1828,N_1658,N_1361);
or U1829 (N_1829,N_1303,N_1566);
and U1830 (N_1830,N_1751,N_1339);
nand U1831 (N_1831,N_1781,N_1599);
or U1832 (N_1832,N_1667,N_1778);
and U1833 (N_1833,N_1706,N_1547);
nand U1834 (N_1834,N_1390,N_1451);
nor U1835 (N_1835,N_1398,N_1712);
nand U1836 (N_1836,N_1298,N_1460);
nor U1837 (N_1837,N_1611,N_1555);
and U1838 (N_1838,N_1413,N_1589);
nand U1839 (N_1839,N_1755,N_1604);
and U1840 (N_1840,N_1578,N_1227);
and U1841 (N_1841,N_1457,N_1513);
or U1842 (N_1842,N_1393,N_1515);
xor U1843 (N_1843,N_1546,N_1317);
nand U1844 (N_1844,N_1719,N_1729);
nand U1845 (N_1845,N_1565,N_1439);
nand U1846 (N_1846,N_1528,N_1418);
nand U1847 (N_1847,N_1375,N_1557);
and U1848 (N_1848,N_1587,N_1402);
nor U1849 (N_1849,N_1664,N_1759);
nor U1850 (N_1850,N_1232,N_1201);
and U1851 (N_1851,N_1274,N_1241);
nand U1852 (N_1852,N_1315,N_1761);
nor U1853 (N_1853,N_1629,N_1279);
or U1854 (N_1854,N_1202,N_1374);
nor U1855 (N_1855,N_1256,N_1247);
and U1856 (N_1856,N_1715,N_1656);
and U1857 (N_1857,N_1388,N_1560);
nand U1858 (N_1858,N_1319,N_1779);
or U1859 (N_1859,N_1230,N_1226);
and U1860 (N_1860,N_1491,N_1307);
or U1861 (N_1861,N_1562,N_1532);
nand U1862 (N_1862,N_1678,N_1214);
nand U1863 (N_1863,N_1647,N_1516);
and U1864 (N_1864,N_1386,N_1379);
nor U1865 (N_1865,N_1639,N_1467);
or U1866 (N_1866,N_1313,N_1591);
nand U1867 (N_1867,N_1748,N_1475);
nand U1868 (N_1868,N_1553,N_1441);
and U1869 (N_1869,N_1449,N_1357);
nand U1870 (N_1870,N_1291,N_1595);
nand U1871 (N_1871,N_1621,N_1747);
or U1872 (N_1872,N_1428,N_1697);
or U1873 (N_1873,N_1321,N_1354);
nor U1874 (N_1874,N_1593,N_1233);
nand U1875 (N_1875,N_1253,N_1634);
nor U1876 (N_1876,N_1383,N_1713);
and U1877 (N_1877,N_1257,N_1576);
and U1878 (N_1878,N_1246,N_1612);
xnor U1879 (N_1879,N_1767,N_1605);
or U1880 (N_1880,N_1580,N_1482);
nand U1881 (N_1881,N_1346,N_1338);
or U1882 (N_1882,N_1682,N_1500);
or U1883 (N_1883,N_1240,N_1262);
or U1884 (N_1884,N_1498,N_1483);
nand U1885 (N_1885,N_1675,N_1704);
or U1886 (N_1886,N_1702,N_1537);
nand U1887 (N_1887,N_1738,N_1267);
and U1888 (N_1888,N_1336,N_1323);
and U1889 (N_1889,N_1584,N_1462);
nor U1890 (N_1890,N_1403,N_1573);
and U1891 (N_1891,N_1623,N_1265);
nor U1892 (N_1892,N_1743,N_1251);
nand U1893 (N_1893,N_1695,N_1327);
nand U1894 (N_1894,N_1447,N_1250);
and U1895 (N_1895,N_1765,N_1261);
nand U1896 (N_1896,N_1348,N_1741);
nor U1897 (N_1897,N_1795,N_1368);
xnor U1898 (N_1898,N_1534,N_1213);
or U1899 (N_1899,N_1501,N_1300);
nor U1900 (N_1900,N_1540,N_1223);
nor U1901 (N_1901,N_1583,N_1597);
xor U1902 (N_1902,N_1495,N_1679);
nor U1903 (N_1903,N_1649,N_1521);
and U1904 (N_1904,N_1480,N_1381);
nor U1905 (N_1905,N_1377,N_1674);
nor U1906 (N_1906,N_1236,N_1364);
and U1907 (N_1907,N_1436,N_1774);
nand U1908 (N_1908,N_1742,N_1598);
or U1909 (N_1909,N_1669,N_1416);
and U1910 (N_1910,N_1688,N_1400);
or U1911 (N_1911,N_1477,N_1756);
and U1912 (N_1912,N_1425,N_1696);
or U1913 (N_1913,N_1620,N_1592);
nor U1914 (N_1914,N_1640,N_1536);
nor U1915 (N_1915,N_1509,N_1399);
nor U1916 (N_1916,N_1613,N_1520);
nand U1917 (N_1917,N_1244,N_1737);
nand U1918 (N_1918,N_1208,N_1788);
nand U1919 (N_1919,N_1296,N_1507);
and U1920 (N_1920,N_1376,N_1369);
nand U1921 (N_1921,N_1796,N_1248);
and U1922 (N_1922,N_1395,N_1458);
and U1923 (N_1923,N_1526,N_1654);
and U1924 (N_1924,N_1341,N_1235);
nand U1925 (N_1925,N_1200,N_1732);
or U1926 (N_1926,N_1284,N_1750);
nand U1927 (N_1927,N_1522,N_1692);
and U1928 (N_1928,N_1220,N_1686);
and U1929 (N_1929,N_1342,N_1269);
nand U1930 (N_1930,N_1299,N_1760);
or U1931 (N_1931,N_1443,N_1275);
nand U1932 (N_1932,N_1419,N_1485);
nor U1933 (N_1933,N_1217,N_1543);
nor U1934 (N_1934,N_1797,N_1739);
or U1935 (N_1935,N_1780,N_1670);
nor U1936 (N_1936,N_1496,N_1266);
or U1937 (N_1937,N_1212,N_1799);
or U1938 (N_1938,N_1655,N_1429);
or U1939 (N_1939,N_1735,N_1632);
nor U1940 (N_1940,N_1207,N_1219);
nor U1941 (N_1941,N_1332,N_1585);
nand U1942 (N_1942,N_1396,N_1616);
nor U1943 (N_1943,N_1740,N_1505);
nor U1944 (N_1944,N_1545,N_1685);
nor U1945 (N_1945,N_1225,N_1359);
and U1946 (N_1946,N_1360,N_1415);
nand U1947 (N_1947,N_1401,N_1312);
nor U1948 (N_1948,N_1619,N_1677);
and U1949 (N_1949,N_1478,N_1417);
nand U1950 (N_1950,N_1681,N_1577);
or U1951 (N_1951,N_1356,N_1318);
nand U1952 (N_1952,N_1340,N_1785);
or U1953 (N_1953,N_1331,N_1437);
nor U1954 (N_1954,N_1744,N_1245);
and U1955 (N_1955,N_1412,N_1610);
and U1956 (N_1956,N_1204,N_1272);
nand U1957 (N_1957,N_1766,N_1504);
or U1958 (N_1958,N_1481,N_1717);
and U1959 (N_1959,N_1487,N_1210);
nor U1960 (N_1960,N_1209,N_1518);
or U1961 (N_1961,N_1716,N_1503);
and U1962 (N_1962,N_1731,N_1636);
or U1963 (N_1963,N_1783,N_1445);
or U1964 (N_1964,N_1493,N_1322);
nor U1965 (N_1965,N_1358,N_1464);
and U1966 (N_1966,N_1793,N_1607);
nor U1967 (N_1967,N_1290,N_1459);
nor U1968 (N_1968,N_1535,N_1730);
or U1969 (N_1969,N_1672,N_1391);
and U1970 (N_1970,N_1588,N_1407);
nor U1971 (N_1971,N_1648,N_1601);
nand U1972 (N_1972,N_1237,N_1628);
nor U1973 (N_1973,N_1263,N_1764);
and U1974 (N_1974,N_1461,N_1351);
or U1975 (N_1975,N_1753,N_1600);
nand U1976 (N_1976,N_1661,N_1494);
and U1977 (N_1977,N_1260,N_1289);
or U1978 (N_1978,N_1635,N_1422);
nor U1979 (N_1979,N_1352,N_1723);
and U1980 (N_1980,N_1693,N_1517);
nand U1981 (N_1981,N_1281,N_1708);
nand U1982 (N_1982,N_1414,N_1470);
and U1983 (N_1983,N_1328,N_1367);
and U1984 (N_1984,N_1242,N_1224);
xor U1985 (N_1985,N_1426,N_1524);
nor U1986 (N_1986,N_1294,N_1718);
or U1987 (N_1987,N_1206,N_1662);
nor U1988 (N_1988,N_1758,N_1471);
or U1989 (N_1989,N_1727,N_1721);
nor U1990 (N_1990,N_1343,N_1657);
or U1991 (N_1991,N_1466,N_1456);
or U1992 (N_1992,N_1699,N_1633);
and U1993 (N_1993,N_1763,N_1455);
nor U1994 (N_1994,N_1448,N_1752);
nor U1995 (N_1995,N_1355,N_1489);
and U1996 (N_1996,N_1310,N_1397);
nand U1997 (N_1997,N_1651,N_1666);
or U1998 (N_1998,N_1782,N_1231);
nand U1999 (N_1999,N_1798,N_1405);
nand U2000 (N_2000,N_1288,N_1408);
or U2001 (N_2001,N_1450,N_1335);
nor U2002 (N_2002,N_1726,N_1722);
or U2003 (N_2003,N_1472,N_1435);
nand U2004 (N_2004,N_1293,N_1365);
nor U2005 (N_2005,N_1794,N_1353);
or U2006 (N_2006,N_1683,N_1549);
nor U2007 (N_2007,N_1215,N_1789);
nor U2008 (N_2008,N_1421,N_1638);
nand U2009 (N_2009,N_1434,N_1680);
nor U2010 (N_2010,N_1652,N_1301);
and U2011 (N_2011,N_1473,N_1684);
or U2012 (N_2012,N_1787,N_1631);
nand U2013 (N_2013,N_1529,N_1304);
or U2014 (N_2014,N_1497,N_1508);
and U2015 (N_2015,N_1302,N_1308);
or U2016 (N_2016,N_1370,N_1575);
nor U2017 (N_2017,N_1325,N_1689);
nand U2018 (N_2018,N_1218,N_1387);
xor U2019 (N_2019,N_1427,N_1410);
nand U2020 (N_2020,N_1625,N_1326);
nand U2021 (N_2021,N_1637,N_1384);
and U2022 (N_2022,N_1530,N_1615);
or U2023 (N_2023,N_1527,N_1488);
and U2024 (N_2024,N_1552,N_1571);
nor U2025 (N_2025,N_1453,N_1349);
nor U2026 (N_2026,N_1564,N_1734);
nor U2027 (N_2027,N_1286,N_1512);
nand U2028 (N_2028,N_1541,N_1641);
or U2029 (N_2029,N_1784,N_1728);
and U2030 (N_2030,N_1770,N_1550);
or U2031 (N_2031,N_1345,N_1618);
nor U2032 (N_2032,N_1791,N_1392);
nor U2033 (N_2033,N_1490,N_1691);
nand U2034 (N_2034,N_1724,N_1586);
nand U2035 (N_2035,N_1603,N_1424);
or U2036 (N_2036,N_1608,N_1394);
or U2037 (N_2037,N_1650,N_1558);
nand U2038 (N_2038,N_1506,N_1701);
and U2039 (N_2039,N_1665,N_1452);
nor U2040 (N_2040,N_1333,N_1773);
xnor U2041 (N_2041,N_1320,N_1222);
or U2042 (N_2042,N_1720,N_1642);
nand U2043 (N_2043,N_1762,N_1433);
and U2044 (N_2044,N_1502,N_1273);
nand U2045 (N_2045,N_1382,N_1249);
nand U2046 (N_2046,N_1769,N_1551);
or U2047 (N_2047,N_1468,N_1538);
nand U2048 (N_2048,N_1306,N_1486);
nand U2049 (N_2049,N_1745,N_1411);
or U2050 (N_2050,N_1736,N_1372);
nor U2051 (N_2051,N_1703,N_1646);
and U2052 (N_2052,N_1757,N_1602);
and U2053 (N_2053,N_1559,N_1644);
nor U2054 (N_2054,N_1484,N_1442);
or U2055 (N_2055,N_1283,N_1252);
and U2056 (N_2056,N_1432,N_1314);
xor U2057 (N_2057,N_1671,N_1568);
xnor U2058 (N_2058,N_1690,N_1627);
nand U2059 (N_2059,N_1211,N_1790);
nor U2060 (N_2060,N_1277,N_1492);
nand U2061 (N_2061,N_1705,N_1371);
nor U2062 (N_2062,N_1548,N_1373);
or U2063 (N_2063,N_1431,N_1556);
nor U2064 (N_2064,N_1594,N_1378);
or U2065 (N_2065,N_1624,N_1660);
and U2066 (N_2066,N_1440,N_1389);
or U2067 (N_2067,N_1687,N_1229);
and U2068 (N_2068,N_1749,N_1366);
nand U2069 (N_2069,N_1772,N_1561);
or U2070 (N_2070,N_1255,N_1771);
or U2071 (N_2071,N_1617,N_1776);
nand U2072 (N_2072,N_1544,N_1754);
and U2073 (N_2073,N_1404,N_1385);
xnor U2074 (N_2074,N_1474,N_1264);
xnor U2075 (N_2075,N_1324,N_1673);
or U2076 (N_2076,N_1519,N_1668);
and U2077 (N_2077,N_1596,N_1539);
or U2078 (N_2078,N_1463,N_1614);
nor U2079 (N_2079,N_1574,N_1330);
nand U2080 (N_2080,N_1465,N_1523);
or U2081 (N_2081,N_1228,N_1786);
and U2082 (N_2082,N_1420,N_1663);
or U2083 (N_2083,N_1280,N_1344);
or U2084 (N_2084,N_1203,N_1622);
and U2085 (N_2085,N_1606,N_1777);
and U2086 (N_2086,N_1337,N_1292);
nor U2087 (N_2087,N_1311,N_1579);
and U2088 (N_2088,N_1239,N_1285);
nand U2089 (N_2089,N_1205,N_1511);
or U2090 (N_2090,N_1643,N_1711);
and U2091 (N_2091,N_1254,N_1287);
nand U2092 (N_2092,N_1409,N_1268);
or U2093 (N_2093,N_1258,N_1533);
or U2094 (N_2094,N_1243,N_1700);
or U2095 (N_2095,N_1362,N_1270);
nand U2096 (N_2096,N_1309,N_1305);
and U2097 (N_2097,N_1350,N_1276);
or U2098 (N_2098,N_1271,N_1590);
or U2099 (N_2099,N_1444,N_1626);
and U2100 (N_2100,N_1631,N_1373);
nand U2101 (N_2101,N_1568,N_1546);
nor U2102 (N_2102,N_1503,N_1276);
or U2103 (N_2103,N_1390,N_1730);
nand U2104 (N_2104,N_1577,N_1329);
nor U2105 (N_2105,N_1689,N_1557);
nand U2106 (N_2106,N_1549,N_1244);
or U2107 (N_2107,N_1471,N_1274);
and U2108 (N_2108,N_1524,N_1611);
and U2109 (N_2109,N_1312,N_1617);
nand U2110 (N_2110,N_1392,N_1278);
and U2111 (N_2111,N_1401,N_1648);
or U2112 (N_2112,N_1402,N_1782);
or U2113 (N_2113,N_1484,N_1478);
nor U2114 (N_2114,N_1233,N_1299);
nor U2115 (N_2115,N_1412,N_1648);
nor U2116 (N_2116,N_1330,N_1788);
and U2117 (N_2117,N_1260,N_1582);
xnor U2118 (N_2118,N_1513,N_1514);
or U2119 (N_2119,N_1329,N_1425);
nor U2120 (N_2120,N_1524,N_1769);
nor U2121 (N_2121,N_1717,N_1355);
and U2122 (N_2122,N_1763,N_1276);
and U2123 (N_2123,N_1732,N_1351);
and U2124 (N_2124,N_1270,N_1208);
or U2125 (N_2125,N_1394,N_1256);
and U2126 (N_2126,N_1609,N_1753);
xor U2127 (N_2127,N_1352,N_1319);
xnor U2128 (N_2128,N_1495,N_1537);
or U2129 (N_2129,N_1379,N_1248);
nand U2130 (N_2130,N_1565,N_1620);
or U2131 (N_2131,N_1452,N_1610);
xnor U2132 (N_2132,N_1766,N_1791);
or U2133 (N_2133,N_1224,N_1383);
and U2134 (N_2134,N_1792,N_1584);
or U2135 (N_2135,N_1785,N_1454);
and U2136 (N_2136,N_1795,N_1745);
or U2137 (N_2137,N_1724,N_1247);
and U2138 (N_2138,N_1480,N_1248);
and U2139 (N_2139,N_1692,N_1770);
or U2140 (N_2140,N_1543,N_1248);
nand U2141 (N_2141,N_1693,N_1289);
or U2142 (N_2142,N_1447,N_1479);
nand U2143 (N_2143,N_1763,N_1777);
and U2144 (N_2144,N_1362,N_1611);
nand U2145 (N_2145,N_1636,N_1787);
nor U2146 (N_2146,N_1771,N_1428);
or U2147 (N_2147,N_1370,N_1413);
or U2148 (N_2148,N_1693,N_1473);
or U2149 (N_2149,N_1651,N_1699);
xnor U2150 (N_2150,N_1379,N_1351);
and U2151 (N_2151,N_1299,N_1672);
nand U2152 (N_2152,N_1609,N_1304);
nor U2153 (N_2153,N_1245,N_1473);
or U2154 (N_2154,N_1250,N_1511);
nor U2155 (N_2155,N_1275,N_1302);
nand U2156 (N_2156,N_1686,N_1638);
and U2157 (N_2157,N_1302,N_1459);
nor U2158 (N_2158,N_1576,N_1205);
and U2159 (N_2159,N_1471,N_1219);
nor U2160 (N_2160,N_1415,N_1759);
nand U2161 (N_2161,N_1727,N_1582);
nand U2162 (N_2162,N_1436,N_1549);
nand U2163 (N_2163,N_1545,N_1402);
or U2164 (N_2164,N_1438,N_1761);
nand U2165 (N_2165,N_1575,N_1376);
nand U2166 (N_2166,N_1737,N_1652);
nand U2167 (N_2167,N_1290,N_1215);
xor U2168 (N_2168,N_1266,N_1241);
and U2169 (N_2169,N_1600,N_1233);
and U2170 (N_2170,N_1408,N_1459);
nor U2171 (N_2171,N_1374,N_1694);
nor U2172 (N_2172,N_1342,N_1344);
xor U2173 (N_2173,N_1456,N_1610);
or U2174 (N_2174,N_1688,N_1236);
xor U2175 (N_2175,N_1348,N_1639);
nor U2176 (N_2176,N_1349,N_1623);
nor U2177 (N_2177,N_1796,N_1653);
and U2178 (N_2178,N_1394,N_1516);
nor U2179 (N_2179,N_1447,N_1348);
nor U2180 (N_2180,N_1335,N_1370);
nand U2181 (N_2181,N_1495,N_1556);
and U2182 (N_2182,N_1547,N_1556);
or U2183 (N_2183,N_1788,N_1582);
nand U2184 (N_2184,N_1307,N_1259);
and U2185 (N_2185,N_1519,N_1714);
nand U2186 (N_2186,N_1565,N_1773);
nor U2187 (N_2187,N_1488,N_1390);
and U2188 (N_2188,N_1793,N_1515);
or U2189 (N_2189,N_1439,N_1491);
nor U2190 (N_2190,N_1260,N_1647);
nand U2191 (N_2191,N_1425,N_1605);
nand U2192 (N_2192,N_1789,N_1446);
xor U2193 (N_2193,N_1605,N_1596);
nand U2194 (N_2194,N_1406,N_1246);
nand U2195 (N_2195,N_1596,N_1675);
nand U2196 (N_2196,N_1528,N_1473);
and U2197 (N_2197,N_1652,N_1698);
nand U2198 (N_2198,N_1621,N_1304);
and U2199 (N_2199,N_1412,N_1342);
and U2200 (N_2200,N_1546,N_1653);
and U2201 (N_2201,N_1383,N_1500);
nand U2202 (N_2202,N_1632,N_1423);
nor U2203 (N_2203,N_1462,N_1206);
or U2204 (N_2204,N_1425,N_1686);
nand U2205 (N_2205,N_1568,N_1663);
nand U2206 (N_2206,N_1796,N_1249);
or U2207 (N_2207,N_1353,N_1533);
nor U2208 (N_2208,N_1749,N_1758);
or U2209 (N_2209,N_1358,N_1720);
and U2210 (N_2210,N_1751,N_1633);
nand U2211 (N_2211,N_1255,N_1730);
nor U2212 (N_2212,N_1454,N_1531);
or U2213 (N_2213,N_1505,N_1644);
and U2214 (N_2214,N_1780,N_1308);
nand U2215 (N_2215,N_1381,N_1529);
or U2216 (N_2216,N_1291,N_1651);
nor U2217 (N_2217,N_1219,N_1681);
or U2218 (N_2218,N_1398,N_1519);
nor U2219 (N_2219,N_1587,N_1303);
nand U2220 (N_2220,N_1506,N_1278);
nor U2221 (N_2221,N_1227,N_1209);
or U2222 (N_2222,N_1660,N_1678);
and U2223 (N_2223,N_1308,N_1455);
nor U2224 (N_2224,N_1393,N_1562);
and U2225 (N_2225,N_1563,N_1409);
nand U2226 (N_2226,N_1722,N_1619);
nor U2227 (N_2227,N_1518,N_1540);
and U2228 (N_2228,N_1412,N_1304);
nor U2229 (N_2229,N_1277,N_1681);
nand U2230 (N_2230,N_1688,N_1541);
nor U2231 (N_2231,N_1713,N_1529);
or U2232 (N_2232,N_1610,N_1736);
or U2233 (N_2233,N_1562,N_1733);
nor U2234 (N_2234,N_1473,N_1568);
and U2235 (N_2235,N_1464,N_1614);
or U2236 (N_2236,N_1694,N_1407);
and U2237 (N_2237,N_1796,N_1555);
and U2238 (N_2238,N_1310,N_1430);
or U2239 (N_2239,N_1511,N_1271);
or U2240 (N_2240,N_1437,N_1472);
nand U2241 (N_2241,N_1421,N_1630);
or U2242 (N_2242,N_1770,N_1512);
and U2243 (N_2243,N_1504,N_1365);
nand U2244 (N_2244,N_1623,N_1526);
and U2245 (N_2245,N_1395,N_1390);
xor U2246 (N_2246,N_1216,N_1745);
nor U2247 (N_2247,N_1642,N_1292);
nand U2248 (N_2248,N_1407,N_1427);
nor U2249 (N_2249,N_1342,N_1231);
and U2250 (N_2250,N_1470,N_1507);
or U2251 (N_2251,N_1545,N_1627);
nand U2252 (N_2252,N_1497,N_1715);
and U2253 (N_2253,N_1729,N_1541);
nor U2254 (N_2254,N_1708,N_1719);
nand U2255 (N_2255,N_1689,N_1233);
or U2256 (N_2256,N_1418,N_1640);
and U2257 (N_2257,N_1544,N_1385);
or U2258 (N_2258,N_1523,N_1789);
and U2259 (N_2259,N_1279,N_1369);
nand U2260 (N_2260,N_1737,N_1231);
nand U2261 (N_2261,N_1761,N_1509);
and U2262 (N_2262,N_1601,N_1433);
and U2263 (N_2263,N_1464,N_1495);
or U2264 (N_2264,N_1748,N_1352);
xnor U2265 (N_2265,N_1235,N_1382);
and U2266 (N_2266,N_1522,N_1298);
or U2267 (N_2267,N_1734,N_1448);
nand U2268 (N_2268,N_1421,N_1764);
and U2269 (N_2269,N_1452,N_1220);
or U2270 (N_2270,N_1420,N_1452);
nor U2271 (N_2271,N_1780,N_1572);
or U2272 (N_2272,N_1646,N_1348);
or U2273 (N_2273,N_1572,N_1294);
or U2274 (N_2274,N_1243,N_1310);
and U2275 (N_2275,N_1215,N_1422);
nand U2276 (N_2276,N_1224,N_1757);
and U2277 (N_2277,N_1742,N_1655);
and U2278 (N_2278,N_1416,N_1689);
nand U2279 (N_2279,N_1721,N_1481);
xor U2280 (N_2280,N_1526,N_1693);
nor U2281 (N_2281,N_1342,N_1716);
xnor U2282 (N_2282,N_1505,N_1440);
nor U2283 (N_2283,N_1530,N_1278);
or U2284 (N_2284,N_1683,N_1483);
nand U2285 (N_2285,N_1217,N_1643);
or U2286 (N_2286,N_1287,N_1479);
nor U2287 (N_2287,N_1221,N_1292);
nand U2288 (N_2288,N_1448,N_1668);
and U2289 (N_2289,N_1770,N_1441);
nand U2290 (N_2290,N_1235,N_1466);
and U2291 (N_2291,N_1584,N_1564);
nand U2292 (N_2292,N_1623,N_1603);
nor U2293 (N_2293,N_1272,N_1335);
or U2294 (N_2294,N_1275,N_1284);
and U2295 (N_2295,N_1425,N_1741);
nand U2296 (N_2296,N_1764,N_1322);
or U2297 (N_2297,N_1266,N_1242);
or U2298 (N_2298,N_1596,N_1613);
nor U2299 (N_2299,N_1727,N_1341);
nor U2300 (N_2300,N_1723,N_1451);
xnor U2301 (N_2301,N_1305,N_1673);
nor U2302 (N_2302,N_1316,N_1694);
nand U2303 (N_2303,N_1500,N_1794);
nor U2304 (N_2304,N_1490,N_1232);
and U2305 (N_2305,N_1703,N_1285);
xor U2306 (N_2306,N_1548,N_1728);
or U2307 (N_2307,N_1222,N_1565);
or U2308 (N_2308,N_1390,N_1701);
nand U2309 (N_2309,N_1717,N_1395);
nand U2310 (N_2310,N_1238,N_1794);
or U2311 (N_2311,N_1363,N_1473);
nor U2312 (N_2312,N_1796,N_1339);
nand U2313 (N_2313,N_1580,N_1624);
nor U2314 (N_2314,N_1207,N_1774);
and U2315 (N_2315,N_1358,N_1717);
and U2316 (N_2316,N_1248,N_1651);
nor U2317 (N_2317,N_1713,N_1395);
or U2318 (N_2318,N_1574,N_1414);
and U2319 (N_2319,N_1255,N_1657);
nand U2320 (N_2320,N_1627,N_1482);
or U2321 (N_2321,N_1291,N_1422);
or U2322 (N_2322,N_1289,N_1538);
nor U2323 (N_2323,N_1290,N_1752);
nand U2324 (N_2324,N_1450,N_1438);
xor U2325 (N_2325,N_1689,N_1441);
xnor U2326 (N_2326,N_1373,N_1300);
nor U2327 (N_2327,N_1218,N_1301);
nor U2328 (N_2328,N_1651,N_1284);
or U2329 (N_2329,N_1241,N_1211);
nor U2330 (N_2330,N_1510,N_1753);
and U2331 (N_2331,N_1373,N_1297);
and U2332 (N_2332,N_1490,N_1733);
xor U2333 (N_2333,N_1575,N_1432);
and U2334 (N_2334,N_1611,N_1248);
nand U2335 (N_2335,N_1505,N_1518);
and U2336 (N_2336,N_1314,N_1242);
nand U2337 (N_2337,N_1205,N_1480);
nand U2338 (N_2338,N_1695,N_1678);
or U2339 (N_2339,N_1767,N_1789);
and U2340 (N_2340,N_1430,N_1329);
and U2341 (N_2341,N_1744,N_1389);
nand U2342 (N_2342,N_1578,N_1208);
nor U2343 (N_2343,N_1361,N_1469);
or U2344 (N_2344,N_1421,N_1375);
and U2345 (N_2345,N_1250,N_1363);
and U2346 (N_2346,N_1268,N_1567);
or U2347 (N_2347,N_1283,N_1203);
nand U2348 (N_2348,N_1437,N_1496);
or U2349 (N_2349,N_1580,N_1504);
nand U2350 (N_2350,N_1414,N_1334);
nand U2351 (N_2351,N_1477,N_1238);
and U2352 (N_2352,N_1481,N_1584);
nor U2353 (N_2353,N_1730,N_1517);
nand U2354 (N_2354,N_1729,N_1630);
nor U2355 (N_2355,N_1657,N_1267);
or U2356 (N_2356,N_1428,N_1474);
nand U2357 (N_2357,N_1542,N_1319);
or U2358 (N_2358,N_1585,N_1439);
xnor U2359 (N_2359,N_1737,N_1553);
nand U2360 (N_2360,N_1786,N_1624);
or U2361 (N_2361,N_1466,N_1717);
nand U2362 (N_2362,N_1314,N_1675);
and U2363 (N_2363,N_1548,N_1352);
or U2364 (N_2364,N_1529,N_1592);
and U2365 (N_2365,N_1363,N_1324);
and U2366 (N_2366,N_1518,N_1572);
or U2367 (N_2367,N_1609,N_1205);
or U2368 (N_2368,N_1272,N_1461);
nor U2369 (N_2369,N_1218,N_1580);
nand U2370 (N_2370,N_1629,N_1323);
and U2371 (N_2371,N_1219,N_1347);
and U2372 (N_2372,N_1771,N_1515);
nor U2373 (N_2373,N_1437,N_1338);
nand U2374 (N_2374,N_1427,N_1632);
or U2375 (N_2375,N_1333,N_1307);
or U2376 (N_2376,N_1533,N_1709);
and U2377 (N_2377,N_1230,N_1284);
or U2378 (N_2378,N_1549,N_1240);
or U2379 (N_2379,N_1530,N_1757);
and U2380 (N_2380,N_1615,N_1704);
nor U2381 (N_2381,N_1691,N_1721);
xor U2382 (N_2382,N_1638,N_1293);
nand U2383 (N_2383,N_1532,N_1639);
nor U2384 (N_2384,N_1420,N_1403);
and U2385 (N_2385,N_1229,N_1500);
or U2386 (N_2386,N_1668,N_1286);
or U2387 (N_2387,N_1693,N_1246);
and U2388 (N_2388,N_1248,N_1201);
nand U2389 (N_2389,N_1346,N_1701);
or U2390 (N_2390,N_1603,N_1721);
nor U2391 (N_2391,N_1242,N_1414);
nor U2392 (N_2392,N_1485,N_1415);
nor U2393 (N_2393,N_1783,N_1378);
nor U2394 (N_2394,N_1466,N_1288);
or U2395 (N_2395,N_1724,N_1662);
and U2396 (N_2396,N_1303,N_1511);
nor U2397 (N_2397,N_1272,N_1566);
nor U2398 (N_2398,N_1424,N_1737);
nand U2399 (N_2399,N_1633,N_1485);
and U2400 (N_2400,N_2338,N_1830);
nand U2401 (N_2401,N_2084,N_1932);
or U2402 (N_2402,N_1893,N_1850);
or U2403 (N_2403,N_2196,N_2036);
xor U2404 (N_2404,N_2110,N_2058);
or U2405 (N_2405,N_2129,N_1909);
nor U2406 (N_2406,N_2151,N_2096);
and U2407 (N_2407,N_2208,N_2283);
nor U2408 (N_2408,N_1875,N_2279);
or U2409 (N_2409,N_2325,N_2165);
or U2410 (N_2410,N_2008,N_2187);
or U2411 (N_2411,N_2015,N_1877);
and U2412 (N_2412,N_1876,N_2305);
or U2413 (N_2413,N_1966,N_2049);
nand U2414 (N_2414,N_1974,N_1904);
or U2415 (N_2415,N_2194,N_2115);
nand U2416 (N_2416,N_1977,N_1922);
nand U2417 (N_2417,N_2169,N_1996);
and U2418 (N_2418,N_1856,N_2144);
and U2419 (N_2419,N_2260,N_2175);
nand U2420 (N_2420,N_2161,N_2121);
or U2421 (N_2421,N_2163,N_2132);
nand U2422 (N_2422,N_2143,N_2339);
nand U2423 (N_2423,N_1957,N_1835);
and U2424 (N_2424,N_2326,N_2383);
and U2425 (N_2425,N_2287,N_2146);
and U2426 (N_2426,N_1886,N_2251);
or U2427 (N_2427,N_2238,N_1841);
or U2428 (N_2428,N_2263,N_1861);
nor U2429 (N_2429,N_1822,N_2273);
and U2430 (N_2430,N_2226,N_2105);
and U2431 (N_2431,N_2356,N_2253);
nand U2432 (N_2432,N_1895,N_2270);
and U2433 (N_2433,N_2331,N_2302);
xnor U2434 (N_2434,N_1855,N_1865);
or U2435 (N_2435,N_2372,N_2373);
and U2436 (N_2436,N_1839,N_2347);
or U2437 (N_2437,N_1967,N_2241);
or U2438 (N_2438,N_2178,N_2073);
xor U2439 (N_2439,N_2289,N_2098);
or U2440 (N_2440,N_2062,N_2292);
xnor U2441 (N_2441,N_2092,N_2301);
or U2442 (N_2442,N_2224,N_1907);
nand U2443 (N_2443,N_2275,N_2294);
or U2444 (N_2444,N_1829,N_1849);
and U2445 (N_2445,N_2154,N_2141);
nor U2446 (N_2446,N_2274,N_1919);
or U2447 (N_2447,N_2171,N_1845);
nor U2448 (N_2448,N_2136,N_1968);
nor U2449 (N_2449,N_1892,N_1965);
or U2450 (N_2450,N_1964,N_2023);
nor U2451 (N_2451,N_2193,N_1947);
nand U2452 (N_2452,N_1900,N_1874);
nor U2453 (N_2453,N_2079,N_2080);
or U2454 (N_2454,N_2106,N_2052);
or U2455 (N_2455,N_2375,N_2192);
nand U2456 (N_2456,N_1990,N_2320);
or U2457 (N_2457,N_1969,N_1978);
nor U2458 (N_2458,N_1954,N_2004);
and U2459 (N_2459,N_2385,N_1920);
nor U2460 (N_2460,N_2122,N_2116);
nor U2461 (N_2461,N_1834,N_2191);
or U2462 (N_2462,N_2035,N_2231);
nor U2463 (N_2463,N_2139,N_2071);
nand U2464 (N_2464,N_2059,N_2362);
nor U2465 (N_2465,N_2321,N_2236);
and U2466 (N_2466,N_1807,N_2019);
or U2467 (N_2467,N_1883,N_2027);
and U2468 (N_2468,N_1854,N_1981);
and U2469 (N_2469,N_1984,N_2237);
nand U2470 (N_2470,N_2046,N_1831);
or U2471 (N_2471,N_1925,N_2316);
nand U2472 (N_2472,N_2177,N_1993);
nand U2473 (N_2473,N_2162,N_2346);
nor U2474 (N_2474,N_2094,N_2038);
nor U2475 (N_2475,N_2135,N_2097);
xor U2476 (N_2476,N_2366,N_2268);
nand U2477 (N_2477,N_2290,N_1915);
and U2478 (N_2478,N_2202,N_2041);
and U2479 (N_2479,N_2160,N_1847);
nor U2480 (N_2480,N_1924,N_2278);
nand U2481 (N_2481,N_2322,N_2078);
or U2482 (N_2482,N_2009,N_1917);
or U2483 (N_2483,N_2376,N_1837);
nand U2484 (N_2484,N_2343,N_2180);
and U2485 (N_2485,N_1959,N_2262);
or U2486 (N_2486,N_1846,N_2367);
and U2487 (N_2487,N_2342,N_1914);
or U2488 (N_2488,N_2108,N_2361);
and U2489 (N_2489,N_1859,N_2051);
or U2490 (N_2490,N_2209,N_2130);
nand U2491 (N_2491,N_2309,N_2182);
nand U2492 (N_2492,N_2107,N_2179);
or U2493 (N_2493,N_2045,N_2284);
or U2494 (N_2494,N_2155,N_2235);
or U2495 (N_2495,N_1818,N_1802);
and U2496 (N_2496,N_2269,N_1963);
nor U2497 (N_2497,N_1833,N_1811);
xnor U2498 (N_2498,N_2215,N_2308);
nand U2499 (N_2499,N_2174,N_2057);
nor U2500 (N_2500,N_1821,N_2371);
or U2501 (N_2501,N_2088,N_1881);
nor U2502 (N_2502,N_2082,N_2021);
and U2503 (N_2503,N_1897,N_1848);
nor U2504 (N_2504,N_2360,N_2254);
or U2505 (N_2505,N_2124,N_1863);
or U2506 (N_2506,N_1955,N_2296);
nor U2507 (N_2507,N_1819,N_2006);
or U2508 (N_2508,N_2298,N_2333);
and U2509 (N_2509,N_2111,N_1916);
xnor U2510 (N_2510,N_1962,N_2134);
nand U2511 (N_2511,N_2386,N_2276);
nand U2512 (N_2512,N_2195,N_2048);
nand U2513 (N_2513,N_1927,N_1952);
or U2514 (N_2514,N_2377,N_2201);
or U2515 (N_2515,N_2340,N_2355);
or U2516 (N_2516,N_1826,N_2207);
or U2517 (N_2517,N_1878,N_2199);
nand U2518 (N_2518,N_1985,N_2040);
nand U2519 (N_2519,N_2087,N_1888);
nand U2520 (N_2520,N_2173,N_2335);
nor U2521 (N_2521,N_1851,N_2222);
and U2522 (N_2522,N_2148,N_1982);
nand U2523 (N_2523,N_2093,N_1940);
and U2524 (N_2524,N_2299,N_2113);
nand U2525 (N_2525,N_2312,N_1801);
nand U2526 (N_2526,N_2128,N_1972);
and U2527 (N_2527,N_2029,N_1884);
or U2528 (N_2528,N_1971,N_2070);
or U2529 (N_2529,N_2198,N_1987);
nor U2530 (N_2530,N_2095,N_2077);
nand U2531 (N_2531,N_2137,N_1999);
or U2532 (N_2532,N_2227,N_2054);
nor U2533 (N_2533,N_2133,N_2131);
and U2534 (N_2534,N_1827,N_2328);
and U2535 (N_2535,N_1808,N_2145);
nand U2536 (N_2536,N_2086,N_2064);
nor U2537 (N_2537,N_2323,N_2240);
and U2538 (N_2538,N_1857,N_2089);
nor U2539 (N_2539,N_1944,N_2074);
nor U2540 (N_2540,N_2358,N_2280);
and U2541 (N_2541,N_2042,N_2158);
nand U2542 (N_2542,N_1891,N_1896);
nor U2543 (N_2543,N_2076,N_1868);
xnor U2544 (N_2544,N_2315,N_2300);
nor U2545 (N_2545,N_2245,N_1858);
nor U2546 (N_2546,N_2282,N_2239);
and U2547 (N_2547,N_2010,N_1899);
nor U2548 (N_2548,N_2392,N_2181);
nand U2549 (N_2549,N_1997,N_2266);
nor U2550 (N_2550,N_1995,N_2390);
or U2551 (N_2551,N_1803,N_1810);
nor U2552 (N_2552,N_1853,N_2391);
and U2553 (N_2553,N_1843,N_1800);
nor U2554 (N_2554,N_2397,N_1873);
nor U2555 (N_2555,N_2291,N_2104);
nand U2556 (N_2556,N_2243,N_2349);
nand U2557 (N_2557,N_2344,N_1836);
xor U2558 (N_2558,N_1950,N_2306);
nor U2559 (N_2559,N_2055,N_2330);
nand U2560 (N_2560,N_2225,N_2378);
and U2561 (N_2561,N_1946,N_1943);
or U2562 (N_2562,N_1961,N_2069);
nand U2563 (N_2563,N_2153,N_2028);
nand U2564 (N_2564,N_2353,N_2318);
nor U2565 (N_2565,N_2341,N_2384);
and U2566 (N_2566,N_2085,N_1832);
and U2567 (N_2567,N_1816,N_1975);
and U2568 (N_2568,N_1825,N_2037);
or U2569 (N_2569,N_2065,N_2102);
and U2570 (N_2570,N_1934,N_2184);
nand U2571 (N_2571,N_2234,N_2394);
and U2572 (N_2572,N_2230,N_2228);
or U2573 (N_2573,N_2011,N_2003);
or U2574 (N_2574,N_2220,N_1933);
nor U2575 (N_2575,N_2001,N_2067);
nor U2576 (N_2576,N_2063,N_2044);
nand U2577 (N_2577,N_2018,N_2150);
nand U2578 (N_2578,N_2396,N_1989);
or U2579 (N_2579,N_1867,N_2060);
nand U2580 (N_2580,N_2017,N_1806);
xnor U2581 (N_2581,N_2248,N_1882);
nor U2582 (N_2582,N_2295,N_2118);
or U2583 (N_2583,N_2348,N_2311);
or U2584 (N_2584,N_2304,N_2370);
nor U2585 (N_2585,N_2256,N_2217);
or U2586 (N_2586,N_2369,N_1901);
or U2587 (N_2587,N_2101,N_2005);
nor U2588 (N_2588,N_2022,N_1903);
or U2589 (N_2589,N_2219,N_2357);
nand U2590 (N_2590,N_1911,N_2168);
nor U2591 (N_2591,N_2147,N_1828);
nor U2592 (N_2592,N_2152,N_1866);
and U2593 (N_2593,N_2127,N_2364);
nor U2594 (N_2594,N_2281,N_2034);
and U2595 (N_2595,N_2388,N_2066);
nand U2596 (N_2596,N_2258,N_1910);
nand U2597 (N_2597,N_1824,N_2307);
or U2598 (N_2598,N_2100,N_2212);
nand U2599 (N_2599,N_1804,N_2334);
and U2600 (N_2600,N_1926,N_2012);
nor U2601 (N_2601,N_1870,N_2170);
and U2602 (N_2602,N_2117,N_2221);
or U2603 (N_2603,N_2345,N_2250);
nor U2604 (N_2604,N_2172,N_2387);
nand U2605 (N_2605,N_2336,N_2293);
nor U2606 (N_2606,N_1838,N_1872);
nor U2607 (N_2607,N_2368,N_2297);
nor U2608 (N_2608,N_2223,N_1937);
and U2609 (N_2609,N_2024,N_2112);
and U2610 (N_2610,N_2288,N_2310);
and U2611 (N_2611,N_2267,N_1898);
nand U2612 (N_2612,N_2379,N_2083);
and U2613 (N_2613,N_1906,N_1942);
and U2614 (N_2614,N_2025,N_2272);
nand U2615 (N_2615,N_2261,N_2002);
nand U2616 (N_2616,N_2203,N_1936);
nand U2617 (N_2617,N_2047,N_2271);
and U2618 (N_2618,N_2286,N_1953);
or U2619 (N_2619,N_1902,N_1885);
nand U2620 (N_2620,N_1921,N_2026);
nor U2621 (N_2621,N_2014,N_2109);
or U2622 (N_2622,N_2125,N_1844);
xnor U2623 (N_2623,N_1918,N_2313);
or U2624 (N_2624,N_1939,N_2381);
or U2625 (N_2625,N_2061,N_2359);
or U2626 (N_2626,N_2398,N_2213);
nor U2627 (N_2627,N_2099,N_1960);
nor U2628 (N_2628,N_2189,N_1923);
nor U2629 (N_2629,N_2166,N_2159);
and U2630 (N_2630,N_2242,N_2197);
and U2631 (N_2631,N_1871,N_2075);
or U2632 (N_2632,N_1864,N_1887);
nand U2633 (N_2633,N_1820,N_1869);
or U2634 (N_2634,N_2249,N_2186);
nor U2635 (N_2635,N_2264,N_2332);
nand U2636 (N_2636,N_1815,N_2324);
and U2637 (N_2637,N_1912,N_2140);
nor U2638 (N_2638,N_2183,N_1992);
nor U2639 (N_2639,N_2252,N_1941);
nor U2640 (N_2640,N_1945,N_1852);
nand U2641 (N_2641,N_1973,N_2176);
nor U2642 (N_2642,N_2232,N_2016);
or U2643 (N_2643,N_2013,N_1809);
or U2644 (N_2644,N_2142,N_1930);
nand U2645 (N_2645,N_2185,N_2216);
and U2646 (N_2646,N_2229,N_1948);
nand U2647 (N_2647,N_2285,N_2319);
nor U2648 (N_2648,N_1994,N_2380);
and U2649 (N_2649,N_1931,N_2205);
nor U2650 (N_2650,N_2149,N_2218);
or U2651 (N_2651,N_2188,N_2257);
nand U2652 (N_2652,N_1949,N_2114);
and U2653 (N_2653,N_2000,N_2382);
nand U2654 (N_2654,N_2317,N_1814);
and U2655 (N_2655,N_1998,N_2393);
or U2656 (N_2656,N_2206,N_2056);
or U2657 (N_2657,N_2351,N_2157);
or U2658 (N_2658,N_1840,N_2277);
nand U2659 (N_2659,N_1908,N_1983);
nand U2660 (N_2660,N_1988,N_2354);
nand U2661 (N_2661,N_2389,N_2050);
and U2662 (N_2662,N_2399,N_1880);
nand U2663 (N_2663,N_2350,N_2126);
or U2664 (N_2664,N_2265,N_2138);
or U2665 (N_2665,N_1951,N_2081);
or U2666 (N_2666,N_1860,N_1813);
nand U2667 (N_2667,N_1929,N_2204);
xnor U2668 (N_2668,N_2255,N_1913);
nor U2669 (N_2669,N_1817,N_2164);
nand U2670 (N_2670,N_1842,N_2211);
nand U2671 (N_2671,N_2020,N_2032);
nand U2672 (N_2672,N_2337,N_2068);
nand U2673 (N_2673,N_2031,N_1890);
nor U2674 (N_2674,N_2214,N_1980);
or U2675 (N_2675,N_2233,N_2007);
or U2676 (N_2676,N_2210,N_2247);
or U2677 (N_2677,N_2303,N_2365);
nand U2678 (N_2678,N_1958,N_1862);
nor U2679 (N_2679,N_2167,N_1805);
nor U2680 (N_2680,N_2119,N_1905);
or U2681 (N_2681,N_1976,N_2091);
nor U2682 (N_2682,N_1935,N_1894);
nand U2683 (N_2683,N_2090,N_2033);
and U2684 (N_2684,N_2103,N_1889);
nand U2685 (N_2685,N_2329,N_2123);
xor U2686 (N_2686,N_2363,N_2190);
and U2687 (N_2687,N_1956,N_2327);
nand U2688 (N_2688,N_1928,N_1970);
or U2689 (N_2689,N_1986,N_2374);
nand U2690 (N_2690,N_2200,N_1812);
or U2691 (N_2691,N_2030,N_2259);
and U2692 (N_2692,N_2314,N_1938);
nor U2693 (N_2693,N_2246,N_2395);
nor U2694 (N_2694,N_1991,N_1823);
and U2695 (N_2695,N_2120,N_2156);
or U2696 (N_2696,N_2072,N_2352);
nor U2697 (N_2697,N_2043,N_2244);
or U2698 (N_2698,N_2053,N_1879);
nor U2699 (N_2699,N_1979,N_2039);
or U2700 (N_2700,N_2003,N_2177);
or U2701 (N_2701,N_1882,N_1957);
or U2702 (N_2702,N_2007,N_1876);
and U2703 (N_2703,N_1861,N_1848);
xnor U2704 (N_2704,N_1842,N_2285);
or U2705 (N_2705,N_1824,N_2059);
nor U2706 (N_2706,N_2325,N_2006);
or U2707 (N_2707,N_2202,N_1897);
nor U2708 (N_2708,N_2100,N_2010);
nor U2709 (N_2709,N_2134,N_1822);
and U2710 (N_2710,N_1975,N_2243);
and U2711 (N_2711,N_1850,N_2269);
and U2712 (N_2712,N_2134,N_1923);
or U2713 (N_2713,N_1890,N_2149);
nor U2714 (N_2714,N_2085,N_2110);
nand U2715 (N_2715,N_2328,N_2134);
or U2716 (N_2716,N_2295,N_1993);
or U2717 (N_2717,N_2074,N_1997);
and U2718 (N_2718,N_1968,N_1805);
nand U2719 (N_2719,N_2019,N_2040);
or U2720 (N_2720,N_2080,N_2336);
xnor U2721 (N_2721,N_2350,N_1930);
nand U2722 (N_2722,N_1920,N_2234);
and U2723 (N_2723,N_1859,N_2391);
nand U2724 (N_2724,N_2337,N_2368);
nor U2725 (N_2725,N_1940,N_2130);
or U2726 (N_2726,N_2045,N_2181);
and U2727 (N_2727,N_2295,N_2168);
or U2728 (N_2728,N_1813,N_2149);
and U2729 (N_2729,N_2061,N_1808);
nand U2730 (N_2730,N_1884,N_1905);
or U2731 (N_2731,N_1959,N_1917);
or U2732 (N_2732,N_2380,N_1882);
nand U2733 (N_2733,N_2226,N_1947);
xnor U2734 (N_2734,N_2163,N_2342);
and U2735 (N_2735,N_2235,N_1853);
and U2736 (N_2736,N_1999,N_2054);
nand U2737 (N_2737,N_2022,N_2036);
or U2738 (N_2738,N_1829,N_1943);
nor U2739 (N_2739,N_1947,N_2113);
xor U2740 (N_2740,N_2314,N_2392);
nand U2741 (N_2741,N_2117,N_2304);
and U2742 (N_2742,N_2221,N_2371);
nor U2743 (N_2743,N_2292,N_2199);
nor U2744 (N_2744,N_2230,N_2144);
nor U2745 (N_2745,N_1852,N_2159);
and U2746 (N_2746,N_1993,N_1990);
or U2747 (N_2747,N_2178,N_2365);
nand U2748 (N_2748,N_2102,N_2392);
or U2749 (N_2749,N_2243,N_1985);
and U2750 (N_2750,N_2364,N_2150);
nand U2751 (N_2751,N_2239,N_2331);
or U2752 (N_2752,N_1923,N_2339);
nor U2753 (N_2753,N_1805,N_2063);
or U2754 (N_2754,N_2155,N_2288);
or U2755 (N_2755,N_2201,N_1893);
and U2756 (N_2756,N_1976,N_1883);
nor U2757 (N_2757,N_2040,N_1819);
and U2758 (N_2758,N_2358,N_2373);
or U2759 (N_2759,N_2003,N_2341);
nor U2760 (N_2760,N_2390,N_2317);
xor U2761 (N_2761,N_2118,N_2376);
and U2762 (N_2762,N_2275,N_1961);
and U2763 (N_2763,N_1812,N_2160);
nor U2764 (N_2764,N_1941,N_1800);
nand U2765 (N_2765,N_2284,N_1826);
and U2766 (N_2766,N_2339,N_2326);
nor U2767 (N_2767,N_1836,N_2335);
or U2768 (N_2768,N_1951,N_2178);
nand U2769 (N_2769,N_1959,N_2320);
nand U2770 (N_2770,N_2264,N_2072);
nor U2771 (N_2771,N_2114,N_2101);
nand U2772 (N_2772,N_2203,N_2131);
nor U2773 (N_2773,N_2031,N_2350);
and U2774 (N_2774,N_1921,N_2280);
or U2775 (N_2775,N_2140,N_2348);
and U2776 (N_2776,N_1971,N_1991);
nand U2777 (N_2777,N_1892,N_1851);
and U2778 (N_2778,N_1805,N_2392);
or U2779 (N_2779,N_1892,N_2100);
nor U2780 (N_2780,N_2012,N_2224);
nand U2781 (N_2781,N_1851,N_2273);
nand U2782 (N_2782,N_2158,N_2122);
or U2783 (N_2783,N_2069,N_2198);
and U2784 (N_2784,N_2108,N_2119);
or U2785 (N_2785,N_1926,N_2325);
and U2786 (N_2786,N_1940,N_1912);
or U2787 (N_2787,N_2108,N_2237);
and U2788 (N_2788,N_2159,N_2339);
or U2789 (N_2789,N_2244,N_1808);
or U2790 (N_2790,N_1989,N_1970);
nor U2791 (N_2791,N_2029,N_2375);
nor U2792 (N_2792,N_2291,N_1858);
nor U2793 (N_2793,N_1932,N_1870);
or U2794 (N_2794,N_2139,N_2060);
nor U2795 (N_2795,N_2337,N_1847);
nand U2796 (N_2796,N_1856,N_2115);
and U2797 (N_2797,N_1883,N_2107);
nor U2798 (N_2798,N_2104,N_1859);
nand U2799 (N_2799,N_2297,N_2299);
and U2800 (N_2800,N_2345,N_2119);
nor U2801 (N_2801,N_1931,N_2311);
xnor U2802 (N_2802,N_2196,N_2080);
and U2803 (N_2803,N_2015,N_2008);
nand U2804 (N_2804,N_2008,N_1880);
and U2805 (N_2805,N_1894,N_2362);
or U2806 (N_2806,N_1863,N_2157);
and U2807 (N_2807,N_2276,N_2274);
or U2808 (N_2808,N_1963,N_1929);
and U2809 (N_2809,N_2161,N_2226);
nor U2810 (N_2810,N_2042,N_2224);
nand U2811 (N_2811,N_1934,N_2050);
nand U2812 (N_2812,N_1978,N_2133);
or U2813 (N_2813,N_1866,N_1951);
and U2814 (N_2814,N_2190,N_1861);
and U2815 (N_2815,N_2246,N_1962);
or U2816 (N_2816,N_2204,N_2313);
and U2817 (N_2817,N_2270,N_2030);
nor U2818 (N_2818,N_2337,N_2367);
and U2819 (N_2819,N_2197,N_2087);
and U2820 (N_2820,N_2261,N_2151);
and U2821 (N_2821,N_2077,N_1954);
or U2822 (N_2822,N_1901,N_2342);
nand U2823 (N_2823,N_1848,N_1984);
or U2824 (N_2824,N_2385,N_1981);
or U2825 (N_2825,N_2105,N_2193);
xnor U2826 (N_2826,N_1841,N_2020);
and U2827 (N_2827,N_1831,N_1952);
or U2828 (N_2828,N_2039,N_1945);
nand U2829 (N_2829,N_2006,N_2357);
or U2830 (N_2830,N_1876,N_2129);
and U2831 (N_2831,N_1898,N_2076);
xnor U2832 (N_2832,N_1972,N_2067);
nor U2833 (N_2833,N_2357,N_1869);
or U2834 (N_2834,N_2004,N_2025);
or U2835 (N_2835,N_2285,N_2216);
xor U2836 (N_2836,N_1991,N_1908);
nor U2837 (N_2837,N_2243,N_2236);
nand U2838 (N_2838,N_2297,N_2259);
and U2839 (N_2839,N_2113,N_1943);
and U2840 (N_2840,N_2080,N_2153);
nor U2841 (N_2841,N_2221,N_1966);
nor U2842 (N_2842,N_2363,N_1905);
nand U2843 (N_2843,N_2186,N_1831);
nand U2844 (N_2844,N_2303,N_2248);
xor U2845 (N_2845,N_1994,N_1967);
nand U2846 (N_2846,N_2222,N_2277);
nor U2847 (N_2847,N_2207,N_1940);
xor U2848 (N_2848,N_2033,N_2012);
or U2849 (N_2849,N_2198,N_2101);
nand U2850 (N_2850,N_2194,N_1899);
nor U2851 (N_2851,N_2116,N_1867);
nor U2852 (N_2852,N_1806,N_1924);
nand U2853 (N_2853,N_1994,N_2000);
and U2854 (N_2854,N_2380,N_2306);
and U2855 (N_2855,N_2264,N_2183);
or U2856 (N_2856,N_2062,N_2181);
nor U2857 (N_2857,N_1967,N_1863);
or U2858 (N_2858,N_2210,N_1820);
nor U2859 (N_2859,N_2055,N_1811);
nor U2860 (N_2860,N_1868,N_2391);
nor U2861 (N_2861,N_2197,N_2264);
or U2862 (N_2862,N_2105,N_2065);
nor U2863 (N_2863,N_2189,N_2365);
nor U2864 (N_2864,N_2209,N_1971);
or U2865 (N_2865,N_2101,N_1836);
and U2866 (N_2866,N_2229,N_2070);
nor U2867 (N_2867,N_2399,N_2142);
or U2868 (N_2868,N_2017,N_2102);
and U2869 (N_2869,N_2005,N_2389);
nor U2870 (N_2870,N_1847,N_2085);
nand U2871 (N_2871,N_2156,N_2293);
nand U2872 (N_2872,N_2268,N_2274);
nand U2873 (N_2873,N_2076,N_1841);
and U2874 (N_2874,N_2017,N_2394);
nor U2875 (N_2875,N_2200,N_2001);
nand U2876 (N_2876,N_1999,N_2187);
or U2877 (N_2877,N_1992,N_2200);
nor U2878 (N_2878,N_2162,N_2200);
nand U2879 (N_2879,N_1987,N_2345);
and U2880 (N_2880,N_2293,N_1926);
and U2881 (N_2881,N_1811,N_2311);
nor U2882 (N_2882,N_2342,N_1918);
or U2883 (N_2883,N_2114,N_2327);
and U2884 (N_2884,N_2026,N_2286);
or U2885 (N_2885,N_1959,N_2189);
nand U2886 (N_2886,N_1853,N_2309);
or U2887 (N_2887,N_1937,N_2354);
or U2888 (N_2888,N_2367,N_2104);
nor U2889 (N_2889,N_1867,N_1830);
and U2890 (N_2890,N_2168,N_2344);
nor U2891 (N_2891,N_1928,N_2070);
xnor U2892 (N_2892,N_2277,N_2146);
nor U2893 (N_2893,N_2138,N_2122);
nand U2894 (N_2894,N_1894,N_2295);
or U2895 (N_2895,N_2010,N_1944);
nand U2896 (N_2896,N_1982,N_2050);
and U2897 (N_2897,N_2361,N_1977);
or U2898 (N_2898,N_2130,N_2113);
nor U2899 (N_2899,N_2145,N_2110);
nor U2900 (N_2900,N_2357,N_2094);
nor U2901 (N_2901,N_2014,N_2229);
and U2902 (N_2902,N_2025,N_1980);
or U2903 (N_2903,N_2331,N_1877);
nand U2904 (N_2904,N_2298,N_2327);
nand U2905 (N_2905,N_2193,N_2312);
and U2906 (N_2906,N_2276,N_2145);
or U2907 (N_2907,N_1916,N_2105);
nand U2908 (N_2908,N_1997,N_2127);
nand U2909 (N_2909,N_1850,N_2194);
or U2910 (N_2910,N_2193,N_2146);
nor U2911 (N_2911,N_2251,N_2363);
nand U2912 (N_2912,N_2049,N_2023);
nor U2913 (N_2913,N_1954,N_2173);
nor U2914 (N_2914,N_2387,N_2396);
and U2915 (N_2915,N_2038,N_1919);
or U2916 (N_2916,N_2099,N_2195);
and U2917 (N_2917,N_2113,N_2260);
and U2918 (N_2918,N_2105,N_1862);
nor U2919 (N_2919,N_1957,N_1836);
nand U2920 (N_2920,N_2327,N_1852);
nand U2921 (N_2921,N_1958,N_1864);
nand U2922 (N_2922,N_2343,N_1916);
and U2923 (N_2923,N_2068,N_1985);
nand U2924 (N_2924,N_2363,N_2067);
or U2925 (N_2925,N_2055,N_2085);
nor U2926 (N_2926,N_2019,N_2201);
nor U2927 (N_2927,N_1951,N_1955);
and U2928 (N_2928,N_2262,N_2077);
nor U2929 (N_2929,N_2021,N_2070);
or U2930 (N_2930,N_2068,N_2169);
xor U2931 (N_2931,N_2242,N_1980);
nor U2932 (N_2932,N_1812,N_1897);
nand U2933 (N_2933,N_1947,N_1816);
nand U2934 (N_2934,N_2146,N_2074);
or U2935 (N_2935,N_1907,N_1909);
nand U2936 (N_2936,N_2308,N_2349);
or U2937 (N_2937,N_2147,N_1903);
nor U2938 (N_2938,N_1968,N_1849);
nand U2939 (N_2939,N_2118,N_2215);
xnor U2940 (N_2940,N_2177,N_2117);
xor U2941 (N_2941,N_1810,N_2259);
nor U2942 (N_2942,N_1862,N_2026);
and U2943 (N_2943,N_2194,N_2187);
or U2944 (N_2944,N_2270,N_2158);
or U2945 (N_2945,N_2197,N_2148);
or U2946 (N_2946,N_1957,N_2086);
and U2947 (N_2947,N_2385,N_1992);
and U2948 (N_2948,N_2174,N_1910);
and U2949 (N_2949,N_2397,N_2053);
nor U2950 (N_2950,N_2101,N_1824);
nor U2951 (N_2951,N_2345,N_2056);
nand U2952 (N_2952,N_2352,N_1876);
and U2953 (N_2953,N_1978,N_1885);
and U2954 (N_2954,N_2030,N_2210);
or U2955 (N_2955,N_2385,N_2382);
or U2956 (N_2956,N_2006,N_1918);
nor U2957 (N_2957,N_2181,N_2312);
nor U2958 (N_2958,N_1813,N_2160);
nand U2959 (N_2959,N_2193,N_1893);
and U2960 (N_2960,N_2294,N_2090);
nor U2961 (N_2961,N_1921,N_2331);
or U2962 (N_2962,N_2338,N_1904);
nor U2963 (N_2963,N_2267,N_2155);
and U2964 (N_2964,N_2382,N_1887);
nor U2965 (N_2965,N_1864,N_2364);
nand U2966 (N_2966,N_1833,N_2310);
nand U2967 (N_2967,N_2272,N_2112);
or U2968 (N_2968,N_2069,N_2108);
or U2969 (N_2969,N_1872,N_2265);
or U2970 (N_2970,N_2206,N_2345);
nand U2971 (N_2971,N_2357,N_1824);
nor U2972 (N_2972,N_2004,N_2006);
nor U2973 (N_2973,N_2161,N_1891);
and U2974 (N_2974,N_1863,N_2182);
nand U2975 (N_2975,N_2386,N_1862);
nor U2976 (N_2976,N_2148,N_1826);
and U2977 (N_2977,N_2320,N_1828);
or U2978 (N_2978,N_2245,N_1911);
nand U2979 (N_2979,N_1844,N_2272);
nor U2980 (N_2980,N_2103,N_1853);
nor U2981 (N_2981,N_2044,N_2364);
nor U2982 (N_2982,N_2188,N_2040);
nor U2983 (N_2983,N_2350,N_1883);
and U2984 (N_2984,N_2093,N_1938);
nor U2985 (N_2985,N_2189,N_2269);
and U2986 (N_2986,N_2193,N_1876);
and U2987 (N_2987,N_2142,N_2187);
and U2988 (N_2988,N_2148,N_2069);
or U2989 (N_2989,N_2350,N_1818);
and U2990 (N_2990,N_2030,N_1915);
xor U2991 (N_2991,N_2092,N_1873);
nor U2992 (N_2992,N_2274,N_2229);
nor U2993 (N_2993,N_2324,N_2123);
nor U2994 (N_2994,N_1955,N_1814);
and U2995 (N_2995,N_1841,N_2183);
and U2996 (N_2996,N_2163,N_2366);
and U2997 (N_2997,N_2193,N_2080);
or U2998 (N_2998,N_2106,N_2394);
or U2999 (N_2999,N_1935,N_2161);
nor UO_0 (O_0,N_2569,N_2815);
nand UO_1 (O_1,N_2767,N_2929);
and UO_2 (O_2,N_2947,N_2449);
or UO_3 (O_3,N_2763,N_2856);
and UO_4 (O_4,N_2958,N_2519);
and UO_5 (O_5,N_2762,N_2965);
nand UO_6 (O_6,N_2685,N_2599);
xor UO_7 (O_7,N_2456,N_2494);
nand UO_8 (O_8,N_2872,N_2499);
and UO_9 (O_9,N_2547,N_2780);
nor UO_10 (O_10,N_2522,N_2918);
xnor UO_11 (O_11,N_2978,N_2884);
nor UO_12 (O_12,N_2657,N_2843);
or UO_13 (O_13,N_2659,N_2718);
nor UO_14 (O_14,N_2980,N_2896);
nand UO_15 (O_15,N_2855,N_2561);
nand UO_16 (O_16,N_2748,N_2905);
and UO_17 (O_17,N_2906,N_2818);
and UO_18 (O_18,N_2832,N_2939);
or UO_19 (O_19,N_2496,N_2675);
and UO_20 (O_20,N_2487,N_2608);
nand UO_21 (O_21,N_2698,N_2482);
nor UO_22 (O_22,N_2422,N_2808);
and UO_23 (O_23,N_2959,N_2418);
nor UO_24 (O_24,N_2756,N_2806);
and UO_25 (O_25,N_2758,N_2969);
nand UO_26 (O_26,N_2535,N_2864);
xor UO_27 (O_27,N_2736,N_2914);
nand UO_28 (O_28,N_2475,N_2798);
and UO_29 (O_29,N_2874,N_2681);
and UO_30 (O_30,N_2515,N_2513);
and UO_31 (O_31,N_2755,N_2684);
nand UO_32 (O_32,N_2474,N_2461);
and UO_33 (O_33,N_2696,N_2904);
or UO_34 (O_34,N_2576,N_2619);
or UO_35 (O_35,N_2689,N_2664);
and UO_36 (O_36,N_2871,N_2699);
nor UO_37 (O_37,N_2478,N_2924);
and UO_38 (O_38,N_2873,N_2531);
nand UO_39 (O_39,N_2586,N_2973);
and UO_40 (O_40,N_2686,N_2641);
nand UO_41 (O_41,N_2403,N_2652);
nor UO_42 (O_42,N_2636,N_2509);
or UO_43 (O_43,N_2618,N_2423);
nor UO_44 (O_44,N_2783,N_2650);
nor UO_45 (O_45,N_2742,N_2824);
and UO_46 (O_46,N_2940,N_2728);
or UO_47 (O_47,N_2447,N_2703);
nor UO_48 (O_48,N_2869,N_2805);
and UO_49 (O_49,N_2598,N_2429);
nor UO_50 (O_50,N_2867,N_2868);
nor UO_51 (O_51,N_2885,N_2745);
or UO_52 (O_52,N_2846,N_2412);
and UO_53 (O_53,N_2663,N_2433);
nor UO_54 (O_54,N_2789,N_2934);
and UO_55 (O_55,N_2770,N_2775);
nor UO_56 (O_56,N_2903,N_2972);
or UO_57 (O_57,N_2889,N_2936);
or UO_58 (O_58,N_2518,N_2524);
or UO_59 (O_59,N_2857,N_2893);
nand UO_60 (O_60,N_2458,N_2485);
xnor UO_61 (O_61,N_2617,N_2723);
nor UO_62 (O_62,N_2845,N_2428);
xnor UO_63 (O_63,N_2788,N_2411);
or UO_64 (O_64,N_2912,N_2951);
or UO_65 (O_65,N_2639,N_2554);
nand UO_66 (O_66,N_2493,N_2455);
or UO_67 (O_67,N_2649,N_2946);
or UO_68 (O_68,N_2457,N_2585);
nor UO_69 (O_69,N_2628,N_2615);
or UO_70 (O_70,N_2716,N_2717);
and UO_71 (O_71,N_2542,N_2920);
nor UO_72 (O_72,N_2690,N_2627);
nand UO_73 (O_73,N_2975,N_2622);
and UO_74 (O_74,N_2407,N_2771);
nor UO_75 (O_75,N_2715,N_2573);
nand UO_76 (O_76,N_2439,N_2931);
nand UO_77 (O_77,N_2996,N_2550);
and UO_78 (O_78,N_2502,N_2833);
nand UO_79 (O_79,N_2838,N_2928);
or UO_80 (O_80,N_2792,N_2667);
nor UO_81 (O_81,N_2452,N_2655);
nand UO_82 (O_82,N_2441,N_2410);
and UO_83 (O_83,N_2956,N_2437);
or UO_84 (O_84,N_2462,N_2529);
nor UO_85 (O_85,N_2436,N_2416);
xnor UO_86 (O_86,N_2647,N_2656);
nor UO_87 (O_87,N_2725,N_2711);
nor UO_88 (O_88,N_2596,N_2621);
nand UO_89 (O_89,N_2720,N_2802);
nand UO_90 (O_90,N_2473,N_2424);
nand UO_91 (O_91,N_2740,N_2630);
nor UO_92 (O_92,N_2691,N_2701);
nand UO_93 (O_93,N_2580,N_2446);
nor UO_94 (O_94,N_2997,N_2523);
or UO_95 (O_95,N_2801,N_2404);
nand UO_96 (O_96,N_2564,N_2993);
nor UO_97 (O_97,N_2707,N_2814);
nand UO_98 (O_98,N_2694,N_2671);
or UO_99 (O_99,N_2527,N_2810);
and UO_100 (O_100,N_2556,N_2614);
nor UO_101 (O_101,N_2638,N_2536);
or UO_102 (O_102,N_2520,N_2776);
and UO_103 (O_103,N_2442,N_2507);
and UO_104 (O_104,N_2425,N_2505);
nor UO_105 (O_105,N_2852,N_2710);
xnor UO_106 (O_106,N_2549,N_2408);
nor UO_107 (O_107,N_2766,N_2480);
xnor UO_108 (O_108,N_2453,N_2730);
and UO_109 (O_109,N_2787,N_2534);
or UO_110 (O_110,N_2445,N_2620);
and UO_111 (O_111,N_2508,N_2779);
or UO_112 (O_112,N_2797,N_2574);
nand UO_113 (O_113,N_2785,N_2584);
xor UO_114 (O_114,N_2477,N_2902);
or UO_115 (O_115,N_2925,N_2577);
or UO_116 (O_116,N_2813,N_2409);
or UO_117 (O_117,N_2858,N_2970);
nor UO_118 (O_118,N_2495,N_2849);
nor UO_119 (O_119,N_2877,N_2603);
nor UO_120 (O_120,N_2963,N_2895);
and UO_121 (O_121,N_2721,N_2605);
nand UO_122 (O_122,N_2420,N_2938);
nor UO_123 (O_123,N_2821,N_2601);
nor UO_124 (O_124,N_2415,N_2668);
nand UO_125 (O_125,N_2962,N_2942);
and UO_126 (O_126,N_2516,N_2413);
and UO_127 (O_127,N_2419,N_2488);
and UO_128 (O_128,N_2559,N_2572);
nor UO_129 (O_129,N_2953,N_2643);
nand UO_130 (O_130,N_2977,N_2911);
or UO_131 (O_131,N_2909,N_2807);
and UO_132 (O_132,N_2537,N_2796);
nor UO_133 (O_133,N_2486,N_2582);
or UO_134 (O_134,N_2553,N_2506);
nor UO_135 (O_135,N_2662,N_2862);
nand UO_136 (O_136,N_2503,N_2632);
nor UO_137 (O_137,N_2994,N_2886);
nor UO_138 (O_138,N_2460,N_2713);
and UO_139 (O_139,N_2570,N_2820);
nand UO_140 (O_140,N_2781,N_2427);
or UO_141 (O_141,N_2830,N_2991);
nand UO_142 (O_142,N_2670,N_2840);
nand UO_143 (O_143,N_2567,N_2592);
nand UO_144 (O_144,N_2539,N_2876);
or UO_145 (O_145,N_2658,N_2944);
nor UO_146 (O_146,N_2459,N_2538);
or UO_147 (O_147,N_2687,N_2930);
and UO_148 (O_148,N_2481,N_2450);
nand UO_149 (O_149,N_2490,N_2901);
xnor UO_150 (O_150,N_2489,N_2752);
and UO_151 (O_151,N_2741,N_2764);
or UO_152 (O_152,N_2544,N_2759);
nand UO_153 (O_153,N_2784,N_2676);
nor UO_154 (O_154,N_2406,N_2402);
nand UO_155 (O_155,N_2882,N_2917);
and UO_156 (O_156,N_2653,N_2602);
and UO_157 (O_157,N_2878,N_2467);
and UO_158 (O_158,N_2811,N_2954);
nor UO_159 (O_159,N_2823,N_2837);
and UO_160 (O_160,N_2774,N_2753);
xor UO_161 (O_161,N_2842,N_2525);
and UO_162 (O_162,N_2955,N_2727);
nor UO_163 (O_163,N_2919,N_2982);
nor UO_164 (O_164,N_2440,N_2678);
and UO_165 (O_165,N_2979,N_2498);
nand UO_166 (O_166,N_2511,N_2479);
nor UO_167 (O_167,N_2483,N_2562);
and UO_168 (O_168,N_2735,N_2985);
nor UO_169 (O_169,N_2695,N_2999);
and UO_170 (O_170,N_2990,N_2624);
xor UO_171 (O_171,N_2637,N_2540);
nor UO_172 (O_172,N_2665,N_2826);
nand UO_173 (O_173,N_2616,N_2644);
nor UO_174 (O_174,N_2921,N_2633);
and UO_175 (O_175,N_2579,N_2654);
nor UO_176 (O_176,N_2754,N_2992);
and UO_177 (O_177,N_2899,N_2916);
nor UO_178 (O_178,N_2952,N_2432);
and UO_179 (O_179,N_2998,N_2631);
nor UO_180 (O_180,N_2848,N_2541);
nor UO_181 (O_181,N_2532,N_2565);
xnor UO_182 (O_182,N_2853,N_2769);
nand UO_183 (O_183,N_2609,N_2746);
nand UO_184 (O_184,N_2545,N_2768);
nand UO_185 (O_185,N_2629,N_2733);
nor UO_186 (O_186,N_2590,N_2860);
or UO_187 (O_187,N_2575,N_2471);
nor UO_188 (O_188,N_2828,N_2894);
nand UO_189 (O_189,N_2708,N_2737);
nand UO_190 (O_190,N_2926,N_2504);
nand UO_191 (O_191,N_2847,N_2812);
nand UO_192 (O_192,N_2533,N_2816);
or UO_193 (O_193,N_2825,N_2760);
nand UO_194 (O_194,N_2484,N_2907);
nand UO_195 (O_195,N_2677,N_2822);
nand UO_196 (O_196,N_2880,N_2438);
or UO_197 (O_197,N_2898,N_2551);
or UO_198 (O_198,N_2600,N_2986);
and UO_199 (O_199,N_2604,N_2400);
and UO_200 (O_200,N_2887,N_2623);
nor UO_201 (O_201,N_2995,N_2714);
nor UO_202 (O_202,N_2957,N_2836);
or UO_203 (O_203,N_2588,N_2786);
nor UO_204 (O_204,N_2530,N_2568);
xor UO_205 (O_205,N_2426,N_2851);
xor UO_206 (O_206,N_2597,N_2431);
nand UO_207 (O_207,N_2750,N_2712);
or UO_208 (O_208,N_2875,N_2772);
or UO_209 (O_209,N_2405,N_2448);
or UO_210 (O_210,N_2839,N_2964);
and UO_211 (O_211,N_2790,N_2470);
nand UO_212 (O_212,N_2866,N_2491);
or UO_213 (O_213,N_2922,N_2645);
or UO_214 (O_214,N_2543,N_2831);
nand UO_215 (O_215,N_2835,N_2510);
and UO_216 (O_216,N_2945,N_2444);
xor UO_217 (O_217,N_2799,N_2625);
nand UO_218 (O_218,N_2626,N_2611);
and UO_219 (O_219,N_2443,N_2651);
nand UO_220 (O_220,N_2581,N_2883);
nor UO_221 (O_221,N_2988,N_2827);
nor UO_222 (O_222,N_2546,N_2900);
nand UO_223 (O_223,N_2782,N_2937);
or UO_224 (O_224,N_2517,N_2960);
or UO_225 (O_225,N_2943,N_2700);
and UO_226 (O_226,N_2476,N_2791);
or UO_227 (O_227,N_2526,N_2558);
and UO_228 (O_228,N_2989,N_2417);
or UO_229 (O_229,N_2738,N_2680);
and UO_230 (O_230,N_2469,N_2591);
nor UO_231 (O_231,N_2892,N_2688);
or UO_232 (O_232,N_2834,N_2679);
nand UO_233 (O_233,N_2646,N_2451);
and UO_234 (O_234,N_2879,N_2589);
nor UO_235 (O_235,N_2583,N_2729);
nand UO_236 (O_236,N_2751,N_2935);
and UO_237 (O_237,N_2706,N_2660);
nor UO_238 (O_238,N_2744,N_2672);
and UO_239 (O_239,N_2793,N_2897);
nor UO_240 (O_240,N_2640,N_2606);
or UO_241 (O_241,N_2910,N_2863);
nor UO_242 (O_242,N_2557,N_2794);
nor UO_243 (O_243,N_2560,N_2739);
xnor UO_244 (O_244,N_2642,N_2414);
or UO_245 (O_245,N_2634,N_2757);
and UO_246 (O_246,N_2865,N_2430);
and UO_247 (O_247,N_2734,N_2492);
and UO_248 (O_248,N_2859,N_2466);
and UO_249 (O_249,N_2724,N_2674);
or UO_250 (O_250,N_2552,N_2464);
nor UO_251 (O_251,N_2731,N_2778);
and UO_252 (O_252,N_2747,N_2610);
nand UO_253 (O_253,N_2468,N_2932);
and UO_254 (O_254,N_2941,N_2661);
and UO_255 (O_255,N_2817,N_2593);
nand UO_256 (O_256,N_2881,N_2613);
nand UO_257 (O_257,N_2773,N_2434);
or UO_258 (O_258,N_2669,N_2974);
or UO_259 (O_259,N_2761,N_2749);
and UO_260 (O_260,N_2578,N_2804);
or UO_261 (O_261,N_2841,N_2971);
and UO_262 (O_262,N_2548,N_2803);
and UO_263 (O_263,N_2709,N_2987);
or UO_264 (O_264,N_2981,N_2497);
nor UO_265 (O_265,N_2850,N_2765);
nand UO_266 (O_266,N_2521,N_2563);
and UO_267 (O_267,N_2692,N_2948);
nor UO_268 (O_268,N_2501,N_2950);
nand UO_269 (O_269,N_2528,N_2933);
and UO_270 (O_270,N_2976,N_2743);
or UO_271 (O_271,N_2683,N_2719);
nor UO_272 (O_272,N_2514,N_2949);
nor UO_273 (O_273,N_2587,N_2682);
nor UO_274 (O_274,N_2612,N_2809);
and UO_275 (O_275,N_2421,N_2891);
nor UO_276 (O_276,N_2777,N_2705);
nor UO_277 (O_277,N_2435,N_2913);
and UO_278 (O_278,N_2961,N_2870);
xor UO_279 (O_279,N_2915,N_2927);
xor UO_280 (O_280,N_2967,N_2968);
nand UO_281 (O_281,N_2854,N_2454);
nor UO_282 (O_282,N_2722,N_2829);
nand UO_283 (O_283,N_2861,N_2607);
nand UO_284 (O_284,N_2702,N_2555);
xnor UO_285 (O_285,N_2693,N_2648);
nor UO_286 (O_286,N_2890,N_2732);
and UO_287 (O_287,N_2726,N_2704);
nor UO_288 (O_288,N_2984,N_2844);
and UO_289 (O_289,N_2666,N_2635);
nand UO_290 (O_290,N_2465,N_2463);
or UO_291 (O_291,N_2673,N_2983);
nand UO_292 (O_292,N_2819,N_2888);
nor UO_293 (O_293,N_2966,N_2923);
nand UO_294 (O_294,N_2512,N_2595);
or UO_295 (O_295,N_2571,N_2401);
and UO_296 (O_296,N_2908,N_2697);
or UO_297 (O_297,N_2795,N_2472);
or UO_298 (O_298,N_2800,N_2594);
or UO_299 (O_299,N_2566,N_2500);
or UO_300 (O_300,N_2902,N_2495);
nor UO_301 (O_301,N_2930,N_2411);
nor UO_302 (O_302,N_2815,N_2760);
nand UO_303 (O_303,N_2620,N_2741);
and UO_304 (O_304,N_2466,N_2575);
and UO_305 (O_305,N_2487,N_2565);
nand UO_306 (O_306,N_2818,N_2771);
nor UO_307 (O_307,N_2660,N_2915);
or UO_308 (O_308,N_2539,N_2486);
nor UO_309 (O_309,N_2583,N_2944);
nor UO_310 (O_310,N_2688,N_2961);
and UO_311 (O_311,N_2814,N_2691);
or UO_312 (O_312,N_2817,N_2711);
nor UO_313 (O_313,N_2403,N_2491);
and UO_314 (O_314,N_2604,N_2421);
and UO_315 (O_315,N_2465,N_2462);
nor UO_316 (O_316,N_2689,N_2866);
or UO_317 (O_317,N_2707,N_2423);
or UO_318 (O_318,N_2459,N_2641);
and UO_319 (O_319,N_2915,N_2649);
nand UO_320 (O_320,N_2585,N_2604);
nor UO_321 (O_321,N_2932,N_2896);
nor UO_322 (O_322,N_2887,N_2500);
nor UO_323 (O_323,N_2822,N_2801);
or UO_324 (O_324,N_2483,N_2724);
or UO_325 (O_325,N_2767,N_2689);
and UO_326 (O_326,N_2977,N_2618);
nor UO_327 (O_327,N_2811,N_2494);
or UO_328 (O_328,N_2613,N_2434);
and UO_329 (O_329,N_2425,N_2656);
nor UO_330 (O_330,N_2866,N_2739);
nand UO_331 (O_331,N_2489,N_2578);
nor UO_332 (O_332,N_2764,N_2894);
and UO_333 (O_333,N_2650,N_2403);
and UO_334 (O_334,N_2430,N_2974);
nor UO_335 (O_335,N_2797,N_2774);
and UO_336 (O_336,N_2926,N_2691);
nor UO_337 (O_337,N_2429,N_2905);
or UO_338 (O_338,N_2683,N_2942);
or UO_339 (O_339,N_2533,N_2997);
or UO_340 (O_340,N_2811,N_2782);
nor UO_341 (O_341,N_2727,N_2488);
or UO_342 (O_342,N_2907,N_2464);
and UO_343 (O_343,N_2762,N_2771);
nand UO_344 (O_344,N_2851,N_2790);
nor UO_345 (O_345,N_2791,N_2917);
or UO_346 (O_346,N_2863,N_2447);
nand UO_347 (O_347,N_2420,N_2648);
nand UO_348 (O_348,N_2584,N_2867);
and UO_349 (O_349,N_2411,N_2952);
nand UO_350 (O_350,N_2897,N_2635);
nand UO_351 (O_351,N_2502,N_2991);
nor UO_352 (O_352,N_2424,N_2548);
and UO_353 (O_353,N_2496,N_2943);
or UO_354 (O_354,N_2408,N_2708);
or UO_355 (O_355,N_2528,N_2594);
or UO_356 (O_356,N_2851,N_2475);
and UO_357 (O_357,N_2511,N_2758);
nor UO_358 (O_358,N_2592,N_2402);
and UO_359 (O_359,N_2651,N_2510);
nand UO_360 (O_360,N_2983,N_2574);
and UO_361 (O_361,N_2766,N_2506);
nand UO_362 (O_362,N_2439,N_2549);
nand UO_363 (O_363,N_2698,N_2609);
or UO_364 (O_364,N_2559,N_2945);
or UO_365 (O_365,N_2777,N_2656);
nand UO_366 (O_366,N_2947,N_2602);
nor UO_367 (O_367,N_2450,N_2932);
nand UO_368 (O_368,N_2624,N_2681);
and UO_369 (O_369,N_2902,N_2879);
or UO_370 (O_370,N_2420,N_2858);
or UO_371 (O_371,N_2439,N_2571);
or UO_372 (O_372,N_2849,N_2863);
xnor UO_373 (O_373,N_2649,N_2569);
nand UO_374 (O_374,N_2860,N_2549);
and UO_375 (O_375,N_2576,N_2671);
and UO_376 (O_376,N_2800,N_2807);
nand UO_377 (O_377,N_2677,N_2831);
nand UO_378 (O_378,N_2502,N_2895);
or UO_379 (O_379,N_2545,N_2405);
and UO_380 (O_380,N_2694,N_2960);
and UO_381 (O_381,N_2753,N_2491);
or UO_382 (O_382,N_2884,N_2880);
nor UO_383 (O_383,N_2975,N_2757);
and UO_384 (O_384,N_2641,N_2571);
nor UO_385 (O_385,N_2891,N_2972);
and UO_386 (O_386,N_2493,N_2676);
or UO_387 (O_387,N_2482,N_2780);
nor UO_388 (O_388,N_2673,N_2755);
nor UO_389 (O_389,N_2803,N_2859);
nor UO_390 (O_390,N_2857,N_2952);
nand UO_391 (O_391,N_2805,N_2904);
nor UO_392 (O_392,N_2945,N_2531);
nand UO_393 (O_393,N_2674,N_2956);
and UO_394 (O_394,N_2744,N_2504);
nor UO_395 (O_395,N_2866,N_2919);
nand UO_396 (O_396,N_2907,N_2565);
nand UO_397 (O_397,N_2470,N_2742);
and UO_398 (O_398,N_2835,N_2971);
nor UO_399 (O_399,N_2786,N_2925);
or UO_400 (O_400,N_2469,N_2965);
or UO_401 (O_401,N_2971,N_2960);
nor UO_402 (O_402,N_2679,N_2860);
nor UO_403 (O_403,N_2622,N_2741);
nor UO_404 (O_404,N_2644,N_2636);
and UO_405 (O_405,N_2981,N_2587);
nor UO_406 (O_406,N_2730,N_2867);
nand UO_407 (O_407,N_2711,N_2931);
nor UO_408 (O_408,N_2923,N_2969);
xor UO_409 (O_409,N_2810,N_2416);
nand UO_410 (O_410,N_2735,N_2484);
and UO_411 (O_411,N_2954,N_2869);
nand UO_412 (O_412,N_2443,N_2926);
and UO_413 (O_413,N_2630,N_2821);
and UO_414 (O_414,N_2468,N_2567);
or UO_415 (O_415,N_2983,N_2840);
nand UO_416 (O_416,N_2554,N_2746);
nand UO_417 (O_417,N_2625,N_2986);
and UO_418 (O_418,N_2701,N_2855);
or UO_419 (O_419,N_2835,N_2748);
or UO_420 (O_420,N_2749,N_2909);
or UO_421 (O_421,N_2737,N_2540);
nor UO_422 (O_422,N_2501,N_2640);
nor UO_423 (O_423,N_2633,N_2594);
or UO_424 (O_424,N_2662,N_2725);
or UO_425 (O_425,N_2550,N_2854);
nor UO_426 (O_426,N_2513,N_2835);
nand UO_427 (O_427,N_2963,N_2746);
or UO_428 (O_428,N_2960,N_2769);
or UO_429 (O_429,N_2599,N_2908);
and UO_430 (O_430,N_2478,N_2407);
or UO_431 (O_431,N_2741,N_2965);
or UO_432 (O_432,N_2962,N_2518);
and UO_433 (O_433,N_2442,N_2409);
or UO_434 (O_434,N_2997,N_2476);
nor UO_435 (O_435,N_2729,N_2815);
nor UO_436 (O_436,N_2409,N_2479);
and UO_437 (O_437,N_2440,N_2495);
nor UO_438 (O_438,N_2669,N_2755);
or UO_439 (O_439,N_2622,N_2660);
and UO_440 (O_440,N_2729,N_2580);
nor UO_441 (O_441,N_2660,N_2537);
or UO_442 (O_442,N_2914,N_2681);
nor UO_443 (O_443,N_2658,N_2759);
nor UO_444 (O_444,N_2568,N_2793);
or UO_445 (O_445,N_2738,N_2976);
or UO_446 (O_446,N_2535,N_2651);
or UO_447 (O_447,N_2577,N_2656);
nand UO_448 (O_448,N_2805,N_2930);
nor UO_449 (O_449,N_2573,N_2901);
or UO_450 (O_450,N_2603,N_2659);
nand UO_451 (O_451,N_2836,N_2469);
and UO_452 (O_452,N_2432,N_2997);
or UO_453 (O_453,N_2466,N_2443);
nand UO_454 (O_454,N_2961,N_2757);
and UO_455 (O_455,N_2869,N_2465);
or UO_456 (O_456,N_2898,N_2778);
and UO_457 (O_457,N_2898,N_2832);
nand UO_458 (O_458,N_2494,N_2800);
or UO_459 (O_459,N_2488,N_2898);
or UO_460 (O_460,N_2570,N_2866);
or UO_461 (O_461,N_2571,N_2409);
nand UO_462 (O_462,N_2651,N_2850);
nand UO_463 (O_463,N_2401,N_2853);
and UO_464 (O_464,N_2957,N_2905);
and UO_465 (O_465,N_2879,N_2839);
nor UO_466 (O_466,N_2473,N_2727);
nor UO_467 (O_467,N_2635,N_2402);
nand UO_468 (O_468,N_2918,N_2587);
and UO_469 (O_469,N_2865,N_2650);
and UO_470 (O_470,N_2759,N_2604);
or UO_471 (O_471,N_2637,N_2542);
nand UO_472 (O_472,N_2707,N_2935);
or UO_473 (O_473,N_2741,N_2841);
nor UO_474 (O_474,N_2914,N_2832);
or UO_475 (O_475,N_2657,N_2584);
or UO_476 (O_476,N_2771,N_2465);
nor UO_477 (O_477,N_2506,N_2634);
or UO_478 (O_478,N_2610,N_2487);
xor UO_479 (O_479,N_2821,N_2459);
nor UO_480 (O_480,N_2538,N_2469);
nor UO_481 (O_481,N_2921,N_2728);
nor UO_482 (O_482,N_2850,N_2862);
nand UO_483 (O_483,N_2671,N_2667);
and UO_484 (O_484,N_2753,N_2428);
or UO_485 (O_485,N_2453,N_2459);
nand UO_486 (O_486,N_2796,N_2917);
and UO_487 (O_487,N_2599,N_2985);
and UO_488 (O_488,N_2949,N_2495);
or UO_489 (O_489,N_2942,N_2725);
and UO_490 (O_490,N_2831,N_2403);
nand UO_491 (O_491,N_2611,N_2844);
or UO_492 (O_492,N_2700,N_2730);
nand UO_493 (O_493,N_2576,N_2914);
or UO_494 (O_494,N_2608,N_2686);
or UO_495 (O_495,N_2669,N_2525);
or UO_496 (O_496,N_2743,N_2877);
xor UO_497 (O_497,N_2837,N_2404);
or UO_498 (O_498,N_2608,N_2654);
and UO_499 (O_499,N_2479,N_2734);
endmodule