module basic_1000_10000_1500_10_levels_1xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_384,In_260);
nor U1 (N_1,In_801,In_388);
nand U2 (N_2,In_910,In_280);
or U3 (N_3,In_201,In_277);
or U4 (N_4,In_752,In_637);
nand U5 (N_5,In_71,In_11);
nand U6 (N_6,In_721,In_414);
nor U7 (N_7,In_290,In_575);
nand U8 (N_8,In_559,In_116);
nor U9 (N_9,In_767,In_429);
or U10 (N_10,In_421,In_86);
nand U11 (N_11,In_122,In_0);
nand U12 (N_12,In_883,In_884);
and U13 (N_13,In_687,In_8);
or U14 (N_14,In_156,In_203);
or U15 (N_15,In_436,In_236);
nand U16 (N_16,In_383,In_413);
and U17 (N_17,In_769,In_862);
and U18 (N_18,In_645,In_165);
or U19 (N_19,In_919,In_706);
or U20 (N_20,In_323,In_219);
nand U21 (N_21,In_90,In_668);
nor U22 (N_22,In_195,In_850);
or U23 (N_23,In_274,In_547);
nand U24 (N_24,In_690,In_155);
and U25 (N_25,In_560,In_617);
nor U26 (N_26,In_716,In_266);
and U27 (N_27,In_856,In_631);
nand U28 (N_28,In_820,In_902);
and U29 (N_29,In_55,In_492);
and U30 (N_30,In_322,In_239);
and U31 (N_31,In_109,In_700);
and U32 (N_32,In_192,In_47);
or U33 (N_33,In_785,In_808);
and U34 (N_34,In_650,In_120);
and U35 (N_35,In_937,In_526);
and U36 (N_36,In_346,In_168);
nor U37 (N_37,In_466,In_273);
or U38 (N_38,In_38,In_476);
or U39 (N_39,In_275,In_283);
nand U40 (N_40,In_362,In_350);
or U41 (N_41,In_479,In_848);
and U42 (N_42,In_488,In_873);
and U43 (N_43,In_939,In_517);
nor U44 (N_44,In_791,In_503);
or U45 (N_45,In_976,In_999);
or U46 (N_46,In_54,In_170);
nor U47 (N_47,In_368,In_740);
nor U48 (N_48,In_226,In_583);
nor U49 (N_49,In_562,In_530);
or U50 (N_50,In_258,In_572);
or U51 (N_51,In_935,In_371);
and U52 (N_52,In_899,In_656);
nor U53 (N_53,In_410,In_215);
or U54 (N_54,In_35,In_874);
and U55 (N_55,In_320,In_345);
nor U56 (N_56,In_119,In_582);
xor U57 (N_57,In_265,In_741);
or U58 (N_58,In_669,In_243);
nor U59 (N_59,In_259,In_132);
nand U60 (N_60,In_3,In_980);
and U61 (N_61,In_692,In_540);
nor U62 (N_62,In_27,In_916);
nor U63 (N_63,In_93,In_361);
or U64 (N_64,In_764,In_748);
nand U65 (N_65,In_638,In_357);
nand U66 (N_66,In_568,In_872);
nand U67 (N_67,In_269,In_197);
or U68 (N_68,In_127,In_111);
or U69 (N_69,In_250,In_257);
nand U70 (N_70,In_888,In_296);
and U71 (N_71,In_146,In_763);
nor U72 (N_72,In_861,In_711);
or U73 (N_73,In_534,In_446);
and U74 (N_74,In_955,In_773);
nand U75 (N_75,In_846,In_697);
or U76 (N_76,In_64,In_954);
or U77 (N_77,In_944,In_768);
or U78 (N_78,In_580,In_489);
and U79 (N_79,In_89,In_126);
and U80 (N_80,In_92,In_536);
nand U81 (N_81,In_851,In_104);
nor U82 (N_82,In_579,In_524);
nor U83 (N_83,In_181,In_807);
nor U84 (N_84,In_314,In_306);
or U85 (N_85,In_609,In_604);
nand U86 (N_86,In_249,In_211);
or U87 (N_87,In_214,In_924);
or U88 (N_88,In_65,In_940);
nor U89 (N_89,In_693,In_304);
or U90 (N_90,In_894,In_490);
and U91 (N_91,In_777,In_480);
or U92 (N_92,In_68,In_847);
nor U93 (N_93,In_589,In_233);
and U94 (N_94,In_738,In_449);
xor U95 (N_95,In_658,In_73);
nor U96 (N_96,In_319,In_284);
nand U97 (N_97,In_806,In_974);
nor U98 (N_98,In_367,In_43);
and U99 (N_99,In_929,In_992);
or U100 (N_100,In_177,In_707);
and U101 (N_101,In_473,In_882);
or U102 (N_102,In_406,In_625);
nor U103 (N_103,In_20,In_61);
and U104 (N_104,In_267,In_810);
nand U105 (N_105,In_673,In_31);
and U106 (N_106,In_981,In_917);
nor U107 (N_107,In_797,In_729);
nand U108 (N_108,In_210,In_506);
or U109 (N_109,In_813,In_46);
or U110 (N_110,In_292,In_230);
and U111 (N_111,In_825,In_863);
nand U112 (N_112,In_375,In_634);
or U113 (N_113,In_427,In_727);
nand U114 (N_114,In_671,In_996);
nand U115 (N_115,In_816,In_455);
nor U116 (N_116,In_196,In_166);
or U117 (N_117,In_291,In_610);
or U118 (N_118,In_930,In_107);
nor U119 (N_119,In_705,In_951);
nor U120 (N_120,In_245,In_461);
nor U121 (N_121,In_184,In_835);
or U122 (N_122,In_643,In_431);
or U123 (N_123,In_584,In_32);
nor U124 (N_124,In_702,In_761);
nand U125 (N_125,In_433,In_42);
nand U126 (N_126,In_853,In_983);
nand U127 (N_127,In_869,In_244);
or U128 (N_128,In_667,In_486);
nand U129 (N_129,In_97,In_636);
and U130 (N_130,In_554,In_264);
nor U131 (N_131,In_337,In_722);
nand U132 (N_132,In_333,In_933);
nor U133 (N_133,In_527,In_922);
and U134 (N_134,In_72,In_784);
and U135 (N_135,In_788,In_703);
or U136 (N_136,In_299,In_733);
nand U137 (N_137,In_392,In_571);
nand U138 (N_138,In_194,In_84);
nand U139 (N_139,In_234,In_499);
nor U140 (N_140,In_6,In_751);
nor U141 (N_141,In_154,In_881);
nor U142 (N_142,In_439,In_659);
nand U143 (N_143,In_648,In_467);
nor U144 (N_144,In_532,In_300);
nor U145 (N_145,In_158,In_223);
nor U146 (N_146,In_485,In_553);
and U147 (N_147,In_642,In_927);
and U148 (N_148,In_897,In_246);
nor U149 (N_149,In_889,In_238);
nand U150 (N_150,In_686,In_440);
nor U151 (N_151,In_521,In_312);
nand U152 (N_152,In_630,In_150);
nand U153 (N_153,In_516,In_484);
and U154 (N_154,In_224,In_815);
nand U155 (N_155,In_188,In_338);
and U156 (N_156,In_321,In_16);
nor U157 (N_157,In_369,In_366);
nor U158 (N_158,In_546,In_41);
or U159 (N_159,In_443,In_652);
and U160 (N_160,In_313,In_528);
or U161 (N_161,In_354,In_399);
nor U162 (N_162,In_207,In_344);
or U163 (N_163,In_900,In_103);
nor U164 (N_164,In_453,In_618);
nand U165 (N_165,In_744,In_670);
or U166 (N_166,In_153,In_593);
nor U167 (N_167,In_858,In_408);
nand U168 (N_168,In_931,In_654);
nand U169 (N_169,In_469,In_404);
nor U170 (N_170,In_533,In_549);
and U171 (N_171,In_890,In_135);
or U172 (N_172,In_370,In_376);
nor U173 (N_173,In_978,In_920);
nand U174 (N_174,In_989,In_566);
or U175 (N_175,In_938,In_918);
nor U176 (N_176,In_735,In_494);
nand U177 (N_177,In_666,In_649);
or U178 (N_178,In_160,In_787);
nand U179 (N_179,In_49,In_493);
nor U180 (N_180,In_576,In_870);
nor U181 (N_181,In_696,In_339);
nor U182 (N_182,In_915,In_843);
and U183 (N_183,In_110,In_204);
or U184 (N_184,In_961,In_471);
or U185 (N_185,In_515,In_48);
and U186 (N_186,In_134,In_783);
and U187 (N_187,In_601,In_475);
nand U188 (N_188,In_830,In_694);
nor U189 (N_189,In_302,In_867);
nor U190 (N_190,In_661,In_298);
and U191 (N_191,In_941,In_24);
nand U192 (N_192,In_749,In_10);
nand U193 (N_193,In_923,In_864);
nor U194 (N_194,In_614,In_993);
and U195 (N_195,In_37,In_912);
nor U196 (N_196,In_823,In_837);
nand U197 (N_197,In_836,In_229);
and U198 (N_198,In_794,In_613);
nor U199 (N_199,In_833,In_151);
nand U200 (N_200,In_611,In_141);
nand U201 (N_201,In_555,In_470);
or U202 (N_202,In_828,In_420);
or U203 (N_203,In_627,In_63);
nor U204 (N_204,In_557,In_422);
nor U205 (N_205,In_180,In_714);
nand U206 (N_206,In_198,In_85);
nor U207 (N_207,In_364,In_419);
nor U208 (N_208,In_795,In_818);
nor U209 (N_209,In_832,In_50);
and U210 (N_210,In_495,In_193);
nand U211 (N_211,In_755,In_209);
and U212 (N_212,In_444,In_7);
nand U213 (N_213,In_909,In_651);
or U214 (N_214,In_569,In_595);
nand U215 (N_215,In_336,In_653);
nor U216 (N_216,In_70,In_950);
nor U217 (N_217,In_854,In_23);
or U218 (N_218,In_871,In_289);
nor U219 (N_219,In_682,In_152);
or U220 (N_220,In_616,In_74);
nor U221 (N_221,In_771,In_908);
nor U222 (N_222,In_56,In_766);
nor U223 (N_223,In_720,In_966);
or U224 (N_224,In_936,In_543);
nand U225 (N_225,In_412,In_615);
or U226 (N_226,In_268,In_728);
or U227 (N_227,In_977,In_281);
xnor U228 (N_228,In_905,In_819);
nor U229 (N_229,In_628,In_647);
nor U230 (N_230,In_734,In_606);
nand U231 (N_231,In_123,In_866);
and U232 (N_232,In_124,In_789);
or U233 (N_233,In_351,In_772);
nand U234 (N_234,In_497,In_82);
nor U235 (N_235,In_952,In_732);
nor U236 (N_236,In_885,In_523);
nand U237 (N_237,In_301,In_365);
nor U238 (N_238,In_891,In_26);
or U239 (N_239,In_505,In_959);
nand U240 (N_240,In_762,In_953);
nand U241 (N_241,In_641,In_674);
and U242 (N_242,In_149,In_254);
or U243 (N_243,In_676,In_498);
or U244 (N_244,In_44,In_307);
or U245 (N_245,In_739,In_675);
and U246 (N_246,In_548,In_665);
and U247 (N_247,In_970,In_102);
and U248 (N_248,In_826,In_445);
nand U249 (N_249,In_802,In_112);
nor U250 (N_250,In_708,In_347);
nor U251 (N_251,In_679,In_33);
and U252 (N_252,In_372,In_512);
nand U253 (N_253,In_220,In_875);
nand U254 (N_254,In_695,In_960);
or U255 (N_255,In_827,In_242);
and U256 (N_256,In_991,In_531);
or U257 (N_257,In_844,In_387);
nor U258 (N_258,In_632,In_441);
nand U259 (N_259,In_926,In_901);
or U260 (N_260,In_459,In_963);
and U261 (N_261,In_293,In_876);
or U262 (N_262,In_639,In_608);
nand U263 (N_263,In_539,In_987);
nor U264 (N_264,In_564,In_684);
and U265 (N_265,In_191,In_162);
and U266 (N_266,In_971,In_263);
nor U267 (N_267,In_348,In_213);
nor U268 (N_268,In_796,In_225);
and U269 (N_269,In_698,In_96);
nor U270 (N_270,In_754,In_432);
and U271 (N_271,In_522,In_745);
and U272 (N_272,In_736,In_57);
nand U273 (N_273,In_776,In_898);
and U274 (N_274,In_261,In_840);
nand U275 (N_275,In_635,In_221);
or U276 (N_276,In_457,In_311);
nor U277 (N_277,In_903,In_774);
and U278 (N_278,In_664,In_680);
nor U279 (N_279,In_94,In_19);
nor U280 (N_280,In_409,In_760);
and U281 (N_281,In_949,In_359);
and U282 (N_282,In_779,In_279);
nor U283 (N_283,In_317,In_398);
nor U284 (N_284,In_513,In_332);
nor U285 (N_285,In_814,In_222);
nor U286 (N_286,In_792,In_435);
nand U287 (N_287,In_585,In_100);
nand U288 (N_288,In_757,In_353);
and U289 (N_289,In_525,In_688);
and U290 (N_290,In_809,In_545);
nor U291 (N_291,In_147,In_510);
nand U292 (N_292,In_770,In_538);
nor U293 (N_293,In_561,In_756);
nand U294 (N_294,In_30,In_262);
or U295 (N_295,In_40,In_437);
or U296 (N_296,In_660,In_859);
nor U297 (N_297,In_15,In_159);
and U298 (N_298,In_701,In_948);
or U299 (N_299,In_21,In_790);
nand U300 (N_300,In_212,In_906);
nand U301 (N_301,In_128,In_13);
nor U302 (N_302,In_169,In_137);
nor U303 (N_303,In_381,In_343);
nand U304 (N_304,In_947,In_130);
or U305 (N_305,In_450,In_276);
nor U306 (N_306,In_986,In_172);
nor U307 (N_307,In_681,In_984);
nand U308 (N_308,In_723,In_330);
and U309 (N_309,In_550,In_623);
and U310 (N_310,In_382,In_468);
or U311 (N_311,In_893,In_185);
nor U312 (N_312,In_29,In_588);
nand U313 (N_313,In_379,In_25);
nand U314 (N_314,In_592,In_759);
and U315 (N_315,In_227,In_535);
nand U316 (N_316,In_442,In_454);
or U317 (N_317,In_886,In_341);
nor U318 (N_318,In_318,In_988);
or U319 (N_319,In_157,In_709);
nand U320 (N_320,In_465,In_904);
nor U321 (N_321,In_45,In_725);
nor U322 (N_322,In_821,In_925);
or U323 (N_323,In_596,In_448);
or U324 (N_324,In_712,In_360);
nand U325 (N_325,In_424,In_115);
nand U326 (N_326,In_782,In_464);
nand U327 (N_327,In_145,In_934);
nand U328 (N_328,In_327,In_985);
or U329 (N_329,In_887,In_75);
nor U330 (N_330,In_303,In_182);
and U331 (N_331,In_140,In_133);
xnor U332 (N_332,In_393,In_143);
nor U333 (N_333,In_52,In_282);
nor U334 (N_334,In_385,In_504);
or U335 (N_335,In_186,In_77);
or U336 (N_336,In_726,In_39);
nand U337 (N_337,In_541,In_101);
nor U338 (N_338,In_520,In_200);
nand U339 (N_339,In_217,In_288);
and U340 (N_340,In_403,In_781);
and U341 (N_341,In_252,In_811);
and U342 (N_342,In_451,In_612);
nor U343 (N_343,In_841,In_619);
or U344 (N_344,In_114,In_163);
or U345 (N_345,In_237,In_928);
nand U346 (N_346,In_817,In_463);
and U347 (N_347,In_753,In_390);
or U348 (N_348,In_849,In_401);
xnor U349 (N_349,In_880,In_509);
xor U350 (N_350,In_199,In_117);
nor U351 (N_351,In_646,In_599);
or U352 (N_352,In_852,In_456);
or U353 (N_353,In_508,In_865);
nor U354 (N_354,In_624,In_106);
and U355 (N_355,In_563,In_793);
nand U356 (N_356,In_98,In_567);
and U357 (N_357,In_747,In_253);
or U358 (N_358,In_683,In_633);
or U359 (N_359,In_374,In_519);
nor U360 (N_360,In_556,In_377);
nand U361 (N_361,In_834,In_724);
and U362 (N_362,In_380,In_205);
or U363 (N_363,In_187,In_895);
and U364 (N_364,In_458,In_53);
nand U365 (N_365,In_12,In_426);
and U366 (N_366,In_689,In_514);
nand U367 (N_367,In_28,In_256);
or U368 (N_368,In_105,In_487);
nand U369 (N_369,In_349,In_621);
nand U370 (N_370,In_60,In_551);
and U371 (N_371,In_231,In_308);
nor U372 (N_372,In_995,In_161);
and U373 (N_373,In_356,In_600);
nand U374 (N_374,In_460,In_743);
nor U375 (N_375,In_310,In_216);
nor U376 (N_376,In_272,In_178);
nor U377 (N_377,In_678,In_324);
nor U378 (N_378,In_95,In_113);
nor U379 (N_379,In_502,In_17);
and U380 (N_380,In_786,In_474);
nand U381 (N_381,In_335,In_968);
and U382 (N_382,In_176,In_241);
and U383 (N_383,In_957,In_483);
or U384 (N_384,In_500,In_425);
nor U385 (N_385,In_879,In_945);
or U386 (N_386,In_423,In_998);
nor U387 (N_387,In_962,In_417);
and U388 (N_388,In_822,In_932);
nor U389 (N_389,In_581,In_956);
nand U390 (N_390,In_62,In_597);
and U391 (N_391,In_389,In_438);
nor U392 (N_392,In_9,In_18);
or U393 (N_393,In_397,In_391);
nand U394 (N_394,In_750,In_921);
nor U395 (N_395,In_358,In_142);
nand U396 (N_396,In_325,In_411);
nand U397 (N_397,In_640,In_573);
nor U398 (N_398,In_737,In_622);
or U399 (N_399,In_78,In_804);
or U400 (N_400,In_713,In_294);
or U401 (N_401,In_644,In_982);
nor U402 (N_402,In_965,In_58);
nor U403 (N_403,In_482,In_208);
or U404 (N_404,In_51,In_537);
and U405 (N_405,In_742,In_251);
and U406 (N_406,In_558,In_395);
nand U407 (N_407,In_340,In_183);
or U408 (N_408,In_481,In_394);
or U409 (N_409,In_67,In_574);
or U410 (N_410,In_407,In_518);
nand U411 (N_411,In_860,In_719);
and U412 (N_412,In_972,In_99);
or U413 (N_413,In_973,In_798);
and U414 (N_414,In_812,In_136);
nor U415 (N_415,In_287,In_842);
nand U416 (N_416,In_430,In_232);
nor U417 (N_417,In_352,In_452);
nor U418 (N_418,In_997,In_175);
or U419 (N_419,In_329,In_87);
and U420 (N_420,In_868,In_434);
or U421 (N_421,In_805,In_76);
nand U422 (N_422,In_778,In_295);
nor U423 (N_423,In_108,In_594);
and U424 (N_424,In_730,In_590);
and U425 (N_425,In_800,In_829);
nand U426 (N_426,In_131,In_447);
nor U427 (N_427,In_171,In_586);
nor U428 (N_428,In_602,In_378);
nand U429 (N_429,In_507,In_577);
nor U430 (N_430,In_942,In_240);
nand U431 (N_431,In_799,In_418);
nand U432 (N_432,In_305,In_315);
nand U433 (N_433,In_478,In_655);
and U434 (N_434,In_278,In_271);
and U435 (N_435,In_838,In_248);
nand U436 (N_436,In_309,In_699);
nand U437 (N_437,In_235,In_190);
nor U438 (N_438,In_121,In_402);
or U439 (N_439,In_80,In_255);
or U440 (N_440,In_363,In_2);
nand U441 (N_441,In_328,In_578);
or U442 (N_442,In_907,In_491);
or U443 (N_443,In_994,In_148);
nor U444 (N_444,In_570,In_496);
and U445 (N_445,In_958,In_710);
and U446 (N_446,In_1,In_677);
nor U447 (N_447,In_36,In_144);
or U448 (N_448,In_228,In_845);
and U449 (N_449,In_331,In_138);
nor U450 (N_450,In_911,In_598);
and U451 (N_451,In_626,In_943);
and U452 (N_452,In_975,In_342);
nand U453 (N_453,In_66,In_780);
and U454 (N_454,In_206,In_59);
nand U455 (N_455,In_218,In_81);
nor U456 (N_456,In_607,In_839);
nand U457 (N_457,In_316,In_591);
xnor U458 (N_458,In_202,In_529);
nor U459 (N_459,In_139,In_717);
nor U460 (N_460,In_22,In_662);
and U461 (N_461,In_5,In_34);
nand U462 (N_462,In_542,In_189);
or U463 (N_463,In_565,In_857);
nor U464 (N_464,In_685,In_913);
nor U465 (N_465,In_831,In_587);
nor U466 (N_466,In_855,In_715);
nand U467 (N_467,In_88,In_285);
and U468 (N_468,In_472,In_462);
or U469 (N_469,In_620,In_731);
nand U470 (N_470,In_326,In_501);
nor U471 (N_471,In_824,In_544);
nor U472 (N_472,In_400,In_428);
xnor U473 (N_473,In_896,In_286);
nand U474 (N_474,In_14,In_83);
and U475 (N_475,In_129,In_672);
nor U476 (N_476,In_552,In_979);
or U477 (N_477,In_629,In_691);
or U478 (N_478,In_415,In_79);
or U479 (N_479,In_511,In_405);
nand U480 (N_480,In_969,In_416);
or U481 (N_481,In_164,In_334);
and U482 (N_482,In_167,In_373);
and U483 (N_483,In_386,In_270);
nand U484 (N_484,In_892,In_125);
nor U485 (N_485,In_718,In_91);
nor U486 (N_486,In_603,In_964);
nand U487 (N_487,In_179,In_746);
or U488 (N_488,In_247,In_877);
nor U489 (N_489,In_355,In_758);
nor U490 (N_490,In_967,In_657);
nand U491 (N_491,In_477,In_775);
and U492 (N_492,In_765,In_605);
and U493 (N_493,In_69,In_396);
or U494 (N_494,In_704,In_946);
nand U495 (N_495,In_118,In_990);
nor U496 (N_496,In_663,In_297);
or U497 (N_497,In_4,In_878);
and U498 (N_498,In_173,In_914);
nand U499 (N_499,In_174,In_803);
or U500 (N_500,In_712,In_598);
or U501 (N_501,In_285,In_644);
and U502 (N_502,In_454,In_436);
nand U503 (N_503,In_349,In_191);
or U504 (N_504,In_444,In_977);
or U505 (N_505,In_288,In_81);
nand U506 (N_506,In_400,In_103);
nand U507 (N_507,In_710,In_282);
or U508 (N_508,In_34,In_630);
nand U509 (N_509,In_171,In_275);
nor U510 (N_510,In_216,In_26);
and U511 (N_511,In_493,In_31);
nand U512 (N_512,In_806,In_170);
or U513 (N_513,In_255,In_540);
or U514 (N_514,In_905,In_716);
nand U515 (N_515,In_577,In_648);
and U516 (N_516,In_37,In_123);
and U517 (N_517,In_697,In_430);
nor U518 (N_518,In_804,In_322);
or U519 (N_519,In_51,In_398);
nand U520 (N_520,In_795,In_270);
nor U521 (N_521,In_522,In_275);
nand U522 (N_522,In_912,In_63);
nand U523 (N_523,In_758,In_788);
nand U524 (N_524,In_256,In_890);
nand U525 (N_525,In_320,In_585);
or U526 (N_526,In_516,In_802);
and U527 (N_527,In_835,In_671);
nor U528 (N_528,In_199,In_130);
or U529 (N_529,In_975,In_201);
nor U530 (N_530,In_824,In_929);
nor U531 (N_531,In_17,In_987);
or U532 (N_532,In_645,In_251);
and U533 (N_533,In_584,In_837);
nor U534 (N_534,In_436,In_561);
nor U535 (N_535,In_365,In_146);
or U536 (N_536,In_955,In_106);
nand U537 (N_537,In_627,In_914);
and U538 (N_538,In_55,In_41);
nand U539 (N_539,In_59,In_614);
and U540 (N_540,In_692,In_376);
and U541 (N_541,In_336,In_236);
or U542 (N_542,In_708,In_390);
nand U543 (N_543,In_896,In_973);
xnor U544 (N_544,In_162,In_178);
or U545 (N_545,In_507,In_145);
or U546 (N_546,In_26,In_551);
nor U547 (N_547,In_21,In_914);
or U548 (N_548,In_119,In_856);
nand U549 (N_549,In_854,In_815);
or U550 (N_550,In_671,In_850);
and U551 (N_551,In_192,In_647);
nand U552 (N_552,In_145,In_640);
nor U553 (N_553,In_137,In_555);
and U554 (N_554,In_536,In_828);
nand U555 (N_555,In_871,In_586);
nor U556 (N_556,In_984,In_78);
or U557 (N_557,In_417,In_491);
nor U558 (N_558,In_418,In_342);
or U559 (N_559,In_974,In_675);
or U560 (N_560,In_289,In_293);
or U561 (N_561,In_396,In_666);
nand U562 (N_562,In_444,In_211);
and U563 (N_563,In_737,In_536);
nand U564 (N_564,In_560,In_649);
and U565 (N_565,In_736,In_456);
and U566 (N_566,In_693,In_299);
nor U567 (N_567,In_861,In_279);
and U568 (N_568,In_642,In_85);
and U569 (N_569,In_949,In_601);
and U570 (N_570,In_877,In_889);
or U571 (N_571,In_321,In_804);
nand U572 (N_572,In_85,In_77);
nor U573 (N_573,In_217,In_198);
or U574 (N_574,In_586,In_705);
or U575 (N_575,In_30,In_374);
nor U576 (N_576,In_78,In_608);
nor U577 (N_577,In_732,In_30);
nor U578 (N_578,In_647,In_583);
nor U579 (N_579,In_920,In_711);
nand U580 (N_580,In_922,In_1);
nor U581 (N_581,In_662,In_782);
nand U582 (N_582,In_373,In_773);
or U583 (N_583,In_452,In_818);
nand U584 (N_584,In_175,In_918);
nor U585 (N_585,In_276,In_560);
nor U586 (N_586,In_601,In_428);
and U587 (N_587,In_757,In_974);
nand U588 (N_588,In_924,In_596);
or U589 (N_589,In_197,In_926);
nand U590 (N_590,In_846,In_106);
nand U591 (N_591,In_527,In_903);
and U592 (N_592,In_487,In_858);
nand U593 (N_593,In_418,In_560);
or U594 (N_594,In_410,In_145);
nand U595 (N_595,In_80,In_430);
nor U596 (N_596,In_810,In_221);
and U597 (N_597,In_476,In_266);
nand U598 (N_598,In_595,In_685);
and U599 (N_599,In_328,In_626);
nor U600 (N_600,In_698,In_178);
or U601 (N_601,In_723,In_446);
and U602 (N_602,In_429,In_742);
nand U603 (N_603,In_13,In_971);
and U604 (N_604,In_665,In_230);
nor U605 (N_605,In_191,In_180);
nor U606 (N_606,In_801,In_653);
and U607 (N_607,In_875,In_995);
xor U608 (N_608,In_406,In_2);
nor U609 (N_609,In_917,In_872);
nand U610 (N_610,In_963,In_397);
and U611 (N_611,In_541,In_648);
nor U612 (N_612,In_567,In_542);
and U613 (N_613,In_677,In_241);
or U614 (N_614,In_693,In_165);
nand U615 (N_615,In_186,In_915);
or U616 (N_616,In_544,In_963);
or U617 (N_617,In_462,In_781);
nand U618 (N_618,In_990,In_502);
or U619 (N_619,In_156,In_658);
nor U620 (N_620,In_824,In_212);
and U621 (N_621,In_70,In_322);
nand U622 (N_622,In_358,In_739);
nand U623 (N_623,In_188,In_856);
nor U624 (N_624,In_61,In_315);
nand U625 (N_625,In_209,In_689);
nand U626 (N_626,In_282,In_826);
nor U627 (N_627,In_344,In_52);
nand U628 (N_628,In_152,In_162);
nand U629 (N_629,In_401,In_892);
nor U630 (N_630,In_220,In_302);
nor U631 (N_631,In_379,In_122);
nor U632 (N_632,In_115,In_391);
nor U633 (N_633,In_495,In_800);
nor U634 (N_634,In_552,In_628);
and U635 (N_635,In_282,In_879);
nor U636 (N_636,In_783,In_499);
or U637 (N_637,In_988,In_829);
nand U638 (N_638,In_501,In_347);
or U639 (N_639,In_822,In_139);
or U640 (N_640,In_145,In_593);
nand U641 (N_641,In_684,In_365);
nand U642 (N_642,In_96,In_855);
and U643 (N_643,In_526,In_847);
or U644 (N_644,In_723,In_545);
nor U645 (N_645,In_446,In_883);
nor U646 (N_646,In_571,In_192);
and U647 (N_647,In_118,In_210);
nand U648 (N_648,In_550,In_994);
and U649 (N_649,In_779,In_853);
and U650 (N_650,In_837,In_836);
or U651 (N_651,In_302,In_758);
or U652 (N_652,In_222,In_260);
nand U653 (N_653,In_668,In_94);
nor U654 (N_654,In_828,In_519);
nor U655 (N_655,In_944,In_715);
and U656 (N_656,In_844,In_448);
nand U657 (N_657,In_687,In_769);
or U658 (N_658,In_122,In_271);
or U659 (N_659,In_248,In_117);
or U660 (N_660,In_207,In_249);
and U661 (N_661,In_569,In_672);
nor U662 (N_662,In_510,In_971);
nor U663 (N_663,In_108,In_754);
nor U664 (N_664,In_45,In_506);
or U665 (N_665,In_502,In_484);
or U666 (N_666,In_61,In_800);
and U667 (N_667,In_728,In_399);
nand U668 (N_668,In_380,In_802);
nand U669 (N_669,In_750,In_154);
and U670 (N_670,In_387,In_301);
and U671 (N_671,In_197,In_281);
nand U672 (N_672,In_646,In_554);
or U673 (N_673,In_419,In_248);
or U674 (N_674,In_349,In_503);
nand U675 (N_675,In_801,In_278);
and U676 (N_676,In_758,In_886);
nor U677 (N_677,In_323,In_105);
or U678 (N_678,In_605,In_436);
nand U679 (N_679,In_808,In_819);
nand U680 (N_680,In_346,In_432);
nand U681 (N_681,In_277,In_685);
or U682 (N_682,In_747,In_859);
and U683 (N_683,In_628,In_848);
and U684 (N_684,In_587,In_187);
nand U685 (N_685,In_794,In_645);
nor U686 (N_686,In_198,In_751);
and U687 (N_687,In_701,In_399);
and U688 (N_688,In_920,In_441);
and U689 (N_689,In_336,In_798);
or U690 (N_690,In_820,In_660);
and U691 (N_691,In_750,In_941);
nor U692 (N_692,In_877,In_221);
and U693 (N_693,In_685,In_844);
nand U694 (N_694,In_487,In_110);
nand U695 (N_695,In_355,In_997);
or U696 (N_696,In_7,In_251);
nand U697 (N_697,In_315,In_149);
and U698 (N_698,In_272,In_34);
and U699 (N_699,In_207,In_729);
nor U700 (N_700,In_603,In_422);
or U701 (N_701,In_428,In_916);
and U702 (N_702,In_100,In_496);
or U703 (N_703,In_759,In_66);
nand U704 (N_704,In_5,In_344);
and U705 (N_705,In_743,In_648);
and U706 (N_706,In_885,In_603);
and U707 (N_707,In_705,In_24);
nand U708 (N_708,In_193,In_673);
or U709 (N_709,In_217,In_278);
or U710 (N_710,In_481,In_650);
or U711 (N_711,In_600,In_681);
nand U712 (N_712,In_459,In_648);
nor U713 (N_713,In_428,In_91);
or U714 (N_714,In_88,In_364);
and U715 (N_715,In_90,In_380);
and U716 (N_716,In_941,In_723);
or U717 (N_717,In_832,In_476);
or U718 (N_718,In_216,In_345);
or U719 (N_719,In_55,In_791);
or U720 (N_720,In_585,In_339);
nor U721 (N_721,In_40,In_715);
and U722 (N_722,In_855,In_124);
nor U723 (N_723,In_440,In_323);
and U724 (N_724,In_559,In_757);
nor U725 (N_725,In_354,In_264);
or U726 (N_726,In_806,In_864);
xor U727 (N_727,In_392,In_350);
and U728 (N_728,In_30,In_252);
nand U729 (N_729,In_75,In_937);
or U730 (N_730,In_168,In_422);
nor U731 (N_731,In_625,In_465);
nor U732 (N_732,In_399,In_68);
or U733 (N_733,In_642,In_138);
nor U734 (N_734,In_185,In_308);
and U735 (N_735,In_909,In_770);
nor U736 (N_736,In_615,In_107);
or U737 (N_737,In_386,In_681);
or U738 (N_738,In_886,In_305);
or U739 (N_739,In_499,In_687);
and U740 (N_740,In_285,In_358);
nand U741 (N_741,In_862,In_537);
or U742 (N_742,In_550,In_95);
nor U743 (N_743,In_154,In_288);
or U744 (N_744,In_364,In_789);
xor U745 (N_745,In_438,In_948);
and U746 (N_746,In_226,In_500);
and U747 (N_747,In_510,In_790);
nand U748 (N_748,In_534,In_750);
nand U749 (N_749,In_814,In_741);
and U750 (N_750,In_480,In_999);
nor U751 (N_751,In_40,In_747);
and U752 (N_752,In_855,In_871);
nor U753 (N_753,In_326,In_90);
nand U754 (N_754,In_530,In_162);
and U755 (N_755,In_750,In_989);
and U756 (N_756,In_331,In_413);
nor U757 (N_757,In_713,In_759);
and U758 (N_758,In_397,In_5);
nand U759 (N_759,In_992,In_507);
nor U760 (N_760,In_489,In_937);
or U761 (N_761,In_839,In_185);
nor U762 (N_762,In_531,In_349);
nand U763 (N_763,In_239,In_293);
and U764 (N_764,In_629,In_237);
nor U765 (N_765,In_884,In_364);
nor U766 (N_766,In_776,In_341);
nor U767 (N_767,In_489,In_436);
or U768 (N_768,In_948,In_609);
or U769 (N_769,In_571,In_871);
nand U770 (N_770,In_18,In_553);
and U771 (N_771,In_429,In_462);
and U772 (N_772,In_517,In_935);
or U773 (N_773,In_780,In_572);
nand U774 (N_774,In_554,In_291);
or U775 (N_775,In_289,In_163);
nand U776 (N_776,In_352,In_50);
nor U777 (N_777,In_185,In_823);
nor U778 (N_778,In_998,In_589);
nand U779 (N_779,In_560,In_874);
nor U780 (N_780,In_168,In_919);
or U781 (N_781,In_955,In_224);
nand U782 (N_782,In_222,In_950);
or U783 (N_783,In_431,In_280);
or U784 (N_784,In_350,In_909);
and U785 (N_785,In_313,In_692);
nor U786 (N_786,In_235,In_506);
and U787 (N_787,In_760,In_668);
nand U788 (N_788,In_60,In_84);
and U789 (N_789,In_99,In_535);
or U790 (N_790,In_328,In_22);
or U791 (N_791,In_748,In_686);
and U792 (N_792,In_865,In_307);
or U793 (N_793,In_310,In_722);
nor U794 (N_794,In_879,In_624);
or U795 (N_795,In_559,In_844);
nand U796 (N_796,In_0,In_522);
nand U797 (N_797,In_435,In_978);
or U798 (N_798,In_842,In_438);
and U799 (N_799,In_582,In_820);
or U800 (N_800,In_571,In_504);
nor U801 (N_801,In_138,In_621);
nand U802 (N_802,In_724,In_635);
and U803 (N_803,In_870,In_945);
and U804 (N_804,In_964,In_521);
nor U805 (N_805,In_417,In_392);
or U806 (N_806,In_631,In_912);
or U807 (N_807,In_520,In_198);
nor U808 (N_808,In_639,In_920);
nor U809 (N_809,In_721,In_615);
or U810 (N_810,In_163,In_760);
nand U811 (N_811,In_77,In_881);
and U812 (N_812,In_725,In_554);
or U813 (N_813,In_779,In_8);
nor U814 (N_814,In_851,In_517);
and U815 (N_815,In_646,In_784);
nor U816 (N_816,In_917,In_649);
and U817 (N_817,In_307,In_133);
nor U818 (N_818,In_746,In_750);
nand U819 (N_819,In_476,In_763);
nand U820 (N_820,In_458,In_759);
and U821 (N_821,In_854,In_521);
or U822 (N_822,In_59,In_809);
and U823 (N_823,In_832,In_389);
nand U824 (N_824,In_518,In_452);
or U825 (N_825,In_648,In_634);
and U826 (N_826,In_866,In_494);
nand U827 (N_827,In_296,In_841);
nand U828 (N_828,In_997,In_699);
nor U829 (N_829,In_935,In_166);
nand U830 (N_830,In_973,In_792);
and U831 (N_831,In_607,In_561);
or U832 (N_832,In_789,In_299);
nand U833 (N_833,In_130,In_557);
or U834 (N_834,In_512,In_947);
and U835 (N_835,In_973,In_605);
nor U836 (N_836,In_721,In_532);
or U837 (N_837,In_991,In_375);
nor U838 (N_838,In_505,In_42);
nor U839 (N_839,In_836,In_468);
nor U840 (N_840,In_191,In_494);
or U841 (N_841,In_831,In_69);
nor U842 (N_842,In_650,In_521);
and U843 (N_843,In_856,In_395);
and U844 (N_844,In_163,In_780);
or U845 (N_845,In_469,In_933);
nand U846 (N_846,In_469,In_386);
nand U847 (N_847,In_588,In_290);
and U848 (N_848,In_318,In_757);
nor U849 (N_849,In_730,In_986);
nor U850 (N_850,In_556,In_72);
and U851 (N_851,In_615,In_969);
nand U852 (N_852,In_426,In_152);
nand U853 (N_853,In_215,In_701);
nand U854 (N_854,In_738,In_257);
or U855 (N_855,In_883,In_650);
nor U856 (N_856,In_484,In_956);
and U857 (N_857,In_792,In_811);
nor U858 (N_858,In_639,In_656);
nand U859 (N_859,In_954,In_226);
nor U860 (N_860,In_832,In_903);
or U861 (N_861,In_176,In_296);
nor U862 (N_862,In_92,In_337);
or U863 (N_863,In_804,In_928);
nor U864 (N_864,In_965,In_216);
nand U865 (N_865,In_106,In_35);
nor U866 (N_866,In_6,In_220);
or U867 (N_867,In_464,In_913);
nand U868 (N_868,In_521,In_289);
nand U869 (N_869,In_491,In_268);
nand U870 (N_870,In_671,In_304);
nand U871 (N_871,In_901,In_785);
nor U872 (N_872,In_977,In_227);
nand U873 (N_873,In_436,In_252);
or U874 (N_874,In_401,In_81);
nand U875 (N_875,In_988,In_828);
or U876 (N_876,In_624,In_972);
nor U877 (N_877,In_340,In_202);
and U878 (N_878,In_928,In_996);
nand U879 (N_879,In_361,In_931);
nand U880 (N_880,In_959,In_781);
nand U881 (N_881,In_730,In_523);
nand U882 (N_882,In_619,In_134);
nand U883 (N_883,In_383,In_0);
nor U884 (N_884,In_426,In_200);
nor U885 (N_885,In_665,In_324);
or U886 (N_886,In_995,In_745);
and U887 (N_887,In_493,In_808);
and U888 (N_888,In_569,In_572);
and U889 (N_889,In_159,In_870);
or U890 (N_890,In_656,In_27);
nor U891 (N_891,In_307,In_448);
or U892 (N_892,In_714,In_719);
nor U893 (N_893,In_974,In_758);
nor U894 (N_894,In_565,In_404);
nand U895 (N_895,In_562,In_840);
nor U896 (N_896,In_442,In_214);
or U897 (N_897,In_342,In_21);
nor U898 (N_898,In_328,In_908);
nor U899 (N_899,In_846,In_920);
nand U900 (N_900,In_324,In_607);
nand U901 (N_901,In_644,In_972);
or U902 (N_902,In_484,In_172);
and U903 (N_903,In_634,In_186);
nor U904 (N_904,In_86,In_502);
and U905 (N_905,In_423,In_885);
or U906 (N_906,In_38,In_677);
or U907 (N_907,In_850,In_476);
and U908 (N_908,In_658,In_418);
or U909 (N_909,In_792,In_934);
or U910 (N_910,In_46,In_457);
nor U911 (N_911,In_205,In_182);
or U912 (N_912,In_943,In_130);
or U913 (N_913,In_514,In_442);
and U914 (N_914,In_94,In_726);
or U915 (N_915,In_601,In_871);
or U916 (N_916,In_484,In_83);
nand U917 (N_917,In_363,In_802);
and U918 (N_918,In_398,In_87);
or U919 (N_919,In_868,In_385);
nor U920 (N_920,In_359,In_941);
nor U921 (N_921,In_111,In_204);
or U922 (N_922,In_603,In_22);
nor U923 (N_923,In_169,In_683);
or U924 (N_924,In_57,In_21);
and U925 (N_925,In_364,In_907);
or U926 (N_926,In_692,In_913);
nand U927 (N_927,In_560,In_957);
and U928 (N_928,In_790,In_38);
nand U929 (N_929,In_515,In_399);
nor U930 (N_930,In_598,In_261);
nor U931 (N_931,In_355,In_274);
and U932 (N_932,In_551,In_244);
nand U933 (N_933,In_104,In_724);
or U934 (N_934,In_406,In_359);
nor U935 (N_935,In_169,In_420);
and U936 (N_936,In_701,In_205);
nor U937 (N_937,In_710,In_612);
or U938 (N_938,In_674,In_963);
or U939 (N_939,In_318,In_607);
and U940 (N_940,In_579,In_715);
nand U941 (N_941,In_205,In_743);
and U942 (N_942,In_710,In_227);
nor U943 (N_943,In_654,In_978);
or U944 (N_944,In_492,In_277);
nand U945 (N_945,In_547,In_179);
nand U946 (N_946,In_506,In_497);
and U947 (N_947,In_548,In_332);
nor U948 (N_948,In_230,In_917);
and U949 (N_949,In_937,In_484);
or U950 (N_950,In_930,In_193);
or U951 (N_951,In_226,In_462);
and U952 (N_952,In_640,In_375);
nor U953 (N_953,In_927,In_446);
xnor U954 (N_954,In_18,In_713);
and U955 (N_955,In_19,In_385);
nand U956 (N_956,In_690,In_383);
nor U957 (N_957,In_614,In_635);
or U958 (N_958,In_820,In_926);
nand U959 (N_959,In_823,In_63);
nor U960 (N_960,In_858,In_532);
nor U961 (N_961,In_404,In_699);
and U962 (N_962,In_299,In_95);
nor U963 (N_963,In_482,In_368);
or U964 (N_964,In_557,In_629);
nor U965 (N_965,In_713,In_442);
and U966 (N_966,In_314,In_439);
or U967 (N_967,In_308,In_484);
and U968 (N_968,In_332,In_707);
and U969 (N_969,In_627,In_143);
and U970 (N_970,In_67,In_567);
or U971 (N_971,In_250,In_942);
or U972 (N_972,In_6,In_550);
nor U973 (N_973,In_358,In_303);
and U974 (N_974,In_344,In_890);
or U975 (N_975,In_300,In_5);
nand U976 (N_976,In_789,In_693);
nor U977 (N_977,In_915,In_618);
nand U978 (N_978,In_342,In_447);
or U979 (N_979,In_574,In_327);
or U980 (N_980,In_12,In_792);
or U981 (N_981,In_704,In_905);
or U982 (N_982,In_16,In_90);
and U983 (N_983,In_695,In_228);
nor U984 (N_984,In_661,In_50);
nand U985 (N_985,In_676,In_718);
xnor U986 (N_986,In_277,In_1);
and U987 (N_987,In_328,In_649);
and U988 (N_988,In_532,In_121);
nand U989 (N_989,In_521,In_551);
or U990 (N_990,In_261,In_763);
and U991 (N_991,In_360,In_609);
or U992 (N_992,In_791,In_706);
nand U993 (N_993,In_369,In_285);
and U994 (N_994,In_301,In_436);
or U995 (N_995,In_268,In_253);
or U996 (N_996,In_808,In_136);
nor U997 (N_997,In_518,In_35);
and U998 (N_998,In_228,In_130);
nor U999 (N_999,In_260,In_764);
or U1000 (N_1000,N_136,N_101);
nor U1001 (N_1001,N_871,N_691);
and U1002 (N_1002,N_803,N_397);
or U1003 (N_1003,N_353,N_654);
or U1004 (N_1004,N_374,N_234);
nor U1005 (N_1005,N_288,N_566);
nand U1006 (N_1006,N_729,N_9);
or U1007 (N_1007,N_138,N_980);
or U1008 (N_1008,N_994,N_559);
and U1009 (N_1009,N_960,N_200);
or U1010 (N_1010,N_574,N_61);
nand U1011 (N_1011,N_121,N_235);
nor U1012 (N_1012,N_689,N_528);
and U1013 (N_1013,N_529,N_252);
and U1014 (N_1014,N_216,N_752);
nand U1015 (N_1015,N_755,N_798);
or U1016 (N_1016,N_360,N_790);
nand U1017 (N_1017,N_756,N_440);
and U1018 (N_1018,N_761,N_912);
or U1019 (N_1019,N_572,N_351);
nor U1020 (N_1020,N_464,N_457);
and U1021 (N_1021,N_509,N_700);
nand U1022 (N_1022,N_639,N_818);
nand U1023 (N_1023,N_857,N_497);
nand U1024 (N_1024,N_77,N_88);
and U1025 (N_1025,N_224,N_949);
nand U1026 (N_1026,N_714,N_342);
nand U1027 (N_1027,N_106,N_609);
nand U1028 (N_1028,N_316,N_968);
nand U1029 (N_1029,N_807,N_370);
or U1030 (N_1030,N_791,N_105);
nand U1031 (N_1031,N_918,N_786);
nand U1032 (N_1032,N_157,N_991);
nand U1033 (N_1033,N_815,N_206);
nand U1034 (N_1034,N_886,N_21);
nand U1035 (N_1035,N_652,N_112);
nand U1036 (N_1036,N_178,N_45);
nand U1037 (N_1037,N_180,N_927);
or U1038 (N_1038,N_621,N_712);
and U1039 (N_1039,N_511,N_296);
nor U1040 (N_1040,N_472,N_820);
nor U1041 (N_1041,N_100,N_281);
nor U1042 (N_1042,N_211,N_212);
or U1043 (N_1043,N_760,N_867);
nor U1044 (N_1044,N_576,N_685);
nor U1045 (N_1045,N_114,N_615);
and U1046 (N_1046,N_40,N_320);
and U1047 (N_1047,N_856,N_629);
or U1048 (N_1048,N_631,N_148);
and U1049 (N_1049,N_362,N_801);
and U1050 (N_1050,N_185,N_644);
nand U1051 (N_1051,N_293,N_723);
and U1052 (N_1052,N_618,N_154);
or U1053 (N_1053,N_119,N_451);
and U1054 (N_1054,N_295,N_116);
or U1055 (N_1055,N_976,N_52);
nand U1056 (N_1056,N_584,N_699);
or U1057 (N_1057,N_326,N_606);
nor U1058 (N_1058,N_196,N_42);
or U1059 (N_1059,N_787,N_648);
or U1060 (N_1060,N_66,N_108);
nor U1061 (N_1061,N_27,N_89);
nand U1062 (N_1062,N_910,N_744);
or U1063 (N_1063,N_226,N_171);
or U1064 (N_1064,N_785,N_569);
nand U1065 (N_1065,N_284,N_937);
nand U1066 (N_1066,N_13,N_941);
or U1067 (N_1067,N_44,N_864);
and U1068 (N_1068,N_58,N_53);
and U1069 (N_1069,N_407,N_974);
or U1070 (N_1070,N_487,N_633);
nor U1071 (N_1071,N_596,N_953);
nand U1072 (N_1072,N_297,N_827);
nor U1073 (N_1073,N_728,N_20);
nor U1074 (N_1074,N_298,N_898);
nand U1075 (N_1075,N_907,N_388);
or U1076 (N_1076,N_855,N_726);
or U1077 (N_1077,N_406,N_670);
nand U1078 (N_1078,N_470,N_55);
nand U1079 (N_1079,N_938,N_378);
nor U1080 (N_1080,N_274,N_930);
and U1081 (N_1081,N_562,N_6);
or U1082 (N_1082,N_198,N_682);
nor U1083 (N_1083,N_462,N_738);
nand U1084 (N_1084,N_539,N_706);
nand U1085 (N_1085,N_425,N_436);
nand U1086 (N_1086,N_306,N_789);
and U1087 (N_1087,N_776,N_543);
nand U1088 (N_1088,N_804,N_906);
nor U1089 (N_1089,N_30,N_376);
and U1090 (N_1090,N_613,N_107);
or U1091 (N_1091,N_813,N_750);
and U1092 (N_1092,N_858,N_504);
nand U1093 (N_1093,N_533,N_552);
nand U1094 (N_1094,N_225,N_421);
and U1095 (N_1095,N_872,N_315);
and U1096 (N_1096,N_167,N_901);
and U1097 (N_1097,N_241,N_364);
or U1098 (N_1098,N_514,N_467);
and U1099 (N_1099,N_985,N_261);
nor U1100 (N_1100,N_657,N_430);
nand U1101 (N_1101,N_477,N_483);
nand U1102 (N_1102,N_76,N_242);
or U1103 (N_1103,N_173,N_501);
xnor U1104 (N_1104,N_109,N_35);
nand U1105 (N_1105,N_361,N_238);
nor U1106 (N_1106,N_961,N_939);
xor U1107 (N_1107,N_142,N_120);
xor U1108 (N_1108,N_377,N_730);
or U1109 (N_1109,N_704,N_630);
and U1110 (N_1110,N_493,N_190);
nor U1111 (N_1111,N_512,N_248);
nor U1112 (N_1112,N_160,N_184);
and U1113 (N_1113,N_954,N_589);
nand U1114 (N_1114,N_266,N_696);
nand U1115 (N_1115,N_688,N_932);
nor U1116 (N_1116,N_643,N_439);
or U1117 (N_1117,N_99,N_47);
nor U1118 (N_1118,N_545,N_159);
or U1119 (N_1119,N_127,N_597);
and U1120 (N_1120,N_193,N_846);
or U1121 (N_1121,N_135,N_740);
nor U1122 (N_1122,N_947,N_658);
or U1123 (N_1123,N_978,N_746);
and U1124 (N_1124,N_824,N_551);
nand U1125 (N_1125,N_967,N_302);
nand U1126 (N_1126,N_946,N_179);
or U1127 (N_1127,N_134,N_683);
or U1128 (N_1128,N_399,N_446);
and U1129 (N_1129,N_338,N_363);
nand U1130 (N_1130,N_331,N_877);
nor U1131 (N_1131,N_608,N_460);
nor U1132 (N_1132,N_458,N_664);
nor U1133 (N_1133,N_902,N_747);
xnor U1134 (N_1134,N_951,N_697);
nor U1135 (N_1135,N_94,N_117);
nor U1136 (N_1136,N_349,N_301);
nor U1137 (N_1137,N_911,N_727);
and U1138 (N_1138,N_384,N_510);
nand U1139 (N_1139,N_246,N_369);
or U1140 (N_1140,N_853,N_152);
nor U1141 (N_1141,N_847,N_616);
nand U1142 (N_1142,N_133,N_659);
and U1143 (N_1143,N_928,N_229);
and U1144 (N_1144,N_395,N_716);
nand U1145 (N_1145,N_817,N_161);
nand U1146 (N_1146,N_259,N_802);
or U1147 (N_1147,N_2,N_531);
xor U1148 (N_1148,N_565,N_836);
nand U1149 (N_1149,N_808,N_724);
nand U1150 (N_1150,N_526,N_656);
nor U1151 (N_1151,N_278,N_764);
nor U1152 (N_1152,N_110,N_422);
and U1153 (N_1153,N_23,N_972);
or U1154 (N_1154,N_347,N_41);
or U1155 (N_1155,N_875,N_577);
and U1156 (N_1156,N_359,N_917);
nand U1157 (N_1157,N_158,N_903);
and U1158 (N_1158,N_722,N_299);
and U1159 (N_1159,N_948,N_769);
nand U1160 (N_1160,N_390,N_313);
nor U1161 (N_1161,N_494,N_758);
nand U1162 (N_1162,N_996,N_309);
nor U1163 (N_1163,N_908,N_254);
nor U1164 (N_1164,N_228,N_516);
nor U1165 (N_1165,N_892,N_197);
nand U1166 (N_1166,N_168,N_38);
and U1167 (N_1167,N_703,N_93);
or U1168 (N_1168,N_524,N_926);
nand U1169 (N_1169,N_289,N_398);
nor U1170 (N_1170,N_29,N_610);
or U1171 (N_1171,N_128,N_486);
and U1172 (N_1172,N_835,N_262);
nand U1173 (N_1173,N_466,N_191);
and U1174 (N_1174,N_219,N_794);
or U1175 (N_1175,N_805,N_253);
nor U1176 (N_1176,N_50,N_721);
nand U1177 (N_1177,N_78,N_247);
nand U1178 (N_1178,N_417,N_409);
nor U1179 (N_1179,N_651,N_371);
or U1180 (N_1180,N_445,N_999);
nand U1181 (N_1181,N_595,N_325);
or U1182 (N_1182,N_958,N_263);
and U1183 (N_1183,N_777,N_373);
nor U1184 (N_1184,N_209,N_952);
or U1185 (N_1185,N_593,N_291);
nand U1186 (N_1186,N_251,N_690);
or U1187 (N_1187,N_957,N_583);
nor U1188 (N_1188,N_12,N_594);
nand U1189 (N_1189,N_336,N_736);
nor U1190 (N_1190,N_669,N_43);
or U1191 (N_1191,N_970,N_969);
nor U1192 (N_1192,N_207,N_715);
or U1193 (N_1193,N_640,N_602);
nand U1194 (N_1194,N_98,N_324);
and U1195 (N_1195,N_662,N_232);
and U1196 (N_1196,N_626,N_201);
and U1197 (N_1197,N_69,N_268);
nor U1198 (N_1198,N_186,N_205);
or U1199 (N_1199,N_177,N_753);
nor U1200 (N_1200,N_541,N_144);
and U1201 (N_1201,N_895,N_64);
nor U1202 (N_1202,N_402,N_778);
and U1203 (N_1203,N_290,N_357);
or U1204 (N_1204,N_122,N_863);
or U1205 (N_1205,N_677,N_940);
or U1206 (N_1206,N_719,N_468);
nor U1207 (N_1207,N_694,N_904);
nand U1208 (N_1208,N_146,N_705);
nor U1209 (N_1209,N_775,N_459);
and U1210 (N_1210,N_202,N_894);
nor U1211 (N_1211,N_702,N_540);
and U1212 (N_1212,N_893,N_661);
nor U1213 (N_1213,N_498,N_544);
or U1214 (N_1214,N_304,N_327);
and U1215 (N_1215,N_882,N_739);
and U1216 (N_1216,N_950,N_708);
nand U1217 (N_1217,N_768,N_95);
nor U1218 (N_1218,N_427,N_646);
or U1219 (N_1219,N_341,N_18);
nor U1220 (N_1220,N_401,N_575);
and U1221 (N_1221,N_878,N_812);
or U1222 (N_1222,N_271,N_130);
or U1223 (N_1223,N_772,N_84);
nand U1224 (N_1224,N_375,N_998);
nor U1225 (N_1225,N_624,N_264);
or U1226 (N_1226,N_780,N_392);
nor U1227 (N_1227,N_558,N_774);
nor U1228 (N_1228,N_617,N_51);
or U1229 (N_1229,N_779,N_33);
and U1230 (N_1230,N_233,N_461);
nor U1231 (N_1231,N_665,N_346);
nor U1232 (N_1232,N_517,N_275);
nor U1233 (N_1233,N_17,N_308);
and U1234 (N_1234,N_332,N_506);
nor U1235 (N_1235,N_410,N_891);
or U1236 (N_1236,N_834,N_428);
or U1237 (N_1237,N_416,N_46);
nor U1238 (N_1238,N_356,N_3);
nand U1239 (N_1239,N_538,N_150);
nand U1240 (N_1240,N_424,N_86);
nand U1241 (N_1241,N_698,N_632);
nand U1242 (N_1242,N_366,N_455);
and U1243 (N_1243,N_34,N_580);
and U1244 (N_1244,N_75,N_521);
or U1245 (N_1245,N_623,N_300);
or U1246 (N_1246,N_438,N_591);
and U1247 (N_1247,N_634,N_605);
nand U1248 (N_1248,N_496,N_387);
nor U1249 (N_1249,N_260,N_124);
or U1250 (N_1250,N_979,N_345);
nand U1251 (N_1251,N_841,N_273);
or U1252 (N_1252,N_221,N_965);
or U1253 (N_1253,N_490,N_434);
or U1254 (N_1254,N_245,N_710);
or U1255 (N_1255,N_426,N_879);
and U1256 (N_1256,N_563,N_63);
nor U1257 (N_1257,N_667,N_125);
nand U1258 (N_1258,N_203,N_810);
or U1259 (N_1259,N_170,N_82);
nand U1260 (N_1260,N_435,N_310);
or U1261 (N_1261,N_4,N_389);
nand U1262 (N_1262,N_329,N_492);
or U1263 (N_1263,N_905,N_537);
nand U1264 (N_1264,N_223,N_687);
and U1265 (N_1265,N_335,N_862);
or U1266 (N_1266,N_535,N_213);
and U1267 (N_1267,N_548,N_874);
nor U1268 (N_1268,N_480,N_60);
or U1269 (N_1269,N_317,N_581);
and U1270 (N_1270,N_532,N_307);
or U1271 (N_1271,N_321,N_782);
nand U1272 (N_1272,N_485,N_649);
and U1273 (N_1273,N_311,N_408);
and U1274 (N_1274,N_79,N_603);
nor U1275 (N_1275,N_981,N_720);
nand U1276 (N_1276,N_837,N_823);
nand U1277 (N_1277,N_795,N_731);
nand U1278 (N_1278,N_192,N_352);
nor U1279 (N_1279,N_151,N_411);
or U1280 (N_1280,N_230,N_187);
nor U1281 (N_1281,N_169,N_627);
nor U1282 (N_1282,N_391,N_783);
or U1283 (N_1283,N_312,N_448);
or U1284 (N_1284,N_607,N_923);
or U1285 (N_1285,N_70,N_92);
or U1286 (N_1286,N_734,N_415);
nand U1287 (N_1287,N_842,N_884);
nand U1288 (N_1288,N_925,N_239);
xor U1289 (N_1289,N_866,N_921);
nand U1290 (N_1290,N_592,N_97);
nor U1291 (N_1291,N_896,N_934);
and U1292 (N_1292,N_636,N_612);
and U1293 (N_1293,N_816,N_141);
xor U1294 (N_1294,N_587,N_959);
nand U1295 (N_1295,N_412,N_989);
nand U1296 (N_1296,N_484,N_619);
and U1297 (N_1297,N_887,N_358);
and U1298 (N_1298,N_839,N_379);
or U1299 (N_1299,N_255,N_85);
nand U1300 (N_1300,N_437,N_220);
and U1301 (N_1301,N_956,N_249);
and U1302 (N_1302,N_527,N_81);
nand U1303 (N_1303,N_936,N_383);
nand U1304 (N_1304,N_11,N_145);
nor U1305 (N_1305,N_328,N_831);
nor U1306 (N_1306,N_67,N_5);
and U1307 (N_1307,N_14,N_573);
nor U1308 (N_1308,N_876,N_988);
and U1309 (N_1309,N_924,N_671);
and U1310 (N_1310,N_861,N_215);
or U1311 (N_1311,N_733,N_265);
nand U1312 (N_1312,N_294,N_505);
and U1313 (N_1313,N_10,N_344);
nor U1314 (N_1314,N_873,N_172);
nor U1315 (N_1315,N_993,N_681);
and U1316 (N_1316,N_919,N_943);
or U1317 (N_1317,N_256,N_1);
or U1318 (N_1318,N_986,N_258);
or U1319 (N_1319,N_793,N_821);
or U1320 (N_1320,N_515,N_56);
nor U1321 (N_1321,N_285,N_319);
and U1322 (N_1322,N_393,N_257);
nor U1323 (N_1323,N_323,N_741);
nand U1324 (N_1324,N_851,N_453);
or U1325 (N_1325,N_982,N_865);
or U1326 (N_1326,N_582,N_870);
nand U1327 (N_1327,N_564,N_642);
or U1328 (N_1328,N_24,N_104);
or U1329 (N_1329,N_784,N_814);
nand U1330 (N_1330,N_118,N_554);
or U1331 (N_1331,N_183,N_72);
or U1332 (N_1332,N_600,N_549);
nor U1333 (N_1333,N_975,N_711);
nor U1334 (N_1334,N_195,N_123);
or U1335 (N_1335,N_641,N_394);
and U1336 (N_1336,N_611,N_149);
nand U1337 (N_1337,N_707,N_550);
nand U1338 (N_1338,N_713,N_513);
or U1339 (N_1339,N_181,N_604);
nand U1340 (N_1340,N_447,N_718);
or U1341 (N_1341,N_236,N_165);
or U1342 (N_1342,N_175,N_748);
nor U1343 (N_1343,N_396,N_49);
or U1344 (N_1344,N_283,N_279);
nor U1345 (N_1345,N_983,N_920);
nand U1346 (N_1346,N_588,N_287);
nand U1347 (N_1347,N_162,N_322);
nor U1348 (N_1348,N_337,N_508);
or U1349 (N_1349,N_267,N_931);
and U1350 (N_1350,N_742,N_343);
and U1351 (N_1351,N_71,N_432);
nor U1352 (N_1352,N_751,N_303);
nor U1353 (N_1353,N_773,N_759);
nor U1354 (N_1354,N_19,N_809);
nor U1355 (N_1355,N_429,N_922);
and U1356 (N_1356,N_869,N_822);
nor U1357 (N_1357,N_139,N_800);
nand U1358 (N_1358,N_479,N_59);
or U1359 (N_1359,N_771,N_502);
and U1360 (N_1360,N_111,N_914);
nand U1361 (N_1361,N_990,N_971);
nand U1362 (N_1362,N_8,N_880);
or U1363 (N_1363,N_163,N_227);
nand U1364 (N_1364,N_96,N_889);
and U1365 (N_1365,N_717,N_944);
or U1366 (N_1366,N_153,N_339);
nand U1367 (N_1367,N_763,N_860);
and U1368 (N_1368,N_26,N_405);
nand U1369 (N_1369,N_614,N_481);
or U1370 (N_1370,N_214,N_80);
and U1371 (N_1371,N_767,N_292);
nor U1372 (N_1372,N_132,N_489);
or U1373 (N_1373,N_156,N_131);
nor U1374 (N_1374,N_385,N_825);
nand U1375 (N_1375,N_330,N_828);
and U1376 (N_1376,N_442,N_909);
and U1377 (N_1377,N_579,N_663);
nand U1378 (N_1378,N_799,N_672);
nor U1379 (N_1379,N_680,N_964);
or U1380 (N_1380,N_868,N_849);
or U1381 (N_1381,N_913,N_272);
or U1382 (N_1382,N_546,N_792);
nand U1383 (N_1383,N_68,N_276);
or U1384 (N_1384,N_334,N_126);
xor U1385 (N_1385,N_547,N_571);
nand U1386 (N_1386,N_354,N_585);
nor U1387 (N_1387,N_91,N_586);
nor U1388 (N_1388,N_456,N_890);
and U1389 (N_1389,N_386,N_113);
nand U1390 (N_1390,N_244,N_622);
nor U1391 (N_1391,N_984,N_955);
nor U1392 (N_1392,N_743,N_668);
nand U1393 (N_1393,N_25,N_557);
and U1394 (N_1394,N_188,N_488);
and U1395 (N_1395,N_819,N_655);
and U1396 (N_1396,N_250,N_83);
and U1397 (N_1397,N_977,N_348);
nor U1398 (N_1398,N_693,N_507);
and U1399 (N_1399,N_525,N_843);
or U1400 (N_1400,N_852,N_666);
or U1401 (N_1401,N_590,N_478);
nor U1402 (N_1402,N_473,N_567);
nor U1403 (N_1403,N_465,N_482);
or U1404 (N_1404,N_73,N_915);
nor U1405 (N_1405,N_598,N_217);
and U1406 (N_1406,N_555,N_520);
nor U1407 (N_1407,N_176,N_844);
or U1408 (N_1408,N_491,N_676);
nand U1409 (N_1409,N_218,N_103);
nor U1410 (N_1410,N_935,N_553);
nor U1411 (N_1411,N_945,N_845);
nand U1412 (N_1412,N_305,N_471);
nor U1413 (N_1413,N_403,N_37);
nor U1414 (N_1414,N_899,N_32);
nand U1415 (N_1415,N_365,N_916);
and U1416 (N_1416,N_423,N_859);
and U1417 (N_1417,N_413,N_647);
and U1418 (N_1418,N_174,N_854);
or U1419 (N_1419,N_499,N_966);
nand U1420 (N_1420,N_270,N_282);
nand U1421 (N_1421,N_709,N_770);
nand U1422 (N_1422,N_942,N_765);
and U1423 (N_1423,N_420,N_692);
and U1424 (N_1424,N_443,N_645);
nand U1425 (N_1425,N_635,N_476);
and U1426 (N_1426,N_686,N_962);
or U1427 (N_1427,N_65,N_102);
and U1428 (N_1428,N_660,N_137);
nand U1429 (N_1429,N_54,N_237);
and U1430 (N_1430,N_368,N_995);
nor U1431 (N_1431,N_380,N_929);
nand U1432 (N_1432,N_382,N_796);
nand U1433 (N_1433,N_519,N_829);
or U1434 (N_1434,N_637,N_15);
nand U1435 (N_1435,N_367,N_673);
or U1436 (N_1436,N_140,N_208);
nor U1437 (N_1437,N_900,N_431);
nor U1438 (N_1438,N_333,N_701);
and U1439 (N_1439,N_28,N_318);
and U1440 (N_1440,N_556,N_534);
and U1441 (N_1441,N_450,N_240);
nand U1442 (N_1442,N_599,N_749);
nand U1443 (N_1443,N_36,N_523);
nor U1444 (N_1444,N_62,N_39);
nor U1445 (N_1445,N_474,N_650);
nand U1446 (N_1446,N_832,N_675);
and U1447 (N_1447,N_90,N_269);
nand U1448 (N_1448,N_578,N_848);
or U1449 (N_1449,N_57,N_143);
nor U1450 (N_1450,N_570,N_452);
nand U1451 (N_1451,N_475,N_0);
or U1452 (N_1452,N_314,N_204);
and U1453 (N_1453,N_48,N_419);
nand U1454 (N_1454,N_115,N_530);
and U1455 (N_1455,N_222,N_781);
nand U1456 (N_1456,N_963,N_826);
or U1457 (N_1457,N_933,N_883);
or U1458 (N_1458,N_638,N_766);
nor U1459 (N_1459,N_418,N_286);
or U1460 (N_1460,N_400,N_164);
nor U1461 (N_1461,N_735,N_74);
or U1462 (N_1462,N_7,N_561);
nor U1463 (N_1463,N_355,N_987);
nor U1464 (N_1464,N_973,N_381);
and U1465 (N_1465,N_732,N_850);
nor U1466 (N_1466,N_87,N_155);
and U1467 (N_1467,N_182,N_881);
or U1468 (N_1468,N_189,N_522);
nor U1469 (N_1469,N_147,N_463);
and U1470 (N_1470,N_754,N_811);
nor U1471 (N_1471,N_725,N_16);
xnor U1472 (N_1472,N_568,N_678);
or U1473 (N_1473,N_830,N_231);
or U1474 (N_1474,N_684,N_806);
and U1475 (N_1475,N_199,N_674);
and U1476 (N_1476,N_620,N_454);
or U1477 (N_1477,N_992,N_441);
or U1478 (N_1478,N_840,N_745);
and U1479 (N_1479,N_757,N_838);
and U1480 (N_1480,N_166,N_449);
or U1481 (N_1481,N_194,N_737);
and U1482 (N_1482,N_762,N_536);
nand U1483 (N_1483,N_560,N_129);
nand U1484 (N_1484,N_503,N_833);
nand U1485 (N_1485,N_625,N_679);
nand U1486 (N_1486,N_695,N_797);
and U1487 (N_1487,N_518,N_22);
and U1488 (N_1488,N_210,N_500);
nor U1489 (N_1489,N_888,N_444);
and U1490 (N_1490,N_601,N_885);
or U1491 (N_1491,N_414,N_243);
or U1492 (N_1492,N_277,N_372);
or U1493 (N_1493,N_542,N_495);
and U1494 (N_1494,N_404,N_628);
nand U1495 (N_1495,N_433,N_31);
or U1496 (N_1496,N_469,N_340);
nor U1497 (N_1497,N_897,N_280);
nor U1498 (N_1498,N_653,N_788);
and U1499 (N_1499,N_997,N_350);
nor U1500 (N_1500,N_85,N_734);
nor U1501 (N_1501,N_258,N_444);
nor U1502 (N_1502,N_836,N_537);
and U1503 (N_1503,N_514,N_763);
and U1504 (N_1504,N_555,N_515);
and U1505 (N_1505,N_958,N_347);
nand U1506 (N_1506,N_200,N_996);
or U1507 (N_1507,N_609,N_136);
and U1508 (N_1508,N_426,N_847);
nand U1509 (N_1509,N_463,N_772);
nor U1510 (N_1510,N_806,N_328);
nand U1511 (N_1511,N_304,N_363);
or U1512 (N_1512,N_245,N_165);
and U1513 (N_1513,N_519,N_112);
and U1514 (N_1514,N_822,N_683);
and U1515 (N_1515,N_524,N_157);
nor U1516 (N_1516,N_617,N_395);
nand U1517 (N_1517,N_522,N_20);
nand U1518 (N_1518,N_455,N_546);
and U1519 (N_1519,N_570,N_723);
nand U1520 (N_1520,N_128,N_672);
nor U1521 (N_1521,N_291,N_167);
nand U1522 (N_1522,N_162,N_782);
or U1523 (N_1523,N_549,N_350);
and U1524 (N_1524,N_94,N_992);
nand U1525 (N_1525,N_564,N_986);
xor U1526 (N_1526,N_293,N_848);
or U1527 (N_1527,N_394,N_246);
or U1528 (N_1528,N_362,N_593);
nand U1529 (N_1529,N_670,N_177);
xnor U1530 (N_1530,N_409,N_941);
nor U1531 (N_1531,N_403,N_247);
nand U1532 (N_1532,N_96,N_814);
or U1533 (N_1533,N_793,N_152);
and U1534 (N_1534,N_202,N_984);
and U1535 (N_1535,N_186,N_766);
and U1536 (N_1536,N_722,N_889);
or U1537 (N_1537,N_196,N_741);
and U1538 (N_1538,N_43,N_564);
or U1539 (N_1539,N_112,N_753);
nor U1540 (N_1540,N_657,N_313);
nor U1541 (N_1541,N_10,N_269);
nor U1542 (N_1542,N_606,N_380);
and U1543 (N_1543,N_505,N_105);
or U1544 (N_1544,N_412,N_818);
or U1545 (N_1545,N_878,N_165);
nand U1546 (N_1546,N_698,N_343);
nand U1547 (N_1547,N_792,N_364);
and U1548 (N_1548,N_637,N_405);
and U1549 (N_1549,N_115,N_583);
and U1550 (N_1550,N_268,N_82);
nor U1551 (N_1551,N_693,N_813);
or U1552 (N_1552,N_460,N_595);
nand U1553 (N_1553,N_220,N_851);
xnor U1554 (N_1554,N_148,N_412);
xor U1555 (N_1555,N_531,N_730);
nand U1556 (N_1556,N_921,N_492);
or U1557 (N_1557,N_924,N_351);
and U1558 (N_1558,N_416,N_330);
nor U1559 (N_1559,N_721,N_479);
and U1560 (N_1560,N_498,N_604);
or U1561 (N_1561,N_272,N_698);
nor U1562 (N_1562,N_113,N_806);
nand U1563 (N_1563,N_739,N_359);
and U1564 (N_1564,N_899,N_644);
or U1565 (N_1565,N_174,N_375);
and U1566 (N_1566,N_839,N_206);
nand U1567 (N_1567,N_494,N_482);
and U1568 (N_1568,N_293,N_692);
nand U1569 (N_1569,N_451,N_351);
nor U1570 (N_1570,N_501,N_892);
or U1571 (N_1571,N_254,N_51);
and U1572 (N_1572,N_425,N_846);
nor U1573 (N_1573,N_2,N_232);
nand U1574 (N_1574,N_699,N_852);
nand U1575 (N_1575,N_630,N_857);
or U1576 (N_1576,N_735,N_424);
and U1577 (N_1577,N_545,N_1);
and U1578 (N_1578,N_783,N_408);
nor U1579 (N_1579,N_451,N_343);
nand U1580 (N_1580,N_255,N_781);
nor U1581 (N_1581,N_22,N_491);
or U1582 (N_1582,N_875,N_785);
nor U1583 (N_1583,N_926,N_433);
or U1584 (N_1584,N_955,N_63);
and U1585 (N_1585,N_86,N_183);
or U1586 (N_1586,N_340,N_314);
nor U1587 (N_1587,N_576,N_200);
nor U1588 (N_1588,N_320,N_415);
or U1589 (N_1589,N_258,N_498);
nand U1590 (N_1590,N_449,N_520);
or U1591 (N_1591,N_404,N_597);
nand U1592 (N_1592,N_818,N_63);
nand U1593 (N_1593,N_259,N_438);
and U1594 (N_1594,N_734,N_440);
or U1595 (N_1595,N_486,N_310);
or U1596 (N_1596,N_203,N_283);
and U1597 (N_1597,N_354,N_191);
or U1598 (N_1598,N_362,N_348);
nand U1599 (N_1599,N_681,N_965);
or U1600 (N_1600,N_288,N_865);
nand U1601 (N_1601,N_310,N_398);
and U1602 (N_1602,N_817,N_364);
nand U1603 (N_1603,N_316,N_249);
xor U1604 (N_1604,N_130,N_125);
nand U1605 (N_1605,N_878,N_919);
and U1606 (N_1606,N_830,N_753);
nand U1607 (N_1607,N_286,N_846);
and U1608 (N_1608,N_844,N_23);
nand U1609 (N_1609,N_925,N_686);
nand U1610 (N_1610,N_866,N_433);
nor U1611 (N_1611,N_616,N_838);
or U1612 (N_1612,N_125,N_320);
nor U1613 (N_1613,N_138,N_584);
and U1614 (N_1614,N_417,N_820);
and U1615 (N_1615,N_788,N_873);
and U1616 (N_1616,N_124,N_658);
and U1617 (N_1617,N_776,N_542);
or U1618 (N_1618,N_322,N_791);
nand U1619 (N_1619,N_321,N_144);
and U1620 (N_1620,N_781,N_551);
nor U1621 (N_1621,N_707,N_250);
or U1622 (N_1622,N_657,N_532);
nand U1623 (N_1623,N_823,N_55);
or U1624 (N_1624,N_278,N_753);
and U1625 (N_1625,N_395,N_892);
or U1626 (N_1626,N_764,N_723);
nand U1627 (N_1627,N_674,N_284);
nand U1628 (N_1628,N_974,N_871);
or U1629 (N_1629,N_952,N_509);
nand U1630 (N_1630,N_430,N_172);
nand U1631 (N_1631,N_564,N_546);
nand U1632 (N_1632,N_425,N_774);
nor U1633 (N_1633,N_402,N_109);
and U1634 (N_1634,N_579,N_234);
and U1635 (N_1635,N_58,N_633);
xnor U1636 (N_1636,N_559,N_537);
nand U1637 (N_1637,N_517,N_767);
or U1638 (N_1638,N_651,N_899);
nor U1639 (N_1639,N_0,N_685);
and U1640 (N_1640,N_54,N_945);
and U1641 (N_1641,N_577,N_597);
nand U1642 (N_1642,N_912,N_144);
or U1643 (N_1643,N_104,N_849);
or U1644 (N_1644,N_838,N_124);
and U1645 (N_1645,N_630,N_135);
nand U1646 (N_1646,N_511,N_891);
or U1647 (N_1647,N_429,N_97);
and U1648 (N_1648,N_927,N_895);
and U1649 (N_1649,N_723,N_558);
nor U1650 (N_1650,N_179,N_420);
nand U1651 (N_1651,N_268,N_259);
nor U1652 (N_1652,N_294,N_677);
and U1653 (N_1653,N_364,N_655);
and U1654 (N_1654,N_671,N_852);
and U1655 (N_1655,N_626,N_384);
xnor U1656 (N_1656,N_853,N_32);
or U1657 (N_1657,N_694,N_996);
nand U1658 (N_1658,N_427,N_134);
and U1659 (N_1659,N_23,N_633);
and U1660 (N_1660,N_481,N_887);
and U1661 (N_1661,N_158,N_572);
or U1662 (N_1662,N_760,N_223);
and U1663 (N_1663,N_91,N_4);
and U1664 (N_1664,N_120,N_143);
and U1665 (N_1665,N_959,N_613);
and U1666 (N_1666,N_787,N_243);
and U1667 (N_1667,N_403,N_628);
and U1668 (N_1668,N_123,N_3);
nor U1669 (N_1669,N_212,N_766);
nand U1670 (N_1670,N_0,N_656);
nand U1671 (N_1671,N_362,N_122);
nor U1672 (N_1672,N_121,N_457);
nor U1673 (N_1673,N_961,N_417);
or U1674 (N_1674,N_773,N_626);
or U1675 (N_1675,N_839,N_382);
and U1676 (N_1676,N_114,N_542);
or U1677 (N_1677,N_649,N_110);
xor U1678 (N_1678,N_529,N_461);
xor U1679 (N_1679,N_139,N_707);
nor U1680 (N_1680,N_572,N_209);
or U1681 (N_1681,N_785,N_867);
or U1682 (N_1682,N_949,N_73);
or U1683 (N_1683,N_336,N_816);
or U1684 (N_1684,N_278,N_15);
nand U1685 (N_1685,N_427,N_530);
and U1686 (N_1686,N_331,N_814);
or U1687 (N_1687,N_583,N_292);
or U1688 (N_1688,N_0,N_841);
and U1689 (N_1689,N_404,N_746);
or U1690 (N_1690,N_914,N_298);
nor U1691 (N_1691,N_628,N_618);
or U1692 (N_1692,N_340,N_632);
and U1693 (N_1693,N_779,N_57);
and U1694 (N_1694,N_527,N_861);
nand U1695 (N_1695,N_988,N_751);
or U1696 (N_1696,N_386,N_191);
or U1697 (N_1697,N_113,N_104);
or U1698 (N_1698,N_891,N_50);
and U1699 (N_1699,N_217,N_814);
nor U1700 (N_1700,N_205,N_227);
nand U1701 (N_1701,N_377,N_670);
nor U1702 (N_1702,N_65,N_478);
and U1703 (N_1703,N_361,N_523);
nor U1704 (N_1704,N_234,N_178);
or U1705 (N_1705,N_414,N_900);
and U1706 (N_1706,N_681,N_39);
and U1707 (N_1707,N_728,N_775);
and U1708 (N_1708,N_486,N_847);
or U1709 (N_1709,N_244,N_524);
or U1710 (N_1710,N_808,N_226);
nor U1711 (N_1711,N_255,N_390);
nor U1712 (N_1712,N_880,N_403);
nand U1713 (N_1713,N_158,N_524);
nor U1714 (N_1714,N_250,N_382);
nor U1715 (N_1715,N_618,N_551);
nand U1716 (N_1716,N_218,N_828);
and U1717 (N_1717,N_169,N_780);
and U1718 (N_1718,N_291,N_491);
nor U1719 (N_1719,N_894,N_742);
and U1720 (N_1720,N_551,N_730);
nand U1721 (N_1721,N_54,N_450);
nor U1722 (N_1722,N_312,N_774);
nor U1723 (N_1723,N_987,N_301);
nor U1724 (N_1724,N_956,N_5);
and U1725 (N_1725,N_726,N_731);
and U1726 (N_1726,N_817,N_747);
nand U1727 (N_1727,N_380,N_432);
nor U1728 (N_1728,N_95,N_576);
or U1729 (N_1729,N_312,N_550);
or U1730 (N_1730,N_73,N_666);
nand U1731 (N_1731,N_191,N_142);
or U1732 (N_1732,N_373,N_709);
and U1733 (N_1733,N_845,N_853);
nand U1734 (N_1734,N_95,N_347);
and U1735 (N_1735,N_289,N_880);
nor U1736 (N_1736,N_721,N_251);
nand U1737 (N_1737,N_802,N_780);
and U1738 (N_1738,N_90,N_666);
nor U1739 (N_1739,N_104,N_588);
or U1740 (N_1740,N_585,N_417);
xor U1741 (N_1741,N_881,N_556);
and U1742 (N_1742,N_454,N_524);
or U1743 (N_1743,N_59,N_252);
or U1744 (N_1744,N_106,N_306);
or U1745 (N_1745,N_253,N_270);
nand U1746 (N_1746,N_987,N_19);
nor U1747 (N_1747,N_961,N_562);
and U1748 (N_1748,N_570,N_1);
and U1749 (N_1749,N_901,N_470);
nand U1750 (N_1750,N_69,N_832);
and U1751 (N_1751,N_374,N_121);
nand U1752 (N_1752,N_255,N_89);
and U1753 (N_1753,N_388,N_6);
or U1754 (N_1754,N_421,N_140);
and U1755 (N_1755,N_382,N_887);
nor U1756 (N_1756,N_978,N_290);
and U1757 (N_1757,N_543,N_24);
and U1758 (N_1758,N_255,N_254);
or U1759 (N_1759,N_246,N_30);
nand U1760 (N_1760,N_214,N_530);
or U1761 (N_1761,N_1,N_100);
nand U1762 (N_1762,N_945,N_171);
nor U1763 (N_1763,N_990,N_561);
and U1764 (N_1764,N_154,N_977);
or U1765 (N_1765,N_518,N_379);
nor U1766 (N_1766,N_9,N_258);
nand U1767 (N_1767,N_648,N_858);
nor U1768 (N_1768,N_663,N_730);
nor U1769 (N_1769,N_753,N_737);
or U1770 (N_1770,N_950,N_99);
or U1771 (N_1771,N_806,N_787);
or U1772 (N_1772,N_409,N_381);
and U1773 (N_1773,N_586,N_361);
or U1774 (N_1774,N_771,N_566);
nor U1775 (N_1775,N_444,N_260);
nor U1776 (N_1776,N_240,N_564);
or U1777 (N_1777,N_288,N_998);
nor U1778 (N_1778,N_801,N_169);
or U1779 (N_1779,N_846,N_53);
or U1780 (N_1780,N_594,N_966);
nand U1781 (N_1781,N_944,N_158);
nand U1782 (N_1782,N_495,N_46);
nor U1783 (N_1783,N_385,N_502);
nand U1784 (N_1784,N_330,N_619);
and U1785 (N_1785,N_817,N_124);
or U1786 (N_1786,N_857,N_400);
nand U1787 (N_1787,N_992,N_857);
nand U1788 (N_1788,N_469,N_719);
nand U1789 (N_1789,N_829,N_982);
nor U1790 (N_1790,N_507,N_398);
nor U1791 (N_1791,N_704,N_956);
or U1792 (N_1792,N_699,N_331);
and U1793 (N_1793,N_151,N_767);
nand U1794 (N_1794,N_469,N_255);
nand U1795 (N_1795,N_384,N_133);
nand U1796 (N_1796,N_833,N_228);
or U1797 (N_1797,N_179,N_688);
nor U1798 (N_1798,N_777,N_548);
and U1799 (N_1799,N_735,N_877);
nand U1800 (N_1800,N_36,N_688);
nand U1801 (N_1801,N_208,N_38);
nor U1802 (N_1802,N_865,N_515);
or U1803 (N_1803,N_280,N_523);
and U1804 (N_1804,N_892,N_734);
nand U1805 (N_1805,N_759,N_208);
nor U1806 (N_1806,N_99,N_827);
and U1807 (N_1807,N_71,N_222);
or U1808 (N_1808,N_695,N_237);
and U1809 (N_1809,N_616,N_899);
or U1810 (N_1810,N_259,N_700);
nand U1811 (N_1811,N_359,N_591);
or U1812 (N_1812,N_839,N_840);
nor U1813 (N_1813,N_53,N_487);
nor U1814 (N_1814,N_495,N_657);
nor U1815 (N_1815,N_684,N_935);
nand U1816 (N_1816,N_209,N_355);
nand U1817 (N_1817,N_455,N_909);
nand U1818 (N_1818,N_624,N_102);
or U1819 (N_1819,N_588,N_596);
nor U1820 (N_1820,N_57,N_772);
or U1821 (N_1821,N_903,N_528);
or U1822 (N_1822,N_166,N_332);
nor U1823 (N_1823,N_164,N_676);
nand U1824 (N_1824,N_140,N_25);
and U1825 (N_1825,N_754,N_221);
and U1826 (N_1826,N_555,N_989);
and U1827 (N_1827,N_175,N_568);
and U1828 (N_1828,N_11,N_884);
or U1829 (N_1829,N_735,N_931);
nor U1830 (N_1830,N_255,N_202);
or U1831 (N_1831,N_270,N_65);
or U1832 (N_1832,N_482,N_522);
and U1833 (N_1833,N_549,N_253);
or U1834 (N_1834,N_811,N_896);
or U1835 (N_1835,N_999,N_239);
nor U1836 (N_1836,N_1,N_984);
or U1837 (N_1837,N_96,N_671);
nor U1838 (N_1838,N_327,N_43);
nand U1839 (N_1839,N_662,N_257);
nand U1840 (N_1840,N_608,N_973);
or U1841 (N_1841,N_582,N_635);
and U1842 (N_1842,N_440,N_397);
nand U1843 (N_1843,N_33,N_448);
nor U1844 (N_1844,N_61,N_463);
or U1845 (N_1845,N_936,N_374);
and U1846 (N_1846,N_548,N_814);
nor U1847 (N_1847,N_319,N_981);
and U1848 (N_1848,N_575,N_105);
nand U1849 (N_1849,N_682,N_329);
or U1850 (N_1850,N_789,N_86);
nand U1851 (N_1851,N_775,N_66);
nand U1852 (N_1852,N_365,N_617);
nand U1853 (N_1853,N_111,N_813);
nor U1854 (N_1854,N_202,N_340);
nor U1855 (N_1855,N_397,N_595);
nor U1856 (N_1856,N_898,N_498);
nor U1857 (N_1857,N_331,N_974);
nor U1858 (N_1858,N_173,N_913);
and U1859 (N_1859,N_899,N_940);
and U1860 (N_1860,N_570,N_167);
and U1861 (N_1861,N_531,N_133);
and U1862 (N_1862,N_147,N_605);
and U1863 (N_1863,N_41,N_741);
and U1864 (N_1864,N_177,N_750);
or U1865 (N_1865,N_848,N_797);
nor U1866 (N_1866,N_275,N_790);
and U1867 (N_1867,N_203,N_3);
or U1868 (N_1868,N_50,N_854);
and U1869 (N_1869,N_382,N_268);
nor U1870 (N_1870,N_700,N_752);
nor U1871 (N_1871,N_66,N_772);
and U1872 (N_1872,N_68,N_636);
or U1873 (N_1873,N_791,N_464);
nand U1874 (N_1874,N_905,N_756);
nor U1875 (N_1875,N_323,N_507);
nand U1876 (N_1876,N_571,N_484);
nand U1877 (N_1877,N_141,N_115);
and U1878 (N_1878,N_131,N_465);
nor U1879 (N_1879,N_733,N_236);
and U1880 (N_1880,N_915,N_688);
and U1881 (N_1881,N_0,N_736);
and U1882 (N_1882,N_289,N_81);
nor U1883 (N_1883,N_215,N_493);
nor U1884 (N_1884,N_694,N_726);
xnor U1885 (N_1885,N_169,N_211);
or U1886 (N_1886,N_834,N_777);
or U1887 (N_1887,N_695,N_751);
nor U1888 (N_1888,N_492,N_872);
nand U1889 (N_1889,N_823,N_264);
nand U1890 (N_1890,N_105,N_770);
and U1891 (N_1891,N_828,N_617);
or U1892 (N_1892,N_110,N_550);
and U1893 (N_1893,N_489,N_652);
and U1894 (N_1894,N_385,N_717);
and U1895 (N_1895,N_407,N_165);
nor U1896 (N_1896,N_767,N_438);
nand U1897 (N_1897,N_462,N_879);
nor U1898 (N_1898,N_414,N_632);
nand U1899 (N_1899,N_810,N_334);
or U1900 (N_1900,N_712,N_384);
nor U1901 (N_1901,N_647,N_482);
or U1902 (N_1902,N_328,N_982);
or U1903 (N_1903,N_982,N_479);
nor U1904 (N_1904,N_857,N_282);
nand U1905 (N_1905,N_676,N_567);
nand U1906 (N_1906,N_372,N_993);
nand U1907 (N_1907,N_86,N_515);
or U1908 (N_1908,N_360,N_714);
nor U1909 (N_1909,N_927,N_541);
and U1910 (N_1910,N_643,N_422);
nor U1911 (N_1911,N_511,N_588);
and U1912 (N_1912,N_194,N_276);
nor U1913 (N_1913,N_146,N_728);
nand U1914 (N_1914,N_598,N_895);
nor U1915 (N_1915,N_249,N_700);
nand U1916 (N_1916,N_30,N_989);
and U1917 (N_1917,N_938,N_640);
or U1918 (N_1918,N_268,N_439);
nand U1919 (N_1919,N_92,N_267);
or U1920 (N_1920,N_657,N_429);
and U1921 (N_1921,N_120,N_937);
and U1922 (N_1922,N_146,N_138);
and U1923 (N_1923,N_927,N_585);
or U1924 (N_1924,N_744,N_568);
or U1925 (N_1925,N_540,N_475);
nand U1926 (N_1926,N_662,N_36);
or U1927 (N_1927,N_260,N_853);
and U1928 (N_1928,N_725,N_59);
and U1929 (N_1929,N_767,N_759);
nor U1930 (N_1930,N_552,N_982);
nand U1931 (N_1931,N_439,N_522);
nand U1932 (N_1932,N_528,N_877);
and U1933 (N_1933,N_487,N_368);
nor U1934 (N_1934,N_627,N_814);
or U1935 (N_1935,N_205,N_965);
nor U1936 (N_1936,N_342,N_579);
nand U1937 (N_1937,N_247,N_111);
nor U1938 (N_1938,N_585,N_604);
or U1939 (N_1939,N_42,N_513);
nor U1940 (N_1940,N_380,N_155);
nor U1941 (N_1941,N_182,N_464);
nand U1942 (N_1942,N_592,N_717);
and U1943 (N_1943,N_822,N_176);
or U1944 (N_1944,N_90,N_827);
nand U1945 (N_1945,N_316,N_712);
nor U1946 (N_1946,N_337,N_402);
and U1947 (N_1947,N_993,N_720);
or U1948 (N_1948,N_969,N_23);
and U1949 (N_1949,N_388,N_536);
nor U1950 (N_1950,N_328,N_218);
nand U1951 (N_1951,N_849,N_19);
or U1952 (N_1952,N_201,N_81);
or U1953 (N_1953,N_217,N_804);
or U1954 (N_1954,N_497,N_752);
nand U1955 (N_1955,N_131,N_134);
or U1956 (N_1956,N_586,N_797);
and U1957 (N_1957,N_235,N_46);
and U1958 (N_1958,N_425,N_862);
nand U1959 (N_1959,N_479,N_96);
or U1960 (N_1960,N_175,N_639);
and U1961 (N_1961,N_534,N_946);
or U1962 (N_1962,N_825,N_873);
or U1963 (N_1963,N_99,N_533);
or U1964 (N_1964,N_917,N_834);
nand U1965 (N_1965,N_506,N_949);
nand U1966 (N_1966,N_294,N_864);
nand U1967 (N_1967,N_460,N_149);
nand U1968 (N_1968,N_824,N_266);
and U1969 (N_1969,N_191,N_597);
or U1970 (N_1970,N_943,N_767);
and U1971 (N_1971,N_504,N_971);
and U1972 (N_1972,N_742,N_969);
nand U1973 (N_1973,N_360,N_201);
nand U1974 (N_1974,N_468,N_915);
and U1975 (N_1975,N_620,N_758);
and U1976 (N_1976,N_826,N_41);
and U1977 (N_1977,N_610,N_442);
and U1978 (N_1978,N_520,N_108);
nand U1979 (N_1979,N_154,N_575);
nand U1980 (N_1980,N_172,N_395);
nor U1981 (N_1981,N_335,N_755);
and U1982 (N_1982,N_644,N_850);
or U1983 (N_1983,N_861,N_201);
or U1984 (N_1984,N_170,N_599);
nand U1985 (N_1985,N_353,N_709);
nand U1986 (N_1986,N_689,N_973);
nand U1987 (N_1987,N_723,N_732);
nand U1988 (N_1988,N_406,N_913);
nor U1989 (N_1989,N_818,N_67);
or U1990 (N_1990,N_10,N_971);
nor U1991 (N_1991,N_678,N_256);
and U1992 (N_1992,N_117,N_797);
nand U1993 (N_1993,N_524,N_180);
and U1994 (N_1994,N_800,N_927);
nor U1995 (N_1995,N_728,N_509);
and U1996 (N_1996,N_67,N_373);
or U1997 (N_1997,N_906,N_98);
nor U1998 (N_1998,N_740,N_169);
and U1999 (N_1999,N_535,N_118);
or U2000 (N_2000,N_1036,N_1178);
or U2001 (N_2001,N_1809,N_1918);
nand U2002 (N_2002,N_1974,N_1104);
or U2003 (N_2003,N_1502,N_1777);
and U2004 (N_2004,N_1078,N_1568);
and U2005 (N_2005,N_1721,N_1558);
nor U2006 (N_2006,N_1647,N_1847);
or U2007 (N_2007,N_1322,N_1472);
nor U2008 (N_2008,N_1842,N_1066);
and U2009 (N_2009,N_1469,N_1949);
or U2010 (N_2010,N_1826,N_1642);
or U2011 (N_2011,N_1088,N_1992);
and U2012 (N_2012,N_1661,N_1493);
and U2013 (N_2013,N_1391,N_1863);
or U2014 (N_2014,N_1432,N_1175);
nor U2015 (N_2015,N_1085,N_1486);
or U2016 (N_2016,N_1941,N_1629);
or U2017 (N_2017,N_1789,N_1467);
or U2018 (N_2018,N_1621,N_1287);
nor U2019 (N_2019,N_1099,N_1180);
nand U2020 (N_2020,N_1732,N_1640);
and U2021 (N_2021,N_1892,N_1478);
and U2022 (N_2022,N_1654,N_1044);
nand U2023 (N_2023,N_1998,N_1367);
nor U2024 (N_2024,N_1716,N_1622);
nand U2025 (N_2025,N_1908,N_1083);
and U2026 (N_2026,N_1098,N_1375);
nand U2027 (N_2027,N_1989,N_1094);
nor U2028 (N_2028,N_1805,N_1966);
nor U2029 (N_2029,N_1215,N_1386);
or U2030 (N_2030,N_1578,N_1143);
or U2031 (N_2031,N_1070,N_1501);
and U2032 (N_2032,N_1565,N_1172);
and U2033 (N_2033,N_1906,N_1818);
or U2034 (N_2034,N_1903,N_1672);
nor U2035 (N_2035,N_1026,N_1772);
nor U2036 (N_2036,N_1293,N_1829);
or U2037 (N_2037,N_1579,N_1228);
nor U2038 (N_2038,N_1910,N_1510);
or U2039 (N_2039,N_1631,N_1177);
or U2040 (N_2040,N_1373,N_1990);
nand U2041 (N_2041,N_1313,N_1873);
nor U2042 (N_2042,N_1308,N_1054);
nand U2043 (N_2043,N_1552,N_1162);
nand U2044 (N_2044,N_1820,N_1576);
nand U2045 (N_2045,N_1471,N_1118);
or U2046 (N_2046,N_1267,N_1075);
and U2047 (N_2047,N_1755,N_1024);
or U2048 (N_2048,N_1276,N_1141);
nor U2049 (N_2049,N_1874,N_1484);
or U2050 (N_2050,N_1278,N_1554);
nand U2051 (N_2051,N_1802,N_1042);
nand U2052 (N_2052,N_1255,N_1316);
or U2053 (N_2053,N_1438,N_1244);
nand U2054 (N_2054,N_1403,N_1776);
or U2055 (N_2055,N_1630,N_1972);
nor U2056 (N_2056,N_1766,N_1524);
or U2057 (N_2057,N_1294,N_1334);
nand U2058 (N_2058,N_1182,N_1010);
or U2059 (N_2059,N_1982,N_1871);
and U2060 (N_2060,N_1106,N_1005);
and U2061 (N_2061,N_1535,N_1167);
or U2062 (N_2062,N_1600,N_1900);
nor U2063 (N_2063,N_1979,N_1832);
or U2064 (N_2064,N_1147,N_1796);
or U2065 (N_2065,N_1213,N_1381);
and U2066 (N_2066,N_1342,N_1016);
and U2067 (N_2067,N_1254,N_1679);
or U2068 (N_2068,N_1206,N_1607);
or U2069 (N_2069,N_1555,N_1623);
or U2070 (N_2070,N_1378,N_1030);
or U2071 (N_2071,N_1503,N_1132);
and U2072 (N_2072,N_1529,N_1929);
nand U2073 (N_2073,N_1304,N_1319);
nor U2074 (N_2074,N_1123,N_1664);
or U2075 (N_2075,N_1298,N_1436);
nand U2076 (N_2076,N_1077,N_1318);
nor U2077 (N_2077,N_1814,N_1539);
or U2078 (N_2078,N_1780,N_1186);
or U2079 (N_2079,N_1144,N_1131);
or U2080 (N_2080,N_1053,N_1179);
nand U2081 (N_2081,N_1210,N_1650);
nor U2082 (N_2082,N_1142,N_1007);
and U2083 (N_2083,N_1008,N_1023);
nand U2084 (N_2084,N_1928,N_1091);
nand U2085 (N_2085,N_1233,N_1598);
and U2086 (N_2086,N_1051,N_1810);
and U2087 (N_2087,N_1111,N_1546);
or U2088 (N_2088,N_1522,N_1133);
or U2089 (N_2089,N_1136,N_1082);
or U2090 (N_2090,N_1626,N_1317);
or U2091 (N_2091,N_1747,N_1382);
nor U2092 (N_2092,N_1680,N_1314);
or U2093 (N_2093,N_1272,N_1663);
nor U2094 (N_2094,N_1997,N_1656);
or U2095 (N_2095,N_1341,N_1139);
nand U2096 (N_2096,N_1209,N_1056);
or U2097 (N_2097,N_1473,N_1475);
and U2098 (N_2098,N_1790,N_1920);
nand U2099 (N_2099,N_1572,N_1935);
or U2100 (N_2100,N_1303,N_1859);
nor U2101 (N_2101,N_1084,N_1216);
or U2102 (N_2102,N_1618,N_1913);
and U2103 (N_2103,N_1039,N_1156);
or U2104 (N_2104,N_1909,N_1839);
nand U2105 (N_2105,N_1715,N_1669);
nand U2106 (N_2106,N_1069,N_1547);
nand U2107 (N_2107,N_1414,N_1065);
or U2108 (N_2108,N_1490,N_1823);
nand U2109 (N_2109,N_1052,N_1761);
or U2110 (N_2110,N_1916,N_1114);
nor U2111 (N_2111,N_1466,N_1037);
nand U2112 (N_2112,N_1852,N_1975);
and U2113 (N_2113,N_1794,N_1028);
and U2114 (N_2114,N_1251,N_1521);
nor U2115 (N_2115,N_1924,N_1987);
nand U2116 (N_2116,N_1290,N_1076);
or U2117 (N_2117,N_1333,N_1343);
nand U2118 (N_2118,N_1337,N_1212);
xnor U2119 (N_2119,N_1281,N_1574);
nor U2120 (N_2120,N_1923,N_1459);
nand U2121 (N_2121,N_1161,N_1116);
nor U2122 (N_2122,N_1635,N_1006);
nand U2123 (N_2123,N_1160,N_1691);
and U2124 (N_2124,N_1628,N_1737);
nand U2125 (N_2125,N_1087,N_1634);
or U2126 (N_2126,N_1100,N_1043);
nand U2127 (N_2127,N_1557,N_1017);
or U2128 (N_2128,N_1881,N_1494);
nand U2129 (N_2129,N_1135,N_1690);
or U2130 (N_2130,N_1932,N_1401);
nand U2131 (N_2131,N_1697,N_1020);
and U2132 (N_2132,N_1451,N_1921);
or U2133 (N_2133,N_1841,N_1659);
nor U2134 (N_2134,N_1402,N_1000);
nor U2135 (N_2135,N_1709,N_1108);
nand U2136 (N_2136,N_1678,N_1811);
nor U2137 (N_2137,N_1528,N_1687);
nand U2138 (N_2138,N_1785,N_1442);
or U2139 (N_2139,N_1046,N_1041);
nand U2140 (N_2140,N_1433,N_1309);
and U2141 (N_2141,N_1201,N_1090);
nand U2142 (N_2142,N_1384,N_1682);
and U2143 (N_2143,N_1954,N_1035);
or U2144 (N_2144,N_1925,N_1788);
or U2145 (N_2145,N_1627,N_1221);
or U2146 (N_2146,N_1795,N_1335);
and U2147 (N_2147,N_1936,N_1413);
and U2148 (N_2148,N_1173,N_1371);
nand U2149 (N_2149,N_1651,N_1567);
nand U2150 (N_2150,N_1944,N_1828);
nor U2151 (N_2151,N_1880,N_1739);
and U2152 (N_2152,N_1243,N_1980);
or U2153 (N_2153,N_1886,N_1032);
and U2154 (N_2154,N_1348,N_1988);
and U2155 (N_2155,N_1655,N_1191);
and U2156 (N_2156,N_1877,N_1109);
and U2157 (N_2157,N_1025,N_1349);
or U2158 (N_2158,N_1418,N_1813);
or U2159 (N_2159,N_1347,N_1279);
and U2160 (N_2160,N_1843,N_1235);
nand U2161 (N_2161,N_1389,N_1962);
nand U2162 (N_2162,N_1211,N_1038);
or U2163 (N_2163,N_1756,N_1400);
nand U2164 (N_2164,N_1550,N_1538);
nand U2165 (N_2165,N_1107,N_1733);
and U2166 (N_2166,N_1580,N_1245);
nand U2167 (N_2167,N_1985,N_1014);
or U2168 (N_2168,N_1029,N_1745);
and U2169 (N_2169,N_1345,N_1280);
nand U2170 (N_2170,N_1291,N_1080);
nor U2171 (N_2171,N_1945,N_1508);
nand U2172 (N_2172,N_1189,N_1658);
nor U2173 (N_2173,N_1002,N_1942);
or U2174 (N_2174,N_1410,N_1986);
xor U2175 (N_2175,N_1190,N_1560);
nand U2176 (N_2176,N_1882,N_1089);
nand U2177 (N_2177,N_1284,N_1458);
or U2178 (N_2178,N_1649,N_1968);
nand U2179 (N_2179,N_1417,N_1463);
and U2180 (N_2180,N_1012,N_1454);
or U2181 (N_2181,N_1549,N_1018);
nor U2182 (N_2182,N_1232,N_1031);
nand U2183 (N_2183,N_1613,N_1507);
or U2184 (N_2184,N_1612,N_1950);
and U2185 (N_2185,N_1984,N_1079);
nor U2186 (N_2186,N_1896,N_1778);
nand U2187 (N_2187,N_1500,N_1205);
and U2188 (N_2188,N_1581,N_1851);
and U2189 (N_2189,N_1525,N_1520);
nand U2190 (N_2190,N_1127,N_1264);
or U2191 (N_2191,N_1257,N_1444);
and U2192 (N_2192,N_1328,N_1887);
or U2193 (N_2193,N_1351,N_1657);
and U2194 (N_2194,N_1352,N_1259);
and U2195 (N_2195,N_1450,N_1515);
and U2196 (N_2196,N_1406,N_1196);
nand U2197 (N_2197,N_1773,N_1312);
xnor U2198 (N_2198,N_1676,N_1670);
or U2199 (N_2199,N_1853,N_1121);
nand U2200 (N_2200,N_1258,N_1643);
or U2201 (N_2201,N_1140,N_1226);
nor U2202 (N_2202,N_1262,N_1261);
or U2203 (N_2203,N_1237,N_1804);
or U2204 (N_2204,N_1854,N_1462);
xnor U2205 (N_2205,N_1838,N_1285);
xnor U2206 (N_2206,N_1126,N_1542);
nor U2207 (N_2207,N_1736,N_1128);
nand U2208 (N_2208,N_1155,N_1566);
or U2209 (N_2209,N_1693,N_1457);
and U2210 (N_2210,N_1145,N_1927);
nor U2211 (N_2211,N_1953,N_1222);
or U2212 (N_2212,N_1274,N_1383);
or U2213 (N_2213,N_1427,N_1531);
or U2214 (N_2214,N_1797,N_1963);
and U2215 (N_2215,N_1122,N_1995);
and U2216 (N_2216,N_1397,N_1708);
and U2217 (N_2217,N_1071,N_1166);
nand U2218 (N_2218,N_1591,N_1398);
nand U2219 (N_2219,N_1372,N_1058);
nor U2220 (N_2220,N_1188,N_1482);
nor U2221 (N_2221,N_1376,N_1359);
nand U2222 (N_2222,N_1798,N_1978);
or U2223 (N_2223,N_1907,N_1860);
and U2224 (N_2224,N_1835,N_1964);
nor U2225 (N_2225,N_1117,N_1488);
or U2226 (N_2226,N_1719,N_1068);
or U2227 (N_2227,N_1353,N_1545);
nor U2228 (N_2228,N_1636,N_1884);
and U2229 (N_2229,N_1686,N_1605);
nor U2230 (N_2230,N_1575,N_1774);
and U2231 (N_2231,N_1699,N_1369);
and U2232 (N_2232,N_1153,N_1004);
or U2233 (N_2233,N_1445,N_1492);
nor U2234 (N_2234,N_1677,N_1022);
or U2235 (N_2235,N_1050,N_1229);
or U2236 (N_2236,N_1412,N_1668);
and U2237 (N_2237,N_1991,N_1409);
nand U2238 (N_2238,N_1385,N_1878);
xor U2239 (N_2239,N_1356,N_1564);
nand U2240 (N_2240,N_1405,N_1247);
and U2241 (N_2241,N_1711,N_1019);
and U2242 (N_2242,N_1955,N_1277);
or U2243 (N_2243,N_1416,N_1781);
and U2244 (N_2244,N_1562,N_1606);
nor U2245 (N_2245,N_1969,N_1919);
and U2246 (N_2246,N_1425,N_1812);
nand U2247 (N_2247,N_1762,N_1758);
or U2248 (N_2248,N_1207,N_1465);
or U2249 (N_2249,N_1750,N_1112);
nor U2250 (N_2250,N_1270,N_1738);
or U2251 (N_2251,N_1366,N_1374);
or U2252 (N_2252,N_1653,N_1148);
xnor U2253 (N_2253,N_1495,N_1393);
and U2254 (N_2254,N_1705,N_1748);
or U2255 (N_2255,N_1480,N_1346);
nand U2256 (N_2256,N_1396,N_1571);
nor U2257 (N_2257,N_1115,N_1086);
nand U2258 (N_2258,N_1577,N_1675);
nand U2259 (N_2259,N_1729,N_1742);
and U2260 (N_2260,N_1849,N_1931);
nand U2261 (N_2261,N_1725,N_1722);
nand U2262 (N_2262,N_1844,N_1633);
and U2263 (N_2263,N_1741,N_1430);
or U2264 (N_2264,N_1517,N_1526);
nor U2265 (N_2265,N_1751,N_1946);
or U2266 (N_2266,N_1559,N_1198);
nand U2267 (N_2267,N_1074,N_1596);
and U2268 (N_2268,N_1326,N_1787);
or U2269 (N_2269,N_1671,N_1227);
nor U2270 (N_2270,N_1464,N_1889);
nor U2271 (N_2271,N_1461,N_1983);
nor U2272 (N_2272,N_1867,N_1271);
nand U2273 (N_2273,N_1893,N_1283);
nand U2274 (N_2274,N_1723,N_1063);
nand U2275 (N_2275,N_1040,N_1302);
nor U2276 (N_2276,N_1771,N_1740);
and U2277 (N_2277,N_1336,N_1169);
or U2278 (N_2278,N_1256,N_1960);
nand U2279 (N_2279,N_1370,N_1420);
nor U2280 (N_2280,N_1350,N_1263);
and U2281 (N_2281,N_1994,N_1674);
or U2282 (N_2282,N_1840,N_1563);
or U2283 (N_2283,N_1157,N_1735);
nor U2284 (N_2284,N_1976,N_1435);
nor U2285 (N_2285,N_1866,N_1176);
nor U2286 (N_2286,N_1377,N_1292);
or U2287 (N_2287,N_1648,N_1363);
nand U2288 (N_2288,N_1223,N_1752);
and U2289 (N_2289,N_1193,N_1553);
or U2290 (N_2290,N_1119,N_1214);
nor U2291 (N_2291,N_1236,N_1712);
nand U2292 (N_2292,N_1573,N_1231);
nand U2293 (N_2293,N_1718,N_1163);
or U2294 (N_2294,N_1540,N_1816);
or U2295 (N_2295,N_1685,N_1704);
and U2296 (N_2296,N_1249,N_1183);
or U2297 (N_2297,N_1230,N_1300);
and U2298 (N_2298,N_1834,N_1394);
nand U2299 (N_2299,N_1034,N_1124);
or U2300 (N_2300,N_1617,N_1282);
or U2301 (N_2301,N_1746,N_1057);
nor U2302 (N_2302,N_1202,N_1504);
nand U2303 (N_2303,N_1831,N_1491);
and U2304 (N_2304,N_1999,N_1977);
or U2305 (N_2305,N_1523,N_1786);
nand U2306 (N_2306,N_1888,N_1996);
and U2307 (N_2307,N_1822,N_1513);
or U2308 (N_2308,N_1305,N_1073);
nor U2309 (N_2309,N_1731,N_1958);
nand U2310 (N_2310,N_1897,N_1130);
or U2311 (N_2311,N_1551,N_1062);
nor U2312 (N_2312,N_1602,N_1593);
nand U2313 (N_2313,N_1364,N_1092);
and U2314 (N_2314,N_1971,N_1701);
nand U2315 (N_2315,N_1242,N_1361);
and U2316 (N_2316,N_1240,N_1011);
or U2317 (N_2317,N_1399,N_1695);
or U2318 (N_2318,N_1876,N_1447);
and U2319 (N_2319,N_1608,N_1692);
or U2320 (N_2320,N_1534,N_1476);
nor U2321 (N_2321,N_1422,N_1224);
nor U2322 (N_2322,N_1779,N_1943);
or U2323 (N_2323,N_1743,N_1597);
nand U2324 (N_2324,N_1097,N_1898);
nand U2325 (N_2325,N_1033,N_1516);
and U2326 (N_2326,N_1047,N_1846);
nor U2327 (N_2327,N_1159,N_1379);
nand U2328 (N_2328,N_1453,N_1836);
nand U2329 (N_2329,N_1710,N_1358);
nor U2330 (N_2330,N_1429,N_1940);
and U2331 (N_2331,N_1061,N_1939);
and U2332 (N_2332,N_1269,N_1603);
nand U2333 (N_2333,N_1174,N_1864);
or U2334 (N_2334,N_1775,N_1434);
nor U2335 (N_2335,N_1489,N_1171);
or U2336 (N_2336,N_1275,N_1067);
or U2337 (N_2337,N_1757,N_1714);
nand U2338 (N_2338,N_1120,N_1194);
xor U2339 (N_2339,N_1611,N_1800);
and U2340 (N_2340,N_1614,N_1101);
or U2341 (N_2341,N_1129,N_1059);
nor U2342 (N_2342,N_1696,N_1641);
or U2343 (N_2343,N_1544,N_1933);
or U2344 (N_2344,N_1509,N_1934);
and U2345 (N_2345,N_1753,N_1754);
or U2346 (N_2346,N_1681,N_1744);
or U2347 (N_2347,N_1717,N_1537);
nor U2348 (N_2348,N_1325,N_1625);
nor U2349 (N_2349,N_1519,N_1357);
nor U2350 (N_2350,N_1703,N_1217);
nand U2351 (N_2351,N_1477,N_1437);
and U2352 (N_2352,N_1764,N_1360);
nor U2353 (N_2353,N_1021,N_1220);
nand U2354 (N_2354,N_1408,N_1499);
and U2355 (N_2355,N_1260,N_1168);
nor U2356 (N_2356,N_1288,N_1297);
nand U2357 (N_2357,N_1295,N_1922);
or U2358 (N_2358,N_1895,N_1095);
nand U2359 (N_2359,N_1252,N_1904);
nand U2360 (N_2360,N_1981,N_1856);
nor U2361 (N_2361,N_1827,N_1355);
or U2362 (N_2362,N_1837,N_1362);
or U2363 (N_2363,N_1421,N_1765);
nand U2364 (N_2364,N_1915,N_1824);
or U2365 (N_2365,N_1137,N_1792);
or U2366 (N_2366,N_1582,N_1961);
or U2367 (N_2367,N_1730,N_1380);
nand U2368 (N_2368,N_1248,N_1203);
and U2369 (N_2369,N_1165,N_1947);
nor U2370 (N_2370,N_1110,N_1446);
and U2371 (N_2371,N_1072,N_1340);
or U2372 (N_2372,N_1511,N_1861);
and U2373 (N_2373,N_1185,N_1957);
nand U2374 (N_2374,N_1392,N_1428);
or U2375 (N_2375,N_1624,N_1590);
nor U2376 (N_2376,N_1973,N_1150);
and U2377 (N_2377,N_1956,N_1315);
nor U2378 (N_2378,N_1587,N_1720);
or U2379 (N_2379,N_1784,N_1533);
nor U2380 (N_2380,N_1665,N_1266);
or U2381 (N_2381,N_1234,N_1530);
or U2382 (N_2382,N_1917,N_1894);
or U2383 (N_2383,N_1105,N_1803);
and U2384 (N_2384,N_1184,N_1684);
nor U2385 (N_2385,N_1113,N_1485);
nand U2386 (N_2386,N_1411,N_1707);
nand U2387 (N_2387,N_1639,N_1138);
and U2388 (N_2388,N_1645,N_1799);
and U2389 (N_2389,N_1419,N_1937);
or U2390 (N_2390,N_1324,N_1899);
nand U2391 (N_2391,N_1299,N_1456);
or U2392 (N_2392,N_1855,N_1702);
nand U2393 (N_2393,N_1660,N_1620);
nor U2394 (N_2394,N_1594,N_1768);
and U2395 (N_2395,N_1646,N_1505);
nor U2396 (N_2396,N_1149,N_1219);
or U2397 (N_2397,N_1239,N_1468);
nor U2398 (N_2398,N_1783,N_1870);
nor U2399 (N_2399,N_1158,N_1698);
and U2400 (N_2400,N_1265,N_1204);
nand U2401 (N_2401,N_1331,N_1200);
or U2402 (N_2402,N_1439,N_1246);
or U2403 (N_2403,N_1589,N_1819);
or U2404 (N_2404,N_1914,N_1443);
and U2405 (N_2405,N_1912,N_1632);
and U2406 (N_2406,N_1015,N_1993);
xnor U2407 (N_2407,N_1387,N_1474);
and U2408 (N_2408,N_1483,N_1588);
nor U2409 (N_2409,N_1902,N_1518);
or U2410 (N_2410,N_1817,N_1009);
nand U2411 (N_2411,N_1638,N_1713);
nand U2412 (N_2412,N_1688,N_1806);
and U2413 (N_2413,N_1673,N_1096);
nor U2414 (N_2414,N_1125,N_1782);
nand U2415 (N_2415,N_1296,N_1487);
and U2416 (N_2416,N_1850,N_1448);
nor U2417 (N_2417,N_1930,N_1481);
and U2418 (N_2418,N_1890,N_1891);
or U2419 (N_2419,N_1354,N_1760);
nor U2420 (N_2420,N_1289,N_1506);
and U2421 (N_2421,N_1332,N_1875);
or U2422 (N_2422,N_1667,N_1767);
nand U2423 (N_2423,N_1543,N_1585);
and U2424 (N_2424,N_1306,N_1848);
nand U2425 (N_2425,N_1694,N_1479);
or U2426 (N_2426,N_1218,N_1965);
or U2427 (N_2427,N_1423,N_1601);
nand U2428 (N_2428,N_1791,N_1883);
nand U2429 (N_2429,N_1911,N_1441);
nand U2430 (N_2430,N_1662,N_1339);
nor U2431 (N_2431,N_1583,N_1151);
xnor U2432 (N_2432,N_1734,N_1407);
or U2433 (N_2433,N_1959,N_1307);
and U2434 (N_2434,N_1683,N_1644);
and U2435 (N_2435,N_1013,N_1365);
nand U2436 (N_2436,N_1310,N_1498);
or U2437 (N_2437,N_1865,N_1970);
nand U2438 (N_2438,N_1609,N_1905);
and U2439 (N_2439,N_1208,N_1967);
nand U2440 (N_2440,N_1793,N_1388);
or U2441 (N_2441,N_1081,N_1586);
nand U2442 (N_2442,N_1045,N_1514);
nor U2443 (N_2443,N_1241,N_1512);
nor U2444 (N_2444,N_1368,N_1869);
or U2445 (N_2445,N_1181,N_1556);
nor U2446 (N_2446,N_1460,N_1253);
nand U2447 (N_2447,N_1170,N_1862);
and U2448 (N_2448,N_1327,N_1395);
or U2449 (N_2449,N_1595,N_1727);
or U2450 (N_2450,N_1301,N_1536);
or U2451 (N_2451,N_1724,N_1329);
nand U2452 (N_2452,N_1821,N_1225);
nand U2453 (N_2453,N_1615,N_1952);
and U2454 (N_2454,N_1868,N_1570);
nand U2455 (N_2455,N_1637,N_1759);
or U2456 (N_2456,N_1415,N_1561);
nor U2457 (N_2457,N_1706,N_1093);
nand U2458 (N_2458,N_1003,N_1470);
and U2459 (N_2459,N_1102,N_1830);
nor U2460 (N_2460,N_1807,N_1569);
nor U2461 (N_2461,N_1103,N_1584);
nand U2462 (N_2462,N_1619,N_1192);
or U2463 (N_2463,N_1592,N_1187);
and U2464 (N_2464,N_1154,N_1048);
nand U2465 (N_2465,N_1749,N_1055);
nand U2466 (N_2466,N_1195,N_1845);
and U2467 (N_2467,N_1728,N_1548);
nand U2468 (N_2468,N_1321,N_1311);
nor U2469 (N_2469,N_1951,N_1700);
and U2470 (N_2470,N_1616,N_1857);
and U2471 (N_2471,N_1527,N_1763);
nor U2472 (N_2472,N_1390,N_1027);
or U2473 (N_2473,N_1452,N_1250);
nor U2474 (N_2474,N_1440,N_1152);
and U2475 (N_2475,N_1858,N_1885);
or U2476 (N_2476,N_1060,N_1268);
nor U2477 (N_2477,N_1197,N_1404);
nor U2478 (N_2478,N_1431,N_1901);
nor U2479 (N_2479,N_1164,N_1726);
and U2480 (N_2480,N_1146,N_1599);
nor U2481 (N_2481,N_1833,N_1338);
and U2482 (N_2482,N_1879,N_1199);
nand U2483 (N_2483,N_1689,N_1825);
nor U2484 (N_2484,N_1496,N_1049);
and U2485 (N_2485,N_1344,N_1666);
nand U2486 (N_2486,N_1426,N_1808);
nor U2487 (N_2487,N_1801,N_1948);
and U2488 (N_2488,N_1815,N_1320);
nand U2489 (N_2489,N_1424,N_1449);
or U2490 (N_2490,N_1323,N_1532);
and U2491 (N_2491,N_1238,N_1770);
nor U2492 (N_2492,N_1610,N_1330);
nor U2493 (N_2493,N_1134,N_1497);
or U2494 (N_2494,N_1064,N_1286);
nor U2495 (N_2495,N_1926,N_1604);
and U2496 (N_2496,N_1455,N_1273);
or U2497 (N_2497,N_1872,N_1001);
and U2498 (N_2498,N_1652,N_1541);
or U2499 (N_2499,N_1938,N_1769);
or U2500 (N_2500,N_1785,N_1359);
nor U2501 (N_2501,N_1342,N_1754);
nor U2502 (N_2502,N_1185,N_1815);
nand U2503 (N_2503,N_1928,N_1053);
nor U2504 (N_2504,N_1532,N_1618);
and U2505 (N_2505,N_1445,N_1221);
nor U2506 (N_2506,N_1258,N_1946);
nor U2507 (N_2507,N_1108,N_1648);
and U2508 (N_2508,N_1654,N_1464);
and U2509 (N_2509,N_1395,N_1907);
nand U2510 (N_2510,N_1365,N_1800);
and U2511 (N_2511,N_1623,N_1126);
and U2512 (N_2512,N_1755,N_1304);
nand U2513 (N_2513,N_1587,N_1570);
and U2514 (N_2514,N_1760,N_1843);
nand U2515 (N_2515,N_1062,N_1549);
and U2516 (N_2516,N_1933,N_1277);
or U2517 (N_2517,N_1990,N_1191);
and U2518 (N_2518,N_1894,N_1744);
nand U2519 (N_2519,N_1917,N_1218);
or U2520 (N_2520,N_1369,N_1217);
xnor U2521 (N_2521,N_1839,N_1836);
nand U2522 (N_2522,N_1253,N_1719);
or U2523 (N_2523,N_1062,N_1766);
xor U2524 (N_2524,N_1593,N_1919);
nor U2525 (N_2525,N_1538,N_1183);
nor U2526 (N_2526,N_1519,N_1597);
or U2527 (N_2527,N_1899,N_1405);
nor U2528 (N_2528,N_1091,N_1816);
and U2529 (N_2529,N_1674,N_1502);
or U2530 (N_2530,N_1711,N_1322);
or U2531 (N_2531,N_1369,N_1085);
or U2532 (N_2532,N_1173,N_1157);
nand U2533 (N_2533,N_1946,N_1208);
nor U2534 (N_2534,N_1439,N_1849);
or U2535 (N_2535,N_1821,N_1696);
or U2536 (N_2536,N_1553,N_1317);
or U2537 (N_2537,N_1837,N_1485);
or U2538 (N_2538,N_1645,N_1455);
or U2539 (N_2539,N_1974,N_1487);
nor U2540 (N_2540,N_1122,N_1818);
or U2541 (N_2541,N_1124,N_1515);
nor U2542 (N_2542,N_1639,N_1611);
and U2543 (N_2543,N_1727,N_1580);
nor U2544 (N_2544,N_1347,N_1531);
and U2545 (N_2545,N_1432,N_1522);
or U2546 (N_2546,N_1536,N_1408);
or U2547 (N_2547,N_1346,N_1284);
and U2548 (N_2548,N_1546,N_1962);
or U2549 (N_2549,N_1560,N_1725);
nor U2550 (N_2550,N_1940,N_1387);
or U2551 (N_2551,N_1511,N_1964);
and U2552 (N_2552,N_1833,N_1699);
and U2553 (N_2553,N_1127,N_1727);
and U2554 (N_2554,N_1728,N_1136);
or U2555 (N_2555,N_1279,N_1277);
nor U2556 (N_2556,N_1683,N_1878);
nor U2557 (N_2557,N_1144,N_1964);
and U2558 (N_2558,N_1847,N_1565);
nor U2559 (N_2559,N_1199,N_1374);
nand U2560 (N_2560,N_1766,N_1063);
nor U2561 (N_2561,N_1786,N_1057);
nor U2562 (N_2562,N_1598,N_1398);
or U2563 (N_2563,N_1243,N_1572);
and U2564 (N_2564,N_1878,N_1028);
and U2565 (N_2565,N_1069,N_1161);
and U2566 (N_2566,N_1552,N_1987);
nor U2567 (N_2567,N_1833,N_1452);
nor U2568 (N_2568,N_1769,N_1054);
or U2569 (N_2569,N_1263,N_1782);
nor U2570 (N_2570,N_1803,N_1931);
or U2571 (N_2571,N_1422,N_1984);
and U2572 (N_2572,N_1958,N_1009);
and U2573 (N_2573,N_1479,N_1275);
nand U2574 (N_2574,N_1948,N_1723);
or U2575 (N_2575,N_1400,N_1655);
nand U2576 (N_2576,N_1300,N_1935);
and U2577 (N_2577,N_1188,N_1984);
nand U2578 (N_2578,N_1477,N_1349);
nor U2579 (N_2579,N_1414,N_1913);
nor U2580 (N_2580,N_1733,N_1330);
nand U2581 (N_2581,N_1900,N_1722);
or U2582 (N_2582,N_1868,N_1804);
nor U2583 (N_2583,N_1890,N_1044);
nor U2584 (N_2584,N_1557,N_1289);
nor U2585 (N_2585,N_1519,N_1023);
and U2586 (N_2586,N_1794,N_1929);
nand U2587 (N_2587,N_1284,N_1725);
nand U2588 (N_2588,N_1097,N_1909);
and U2589 (N_2589,N_1816,N_1513);
nor U2590 (N_2590,N_1539,N_1476);
nor U2591 (N_2591,N_1265,N_1678);
or U2592 (N_2592,N_1774,N_1101);
and U2593 (N_2593,N_1207,N_1131);
nand U2594 (N_2594,N_1261,N_1828);
nor U2595 (N_2595,N_1590,N_1168);
nand U2596 (N_2596,N_1257,N_1966);
and U2597 (N_2597,N_1569,N_1657);
and U2598 (N_2598,N_1930,N_1432);
and U2599 (N_2599,N_1874,N_1470);
nand U2600 (N_2600,N_1539,N_1374);
nand U2601 (N_2601,N_1847,N_1507);
or U2602 (N_2602,N_1168,N_1475);
or U2603 (N_2603,N_1944,N_1491);
and U2604 (N_2604,N_1665,N_1752);
nor U2605 (N_2605,N_1400,N_1601);
nand U2606 (N_2606,N_1131,N_1317);
and U2607 (N_2607,N_1969,N_1459);
and U2608 (N_2608,N_1089,N_1205);
or U2609 (N_2609,N_1020,N_1909);
or U2610 (N_2610,N_1289,N_1797);
or U2611 (N_2611,N_1159,N_1347);
and U2612 (N_2612,N_1262,N_1480);
nor U2613 (N_2613,N_1146,N_1502);
or U2614 (N_2614,N_1534,N_1624);
and U2615 (N_2615,N_1234,N_1424);
nor U2616 (N_2616,N_1894,N_1506);
nor U2617 (N_2617,N_1261,N_1223);
nor U2618 (N_2618,N_1782,N_1535);
nand U2619 (N_2619,N_1029,N_1918);
nand U2620 (N_2620,N_1916,N_1854);
nand U2621 (N_2621,N_1639,N_1600);
or U2622 (N_2622,N_1826,N_1293);
nor U2623 (N_2623,N_1341,N_1422);
and U2624 (N_2624,N_1194,N_1404);
or U2625 (N_2625,N_1085,N_1435);
and U2626 (N_2626,N_1477,N_1744);
nand U2627 (N_2627,N_1790,N_1587);
nor U2628 (N_2628,N_1185,N_1159);
nand U2629 (N_2629,N_1299,N_1287);
nand U2630 (N_2630,N_1458,N_1751);
nor U2631 (N_2631,N_1930,N_1653);
nor U2632 (N_2632,N_1106,N_1349);
or U2633 (N_2633,N_1771,N_1989);
nor U2634 (N_2634,N_1809,N_1076);
nand U2635 (N_2635,N_1778,N_1082);
nand U2636 (N_2636,N_1733,N_1765);
nor U2637 (N_2637,N_1694,N_1090);
nand U2638 (N_2638,N_1627,N_1102);
nand U2639 (N_2639,N_1646,N_1794);
or U2640 (N_2640,N_1389,N_1488);
and U2641 (N_2641,N_1671,N_1530);
nor U2642 (N_2642,N_1821,N_1173);
and U2643 (N_2643,N_1624,N_1368);
and U2644 (N_2644,N_1008,N_1934);
nand U2645 (N_2645,N_1964,N_1669);
nand U2646 (N_2646,N_1436,N_1562);
and U2647 (N_2647,N_1502,N_1258);
nand U2648 (N_2648,N_1673,N_1105);
nor U2649 (N_2649,N_1949,N_1550);
or U2650 (N_2650,N_1943,N_1399);
and U2651 (N_2651,N_1208,N_1765);
and U2652 (N_2652,N_1973,N_1923);
and U2653 (N_2653,N_1711,N_1609);
and U2654 (N_2654,N_1579,N_1004);
nand U2655 (N_2655,N_1326,N_1477);
nand U2656 (N_2656,N_1024,N_1794);
nor U2657 (N_2657,N_1097,N_1537);
nand U2658 (N_2658,N_1190,N_1369);
nand U2659 (N_2659,N_1547,N_1545);
and U2660 (N_2660,N_1276,N_1517);
or U2661 (N_2661,N_1169,N_1673);
nor U2662 (N_2662,N_1219,N_1506);
nand U2663 (N_2663,N_1567,N_1038);
and U2664 (N_2664,N_1988,N_1243);
nand U2665 (N_2665,N_1821,N_1358);
nor U2666 (N_2666,N_1279,N_1797);
and U2667 (N_2667,N_1403,N_1629);
nand U2668 (N_2668,N_1781,N_1029);
nand U2669 (N_2669,N_1738,N_1901);
nor U2670 (N_2670,N_1228,N_1657);
or U2671 (N_2671,N_1671,N_1852);
and U2672 (N_2672,N_1792,N_1942);
or U2673 (N_2673,N_1573,N_1748);
nand U2674 (N_2674,N_1359,N_1148);
nor U2675 (N_2675,N_1578,N_1588);
or U2676 (N_2676,N_1410,N_1382);
nand U2677 (N_2677,N_1700,N_1983);
or U2678 (N_2678,N_1906,N_1090);
nand U2679 (N_2679,N_1942,N_1278);
nand U2680 (N_2680,N_1290,N_1654);
or U2681 (N_2681,N_1172,N_1888);
nand U2682 (N_2682,N_1549,N_1577);
nand U2683 (N_2683,N_1159,N_1953);
nor U2684 (N_2684,N_1370,N_1148);
and U2685 (N_2685,N_1464,N_1992);
nand U2686 (N_2686,N_1483,N_1514);
or U2687 (N_2687,N_1105,N_1552);
and U2688 (N_2688,N_1264,N_1648);
and U2689 (N_2689,N_1536,N_1225);
or U2690 (N_2690,N_1033,N_1780);
nand U2691 (N_2691,N_1743,N_1599);
and U2692 (N_2692,N_1867,N_1788);
nor U2693 (N_2693,N_1329,N_1941);
and U2694 (N_2694,N_1125,N_1766);
nand U2695 (N_2695,N_1637,N_1670);
and U2696 (N_2696,N_1710,N_1446);
nand U2697 (N_2697,N_1881,N_1087);
nor U2698 (N_2698,N_1976,N_1150);
nor U2699 (N_2699,N_1201,N_1907);
nand U2700 (N_2700,N_1356,N_1355);
nor U2701 (N_2701,N_1037,N_1304);
nor U2702 (N_2702,N_1015,N_1595);
nor U2703 (N_2703,N_1809,N_1929);
and U2704 (N_2704,N_1798,N_1572);
and U2705 (N_2705,N_1935,N_1476);
or U2706 (N_2706,N_1000,N_1931);
and U2707 (N_2707,N_1987,N_1284);
and U2708 (N_2708,N_1122,N_1342);
nand U2709 (N_2709,N_1390,N_1264);
and U2710 (N_2710,N_1090,N_1946);
or U2711 (N_2711,N_1924,N_1240);
nand U2712 (N_2712,N_1744,N_1276);
or U2713 (N_2713,N_1560,N_1143);
nand U2714 (N_2714,N_1479,N_1581);
nor U2715 (N_2715,N_1854,N_1117);
or U2716 (N_2716,N_1401,N_1792);
and U2717 (N_2717,N_1825,N_1739);
nand U2718 (N_2718,N_1528,N_1375);
nand U2719 (N_2719,N_1594,N_1022);
nor U2720 (N_2720,N_1797,N_1873);
or U2721 (N_2721,N_1962,N_1137);
nor U2722 (N_2722,N_1615,N_1755);
nor U2723 (N_2723,N_1848,N_1709);
nor U2724 (N_2724,N_1460,N_1792);
nand U2725 (N_2725,N_1514,N_1017);
or U2726 (N_2726,N_1910,N_1014);
or U2727 (N_2727,N_1387,N_1717);
nor U2728 (N_2728,N_1367,N_1206);
or U2729 (N_2729,N_1819,N_1146);
and U2730 (N_2730,N_1448,N_1609);
nor U2731 (N_2731,N_1297,N_1038);
nor U2732 (N_2732,N_1702,N_1707);
and U2733 (N_2733,N_1367,N_1056);
and U2734 (N_2734,N_1666,N_1086);
nor U2735 (N_2735,N_1587,N_1855);
nor U2736 (N_2736,N_1360,N_1164);
and U2737 (N_2737,N_1874,N_1343);
and U2738 (N_2738,N_1993,N_1343);
nand U2739 (N_2739,N_1508,N_1196);
nor U2740 (N_2740,N_1287,N_1916);
or U2741 (N_2741,N_1669,N_1157);
or U2742 (N_2742,N_1065,N_1217);
nand U2743 (N_2743,N_1378,N_1359);
xor U2744 (N_2744,N_1599,N_1594);
and U2745 (N_2745,N_1551,N_1796);
nor U2746 (N_2746,N_1107,N_1257);
or U2747 (N_2747,N_1415,N_1203);
or U2748 (N_2748,N_1105,N_1490);
and U2749 (N_2749,N_1051,N_1703);
nand U2750 (N_2750,N_1102,N_1482);
or U2751 (N_2751,N_1602,N_1586);
and U2752 (N_2752,N_1190,N_1833);
and U2753 (N_2753,N_1800,N_1770);
or U2754 (N_2754,N_1961,N_1949);
or U2755 (N_2755,N_1591,N_1081);
nor U2756 (N_2756,N_1655,N_1612);
nor U2757 (N_2757,N_1156,N_1613);
and U2758 (N_2758,N_1817,N_1661);
nand U2759 (N_2759,N_1107,N_1165);
nor U2760 (N_2760,N_1364,N_1363);
nor U2761 (N_2761,N_1348,N_1152);
or U2762 (N_2762,N_1130,N_1210);
nand U2763 (N_2763,N_1912,N_1031);
nor U2764 (N_2764,N_1277,N_1164);
nand U2765 (N_2765,N_1733,N_1544);
and U2766 (N_2766,N_1834,N_1003);
nand U2767 (N_2767,N_1696,N_1348);
and U2768 (N_2768,N_1503,N_1627);
nor U2769 (N_2769,N_1339,N_1713);
nand U2770 (N_2770,N_1970,N_1470);
nor U2771 (N_2771,N_1714,N_1710);
or U2772 (N_2772,N_1097,N_1781);
or U2773 (N_2773,N_1910,N_1251);
and U2774 (N_2774,N_1545,N_1593);
and U2775 (N_2775,N_1469,N_1977);
nand U2776 (N_2776,N_1632,N_1506);
nor U2777 (N_2777,N_1633,N_1456);
or U2778 (N_2778,N_1981,N_1098);
nand U2779 (N_2779,N_1419,N_1324);
nand U2780 (N_2780,N_1355,N_1252);
or U2781 (N_2781,N_1507,N_1200);
and U2782 (N_2782,N_1189,N_1299);
nand U2783 (N_2783,N_1185,N_1570);
nand U2784 (N_2784,N_1055,N_1563);
nand U2785 (N_2785,N_1026,N_1103);
or U2786 (N_2786,N_1538,N_1674);
and U2787 (N_2787,N_1973,N_1943);
nand U2788 (N_2788,N_1843,N_1416);
and U2789 (N_2789,N_1069,N_1514);
and U2790 (N_2790,N_1328,N_1337);
nand U2791 (N_2791,N_1740,N_1581);
nand U2792 (N_2792,N_1082,N_1923);
nand U2793 (N_2793,N_1978,N_1572);
nand U2794 (N_2794,N_1733,N_1652);
or U2795 (N_2795,N_1425,N_1330);
or U2796 (N_2796,N_1912,N_1934);
nand U2797 (N_2797,N_1650,N_1247);
nor U2798 (N_2798,N_1661,N_1943);
or U2799 (N_2799,N_1379,N_1526);
or U2800 (N_2800,N_1532,N_1844);
and U2801 (N_2801,N_1052,N_1640);
nand U2802 (N_2802,N_1141,N_1938);
and U2803 (N_2803,N_1700,N_1281);
and U2804 (N_2804,N_1411,N_1957);
nor U2805 (N_2805,N_1989,N_1753);
or U2806 (N_2806,N_1932,N_1065);
nor U2807 (N_2807,N_1673,N_1727);
nand U2808 (N_2808,N_1086,N_1431);
nor U2809 (N_2809,N_1572,N_1121);
and U2810 (N_2810,N_1874,N_1065);
or U2811 (N_2811,N_1646,N_1092);
nor U2812 (N_2812,N_1942,N_1357);
or U2813 (N_2813,N_1648,N_1963);
nor U2814 (N_2814,N_1181,N_1129);
and U2815 (N_2815,N_1647,N_1177);
nor U2816 (N_2816,N_1421,N_1383);
nor U2817 (N_2817,N_1566,N_1777);
and U2818 (N_2818,N_1698,N_1569);
nand U2819 (N_2819,N_1954,N_1045);
or U2820 (N_2820,N_1165,N_1819);
nor U2821 (N_2821,N_1790,N_1046);
or U2822 (N_2822,N_1168,N_1680);
and U2823 (N_2823,N_1692,N_1804);
nor U2824 (N_2824,N_1088,N_1494);
or U2825 (N_2825,N_1412,N_1453);
and U2826 (N_2826,N_1683,N_1833);
and U2827 (N_2827,N_1400,N_1056);
and U2828 (N_2828,N_1362,N_1599);
nand U2829 (N_2829,N_1352,N_1324);
nand U2830 (N_2830,N_1949,N_1926);
or U2831 (N_2831,N_1857,N_1408);
nand U2832 (N_2832,N_1402,N_1341);
nand U2833 (N_2833,N_1711,N_1694);
nor U2834 (N_2834,N_1614,N_1156);
nor U2835 (N_2835,N_1622,N_1303);
or U2836 (N_2836,N_1315,N_1971);
nand U2837 (N_2837,N_1390,N_1781);
nand U2838 (N_2838,N_1140,N_1651);
and U2839 (N_2839,N_1787,N_1974);
and U2840 (N_2840,N_1019,N_1563);
nand U2841 (N_2841,N_1512,N_1874);
nand U2842 (N_2842,N_1503,N_1226);
and U2843 (N_2843,N_1404,N_1643);
or U2844 (N_2844,N_1009,N_1409);
or U2845 (N_2845,N_1768,N_1317);
or U2846 (N_2846,N_1308,N_1846);
or U2847 (N_2847,N_1062,N_1429);
nor U2848 (N_2848,N_1033,N_1171);
and U2849 (N_2849,N_1773,N_1466);
and U2850 (N_2850,N_1021,N_1496);
or U2851 (N_2851,N_1718,N_1087);
nand U2852 (N_2852,N_1905,N_1187);
nor U2853 (N_2853,N_1992,N_1508);
and U2854 (N_2854,N_1573,N_1610);
nor U2855 (N_2855,N_1384,N_1053);
or U2856 (N_2856,N_1487,N_1479);
nand U2857 (N_2857,N_1623,N_1153);
nor U2858 (N_2858,N_1974,N_1124);
and U2859 (N_2859,N_1804,N_1361);
and U2860 (N_2860,N_1297,N_1594);
nor U2861 (N_2861,N_1808,N_1650);
or U2862 (N_2862,N_1563,N_1985);
and U2863 (N_2863,N_1495,N_1590);
and U2864 (N_2864,N_1962,N_1108);
nor U2865 (N_2865,N_1835,N_1504);
or U2866 (N_2866,N_1184,N_1944);
nand U2867 (N_2867,N_1077,N_1189);
and U2868 (N_2868,N_1599,N_1051);
nand U2869 (N_2869,N_1519,N_1281);
nand U2870 (N_2870,N_1475,N_1418);
and U2871 (N_2871,N_1341,N_1867);
nor U2872 (N_2872,N_1353,N_1541);
nor U2873 (N_2873,N_1872,N_1665);
and U2874 (N_2874,N_1811,N_1167);
nand U2875 (N_2875,N_1343,N_1125);
or U2876 (N_2876,N_1195,N_1866);
or U2877 (N_2877,N_1899,N_1319);
and U2878 (N_2878,N_1745,N_1087);
and U2879 (N_2879,N_1338,N_1214);
nor U2880 (N_2880,N_1310,N_1798);
or U2881 (N_2881,N_1624,N_1424);
nor U2882 (N_2882,N_1891,N_1393);
nor U2883 (N_2883,N_1700,N_1104);
nor U2884 (N_2884,N_1591,N_1137);
nand U2885 (N_2885,N_1127,N_1322);
and U2886 (N_2886,N_1058,N_1159);
or U2887 (N_2887,N_1371,N_1648);
nand U2888 (N_2888,N_1066,N_1364);
nand U2889 (N_2889,N_1812,N_1488);
nor U2890 (N_2890,N_1018,N_1406);
and U2891 (N_2891,N_1383,N_1946);
or U2892 (N_2892,N_1694,N_1774);
or U2893 (N_2893,N_1579,N_1526);
or U2894 (N_2894,N_1439,N_1549);
and U2895 (N_2895,N_1761,N_1420);
or U2896 (N_2896,N_1215,N_1542);
nand U2897 (N_2897,N_1159,N_1001);
or U2898 (N_2898,N_1027,N_1249);
nand U2899 (N_2899,N_1713,N_1232);
and U2900 (N_2900,N_1421,N_1289);
or U2901 (N_2901,N_1002,N_1326);
and U2902 (N_2902,N_1051,N_1765);
and U2903 (N_2903,N_1232,N_1978);
or U2904 (N_2904,N_1640,N_1229);
and U2905 (N_2905,N_1766,N_1513);
or U2906 (N_2906,N_1440,N_1388);
and U2907 (N_2907,N_1434,N_1879);
or U2908 (N_2908,N_1547,N_1216);
or U2909 (N_2909,N_1792,N_1851);
and U2910 (N_2910,N_1830,N_1268);
nand U2911 (N_2911,N_1935,N_1638);
nor U2912 (N_2912,N_1178,N_1072);
or U2913 (N_2913,N_1356,N_1200);
or U2914 (N_2914,N_1662,N_1956);
or U2915 (N_2915,N_1680,N_1916);
nand U2916 (N_2916,N_1972,N_1709);
nand U2917 (N_2917,N_1185,N_1753);
or U2918 (N_2918,N_1084,N_1901);
or U2919 (N_2919,N_1112,N_1945);
nand U2920 (N_2920,N_1044,N_1627);
and U2921 (N_2921,N_1921,N_1133);
nor U2922 (N_2922,N_1114,N_1043);
and U2923 (N_2923,N_1451,N_1896);
or U2924 (N_2924,N_1871,N_1811);
nand U2925 (N_2925,N_1525,N_1974);
nand U2926 (N_2926,N_1515,N_1613);
and U2927 (N_2927,N_1220,N_1821);
nor U2928 (N_2928,N_1914,N_1911);
and U2929 (N_2929,N_1419,N_1589);
nand U2930 (N_2930,N_1932,N_1084);
or U2931 (N_2931,N_1998,N_1239);
or U2932 (N_2932,N_1705,N_1484);
nand U2933 (N_2933,N_1174,N_1607);
or U2934 (N_2934,N_1292,N_1358);
nor U2935 (N_2935,N_1818,N_1579);
or U2936 (N_2936,N_1840,N_1422);
and U2937 (N_2937,N_1122,N_1053);
nand U2938 (N_2938,N_1616,N_1990);
nand U2939 (N_2939,N_1748,N_1763);
nor U2940 (N_2940,N_1572,N_1993);
nor U2941 (N_2941,N_1232,N_1181);
or U2942 (N_2942,N_1137,N_1665);
nand U2943 (N_2943,N_1246,N_1421);
and U2944 (N_2944,N_1001,N_1061);
nor U2945 (N_2945,N_1542,N_1645);
and U2946 (N_2946,N_1150,N_1018);
nor U2947 (N_2947,N_1288,N_1676);
or U2948 (N_2948,N_1269,N_1259);
and U2949 (N_2949,N_1097,N_1293);
nor U2950 (N_2950,N_1142,N_1386);
and U2951 (N_2951,N_1758,N_1259);
or U2952 (N_2952,N_1736,N_1510);
and U2953 (N_2953,N_1444,N_1941);
nor U2954 (N_2954,N_1463,N_1819);
and U2955 (N_2955,N_1276,N_1469);
nand U2956 (N_2956,N_1112,N_1047);
nand U2957 (N_2957,N_1659,N_1050);
and U2958 (N_2958,N_1025,N_1409);
xor U2959 (N_2959,N_1193,N_1517);
or U2960 (N_2960,N_1764,N_1740);
or U2961 (N_2961,N_1834,N_1932);
or U2962 (N_2962,N_1844,N_1565);
nor U2963 (N_2963,N_1387,N_1578);
or U2964 (N_2964,N_1415,N_1401);
or U2965 (N_2965,N_1727,N_1903);
nand U2966 (N_2966,N_1817,N_1903);
nand U2967 (N_2967,N_1601,N_1864);
nand U2968 (N_2968,N_1039,N_1197);
nand U2969 (N_2969,N_1908,N_1240);
xor U2970 (N_2970,N_1492,N_1886);
and U2971 (N_2971,N_1887,N_1956);
nor U2972 (N_2972,N_1158,N_1606);
nor U2973 (N_2973,N_1966,N_1955);
or U2974 (N_2974,N_1506,N_1747);
nor U2975 (N_2975,N_1059,N_1902);
nand U2976 (N_2976,N_1476,N_1743);
or U2977 (N_2977,N_1431,N_1692);
or U2978 (N_2978,N_1132,N_1386);
and U2979 (N_2979,N_1757,N_1417);
nand U2980 (N_2980,N_1299,N_1121);
or U2981 (N_2981,N_1756,N_1297);
nand U2982 (N_2982,N_1747,N_1826);
nor U2983 (N_2983,N_1886,N_1112);
or U2984 (N_2984,N_1036,N_1287);
nor U2985 (N_2985,N_1682,N_1731);
xnor U2986 (N_2986,N_1885,N_1070);
and U2987 (N_2987,N_1333,N_1407);
nand U2988 (N_2988,N_1726,N_1913);
or U2989 (N_2989,N_1276,N_1643);
nor U2990 (N_2990,N_1431,N_1847);
and U2991 (N_2991,N_1725,N_1916);
nor U2992 (N_2992,N_1494,N_1044);
and U2993 (N_2993,N_1168,N_1461);
or U2994 (N_2994,N_1200,N_1503);
and U2995 (N_2995,N_1908,N_1392);
and U2996 (N_2996,N_1826,N_1573);
nand U2997 (N_2997,N_1082,N_1267);
or U2998 (N_2998,N_1272,N_1533);
and U2999 (N_2999,N_1908,N_1628);
or U3000 (N_3000,N_2084,N_2568);
or U3001 (N_3001,N_2092,N_2427);
and U3002 (N_3002,N_2796,N_2836);
nor U3003 (N_3003,N_2213,N_2718);
and U3004 (N_3004,N_2663,N_2336);
nor U3005 (N_3005,N_2957,N_2494);
and U3006 (N_3006,N_2536,N_2126);
nand U3007 (N_3007,N_2540,N_2178);
nor U3008 (N_3008,N_2408,N_2260);
nor U3009 (N_3009,N_2877,N_2592);
or U3010 (N_3010,N_2095,N_2969);
nor U3011 (N_3011,N_2374,N_2087);
nand U3012 (N_3012,N_2563,N_2973);
and U3013 (N_3013,N_2338,N_2489);
or U3014 (N_3014,N_2464,N_2797);
or U3015 (N_3015,N_2813,N_2546);
and U3016 (N_3016,N_2460,N_2693);
nor U3017 (N_3017,N_2418,N_2934);
nand U3018 (N_3018,N_2500,N_2620);
and U3019 (N_3019,N_2597,N_2520);
or U3020 (N_3020,N_2284,N_2577);
nor U3021 (N_3021,N_2586,N_2791);
or U3022 (N_3022,N_2595,N_2628);
nand U3023 (N_3023,N_2208,N_2661);
nand U3024 (N_3024,N_2274,N_2676);
or U3025 (N_3025,N_2825,N_2267);
and U3026 (N_3026,N_2329,N_2962);
nand U3027 (N_3027,N_2647,N_2868);
or U3028 (N_3028,N_2901,N_2051);
nand U3029 (N_3029,N_2006,N_2042);
or U3030 (N_3030,N_2701,N_2148);
nand U3031 (N_3031,N_2780,N_2610);
nor U3032 (N_3032,N_2776,N_2856);
nand U3033 (N_3033,N_2379,N_2264);
or U3034 (N_3034,N_2930,N_2407);
nor U3035 (N_3035,N_2687,N_2063);
nor U3036 (N_3036,N_2085,N_2448);
nor U3037 (N_3037,N_2712,N_2668);
nand U3038 (N_3038,N_2831,N_2872);
nor U3039 (N_3039,N_2059,N_2483);
or U3040 (N_3040,N_2176,N_2435);
and U3041 (N_3041,N_2392,N_2140);
or U3042 (N_3042,N_2649,N_2562);
or U3043 (N_3043,N_2220,N_2139);
nand U3044 (N_3044,N_2508,N_2088);
nand U3045 (N_3045,N_2770,N_2972);
or U3046 (N_3046,N_2576,N_2943);
nand U3047 (N_3047,N_2565,N_2533);
nor U3048 (N_3048,N_2790,N_2522);
or U3049 (N_3049,N_2204,N_2294);
nor U3050 (N_3050,N_2710,N_2600);
nand U3051 (N_3051,N_2990,N_2099);
and U3052 (N_3052,N_2775,N_2293);
and U3053 (N_3053,N_2297,N_2918);
and U3054 (N_3054,N_2240,N_2965);
nor U3055 (N_3055,N_2823,N_2396);
nor U3056 (N_3056,N_2230,N_2206);
nor U3057 (N_3057,N_2870,N_2594);
and U3058 (N_3058,N_2763,N_2190);
nor U3059 (N_3059,N_2587,N_2133);
and U3060 (N_3060,N_2585,N_2377);
or U3061 (N_3061,N_2802,N_2300);
and U3062 (N_3062,N_2409,N_2228);
and U3063 (N_3063,N_2781,N_2584);
or U3064 (N_3064,N_2094,N_2170);
nor U3065 (N_3065,N_2955,N_2517);
or U3066 (N_3066,N_2681,N_2008);
nor U3067 (N_3067,N_2765,N_2837);
nand U3068 (N_3068,N_2547,N_2299);
or U3069 (N_3069,N_2977,N_2337);
nor U3070 (N_3070,N_2175,N_2469);
xor U3071 (N_3071,N_2147,N_2201);
nor U3072 (N_3072,N_2015,N_2214);
or U3073 (N_3073,N_2524,N_2958);
nand U3074 (N_3074,N_2160,N_2513);
nor U3075 (N_3075,N_2224,N_2075);
nor U3076 (N_3076,N_2366,N_2673);
and U3077 (N_3077,N_2455,N_2196);
or U3078 (N_3078,N_2321,N_2864);
nand U3079 (N_3079,N_2161,N_2983);
and U3080 (N_3080,N_2376,N_2117);
or U3081 (N_3081,N_2182,N_2618);
and U3082 (N_3082,N_2428,N_2716);
nand U3083 (N_3083,N_2675,N_2027);
nor U3084 (N_3084,N_2128,N_2330);
or U3085 (N_3085,N_2940,N_2458);
nand U3086 (N_3086,N_2726,N_2028);
or U3087 (N_3087,N_2165,N_2475);
nand U3088 (N_3088,N_2273,N_2920);
nor U3089 (N_3089,N_2159,N_2662);
nand U3090 (N_3090,N_2880,N_2899);
or U3091 (N_3091,N_2022,N_2558);
or U3092 (N_3092,N_2306,N_2660);
and U3093 (N_3093,N_2553,N_2760);
and U3094 (N_3094,N_2741,N_2793);
nor U3095 (N_3095,N_2077,N_2656);
or U3096 (N_3096,N_2890,N_2310);
nand U3097 (N_3097,N_2941,N_2733);
nand U3098 (N_3098,N_2646,N_2949);
nand U3099 (N_3099,N_2689,N_2367);
nand U3100 (N_3100,N_2682,N_2002);
nor U3101 (N_3101,N_2185,N_2272);
nand U3102 (N_3102,N_2739,N_2542);
nand U3103 (N_3103,N_2303,N_2071);
and U3104 (N_3104,N_2928,N_2501);
nor U3105 (N_3105,N_2617,N_2061);
nor U3106 (N_3106,N_2976,N_2188);
and U3107 (N_3107,N_2218,N_2664);
nand U3108 (N_3108,N_2679,N_2242);
nand U3109 (N_3109,N_2420,N_2353);
nor U3110 (N_3110,N_2065,N_2062);
and U3111 (N_3111,N_2704,N_2232);
nor U3112 (N_3112,N_2745,N_2179);
xnor U3113 (N_3113,N_2578,N_2343);
and U3114 (N_3114,N_2157,N_2609);
nand U3115 (N_3115,N_2912,N_2442);
nand U3116 (N_3116,N_2657,N_2688);
nand U3117 (N_3117,N_2554,N_2270);
nor U3118 (N_3118,N_2491,N_2351);
and U3119 (N_3119,N_2531,N_2634);
nand U3120 (N_3120,N_2740,N_2108);
and U3121 (N_3121,N_2255,N_2843);
and U3122 (N_3122,N_2807,N_2285);
nand U3123 (N_3123,N_2691,N_2527);
or U3124 (N_3124,N_2980,N_2871);
nand U3125 (N_3125,N_2699,N_2951);
or U3126 (N_3126,N_2219,N_2380);
and U3127 (N_3127,N_2607,N_2915);
nand U3128 (N_3128,N_2332,N_2695);
nand U3129 (N_3129,N_2486,N_2938);
or U3130 (N_3130,N_2979,N_2080);
nor U3131 (N_3131,N_2044,N_2583);
nor U3132 (N_3132,N_2144,N_2093);
nand U3133 (N_3133,N_2750,N_2589);
or U3134 (N_3134,N_2867,N_2068);
nand U3135 (N_3135,N_2417,N_2411);
or U3136 (N_3136,N_2234,N_2452);
or U3137 (N_3137,N_2598,N_2164);
or U3138 (N_3138,N_2150,N_2771);
xor U3139 (N_3139,N_2963,N_2368);
nor U3140 (N_3140,N_2993,N_2569);
and U3141 (N_3141,N_2119,N_2623);
and U3142 (N_3142,N_2987,N_2324);
nor U3143 (N_3143,N_2423,N_2279);
nor U3144 (N_3144,N_2091,N_2838);
and U3145 (N_3145,N_2395,N_2443);
and U3146 (N_3146,N_2801,N_2152);
nor U3147 (N_3147,N_2064,N_2961);
and U3148 (N_3148,N_2249,N_2195);
nor U3149 (N_3149,N_2855,N_2142);
and U3150 (N_3150,N_2803,N_2528);
and U3151 (N_3151,N_2764,N_2111);
nor U3152 (N_3152,N_2135,N_2895);
nor U3153 (N_3153,N_2734,N_2629);
and U3154 (N_3154,N_2282,N_2931);
and U3155 (N_3155,N_2136,N_2824);
and U3156 (N_3156,N_2419,N_2535);
and U3157 (N_3157,N_2809,N_2852);
nand U3158 (N_3158,N_2308,N_2298);
and U3159 (N_3159,N_2177,N_2007);
and U3160 (N_3160,N_2606,N_2919);
or U3161 (N_3161,N_2341,N_2069);
nor U3162 (N_3162,N_2883,N_2317);
and U3163 (N_3163,N_2821,N_2881);
nand U3164 (N_3164,N_2907,N_2143);
and U3165 (N_3165,N_2348,N_2205);
and U3166 (N_3166,N_2914,N_2118);
and U3167 (N_3167,N_2327,N_2216);
or U3168 (N_3168,N_2480,N_2888);
or U3169 (N_3169,N_2451,N_2197);
or U3170 (N_3170,N_2243,N_2638);
nor U3171 (N_3171,N_2252,N_2616);
or U3172 (N_3172,N_2596,N_2670);
nand U3173 (N_3173,N_2246,N_2104);
nand U3174 (N_3174,N_2459,N_2581);
or U3175 (N_3175,N_2039,N_2835);
and U3176 (N_3176,N_2658,N_2354);
and U3177 (N_3177,N_2677,N_2371);
and U3178 (N_3178,N_2253,N_2643);
nand U3179 (N_3179,N_2544,N_2081);
or U3180 (N_3180,N_2356,N_2570);
or U3181 (N_3181,N_2806,N_2373);
or U3182 (N_3182,N_2112,N_2916);
or U3183 (N_3183,N_2711,N_2946);
and U3184 (N_3184,N_2456,N_2241);
nor U3185 (N_3185,N_2192,N_2873);
nor U3186 (N_3186,N_2405,N_2302);
or U3187 (N_3187,N_2262,N_2360);
or U3188 (N_3188,N_2259,N_2786);
and U3189 (N_3189,N_2706,N_2991);
or U3190 (N_3190,N_2614,N_2625);
or U3191 (N_3191,N_2653,N_2060);
and U3192 (N_3192,N_2278,N_2678);
or U3193 (N_3193,N_2684,N_2445);
nor U3194 (N_3194,N_2511,N_2738);
or U3195 (N_3195,N_2903,N_2097);
nor U3196 (N_3196,N_2257,N_2275);
nor U3197 (N_3197,N_2296,N_2690);
nand U3198 (N_3198,N_2572,N_2212);
nand U3199 (N_3199,N_2326,N_2879);
nor U3200 (N_3200,N_2277,N_2495);
and U3201 (N_3201,N_2359,N_2410);
nor U3202 (N_3202,N_2818,N_2424);
and U3203 (N_3203,N_2441,N_2107);
and U3204 (N_3204,N_2050,N_2548);
or U3205 (N_3205,N_2847,N_2258);
nand U3206 (N_3206,N_2537,N_2902);
and U3207 (N_3207,N_2530,N_2462);
or U3208 (N_3208,N_2265,N_2842);
nand U3209 (N_3209,N_2030,N_2925);
or U3210 (N_3210,N_2320,N_2696);
or U3211 (N_3211,N_2671,N_2913);
nand U3212 (N_3212,N_2636,N_2101);
nor U3213 (N_3213,N_2023,N_2429);
and U3214 (N_3214,N_2156,N_2444);
and U3215 (N_3215,N_2454,N_2287);
nand U3216 (N_3216,N_2950,N_2053);
or U3217 (N_3217,N_2848,N_2523);
nor U3218 (N_3218,N_2100,N_2134);
nand U3219 (N_3219,N_2127,N_2897);
and U3220 (N_3220,N_2431,N_2947);
or U3221 (N_3221,N_2624,N_2552);
nor U3222 (N_3222,N_2519,N_2762);
and U3223 (N_3223,N_2072,N_2013);
or U3224 (N_3224,N_2492,N_2685);
or U3225 (N_3225,N_2404,N_2295);
nor U3226 (N_3226,N_2882,N_2816);
nor U3227 (N_3227,N_2635,N_2334);
nor U3228 (N_3228,N_2398,N_2922);
and U3229 (N_3229,N_2948,N_2884);
nand U3230 (N_3230,N_2729,N_2966);
and U3231 (N_3231,N_2244,N_2892);
or U3232 (N_3232,N_2854,N_2439);
nor U3233 (N_3233,N_2309,N_2438);
and U3234 (N_3234,N_2481,N_2998);
or U3235 (N_3235,N_2588,N_2952);
and U3236 (N_3236,N_2774,N_2102);
or U3237 (N_3237,N_2611,N_2056);
and U3238 (N_3238,N_2746,N_2844);
and U3239 (N_3239,N_2543,N_2939);
nand U3240 (N_3240,N_2680,N_2782);
nand U3241 (N_3241,N_2927,N_2840);
nor U3242 (N_3242,N_2271,N_2832);
and U3243 (N_3243,N_2217,N_2488);
and U3244 (N_3244,N_2288,N_2981);
nand U3245 (N_3245,N_2619,N_2043);
nor U3246 (N_3246,N_2394,N_2123);
and U3247 (N_3247,N_2613,N_2414);
or U3248 (N_3248,N_2532,N_2659);
or U3249 (N_3249,N_2505,N_2328);
or U3250 (N_3250,N_2942,N_2978);
or U3251 (N_3251,N_2667,N_2034);
nand U3252 (N_3252,N_2145,N_2999);
or U3253 (N_3253,N_2186,N_2346);
nand U3254 (N_3254,N_2052,N_2026);
and U3255 (N_3255,N_2250,N_2732);
and U3256 (N_3256,N_2518,N_2471);
nand U3257 (N_3257,N_2316,N_2383);
or U3258 (N_3258,N_2105,N_2058);
nor U3259 (N_3259,N_2057,N_2453);
or U3260 (N_3260,N_2132,N_2385);
and U3261 (N_3261,N_2450,N_2375);
or U3262 (N_3262,N_2603,N_2526);
nand U3263 (N_3263,N_2485,N_2342);
nand U3264 (N_3264,N_2361,N_2564);
nand U3265 (N_3265,N_2633,N_2698);
nor U3266 (N_3266,N_2004,N_2365);
and U3267 (N_3267,N_2432,N_2792);
nand U3268 (N_3268,N_2210,N_2207);
or U3269 (N_3269,N_2641,N_2289);
and U3270 (N_3270,N_2755,N_2041);
or U3271 (N_3271,N_2756,N_2974);
nand U3272 (N_3272,N_2810,N_2074);
and U3273 (N_3273,N_2067,N_2758);
and U3274 (N_3274,N_2735,N_2031);
or U3275 (N_3275,N_2312,N_2369);
nor U3276 (N_3276,N_2109,N_2171);
or U3277 (N_3277,N_2124,N_2715);
or U3278 (N_3278,N_2778,N_2233);
nand U3279 (N_3279,N_2968,N_2163);
and U3280 (N_3280,N_2672,N_2499);
nor U3281 (N_3281,N_2509,N_2425);
or U3282 (N_3282,N_2358,N_2650);
or U3283 (N_3283,N_2223,N_2665);
or U3284 (N_3284,N_2291,N_2339);
nand U3285 (N_3285,N_2637,N_2076);
nor U3286 (N_3286,N_2751,N_2169);
nor U3287 (N_3287,N_2073,N_2545);
nand U3288 (N_3288,N_2040,N_2640);
or U3289 (N_3289,N_2988,N_2604);
nand U3290 (N_3290,N_2994,N_2386);
nor U3291 (N_3291,N_2493,N_2944);
or U3292 (N_3292,N_2904,N_2929);
nand U3293 (N_3293,N_2245,N_2773);
and U3294 (N_3294,N_2335,N_2263);
and U3295 (N_3295,N_2231,N_2347);
nand U3296 (N_3296,N_2183,N_2322);
and U3297 (N_3297,N_2754,N_2166);
and U3298 (N_3298,N_2016,N_2221);
or U3299 (N_3299,N_2959,N_2477);
nand U3300 (N_3300,N_2730,N_2029);
nor U3301 (N_3301,N_2211,N_2534);
or U3302 (N_3302,N_2490,N_2630);
and U3303 (N_3303,N_2997,N_2413);
nor U3304 (N_3304,N_2567,N_2817);
and U3305 (N_3305,N_2827,N_2591);
or U3306 (N_3306,N_2984,N_2047);
and U3307 (N_3307,N_2184,N_2719);
or U3308 (N_3308,N_2794,N_2172);
nand U3309 (N_3309,N_2005,N_2116);
or U3310 (N_3310,N_2174,N_2839);
or U3311 (N_3311,N_2858,N_2503);
nand U3312 (N_3312,N_2372,N_2752);
xor U3313 (N_3313,N_2612,N_2971);
nand U3314 (N_3314,N_2024,N_2953);
or U3315 (N_3315,N_2467,N_2686);
or U3316 (N_3316,N_2727,N_2149);
or U3317 (N_3317,N_2412,N_2254);
nor U3318 (N_3318,N_2402,N_2125);
xor U3319 (N_3319,N_2011,N_2502);
or U3320 (N_3320,N_2151,N_2863);
nor U3321 (N_3321,N_2787,N_2642);
and U3322 (N_3322,N_2122,N_2349);
nor U3323 (N_3323,N_2845,N_2020);
or U3324 (N_3324,N_2323,N_2602);
and U3325 (N_3325,N_2364,N_2639);
or U3326 (N_3326,N_2560,N_2559);
and U3327 (N_3327,N_2853,N_2648);
nor U3328 (N_3328,N_2860,N_2906);
or U3329 (N_3329,N_2666,N_2158);
nand U3330 (N_3330,N_2767,N_2785);
nand U3331 (N_3331,N_2894,N_2724);
nor U3332 (N_3332,N_2266,N_2399);
nor U3333 (N_3333,N_2580,N_2932);
nand U3334 (N_3334,N_2815,N_2021);
or U3335 (N_3335,N_2191,N_2292);
or U3336 (N_3336,N_2574,N_2311);
nand U3337 (N_3337,N_2910,N_2449);
or U3338 (N_3338,N_2889,N_2478);
and U3339 (N_3339,N_2822,N_2086);
and U3340 (N_3340,N_2593,N_2146);
and U3341 (N_3341,N_2761,N_2632);
nand U3342 (N_3342,N_2400,N_2529);
nor U3343 (N_3343,N_2886,N_2728);
or U3344 (N_3344,N_2748,N_2473);
nand U3345 (N_3345,N_2268,N_2301);
nor U3346 (N_3346,N_2304,N_2436);
nand U3347 (N_3347,N_2707,N_2115);
nor U3348 (N_3348,N_2887,N_2437);
nand U3349 (N_3349,N_2484,N_2226);
and U3350 (N_3350,N_2700,N_2089);
or U3351 (N_3351,N_2019,N_2601);
nand U3352 (N_3352,N_2120,N_2098);
nand U3353 (N_3353,N_2812,N_2238);
or U3354 (N_3354,N_2736,N_2430);
nand U3355 (N_3355,N_2645,N_2996);
nand U3356 (N_3356,N_2363,N_2964);
and U3357 (N_3357,N_2561,N_2202);
nand U3358 (N_3358,N_2970,N_2199);
or U3359 (N_3359,N_2256,N_2722);
nor U3360 (N_3360,N_2319,N_2893);
and U3361 (N_3361,N_2833,N_2237);
or U3362 (N_3362,N_2541,N_2849);
nor U3363 (N_3363,N_2391,N_2992);
nor U3364 (N_3364,N_2669,N_2819);
nor U3365 (N_3365,N_2539,N_2960);
or U3366 (N_3366,N_2384,N_2000);
nand U3367 (N_3367,N_2247,N_2236);
or U3368 (N_3368,N_2482,N_2422);
nand U3369 (N_3369,N_2851,N_2200);
or U3370 (N_3370,N_2744,N_2985);
or U3371 (N_3371,N_2433,N_2936);
or U3372 (N_3372,N_2113,N_2036);
nor U3373 (N_3373,N_2525,N_2045);
nand U3374 (N_3374,N_2440,N_2154);
nor U3375 (N_3375,N_2521,N_2713);
nor U3376 (N_3376,N_2516,N_2313);
or U3377 (N_3377,N_2721,N_2766);
or U3378 (N_3378,N_2605,N_2345);
nor U3379 (N_3379,N_2397,N_2788);
nor U3380 (N_3380,N_2350,N_2908);
nor U3381 (N_3381,N_2141,N_2155);
nor U3382 (N_3382,N_2479,N_2181);
nor U3383 (N_3383,N_2110,N_2504);
or U3384 (N_3384,N_2573,N_2498);
nor U3385 (N_3385,N_2194,N_2130);
and U3386 (N_3386,N_2869,N_2510);
nand U3387 (N_3387,N_2466,N_2193);
and U3388 (N_3388,N_2340,N_2674);
nor U3389 (N_3389,N_2911,N_2694);
nand U3390 (N_3390,N_2131,N_2079);
and U3391 (N_3391,N_2283,N_2692);
or U3392 (N_3392,N_2010,N_2626);
or U3393 (N_3393,N_2731,N_2401);
nand U3394 (N_3394,N_2239,N_2608);
nand U3395 (N_3395,N_2162,N_2697);
or U3396 (N_3396,N_2749,N_2468);
nand U3397 (N_3397,N_2012,N_2723);
nand U3398 (N_3398,N_2865,N_2954);
nor U3399 (N_3399,N_2875,N_2496);
and U3400 (N_3400,N_2702,N_2406);
nand U3401 (N_3401,N_2967,N_2476);
nand U3402 (N_3402,N_2579,N_2090);
and U3403 (N_3403,N_2917,N_2180);
or U3404 (N_3404,N_2269,N_2945);
nand U3405 (N_3405,N_2808,N_2106);
and U3406 (N_3406,N_2814,N_2209);
and U3407 (N_3407,N_2114,N_2924);
or U3408 (N_3408,N_2717,N_2507);
nand U3409 (N_3409,N_2261,N_2235);
nor U3410 (N_3410,N_2514,N_2286);
nor U3411 (N_3411,N_2862,N_2129);
or U3412 (N_3412,N_2599,N_2331);
nor U3413 (N_3413,N_2811,N_2307);
and U3414 (N_3414,N_2757,N_2557);
xnor U3415 (N_3415,N_2850,N_2001);
nand U3416 (N_3416,N_2772,N_2333);
or U3417 (N_3417,N_2829,N_2779);
nand U3418 (N_3418,N_2314,N_2229);
and U3419 (N_3419,N_2512,N_2550);
nand U3420 (N_3420,N_2820,N_2121);
and U3421 (N_3421,N_2644,N_2225);
or U3422 (N_3422,N_2470,N_2276);
nor U3423 (N_3423,N_2426,N_2248);
or U3424 (N_3424,N_2956,N_2742);
nor U3425 (N_3425,N_2168,N_2389);
nand U3426 (N_3426,N_2709,N_2070);
nand U3427 (N_3427,N_2382,N_2759);
nor U3428 (N_3428,N_2866,N_2403);
and U3429 (N_3429,N_2463,N_2048);
or U3430 (N_3430,N_2846,N_2800);
or U3431 (N_3431,N_2769,N_2859);
nand U3432 (N_3432,N_2357,N_2082);
or U3433 (N_3433,N_2799,N_2315);
and U3434 (N_3434,N_2447,N_2078);
or U3435 (N_3435,N_2390,N_2017);
nand U3436 (N_3436,N_2415,N_2898);
and U3437 (N_3437,N_2003,N_2487);
or U3438 (N_3438,N_2018,N_2655);
and U3439 (N_3439,N_2009,N_2652);
nand U3440 (N_3440,N_2777,N_2153);
nor U3441 (N_3441,N_2054,N_2874);
nand U3442 (N_3442,N_2798,N_2167);
xor U3443 (N_3443,N_2582,N_2055);
or U3444 (N_3444,N_2038,N_2506);
and U3445 (N_3445,N_2280,N_2861);
nor U3446 (N_3446,N_2651,N_2590);
and U3447 (N_3447,N_2986,N_2381);
nor U3448 (N_3448,N_2434,N_2876);
or U3449 (N_3449,N_2388,N_2137);
or U3450 (N_3450,N_2538,N_2352);
or U3451 (N_3451,N_2037,N_2621);
nand U3452 (N_3452,N_2631,N_2416);
and U3453 (N_3453,N_2905,N_2935);
or U3454 (N_3454,N_2215,N_2549);
nand U3455 (N_3455,N_2995,N_2189);
or U3456 (N_3456,N_2705,N_2753);
nand U3457 (N_3457,N_2203,N_2227);
or U3458 (N_3458,N_2923,N_2857);
or U3459 (N_3459,N_2515,N_2378);
or U3460 (N_3460,N_2251,N_2472);
nor U3461 (N_3461,N_2446,N_2325);
xor U3462 (N_3462,N_2461,N_2720);
or U3463 (N_3463,N_2066,N_2362);
and U3464 (N_3464,N_2556,N_2622);
nand U3465 (N_3465,N_2834,N_2355);
and U3466 (N_3466,N_2497,N_2198);
nor U3467 (N_3467,N_2222,N_2032);
nand U3468 (N_3468,N_2457,N_2465);
and U3469 (N_3469,N_2828,N_2937);
nand U3470 (N_3470,N_2900,N_2318);
and U3471 (N_3471,N_2138,N_2795);
and U3472 (N_3472,N_2784,N_2747);
xor U3473 (N_3473,N_2789,N_2344);
nor U3474 (N_3474,N_2387,N_2885);
and U3475 (N_3475,N_2708,N_2725);
nand U3476 (N_3476,N_2305,N_2896);
xor U3477 (N_3477,N_2683,N_2421);
nor U3478 (N_3478,N_2083,N_2025);
or U3479 (N_3479,N_2281,N_2049);
and U3480 (N_3480,N_2909,N_2737);
nand U3481 (N_3481,N_2783,N_2654);
and U3482 (N_3482,N_2551,N_2841);
or U3483 (N_3483,N_2370,N_2096);
nor U3484 (N_3484,N_2826,N_2555);
and U3485 (N_3485,N_2615,N_2891);
or U3486 (N_3486,N_2187,N_2703);
or U3487 (N_3487,N_2046,N_2173);
and U3488 (N_3488,N_2290,N_2933);
and U3489 (N_3489,N_2830,N_2627);
nand U3490 (N_3490,N_2982,N_2014);
or U3491 (N_3491,N_2575,N_2393);
nor U3492 (N_3492,N_2743,N_2989);
nor U3493 (N_3493,N_2975,N_2035);
nand U3494 (N_3494,N_2805,N_2804);
nor U3495 (N_3495,N_2878,N_2768);
nand U3496 (N_3496,N_2571,N_2921);
nand U3497 (N_3497,N_2103,N_2714);
or U3498 (N_3498,N_2474,N_2926);
nor U3499 (N_3499,N_2566,N_2033);
and U3500 (N_3500,N_2364,N_2282);
nand U3501 (N_3501,N_2483,N_2023);
and U3502 (N_3502,N_2887,N_2960);
xnor U3503 (N_3503,N_2125,N_2786);
or U3504 (N_3504,N_2129,N_2991);
nor U3505 (N_3505,N_2495,N_2498);
nand U3506 (N_3506,N_2640,N_2545);
and U3507 (N_3507,N_2726,N_2376);
nor U3508 (N_3508,N_2538,N_2753);
and U3509 (N_3509,N_2172,N_2829);
and U3510 (N_3510,N_2286,N_2557);
and U3511 (N_3511,N_2080,N_2686);
nand U3512 (N_3512,N_2292,N_2314);
and U3513 (N_3513,N_2327,N_2332);
and U3514 (N_3514,N_2721,N_2148);
or U3515 (N_3515,N_2758,N_2804);
or U3516 (N_3516,N_2793,N_2980);
nor U3517 (N_3517,N_2097,N_2175);
nor U3518 (N_3518,N_2274,N_2873);
nand U3519 (N_3519,N_2270,N_2275);
and U3520 (N_3520,N_2668,N_2158);
nor U3521 (N_3521,N_2547,N_2852);
nor U3522 (N_3522,N_2136,N_2692);
nor U3523 (N_3523,N_2267,N_2860);
nor U3524 (N_3524,N_2989,N_2389);
nor U3525 (N_3525,N_2421,N_2344);
or U3526 (N_3526,N_2554,N_2498);
or U3527 (N_3527,N_2512,N_2800);
nand U3528 (N_3528,N_2716,N_2174);
and U3529 (N_3529,N_2333,N_2233);
nor U3530 (N_3530,N_2335,N_2208);
nor U3531 (N_3531,N_2260,N_2863);
or U3532 (N_3532,N_2580,N_2341);
or U3533 (N_3533,N_2593,N_2113);
nand U3534 (N_3534,N_2892,N_2337);
nand U3535 (N_3535,N_2357,N_2555);
or U3536 (N_3536,N_2153,N_2665);
nand U3537 (N_3537,N_2235,N_2714);
and U3538 (N_3538,N_2307,N_2257);
or U3539 (N_3539,N_2294,N_2782);
nor U3540 (N_3540,N_2277,N_2031);
nand U3541 (N_3541,N_2056,N_2239);
and U3542 (N_3542,N_2660,N_2359);
xor U3543 (N_3543,N_2034,N_2502);
nand U3544 (N_3544,N_2816,N_2118);
nand U3545 (N_3545,N_2827,N_2556);
nor U3546 (N_3546,N_2140,N_2636);
nor U3547 (N_3547,N_2484,N_2379);
xor U3548 (N_3548,N_2482,N_2534);
nand U3549 (N_3549,N_2517,N_2255);
and U3550 (N_3550,N_2400,N_2954);
nand U3551 (N_3551,N_2180,N_2714);
nand U3552 (N_3552,N_2504,N_2522);
and U3553 (N_3553,N_2617,N_2654);
or U3554 (N_3554,N_2661,N_2123);
or U3555 (N_3555,N_2396,N_2438);
or U3556 (N_3556,N_2132,N_2039);
nor U3557 (N_3557,N_2812,N_2900);
nand U3558 (N_3558,N_2001,N_2716);
or U3559 (N_3559,N_2011,N_2900);
nand U3560 (N_3560,N_2402,N_2871);
or U3561 (N_3561,N_2614,N_2551);
nor U3562 (N_3562,N_2857,N_2026);
nand U3563 (N_3563,N_2308,N_2068);
and U3564 (N_3564,N_2031,N_2685);
xnor U3565 (N_3565,N_2446,N_2350);
nand U3566 (N_3566,N_2075,N_2938);
nor U3567 (N_3567,N_2572,N_2289);
nand U3568 (N_3568,N_2872,N_2498);
or U3569 (N_3569,N_2765,N_2212);
and U3570 (N_3570,N_2674,N_2292);
nand U3571 (N_3571,N_2671,N_2134);
and U3572 (N_3572,N_2624,N_2198);
or U3573 (N_3573,N_2164,N_2289);
or U3574 (N_3574,N_2399,N_2001);
nand U3575 (N_3575,N_2921,N_2445);
and U3576 (N_3576,N_2552,N_2229);
or U3577 (N_3577,N_2360,N_2208);
nor U3578 (N_3578,N_2771,N_2926);
and U3579 (N_3579,N_2763,N_2159);
nand U3580 (N_3580,N_2827,N_2293);
or U3581 (N_3581,N_2005,N_2001);
nor U3582 (N_3582,N_2762,N_2016);
nand U3583 (N_3583,N_2984,N_2306);
nor U3584 (N_3584,N_2401,N_2899);
nand U3585 (N_3585,N_2208,N_2784);
nand U3586 (N_3586,N_2137,N_2319);
and U3587 (N_3587,N_2621,N_2326);
or U3588 (N_3588,N_2654,N_2845);
nor U3589 (N_3589,N_2620,N_2564);
nand U3590 (N_3590,N_2065,N_2499);
nand U3591 (N_3591,N_2868,N_2729);
and U3592 (N_3592,N_2356,N_2827);
and U3593 (N_3593,N_2551,N_2225);
or U3594 (N_3594,N_2483,N_2455);
nor U3595 (N_3595,N_2333,N_2915);
or U3596 (N_3596,N_2268,N_2244);
nor U3597 (N_3597,N_2869,N_2922);
and U3598 (N_3598,N_2385,N_2480);
and U3599 (N_3599,N_2149,N_2197);
nand U3600 (N_3600,N_2883,N_2682);
nor U3601 (N_3601,N_2786,N_2062);
xnor U3602 (N_3602,N_2784,N_2214);
and U3603 (N_3603,N_2669,N_2682);
nor U3604 (N_3604,N_2671,N_2310);
nor U3605 (N_3605,N_2238,N_2690);
or U3606 (N_3606,N_2087,N_2397);
nand U3607 (N_3607,N_2379,N_2335);
xor U3608 (N_3608,N_2738,N_2213);
or U3609 (N_3609,N_2806,N_2764);
nand U3610 (N_3610,N_2308,N_2830);
and U3611 (N_3611,N_2645,N_2448);
or U3612 (N_3612,N_2488,N_2887);
and U3613 (N_3613,N_2381,N_2980);
xor U3614 (N_3614,N_2256,N_2414);
and U3615 (N_3615,N_2196,N_2873);
or U3616 (N_3616,N_2902,N_2291);
nor U3617 (N_3617,N_2456,N_2674);
or U3618 (N_3618,N_2101,N_2478);
or U3619 (N_3619,N_2336,N_2287);
nor U3620 (N_3620,N_2806,N_2011);
or U3621 (N_3621,N_2596,N_2569);
or U3622 (N_3622,N_2544,N_2112);
nor U3623 (N_3623,N_2741,N_2476);
nand U3624 (N_3624,N_2371,N_2303);
and U3625 (N_3625,N_2788,N_2254);
and U3626 (N_3626,N_2209,N_2572);
and U3627 (N_3627,N_2092,N_2429);
nor U3628 (N_3628,N_2347,N_2358);
nor U3629 (N_3629,N_2290,N_2161);
nand U3630 (N_3630,N_2359,N_2802);
and U3631 (N_3631,N_2787,N_2509);
nand U3632 (N_3632,N_2935,N_2097);
and U3633 (N_3633,N_2306,N_2378);
or U3634 (N_3634,N_2596,N_2010);
and U3635 (N_3635,N_2639,N_2700);
nand U3636 (N_3636,N_2428,N_2927);
and U3637 (N_3637,N_2087,N_2506);
nand U3638 (N_3638,N_2964,N_2174);
nor U3639 (N_3639,N_2012,N_2690);
or U3640 (N_3640,N_2562,N_2172);
and U3641 (N_3641,N_2221,N_2731);
nand U3642 (N_3642,N_2680,N_2023);
xor U3643 (N_3643,N_2187,N_2580);
and U3644 (N_3644,N_2334,N_2752);
and U3645 (N_3645,N_2103,N_2470);
and U3646 (N_3646,N_2145,N_2823);
or U3647 (N_3647,N_2246,N_2233);
or U3648 (N_3648,N_2125,N_2597);
and U3649 (N_3649,N_2489,N_2755);
nor U3650 (N_3650,N_2480,N_2372);
nor U3651 (N_3651,N_2843,N_2332);
nand U3652 (N_3652,N_2733,N_2913);
and U3653 (N_3653,N_2642,N_2041);
nand U3654 (N_3654,N_2108,N_2202);
nand U3655 (N_3655,N_2652,N_2083);
or U3656 (N_3656,N_2835,N_2063);
nand U3657 (N_3657,N_2370,N_2320);
and U3658 (N_3658,N_2601,N_2069);
nand U3659 (N_3659,N_2132,N_2694);
nor U3660 (N_3660,N_2736,N_2318);
or U3661 (N_3661,N_2154,N_2110);
nor U3662 (N_3662,N_2856,N_2416);
or U3663 (N_3663,N_2977,N_2263);
nor U3664 (N_3664,N_2311,N_2931);
nand U3665 (N_3665,N_2990,N_2133);
and U3666 (N_3666,N_2406,N_2913);
and U3667 (N_3667,N_2773,N_2000);
and U3668 (N_3668,N_2934,N_2260);
nand U3669 (N_3669,N_2896,N_2806);
and U3670 (N_3670,N_2886,N_2208);
and U3671 (N_3671,N_2637,N_2828);
nand U3672 (N_3672,N_2464,N_2627);
nand U3673 (N_3673,N_2875,N_2933);
nand U3674 (N_3674,N_2364,N_2349);
and U3675 (N_3675,N_2721,N_2722);
nor U3676 (N_3676,N_2130,N_2356);
nand U3677 (N_3677,N_2593,N_2904);
and U3678 (N_3678,N_2233,N_2813);
and U3679 (N_3679,N_2547,N_2713);
nor U3680 (N_3680,N_2301,N_2891);
nor U3681 (N_3681,N_2906,N_2450);
nand U3682 (N_3682,N_2054,N_2970);
and U3683 (N_3683,N_2123,N_2830);
nor U3684 (N_3684,N_2117,N_2059);
and U3685 (N_3685,N_2633,N_2370);
and U3686 (N_3686,N_2285,N_2468);
and U3687 (N_3687,N_2944,N_2256);
nand U3688 (N_3688,N_2818,N_2546);
or U3689 (N_3689,N_2773,N_2307);
nand U3690 (N_3690,N_2257,N_2574);
nand U3691 (N_3691,N_2822,N_2170);
or U3692 (N_3692,N_2537,N_2376);
nor U3693 (N_3693,N_2258,N_2015);
or U3694 (N_3694,N_2304,N_2659);
nand U3695 (N_3695,N_2049,N_2819);
and U3696 (N_3696,N_2268,N_2944);
nand U3697 (N_3697,N_2027,N_2525);
nand U3698 (N_3698,N_2063,N_2090);
nor U3699 (N_3699,N_2451,N_2358);
or U3700 (N_3700,N_2952,N_2126);
nor U3701 (N_3701,N_2528,N_2559);
or U3702 (N_3702,N_2617,N_2538);
and U3703 (N_3703,N_2273,N_2657);
and U3704 (N_3704,N_2970,N_2494);
nand U3705 (N_3705,N_2102,N_2757);
and U3706 (N_3706,N_2249,N_2546);
and U3707 (N_3707,N_2714,N_2660);
and U3708 (N_3708,N_2665,N_2177);
or U3709 (N_3709,N_2652,N_2359);
or U3710 (N_3710,N_2418,N_2555);
or U3711 (N_3711,N_2908,N_2038);
nand U3712 (N_3712,N_2422,N_2024);
nor U3713 (N_3713,N_2544,N_2180);
or U3714 (N_3714,N_2169,N_2851);
nand U3715 (N_3715,N_2709,N_2863);
nand U3716 (N_3716,N_2786,N_2708);
nor U3717 (N_3717,N_2092,N_2766);
or U3718 (N_3718,N_2676,N_2202);
nor U3719 (N_3719,N_2971,N_2916);
nand U3720 (N_3720,N_2335,N_2842);
nor U3721 (N_3721,N_2118,N_2721);
nand U3722 (N_3722,N_2319,N_2875);
or U3723 (N_3723,N_2821,N_2865);
nor U3724 (N_3724,N_2260,N_2008);
and U3725 (N_3725,N_2245,N_2159);
and U3726 (N_3726,N_2481,N_2940);
and U3727 (N_3727,N_2655,N_2753);
nor U3728 (N_3728,N_2262,N_2123);
nor U3729 (N_3729,N_2231,N_2355);
or U3730 (N_3730,N_2028,N_2766);
and U3731 (N_3731,N_2320,N_2451);
nand U3732 (N_3732,N_2052,N_2321);
and U3733 (N_3733,N_2390,N_2751);
or U3734 (N_3734,N_2183,N_2318);
and U3735 (N_3735,N_2437,N_2266);
nor U3736 (N_3736,N_2573,N_2310);
nor U3737 (N_3737,N_2422,N_2903);
nand U3738 (N_3738,N_2199,N_2048);
nand U3739 (N_3739,N_2379,N_2757);
or U3740 (N_3740,N_2790,N_2531);
nand U3741 (N_3741,N_2390,N_2333);
nand U3742 (N_3742,N_2714,N_2917);
and U3743 (N_3743,N_2480,N_2843);
nor U3744 (N_3744,N_2591,N_2678);
nor U3745 (N_3745,N_2244,N_2347);
or U3746 (N_3746,N_2626,N_2163);
nor U3747 (N_3747,N_2261,N_2466);
or U3748 (N_3748,N_2194,N_2339);
or U3749 (N_3749,N_2802,N_2494);
nand U3750 (N_3750,N_2767,N_2922);
and U3751 (N_3751,N_2357,N_2620);
nor U3752 (N_3752,N_2232,N_2327);
nor U3753 (N_3753,N_2226,N_2857);
nand U3754 (N_3754,N_2827,N_2263);
or U3755 (N_3755,N_2776,N_2633);
and U3756 (N_3756,N_2014,N_2940);
nand U3757 (N_3757,N_2856,N_2517);
nor U3758 (N_3758,N_2734,N_2969);
nand U3759 (N_3759,N_2126,N_2469);
nand U3760 (N_3760,N_2048,N_2793);
and U3761 (N_3761,N_2192,N_2096);
or U3762 (N_3762,N_2588,N_2887);
or U3763 (N_3763,N_2810,N_2880);
and U3764 (N_3764,N_2590,N_2147);
nor U3765 (N_3765,N_2077,N_2687);
and U3766 (N_3766,N_2256,N_2572);
or U3767 (N_3767,N_2912,N_2203);
nor U3768 (N_3768,N_2089,N_2032);
or U3769 (N_3769,N_2274,N_2672);
and U3770 (N_3770,N_2687,N_2545);
nor U3771 (N_3771,N_2338,N_2516);
nand U3772 (N_3772,N_2347,N_2260);
nor U3773 (N_3773,N_2293,N_2856);
nor U3774 (N_3774,N_2506,N_2717);
nor U3775 (N_3775,N_2111,N_2969);
and U3776 (N_3776,N_2997,N_2114);
nand U3777 (N_3777,N_2139,N_2124);
nor U3778 (N_3778,N_2937,N_2201);
nor U3779 (N_3779,N_2449,N_2037);
nor U3780 (N_3780,N_2771,N_2388);
and U3781 (N_3781,N_2199,N_2460);
nor U3782 (N_3782,N_2596,N_2115);
nor U3783 (N_3783,N_2347,N_2728);
and U3784 (N_3784,N_2183,N_2686);
nor U3785 (N_3785,N_2415,N_2919);
nor U3786 (N_3786,N_2487,N_2586);
nand U3787 (N_3787,N_2397,N_2855);
and U3788 (N_3788,N_2534,N_2576);
and U3789 (N_3789,N_2345,N_2011);
and U3790 (N_3790,N_2569,N_2872);
nand U3791 (N_3791,N_2662,N_2890);
and U3792 (N_3792,N_2712,N_2003);
or U3793 (N_3793,N_2900,N_2829);
nor U3794 (N_3794,N_2071,N_2364);
nand U3795 (N_3795,N_2401,N_2540);
nor U3796 (N_3796,N_2674,N_2210);
nor U3797 (N_3797,N_2475,N_2304);
or U3798 (N_3798,N_2860,N_2164);
nand U3799 (N_3799,N_2047,N_2704);
nand U3800 (N_3800,N_2742,N_2071);
or U3801 (N_3801,N_2768,N_2594);
nand U3802 (N_3802,N_2684,N_2504);
nor U3803 (N_3803,N_2149,N_2455);
nand U3804 (N_3804,N_2611,N_2135);
nand U3805 (N_3805,N_2090,N_2238);
or U3806 (N_3806,N_2365,N_2294);
or U3807 (N_3807,N_2349,N_2496);
or U3808 (N_3808,N_2058,N_2516);
nand U3809 (N_3809,N_2798,N_2254);
nor U3810 (N_3810,N_2956,N_2655);
nor U3811 (N_3811,N_2339,N_2011);
nand U3812 (N_3812,N_2067,N_2307);
nor U3813 (N_3813,N_2313,N_2937);
nand U3814 (N_3814,N_2962,N_2497);
and U3815 (N_3815,N_2543,N_2653);
and U3816 (N_3816,N_2204,N_2357);
nand U3817 (N_3817,N_2415,N_2701);
and U3818 (N_3818,N_2179,N_2308);
nand U3819 (N_3819,N_2056,N_2702);
and U3820 (N_3820,N_2015,N_2627);
nand U3821 (N_3821,N_2766,N_2689);
nor U3822 (N_3822,N_2227,N_2219);
nand U3823 (N_3823,N_2878,N_2191);
and U3824 (N_3824,N_2373,N_2969);
nor U3825 (N_3825,N_2143,N_2237);
and U3826 (N_3826,N_2394,N_2890);
nor U3827 (N_3827,N_2358,N_2825);
nor U3828 (N_3828,N_2348,N_2181);
or U3829 (N_3829,N_2863,N_2944);
and U3830 (N_3830,N_2791,N_2564);
and U3831 (N_3831,N_2807,N_2925);
nor U3832 (N_3832,N_2577,N_2959);
nand U3833 (N_3833,N_2660,N_2542);
and U3834 (N_3834,N_2827,N_2810);
nand U3835 (N_3835,N_2151,N_2120);
nand U3836 (N_3836,N_2541,N_2884);
nor U3837 (N_3837,N_2412,N_2289);
or U3838 (N_3838,N_2395,N_2217);
or U3839 (N_3839,N_2989,N_2910);
or U3840 (N_3840,N_2418,N_2615);
nor U3841 (N_3841,N_2734,N_2147);
nor U3842 (N_3842,N_2397,N_2911);
nor U3843 (N_3843,N_2505,N_2737);
nor U3844 (N_3844,N_2591,N_2700);
and U3845 (N_3845,N_2418,N_2769);
nor U3846 (N_3846,N_2564,N_2622);
and U3847 (N_3847,N_2645,N_2456);
and U3848 (N_3848,N_2352,N_2514);
nor U3849 (N_3849,N_2815,N_2561);
nand U3850 (N_3850,N_2823,N_2814);
nand U3851 (N_3851,N_2572,N_2097);
or U3852 (N_3852,N_2455,N_2395);
or U3853 (N_3853,N_2147,N_2343);
or U3854 (N_3854,N_2198,N_2501);
and U3855 (N_3855,N_2342,N_2659);
and U3856 (N_3856,N_2786,N_2356);
nand U3857 (N_3857,N_2567,N_2383);
nand U3858 (N_3858,N_2178,N_2049);
and U3859 (N_3859,N_2934,N_2003);
and U3860 (N_3860,N_2495,N_2686);
or U3861 (N_3861,N_2261,N_2338);
nor U3862 (N_3862,N_2220,N_2576);
nand U3863 (N_3863,N_2038,N_2861);
nand U3864 (N_3864,N_2718,N_2360);
nor U3865 (N_3865,N_2268,N_2212);
nor U3866 (N_3866,N_2803,N_2543);
nor U3867 (N_3867,N_2150,N_2651);
nor U3868 (N_3868,N_2445,N_2156);
or U3869 (N_3869,N_2377,N_2367);
nand U3870 (N_3870,N_2584,N_2346);
or U3871 (N_3871,N_2673,N_2440);
or U3872 (N_3872,N_2081,N_2304);
and U3873 (N_3873,N_2056,N_2991);
nor U3874 (N_3874,N_2588,N_2540);
nand U3875 (N_3875,N_2690,N_2595);
or U3876 (N_3876,N_2097,N_2910);
and U3877 (N_3877,N_2649,N_2458);
or U3878 (N_3878,N_2514,N_2133);
or U3879 (N_3879,N_2832,N_2332);
or U3880 (N_3880,N_2051,N_2632);
and U3881 (N_3881,N_2624,N_2867);
nand U3882 (N_3882,N_2074,N_2545);
nor U3883 (N_3883,N_2642,N_2619);
nand U3884 (N_3884,N_2261,N_2730);
and U3885 (N_3885,N_2019,N_2953);
and U3886 (N_3886,N_2572,N_2487);
nor U3887 (N_3887,N_2985,N_2017);
nor U3888 (N_3888,N_2608,N_2691);
nor U3889 (N_3889,N_2217,N_2187);
nor U3890 (N_3890,N_2710,N_2940);
or U3891 (N_3891,N_2502,N_2922);
nor U3892 (N_3892,N_2011,N_2343);
or U3893 (N_3893,N_2870,N_2764);
nand U3894 (N_3894,N_2846,N_2058);
and U3895 (N_3895,N_2337,N_2176);
or U3896 (N_3896,N_2016,N_2496);
and U3897 (N_3897,N_2830,N_2914);
or U3898 (N_3898,N_2678,N_2950);
and U3899 (N_3899,N_2257,N_2975);
or U3900 (N_3900,N_2735,N_2307);
nor U3901 (N_3901,N_2003,N_2732);
nor U3902 (N_3902,N_2611,N_2793);
nor U3903 (N_3903,N_2700,N_2887);
nor U3904 (N_3904,N_2698,N_2002);
nand U3905 (N_3905,N_2252,N_2871);
and U3906 (N_3906,N_2418,N_2914);
and U3907 (N_3907,N_2432,N_2104);
nand U3908 (N_3908,N_2085,N_2991);
or U3909 (N_3909,N_2157,N_2786);
and U3910 (N_3910,N_2891,N_2582);
nand U3911 (N_3911,N_2578,N_2229);
nand U3912 (N_3912,N_2000,N_2618);
and U3913 (N_3913,N_2978,N_2341);
or U3914 (N_3914,N_2001,N_2184);
nand U3915 (N_3915,N_2870,N_2877);
nand U3916 (N_3916,N_2707,N_2569);
nand U3917 (N_3917,N_2686,N_2059);
and U3918 (N_3918,N_2222,N_2517);
nand U3919 (N_3919,N_2493,N_2714);
xor U3920 (N_3920,N_2474,N_2463);
nand U3921 (N_3921,N_2297,N_2375);
or U3922 (N_3922,N_2941,N_2126);
nor U3923 (N_3923,N_2927,N_2514);
nand U3924 (N_3924,N_2478,N_2135);
nor U3925 (N_3925,N_2472,N_2512);
nor U3926 (N_3926,N_2317,N_2440);
nand U3927 (N_3927,N_2670,N_2250);
nor U3928 (N_3928,N_2856,N_2508);
nor U3929 (N_3929,N_2861,N_2488);
and U3930 (N_3930,N_2837,N_2619);
or U3931 (N_3931,N_2414,N_2513);
nand U3932 (N_3932,N_2637,N_2988);
nor U3933 (N_3933,N_2978,N_2317);
and U3934 (N_3934,N_2931,N_2491);
and U3935 (N_3935,N_2853,N_2003);
nand U3936 (N_3936,N_2724,N_2348);
nand U3937 (N_3937,N_2407,N_2912);
nor U3938 (N_3938,N_2027,N_2738);
nand U3939 (N_3939,N_2705,N_2997);
or U3940 (N_3940,N_2486,N_2200);
and U3941 (N_3941,N_2849,N_2706);
nor U3942 (N_3942,N_2754,N_2511);
and U3943 (N_3943,N_2085,N_2257);
nand U3944 (N_3944,N_2808,N_2816);
nor U3945 (N_3945,N_2468,N_2454);
nor U3946 (N_3946,N_2558,N_2362);
nand U3947 (N_3947,N_2745,N_2568);
or U3948 (N_3948,N_2773,N_2111);
and U3949 (N_3949,N_2117,N_2114);
or U3950 (N_3950,N_2374,N_2603);
or U3951 (N_3951,N_2404,N_2485);
or U3952 (N_3952,N_2809,N_2442);
nand U3953 (N_3953,N_2672,N_2402);
or U3954 (N_3954,N_2890,N_2332);
nor U3955 (N_3955,N_2704,N_2903);
nor U3956 (N_3956,N_2298,N_2025);
and U3957 (N_3957,N_2813,N_2512);
nor U3958 (N_3958,N_2886,N_2168);
nand U3959 (N_3959,N_2433,N_2162);
and U3960 (N_3960,N_2385,N_2135);
or U3961 (N_3961,N_2770,N_2124);
and U3962 (N_3962,N_2285,N_2262);
nor U3963 (N_3963,N_2500,N_2560);
nand U3964 (N_3964,N_2815,N_2250);
and U3965 (N_3965,N_2111,N_2771);
nor U3966 (N_3966,N_2025,N_2683);
and U3967 (N_3967,N_2773,N_2280);
or U3968 (N_3968,N_2381,N_2359);
nand U3969 (N_3969,N_2096,N_2308);
nor U3970 (N_3970,N_2173,N_2974);
nor U3971 (N_3971,N_2565,N_2814);
nand U3972 (N_3972,N_2651,N_2224);
nor U3973 (N_3973,N_2788,N_2024);
and U3974 (N_3974,N_2641,N_2805);
nor U3975 (N_3975,N_2522,N_2734);
and U3976 (N_3976,N_2893,N_2670);
nand U3977 (N_3977,N_2182,N_2230);
or U3978 (N_3978,N_2787,N_2227);
and U3979 (N_3979,N_2710,N_2492);
and U3980 (N_3980,N_2383,N_2974);
and U3981 (N_3981,N_2832,N_2239);
or U3982 (N_3982,N_2687,N_2695);
and U3983 (N_3983,N_2207,N_2368);
nor U3984 (N_3984,N_2260,N_2220);
and U3985 (N_3985,N_2809,N_2573);
nand U3986 (N_3986,N_2000,N_2942);
and U3987 (N_3987,N_2422,N_2094);
or U3988 (N_3988,N_2831,N_2051);
nor U3989 (N_3989,N_2460,N_2043);
nor U3990 (N_3990,N_2915,N_2591);
nor U3991 (N_3991,N_2299,N_2794);
nor U3992 (N_3992,N_2169,N_2612);
and U3993 (N_3993,N_2844,N_2036);
nor U3994 (N_3994,N_2947,N_2217);
nor U3995 (N_3995,N_2915,N_2455);
and U3996 (N_3996,N_2681,N_2873);
and U3997 (N_3997,N_2967,N_2947);
and U3998 (N_3998,N_2310,N_2629);
nand U3999 (N_3999,N_2199,N_2410);
nand U4000 (N_4000,N_3714,N_3835);
or U4001 (N_4001,N_3285,N_3863);
and U4002 (N_4002,N_3214,N_3810);
nor U4003 (N_4003,N_3941,N_3851);
xnor U4004 (N_4004,N_3157,N_3132);
nand U4005 (N_4005,N_3046,N_3592);
nand U4006 (N_4006,N_3893,N_3009);
nand U4007 (N_4007,N_3420,N_3746);
or U4008 (N_4008,N_3692,N_3717);
nand U4009 (N_4009,N_3805,N_3301);
nand U4010 (N_4010,N_3092,N_3059);
nor U4011 (N_4011,N_3277,N_3346);
or U4012 (N_4012,N_3077,N_3398);
nor U4013 (N_4013,N_3284,N_3133);
and U4014 (N_4014,N_3883,N_3821);
nor U4015 (N_4015,N_3709,N_3027);
nand U4016 (N_4016,N_3425,N_3933);
nand U4017 (N_4017,N_3704,N_3313);
or U4018 (N_4018,N_3584,N_3418);
or U4019 (N_4019,N_3292,N_3181);
and U4020 (N_4020,N_3140,N_3889);
and U4021 (N_4021,N_3200,N_3345);
nor U4022 (N_4022,N_3050,N_3256);
nor U4023 (N_4023,N_3659,N_3267);
or U4024 (N_4024,N_3696,N_3466);
xnor U4025 (N_4025,N_3397,N_3366);
nor U4026 (N_4026,N_3251,N_3839);
and U4027 (N_4027,N_3569,N_3379);
nor U4028 (N_4028,N_3886,N_3975);
or U4029 (N_4029,N_3706,N_3006);
nor U4030 (N_4030,N_3287,N_3739);
nor U4031 (N_4031,N_3773,N_3192);
nor U4032 (N_4032,N_3171,N_3517);
nand U4033 (N_4033,N_3344,N_3529);
nand U4034 (N_4034,N_3128,N_3608);
or U4035 (N_4035,N_3723,N_3678);
nor U4036 (N_4036,N_3900,N_3385);
nand U4037 (N_4037,N_3943,N_3628);
or U4038 (N_4038,N_3074,N_3088);
and U4039 (N_4039,N_3135,N_3813);
nand U4040 (N_4040,N_3745,N_3433);
or U4041 (N_4041,N_3486,N_3934);
or U4042 (N_4042,N_3511,N_3021);
xor U4043 (N_4043,N_3311,N_3986);
or U4044 (N_4044,N_3837,N_3896);
nand U4045 (N_4045,N_3514,N_3415);
nor U4046 (N_4046,N_3047,N_3829);
nand U4047 (N_4047,N_3333,N_3327);
nor U4048 (N_4048,N_3772,N_3364);
nor U4049 (N_4049,N_3349,N_3034);
or U4050 (N_4050,N_3208,N_3483);
and U4051 (N_4051,N_3743,N_3417);
or U4052 (N_4052,N_3775,N_3120);
and U4053 (N_4053,N_3556,N_3547);
or U4054 (N_4054,N_3961,N_3029);
nand U4055 (N_4055,N_3014,N_3347);
nor U4056 (N_4056,N_3676,N_3985);
or U4057 (N_4057,N_3968,N_3150);
or U4058 (N_4058,N_3023,N_3590);
nand U4059 (N_4059,N_3639,N_3010);
and U4060 (N_4060,N_3626,N_3165);
and U4061 (N_4061,N_3924,N_3691);
and U4062 (N_4062,N_3809,N_3532);
and U4063 (N_4063,N_3353,N_3081);
nand U4064 (N_4064,N_3158,N_3687);
nor U4065 (N_4065,N_3502,N_3155);
or U4066 (N_4066,N_3615,N_3020);
and U4067 (N_4067,N_3358,N_3248);
and U4068 (N_4068,N_3954,N_3348);
or U4069 (N_4069,N_3621,N_3847);
nor U4070 (N_4070,N_3053,N_3664);
and U4071 (N_4071,N_3751,N_3749);
nor U4072 (N_4072,N_3721,N_3573);
or U4073 (N_4073,N_3445,N_3151);
and U4074 (N_4074,N_3656,N_3060);
nand U4075 (N_4075,N_3784,N_3280);
nor U4076 (N_4076,N_3026,N_3808);
nand U4077 (N_4077,N_3763,N_3812);
nor U4078 (N_4078,N_3666,N_3949);
or U4079 (N_4079,N_3377,N_3310);
and U4080 (N_4080,N_3764,N_3295);
nor U4081 (N_4081,N_3566,N_3728);
and U4082 (N_4082,N_3903,N_3747);
nor U4083 (N_4083,N_3463,N_3218);
and U4084 (N_4084,N_3652,N_3734);
or U4085 (N_4085,N_3510,N_3370);
nor U4086 (N_4086,N_3507,N_3384);
or U4087 (N_4087,N_3634,N_3354);
nor U4088 (N_4088,N_3735,N_3738);
or U4089 (N_4089,N_3591,N_3530);
nand U4090 (N_4090,N_3874,N_3435);
nor U4091 (N_4091,N_3557,N_3799);
and U4092 (N_4092,N_3375,N_3552);
or U4093 (N_4093,N_3095,N_3603);
and U4094 (N_4094,N_3381,N_3176);
and U4095 (N_4095,N_3138,N_3712);
nand U4096 (N_4096,N_3841,N_3005);
nand U4097 (N_4097,N_3314,N_3802);
nor U4098 (N_4098,N_3336,N_3859);
nor U4099 (N_4099,N_3703,N_3307);
nor U4100 (N_4100,N_3493,N_3882);
nor U4101 (N_4101,N_3996,N_3660);
or U4102 (N_4102,N_3290,N_3054);
or U4103 (N_4103,N_3097,N_3693);
and U4104 (N_4104,N_3306,N_3167);
or U4105 (N_4105,N_3066,N_3318);
nand U4106 (N_4106,N_3561,N_3117);
nand U4107 (N_4107,N_3711,N_3250);
or U4108 (N_4108,N_3451,N_3540);
xor U4109 (N_4109,N_3684,N_3665);
nor U4110 (N_4110,N_3411,N_3645);
or U4111 (N_4111,N_3604,N_3786);
and U4112 (N_4112,N_3589,N_3689);
and U4113 (N_4113,N_3270,N_3672);
nor U4114 (N_4114,N_3679,N_3601);
or U4115 (N_4115,N_3793,N_3175);
or U4116 (N_4116,N_3559,N_3210);
and U4117 (N_4117,N_3025,N_3145);
nand U4118 (N_4118,N_3825,N_3118);
or U4119 (N_4119,N_3423,N_3362);
or U4120 (N_4120,N_3614,N_3106);
nand U4121 (N_4121,N_3455,N_3823);
or U4122 (N_4122,N_3472,N_3405);
and U4123 (N_4123,N_3112,N_3981);
nor U4124 (N_4124,N_3068,N_3154);
or U4125 (N_4125,N_3650,N_3352);
nor U4126 (N_4126,N_3441,N_3207);
and U4127 (N_4127,N_3962,N_3651);
nor U4128 (N_4128,N_3866,N_3197);
xor U4129 (N_4129,N_3759,N_3387);
xnor U4130 (N_4130,N_3035,N_3636);
and U4131 (N_4131,N_3419,N_3462);
nand U4132 (N_4132,N_3765,N_3555);
nor U4133 (N_4133,N_3072,N_3733);
or U4134 (N_4134,N_3872,N_3897);
nor U4135 (N_4135,N_3048,N_3906);
nand U4136 (N_4136,N_3550,N_3931);
or U4137 (N_4137,N_3811,N_3754);
nor U4138 (N_4138,N_3972,N_3041);
nand U4139 (N_4139,N_3350,N_3320);
and U4140 (N_4140,N_3568,N_3548);
nor U4141 (N_4141,N_3243,N_3824);
nand U4142 (N_4142,N_3663,N_3796);
and U4143 (N_4143,N_3259,N_3792);
nand U4144 (N_4144,N_3474,N_3096);
nand U4145 (N_4145,N_3803,N_3244);
and U4146 (N_4146,N_3351,N_3178);
or U4147 (N_4147,N_3720,N_3777);
nor U4148 (N_4148,N_3093,N_3580);
or U4149 (N_4149,N_3073,N_3952);
nand U4150 (N_4150,N_3944,N_3235);
nand U4151 (N_4151,N_3729,N_3432);
and U4152 (N_4152,N_3618,N_3141);
and U4153 (N_4153,N_3710,N_3646);
nand U4154 (N_4154,N_3281,N_3727);
nor U4155 (N_4155,N_3613,N_3399);
nor U4156 (N_4156,N_3937,N_3334);
nand U4157 (N_4157,N_3257,N_3667);
nor U4158 (N_4158,N_3518,N_3058);
and U4159 (N_4159,N_3031,N_3011);
nand U4160 (N_4160,N_3316,N_3448);
nor U4161 (N_4161,N_3304,N_3554);
nor U4162 (N_4162,N_3905,N_3857);
nand U4163 (N_4163,N_3409,N_3305);
nor U4164 (N_4164,N_3085,N_3459);
nand U4165 (N_4165,N_3852,N_3209);
nor U4166 (N_4166,N_3884,N_3674);
nand U4167 (N_4167,N_3766,N_3215);
or U4168 (N_4168,N_3774,N_3390);
nand U4169 (N_4169,N_3376,N_3083);
and U4170 (N_4170,N_3928,N_3907);
nand U4171 (N_4171,N_3715,N_3546);
nand U4172 (N_4172,N_3683,N_3232);
nor U4173 (N_4173,N_3216,N_3551);
or U4174 (N_4174,N_3583,N_3164);
xnor U4175 (N_4175,N_3702,N_3950);
and U4176 (N_4176,N_3076,N_3909);
nand U4177 (N_4177,N_3669,N_3482);
and U4178 (N_4178,N_3392,N_3910);
and U4179 (N_4179,N_3363,N_3960);
or U4180 (N_4180,N_3194,N_3948);
nor U4181 (N_4181,N_3951,N_3080);
and U4182 (N_4182,N_3084,N_3007);
nand U4183 (N_4183,N_3315,N_3129);
or U4184 (N_4184,N_3137,N_3170);
or U4185 (N_4185,N_3581,N_3586);
or U4186 (N_4186,N_3853,N_3637);
or U4187 (N_4187,N_3094,N_3144);
and U4188 (N_4188,N_3015,N_3625);
or U4189 (N_4189,N_3585,N_3266);
nand U4190 (N_4190,N_3069,N_3974);
or U4191 (N_4191,N_3848,N_3912);
and U4192 (N_4192,N_3204,N_3778);
nand U4193 (N_4193,N_3644,N_3606);
nand U4194 (N_4194,N_3291,N_3495);
or U4195 (N_4195,N_3797,N_3654);
and U4196 (N_4196,N_3785,N_3403);
nor U4197 (N_4197,N_3649,N_3515);
nand U4198 (N_4198,N_3492,N_3869);
or U4199 (N_4199,N_3588,N_3453);
xor U4200 (N_4200,N_3271,N_3434);
or U4201 (N_4201,N_3560,N_3494);
and U4202 (N_4202,N_3575,N_3541);
nor U4203 (N_4203,N_3885,N_3877);
nor U4204 (N_4204,N_3226,N_3187);
or U4205 (N_4205,N_3436,N_3919);
or U4206 (N_4206,N_3719,N_3052);
or U4207 (N_4207,N_3925,N_3373);
or U4208 (N_4208,N_3838,N_3282);
nand U4209 (N_4209,N_3758,N_3146);
nand U4210 (N_4210,N_3365,N_3534);
and U4211 (N_4211,N_3324,N_3806);
nor U4212 (N_4212,N_3776,N_3177);
and U4213 (N_4213,N_3255,N_3460);
and U4214 (N_4214,N_3718,N_3816);
and U4215 (N_4215,N_3481,N_3261);
nor U4216 (N_4216,N_3018,N_3378);
and U4217 (N_4217,N_3844,N_3283);
and U4218 (N_4218,N_3682,N_3891);
nor U4219 (N_4219,N_3597,N_3039);
or U4220 (N_4220,N_3990,N_3902);
nor U4221 (N_4221,N_3543,N_3973);
nand U4222 (N_4222,N_3220,N_3219);
and U4223 (N_4223,N_3182,N_3755);
nand U4224 (N_4224,N_3527,N_3211);
or U4225 (N_4225,N_3890,N_3576);
or U4226 (N_4226,N_3431,N_3622);
nor U4227 (N_4227,N_3500,N_3791);
and U4228 (N_4228,N_3268,N_3690);
or U4229 (N_4229,N_3713,N_3438);
and U4230 (N_4230,N_3173,N_3523);
or U4231 (N_4231,N_3807,N_3499);
and U4232 (N_4232,N_3553,N_3198);
or U4233 (N_4233,N_3265,N_3564);
or U4234 (N_4234,N_3593,N_3800);
nand U4235 (N_4235,N_3190,N_3850);
nand U4236 (N_4236,N_3075,N_3461);
nand U4237 (N_4237,N_3976,N_3013);
nor U4238 (N_4238,N_3180,N_3503);
nand U4239 (N_4239,N_3750,N_3865);
and U4240 (N_4240,N_3955,N_3328);
nor U4241 (N_4241,N_3380,N_3446);
nand U4242 (N_4242,N_3966,N_3478);
or U4243 (N_4243,N_3685,N_3741);
nor U4244 (N_4244,N_3159,N_3971);
nor U4245 (N_4245,N_3309,N_3531);
and U4246 (N_4246,N_3927,N_3108);
or U4247 (N_4247,N_3982,N_3104);
nand U4248 (N_4248,N_3587,N_3744);
nor U4249 (N_4249,N_3030,N_3428);
nand U4250 (N_4250,N_3203,N_3509);
and U4251 (N_4251,N_3071,N_3496);
nand U4252 (N_4252,N_3294,N_3828);
xor U4253 (N_4253,N_3525,N_3875);
and U4254 (N_4254,N_3545,N_3999);
nor U4255 (N_4255,N_3779,N_3632);
or U4256 (N_4256,N_3675,N_3657);
or U4257 (N_4257,N_3458,N_3161);
nand U4258 (N_4258,N_3947,N_3061);
and U4259 (N_4259,N_3922,N_3049);
nand U4260 (N_4260,N_3570,N_3914);
and U4261 (N_4261,N_3762,N_3168);
or U4262 (N_4262,N_3470,N_3439);
and U4263 (N_4263,N_3607,N_3724);
or U4264 (N_4264,N_3901,N_3402);
or U4265 (N_4265,N_3412,N_3491);
nor U4266 (N_4266,N_3464,N_3864);
nand U4267 (N_4267,N_3465,N_3342);
nand U4268 (N_4268,N_3957,N_3640);
nand U4269 (N_4269,N_3148,N_3245);
nor U4270 (N_4270,N_3089,N_3508);
nor U4271 (N_4271,N_3787,N_3705);
nor U4272 (N_4272,N_3736,N_3329);
or U4273 (N_4273,N_3630,N_3183);
or U4274 (N_4274,N_3374,N_3598);
nor U4275 (N_4275,N_3456,N_3643);
nand U4276 (N_4276,N_3253,N_3343);
nor U4277 (N_4277,N_3707,N_3401);
nor U4278 (N_4278,N_3332,N_3228);
nor U4279 (N_4279,N_3959,N_3610);
or U4280 (N_4280,N_3427,N_3680);
nand U4281 (N_4281,N_3526,N_3833);
nand U4282 (N_4282,N_3567,N_3449);
nor U4283 (N_4283,N_3742,N_3558);
nor U4284 (N_4284,N_3770,N_3372);
and U4285 (N_4285,N_3330,N_3388);
nor U4286 (N_4286,N_3921,N_3040);
nor U4287 (N_4287,N_3641,N_3444);
nor U4288 (N_4288,N_3609,N_3781);
nor U4289 (N_4289,N_3963,N_3000);
nor U4290 (N_4290,N_3367,N_3252);
nand U4291 (N_4291,N_3239,N_3227);
and U4292 (N_4292,N_3156,N_3498);
nor U4293 (N_4293,N_3440,N_3231);
nand U4294 (N_4294,N_3473,N_3426);
and U4295 (N_4295,N_3065,N_3312);
nand U4296 (N_4296,N_3443,N_3217);
nand U4297 (N_4297,N_3845,N_3655);
and U4298 (N_4298,N_3143,N_3229);
or U4299 (N_4299,N_3188,N_3991);
and U4300 (N_4300,N_3822,N_3289);
and U4301 (N_4301,N_3730,N_3174);
nand U4302 (N_4302,N_3769,N_3430);
and U4303 (N_4303,N_3623,N_3331);
nand U4304 (N_4304,N_3668,N_3832);
or U4305 (N_4305,N_3688,N_3236);
nor U4306 (N_4306,N_3340,N_3894);
nand U4307 (N_4307,N_3238,N_3528);
nand U4308 (N_4308,N_3695,N_3814);
or U4309 (N_4309,N_3524,N_3263);
nor U4310 (N_4310,N_3868,N_3856);
or U4311 (N_4311,N_3127,N_3036);
nand U4312 (N_4312,N_3497,N_3408);
or U4313 (N_4313,N_3748,N_3522);
or U4314 (N_4314,N_3782,N_3471);
and U4315 (N_4315,N_3099,N_3160);
and U4316 (N_4316,N_3485,N_3780);
nand U4317 (N_4317,N_3633,N_3087);
nand U4318 (N_4318,N_3516,N_3098);
nor U4319 (N_4319,N_3908,N_3670);
nor U4320 (N_4320,N_3450,N_3212);
or U4321 (N_4321,N_3337,N_3572);
nor U4322 (N_4322,N_3624,N_3067);
nor U4323 (N_4323,N_3979,N_3870);
or U4324 (N_4324,N_3163,N_3191);
and U4325 (N_4325,N_3977,N_3574);
and U4326 (N_4326,N_3126,N_3279);
nor U4327 (N_4327,N_3202,N_3359);
nand U4328 (N_4328,N_3442,N_3467);
or U4329 (N_4329,N_3965,N_3519);
or U4330 (N_4330,N_3945,N_3817);
and U4331 (N_4331,N_3414,N_3956);
nand U4332 (N_4332,N_3119,N_3276);
or U4333 (N_4333,N_3876,N_3233);
and U4334 (N_4334,N_3424,N_3260);
and U4335 (N_4335,N_3091,N_3843);
or U4336 (N_4336,N_3407,N_3867);
nor U4337 (N_4337,N_3579,N_3760);
and U4338 (N_4338,N_3726,N_3421);
and U4339 (N_4339,N_3504,N_3109);
nand U4340 (N_4340,N_3131,N_3100);
or U4341 (N_4341,N_3051,N_3079);
nand U4342 (N_4342,N_3122,N_3062);
or U4343 (N_4343,N_3936,N_3539);
and U4344 (N_4344,N_3542,N_3394);
nand U4345 (N_4345,N_3946,N_3533);
and U4346 (N_4346,N_3830,N_3888);
and U4347 (N_4347,N_3513,N_3677);
or U4348 (N_4348,N_3701,N_3166);
nor U4349 (N_4349,N_3898,N_3272);
or U4350 (N_4350,N_3479,N_3771);
nor U4351 (N_4351,N_3139,N_3299);
and U4352 (N_4352,N_3241,N_3317);
or U4353 (N_4353,N_3234,N_3562);
or U4354 (N_4354,N_3468,N_3929);
nor U4355 (N_4355,N_3114,N_3834);
nand U4356 (N_4356,N_3186,N_3185);
nand U4357 (N_4357,N_3396,N_3278);
and U4358 (N_4358,N_3804,N_3339);
nand U4359 (N_4359,N_3854,N_3386);
nand U4360 (N_4360,N_3917,N_3325);
and U4361 (N_4361,N_3082,N_3286);
nor U4362 (N_4362,N_3994,N_3037);
nand U4363 (N_4363,N_3501,N_3162);
or U4364 (N_4364,N_3296,N_3149);
or U4365 (N_4365,N_3795,N_3323);
nor U4366 (N_4366,N_3406,N_3995);
nor U4367 (N_4367,N_3070,N_3767);
nand U4368 (N_4368,N_3855,N_3967);
and U4369 (N_4369,N_3264,N_3258);
or U4370 (N_4370,N_3916,N_3647);
or U4371 (N_4371,N_3136,N_3404);
nand U4372 (N_4372,N_3221,N_3997);
and U4373 (N_4373,N_3798,N_3873);
nand U4374 (N_4374,N_3476,N_3356);
nor U4375 (N_4375,N_3043,N_3413);
nor U4376 (N_4376,N_3642,N_3369);
nand U4377 (N_4377,N_3801,N_3338);
nor U4378 (N_4378,N_3383,N_3904);
and U4379 (N_4379,N_3395,N_3860);
and U4380 (N_4380,N_3019,N_3699);
or U4381 (N_4381,N_3708,N_3293);
nor U4382 (N_4382,N_3536,N_3520);
and U4383 (N_4383,N_3836,N_3998);
and U4384 (N_4384,N_3565,N_3638);
and U4385 (N_4385,N_3003,N_3661);
and U4386 (N_4386,N_3980,N_3321);
nor U4387 (N_4387,N_3698,N_3057);
or U4388 (N_4388,N_3629,N_3262);
and U4389 (N_4389,N_3237,N_3549);
and U4390 (N_4390,N_3969,N_3987);
nand U4391 (N_4391,N_3595,N_3022);
and U4392 (N_4392,N_3616,N_3819);
or U4393 (N_4393,N_3032,N_3179);
nand U4394 (N_4394,N_3731,N_3849);
and U4395 (N_4395,N_3732,N_3172);
and U4396 (N_4396,N_3447,N_3892);
or U4397 (N_4397,N_3862,N_3134);
or U4398 (N_4398,N_3008,N_3086);
and U4399 (N_4399,N_3242,N_3619);
nor U4400 (N_4400,N_3038,N_3938);
nand U4401 (N_4401,N_3147,N_3105);
nand U4402 (N_4402,N_3571,N_3489);
nand U4403 (N_4403,N_3887,N_3577);
nand U4404 (N_4404,N_3142,N_3152);
or U4405 (N_4405,N_3861,N_3254);
or U4406 (N_4406,N_3846,N_3989);
or U4407 (N_4407,N_3752,N_3697);
nand U4408 (N_4408,N_3288,N_3895);
or U4409 (N_4409,N_3858,N_3820);
or U4410 (N_4410,N_3319,N_3789);
and U4411 (N_4411,N_3631,N_3635);
or U4412 (N_4412,N_3578,N_3620);
and U4413 (N_4413,N_3196,N_3662);
nor U4414 (N_4414,N_3247,N_3102);
xor U4415 (N_4415,N_3341,N_3107);
and U4416 (N_4416,N_3002,N_3322);
nand U4417 (N_4417,N_3116,N_3193);
and U4418 (N_4418,N_3880,N_3437);
nand U4419 (N_4419,N_3988,N_3694);
nor U4420 (N_4420,N_3125,N_3926);
or U4421 (N_4421,N_3612,N_3671);
nand U4422 (N_4422,N_3429,N_3521);
nand U4423 (N_4423,N_3115,N_3297);
or U4424 (N_4424,N_3535,N_3355);
or U4425 (N_4425,N_3269,N_3911);
xnor U4426 (N_4426,N_3878,N_3056);
and U4427 (N_4427,N_3879,N_3457);
or U4428 (N_4428,N_3506,N_3658);
nand U4429 (N_4429,N_3993,N_3273);
or U4430 (N_4430,N_3881,N_3078);
or U4431 (N_4431,N_3488,N_3393);
or U4432 (N_4432,N_3184,N_3213);
or U4433 (N_4433,N_3602,N_3484);
nand U4434 (N_4434,N_3899,N_3827);
and U4435 (N_4435,N_3826,N_3725);
nor U4436 (N_4436,N_3335,N_3064);
or U4437 (N_4437,N_3992,N_3537);
xor U4438 (N_4438,N_3368,N_3001);
nor U4439 (N_4439,N_3249,N_3410);
nor U4440 (N_4440,N_3044,N_3563);
and U4441 (N_4441,N_3101,N_3195);
nand U4442 (N_4442,N_3224,N_3110);
nand U4443 (N_4443,N_3222,N_3206);
nor U4444 (N_4444,N_3753,N_3016);
nand U4445 (N_4445,N_3842,N_3648);
or U4446 (N_4446,N_3391,N_3246);
nor U4447 (N_4447,N_3028,N_3716);
nor U4448 (N_4448,N_3469,N_3544);
nor U4449 (N_4449,N_3600,N_3920);
and U4450 (N_4450,N_3382,N_3205);
and U4451 (N_4451,N_3361,N_3686);
nand U4452 (N_4452,N_3942,N_3840);
or U4453 (N_4453,N_3737,N_3090);
nor U4454 (N_4454,N_3932,N_3130);
nor U4455 (N_4455,N_3371,N_3487);
nand U4456 (N_4456,N_3617,N_3964);
nand U4457 (N_4457,N_3480,N_3505);
or U4458 (N_4458,N_3199,N_3915);
nand U4459 (N_4459,N_3627,N_3124);
nor U4460 (N_4460,N_3230,N_3275);
and U4461 (N_4461,N_3512,N_3788);
nor U4462 (N_4462,N_3815,N_3012);
or U4463 (N_4463,N_3490,N_3225);
nand U4464 (N_4464,N_3189,N_3582);
nand U4465 (N_4465,N_3538,N_3831);
nor U4466 (N_4466,N_3042,N_3923);
nand U4467 (N_4467,N_3596,N_3113);
nor U4468 (N_4468,N_3871,N_3389);
or U4469 (N_4469,N_3611,N_3599);
nand U4470 (N_4470,N_3605,N_3757);
nand U4471 (N_4471,N_3761,N_3970);
and U4472 (N_4472,N_3930,N_3984);
nand U4473 (N_4473,N_3681,N_3121);
nand U4474 (N_4474,N_3475,N_3913);
nor U4475 (N_4475,N_3024,N_3357);
nand U4476 (N_4476,N_3818,N_3300);
nand U4477 (N_4477,N_3004,N_3298);
and U4478 (N_4478,N_3452,N_3794);
nand U4479 (N_4479,N_3653,N_3722);
or U4480 (N_4480,N_3416,N_3240);
xor U4481 (N_4481,N_3783,N_3274);
nor U4482 (N_4482,N_3017,N_3958);
and U4483 (N_4483,N_3153,N_3063);
xnor U4484 (N_4484,N_3768,N_3303);
nand U4485 (N_4485,N_3454,N_3045);
nor U4486 (N_4486,N_3223,N_3756);
nand U4487 (N_4487,N_3983,N_3308);
or U4488 (N_4488,N_3111,N_3700);
nor U4489 (N_4489,N_3055,N_3326);
nor U4490 (N_4490,N_3400,N_3169);
nor U4491 (N_4491,N_3103,N_3033);
nand U4492 (N_4492,N_3594,N_3940);
and U4493 (N_4493,N_3422,N_3790);
nand U4494 (N_4494,N_3740,N_3201);
or U4495 (N_4495,N_3123,N_3673);
and U4496 (N_4496,N_3953,N_3360);
and U4497 (N_4497,N_3477,N_3302);
nor U4498 (N_4498,N_3939,N_3918);
nor U4499 (N_4499,N_3935,N_3978);
nand U4500 (N_4500,N_3999,N_3265);
and U4501 (N_4501,N_3162,N_3852);
and U4502 (N_4502,N_3905,N_3964);
or U4503 (N_4503,N_3169,N_3048);
or U4504 (N_4504,N_3776,N_3048);
nor U4505 (N_4505,N_3960,N_3062);
nor U4506 (N_4506,N_3159,N_3396);
or U4507 (N_4507,N_3288,N_3470);
or U4508 (N_4508,N_3561,N_3611);
nor U4509 (N_4509,N_3196,N_3149);
nor U4510 (N_4510,N_3370,N_3226);
or U4511 (N_4511,N_3210,N_3925);
or U4512 (N_4512,N_3321,N_3108);
nor U4513 (N_4513,N_3860,N_3389);
xnor U4514 (N_4514,N_3647,N_3620);
nand U4515 (N_4515,N_3821,N_3454);
nor U4516 (N_4516,N_3501,N_3847);
nand U4517 (N_4517,N_3774,N_3736);
and U4518 (N_4518,N_3265,N_3064);
nor U4519 (N_4519,N_3898,N_3478);
nor U4520 (N_4520,N_3847,N_3214);
and U4521 (N_4521,N_3678,N_3480);
nor U4522 (N_4522,N_3486,N_3585);
or U4523 (N_4523,N_3812,N_3235);
nand U4524 (N_4524,N_3296,N_3644);
or U4525 (N_4525,N_3750,N_3287);
nand U4526 (N_4526,N_3045,N_3583);
nand U4527 (N_4527,N_3665,N_3013);
and U4528 (N_4528,N_3108,N_3672);
nor U4529 (N_4529,N_3334,N_3235);
and U4530 (N_4530,N_3667,N_3017);
nor U4531 (N_4531,N_3443,N_3290);
and U4532 (N_4532,N_3925,N_3775);
nand U4533 (N_4533,N_3695,N_3714);
or U4534 (N_4534,N_3577,N_3672);
or U4535 (N_4535,N_3897,N_3726);
and U4536 (N_4536,N_3347,N_3973);
nor U4537 (N_4537,N_3255,N_3944);
and U4538 (N_4538,N_3160,N_3045);
nand U4539 (N_4539,N_3196,N_3458);
or U4540 (N_4540,N_3926,N_3472);
or U4541 (N_4541,N_3736,N_3355);
nand U4542 (N_4542,N_3776,N_3215);
nand U4543 (N_4543,N_3689,N_3663);
and U4544 (N_4544,N_3062,N_3569);
nand U4545 (N_4545,N_3770,N_3667);
nor U4546 (N_4546,N_3058,N_3752);
and U4547 (N_4547,N_3915,N_3108);
or U4548 (N_4548,N_3106,N_3244);
and U4549 (N_4549,N_3068,N_3881);
nor U4550 (N_4550,N_3384,N_3551);
and U4551 (N_4551,N_3975,N_3530);
and U4552 (N_4552,N_3346,N_3928);
nor U4553 (N_4553,N_3674,N_3438);
and U4554 (N_4554,N_3117,N_3010);
nor U4555 (N_4555,N_3700,N_3903);
nand U4556 (N_4556,N_3455,N_3231);
or U4557 (N_4557,N_3931,N_3146);
and U4558 (N_4558,N_3762,N_3450);
and U4559 (N_4559,N_3197,N_3923);
nor U4560 (N_4560,N_3091,N_3839);
nand U4561 (N_4561,N_3169,N_3745);
nand U4562 (N_4562,N_3005,N_3530);
or U4563 (N_4563,N_3017,N_3815);
nor U4564 (N_4564,N_3117,N_3356);
or U4565 (N_4565,N_3075,N_3608);
xor U4566 (N_4566,N_3597,N_3444);
and U4567 (N_4567,N_3064,N_3565);
and U4568 (N_4568,N_3626,N_3491);
nor U4569 (N_4569,N_3086,N_3781);
nand U4570 (N_4570,N_3152,N_3920);
or U4571 (N_4571,N_3779,N_3352);
nor U4572 (N_4572,N_3290,N_3763);
and U4573 (N_4573,N_3301,N_3013);
xnor U4574 (N_4574,N_3209,N_3578);
nand U4575 (N_4575,N_3874,N_3484);
nand U4576 (N_4576,N_3810,N_3603);
nand U4577 (N_4577,N_3755,N_3850);
nor U4578 (N_4578,N_3585,N_3973);
or U4579 (N_4579,N_3478,N_3551);
nand U4580 (N_4580,N_3238,N_3530);
and U4581 (N_4581,N_3259,N_3191);
nand U4582 (N_4582,N_3911,N_3116);
and U4583 (N_4583,N_3865,N_3973);
nand U4584 (N_4584,N_3658,N_3875);
and U4585 (N_4585,N_3295,N_3392);
nor U4586 (N_4586,N_3097,N_3242);
and U4587 (N_4587,N_3592,N_3295);
and U4588 (N_4588,N_3253,N_3546);
and U4589 (N_4589,N_3799,N_3570);
nand U4590 (N_4590,N_3733,N_3298);
or U4591 (N_4591,N_3147,N_3515);
and U4592 (N_4592,N_3005,N_3087);
and U4593 (N_4593,N_3463,N_3214);
nand U4594 (N_4594,N_3045,N_3242);
or U4595 (N_4595,N_3925,N_3353);
nand U4596 (N_4596,N_3451,N_3947);
xnor U4597 (N_4597,N_3056,N_3172);
and U4598 (N_4598,N_3944,N_3212);
or U4599 (N_4599,N_3132,N_3334);
nor U4600 (N_4600,N_3517,N_3349);
nand U4601 (N_4601,N_3200,N_3166);
nor U4602 (N_4602,N_3128,N_3668);
or U4603 (N_4603,N_3500,N_3619);
and U4604 (N_4604,N_3545,N_3730);
or U4605 (N_4605,N_3165,N_3561);
or U4606 (N_4606,N_3165,N_3404);
and U4607 (N_4607,N_3027,N_3506);
nor U4608 (N_4608,N_3910,N_3646);
nor U4609 (N_4609,N_3363,N_3479);
and U4610 (N_4610,N_3219,N_3218);
and U4611 (N_4611,N_3657,N_3515);
nand U4612 (N_4612,N_3706,N_3001);
nor U4613 (N_4613,N_3026,N_3492);
nand U4614 (N_4614,N_3672,N_3860);
nand U4615 (N_4615,N_3270,N_3013);
and U4616 (N_4616,N_3934,N_3632);
and U4617 (N_4617,N_3338,N_3600);
or U4618 (N_4618,N_3059,N_3190);
and U4619 (N_4619,N_3890,N_3427);
or U4620 (N_4620,N_3541,N_3237);
and U4621 (N_4621,N_3306,N_3409);
nor U4622 (N_4622,N_3443,N_3576);
nand U4623 (N_4623,N_3945,N_3856);
nand U4624 (N_4624,N_3488,N_3495);
and U4625 (N_4625,N_3013,N_3589);
and U4626 (N_4626,N_3294,N_3650);
and U4627 (N_4627,N_3350,N_3063);
or U4628 (N_4628,N_3339,N_3607);
and U4629 (N_4629,N_3578,N_3604);
nand U4630 (N_4630,N_3293,N_3913);
nand U4631 (N_4631,N_3449,N_3155);
or U4632 (N_4632,N_3829,N_3510);
nor U4633 (N_4633,N_3661,N_3472);
or U4634 (N_4634,N_3165,N_3305);
and U4635 (N_4635,N_3457,N_3667);
nand U4636 (N_4636,N_3992,N_3627);
and U4637 (N_4637,N_3001,N_3566);
and U4638 (N_4638,N_3276,N_3856);
nor U4639 (N_4639,N_3202,N_3875);
and U4640 (N_4640,N_3793,N_3535);
xor U4641 (N_4641,N_3819,N_3065);
or U4642 (N_4642,N_3965,N_3055);
or U4643 (N_4643,N_3543,N_3394);
or U4644 (N_4644,N_3365,N_3470);
or U4645 (N_4645,N_3306,N_3931);
nand U4646 (N_4646,N_3113,N_3916);
and U4647 (N_4647,N_3929,N_3452);
nor U4648 (N_4648,N_3966,N_3495);
or U4649 (N_4649,N_3159,N_3935);
nand U4650 (N_4650,N_3526,N_3186);
nor U4651 (N_4651,N_3970,N_3012);
nand U4652 (N_4652,N_3210,N_3675);
and U4653 (N_4653,N_3446,N_3563);
or U4654 (N_4654,N_3284,N_3963);
and U4655 (N_4655,N_3871,N_3504);
and U4656 (N_4656,N_3461,N_3809);
nand U4657 (N_4657,N_3125,N_3719);
and U4658 (N_4658,N_3094,N_3225);
nor U4659 (N_4659,N_3505,N_3044);
or U4660 (N_4660,N_3134,N_3691);
and U4661 (N_4661,N_3814,N_3591);
nor U4662 (N_4662,N_3470,N_3876);
or U4663 (N_4663,N_3675,N_3198);
and U4664 (N_4664,N_3367,N_3862);
nand U4665 (N_4665,N_3866,N_3493);
or U4666 (N_4666,N_3343,N_3557);
or U4667 (N_4667,N_3831,N_3542);
nand U4668 (N_4668,N_3043,N_3845);
or U4669 (N_4669,N_3648,N_3165);
or U4670 (N_4670,N_3298,N_3620);
or U4671 (N_4671,N_3151,N_3033);
or U4672 (N_4672,N_3794,N_3031);
nor U4673 (N_4673,N_3221,N_3424);
nand U4674 (N_4674,N_3553,N_3106);
nor U4675 (N_4675,N_3440,N_3447);
or U4676 (N_4676,N_3039,N_3433);
and U4677 (N_4677,N_3872,N_3851);
or U4678 (N_4678,N_3484,N_3549);
or U4679 (N_4679,N_3828,N_3706);
or U4680 (N_4680,N_3267,N_3741);
and U4681 (N_4681,N_3530,N_3875);
nor U4682 (N_4682,N_3146,N_3601);
nor U4683 (N_4683,N_3092,N_3056);
nand U4684 (N_4684,N_3658,N_3142);
or U4685 (N_4685,N_3450,N_3097);
nor U4686 (N_4686,N_3830,N_3111);
and U4687 (N_4687,N_3309,N_3439);
nand U4688 (N_4688,N_3236,N_3223);
and U4689 (N_4689,N_3519,N_3998);
and U4690 (N_4690,N_3208,N_3895);
nand U4691 (N_4691,N_3408,N_3327);
and U4692 (N_4692,N_3957,N_3863);
nand U4693 (N_4693,N_3349,N_3728);
and U4694 (N_4694,N_3600,N_3515);
nand U4695 (N_4695,N_3679,N_3023);
nand U4696 (N_4696,N_3090,N_3153);
nor U4697 (N_4697,N_3355,N_3082);
nor U4698 (N_4698,N_3416,N_3554);
nor U4699 (N_4699,N_3747,N_3779);
or U4700 (N_4700,N_3208,N_3802);
nor U4701 (N_4701,N_3796,N_3817);
and U4702 (N_4702,N_3260,N_3473);
nand U4703 (N_4703,N_3891,N_3442);
nand U4704 (N_4704,N_3295,N_3518);
nand U4705 (N_4705,N_3992,N_3717);
and U4706 (N_4706,N_3082,N_3894);
or U4707 (N_4707,N_3645,N_3186);
nand U4708 (N_4708,N_3098,N_3274);
nand U4709 (N_4709,N_3494,N_3183);
xnor U4710 (N_4710,N_3307,N_3763);
or U4711 (N_4711,N_3107,N_3431);
or U4712 (N_4712,N_3537,N_3863);
nand U4713 (N_4713,N_3722,N_3878);
and U4714 (N_4714,N_3876,N_3914);
and U4715 (N_4715,N_3727,N_3639);
nor U4716 (N_4716,N_3578,N_3133);
nor U4717 (N_4717,N_3885,N_3685);
and U4718 (N_4718,N_3598,N_3757);
nor U4719 (N_4719,N_3457,N_3939);
nor U4720 (N_4720,N_3511,N_3212);
or U4721 (N_4721,N_3884,N_3185);
nor U4722 (N_4722,N_3794,N_3617);
or U4723 (N_4723,N_3146,N_3219);
nor U4724 (N_4724,N_3464,N_3009);
and U4725 (N_4725,N_3152,N_3455);
or U4726 (N_4726,N_3033,N_3216);
or U4727 (N_4727,N_3007,N_3265);
and U4728 (N_4728,N_3726,N_3144);
and U4729 (N_4729,N_3600,N_3304);
nand U4730 (N_4730,N_3874,N_3469);
and U4731 (N_4731,N_3624,N_3524);
or U4732 (N_4732,N_3857,N_3847);
and U4733 (N_4733,N_3181,N_3508);
nor U4734 (N_4734,N_3785,N_3774);
and U4735 (N_4735,N_3072,N_3642);
nor U4736 (N_4736,N_3380,N_3415);
or U4737 (N_4737,N_3395,N_3992);
nand U4738 (N_4738,N_3026,N_3699);
or U4739 (N_4739,N_3845,N_3246);
nor U4740 (N_4740,N_3392,N_3239);
and U4741 (N_4741,N_3628,N_3563);
nor U4742 (N_4742,N_3357,N_3897);
nand U4743 (N_4743,N_3059,N_3445);
or U4744 (N_4744,N_3524,N_3028);
and U4745 (N_4745,N_3759,N_3736);
and U4746 (N_4746,N_3732,N_3316);
nor U4747 (N_4747,N_3085,N_3239);
nand U4748 (N_4748,N_3422,N_3509);
nand U4749 (N_4749,N_3531,N_3114);
or U4750 (N_4750,N_3295,N_3566);
nand U4751 (N_4751,N_3203,N_3137);
and U4752 (N_4752,N_3314,N_3471);
or U4753 (N_4753,N_3742,N_3214);
or U4754 (N_4754,N_3477,N_3897);
or U4755 (N_4755,N_3816,N_3290);
or U4756 (N_4756,N_3154,N_3638);
nor U4757 (N_4757,N_3357,N_3336);
and U4758 (N_4758,N_3468,N_3852);
and U4759 (N_4759,N_3052,N_3695);
nor U4760 (N_4760,N_3904,N_3013);
nand U4761 (N_4761,N_3474,N_3061);
or U4762 (N_4762,N_3256,N_3478);
or U4763 (N_4763,N_3521,N_3060);
nor U4764 (N_4764,N_3735,N_3308);
and U4765 (N_4765,N_3632,N_3715);
nand U4766 (N_4766,N_3974,N_3123);
and U4767 (N_4767,N_3831,N_3485);
or U4768 (N_4768,N_3636,N_3476);
and U4769 (N_4769,N_3721,N_3558);
nor U4770 (N_4770,N_3670,N_3482);
or U4771 (N_4771,N_3055,N_3778);
and U4772 (N_4772,N_3250,N_3137);
nand U4773 (N_4773,N_3129,N_3460);
or U4774 (N_4774,N_3678,N_3779);
and U4775 (N_4775,N_3651,N_3251);
and U4776 (N_4776,N_3340,N_3367);
nand U4777 (N_4777,N_3758,N_3047);
and U4778 (N_4778,N_3298,N_3303);
and U4779 (N_4779,N_3708,N_3376);
and U4780 (N_4780,N_3616,N_3253);
nand U4781 (N_4781,N_3252,N_3187);
or U4782 (N_4782,N_3423,N_3826);
or U4783 (N_4783,N_3145,N_3316);
nor U4784 (N_4784,N_3337,N_3534);
nor U4785 (N_4785,N_3161,N_3762);
nor U4786 (N_4786,N_3988,N_3434);
nor U4787 (N_4787,N_3479,N_3844);
and U4788 (N_4788,N_3508,N_3021);
nand U4789 (N_4789,N_3232,N_3195);
nor U4790 (N_4790,N_3709,N_3179);
or U4791 (N_4791,N_3403,N_3457);
or U4792 (N_4792,N_3280,N_3420);
nor U4793 (N_4793,N_3303,N_3160);
and U4794 (N_4794,N_3058,N_3732);
nand U4795 (N_4795,N_3264,N_3907);
and U4796 (N_4796,N_3777,N_3564);
or U4797 (N_4797,N_3198,N_3427);
nand U4798 (N_4798,N_3150,N_3570);
nand U4799 (N_4799,N_3869,N_3557);
nand U4800 (N_4800,N_3976,N_3102);
nor U4801 (N_4801,N_3755,N_3878);
and U4802 (N_4802,N_3286,N_3383);
nand U4803 (N_4803,N_3521,N_3927);
or U4804 (N_4804,N_3806,N_3457);
nor U4805 (N_4805,N_3524,N_3654);
nand U4806 (N_4806,N_3607,N_3857);
or U4807 (N_4807,N_3370,N_3467);
and U4808 (N_4808,N_3344,N_3097);
or U4809 (N_4809,N_3758,N_3409);
and U4810 (N_4810,N_3421,N_3827);
nand U4811 (N_4811,N_3021,N_3961);
nor U4812 (N_4812,N_3778,N_3192);
and U4813 (N_4813,N_3001,N_3079);
or U4814 (N_4814,N_3459,N_3593);
nor U4815 (N_4815,N_3599,N_3816);
nor U4816 (N_4816,N_3330,N_3304);
and U4817 (N_4817,N_3310,N_3286);
and U4818 (N_4818,N_3780,N_3670);
or U4819 (N_4819,N_3630,N_3485);
nand U4820 (N_4820,N_3664,N_3229);
nand U4821 (N_4821,N_3132,N_3781);
nor U4822 (N_4822,N_3712,N_3475);
nand U4823 (N_4823,N_3797,N_3548);
or U4824 (N_4824,N_3635,N_3536);
nand U4825 (N_4825,N_3186,N_3557);
or U4826 (N_4826,N_3229,N_3699);
nor U4827 (N_4827,N_3592,N_3624);
or U4828 (N_4828,N_3394,N_3941);
nor U4829 (N_4829,N_3297,N_3914);
and U4830 (N_4830,N_3520,N_3434);
and U4831 (N_4831,N_3632,N_3230);
or U4832 (N_4832,N_3637,N_3059);
and U4833 (N_4833,N_3117,N_3349);
or U4834 (N_4834,N_3321,N_3243);
or U4835 (N_4835,N_3694,N_3073);
nor U4836 (N_4836,N_3076,N_3878);
or U4837 (N_4837,N_3177,N_3310);
and U4838 (N_4838,N_3408,N_3037);
nand U4839 (N_4839,N_3629,N_3515);
nor U4840 (N_4840,N_3033,N_3611);
or U4841 (N_4841,N_3663,N_3876);
nand U4842 (N_4842,N_3881,N_3439);
and U4843 (N_4843,N_3755,N_3453);
nand U4844 (N_4844,N_3166,N_3673);
or U4845 (N_4845,N_3718,N_3263);
nand U4846 (N_4846,N_3022,N_3062);
nor U4847 (N_4847,N_3181,N_3954);
nor U4848 (N_4848,N_3317,N_3044);
and U4849 (N_4849,N_3032,N_3888);
nor U4850 (N_4850,N_3731,N_3983);
and U4851 (N_4851,N_3339,N_3380);
or U4852 (N_4852,N_3115,N_3259);
nor U4853 (N_4853,N_3570,N_3346);
nand U4854 (N_4854,N_3029,N_3938);
nand U4855 (N_4855,N_3192,N_3540);
or U4856 (N_4856,N_3104,N_3881);
nor U4857 (N_4857,N_3000,N_3781);
or U4858 (N_4858,N_3230,N_3475);
or U4859 (N_4859,N_3345,N_3571);
nand U4860 (N_4860,N_3846,N_3461);
or U4861 (N_4861,N_3848,N_3651);
nor U4862 (N_4862,N_3094,N_3017);
nor U4863 (N_4863,N_3969,N_3139);
nand U4864 (N_4864,N_3467,N_3883);
nand U4865 (N_4865,N_3135,N_3492);
nor U4866 (N_4866,N_3447,N_3361);
nand U4867 (N_4867,N_3701,N_3533);
or U4868 (N_4868,N_3495,N_3443);
and U4869 (N_4869,N_3715,N_3761);
nor U4870 (N_4870,N_3818,N_3841);
nor U4871 (N_4871,N_3737,N_3742);
nor U4872 (N_4872,N_3158,N_3688);
and U4873 (N_4873,N_3806,N_3420);
nor U4874 (N_4874,N_3574,N_3948);
nor U4875 (N_4875,N_3938,N_3638);
or U4876 (N_4876,N_3960,N_3408);
and U4877 (N_4877,N_3515,N_3725);
nor U4878 (N_4878,N_3105,N_3573);
and U4879 (N_4879,N_3282,N_3923);
and U4880 (N_4880,N_3963,N_3588);
and U4881 (N_4881,N_3711,N_3773);
and U4882 (N_4882,N_3364,N_3089);
or U4883 (N_4883,N_3801,N_3282);
nand U4884 (N_4884,N_3875,N_3825);
and U4885 (N_4885,N_3226,N_3335);
nand U4886 (N_4886,N_3424,N_3374);
nor U4887 (N_4887,N_3394,N_3624);
and U4888 (N_4888,N_3427,N_3600);
nor U4889 (N_4889,N_3562,N_3333);
nand U4890 (N_4890,N_3356,N_3612);
and U4891 (N_4891,N_3110,N_3069);
nand U4892 (N_4892,N_3846,N_3632);
nand U4893 (N_4893,N_3997,N_3433);
nor U4894 (N_4894,N_3155,N_3612);
or U4895 (N_4895,N_3818,N_3705);
or U4896 (N_4896,N_3271,N_3192);
or U4897 (N_4897,N_3706,N_3743);
and U4898 (N_4898,N_3111,N_3100);
nor U4899 (N_4899,N_3912,N_3599);
or U4900 (N_4900,N_3532,N_3081);
nand U4901 (N_4901,N_3190,N_3259);
and U4902 (N_4902,N_3867,N_3269);
nor U4903 (N_4903,N_3613,N_3867);
nor U4904 (N_4904,N_3374,N_3860);
nand U4905 (N_4905,N_3116,N_3432);
nor U4906 (N_4906,N_3780,N_3528);
or U4907 (N_4907,N_3486,N_3129);
xor U4908 (N_4908,N_3553,N_3527);
nand U4909 (N_4909,N_3075,N_3498);
nand U4910 (N_4910,N_3196,N_3250);
or U4911 (N_4911,N_3643,N_3642);
nor U4912 (N_4912,N_3524,N_3658);
nand U4913 (N_4913,N_3134,N_3221);
nand U4914 (N_4914,N_3680,N_3031);
nor U4915 (N_4915,N_3616,N_3679);
nor U4916 (N_4916,N_3349,N_3682);
nand U4917 (N_4917,N_3864,N_3456);
nand U4918 (N_4918,N_3380,N_3091);
nor U4919 (N_4919,N_3053,N_3948);
nand U4920 (N_4920,N_3978,N_3612);
or U4921 (N_4921,N_3102,N_3970);
nor U4922 (N_4922,N_3341,N_3456);
and U4923 (N_4923,N_3697,N_3772);
nor U4924 (N_4924,N_3869,N_3901);
or U4925 (N_4925,N_3324,N_3868);
nor U4926 (N_4926,N_3507,N_3229);
nand U4927 (N_4927,N_3782,N_3701);
and U4928 (N_4928,N_3161,N_3375);
and U4929 (N_4929,N_3266,N_3773);
or U4930 (N_4930,N_3870,N_3738);
or U4931 (N_4931,N_3368,N_3410);
or U4932 (N_4932,N_3520,N_3870);
nand U4933 (N_4933,N_3730,N_3533);
or U4934 (N_4934,N_3600,N_3756);
nand U4935 (N_4935,N_3688,N_3523);
nor U4936 (N_4936,N_3688,N_3208);
nand U4937 (N_4937,N_3507,N_3323);
nor U4938 (N_4938,N_3629,N_3738);
nand U4939 (N_4939,N_3738,N_3700);
nor U4940 (N_4940,N_3599,N_3329);
nand U4941 (N_4941,N_3015,N_3369);
nand U4942 (N_4942,N_3127,N_3075);
and U4943 (N_4943,N_3863,N_3522);
and U4944 (N_4944,N_3793,N_3000);
or U4945 (N_4945,N_3531,N_3298);
nor U4946 (N_4946,N_3562,N_3496);
nand U4947 (N_4947,N_3952,N_3144);
and U4948 (N_4948,N_3600,N_3360);
xor U4949 (N_4949,N_3297,N_3493);
and U4950 (N_4950,N_3475,N_3510);
nor U4951 (N_4951,N_3845,N_3034);
nand U4952 (N_4952,N_3233,N_3266);
nor U4953 (N_4953,N_3294,N_3551);
nand U4954 (N_4954,N_3371,N_3657);
or U4955 (N_4955,N_3400,N_3578);
or U4956 (N_4956,N_3184,N_3215);
nand U4957 (N_4957,N_3177,N_3259);
or U4958 (N_4958,N_3317,N_3285);
nor U4959 (N_4959,N_3684,N_3362);
and U4960 (N_4960,N_3097,N_3718);
nand U4961 (N_4961,N_3103,N_3426);
and U4962 (N_4962,N_3255,N_3147);
nand U4963 (N_4963,N_3351,N_3208);
nor U4964 (N_4964,N_3060,N_3226);
nor U4965 (N_4965,N_3731,N_3443);
nor U4966 (N_4966,N_3513,N_3171);
or U4967 (N_4967,N_3057,N_3070);
nand U4968 (N_4968,N_3341,N_3997);
or U4969 (N_4969,N_3509,N_3837);
nand U4970 (N_4970,N_3875,N_3731);
nor U4971 (N_4971,N_3342,N_3751);
nor U4972 (N_4972,N_3019,N_3908);
nand U4973 (N_4973,N_3928,N_3288);
xor U4974 (N_4974,N_3637,N_3035);
nand U4975 (N_4975,N_3393,N_3384);
nor U4976 (N_4976,N_3458,N_3817);
nor U4977 (N_4977,N_3028,N_3163);
nor U4978 (N_4978,N_3196,N_3962);
nor U4979 (N_4979,N_3203,N_3140);
nor U4980 (N_4980,N_3314,N_3345);
and U4981 (N_4981,N_3349,N_3318);
and U4982 (N_4982,N_3360,N_3918);
nor U4983 (N_4983,N_3831,N_3615);
nor U4984 (N_4984,N_3235,N_3234);
nor U4985 (N_4985,N_3890,N_3345);
or U4986 (N_4986,N_3611,N_3558);
nor U4987 (N_4987,N_3078,N_3194);
nor U4988 (N_4988,N_3442,N_3289);
nand U4989 (N_4989,N_3933,N_3024);
and U4990 (N_4990,N_3683,N_3865);
and U4991 (N_4991,N_3529,N_3507);
nor U4992 (N_4992,N_3159,N_3150);
nand U4993 (N_4993,N_3691,N_3415);
nor U4994 (N_4994,N_3556,N_3270);
nand U4995 (N_4995,N_3051,N_3698);
nand U4996 (N_4996,N_3396,N_3097);
nor U4997 (N_4997,N_3037,N_3729);
and U4998 (N_4998,N_3978,N_3548);
or U4999 (N_4999,N_3840,N_3004);
nand U5000 (N_5000,N_4678,N_4153);
and U5001 (N_5001,N_4454,N_4638);
nand U5002 (N_5002,N_4098,N_4789);
and U5003 (N_5003,N_4597,N_4489);
and U5004 (N_5004,N_4302,N_4307);
or U5005 (N_5005,N_4719,N_4121);
nor U5006 (N_5006,N_4372,N_4116);
nand U5007 (N_5007,N_4024,N_4931);
nor U5008 (N_5008,N_4217,N_4775);
and U5009 (N_5009,N_4171,N_4874);
nor U5010 (N_5010,N_4283,N_4130);
and U5011 (N_5011,N_4025,N_4947);
or U5012 (N_5012,N_4318,N_4886);
or U5013 (N_5013,N_4268,N_4215);
and U5014 (N_5014,N_4077,N_4309);
nor U5015 (N_5015,N_4788,N_4261);
nor U5016 (N_5016,N_4009,N_4576);
nor U5017 (N_5017,N_4708,N_4816);
or U5018 (N_5018,N_4831,N_4490);
nor U5019 (N_5019,N_4562,N_4999);
and U5020 (N_5020,N_4817,N_4698);
or U5021 (N_5021,N_4974,N_4300);
and U5022 (N_5022,N_4688,N_4715);
nor U5023 (N_5023,N_4236,N_4990);
or U5024 (N_5024,N_4131,N_4053);
or U5025 (N_5025,N_4328,N_4552);
and U5026 (N_5026,N_4257,N_4159);
nand U5027 (N_5027,N_4804,N_4881);
and U5028 (N_5028,N_4457,N_4961);
or U5029 (N_5029,N_4900,N_4614);
and U5030 (N_5030,N_4436,N_4085);
nand U5031 (N_5031,N_4369,N_4665);
or U5032 (N_5032,N_4593,N_4448);
and U5033 (N_5033,N_4579,N_4679);
nor U5034 (N_5034,N_4557,N_4212);
nor U5035 (N_5035,N_4342,N_4591);
and U5036 (N_5036,N_4943,N_4118);
or U5037 (N_5037,N_4882,N_4966);
or U5038 (N_5038,N_4287,N_4043);
or U5039 (N_5039,N_4237,N_4428);
nor U5040 (N_5040,N_4983,N_4808);
and U5041 (N_5041,N_4850,N_4909);
or U5042 (N_5042,N_4339,N_4516);
and U5043 (N_5043,N_4948,N_4035);
or U5044 (N_5044,N_4365,N_4381);
or U5045 (N_5045,N_4202,N_4356);
nand U5046 (N_5046,N_4327,N_4537);
nand U5047 (N_5047,N_4613,N_4656);
and U5048 (N_5048,N_4050,N_4061);
or U5049 (N_5049,N_4226,N_4308);
nand U5050 (N_5050,N_4336,N_4600);
or U5051 (N_5051,N_4924,N_4921);
and U5052 (N_5052,N_4723,N_4539);
nand U5053 (N_5053,N_4806,N_4620);
or U5054 (N_5054,N_4861,N_4640);
nand U5055 (N_5055,N_4542,N_4774);
or U5056 (N_5056,N_4623,N_4524);
nor U5057 (N_5057,N_4015,N_4271);
nand U5058 (N_5058,N_4345,N_4791);
nor U5059 (N_5059,N_4293,N_4841);
and U5060 (N_5060,N_4496,N_4707);
or U5061 (N_5061,N_4721,N_4095);
and U5062 (N_5062,N_4568,N_4086);
and U5063 (N_5063,N_4695,N_4389);
and U5064 (N_5064,N_4891,N_4151);
nor U5065 (N_5065,N_4464,N_4472);
and U5066 (N_5066,N_4144,N_4439);
xor U5067 (N_5067,N_4556,N_4809);
and U5068 (N_5068,N_4396,N_4757);
and U5069 (N_5069,N_4184,N_4361);
or U5070 (N_5070,N_4631,N_4001);
or U5071 (N_5071,N_4670,N_4551);
and U5072 (N_5072,N_4330,N_4824);
nand U5073 (N_5073,N_4957,N_4278);
and U5074 (N_5074,N_4923,N_4857);
and U5075 (N_5075,N_4741,N_4155);
or U5076 (N_5076,N_4852,N_4701);
or U5077 (N_5077,N_4682,N_4334);
nor U5078 (N_5078,N_4792,N_4559);
nand U5079 (N_5079,N_4965,N_4451);
nor U5080 (N_5080,N_4069,N_4262);
nand U5081 (N_5081,N_4223,N_4126);
and U5082 (N_5082,N_4219,N_4067);
nor U5083 (N_5083,N_4853,N_4865);
or U5084 (N_5084,N_4054,N_4952);
or U5085 (N_5085,N_4863,N_4437);
nor U5086 (N_5086,N_4843,N_4578);
nand U5087 (N_5087,N_4916,N_4522);
nand U5088 (N_5088,N_4773,N_4398);
nand U5089 (N_5089,N_4798,N_4628);
nor U5090 (N_5090,N_4145,N_4822);
and U5091 (N_5091,N_4705,N_4718);
nor U5092 (N_5092,N_4094,N_4913);
nand U5093 (N_5093,N_4956,N_4739);
nor U5094 (N_5094,N_4344,N_4927);
and U5095 (N_5095,N_4662,N_4232);
nand U5096 (N_5096,N_4373,N_4500);
nand U5097 (N_5097,N_4580,N_4427);
and U5098 (N_5098,N_4049,N_4429);
or U5099 (N_5099,N_4512,N_4088);
and U5100 (N_5100,N_4146,N_4897);
nand U5101 (N_5101,N_4386,N_4058);
nor U5102 (N_5102,N_4477,N_4851);
or U5103 (N_5103,N_4609,N_4107);
or U5104 (N_5104,N_4141,N_4314);
nor U5105 (N_5105,N_4848,N_4374);
and U5106 (N_5106,N_4823,N_4685);
or U5107 (N_5107,N_4795,N_4080);
or U5108 (N_5108,N_4972,N_4175);
or U5109 (N_5109,N_4438,N_4097);
and U5110 (N_5110,N_4370,N_4284);
nand U5111 (N_5111,N_4412,N_4960);
and U5112 (N_5112,N_4127,N_4581);
and U5113 (N_5113,N_4915,N_4790);
nand U5114 (N_5114,N_4363,N_4855);
nand U5115 (N_5115,N_4978,N_4819);
nand U5116 (N_5116,N_4598,N_4986);
nor U5117 (N_5117,N_4945,N_4286);
nor U5118 (N_5118,N_4291,N_4243);
or U5119 (N_5119,N_4977,N_4310);
nand U5120 (N_5120,N_4265,N_4020);
nor U5121 (N_5121,N_4198,N_4266);
nor U5122 (N_5122,N_4583,N_4519);
nand U5123 (N_5123,N_4811,N_4486);
nor U5124 (N_5124,N_4743,N_4332);
nand U5125 (N_5125,N_4611,N_4919);
nor U5126 (N_5126,N_4488,N_4117);
or U5127 (N_5127,N_4892,N_4466);
nor U5128 (N_5128,N_4717,N_4696);
nor U5129 (N_5129,N_4324,N_4964);
or U5130 (N_5130,N_4836,N_4197);
xor U5131 (N_5131,N_4734,N_4469);
and U5132 (N_5132,N_4419,N_4164);
or U5133 (N_5133,N_4047,N_4549);
nand U5134 (N_5134,N_4733,N_4526);
nand U5135 (N_5135,N_4442,N_4148);
nor U5136 (N_5136,N_4112,N_4962);
nand U5137 (N_5137,N_4358,N_4125);
or U5138 (N_5138,N_4289,N_4675);
nor U5139 (N_5139,N_4042,N_4989);
nor U5140 (N_5140,N_4652,N_4478);
and U5141 (N_5141,N_4585,N_4725);
and U5142 (N_5142,N_4220,N_4895);
nor U5143 (N_5143,N_4239,N_4747);
nor U5144 (N_5144,N_4993,N_4235);
and U5145 (N_5145,N_4668,N_4258);
and U5146 (N_5146,N_4941,N_4632);
and U5147 (N_5147,N_4218,N_4254);
nor U5148 (N_5148,N_4390,N_4746);
nand U5149 (N_5149,N_4608,N_4564);
or U5150 (N_5150,N_4311,N_4022);
nor U5151 (N_5151,N_4584,N_4250);
or U5152 (N_5152,N_4996,N_4432);
nand U5153 (N_5153,N_4654,N_4535);
nand U5154 (N_5154,N_4669,N_4818);
nor U5155 (N_5155,N_4301,N_4887);
or U5156 (N_5156,N_4446,N_4060);
nor U5157 (N_5157,N_4749,N_4622);
nor U5158 (N_5158,N_4907,N_4498);
and U5159 (N_5159,N_4099,N_4994);
nand U5160 (N_5160,N_4742,N_4767);
and U5161 (N_5161,N_4636,N_4511);
nor U5162 (N_5162,N_4615,N_4967);
and U5163 (N_5163,N_4467,N_4105);
nand U5164 (N_5164,N_4082,N_4862);
nand U5165 (N_5165,N_4177,N_4329);
or U5166 (N_5166,N_4513,N_4573);
nand U5167 (N_5167,N_4109,N_4182);
nand U5168 (N_5168,N_4671,N_4313);
nand U5169 (N_5169,N_4722,N_4139);
or U5170 (N_5170,N_4248,N_4596);
nand U5171 (N_5171,N_4482,N_4737);
nor U5172 (N_5172,N_4771,N_4812);
nand U5173 (N_5173,N_4027,N_4303);
or U5174 (N_5174,N_4637,N_4758);
and U5175 (N_5175,N_4331,N_4917);
nor U5176 (N_5176,N_4461,N_4735);
nor U5177 (N_5177,N_4465,N_4922);
or U5178 (N_5178,N_4201,N_4487);
and U5179 (N_5179,N_4252,N_4355);
nand U5180 (N_5180,N_4221,N_4294);
nand U5181 (N_5181,N_4713,N_4242);
nand U5182 (N_5182,N_4877,N_4506);
and U5183 (N_5183,N_4878,N_4902);
nand U5184 (N_5184,N_4306,N_4190);
or U5185 (N_5185,N_4660,N_4980);
nand U5186 (N_5186,N_4971,N_4642);
nor U5187 (N_5187,N_4021,N_4794);
nor U5188 (N_5188,N_4727,N_4188);
nand U5189 (N_5189,N_4485,N_4147);
or U5190 (N_5190,N_4091,N_4343);
nand U5191 (N_5191,N_4183,N_4434);
nand U5192 (N_5192,N_4264,N_4920);
and U5193 (N_5193,N_4114,N_4548);
or U5194 (N_5194,N_4435,N_4592);
or U5195 (N_5195,N_4787,N_4859);
nand U5196 (N_5196,N_4969,N_4203);
nand U5197 (N_5197,N_4532,N_4784);
and U5198 (N_5198,N_4894,N_4152);
or U5199 (N_5199,N_4325,N_4193);
or U5200 (N_5200,N_4534,N_4899);
nor U5201 (N_5201,N_4450,N_4383);
and U5202 (N_5202,N_4233,N_4425);
and U5203 (N_5203,N_4906,N_4992);
nand U5204 (N_5204,N_4453,N_4167);
nor U5205 (N_5205,N_4693,N_4520);
and U5206 (N_5206,N_4805,N_4686);
nor U5207 (N_5207,N_4814,N_4936);
nand U5208 (N_5208,N_4449,N_4418);
nand U5209 (N_5209,N_4738,N_4333);
or U5210 (N_5210,N_4560,N_4316);
nor U5211 (N_5211,N_4647,N_4627);
nor U5212 (N_5212,N_4068,N_4904);
and U5213 (N_5213,N_4244,N_4351);
nand U5214 (N_5214,N_4483,N_4277);
or U5215 (N_5215,N_4540,N_4426);
nor U5216 (N_5216,N_4801,N_4828);
nand U5217 (N_5217,N_4006,N_4950);
or U5218 (N_5218,N_4566,N_4528);
or U5219 (N_5219,N_4111,N_4644);
nand U5220 (N_5220,N_4388,N_4910);
nand U5221 (N_5221,N_4658,N_4903);
nor U5222 (N_5222,N_4140,N_4555);
or U5223 (N_5223,N_4104,N_4588);
or U5224 (N_5224,N_4399,N_4765);
nor U5225 (N_5225,N_4751,N_4543);
or U5226 (N_5226,N_4803,N_4603);
nor U5227 (N_5227,N_4700,N_4259);
nor U5228 (N_5228,N_4222,N_4527);
and U5229 (N_5229,N_4982,N_4946);
nor U5230 (N_5230,N_4157,N_4406);
xnor U5231 (N_5231,N_4247,N_4234);
nand U5232 (N_5232,N_4869,N_4979);
nand U5233 (N_5233,N_4835,N_4995);
and U5234 (N_5234,N_4174,N_4447);
nor U5235 (N_5235,N_4181,N_4100);
nand U5236 (N_5236,N_4200,N_4275);
nor U5237 (N_5237,N_4711,N_4650);
or U5238 (N_5238,N_4829,N_4769);
or U5239 (N_5239,N_4832,N_4624);
and U5240 (N_5240,N_4031,N_4504);
nor U5241 (N_5241,N_4224,N_4297);
or U5242 (N_5242,N_4000,N_4845);
and U5243 (N_5243,N_4868,N_4376);
nand U5244 (N_5244,N_4385,N_4322);
nor U5245 (N_5245,N_4770,N_4230);
or U5246 (N_5246,N_4616,N_4057);
or U5247 (N_5247,N_4606,N_4797);
and U5248 (N_5248,N_4856,N_4393);
or U5249 (N_5249,N_4368,N_4028);
and U5250 (N_5250,N_4612,N_4976);
and U5251 (N_5251,N_4176,N_4002);
nand U5252 (N_5252,N_4825,N_4350);
nand U5253 (N_5253,N_4191,N_4371);
or U5254 (N_5254,N_4505,N_4984);
nor U5255 (N_5255,N_4462,N_4626);
nor U5256 (N_5256,N_4410,N_4925);
or U5257 (N_5257,N_4546,N_4607);
and U5258 (N_5258,N_4629,N_4380);
or U5259 (N_5259,N_4893,N_4347);
and U5260 (N_5260,N_4037,N_4531);
nand U5261 (N_5261,N_4052,N_4321);
nor U5262 (N_5262,N_4677,N_4515);
nand U5263 (N_5263,N_4096,N_4137);
nor U5264 (N_5264,N_4110,N_4003);
nand U5265 (N_5265,N_4683,N_4392);
nor U5266 (N_5266,N_4459,N_4366);
or U5267 (N_5267,N_4760,N_4064);
or U5268 (N_5268,N_4409,N_4023);
nand U5269 (N_5269,N_4170,N_4680);
and U5270 (N_5270,N_4860,N_4225);
nand U5271 (N_5271,N_4208,N_4720);
nor U5272 (N_5272,N_4988,N_4569);
nand U5273 (N_5273,N_4864,N_4959);
or U5274 (N_5274,N_4352,N_4502);
or U5275 (N_5275,N_4838,N_4673);
nor U5276 (N_5276,N_4648,N_4076);
nand U5277 (N_5277,N_4227,N_4231);
and U5278 (N_5278,N_4414,N_4518);
or U5279 (N_5279,N_4038,N_4158);
and U5280 (N_5280,N_4128,N_4731);
nor U5281 (N_5281,N_4207,N_4292);
nand U5282 (N_5282,N_4185,N_4776);
nor U5283 (N_5283,N_4149,N_4589);
and U5284 (N_5284,N_4530,N_4282);
nor U5285 (N_5285,N_4016,N_4525);
nor U5286 (N_5286,N_4196,N_4684);
nand U5287 (N_5287,N_4763,N_4572);
or U5288 (N_5288,N_4699,N_4541);
or U5289 (N_5289,N_4544,N_4093);
nand U5290 (N_5290,N_4103,N_4382);
nand U5291 (N_5291,N_4092,N_4229);
or U5292 (N_5292,N_4929,N_4470);
nand U5293 (N_5293,N_4211,N_4353);
or U5294 (N_5294,N_4712,N_4529);
or U5295 (N_5295,N_4618,N_4667);
nand U5296 (N_5296,N_4348,N_4844);
and U5297 (N_5297,N_4367,N_4270);
nand U5298 (N_5298,N_4846,N_4694);
nand U5299 (N_5299,N_4926,N_4349);
nor U5300 (N_5300,N_4172,N_4858);
and U5301 (N_5301,N_4681,N_4499);
and U5302 (N_5302,N_4168,N_4113);
and U5303 (N_5303,N_4046,N_4178);
nand U5304 (N_5304,N_4587,N_4768);
nor U5305 (N_5305,N_4827,N_4317);
and U5306 (N_5306,N_4026,N_4195);
nor U5307 (N_5307,N_4143,N_4663);
nor U5308 (N_5308,N_4871,N_4084);
nand U5309 (N_5309,N_4692,N_4337);
and U5310 (N_5310,N_4752,N_4884);
nand U5311 (N_5311,N_4228,N_4610);
or U5312 (N_5312,N_4165,N_4879);
or U5313 (N_5313,N_4444,N_4617);
nand U5314 (N_5314,N_4565,N_4762);
nand U5315 (N_5315,N_4558,N_4704);
or U5316 (N_5316,N_4004,N_4173);
or U5317 (N_5317,N_4796,N_4605);
nor U5318 (N_5318,N_4411,N_4471);
and U5319 (N_5319,N_4189,N_4997);
or U5320 (N_5320,N_4599,N_4839);
nand U5321 (N_5321,N_4378,N_4199);
or U5322 (N_5322,N_4070,N_4575);
or U5323 (N_5323,N_4998,N_4408);
or U5324 (N_5324,N_4550,N_4205);
nor U5325 (N_5325,N_4706,N_4940);
nor U5326 (N_5326,N_4420,N_4475);
and U5327 (N_5327,N_4582,N_4187);
or U5328 (N_5328,N_4071,N_4341);
and U5329 (N_5329,N_4645,N_4073);
nand U5330 (N_5330,N_4161,N_4304);
or U5331 (N_5331,N_4338,N_4641);
nand U5332 (N_5332,N_4981,N_4033);
or U5333 (N_5333,N_4285,N_4780);
and U5334 (N_5334,N_4008,N_4933);
or U5335 (N_5335,N_4753,N_4820);
and U5336 (N_5336,N_4075,N_4290);
nor U5337 (N_5337,N_4346,N_4013);
nor U5338 (N_5338,N_4586,N_4842);
nor U5339 (N_5339,N_4666,N_4837);
nor U5340 (N_5340,N_4423,N_4281);
nor U5341 (N_5341,N_4040,N_4280);
and U5342 (N_5342,N_4521,N_4441);
nor U5343 (N_5343,N_4039,N_4400);
nand U5344 (N_5344,N_4594,N_4276);
nand U5345 (N_5345,N_4810,N_4873);
nor U5346 (N_5346,N_4206,N_4570);
or U5347 (N_5347,N_4431,N_4005);
or U5348 (N_5348,N_4975,N_4918);
nor U5349 (N_5349,N_4405,N_4779);
nand U5350 (N_5350,N_4413,N_4826);
nor U5351 (N_5351,N_4939,N_4326);
nor U5352 (N_5352,N_4030,N_4876);
nand U5353 (N_5353,N_4364,N_4036);
and U5354 (N_5354,N_4942,N_4253);
nor U5355 (N_5355,N_4136,N_4938);
or U5356 (N_5356,N_4934,N_4689);
and U5357 (N_5357,N_4362,N_4194);
nor U5358 (N_5358,N_4204,N_4951);
nor U5359 (N_5359,N_4571,N_4017);
or U5360 (N_5360,N_4401,N_4510);
xor U5361 (N_5361,N_4452,N_4416);
nand U5362 (N_5362,N_4090,N_4260);
or U5363 (N_5363,N_4209,N_4012);
and U5364 (N_5364,N_4299,N_4690);
and U5365 (N_5365,N_4056,N_4384);
or U5366 (N_5366,N_4653,N_4422);
or U5367 (N_5367,N_4460,N_4655);
and U5368 (N_5368,N_4911,N_4034);
and U5369 (N_5369,N_4639,N_4724);
nand U5370 (N_5370,N_4732,N_4750);
and U5371 (N_5371,N_4163,N_4273);
nand U5372 (N_5372,N_4192,N_4872);
nor U5373 (N_5373,N_4710,N_4272);
and U5374 (N_5374,N_4935,N_4083);
nor U5375 (N_5375,N_4468,N_4079);
nand U5376 (N_5376,N_4885,N_4256);
and U5377 (N_5377,N_4119,N_4968);
nor U5378 (N_5378,N_4072,N_4875);
nor U5379 (N_5379,N_4415,N_4799);
nor U5380 (N_5380,N_4937,N_4736);
and U5381 (N_5381,N_4595,N_4987);
or U5382 (N_5382,N_4440,N_4395);
nor U5383 (N_5383,N_4007,N_4404);
nor U5384 (N_5384,N_4778,N_4577);
and U5385 (N_5385,N_4240,N_4180);
nor U5386 (N_5386,N_4379,N_4766);
and U5387 (N_5387,N_4357,N_4635);
or U5388 (N_5388,N_4150,N_4932);
and U5389 (N_5389,N_4377,N_4407);
nor U5390 (N_5390,N_4402,N_4169);
nand U5391 (N_5391,N_4269,N_4755);
nor U5392 (N_5392,N_4786,N_4296);
or U5393 (N_5393,N_4538,N_4867);
or U5394 (N_5394,N_4726,N_4970);
or U5395 (N_5395,N_4728,N_4928);
nand U5396 (N_5396,N_4359,N_4702);
or U5397 (N_5397,N_4691,N_4066);
or U5398 (N_5398,N_4800,N_4456);
nand U5399 (N_5399,N_4661,N_4509);
nor U5400 (N_5400,N_4883,N_4563);
nand U5401 (N_5401,N_4953,N_4081);
and U5402 (N_5402,N_4649,N_4714);
and U5403 (N_5403,N_4602,N_4898);
or U5404 (N_5404,N_4754,N_4479);
nor U5405 (N_5405,N_4101,N_4394);
or U5406 (N_5406,N_4055,N_4032);
nand U5407 (N_5407,N_4497,N_4315);
nand U5408 (N_5408,N_4888,N_4847);
or U5409 (N_5409,N_4387,N_4089);
nand U5410 (N_5410,N_4455,N_4687);
or U5411 (N_5411,N_4764,N_4604);
or U5412 (N_5412,N_4323,N_4912);
or U5413 (N_5413,N_4672,N_4134);
or U5414 (N_5414,N_4651,N_4866);
and U5415 (N_5415,N_4621,N_4476);
nand U5416 (N_5416,N_4115,N_4295);
nand U5417 (N_5417,N_4397,N_4123);
and U5418 (N_5418,N_4914,N_4263);
nand U5419 (N_5419,N_4703,N_4458);
or U5420 (N_5420,N_4319,N_4051);
nor U5421 (N_5421,N_4840,N_4944);
nor U5422 (N_5422,N_4484,N_4014);
nand U5423 (N_5423,N_4833,N_4106);
or U5424 (N_5424,N_4010,N_4730);
and U5425 (N_5425,N_4508,N_4494);
and U5426 (N_5426,N_4954,N_4501);
or U5427 (N_5427,N_4716,N_4124);
xnor U5428 (N_5428,N_4930,N_4491);
nor U5429 (N_5429,N_4102,N_4756);
or U5430 (N_5430,N_4241,N_4213);
or U5431 (N_5431,N_4391,N_4740);
nand U5432 (N_5432,N_4044,N_4630);
or U5433 (N_5433,N_4821,N_4246);
and U5434 (N_5434,N_4949,N_4011);
nand U5435 (N_5435,N_4288,N_4065);
nor U5436 (N_5436,N_4154,N_4298);
nand U5437 (N_5437,N_4305,N_4545);
nor U5438 (N_5438,N_4421,N_4216);
nand U5439 (N_5439,N_4813,N_4815);
or U5440 (N_5440,N_4514,N_4772);
nand U5441 (N_5441,N_4433,N_4019);
nor U5442 (N_5442,N_4517,N_4781);
nand U5443 (N_5443,N_4179,N_4495);
and U5444 (N_5444,N_4880,N_4601);
nand U5445 (N_5445,N_4210,N_4958);
or U5446 (N_5446,N_4785,N_4676);
nand U5447 (N_5447,N_4729,N_4963);
or U5448 (N_5448,N_4463,N_4255);
or U5449 (N_5449,N_4709,N_4360);
nor U5450 (N_5450,N_4133,N_4554);
nand U5451 (N_5451,N_4138,N_4120);
or U5452 (N_5452,N_4312,N_4783);
and U5453 (N_5453,N_4547,N_4238);
and U5454 (N_5454,N_4507,N_4633);
and U5455 (N_5455,N_4973,N_4074);
and U5456 (N_5456,N_4041,N_4267);
nand U5457 (N_5457,N_4063,N_4166);
nand U5458 (N_5458,N_4748,N_4129);
and U5459 (N_5459,N_4424,N_4782);
and U5460 (N_5460,N_4745,N_4048);
and U5461 (N_5461,N_4492,N_4759);
or U5462 (N_5462,N_4674,N_4646);
or U5463 (N_5463,N_4132,N_4634);
nor U5464 (N_5464,N_4135,N_4417);
nor U5465 (N_5465,N_4480,N_4830);
and U5466 (N_5466,N_4567,N_4335);
or U5467 (N_5467,N_4445,N_4802);
nor U5468 (N_5468,N_4889,N_4896);
nand U5469 (N_5469,N_4062,N_4214);
nand U5470 (N_5470,N_4870,N_4523);
or U5471 (N_5471,N_4503,N_4320);
nand U5472 (N_5472,N_4443,N_4274);
nand U5473 (N_5473,N_4793,N_4160);
and U5474 (N_5474,N_4659,N_4018);
or U5475 (N_5475,N_4354,N_4643);
and U5476 (N_5476,N_4279,N_4985);
and U5477 (N_5477,N_4991,N_4697);
or U5478 (N_5478,N_4908,N_4430);
nor U5479 (N_5479,N_4403,N_4777);
nor U5480 (N_5480,N_4108,N_4854);
and U5481 (N_5481,N_4619,N_4553);
nor U5482 (N_5482,N_4087,N_4849);
or U5483 (N_5483,N_4251,N_4834);
nand U5484 (N_5484,N_4901,N_4162);
and U5485 (N_5485,N_4890,N_4375);
and U5486 (N_5486,N_4493,N_4955);
and U5487 (N_5487,N_4536,N_4533);
or U5488 (N_5488,N_4245,N_4474);
nand U5489 (N_5489,N_4186,N_4481);
or U5490 (N_5490,N_4142,N_4045);
and U5491 (N_5491,N_4078,N_4561);
or U5492 (N_5492,N_4664,N_4625);
nor U5493 (N_5493,N_4249,N_4761);
nand U5494 (N_5494,N_4122,N_4029);
and U5495 (N_5495,N_4059,N_4473);
or U5496 (N_5496,N_4657,N_4340);
nand U5497 (N_5497,N_4807,N_4574);
xor U5498 (N_5498,N_4590,N_4156);
nand U5499 (N_5499,N_4744,N_4905);
or U5500 (N_5500,N_4542,N_4016);
nor U5501 (N_5501,N_4663,N_4865);
or U5502 (N_5502,N_4372,N_4678);
or U5503 (N_5503,N_4281,N_4181);
nand U5504 (N_5504,N_4769,N_4511);
or U5505 (N_5505,N_4105,N_4938);
and U5506 (N_5506,N_4418,N_4885);
or U5507 (N_5507,N_4113,N_4891);
nor U5508 (N_5508,N_4809,N_4908);
nor U5509 (N_5509,N_4911,N_4582);
nand U5510 (N_5510,N_4939,N_4253);
nand U5511 (N_5511,N_4050,N_4663);
nand U5512 (N_5512,N_4113,N_4145);
or U5513 (N_5513,N_4570,N_4582);
nand U5514 (N_5514,N_4480,N_4821);
or U5515 (N_5515,N_4635,N_4536);
nor U5516 (N_5516,N_4010,N_4038);
and U5517 (N_5517,N_4330,N_4387);
nor U5518 (N_5518,N_4591,N_4493);
or U5519 (N_5519,N_4836,N_4609);
or U5520 (N_5520,N_4199,N_4249);
or U5521 (N_5521,N_4830,N_4651);
or U5522 (N_5522,N_4753,N_4030);
xnor U5523 (N_5523,N_4502,N_4224);
and U5524 (N_5524,N_4271,N_4201);
or U5525 (N_5525,N_4738,N_4222);
nor U5526 (N_5526,N_4694,N_4130);
and U5527 (N_5527,N_4732,N_4370);
or U5528 (N_5528,N_4935,N_4991);
and U5529 (N_5529,N_4771,N_4393);
or U5530 (N_5530,N_4116,N_4861);
nor U5531 (N_5531,N_4530,N_4143);
nor U5532 (N_5532,N_4211,N_4093);
or U5533 (N_5533,N_4613,N_4675);
or U5534 (N_5534,N_4080,N_4648);
nor U5535 (N_5535,N_4735,N_4331);
nand U5536 (N_5536,N_4362,N_4926);
or U5537 (N_5537,N_4987,N_4094);
or U5538 (N_5538,N_4656,N_4832);
nand U5539 (N_5539,N_4289,N_4367);
nand U5540 (N_5540,N_4628,N_4203);
nor U5541 (N_5541,N_4767,N_4092);
or U5542 (N_5542,N_4618,N_4836);
nand U5543 (N_5543,N_4915,N_4527);
and U5544 (N_5544,N_4170,N_4700);
and U5545 (N_5545,N_4424,N_4039);
or U5546 (N_5546,N_4174,N_4932);
and U5547 (N_5547,N_4688,N_4977);
and U5548 (N_5548,N_4547,N_4253);
nand U5549 (N_5549,N_4652,N_4286);
and U5550 (N_5550,N_4849,N_4009);
nand U5551 (N_5551,N_4029,N_4800);
or U5552 (N_5552,N_4373,N_4572);
and U5553 (N_5553,N_4907,N_4233);
or U5554 (N_5554,N_4265,N_4989);
nand U5555 (N_5555,N_4147,N_4220);
nand U5556 (N_5556,N_4067,N_4883);
nor U5557 (N_5557,N_4766,N_4087);
xor U5558 (N_5558,N_4864,N_4160);
and U5559 (N_5559,N_4967,N_4935);
and U5560 (N_5560,N_4860,N_4547);
and U5561 (N_5561,N_4237,N_4640);
or U5562 (N_5562,N_4690,N_4843);
nand U5563 (N_5563,N_4101,N_4927);
nand U5564 (N_5564,N_4073,N_4052);
and U5565 (N_5565,N_4750,N_4567);
or U5566 (N_5566,N_4680,N_4901);
nand U5567 (N_5567,N_4107,N_4183);
nand U5568 (N_5568,N_4978,N_4091);
and U5569 (N_5569,N_4628,N_4958);
or U5570 (N_5570,N_4200,N_4731);
and U5571 (N_5571,N_4007,N_4469);
and U5572 (N_5572,N_4185,N_4086);
and U5573 (N_5573,N_4830,N_4201);
nor U5574 (N_5574,N_4181,N_4893);
nand U5575 (N_5575,N_4733,N_4509);
nand U5576 (N_5576,N_4572,N_4552);
and U5577 (N_5577,N_4307,N_4921);
or U5578 (N_5578,N_4321,N_4707);
nor U5579 (N_5579,N_4062,N_4091);
nor U5580 (N_5580,N_4497,N_4709);
or U5581 (N_5581,N_4286,N_4506);
nand U5582 (N_5582,N_4992,N_4338);
nand U5583 (N_5583,N_4142,N_4673);
and U5584 (N_5584,N_4224,N_4012);
nand U5585 (N_5585,N_4101,N_4979);
nor U5586 (N_5586,N_4005,N_4572);
or U5587 (N_5587,N_4233,N_4186);
nand U5588 (N_5588,N_4374,N_4518);
and U5589 (N_5589,N_4191,N_4850);
or U5590 (N_5590,N_4204,N_4264);
nand U5591 (N_5591,N_4346,N_4010);
nor U5592 (N_5592,N_4658,N_4387);
and U5593 (N_5593,N_4061,N_4363);
nor U5594 (N_5594,N_4825,N_4288);
or U5595 (N_5595,N_4097,N_4411);
and U5596 (N_5596,N_4529,N_4332);
nor U5597 (N_5597,N_4429,N_4643);
nor U5598 (N_5598,N_4832,N_4445);
or U5599 (N_5599,N_4520,N_4739);
or U5600 (N_5600,N_4485,N_4207);
and U5601 (N_5601,N_4392,N_4621);
nand U5602 (N_5602,N_4895,N_4133);
nand U5603 (N_5603,N_4352,N_4748);
or U5604 (N_5604,N_4311,N_4218);
and U5605 (N_5605,N_4337,N_4585);
nand U5606 (N_5606,N_4393,N_4256);
and U5607 (N_5607,N_4399,N_4743);
nand U5608 (N_5608,N_4583,N_4253);
or U5609 (N_5609,N_4400,N_4648);
nand U5610 (N_5610,N_4504,N_4205);
xnor U5611 (N_5611,N_4036,N_4981);
nand U5612 (N_5612,N_4792,N_4533);
or U5613 (N_5613,N_4888,N_4485);
nor U5614 (N_5614,N_4872,N_4490);
nor U5615 (N_5615,N_4455,N_4716);
and U5616 (N_5616,N_4696,N_4465);
nor U5617 (N_5617,N_4294,N_4366);
and U5618 (N_5618,N_4945,N_4869);
nor U5619 (N_5619,N_4226,N_4314);
and U5620 (N_5620,N_4865,N_4306);
nand U5621 (N_5621,N_4621,N_4140);
or U5622 (N_5622,N_4150,N_4795);
nor U5623 (N_5623,N_4986,N_4422);
nor U5624 (N_5624,N_4570,N_4228);
or U5625 (N_5625,N_4110,N_4840);
or U5626 (N_5626,N_4024,N_4618);
nand U5627 (N_5627,N_4576,N_4073);
nor U5628 (N_5628,N_4873,N_4897);
or U5629 (N_5629,N_4744,N_4422);
nor U5630 (N_5630,N_4454,N_4754);
or U5631 (N_5631,N_4626,N_4924);
or U5632 (N_5632,N_4471,N_4632);
or U5633 (N_5633,N_4218,N_4918);
or U5634 (N_5634,N_4541,N_4756);
and U5635 (N_5635,N_4379,N_4011);
nor U5636 (N_5636,N_4339,N_4093);
and U5637 (N_5637,N_4002,N_4461);
or U5638 (N_5638,N_4056,N_4889);
nand U5639 (N_5639,N_4813,N_4604);
or U5640 (N_5640,N_4151,N_4370);
nand U5641 (N_5641,N_4612,N_4930);
nand U5642 (N_5642,N_4286,N_4160);
or U5643 (N_5643,N_4565,N_4251);
and U5644 (N_5644,N_4826,N_4496);
and U5645 (N_5645,N_4023,N_4332);
and U5646 (N_5646,N_4485,N_4262);
nand U5647 (N_5647,N_4869,N_4069);
and U5648 (N_5648,N_4322,N_4441);
nor U5649 (N_5649,N_4421,N_4798);
or U5650 (N_5650,N_4530,N_4797);
or U5651 (N_5651,N_4043,N_4744);
nor U5652 (N_5652,N_4495,N_4566);
nand U5653 (N_5653,N_4003,N_4281);
and U5654 (N_5654,N_4517,N_4714);
nor U5655 (N_5655,N_4390,N_4687);
nand U5656 (N_5656,N_4527,N_4515);
nor U5657 (N_5657,N_4482,N_4151);
and U5658 (N_5658,N_4245,N_4338);
and U5659 (N_5659,N_4984,N_4552);
nor U5660 (N_5660,N_4758,N_4145);
and U5661 (N_5661,N_4467,N_4832);
or U5662 (N_5662,N_4246,N_4252);
and U5663 (N_5663,N_4422,N_4297);
nand U5664 (N_5664,N_4290,N_4436);
nand U5665 (N_5665,N_4911,N_4212);
nand U5666 (N_5666,N_4038,N_4865);
or U5667 (N_5667,N_4506,N_4685);
nor U5668 (N_5668,N_4639,N_4016);
nor U5669 (N_5669,N_4412,N_4283);
and U5670 (N_5670,N_4198,N_4181);
and U5671 (N_5671,N_4883,N_4986);
or U5672 (N_5672,N_4041,N_4445);
or U5673 (N_5673,N_4884,N_4349);
nor U5674 (N_5674,N_4472,N_4886);
nor U5675 (N_5675,N_4409,N_4845);
nand U5676 (N_5676,N_4235,N_4513);
or U5677 (N_5677,N_4348,N_4545);
nand U5678 (N_5678,N_4205,N_4875);
nand U5679 (N_5679,N_4960,N_4270);
or U5680 (N_5680,N_4709,N_4441);
or U5681 (N_5681,N_4387,N_4619);
or U5682 (N_5682,N_4505,N_4555);
nor U5683 (N_5683,N_4702,N_4394);
nor U5684 (N_5684,N_4153,N_4092);
and U5685 (N_5685,N_4833,N_4981);
nor U5686 (N_5686,N_4645,N_4147);
nor U5687 (N_5687,N_4556,N_4756);
and U5688 (N_5688,N_4376,N_4724);
or U5689 (N_5689,N_4991,N_4424);
and U5690 (N_5690,N_4033,N_4748);
nor U5691 (N_5691,N_4948,N_4596);
nor U5692 (N_5692,N_4858,N_4614);
or U5693 (N_5693,N_4626,N_4604);
and U5694 (N_5694,N_4758,N_4871);
nor U5695 (N_5695,N_4633,N_4140);
or U5696 (N_5696,N_4888,N_4570);
nor U5697 (N_5697,N_4765,N_4660);
and U5698 (N_5698,N_4054,N_4394);
and U5699 (N_5699,N_4366,N_4839);
nor U5700 (N_5700,N_4026,N_4919);
nand U5701 (N_5701,N_4923,N_4768);
nor U5702 (N_5702,N_4446,N_4467);
nor U5703 (N_5703,N_4544,N_4498);
and U5704 (N_5704,N_4291,N_4206);
nor U5705 (N_5705,N_4583,N_4538);
and U5706 (N_5706,N_4091,N_4736);
nor U5707 (N_5707,N_4979,N_4673);
nand U5708 (N_5708,N_4645,N_4630);
nand U5709 (N_5709,N_4770,N_4942);
nand U5710 (N_5710,N_4213,N_4089);
nand U5711 (N_5711,N_4811,N_4271);
and U5712 (N_5712,N_4184,N_4672);
nor U5713 (N_5713,N_4351,N_4401);
or U5714 (N_5714,N_4543,N_4285);
nand U5715 (N_5715,N_4672,N_4172);
or U5716 (N_5716,N_4381,N_4257);
and U5717 (N_5717,N_4985,N_4290);
or U5718 (N_5718,N_4404,N_4960);
and U5719 (N_5719,N_4296,N_4967);
nor U5720 (N_5720,N_4080,N_4915);
or U5721 (N_5721,N_4934,N_4587);
nor U5722 (N_5722,N_4016,N_4841);
and U5723 (N_5723,N_4608,N_4325);
and U5724 (N_5724,N_4382,N_4337);
nor U5725 (N_5725,N_4319,N_4275);
nor U5726 (N_5726,N_4277,N_4898);
nor U5727 (N_5727,N_4380,N_4338);
nand U5728 (N_5728,N_4111,N_4106);
nand U5729 (N_5729,N_4224,N_4769);
nor U5730 (N_5730,N_4197,N_4390);
nor U5731 (N_5731,N_4314,N_4875);
nor U5732 (N_5732,N_4082,N_4117);
or U5733 (N_5733,N_4855,N_4627);
nand U5734 (N_5734,N_4857,N_4221);
or U5735 (N_5735,N_4754,N_4963);
or U5736 (N_5736,N_4095,N_4624);
nand U5737 (N_5737,N_4325,N_4334);
and U5738 (N_5738,N_4029,N_4854);
and U5739 (N_5739,N_4300,N_4867);
and U5740 (N_5740,N_4877,N_4236);
and U5741 (N_5741,N_4524,N_4260);
xnor U5742 (N_5742,N_4289,N_4834);
nor U5743 (N_5743,N_4248,N_4860);
and U5744 (N_5744,N_4812,N_4293);
and U5745 (N_5745,N_4091,N_4632);
and U5746 (N_5746,N_4037,N_4161);
and U5747 (N_5747,N_4202,N_4369);
nor U5748 (N_5748,N_4588,N_4795);
nor U5749 (N_5749,N_4082,N_4572);
nand U5750 (N_5750,N_4930,N_4905);
nor U5751 (N_5751,N_4496,N_4075);
nor U5752 (N_5752,N_4478,N_4039);
nor U5753 (N_5753,N_4858,N_4926);
nor U5754 (N_5754,N_4820,N_4773);
nor U5755 (N_5755,N_4967,N_4488);
and U5756 (N_5756,N_4053,N_4000);
and U5757 (N_5757,N_4252,N_4572);
or U5758 (N_5758,N_4886,N_4020);
and U5759 (N_5759,N_4840,N_4054);
nor U5760 (N_5760,N_4971,N_4577);
nor U5761 (N_5761,N_4710,N_4105);
xor U5762 (N_5762,N_4823,N_4198);
or U5763 (N_5763,N_4198,N_4352);
nor U5764 (N_5764,N_4407,N_4803);
and U5765 (N_5765,N_4109,N_4690);
or U5766 (N_5766,N_4308,N_4515);
and U5767 (N_5767,N_4346,N_4790);
and U5768 (N_5768,N_4490,N_4605);
nor U5769 (N_5769,N_4545,N_4903);
or U5770 (N_5770,N_4163,N_4159);
nor U5771 (N_5771,N_4993,N_4320);
nand U5772 (N_5772,N_4286,N_4492);
nand U5773 (N_5773,N_4177,N_4617);
nand U5774 (N_5774,N_4895,N_4965);
or U5775 (N_5775,N_4330,N_4320);
or U5776 (N_5776,N_4950,N_4076);
and U5777 (N_5777,N_4998,N_4453);
nand U5778 (N_5778,N_4421,N_4207);
nor U5779 (N_5779,N_4937,N_4070);
nor U5780 (N_5780,N_4382,N_4784);
or U5781 (N_5781,N_4991,N_4333);
nand U5782 (N_5782,N_4111,N_4248);
or U5783 (N_5783,N_4079,N_4219);
nor U5784 (N_5784,N_4788,N_4726);
nand U5785 (N_5785,N_4549,N_4068);
nor U5786 (N_5786,N_4155,N_4245);
or U5787 (N_5787,N_4380,N_4178);
nand U5788 (N_5788,N_4149,N_4669);
and U5789 (N_5789,N_4381,N_4447);
nor U5790 (N_5790,N_4447,N_4200);
nand U5791 (N_5791,N_4688,N_4788);
nor U5792 (N_5792,N_4770,N_4509);
nor U5793 (N_5793,N_4562,N_4475);
and U5794 (N_5794,N_4167,N_4415);
nor U5795 (N_5795,N_4460,N_4638);
or U5796 (N_5796,N_4509,N_4607);
nor U5797 (N_5797,N_4300,N_4794);
or U5798 (N_5798,N_4553,N_4813);
and U5799 (N_5799,N_4812,N_4068);
nor U5800 (N_5800,N_4604,N_4941);
or U5801 (N_5801,N_4129,N_4664);
and U5802 (N_5802,N_4184,N_4545);
nand U5803 (N_5803,N_4775,N_4454);
or U5804 (N_5804,N_4011,N_4154);
nor U5805 (N_5805,N_4895,N_4095);
nor U5806 (N_5806,N_4203,N_4495);
and U5807 (N_5807,N_4298,N_4281);
nor U5808 (N_5808,N_4198,N_4887);
nand U5809 (N_5809,N_4599,N_4279);
nand U5810 (N_5810,N_4728,N_4666);
nand U5811 (N_5811,N_4486,N_4067);
and U5812 (N_5812,N_4088,N_4433);
nand U5813 (N_5813,N_4706,N_4033);
nand U5814 (N_5814,N_4514,N_4721);
or U5815 (N_5815,N_4358,N_4791);
nor U5816 (N_5816,N_4584,N_4311);
nor U5817 (N_5817,N_4404,N_4551);
and U5818 (N_5818,N_4264,N_4663);
or U5819 (N_5819,N_4121,N_4834);
and U5820 (N_5820,N_4318,N_4227);
xnor U5821 (N_5821,N_4950,N_4747);
nor U5822 (N_5822,N_4842,N_4290);
nor U5823 (N_5823,N_4445,N_4786);
nand U5824 (N_5824,N_4481,N_4562);
nor U5825 (N_5825,N_4073,N_4497);
xnor U5826 (N_5826,N_4039,N_4989);
nor U5827 (N_5827,N_4160,N_4317);
or U5828 (N_5828,N_4018,N_4745);
and U5829 (N_5829,N_4417,N_4088);
nor U5830 (N_5830,N_4478,N_4235);
nor U5831 (N_5831,N_4028,N_4890);
and U5832 (N_5832,N_4608,N_4980);
and U5833 (N_5833,N_4198,N_4687);
and U5834 (N_5834,N_4453,N_4936);
and U5835 (N_5835,N_4204,N_4339);
nor U5836 (N_5836,N_4601,N_4914);
nor U5837 (N_5837,N_4731,N_4208);
and U5838 (N_5838,N_4307,N_4091);
and U5839 (N_5839,N_4459,N_4708);
nor U5840 (N_5840,N_4477,N_4376);
and U5841 (N_5841,N_4008,N_4408);
and U5842 (N_5842,N_4719,N_4643);
and U5843 (N_5843,N_4744,N_4416);
or U5844 (N_5844,N_4340,N_4254);
or U5845 (N_5845,N_4266,N_4123);
nand U5846 (N_5846,N_4198,N_4394);
or U5847 (N_5847,N_4747,N_4644);
or U5848 (N_5848,N_4089,N_4108);
or U5849 (N_5849,N_4719,N_4456);
or U5850 (N_5850,N_4823,N_4852);
nor U5851 (N_5851,N_4412,N_4261);
nand U5852 (N_5852,N_4872,N_4597);
or U5853 (N_5853,N_4029,N_4653);
or U5854 (N_5854,N_4159,N_4480);
nand U5855 (N_5855,N_4030,N_4559);
nor U5856 (N_5856,N_4563,N_4805);
and U5857 (N_5857,N_4855,N_4929);
and U5858 (N_5858,N_4718,N_4014);
and U5859 (N_5859,N_4766,N_4243);
or U5860 (N_5860,N_4469,N_4387);
and U5861 (N_5861,N_4613,N_4902);
nand U5862 (N_5862,N_4033,N_4629);
nor U5863 (N_5863,N_4125,N_4602);
nand U5864 (N_5864,N_4810,N_4281);
or U5865 (N_5865,N_4567,N_4318);
nand U5866 (N_5866,N_4276,N_4315);
and U5867 (N_5867,N_4414,N_4012);
or U5868 (N_5868,N_4338,N_4799);
nand U5869 (N_5869,N_4506,N_4670);
nor U5870 (N_5870,N_4063,N_4133);
nand U5871 (N_5871,N_4847,N_4415);
nor U5872 (N_5872,N_4786,N_4501);
and U5873 (N_5873,N_4188,N_4653);
nand U5874 (N_5874,N_4483,N_4778);
nor U5875 (N_5875,N_4884,N_4446);
and U5876 (N_5876,N_4751,N_4252);
or U5877 (N_5877,N_4650,N_4173);
and U5878 (N_5878,N_4441,N_4997);
nor U5879 (N_5879,N_4873,N_4470);
or U5880 (N_5880,N_4588,N_4906);
and U5881 (N_5881,N_4636,N_4633);
and U5882 (N_5882,N_4102,N_4794);
or U5883 (N_5883,N_4982,N_4844);
or U5884 (N_5884,N_4856,N_4585);
nand U5885 (N_5885,N_4033,N_4572);
xnor U5886 (N_5886,N_4901,N_4948);
nand U5887 (N_5887,N_4619,N_4706);
or U5888 (N_5888,N_4860,N_4605);
and U5889 (N_5889,N_4912,N_4388);
nand U5890 (N_5890,N_4725,N_4060);
and U5891 (N_5891,N_4391,N_4611);
nand U5892 (N_5892,N_4616,N_4054);
and U5893 (N_5893,N_4724,N_4102);
nor U5894 (N_5894,N_4737,N_4763);
nor U5895 (N_5895,N_4888,N_4193);
nor U5896 (N_5896,N_4438,N_4286);
nor U5897 (N_5897,N_4828,N_4576);
and U5898 (N_5898,N_4136,N_4142);
or U5899 (N_5899,N_4867,N_4354);
and U5900 (N_5900,N_4122,N_4714);
nor U5901 (N_5901,N_4440,N_4903);
nand U5902 (N_5902,N_4275,N_4133);
and U5903 (N_5903,N_4659,N_4118);
and U5904 (N_5904,N_4335,N_4190);
nand U5905 (N_5905,N_4305,N_4060);
nand U5906 (N_5906,N_4913,N_4183);
and U5907 (N_5907,N_4389,N_4173);
or U5908 (N_5908,N_4451,N_4384);
nand U5909 (N_5909,N_4418,N_4984);
nand U5910 (N_5910,N_4292,N_4371);
xor U5911 (N_5911,N_4725,N_4102);
or U5912 (N_5912,N_4555,N_4429);
nand U5913 (N_5913,N_4770,N_4373);
nand U5914 (N_5914,N_4537,N_4569);
nor U5915 (N_5915,N_4878,N_4148);
nor U5916 (N_5916,N_4746,N_4738);
nor U5917 (N_5917,N_4626,N_4674);
and U5918 (N_5918,N_4169,N_4037);
nand U5919 (N_5919,N_4395,N_4757);
nand U5920 (N_5920,N_4687,N_4239);
and U5921 (N_5921,N_4387,N_4033);
nor U5922 (N_5922,N_4626,N_4595);
or U5923 (N_5923,N_4099,N_4028);
nand U5924 (N_5924,N_4552,N_4058);
nor U5925 (N_5925,N_4824,N_4227);
or U5926 (N_5926,N_4456,N_4713);
and U5927 (N_5927,N_4258,N_4653);
nand U5928 (N_5928,N_4358,N_4735);
nand U5929 (N_5929,N_4140,N_4998);
nor U5930 (N_5930,N_4144,N_4848);
and U5931 (N_5931,N_4275,N_4700);
nor U5932 (N_5932,N_4496,N_4085);
nand U5933 (N_5933,N_4424,N_4241);
nand U5934 (N_5934,N_4631,N_4256);
or U5935 (N_5935,N_4236,N_4677);
or U5936 (N_5936,N_4282,N_4144);
nand U5937 (N_5937,N_4527,N_4427);
nor U5938 (N_5938,N_4800,N_4028);
nor U5939 (N_5939,N_4784,N_4656);
and U5940 (N_5940,N_4840,N_4699);
nor U5941 (N_5941,N_4951,N_4104);
or U5942 (N_5942,N_4240,N_4770);
or U5943 (N_5943,N_4618,N_4276);
or U5944 (N_5944,N_4502,N_4465);
and U5945 (N_5945,N_4527,N_4716);
nor U5946 (N_5946,N_4582,N_4992);
or U5947 (N_5947,N_4223,N_4507);
nor U5948 (N_5948,N_4614,N_4728);
nand U5949 (N_5949,N_4014,N_4488);
nand U5950 (N_5950,N_4842,N_4139);
nor U5951 (N_5951,N_4958,N_4700);
nand U5952 (N_5952,N_4164,N_4094);
nand U5953 (N_5953,N_4437,N_4002);
and U5954 (N_5954,N_4403,N_4998);
and U5955 (N_5955,N_4141,N_4257);
nand U5956 (N_5956,N_4519,N_4912);
nand U5957 (N_5957,N_4525,N_4957);
or U5958 (N_5958,N_4011,N_4547);
xnor U5959 (N_5959,N_4555,N_4006);
or U5960 (N_5960,N_4099,N_4322);
xor U5961 (N_5961,N_4429,N_4534);
and U5962 (N_5962,N_4757,N_4303);
or U5963 (N_5963,N_4399,N_4378);
or U5964 (N_5964,N_4279,N_4185);
nand U5965 (N_5965,N_4303,N_4243);
nand U5966 (N_5966,N_4809,N_4985);
nand U5967 (N_5967,N_4763,N_4713);
nor U5968 (N_5968,N_4976,N_4961);
nand U5969 (N_5969,N_4743,N_4997);
nand U5970 (N_5970,N_4748,N_4777);
or U5971 (N_5971,N_4887,N_4554);
nor U5972 (N_5972,N_4776,N_4177);
nor U5973 (N_5973,N_4713,N_4188);
or U5974 (N_5974,N_4372,N_4499);
nand U5975 (N_5975,N_4373,N_4063);
nor U5976 (N_5976,N_4594,N_4883);
or U5977 (N_5977,N_4995,N_4926);
or U5978 (N_5978,N_4073,N_4986);
and U5979 (N_5979,N_4574,N_4554);
and U5980 (N_5980,N_4089,N_4306);
or U5981 (N_5981,N_4752,N_4340);
or U5982 (N_5982,N_4652,N_4171);
or U5983 (N_5983,N_4496,N_4701);
and U5984 (N_5984,N_4771,N_4147);
xor U5985 (N_5985,N_4023,N_4590);
nor U5986 (N_5986,N_4956,N_4327);
and U5987 (N_5987,N_4104,N_4908);
nand U5988 (N_5988,N_4915,N_4360);
nor U5989 (N_5989,N_4155,N_4264);
nand U5990 (N_5990,N_4666,N_4533);
and U5991 (N_5991,N_4057,N_4615);
and U5992 (N_5992,N_4607,N_4056);
or U5993 (N_5993,N_4416,N_4287);
and U5994 (N_5994,N_4582,N_4700);
or U5995 (N_5995,N_4251,N_4720);
and U5996 (N_5996,N_4662,N_4743);
or U5997 (N_5997,N_4633,N_4655);
nor U5998 (N_5998,N_4725,N_4447);
nor U5999 (N_5999,N_4854,N_4951);
and U6000 (N_6000,N_5328,N_5918);
nand U6001 (N_6001,N_5360,N_5000);
and U6002 (N_6002,N_5712,N_5057);
nand U6003 (N_6003,N_5789,N_5771);
nand U6004 (N_6004,N_5669,N_5302);
and U6005 (N_6005,N_5923,N_5678);
or U6006 (N_6006,N_5530,N_5810);
nand U6007 (N_6007,N_5824,N_5286);
or U6008 (N_6008,N_5606,N_5689);
nor U6009 (N_6009,N_5886,N_5751);
or U6010 (N_6010,N_5592,N_5571);
or U6011 (N_6011,N_5668,N_5921);
or U6012 (N_6012,N_5765,N_5096);
or U6013 (N_6013,N_5058,N_5183);
nand U6014 (N_6014,N_5877,N_5821);
and U6015 (N_6015,N_5456,N_5152);
and U6016 (N_6016,N_5763,N_5777);
nand U6017 (N_6017,N_5326,N_5797);
nand U6018 (N_6018,N_5598,N_5186);
nand U6019 (N_6019,N_5185,N_5426);
nand U6020 (N_6020,N_5820,N_5964);
and U6021 (N_6021,N_5139,N_5078);
and U6022 (N_6022,N_5263,N_5958);
nor U6023 (N_6023,N_5221,N_5550);
or U6024 (N_6024,N_5212,N_5049);
or U6025 (N_6025,N_5093,N_5228);
xnor U6026 (N_6026,N_5932,N_5573);
or U6027 (N_6027,N_5252,N_5053);
nor U6028 (N_6028,N_5738,N_5052);
nor U6029 (N_6029,N_5397,N_5579);
and U6030 (N_6030,N_5853,N_5858);
nor U6031 (N_6031,N_5706,N_5545);
or U6032 (N_6032,N_5719,N_5366);
nor U6033 (N_6033,N_5816,N_5452);
nor U6034 (N_6034,N_5103,N_5213);
and U6035 (N_6035,N_5187,N_5946);
nor U6036 (N_6036,N_5071,N_5069);
and U6037 (N_6037,N_5140,N_5622);
or U6038 (N_6038,N_5233,N_5645);
nand U6039 (N_6039,N_5753,N_5723);
and U6040 (N_6040,N_5247,N_5846);
and U6041 (N_6041,N_5350,N_5818);
nor U6042 (N_6042,N_5888,N_5418);
or U6043 (N_6043,N_5474,N_5640);
or U6044 (N_6044,N_5525,N_5405);
and U6045 (N_6045,N_5192,N_5811);
nor U6046 (N_6046,N_5055,N_5812);
and U6047 (N_6047,N_5108,N_5799);
or U6048 (N_6048,N_5778,N_5869);
or U6049 (N_6049,N_5784,N_5989);
nand U6050 (N_6050,N_5037,N_5859);
nand U6051 (N_6051,N_5515,N_5179);
nor U6052 (N_6052,N_5945,N_5014);
nand U6053 (N_6053,N_5922,N_5795);
or U6054 (N_6054,N_5936,N_5218);
and U6055 (N_6055,N_5968,N_5411);
and U6056 (N_6056,N_5477,N_5283);
and U6057 (N_6057,N_5240,N_5908);
or U6058 (N_6058,N_5162,N_5942);
nand U6059 (N_6059,N_5051,N_5295);
nor U6060 (N_6060,N_5834,N_5660);
nor U6061 (N_6061,N_5632,N_5806);
and U6062 (N_6062,N_5214,N_5371);
or U6063 (N_6063,N_5574,N_5601);
nor U6064 (N_6064,N_5190,N_5017);
and U6065 (N_6065,N_5759,N_5972);
and U6066 (N_6066,N_5890,N_5184);
nand U6067 (N_6067,N_5315,N_5408);
nor U6068 (N_6068,N_5843,N_5102);
and U6069 (N_6069,N_5840,N_5803);
and U6070 (N_6070,N_5073,N_5349);
and U6071 (N_6071,N_5896,N_5265);
nand U6072 (N_6072,N_5623,N_5424);
or U6073 (N_6073,N_5343,N_5937);
nand U6074 (N_6074,N_5458,N_5112);
and U6075 (N_6075,N_5457,N_5624);
or U6076 (N_6076,N_5100,N_5493);
and U6077 (N_6077,N_5970,N_5851);
nand U6078 (N_6078,N_5798,N_5384);
nor U6079 (N_6079,N_5992,N_5871);
nand U6080 (N_6080,N_5375,N_5904);
or U6081 (N_6081,N_5654,N_5650);
or U6082 (N_6082,N_5234,N_5651);
nor U6083 (N_6083,N_5159,N_5526);
or U6084 (N_6084,N_5508,N_5711);
nor U6085 (N_6085,N_5420,N_5437);
or U6086 (N_6086,N_5898,N_5066);
or U6087 (N_6087,N_5012,N_5345);
nor U6088 (N_6088,N_5196,N_5781);
nor U6089 (N_6089,N_5892,N_5236);
nand U6090 (N_6090,N_5098,N_5665);
nand U6091 (N_6091,N_5586,N_5262);
or U6092 (N_6092,N_5064,N_5273);
nand U6093 (N_6093,N_5661,N_5451);
and U6094 (N_6094,N_5311,N_5878);
or U6095 (N_6095,N_5325,N_5754);
or U6096 (N_6096,N_5741,N_5676);
nand U6097 (N_6097,N_5626,N_5028);
and U6098 (N_6098,N_5322,N_5143);
or U6099 (N_6099,N_5721,N_5459);
nor U6100 (N_6100,N_5925,N_5863);
or U6101 (N_6101,N_5591,N_5557);
and U6102 (N_6102,N_5796,N_5607);
nand U6103 (N_6103,N_5074,N_5617);
or U6104 (N_6104,N_5895,N_5001);
nor U6105 (N_6105,N_5046,N_5667);
and U6106 (N_6106,N_5561,N_5841);
or U6107 (N_6107,N_5903,N_5340);
and U6108 (N_6108,N_5900,N_5897);
and U6109 (N_6109,N_5955,N_5278);
nor U6110 (N_6110,N_5790,N_5547);
and U6111 (N_6111,N_5518,N_5764);
xor U6112 (N_6112,N_5177,N_5410);
and U6113 (N_6113,N_5377,N_5612);
nand U6114 (N_6114,N_5484,N_5739);
xor U6115 (N_6115,N_5572,N_5804);
nand U6116 (N_6116,N_5031,N_5709);
and U6117 (N_6117,N_5831,N_5267);
nand U6118 (N_6118,N_5730,N_5308);
or U6119 (N_6119,N_5695,N_5376);
nor U6120 (N_6120,N_5216,N_5982);
nand U6121 (N_6121,N_5027,N_5774);
and U6122 (N_6122,N_5581,N_5748);
nand U6123 (N_6123,N_5680,N_5829);
nand U6124 (N_6124,N_5210,N_5913);
nor U6125 (N_6125,N_5346,N_5994);
nand U6126 (N_6126,N_5542,N_5181);
nor U6127 (N_6127,N_5422,N_5911);
and U6128 (N_6128,N_5427,N_5113);
nand U6129 (N_6129,N_5867,N_5173);
and U6130 (N_6130,N_5081,N_5835);
nand U6131 (N_6131,N_5095,N_5250);
nor U6132 (N_6132,N_5365,N_5060);
or U6133 (N_6133,N_5121,N_5337);
nor U6134 (N_6134,N_5373,N_5637);
and U6135 (N_6135,N_5447,N_5658);
nor U6136 (N_6136,N_5380,N_5125);
and U6137 (N_6137,N_5063,N_5567);
or U6138 (N_6138,N_5013,N_5745);
nand U6139 (N_6139,N_5387,N_5909);
or U6140 (N_6140,N_5011,N_5111);
nand U6141 (N_6141,N_5020,N_5733);
or U6142 (N_6142,N_5865,N_5164);
and U6143 (N_6143,N_5023,N_5110);
nand U6144 (N_6144,N_5061,N_5313);
nor U6145 (N_6145,N_5707,N_5756);
or U6146 (N_6146,N_5644,N_5495);
and U6147 (N_6147,N_5643,N_5305);
nand U6148 (N_6148,N_5423,N_5298);
nor U6149 (N_6149,N_5593,N_5696);
and U6150 (N_6150,N_5649,N_5987);
nor U6151 (N_6151,N_5282,N_5604);
and U6152 (N_6152,N_5594,N_5516);
nor U6153 (N_6153,N_5468,N_5347);
or U6154 (N_6154,N_5862,N_5156);
and U6155 (N_6155,N_5421,N_5438);
nand U6156 (N_6156,N_5091,N_5522);
nand U6157 (N_6157,N_5692,N_5761);
nor U6158 (N_6158,N_5779,N_5808);
nor U6159 (N_6159,N_5901,N_5770);
and U6160 (N_6160,N_5587,N_5406);
nor U6161 (N_6161,N_5681,N_5439);
or U6162 (N_6162,N_5646,N_5442);
nor U6163 (N_6163,N_5369,N_5524);
nand U6164 (N_6164,N_5016,N_5155);
nor U6165 (N_6165,N_5407,N_5294);
or U6166 (N_6166,N_5523,N_5157);
nand U6167 (N_6167,N_5540,N_5342);
nand U6168 (N_6168,N_5819,N_5035);
nor U6169 (N_6169,N_5225,N_5564);
or U6170 (N_6170,N_5202,N_5613);
nand U6171 (N_6171,N_5092,N_5630);
nor U6172 (N_6172,N_5032,N_5166);
and U6173 (N_6173,N_5448,N_5833);
or U6174 (N_6174,N_5967,N_5735);
nand U6175 (N_6175,N_5101,N_5507);
nor U6176 (N_6176,N_5847,N_5755);
nand U6177 (N_6177,N_5289,N_5478);
nor U6178 (N_6178,N_5450,N_5194);
and U6179 (N_6179,N_5631,N_5232);
nor U6180 (N_6180,N_5168,N_5090);
or U6181 (N_6181,N_5546,N_5852);
and U6182 (N_6182,N_5677,N_5076);
or U6183 (N_6183,N_5544,N_5389);
nor U6184 (N_6184,N_5082,N_5512);
and U6185 (N_6185,N_5527,N_5310);
and U6186 (N_6186,N_5378,N_5555);
and U6187 (N_6187,N_5576,N_5290);
and U6188 (N_6188,N_5268,N_5191);
nand U6189 (N_6189,N_5722,N_5473);
or U6190 (N_6190,N_5562,N_5995);
and U6191 (N_6191,N_5568,N_5978);
or U6192 (N_6192,N_5956,N_5400);
or U6193 (N_6193,N_5021,N_5171);
nand U6194 (N_6194,N_5984,N_5940);
and U6195 (N_6195,N_5425,N_5368);
nor U6196 (N_6196,N_5024,N_5827);
nand U6197 (N_6197,N_5610,N_5705);
and U6198 (N_6198,N_5953,N_5698);
nor U6199 (N_6199,N_5237,N_5868);
nand U6200 (N_6200,N_5255,N_5463);
and U6201 (N_6201,N_5548,N_5131);
nand U6202 (N_6202,N_5435,N_5099);
nor U6203 (N_6203,N_5980,N_5404);
nand U6204 (N_6204,N_5396,N_5963);
nand U6205 (N_6205,N_5211,N_5894);
nand U6206 (N_6206,N_5618,N_5876);
and U6207 (N_6207,N_5075,N_5726);
nor U6208 (N_6208,N_5498,N_5879);
nand U6209 (N_6209,N_5907,N_5792);
and U6210 (N_6210,N_5022,N_5386);
nor U6211 (N_6211,N_5485,N_5483);
and U6212 (N_6212,N_5822,N_5358);
and U6213 (N_6213,N_5331,N_5655);
nand U6214 (N_6214,N_5446,N_5089);
or U6215 (N_6215,N_5672,N_5928);
and U6216 (N_6216,N_5204,N_5409);
and U6217 (N_6217,N_5172,N_5319);
or U6218 (N_6218,N_5416,N_5570);
nor U6219 (N_6219,N_5244,N_5971);
and U6220 (N_6220,N_5899,N_5067);
or U6221 (N_6221,N_5614,N_5511);
or U6222 (N_6222,N_5379,N_5575);
nand U6223 (N_6223,N_5150,N_5339);
and U6224 (N_6224,N_5433,N_5817);
or U6225 (N_6225,N_5532,N_5398);
nor U6226 (N_6226,N_5961,N_5284);
or U6227 (N_6227,N_5281,N_5619);
nand U6228 (N_6228,N_5935,N_5264);
or U6229 (N_6229,N_5401,N_5521);
or U6230 (N_6230,N_5809,N_5704);
nand U6231 (N_6231,N_5077,N_5415);
and U6232 (N_6232,N_5916,N_5383);
or U6233 (N_6233,N_5201,N_5702);
nand U6234 (N_6234,N_5837,N_5039);
nor U6235 (N_6235,N_5266,N_5359);
or U6236 (N_6236,N_5679,N_5080);
and U6237 (N_6237,N_5481,N_5788);
nand U6238 (N_6238,N_5627,N_5927);
or U6239 (N_6239,N_5285,N_5697);
nand U6240 (N_6240,N_5043,N_5549);
nor U6241 (N_6241,N_5030,N_5390);
and U6242 (N_6242,N_5222,N_5374);
nand U6243 (N_6243,N_5732,N_5563);
nor U6244 (N_6244,N_5513,N_5634);
and U6245 (N_6245,N_5716,N_5475);
and U6246 (N_6246,N_5314,N_5559);
and U6247 (N_6247,N_5123,N_5487);
and U6248 (N_6248,N_5083,N_5553);
or U6249 (N_6249,N_5154,N_5582);
nand U6250 (N_6250,N_5556,N_5009);
nor U6251 (N_6251,N_5949,N_5496);
and U6252 (N_6252,N_5494,N_5977);
nand U6253 (N_6253,N_5957,N_5850);
nand U6254 (N_6254,N_5392,N_5275);
and U6255 (N_6255,N_5757,N_5905);
nand U6256 (N_6256,N_5462,N_5749);
or U6257 (N_6257,N_5258,N_5472);
nor U6258 (N_6258,N_5208,N_5832);
nor U6259 (N_6259,N_5490,N_5580);
and U6260 (N_6260,N_5455,N_5536);
or U6261 (N_6261,N_5686,N_5363);
nor U6262 (N_6262,N_5119,N_5828);
and U6263 (N_6263,N_5174,N_5167);
or U6264 (N_6264,N_5151,N_5460);
nand U6265 (N_6265,N_5595,N_5019);
nor U6266 (N_6266,N_5324,N_5966);
nand U6267 (N_6267,N_5394,N_5312);
nand U6268 (N_6268,N_5773,N_5094);
and U6269 (N_6269,N_5002,N_5766);
and U6270 (N_6270,N_5710,N_5120);
and U6271 (N_6271,N_5969,N_5038);
nand U6272 (N_6272,N_5772,N_5332);
or U6273 (N_6273,N_5974,N_5588);
nand U6274 (N_6274,N_5694,N_5551);
or U6275 (N_6275,N_5577,N_5983);
or U6276 (N_6276,N_5033,N_5912);
nand U6277 (N_6277,N_5417,N_5029);
or U6278 (N_6278,N_5520,N_5443);
nand U6279 (N_6279,N_5537,N_5178);
or U6280 (N_6280,N_5133,N_5117);
or U6281 (N_6281,N_5261,N_5952);
nand U6282 (N_6282,N_5688,N_5857);
and U6283 (N_6283,N_5464,N_5533);
or U6284 (N_6284,N_5599,N_5480);
or U6285 (N_6285,N_5509,N_5440);
and U6286 (N_6286,N_5620,N_5849);
and U6287 (N_6287,N_5238,N_5354);
or U6288 (N_6288,N_5048,N_5137);
nor U6289 (N_6289,N_5998,N_5200);
and U6290 (N_6290,N_5391,N_5006);
nor U6291 (N_6291,N_5758,N_5670);
or U6292 (N_6292,N_5501,N_5056);
nand U6293 (N_6293,N_5287,N_5780);
nand U6294 (N_6294,N_5786,N_5589);
and U6295 (N_6295,N_5025,N_5445);
nor U6296 (N_6296,N_5638,N_5736);
or U6297 (N_6297,N_5260,N_5647);
nor U6298 (N_6298,N_5303,N_5794);
or U6299 (N_6299,N_5541,N_5335);
and U6300 (N_6300,N_5684,N_5554);
or U6301 (N_6301,N_5469,N_5744);
nor U6302 (N_6302,N_5235,N_5296);
or U6303 (N_6303,N_5505,N_5641);
and U6304 (N_6304,N_5492,N_5466);
nand U6305 (N_6305,N_5118,N_5583);
nor U6306 (N_6306,N_5882,N_5018);
nor U6307 (N_6307,N_5656,N_5915);
or U6308 (N_6308,N_5737,N_5388);
or U6309 (N_6309,N_5253,N_5217);
nand U6310 (N_6310,N_5207,N_5685);
and U6311 (N_6311,N_5403,N_5954);
nor U6312 (N_6312,N_5044,N_5747);
or U6313 (N_6313,N_5815,N_5881);
nor U6314 (N_6314,N_5317,N_5395);
or U6315 (N_6315,N_5944,N_5615);
or U6316 (N_6316,N_5539,N_5902);
nand U6317 (N_6317,N_5413,N_5997);
nand U6318 (N_6318,N_5514,N_5889);
or U6319 (N_6319,N_5291,N_5097);
nor U6320 (N_6320,N_5700,N_5441);
nor U6321 (N_6321,N_5136,N_5652);
or U6322 (N_6322,N_5301,N_5045);
nand U6323 (N_6323,N_5965,N_5239);
or U6324 (N_6324,N_5402,N_5249);
nand U6325 (N_6325,N_5323,N_5979);
and U6326 (N_6326,N_5115,N_5436);
and U6327 (N_6327,N_5693,N_5454);
nor U6328 (N_6328,N_5584,N_5434);
or U6329 (N_6329,N_5662,N_5768);
nor U6330 (N_6330,N_5288,N_5951);
and U6331 (N_6331,N_5813,N_5625);
or U6332 (N_6332,N_5203,N_5504);
nor U6333 (N_6333,N_5683,N_5642);
nor U6334 (N_6334,N_5341,N_5306);
nand U6335 (N_6335,N_5746,N_5875);
and U6336 (N_6336,N_5146,N_5334);
or U6337 (N_6337,N_5842,N_5621);
nand U6338 (N_6338,N_5947,N_5036);
nor U6339 (N_6339,N_5578,N_5412);
nor U6340 (N_6340,N_5034,N_5883);
or U6341 (N_6341,N_5791,N_5141);
and U6342 (N_6342,N_5930,N_5560);
nand U6343 (N_6343,N_5750,N_5393);
or U6344 (N_6344,N_5276,N_5552);
and U6345 (N_6345,N_5482,N_5318);
nor U6346 (N_6346,N_5351,N_5010);
and U6347 (N_6347,N_5499,N_5189);
and U6348 (N_6348,N_5175,N_5991);
nor U6349 (N_6349,N_5742,N_5381);
nor U6350 (N_6350,N_5534,N_5348);
nor U6351 (N_6351,N_5361,N_5767);
and U6352 (N_6352,N_5657,N_5729);
nand U6353 (N_6353,N_5919,N_5648);
nand U6354 (N_6354,N_5040,N_5470);
or U6355 (N_6355,N_5135,N_5535);
nand U6356 (N_6356,N_5251,N_5144);
nor U6357 (N_6357,N_5924,N_5715);
nand U6358 (N_6358,N_5274,N_5673);
nor U6359 (N_6359,N_5243,N_5962);
and U6360 (N_6360,N_5338,N_5370);
nand U6361 (N_6361,N_5107,N_5223);
and U6362 (N_6362,N_5042,N_5372);
nor U6363 (N_6363,N_5206,N_5116);
and U6364 (N_6364,N_5050,N_5981);
and U6365 (N_6365,N_5793,N_5703);
and U6366 (N_6366,N_5941,N_5430);
or U6367 (N_6367,N_5219,N_5724);
nor U6368 (N_6368,N_5356,N_5939);
or U6369 (N_6369,N_5906,N_5713);
nand U6370 (N_6370,N_5124,N_5429);
or U6371 (N_6371,N_5227,N_5752);
nand U6372 (N_6372,N_5209,N_5866);
and U6373 (N_6373,N_5259,N_5874);
and U6374 (N_6374,N_5873,N_5142);
and U6375 (N_6375,N_5887,N_5419);
and U6376 (N_6376,N_5479,N_5510);
or U6377 (N_6377,N_5728,N_5926);
nor U6378 (N_6378,N_5079,N_5605);
or U6379 (N_6379,N_5256,N_5344);
and U6380 (N_6380,N_5432,N_5633);
nor U6381 (N_6381,N_5182,N_5199);
or U6382 (N_6382,N_5280,N_5149);
and U6383 (N_6383,N_5985,N_5254);
nand U6384 (N_6384,N_5976,N_5864);
nand U6385 (N_6385,N_5461,N_5176);
or U6386 (N_6386,N_5609,N_5823);
nor U6387 (N_6387,N_5059,N_5165);
or U6388 (N_6388,N_5327,N_5148);
nand U6389 (N_6389,N_5727,N_5128);
nor U6390 (N_6390,N_5245,N_5127);
nand U6391 (N_6391,N_5893,N_5153);
and U6392 (N_6392,N_5861,N_5585);
and U6393 (N_6393,N_5708,N_5565);
nor U6394 (N_6394,N_5762,N_5986);
and U6395 (N_6395,N_5453,N_5362);
nor U6396 (N_6396,N_5465,N_5960);
or U6397 (N_6397,N_5558,N_5844);
or U6398 (N_6398,N_5333,N_5336);
nor U6399 (N_6399,N_5329,N_5782);
or U6400 (N_6400,N_5848,N_5805);
or U6401 (N_6401,N_5353,N_5718);
nand U6402 (N_6402,N_5538,N_5004);
and U6403 (N_6403,N_5855,N_5220);
and U6404 (N_6404,N_5357,N_5990);
and U6405 (N_6405,N_5880,N_5003);
nor U6406 (N_6406,N_5015,N_5814);
nand U6407 (N_6407,N_5352,N_5528);
or U6408 (N_6408,N_5047,N_5787);
and U6409 (N_6409,N_5699,N_5007);
nand U6410 (N_6410,N_5008,N_5114);
or U6411 (N_6411,N_5731,N_5943);
nand U6412 (N_6412,N_5316,N_5215);
and U6413 (N_6413,N_5775,N_5134);
and U6414 (N_6414,N_5543,N_5271);
nand U6415 (N_6415,N_5743,N_5449);
and U6416 (N_6416,N_5917,N_5230);
or U6417 (N_6417,N_5444,N_5659);
and U6418 (N_6418,N_5734,N_5740);
nand U6419 (N_6419,N_5872,N_5367);
and U6420 (N_6420,N_5664,N_5500);
or U6421 (N_6421,N_5870,N_5860);
or U6422 (N_6422,N_5106,N_5297);
nand U6423 (N_6423,N_5170,N_5720);
or U6424 (N_6424,N_5597,N_5825);
nor U6425 (N_6425,N_5725,N_5938);
and U6426 (N_6426,N_5087,N_5065);
nor U6427 (N_6427,N_5330,N_5180);
or U6428 (N_6428,N_5503,N_5226);
or U6429 (N_6429,N_5355,N_5529);
or U6430 (N_6430,N_5590,N_5636);
or U6431 (N_6431,N_5169,N_5959);
xnor U6432 (N_6432,N_5999,N_5205);
nor U6433 (N_6433,N_5663,N_5800);
nand U6434 (N_6434,N_5611,N_5769);
nor U6435 (N_6435,N_5973,N_5304);
nor U6436 (N_6436,N_5428,N_5130);
nand U6437 (N_6437,N_5242,N_5062);
and U6438 (N_6438,N_5783,N_5502);
xor U6439 (N_6439,N_5070,N_5785);
or U6440 (N_6440,N_5884,N_5671);
and U6441 (N_6441,N_5299,N_5596);
nor U6442 (N_6442,N_5488,N_5188);
nand U6443 (N_6443,N_5229,N_5193);
and U6444 (N_6444,N_5629,N_5929);
and U6445 (N_6445,N_5602,N_5603);
nor U6446 (N_6446,N_5224,N_5414);
nor U6447 (N_6447,N_5801,N_5231);
or U6448 (N_6448,N_5802,N_5497);
or U6449 (N_6449,N_5653,N_5320);
and U6450 (N_6450,N_5910,N_5854);
nand U6451 (N_6451,N_5309,N_5293);
nand U6452 (N_6452,N_5839,N_5005);
and U6453 (N_6453,N_5241,N_5160);
and U6454 (N_6454,N_5701,N_5147);
and U6455 (N_6455,N_5988,N_5687);
nor U6456 (N_6456,N_5195,N_5891);
nor U6457 (N_6457,N_5068,N_5608);
nand U6458 (N_6458,N_5072,N_5856);
and U6459 (N_6459,N_5257,N_5085);
nor U6460 (N_6460,N_5138,N_5682);
and U6461 (N_6461,N_5666,N_5307);
nor U6462 (N_6462,N_5675,N_5531);
nor U6463 (N_6463,N_5277,N_5517);
nor U6464 (N_6464,N_5914,N_5122);
and U6465 (N_6465,N_5489,N_5674);
nand U6466 (N_6466,N_5993,N_5272);
and U6467 (N_6467,N_5269,N_5975);
nand U6468 (N_6468,N_5467,N_5109);
nor U6469 (N_6469,N_5399,N_5084);
nor U6470 (N_6470,N_5948,N_5279);
and U6471 (N_6471,N_5845,N_5714);
or U6472 (N_6472,N_5486,N_5126);
nand U6473 (N_6473,N_5248,N_5931);
or U6474 (N_6474,N_5088,N_5639);
or U6475 (N_6475,N_5246,N_5270);
nand U6476 (N_6476,N_5054,N_5292);
or U6477 (N_6477,N_5717,N_5826);
xor U6478 (N_6478,N_5807,N_5158);
or U6479 (N_6479,N_5616,N_5635);
or U6480 (N_6480,N_5920,N_5933);
nor U6481 (N_6481,N_5385,N_5197);
or U6482 (N_6482,N_5934,N_5830);
or U6483 (N_6483,N_5569,N_5086);
or U6484 (N_6484,N_5041,N_5836);
nand U6485 (N_6485,N_5996,N_5628);
nor U6486 (N_6486,N_5691,N_5950);
and U6487 (N_6487,N_5690,N_5364);
and U6488 (N_6488,N_5776,N_5163);
or U6489 (N_6489,N_5198,N_5506);
nand U6490 (N_6490,N_5321,N_5519);
and U6491 (N_6491,N_5129,N_5145);
and U6492 (N_6492,N_5471,N_5566);
nor U6493 (N_6493,N_5760,N_5104);
nand U6494 (N_6494,N_5382,N_5300);
or U6495 (N_6495,N_5491,N_5885);
or U6496 (N_6496,N_5600,N_5431);
or U6497 (N_6497,N_5161,N_5026);
nand U6498 (N_6498,N_5838,N_5105);
and U6499 (N_6499,N_5132,N_5476);
nor U6500 (N_6500,N_5829,N_5400);
nand U6501 (N_6501,N_5531,N_5975);
and U6502 (N_6502,N_5147,N_5540);
or U6503 (N_6503,N_5208,N_5299);
or U6504 (N_6504,N_5952,N_5794);
nand U6505 (N_6505,N_5340,N_5757);
nand U6506 (N_6506,N_5323,N_5668);
nand U6507 (N_6507,N_5161,N_5795);
or U6508 (N_6508,N_5568,N_5814);
nor U6509 (N_6509,N_5339,N_5335);
nor U6510 (N_6510,N_5627,N_5743);
nand U6511 (N_6511,N_5144,N_5916);
and U6512 (N_6512,N_5644,N_5810);
and U6513 (N_6513,N_5094,N_5945);
nand U6514 (N_6514,N_5876,N_5487);
nor U6515 (N_6515,N_5853,N_5395);
nor U6516 (N_6516,N_5273,N_5333);
and U6517 (N_6517,N_5458,N_5600);
nor U6518 (N_6518,N_5541,N_5693);
and U6519 (N_6519,N_5689,N_5455);
nor U6520 (N_6520,N_5408,N_5615);
nor U6521 (N_6521,N_5081,N_5673);
nor U6522 (N_6522,N_5215,N_5685);
nor U6523 (N_6523,N_5295,N_5839);
nand U6524 (N_6524,N_5115,N_5774);
or U6525 (N_6525,N_5938,N_5672);
and U6526 (N_6526,N_5629,N_5827);
nand U6527 (N_6527,N_5489,N_5546);
and U6528 (N_6528,N_5190,N_5280);
and U6529 (N_6529,N_5056,N_5116);
or U6530 (N_6530,N_5763,N_5254);
nand U6531 (N_6531,N_5764,N_5334);
nor U6532 (N_6532,N_5707,N_5859);
and U6533 (N_6533,N_5971,N_5630);
nand U6534 (N_6534,N_5813,N_5016);
and U6535 (N_6535,N_5113,N_5226);
and U6536 (N_6536,N_5947,N_5689);
or U6537 (N_6537,N_5969,N_5292);
nand U6538 (N_6538,N_5637,N_5828);
or U6539 (N_6539,N_5989,N_5794);
and U6540 (N_6540,N_5443,N_5275);
nand U6541 (N_6541,N_5794,N_5265);
and U6542 (N_6542,N_5188,N_5823);
nand U6543 (N_6543,N_5313,N_5113);
nor U6544 (N_6544,N_5375,N_5417);
nand U6545 (N_6545,N_5873,N_5025);
and U6546 (N_6546,N_5536,N_5269);
nand U6547 (N_6547,N_5125,N_5846);
and U6548 (N_6548,N_5953,N_5354);
or U6549 (N_6549,N_5269,N_5735);
xor U6550 (N_6550,N_5175,N_5320);
and U6551 (N_6551,N_5914,N_5661);
nor U6552 (N_6552,N_5724,N_5305);
nor U6553 (N_6553,N_5703,N_5085);
nand U6554 (N_6554,N_5982,N_5577);
or U6555 (N_6555,N_5187,N_5158);
nand U6556 (N_6556,N_5453,N_5437);
and U6557 (N_6557,N_5670,N_5412);
nor U6558 (N_6558,N_5449,N_5394);
nand U6559 (N_6559,N_5019,N_5679);
or U6560 (N_6560,N_5276,N_5351);
nand U6561 (N_6561,N_5555,N_5083);
nor U6562 (N_6562,N_5462,N_5033);
or U6563 (N_6563,N_5820,N_5016);
nand U6564 (N_6564,N_5201,N_5129);
or U6565 (N_6565,N_5390,N_5097);
or U6566 (N_6566,N_5710,N_5572);
and U6567 (N_6567,N_5266,N_5241);
or U6568 (N_6568,N_5342,N_5343);
nor U6569 (N_6569,N_5612,N_5885);
nand U6570 (N_6570,N_5444,N_5052);
and U6571 (N_6571,N_5829,N_5489);
or U6572 (N_6572,N_5551,N_5508);
nor U6573 (N_6573,N_5570,N_5160);
or U6574 (N_6574,N_5652,N_5134);
nand U6575 (N_6575,N_5014,N_5129);
nand U6576 (N_6576,N_5146,N_5552);
nor U6577 (N_6577,N_5327,N_5666);
nor U6578 (N_6578,N_5714,N_5385);
or U6579 (N_6579,N_5449,N_5127);
nand U6580 (N_6580,N_5360,N_5114);
and U6581 (N_6581,N_5205,N_5720);
nand U6582 (N_6582,N_5973,N_5911);
or U6583 (N_6583,N_5748,N_5618);
nand U6584 (N_6584,N_5792,N_5235);
nor U6585 (N_6585,N_5509,N_5832);
or U6586 (N_6586,N_5400,N_5060);
and U6587 (N_6587,N_5047,N_5676);
or U6588 (N_6588,N_5747,N_5594);
nor U6589 (N_6589,N_5732,N_5094);
xnor U6590 (N_6590,N_5072,N_5566);
nand U6591 (N_6591,N_5138,N_5492);
or U6592 (N_6592,N_5258,N_5309);
xnor U6593 (N_6593,N_5294,N_5622);
or U6594 (N_6594,N_5467,N_5381);
or U6595 (N_6595,N_5769,N_5759);
nand U6596 (N_6596,N_5112,N_5075);
and U6597 (N_6597,N_5315,N_5502);
and U6598 (N_6598,N_5654,N_5644);
and U6599 (N_6599,N_5123,N_5063);
and U6600 (N_6600,N_5171,N_5000);
or U6601 (N_6601,N_5434,N_5647);
or U6602 (N_6602,N_5621,N_5262);
nand U6603 (N_6603,N_5288,N_5683);
or U6604 (N_6604,N_5425,N_5485);
nand U6605 (N_6605,N_5413,N_5463);
or U6606 (N_6606,N_5078,N_5999);
nand U6607 (N_6607,N_5261,N_5968);
nand U6608 (N_6608,N_5088,N_5531);
nand U6609 (N_6609,N_5608,N_5075);
nand U6610 (N_6610,N_5107,N_5553);
or U6611 (N_6611,N_5408,N_5719);
and U6612 (N_6612,N_5719,N_5246);
or U6613 (N_6613,N_5033,N_5611);
nand U6614 (N_6614,N_5522,N_5097);
nor U6615 (N_6615,N_5031,N_5592);
nand U6616 (N_6616,N_5096,N_5817);
or U6617 (N_6617,N_5962,N_5690);
nor U6618 (N_6618,N_5662,N_5121);
nand U6619 (N_6619,N_5407,N_5547);
nor U6620 (N_6620,N_5754,N_5689);
nor U6621 (N_6621,N_5746,N_5169);
nand U6622 (N_6622,N_5670,N_5304);
and U6623 (N_6623,N_5342,N_5935);
or U6624 (N_6624,N_5496,N_5293);
and U6625 (N_6625,N_5701,N_5060);
or U6626 (N_6626,N_5502,N_5115);
nand U6627 (N_6627,N_5304,N_5662);
and U6628 (N_6628,N_5343,N_5163);
or U6629 (N_6629,N_5264,N_5629);
and U6630 (N_6630,N_5829,N_5582);
or U6631 (N_6631,N_5651,N_5722);
nor U6632 (N_6632,N_5069,N_5793);
nor U6633 (N_6633,N_5137,N_5365);
nand U6634 (N_6634,N_5297,N_5391);
nand U6635 (N_6635,N_5259,N_5478);
nand U6636 (N_6636,N_5101,N_5106);
or U6637 (N_6637,N_5096,N_5223);
nor U6638 (N_6638,N_5128,N_5216);
and U6639 (N_6639,N_5822,N_5614);
and U6640 (N_6640,N_5163,N_5031);
nor U6641 (N_6641,N_5385,N_5471);
nand U6642 (N_6642,N_5714,N_5707);
nor U6643 (N_6643,N_5456,N_5162);
nand U6644 (N_6644,N_5190,N_5587);
and U6645 (N_6645,N_5155,N_5832);
nand U6646 (N_6646,N_5449,N_5408);
nand U6647 (N_6647,N_5734,N_5289);
or U6648 (N_6648,N_5166,N_5386);
and U6649 (N_6649,N_5361,N_5297);
nand U6650 (N_6650,N_5861,N_5300);
xnor U6651 (N_6651,N_5541,N_5706);
or U6652 (N_6652,N_5752,N_5059);
nand U6653 (N_6653,N_5583,N_5418);
and U6654 (N_6654,N_5928,N_5733);
or U6655 (N_6655,N_5704,N_5747);
nor U6656 (N_6656,N_5687,N_5691);
or U6657 (N_6657,N_5229,N_5204);
nor U6658 (N_6658,N_5261,N_5482);
nor U6659 (N_6659,N_5381,N_5754);
and U6660 (N_6660,N_5273,N_5456);
nand U6661 (N_6661,N_5531,N_5714);
and U6662 (N_6662,N_5377,N_5435);
and U6663 (N_6663,N_5643,N_5178);
and U6664 (N_6664,N_5988,N_5038);
or U6665 (N_6665,N_5195,N_5645);
nand U6666 (N_6666,N_5637,N_5821);
and U6667 (N_6667,N_5268,N_5714);
or U6668 (N_6668,N_5842,N_5816);
and U6669 (N_6669,N_5771,N_5850);
or U6670 (N_6670,N_5755,N_5340);
or U6671 (N_6671,N_5295,N_5541);
nor U6672 (N_6672,N_5009,N_5285);
and U6673 (N_6673,N_5201,N_5872);
and U6674 (N_6674,N_5868,N_5960);
or U6675 (N_6675,N_5789,N_5177);
and U6676 (N_6676,N_5711,N_5426);
nand U6677 (N_6677,N_5927,N_5570);
nor U6678 (N_6678,N_5278,N_5233);
nor U6679 (N_6679,N_5276,N_5108);
and U6680 (N_6680,N_5479,N_5125);
or U6681 (N_6681,N_5513,N_5787);
nand U6682 (N_6682,N_5508,N_5596);
and U6683 (N_6683,N_5829,N_5354);
and U6684 (N_6684,N_5090,N_5592);
and U6685 (N_6685,N_5911,N_5284);
or U6686 (N_6686,N_5320,N_5633);
or U6687 (N_6687,N_5510,N_5594);
nor U6688 (N_6688,N_5276,N_5803);
and U6689 (N_6689,N_5554,N_5673);
nand U6690 (N_6690,N_5623,N_5744);
xor U6691 (N_6691,N_5491,N_5839);
nor U6692 (N_6692,N_5231,N_5694);
and U6693 (N_6693,N_5861,N_5319);
or U6694 (N_6694,N_5682,N_5879);
or U6695 (N_6695,N_5109,N_5178);
and U6696 (N_6696,N_5795,N_5385);
nor U6697 (N_6697,N_5619,N_5187);
or U6698 (N_6698,N_5431,N_5450);
nand U6699 (N_6699,N_5835,N_5887);
or U6700 (N_6700,N_5042,N_5178);
and U6701 (N_6701,N_5571,N_5952);
nor U6702 (N_6702,N_5121,N_5726);
or U6703 (N_6703,N_5502,N_5901);
and U6704 (N_6704,N_5997,N_5681);
and U6705 (N_6705,N_5464,N_5847);
xor U6706 (N_6706,N_5018,N_5612);
and U6707 (N_6707,N_5048,N_5560);
nand U6708 (N_6708,N_5149,N_5316);
and U6709 (N_6709,N_5729,N_5497);
and U6710 (N_6710,N_5422,N_5894);
and U6711 (N_6711,N_5121,N_5252);
nand U6712 (N_6712,N_5643,N_5280);
xnor U6713 (N_6713,N_5204,N_5428);
nand U6714 (N_6714,N_5855,N_5094);
nand U6715 (N_6715,N_5225,N_5423);
nand U6716 (N_6716,N_5639,N_5780);
and U6717 (N_6717,N_5335,N_5215);
or U6718 (N_6718,N_5860,N_5922);
nand U6719 (N_6719,N_5924,N_5173);
or U6720 (N_6720,N_5257,N_5455);
and U6721 (N_6721,N_5108,N_5943);
nand U6722 (N_6722,N_5123,N_5430);
nand U6723 (N_6723,N_5432,N_5756);
and U6724 (N_6724,N_5424,N_5103);
or U6725 (N_6725,N_5270,N_5000);
nand U6726 (N_6726,N_5508,N_5355);
or U6727 (N_6727,N_5050,N_5034);
or U6728 (N_6728,N_5391,N_5186);
or U6729 (N_6729,N_5099,N_5971);
nor U6730 (N_6730,N_5989,N_5952);
nor U6731 (N_6731,N_5308,N_5788);
and U6732 (N_6732,N_5956,N_5422);
nand U6733 (N_6733,N_5002,N_5520);
nor U6734 (N_6734,N_5119,N_5138);
or U6735 (N_6735,N_5821,N_5204);
nand U6736 (N_6736,N_5267,N_5858);
nand U6737 (N_6737,N_5017,N_5302);
or U6738 (N_6738,N_5329,N_5994);
nand U6739 (N_6739,N_5099,N_5671);
nand U6740 (N_6740,N_5729,N_5686);
nand U6741 (N_6741,N_5044,N_5968);
nor U6742 (N_6742,N_5736,N_5443);
and U6743 (N_6743,N_5859,N_5600);
nand U6744 (N_6744,N_5926,N_5791);
or U6745 (N_6745,N_5632,N_5370);
and U6746 (N_6746,N_5729,N_5309);
and U6747 (N_6747,N_5311,N_5493);
or U6748 (N_6748,N_5737,N_5132);
nand U6749 (N_6749,N_5220,N_5846);
nand U6750 (N_6750,N_5281,N_5064);
nor U6751 (N_6751,N_5990,N_5190);
nand U6752 (N_6752,N_5768,N_5748);
nand U6753 (N_6753,N_5494,N_5382);
or U6754 (N_6754,N_5569,N_5323);
and U6755 (N_6755,N_5266,N_5308);
nor U6756 (N_6756,N_5329,N_5604);
nor U6757 (N_6757,N_5749,N_5645);
or U6758 (N_6758,N_5476,N_5792);
or U6759 (N_6759,N_5829,N_5887);
nand U6760 (N_6760,N_5111,N_5469);
or U6761 (N_6761,N_5206,N_5079);
nand U6762 (N_6762,N_5063,N_5795);
or U6763 (N_6763,N_5769,N_5332);
and U6764 (N_6764,N_5720,N_5160);
nor U6765 (N_6765,N_5608,N_5615);
or U6766 (N_6766,N_5058,N_5114);
nand U6767 (N_6767,N_5039,N_5459);
nor U6768 (N_6768,N_5262,N_5158);
or U6769 (N_6769,N_5567,N_5599);
nand U6770 (N_6770,N_5092,N_5495);
and U6771 (N_6771,N_5925,N_5940);
or U6772 (N_6772,N_5938,N_5000);
nand U6773 (N_6773,N_5515,N_5049);
nand U6774 (N_6774,N_5921,N_5243);
nor U6775 (N_6775,N_5257,N_5596);
or U6776 (N_6776,N_5653,N_5963);
or U6777 (N_6777,N_5493,N_5716);
and U6778 (N_6778,N_5304,N_5220);
nor U6779 (N_6779,N_5275,N_5922);
nor U6780 (N_6780,N_5263,N_5218);
nand U6781 (N_6781,N_5180,N_5549);
or U6782 (N_6782,N_5482,N_5283);
or U6783 (N_6783,N_5397,N_5276);
or U6784 (N_6784,N_5256,N_5041);
nand U6785 (N_6785,N_5618,N_5088);
or U6786 (N_6786,N_5064,N_5963);
or U6787 (N_6787,N_5093,N_5201);
or U6788 (N_6788,N_5650,N_5981);
nand U6789 (N_6789,N_5282,N_5034);
and U6790 (N_6790,N_5267,N_5208);
nor U6791 (N_6791,N_5504,N_5695);
nor U6792 (N_6792,N_5857,N_5062);
nor U6793 (N_6793,N_5086,N_5158);
nand U6794 (N_6794,N_5783,N_5198);
and U6795 (N_6795,N_5680,N_5207);
and U6796 (N_6796,N_5867,N_5187);
nor U6797 (N_6797,N_5304,N_5880);
nand U6798 (N_6798,N_5988,N_5631);
or U6799 (N_6799,N_5357,N_5597);
or U6800 (N_6800,N_5304,N_5190);
nor U6801 (N_6801,N_5293,N_5734);
nor U6802 (N_6802,N_5093,N_5685);
nor U6803 (N_6803,N_5107,N_5261);
or U6804 (N_6804,N_5422,N_5452);
or U6805 (N_6805,N_5366,N_5443);
nand U6806 (N_6806,N_5203,N_5910);
nand U6807 (N_6807,N_5893,N_5391);
and U6808 (N_6808,N_5701,N_5404);
and U6809 (N_6809,N_5258,N_5305);
or U6810 (N_6810,N_5992,N_5662);
or U6811 (N_6811,N_5809,N_5792);
nor U6812 (N_6812,N_5568,N_5931);
and U6813 (N_6813,N_5295,N_5502);
nor U6814 (N_6814,N_5200,N_5385);
nor U6815 (N_6815,N_5128,N_5219);
nor U6816 (N_6816,N_5951,N_5867);
or U6817 (N_6817,N_5507,N_5738);
nor U6818 (N_6818,N_5421,N_5636);
nand U6819 (N_6819,N_5546,N_5273);
nor U6820 (N_6820,N_5048,N_5400);
and U6821 (N_6821,N_5717,N_5323);
or U6822 (N_6822,N_5121,N_5709);
nor U6823 (N_6823,N_5073,N_5737);
nand U6824 (N_6824,N_5432,N_5152);
or U6825 (N_6825,N_5370,N_5663);
nand U6826 (N_6826,N_5870,N_5973);
nand U6827 (N_6827,N_5026,N_5839);
or U6828 (N_6828,N_5559,N_5582);
nor U6829 (N_6829,N_5460,N_5315);
nor U6830 (N_6830,N_5136,N_5200);
nand U6831 (N_6831,N_5256,N_5748);
nand U6832 (N_6832,N_5523,N_5796);
nand U6833 (N_6833,N_5464,N_5743);
nand U6834 (N_6834,N_5832,N_5676);
nor U6835 (N_6835,N_5504,N_5501);
and U6836 (N_6836,N_5865,N_5700);
nand U6837 (N_6837,N_5711,N_5295);
nand U6838 (N_6838,N_5297,N_5041);
nor U6839 (N_6839,N_5306,N_5727);
and U6840 (N_6840,N_5756,N_5884);
nand U6841 (N_6841,N_5612,N_5109);
and U6842 (N_6842,N_5440,N_5180);
and U6843 (N_6843,N_5033,N_5784);
or U6844 (N_6844,N_5921,N_5118);
and U6845 (N_6845,N_5730,N_5697);
nand U6846 (N_6846,N_5575,N_5519);
nand U6847 (N_6847,N_5090,N_5066);
nand U6848 (N_6848,N_5315,N_5687);
nand U6849 (N_6849,N_5729,N_5716);
and U6850 (N_6850,N_5592,N_5476);
or U6851 (N_6851,N_5438,N_5428);
nor U6852 (N_6852,N_5647,N_5118);
and U6853 (N_6853,N_5619,N_5963);
or U6854 (N_6854,N_5778,N_5262);
nand U6855 (N_6855,N_5511,N_5353);
nor U6856 (N_6856,N_5290,N_5997);
and U6857 (N_6857,N_5999,N_5884);
or U6858 (N_6858,N_5448,N_5244);
nand U6859 (N_6859,N_5921,N_5073);
or U6860 (N_6860,N_5124,N_5994);
nor U6861 (N_6861,N_5425,N_5440);
nor U6862 (N_6862,N_5225,N_5924);
and U6863 (N_6863,N_5115,N_5282);
nand U6864 (N_6864,N_5289,N_5667);
nand U6865 (N_6865,N_5886,N_5820);
and U6866 (N_6866,N_5877,N_5725);
or U6867 (N_6867,N_5401,N_5676);
and U6868 (N_6868,N_5033,N_5308);
nor U6869 (N_6869,N_5107,N_5220);
nor U6870 (N_6870,N_5935,N_5090);
and U6871 (N_6871,N_5510,N_5382);
and U6872 (N_6872,N_5118,N_5841);
nor U6873 (N_6873,N_5137,N_5261);
nand U6874 (N_6874,N_5454,N_5295);
nor U6875 (N_6875,N_5314,N_5593);
or U6876 (N_6876,N_5082,N_5504);
and U6877 (N_6877,N_5825,N_5427);
nor U6878 (N_6878,N_5671,N_5385);
nor U6879 (N_6879,N_5604,N_5574);
and U6880 (N_6880,N_5727,N_5205);
and U6881 (N_6881,N_5114,N_5202);
nand U6882 (N_6882,N_5326,N_5833);
nand U6883 (N_6883,N_5373,N_5388);
xor U6884 (N_6884,N_5269,N_5304);
and U6885 (N_6885,N_5059,N_5856);
and U6886 (N_6886,N_5383,N_5652);
nor U6887 (N_6887,N_5085,N_5544);
or U6888 (N_6888,N_5032,N_5398);
or U6889 (N_6889,N_5807,N_5831);
and U6890 (N_6890,N_5176,N_5671);
nand U6891 (N_6891,N_5140,N_5273);
or U6892 (N_6892,N_5205,N_5609);
nor U6893 (N_6893,N_5903,N_5677);
nand U6894 (N_6894,N_5259,N_5430);
nand U6895 (N_6895,N_5161,N_5617);
or U6896 (N_6896,N_5988,N_5206);
and U6897 (N_6897,N_5122,N_5845);
nand U6898 (N_6898,N_5661,N_5812);
nor U6899 (N_6899,N_5309,N_5015);
nand U6900 (N_6900,N_5032,N_5206);
or U6901 (N_6901,N_5740,N_5982);
nand U6902 (N_6902,N_5660,N_5122);
and U6903 (N_6903,N_5158,N_5726);
nor U6904 (N_6904,N_5662,N_5423);
nand U6905 (N_6905,N_5479,N_5733);
nor U6906 (N_6906,N_5895,N_5594);
nand U6907 (N_6907,N_5380,N_5611);
nor U6908 (N_6908,N_5386,N_5202);
nor U6909 (N_6909,N_5170,N_5390);
or U6910 (N_6910,N_5601,N_5671);
nor U6911 (N_6911,N_5304,N_5413);
nor U6912 (N_6912,N_5131,N_5362);
and U6913 (N_6913,N_5134,N_5227);
nand U6914 (N_6914,N_5565,N_5701);
and U6915 (N_6915,N_5044,N_5534);
nor U6916 (N_6916,N_5544,N_5102);
nand U6917 (N_6917,N_5395,N_5239);
nand U6918 (N_6918,N_5920,N_5805);
nor U6919 (N_6919,N_5782,N_5105);
and U6920 (N_6920,N_5003,N_5556);
or U6921 (N_6921,N_5601,N_5963);
nand U6922 (N_6922,N_5644,N_5420);
nand U6923 (N_6923,N_5347,N_5889);
nand U6924 (N_6924,N_5934,N_5039);
nand U6925 (N_6925,N_5786,N_5109);
nand U6926 (N_6926,N_5479,N_5552);
nand U6927 (N_6927,N_5525,N_5758);
and U6928 (N_6928,N_5504,N_5478);
nor U6929 (N_6929,N_5777,N_5846);
nand U6930 (N_6930,N_5819,N_5373);
or U6931 (N_6931,N_5599,N_5716);
or U6932 (N_6932,N_5869,N_5838);
and U6933 (N_6933,N_5433,N_5024);
nand U6934 (N_6934,N_5590,N_5606);
nand U6935 (N_6935,N_5705,N_5224);
nand U6936 (N_6936,N_5580,N_5230);
nand U6937 (N_6937,N_5661,N_5774);
or U6938 (N_6938,N_5185,N_5532);
and U6939 (N_6939,N_5733,N_5578);
xnor U6940 (N_6940,N_5776,N_5810);
nand U6941 (N_6941,N_5795,N_5839);
nor U6942 (N_6942,N_5825,N_5287);
or U6943 (N_6943,N_5814,N_5509);
or U6944 (N_6944,N_5393,N_5185);
nor U6945 (N_6945,N_5977,N_5209);
nor U6946 (N_6946,N_5614,N_5552);
or U6947 (N_6947,N_5499,N_5715);
and U6948 (N_6948,N_5363,N_5295);
or U6949 (N_6949,N_5847,N_5455);
nand U6950 (N_6950,N_5181,N_5867);
and U6951 (N_6951,N_5074,N_5653);
and U6952 (N_6952,N_5252,N_5696);
or U6953 (N_6953,N_5623,N_5673);
or U6954 (N_6954,N_5110,N_5267);
and U6955 (N_6955,N_5534,N_5225);
nand U6956 (N_6956,N_5768,N_5339);
nand U6957 (N_6957,N_5028,N_5282);
and U6958 (N_6958,N_5283,N_5867);
and U6959 (N_6959,N_5743,N_5548);
and U6960 (N_6960,N_5492,N_5099);
and U6961 (N_6961,N_5392,N_5901);
nor U6962 (N_6962,N_5742,N_5111);
nor U6963 (N_6963,N_5402,N_5972);
and U6964 (N_6964,N_5240,N_5532);
or U6965 (N_6965,N_5071,N_5000);
or U6966 (N_6966,N_5803,N_5580);
and U6967 (N_6967,N_5817,N_5217);
or U6968 (N_6968,N_5250,N_5671);
and U6969 (N_6969,N_5109,N_5791);
nor U6970 (N_6970,N_5684,N_5268);
nor U6971 (N_6971,N_5679,N_5258);
and U6972 (N_6972,N_5313,N_5334);
nand U6973 (N_6973,N_5299,N_5436);
nand U6974 (N_6974,N_5236,N_5133);
and U6975 (N_6975,N_5469,N_5866);
and U6976 (N_6976,N_5318,N_5597);
nor U6977 (N_6977,N_5348,N_5212);
nor U6978 (N_6978,N_5025,N_5381);
nand U6979 (N_6979,N_5500,N_5085);
nand U6980 (N_6980,N_5538,N_5993);
nand U6981 (N_6981,N_5882,N_5165);
and U6982 (N_6982,N_5878,N_5871);
nor U6983 (N_6983,N_5433,N_5337);
nand U6984 (N_6984,N_5900,N_5966);
or U6985 (N_6985,N_5140,N_5233);
or U6986 (N_6986,N_5076,N_5807);
nor U6987 (N_6987,N_5232,N_5358);
and U6988 (N_6988,N_5921,N_5710);
nand U6989 (N_6989,N_5088,N_5924);
nand U6990 (N_6990,N_5780,N_5723);
nor U6991 (N_6991,N_5898,N_5095);
nor U6992 (N_6992,N_5963,N_5249);
or U6993 (N_6993,N_5586,N_5335);
nand U6994 (N_6994,N_5239,N_5358);
and U6995 (N_6995,N_5718,N_5195);
nor U6996 (N_6996,N_5563,N_5597);
nor U6997 (N_6997,N_5844,N_5197);
or U6998 (N_6998,N_5887,N_5342);
or U6999 (N_6999,N_5327,N_5757);
and U7000 (N_7000,N_6246,N_6806);
and U7001 (N_7001,N_6749,N_6924);
nand U7002 (N_7002,N_6697,N_6771);
nand U7003 (N_7003,N_6177,N_6028);
and U7004 (N_7004,N_6886,N_6862);
nand U7005 (N_7005,N_6432,N_6292);
nand U7006 (N_7006,N_6724,N_6005);
nand U7007 (N_7007,N_6152,N_6585);
and U7008 (N_7008,N_6860,N_6078);
nor U7009 (N_7009,N_6242,N_6163);
and U7010 (N_7010,N_6944,N_6117);
xor U7011 (N_7011,N_6759,N_6682);
and U7012 (N_7012,N_6065,N_6095);
or U7013 (N_7013,N_6788,N_6981);
and U7014 (N_7014,N_6408,N_6165);
nand U7015 (N_7015,N_6300,N_6146);
nor U7016 (N_7016,N_6138,N_6441);
nand U7017 (N_7017,N_6828,N_6977);
nand U7018 (N_7018,N_6639,N_6086);
and U7019 (N_7019,N_6983,N_6495);
nor U7020 (N_7020,N_6107,N_6079);
nor U7021 (N_7021,N_6700,N_6919);
nand U7022 (N_7022,N_6746,N_6371);
nand U7023 (N_7023,N_6468,N_6511);
and U7024 (N_7024,N_6528,N_6387);
or U7025 (N_7025,N_6849,N_6710);
or U7026 (N_7026,N_6580,N_6265);
nand U7027 (N_7027,N_6046,N_6324);
or U7028 (N_7028,N_6124,N_6933);
nand U7029 (N_7029,N_6023,N_6821);
nand U7030 (N_7030,N_6449,N_6601);
nor U7031 (N_7031,N_6407,N_6956);
nor U7032 (N_7032,N_6647,N_6189);
or U7033 (N_7033,N_6323,N_6606);
nor U7034 (N_7034,N_6636,N_6998);
nand U7035 (N_7035,N_6872,N_6804);
and U7036 (N_7036,N_6794,N_6744);
and U7037 (N_7037,N_6178,N_6176);
and U7038 (N_7038,N_6516,N_6793);
nand U7039 (N_7039,N_6971,N_6876);
nand U7040 (N_7040,N_6121,N_6572);
or U7041 (N_7041,N_6277,N_6627);
or U7042 (N_7042,N_6061,N_6421);
nand U7043 (N_7043,N_6913,N_6846);
nor U7044 (N_7044,N_6181,N_6032);
or U7045 (N_7045,N_6471,N_6366);
or U7046 (N_7046,N_6745,N_6708);
nand U7047 (N_7047,N_6772,N_6409);
and U7048 (N_7048,N_6493,N_6494);
nor U7049 (N_7049,N_6676,N_6762);
or U7050 (N_7050,N_6004,N_6497);
and U7051 (N_7051,N_6444,N_6501);
nor U7052 (N_7052,N_6080,N_6241);
nor U7053 (N_7053,N_6670,N_6765);
nand U7054 (N_7054,N_6056,N_6083);
nand U7055 (N_7055,N_6690,N_6395);
nand U7056 (N_7056,N_6452,N_6049);
or U7057 (N_7057,N_6739,N_6760);
nand U7058 (N_7058,N_6200,N_6466);
nand U7059 (N_7059,N_6375,N_6558);
or U7060 (N_7060,N_6365,N_6225);
nand U7061 (N_7061,N_6029,N_6467);
and U7062 (N_7062,N_6942,N_6964);
nor U7063 (N_7063,N_6819,N_6287);
and U7064 (N_7064,N_6425,N_6472);
nor U7065 (N_7065,N_6605,N_6037);
or U7066 (N_7066,N_6156,N_6115);
or U7067 (N_7067,N_6011,N_6024);
nand U7068 (N_7068,N_6948,N_6677);
or U7069 (N_7069,N_6057,N_6884);
nand U7070 (N_7070,N_6282,N_6003);
and U7071 (N_7071,N_6829,N_6027);
nand U7072 (N_7072,N_6680,N_6747);
or U7073 (N_7073,N_6344,N_6826);
and U7074 (N_7074,N_6638,N_6487);
or U7075 (N_7075,N_6654,N_6322);
nor U7076 (N_7076,N_6135,N_6986);
and U7077 (N_7077,N_6930,N_6567);
nand U7078 (N_7078,N_6073,N_6215);
nand U7079 (N_7079,N_6656,N_6554);
and U7080 (N_7080,N_6419,N_6067);
or U7081 (N_7081,N_6123,N_6085);
or U7082 (N_7082,N_6614,N_6321);
nor U7083 (N_7083,N_6183,N_6608);
nor U7084 (N_7084,N_6485,N_6034);
or U7085 (N_7085,N_6524,N_6458);
nand U7086 (N_7086,N_6349,N_6858);
or U7087 (N_7087,N_6380,N_6573);
nand U7088 (N_7088,N_6811,N_6888);
nand U7089 (N_7089,N_6790,N_6206);
and U7090 (N_7090,N_6920,N_6100);
nand U7091 (N_7091,N_6403,N_6835);
and U7092 (N_7092,N_6119,N_6370);
and U7093 (N_7093,N_6478,N_6768);
and U7094 (N_7094,N_6650,N_6574);
or U7095 (N_7095,N_6069,N_6332);
or U7096 (N_7096,N_6757,N_6263);
nand U7097 (N_7097,N_6801,N_6378);
or U7098 (N_7098,N_6512,N_6127);
or U7099 (N_7099,N_6576,N_6149);
or U7100 (N_7100,N_6847,N_6406);
nor U7101 (N_7101,N_6714,N_6267);
or U7102 (N_7102,N_6338,N_6557);
nand U7103 (N_7103,N_6996,N_6162);
and U7104 (N_7104,N_6489,N_6609);
or U7105 (N_7105,N_6549,N_6326);
nor U7106 (N_7106,N_6743,N_6304);
nand U7107 (N_7107,N_6173,N_6994);
and U7108 (N_7108,N_6210,N_6020);
or U7109 (N_7109,N_6018,N_6686);
nand U7110 (N_7110,N_6988,N_6040);
xnor U7111 (N_7111,N_6174,N_6187);
and U7112 (N_7112,N_6298,N_6632);
nand U7113 (N_7113,N_6274,N_6667);
or U7114 (N_7114,N_6587,N_6684);
nor U7115 (N_7115,N_6613,N_6195);
or U7116 (N_7116,N_6052,N_6653);
nand U7117 (N_7117,N_6240,N_6327);
and U7118 (N_7118,N_6637,N_6373);
nand U7119 (N_7119,N_6498,N_6773);
nor U7120 (N_7120,N_6623,N_6622);
or U7121 (N_7121,N_6553,N_6405);
and U7122 (N_7122,N_6669,N_6892);
xor U7123 (N_7123,N_6541,N_6068);
nor U7124 (N_7124,N_6685,N_6222);
nand U7125 (N_7125,N_6514,N_6674);
nor U7126 (N_7126,N_6130,N_6281);
or U7127 (N_7127,N_6384,N_6188);
xor U7128 (N_7128,N_6354,N_6460);
and U7129 (N_7129,N_6051,N_6232);
or U7130 (N_7130,N_6589,N_6869);
or U7131 (N_7131,N_6715,N_6989);
nand U7132 (N_7132,N_6129,N_6792);
nand U7133 (N_7133,N_6500,N_6503);
and U7134 (N_7134,N_6529,N_6887);
nand U7135 (N_7135,N_6251,N_6523);
or U7136 (N_7136,N_6525,N_6019);
nand U7137 (N_7137,N_6642,N_6730);
nand U7138 (N_7138,N_6249,N_6381);
or U7139 (N_7139,N_6191,N_6278);
nand U7140 (N_7140,N_6470,N_6770);
or U7141 (N_7141,N_6317,N_6615);
nor U7142 (N_7142,N_6959,N_6911);
or U7143 (N_7143,N_6900,N_6170);
or U7144 (N_7144,N_6270,N_6430);
xor U7145 (N_7145,N_6015,N_6054);
and U7146 (N_7146,N_6041,N_6357);
nor U7147 (N_7147,N_6641,N_6390);
nor U7148 (N_7148,N_6290,N_6343);
nand U7149 (N_7149,N_6481,N_6861);
nor U7150 (N_7150,N_6142,N_6379);
and U7151 (N_7151,N_6388,N_6845);
nor U7152 (N_7152,N_6256,N_6031);
or U7153 (N_7153,N_6852,N_6795);
and U7154 (N_7154,N_6644,N_6219);
nor U7155 (N_7155,N_6877,N_6518);
nand U7156 (N_7156,N_6935,N_6209);
and U7157 (N_7157,N_6299,N_6448);
and U7158 (N_7158,N_6698,N_6443);
nor U7159 (N_7159,N_6348,N_6313);
and U7160 (N_7160,N_6979,N_6383);
or U7161 (N_7161,N_6681,N_6372);
nor U7162 (N_7162,N_6036,N_6310);
nand U7163 (N_7163,N_6258,N_6602);
nor U7164 (N_7164,N_6717,N_6668);
nand U7165 (N_7165,N_6253,N_6030);
or U7166 (N_7166,N_6076,N_6537);
nand U7167 (N_7167,N_6937,N_6734);
or U7168 (N_7168,N_6562,N_6917);
nor U7169 (N_7169,N_6486,N_6202);
nand U7170 (N_7170,N_6014,N_6465);
nand U7171 (N_7171,N_6141,N_6314);
nand U7172 (N_7172,N_6890,N_6775);
nor U7173 (N_7173,N_6891,N_6865);
nand U7174 (N_7174,N_6045,N_6837);
nand U7175 (N_7175,N_6473,N_6145);
and U7176 (N_7176,N_6047,N_6547);
nand U7177 (N_7177,N_6205,N_6836);
nor U7178 (N_7178,N_6907,N_6534);
nor U7179 (N_7179,N_6412,N_6955);
nand U7180 (N_7180,N_6429,N_6755);
or U7181 (N_7181,N_6551,N_6185);
nor U7182 (N_7182,N_6564,N_6342);
nor U7183 (N_7183,N_6612,N_6603);
xnor U7184 (N_7184,N_6803,N_6105);
or U7185 (N_7185,N_6198,N_6597);
nor U7186 (N_7186,N_6675,N_6442);
and U7187 (N_7187,N_6131,N_6995);
nor U7188 (N_7188,N_6233,N_6719);
nand U7189 (N_7189,N_6368,N_6306);
xnor U7190 (N_7190,N_6264,N_6160);
or U7191 (N_7191,N_6382,N_6483);
nor U7192 (N_7192,N_6910,N_6113);
or U7193 (N_7193,N_6101,N_6280);
nand U7194 (N_7194,N_6451,N_6112);
nand U7195 (N_7195,N_6231,N_6437);
nor U7196 (N_7196,N_6401,N_6856);
xor U7197 (N_7197,N_6477,N_6611);
or U7198 (N_7198,N_6575,N_6226);
or U7199 (N_7199,N_6659,N_6974);
or U7200 (N_7200,N_6946,N_6905);
and U7201 (N_7201,N_6022,N_6157);
or U7202 (N_7202,N_6752,N_6969);
xor U7203 (N_7203,N_6137,N_6626);
or U7204 (N_7204,N_6586,N_6921);
and U7205 (N_7205,N_6651,N_6218);
and U7206 (N_7206,N_6158,N_6758);
nand U7207 (N_7207,N_6832,N_6873);
nand U7208 (N_7208,N_6293,N_6619);
and U7209 (N_7209,N_6712,N_6392);
and U7210 (N_7210,N_6404,N_6629);
nand U7211 (N_7211,N_6064,N_6201);
and U7212 (N_7212,N_6440,N_6081);
and U7213 (N_7213,N_6997,N_6958);
nand U7214 (N_7214,N_6925,N_6699);
nand U7215 (N_7215,N_6657,N_6221);
or U7216 (N_7216,N_6340,N_6513);
and U7217 (N_7217,N_6017,N_6800);
nand U7218 (N_7218,N_6134,N_6088);
nand U7219 (N_7219,N_6013,N_6914);
or U7220 (N_7220,N_6339,N_6171);
nor U7221 (N_7221,N_6302,N_6376);
nor U7222 (N_7222,N_6199,N_6966);
nand U7223 (N_7223,N_6179,N_6211);
nor U7224 (N_7224,N_6940,N_6866);
or U7225 (N_7225,N_6649,N_6560);
or U7226 (N_7226,N_6662,N_6255);
nand U7227 (N_7227,N_6389,N_6168);
nor U7228 (N_7228,N_6731,N_6797);
nor U7229 (N_7229,N_6791,N_6972);
nor U7230 (N_7230,N_6732,N_6414);
nor U7231 (N_7231,N_6616,N_6630);
nor U7232 (N_7232,N_6620,N_6507);
nor U7233 (N_7233,N_6993,N_6128);
nand U7234 (N_7234,N_6025,N_6672);
nor U7235 (N_7235,N_6026,N_6090);
nand U7236 (N_7236,N_6320,N_6454);
and U7237 (N_7237,N_6318,N_6645);
and U7238 (N_7238,N_6418,N_6631);
nand U7239 (N_7239,N_6583,N_6457);
and U7240 (N_7240,N_6927,N_6953);
and U7241 (N_7241,N_6154,N_6531);
or U7242 (N_7242,N_6542,N_6702);
and U7243 (N_7243,N_6087,N_6802);
or U7244 (N_7244,N_6506,N_6853);
and U7245 (N_7245,N_6782,N_6262);
and U7246 (N_7246,N_6704,N_6661);
nor U7247 (N_7247,N_6439,N_6915);
nor U7248 (N_7248,N_6742,N_6143);
nand U7249 (N_7249,N_6857,N_6035);
nor U7250 (N_7250,N_6545,N_6723);
or U7251 (N_7251,N_6565,N_6254);
nor U7252 (N_7252,N_6526,N_6386);
nand U7253 (N_7253,N_6038,N_6491);
and U7254 (N_7254,N_6823,N_6735);
nand U7255 (N_7255,N_6607,N_6947);
nand U7256 (N_7256,N_6329,N_6398);
nand U7257 (N_7257,N_6520,N_6960);
and U7258 (N_7258,N_6726,N_6266);
nand U7259 (N_7259,N_6519,N_6741);
and U7260 (N_7260,N_6751,N_6346);
or U7261 (N_7261,N_6590,N_6691);
or U7262 (N_7262,N_6875,N_6103);
or U7263 (N_7263,N_6367,N_6785);
nand U7264 (N_7264,N_6713,N_6840);
nand U7265 (N_7265,N_6237,N_6099);
or U7266 (N_7266,N_6968,N_6863);
nand U7267 (N_7267,N_6132,N_6902);
nor U7268 (N_7268,N_6377,N_6396);
or U7269 (N_7269,N_6786,N_6546);
nand U7270 (N_7270,N_6161,N_6217);
nor U7271 (N_7271,N_6753,N_6683);
nand U7272 (N_7272,N_6918,N_6515);
nor U7273 (N_7273,N_6830,N_6147);
and U7274 (N_7274,N_6182,N_6268);
and U7275 (N_7275,N_6008,N_6663);
or U7276 (N_7276,N_6416,N_6220);
and U7277 (N_7277,N_6725,N_6360);
nor U7278 (N_7278,N_6492,N_6315);
or U7279 (N_7279,N_6350,N_6422);
nand U7280 (N_7280,N_6854,N_6707);
nor U7281 (N_7281,N_6949,N_6294);
nor U7282 (N_7282,N_6796,N_6692);
nor U7283 (N_7283,N_6261,N_6729);
nand U7284 (N_7284,N_6279,N_6736);
or U7285 (N_7285,N_6916,N_6144);
nand U7286 (N_7286,N_6756,N_6043);
nor U7287 (N_7287,N_6063,N_6001);
nor U7288 (N_7288,N_6484,N_6559);
nand U7289 (N_7289,N_6943,N_6635);
nor U7290 (N_7290,N_6167,N_6336);
nor U7291 (N_7291,N_6415,N_6588);
and U7292 (N_7292,N_6643,N_6530);
or U7293 (N_7293,N_6312,N_6664);
or U7294 (N_7294,N_6247,N_6070);
or U7295 (N_7295,N_6355,N_6807);
nor U7296 (N_7296,N_6062,N_6563);
nand U7297 (N_7297,N_6550,N_6197);
nand U7298 (N_7298,N_6665,N_6508);
or U7299 (N_7299,N_6783,N_6555);
or U7300 (N_7300,N_6248,N_6307);
nor U7301 (N_7301,N_6438,N_6058);
and U7302 (N_7302,N_6628,N_6999);
nor U7303 (N_7303,N_6108,N_6688);
and U7304 (N_7304,N_6453,N_6000);
or U7305 (N_7305,N_6213,N_6301);
nor U7306 (N_7306,N_6055,N_6505);
or U7307 (N_7307,N_6309,N_6475);
or U7308 (N_7308,N_6878,N_6275);
and U7309 (N_7309,N_6288,N_6991);
and U7310 (N_7310,N_6831,N_6776);
nor U7311 (N_7311,N_6599,N_6071);
nand U7312 (N_7312,N_6976,N_6402);
nand U7313 (N_7313,N_6330,N_6824);
nor U7314 (N_7314,N_6571,N_6196);
nor U7315 (N_7315,N_6718,N_6166);
nor U7316 (N_7316,N_6450,N_6413);
and U7317 (N_7317,N_6952,N_6798);
or U7318 (N_7318,N_6985,N_6906);
and U7319 (N_7319,N_6111,N_6394);
nand U7320 (N_7320,N_6813,N_6042);
nor U7321 (N_7321,N_6136,N_6295);
or U7322 (N_7322,N_6420,N_6252);
and U7323 (N_7323,N_6652,N_6228);
nor U7324 (N_7324,N_6369,N_6738);
nor U7325 (N_7325,N_6552,N_6094);
or U7326 (N_7326,N_6767,N_6456);
and U7327 (N_7327,N_6646,N_6016);
or U7328 (N_7328,N_6291,N_6098);
or U7329 (N_7329,N_6347,N_6694);
or U7330 (N_7330,N_6397,N_6110);
or U7331 (N_7331,N_6864,N_6333);
nand U7332 (N_7332,N_6434,N_6337);
nor U7333 (N_7333,N_6316,N_6479);
nand U7334 (N_7334,N_6893,N_6364);
or U7335 (N_7335,N_6728,N_6216);
nand U7336 (N_7336,N_6581,N_6568);
nor U7337 (N_7337,N_6841,N_6334);
or U7338 (N_7338,N_6400,N_6072);
or U7339 (N_7339,N_6356,N_6950);
nor U7340 (N_7340,N_6737,N_6104);
or U7341 (N_7341,N_6543,N_6303);
or U7342 (N_7342,N_6345,N_6109);
or U7343 (N_7343,N_6781,N_6780);
or U7344 (N_7344,N_6621,N_6848);
nor U7345 (N_7345,N_6490,N_6880);
and U7346 (N_7346,N_6509,N_6850);
nor U7347 (N_7347,N_6992,N_6640);
nand U7348 (N_7348,N_6923,N_6778);
and U7349 (N_7349,N_6810,N_6053);
nand U7350 (N_7350,N_6812,N_6496);
or U7351 (N_7351,N_6727,N_6987);
nor U7352 (N_7352,N_6305,N_6689);
and U7353 (N_7353,N_6150,N_6687);
or U7354 (N_7354,N_6982,N_6633);
nor U7355 (N_7355,N_6363,N_6570);
nand U7356 (N_7356,N_6871,N_6764);
xnor U7357 (N_7357,N_6883,N_6624);
nand U7358 (N_7358,N_6060,N_6148);
nand U7359 (N_7359,N_6223,N_6527);
xnor U7360 (N_7360,N_6351,N_6229);
and U7361 (N_7361,N_6259,N_6705);
and U7362 (N_7362,N_6427,N_6120);
and U7363 (N_7363,N_6816,N_6899);
nor U7364 (N_7364,N_6750,N_6139);
nand U7365 (N_7365,N_6721,N_6469);
nor U7366 (N_7366,N_6391,N_6777);
nor U7367 (N_7367,N_6331,N_6385);
nor U7368 (N_7368,N_6954,N_6593);
xnor U7369 (N_7369,N_6243,N_6561);
nor U7370 (N_7370,N_6010,N_6289);
nand U7371 (N_7371,N_6701,N_6720);
nand U7372 (N_7372,N_6932,N_6180);
nor U7373 (N_7373,N_6926,N_6678);
and U7374 (N_7374,N_6352,N_6897);
nor U7375 (N_7375,N_6814,N_6660);
and U7376 (N_7376,N_6273,N_6285);
nor U7377 (N_7377,N_6361,N_6474);
nor U7378 (N_7378,N_6227,N_6423);
xor U7379 (N_7379,N_6695,N_6193);
nor U7380 (N_7380,N_6990,N_6059);
nor U7381 (N_7381,N_6445,N_6286);
nor U7382 (N_7382,N_6673,N_6787);
and U7383 (N_7383,N_6870,N_6617);
nor U7384 (N_7384,N_6102,N_6815);
and U7385 (N_7385,N_6904,N_6048);
nor U7386 (N_7386,N_6164,N_6433);
nor U7387 (N_7387,N_6125,N_6033);
and U7388 (N_7388,N_6928,N_6766);
nand U7389 (N_7389,N_6186,N_6584);
or U7390 (N_7390,N_6319,N_6885);
nand U7391 (N_7391,N_6140,N_6212);
or U7392 (N_7392,N_6532,N_6431);
or U7393 (N_7393,N_6984,N_6868);
or U7394 (N_7394,N_6244,N_6961);
nand U7395 (N_7395,N_6833,N_6203);
and U7396 (N_7396,N_6963,N_6522);
nand U7397 (N_7397,N_6446,N_6938);
and U7398 (N_7398,N_6598,N_6703);
nor U7399 (N_7399,N_6250,N_6945);
or U7400 (N_7400,N_6133,N_6359);
nor U7401 (N_7401,N_6908,N_6634);
or U7402 (N_7402,N_6151,N_6084);
nor U7403 (N_7403,N_6842,N_6709);
and U7404 (N_7404,N_6825,N_6779);
nand U7405 (N_7405,N_6276,N_6459);
nand U7406 (N_7406,N_6410,N_6239);
nor U7407 (N_7407,N_6012,N_6044);
nor U7408 (N_7408,N_6896,N_6194);
and U7409 (N_7409,N_6435,N_6610);
or U7410 (N_7410,N_6851,N_6510);
nand U7411 (N_7411,N_6358,N_6648);
or U7412 (N_7412,N_6679,N_6957);
nand U7413 (N_7413,N_6962,N_6879);
or U7414 (N_7414,N_6499,N_6399);
or U7415 (N_7415,N_6393,N_6895);
and U7416 (N_7416,N_6096,N_6973);
and U7417 (N_7417,N_6106,N_6855);
or U7418 (N_7418,N_6362,N_6476);
and U7419 (N_7419,N_6426,N_6595);
nor U7420 (N_7420,N_6066,N_6582);
or U7421 (N_7421,N_6172,N_6539);
nand U7422 (N_7422,N_6461,N_6901);
nand U7423 (N_7423,N_6579,N_6578);
nand U7424 (N_7424,N_6834,N_6092);
or U7425 (N_7425,N_6600,N_6074);
nor U7426 (N_7426,N_6941,N_6748);
or U7427 (N_7427,N_6556,N_6592);
nand U7428 (N_7428,N_6844,N_6462);
nor U7429 (N_7429,N_6021,N_6482);
and U7430 (N_7430,N_6536,N_6722);
nor U7431 (N_7431,N_6693,N_6827);
nand U7432 (N_7432,N_6859,N_6909);
nand U7433 (N_7433,N_6591,N_6411);
nor U7434 (N_7434,N_6271,N_6696);
nor U7435 (N_7435,N_6488,N_6839);
nand U7436 (N_7436,N_6082,N_6774);
nor U7437 (N_7437,N_6658,N_6236);
nand U7438 (N_7438,N_6504,N_6789);
nand U7439 (N_7439,N_6296,N_6325);
and U7440 (N_7440,N_6122,N_6596);
and U7441 (N_7441,N_6889,N_6769);
or U7442 (N_7442,N_6533,N_6208);
nand U7443 (N_7443,N_6838,N_6308);
nand U7444 (N_7444,N_6655,N_6666);
and U7445 (N_7445,N_6039,N_6169);
and U7446 (N_7446,N_6799,N_6230);
and U7447 (N_7447,N_6341,N_6951);
nand U7448 (N_7448,N_6257,N_6867);
and U7449 (N_7449,N_6007,N_6009);
nand U7450 (N_7450,N_6238,N_6126);
or U7451 (N_7451,N_6002,N_6894);
nand U7452 (N_7452,N_6538,N_6184);
and U7453 (N_7453,N_6464,N_6335);
or U7454 (N_7454,N_6116,N_6207);
nand U7455 (N_7455,N_6297,N_6091);
nand U7456 (N_7456,N_6214,N_6155);
nand U7457 (N_7457,N_6089,N_6159);
and U7458 (N_7458,N_6874,N_6763);
and U7459 (N_7459,N_6912,N_6328);
nand U7460 (N_7460,N_6929,N_6980);
nor U7461 (N_7461,N_6447,N_6077);
and U7462 (N_7462,N_6153,N_6175);
and U7463 (N_7463,N_6808,N_6843);
nand U7464 (N_7464,N_6939,N_6480);
or U7465 (N_7465,N_6970,N_6548);
xnor U7466 (N_7466,N_6284,N_6006);
and U7467 (N_7467,N_6711,N_6967);
and U7468 (N_7468,N_6118,N_6269);
nand U7469 (N_7469,N_6192,N_6424);
nor U7470 (N_7470,N_6934,N_6881);
or U7471 (N_7471,N_6544,N_6234);
nor U7472 (N_7472,N_6965,N_6204);
or U7473 (N_7473,N_6093,N_6417);
nor U7474 (N_7474,N_6903,N_6820);
and U7475 (N_7475,N_6882,N_6050);
and U7476 (N_7476,N_6260,N_6805);
and U7477 (N_7477,N_6818,N_6978);
or U7478 (N_7478,N_6733,N_6936);
nand U7479 (N_7479,N_6114,N_6569);
or U7480 (N_7480,N_6740,N_6190);
nand U7481 (N_7481,N_6097,N_6235);
nor U7482 (N_7482,N_6625,N_6283);
or U7483 (N_7483,N_6502,N_6566);
nor U7484 (N_7484,N_6374,N_6784);
or U7485 (N_7485,N_6817,N_6809);
nor U7486 (N_7486,N_6521,N_6540);
or U7487 (N_7487,N_6931,N_6594);
or U7488 (N_7488,N_6671,N_6075);
and U7489 (N_7489,N_6463,N_6975);
or U7490 (N_7490,N_6436,N_6455);
nor U7491 (N_7491,N_6311,N_6922);
and U7492 (N_7492,N_6272,N_6577);
nor U7493 (N_7493,N_6224,N_6706);
and U7494 (N_7494,N_6716,N_6353);
and U7495 (N_7495,N_6535,N_6428);
or U7496 (N_7496,N_6517,N_6245);
or U7497 (N_7497,N_6754,N_6822);
and U7498 (N_7498,N_6604,N_6618);
nand U7499 (N_7499,N_6898,N_6761);
and U7500 (N_7500,N_6659,N_6774);
nand U7501 (N_7501,N_6025,N_6106);
or U7502 (N_7502,N_6002,N_6086);
or U7503 (N_7503,N_6734,N_6620);
nand U7504 (N_7504,N_6580,N_6296);
or U7505 (N_7505,N_6468,N_6711);
nand U7506 (N_7506,N_6390,N_6955);
nor U7507 (N_7507,N_6918,N_6093);
nand U7508 (N_7508,N_6993,N_6584);
xor U7509 (N_7509,N_6261,N_6258);
and U7510 (N_7510,N_6876,N_6690);
nand U7511 (N_7511,N_6570,N_6327);
or U7512 (N_7512,N_6879,N_6678);
and U7513 (N_7513,N_6367,N_6221);
nor U7514 (N_7514,N_6660,N_6626);
and U7515 (N_7515,N_6345,N_6567);
nand U7516 (N_7516,N_6031,N_6747);
or U7517 (N_7517,N_6433,N_6898);
and U7518 (N_7518,N_6885,N_6485);
or U7519 (N_7519,N_6677,N_6958);
nand U7520 (N_7520,N_6979,N_6437);
and U7521 (N_7521,N_6233,N_6547);
nor U7522 (N_7522,N_6401,N_6887);
nand U7523 (N_7523,N_6271,N_6283);
and U7524 (N_7524,N_6247,N_6924);
nor U7525 (N_7525,N_6621,N_6873);
and U7526 (N_7526,N_6268,N_6541);
or U7527 (N_7527,N_6709,N_6240);
nand U7528 (N_7528,N_6526,N_6337);
nor U7529 (N_7529,N_6199,N_6159);
and U7530 (N_7530,N_6957,N_6978);
nor U7531 (N_7531,N_6872,N_6716);
and U7532 (N_7532,N_6741,N_6353);
nand U7533 (N_7533,N_6369,N_6849);
and U7534 (N_7534,N_6072,N_6839);
or U7535 (N_7535,N_6471,N_6653);
and U7536 (N_7536,N_6654,N_6407);
nand U7537 (N_7537,N_6271,N_6961);
nand U7538 (N_7538,N_6293,N_6530);
nand U7539 (N_7539,N_6769,N_6458);
nand U7540 (N_7540,N_6092,N_6021);
nor U7541 (N_7541,N_6830,N_6723);
or U7542 (N_7542,N_6893,N_6635);
nor U7543 (N_7543,N_6964,N_6219);
or U7544 (N_7544,N_6741,N_6945);
nor U7545 (N_7545,N_6782,N_6590);
or U7546 (N_7546,N_6109,N_6198);
or U7547 (N_7547,N_6956,N_6049);
nand U7548 (N_7548,N_6336,N_6374);
and U7549 (N_7549,N_6011,N_6131);
and U7550 (N_7550,N_6321,N_6161);
nand U7551 (N_7551,N_6755,N_6627);
nor U7552 (N_7552,N_6820,N_6238);
nor U7553 (N_7553,N_6447,N_6078);
or U7554 (N_7554,N_6960,N_6306);
nand U7555 (N_7555,N_6844,N_6334);
and U7556 (N_7556,N_6485,N_6109);
or U7557 (N_7557,N_6749,N_6909);
nand U7558 (N_7558,N_6418,N_6628);
or U7559 (N_7559,N_6136,N_6681);
and U7560 (N_7560,N_6540,N_6682);
nor U7561 (N_7561,N_6761,N_6006);
and U7562 (N_7562,N_6568,N_6316);
or U7563 (N_7563,N_6778,N_6967);
nand U7564 (N_7564,N_6382,N_6879);
or U7565 (N_7565,N_6955,N_6576);
and U7566 (N_7566,N_6354,N_6428);
nand U7567 (N_7567,N_6932,N_6987);
nor U7568 (N_7568,N_6197,N_6262);
nor U7569 (N_7569,N_6756,N_6284);
nand U7570 (N_7570,N_6857,N_6494);
nor U7571 (N_7571,N_6664,N_6827);
or U7572 (N_7572,N_6508,N_6954);
and U7573 (N_7573,N_6050,N_6884);
and U7574 (N_7574,N_6249,N_6897);
or U7575 (N_7575,N_6347,N_6590);
and U7576 (N_7576,N_6200,N_6866);
or U7577 (N_7577,N_6382,N_6322);
nand U7578 (N_7578,N_6735,N_6149);
nand U7579 (N_7579,N_6372,N_6519);
or U7580 (N_7580,N_6715,N_6882);
nor U7581 (N_7581,N_6715,N_6781);
and U7582 (N_7582,N_6382,N_6428);
nand U7583 (N_7583,N_6642,N_6698);
and U7584 (N_7584,N_6953,N_6384);
nand U7585 (N_7585,N_6784,N_6617);
and U7586 (N_7586,N_6044,N_6801);
nand U7587 (N_7587,N_6770,N_6994);
and U7588 (N_7588,N_6902,N_6083);
nand U7589 (N_7589,N_6043,N_6977);
nor U7590 (N_7590,N_6931,N_6048);
nand U7591 (N_7591,N_6661,N_6250);
or U7592 (N_7592,N_6778,N_6265);
and U7593 (N_7593,N_6289,N_6341);
nand U7594 (N_7594,N_6664,N_6279);
and U7595 (N_7595,N_6394,N_6331);
nor U7596 (N_7596,N_6201,N_6255);
and U7597 (N_7597,N_6823,N_6595);
nand U7598 (N_7598,N_6973,N_6640);
or U7599 (N_7599,N_6618,N_6072);
and U7600 (N_7600,N_6797,N_6741);
and U7601 (N_7601,N_6637,N_6341);
nand U7602 (N_7602,N_6467,N_6992);
or U7603 (N_7603,N_6055,N_6755);
or U7604 (N_7604,N_6512,N_6096);
nand U7605 (N_7605,N_6418,N_6355);
and U7606 (N_7606,N_6977,N_6754);
and U7607 (N_7607,N_6288,N_6725);
or U7608 (N_7608,N_6576,N_6883);
nand U7609 (N_7609,N_6847,N_6457);
and U7610 (N_7610,N_6983,N_6986);
or U7611 (N_7611,N_6888,N_6673);
or U7612 (N_7612,N_6207,N_6694);
and U7613 (N_7613,N_6355,N_6150);
and U7614 (N_7614,N_6315,N_6735);
and U7615 (N_7615,N_6579,N_6421);
or U7616 (N_7616,N_6119,N_6053);
nor U7617 (N_7617,N_6268,N_6161);
nor U7618 (N_7618,N_6193,N_6469);
and U7619 (N_7619,N_6906,N_6789);
and U7620 (N_7620,N_6666,N_6976);
and U7621 (N_7621,N_6653,N_6754);
nand U7622 (N_7622,N_6835,N_6969);
nand U7623 (N_7623,N_6883,N_6566);
or U7624 (N_7624,N_6977,N_6302);
and U7625 (N_7625,N_6126,N_6321);
or U7626 (N_7626,N_6432,N_6150);
nand U7627 (N_7627,N_6787,N_6132);
nand U7628 (N_7628,N_6202,N_6023);
nand U7629 (N_7629,N_6504,N_6436);
nand U7630 (N_7630,N_6292,N_6055);
and U7631 (N_7631,N_6250,N_6078);
and U7632 (N_7632,N_6295,N_6741);
nand U7633 (N_7633,N_6539,N_6408);
nand U7634 (N_7634,N_6222,N_6919);
nor U7635 (N_7635,N_6963,N_6841);
nor U7636 (N_7636,N_6144,N_6031);
nor U7637 (N_7637,N_6568,N_6488);
or U7638 (N_7638,N_6547,N_6614);
nand U7639 (N_7639,N_6793,N_6874);
nor U7640 (N_7640,N_6633,N_6439);
nand U7641 (N_7641,N_6915,N_6685);
or U7642 (N_7642,N_6184,N_6583);
nor U7643 (N_7643,N_6181,N_6821);
and U7644 (N_7644,N_6836,N_6645);
nand U7645 (N_7645,N_6596,N_6637);
or U7646 (N_7646,N_6255,N_6960);
nand U7647 (N_7647,N_6471,N_6531);
nand U7648 (N_7648,N_6490,N_6359);
and U7649 (N_7649,N_6802,N_6555);
and U7650 (N_7650,N_6109,N_6246);
nand U7651 (N_7651,N_6151,N_6285);
and U7652 (N_7652,N_6201,N_6780);
nand U7653 (N_7653,N_6728,N_6673);
nor U7654 (N_7654,N_6454,N_6826);
or U7655 (N_7655,N_6888,N_6156);
or U7656 (N_7656,N_6704,N_6134);
nand U7657 (N_7657,N_6865,N_6787);
or U7658 (N_7658,N_6825,N_6530);
or U7659 (N_7659,N_6692,N_6890);
nand U7660 (N_7660,N_6517,N_6795);
or U7661 (N_7661,N_6401,N_6722);
and U7662 (N_7662,N_6225,N_6257);
and U7663 (N_7663,N_6346,N_6433);
and U7664 (N_7664,N_6157,N_6044);
or U7665 (N_7665,N_6766,N_6431);
nand U7666 (N_7666,N_6067,N_6735);
nor U7667 (N_7667,N_6446,N_6046);
or U7668 (N_7668,N_6625,N_6624);
or U7669 (N_7669,N_6387,N_6907);
and U7670 (N_7670,N_6078,N_6218);
and U7671 (N_7671,N_6365,N_6606);
and U7672 (N_7672,N_6259,N_6292);
nand U7673 (N_7673,N_6244,N_6293);
nor U7674 (N_7674,N_6975,N_6481);
and U7675 (N_7675,N_6567,N_6445);
and U7676 (N_7676,N_6731,N_6427);
nand U7677 (N_7677,N_6474,N_6484);
or U7678 (N_7678,N_6388,N_6138);
and U7679 (N_7679,N_6483,N_6292);
nor U7680 (N_7680,N_6889,N_6032);
nand U7681 (N_7681,N_6510,N_6952);
nand U7682 (N_7682,N_6122,N_6641);
nor U7683 (N_7683,N_6335,N_6276);
nand U7684 (N_7684,N_6522,N_6574);
nand U7685 (N_7685,N_6917,N_6706);
nor U7686 (N_7686,N_6860,N_6439);
nor U7687 (N_7687,N_6819,N_6332);
or U7688 (N_7688,N_6857,N_6825);
nand U7689 (N_7689,N_6685,N_6565);
nor U7690 (N_7690,N_6690,N_6049);
nand U7691 (N_7691,N_6470,N_6103);
or U7692 (N_7692,N_6830,N_6210);
nor U7693 (N_7693,N_6388,N_6411);
or U7694 (N_7694,N_6868,N_6999);
and U7695 (N_7695,N_6814,N_6146);
nor U7696 (N_7696,N_6166,N_6643);
nand U7697 (N_7697,N_6973,N_6295);
or U7698 (N_7698,N_6139,N_6201);
nand U7699 (N_7699,N_6050,N_6976);
nor U7700 (N_7700,N_6033,N_6874);
or U7701 (N_7701,N_6169,N_6873);
or U7702 (N_7702,N_6215,N_6824);
or U7703 (N_7703,N_6651,N_6870);
and U7704 (N_7704,N_6266,N_6957);
nor U7705 (N_7705,N_6253,N_6666);
nand U7706 (N_7706,N_6305,N_6674);
and U7707 (N_7707,N_6713,N_6851);
nor U7708 (N_7708,N_6690,N_6917);
nor U7709 (N_7709,N_6351,N_6172);
nand U7710 (N_7710,N_6968,N_6662);
nand U7711 (N_7711,N_6277,N_6175);
nand U7712 (N_7712,N_6262,N_6875);
nand U7713 (N_7713,N_6852,N_6618);
or U7714 (N_7714,N_6239,N_6057);
nand U7715 (N_7715,N_6824,N_6123);
nand U7716 (N_7716,N_6628,N_6775);
nand U7717 (N_7717,N_6676,N_6677);
or U7718 (N_7718,N_6184,N_6279);
or U7719 (N_7719,N_6843,N_6366);
nor U7720 (N_7720,N_6847,N_6888);
nor U7721 (N_7721,N_6018,N_6957);
nor U7722 (N_7722,N_6357,N_6514);
and U7723 (N_7723,N_6178,N_6677);
and U7724 (N_7724,N_6021,N_6179);
and U7725 (N_7725,N_6879,N_6200);
nand U7726 (N_7726,N_6236,N_6736);
or U7727 (N_7727,N_6075,N_6009);
nor U7728 (N_7728,N_6597,N_6134);
nand U7729 (N_7729,N_6032,N_6824);
and U7730 (N_7730,N_6885,N_6191);
or U7731 (N_7731,N_6394,N_6743);
and U7732 (N_7732,N_6633,N_6389);
nor U7733 (N_7733,N_6578,N_6424);
nor U7734 (N_7734,N_6427,N_6010);
nor U7735 (N_7735,N_6133,N_6552);
or U7736 (N_7736,N_6006,N_6219);
nand U7737 (N_7737,N_6049,N_6900);
nor U7738 (N_7738,N_6531,N_6042);
nand U7739 (N_7739,N_6993,N_6231);
nor U7740 (N_7740,N_6546,N_6221);
nand U7741 (N_7741,N_6370,N_6090);
and U7742 (N_7742,N_6752,N_6710);
and U7743 (N_7743,N_6297,N_6837);
nor U7744 (N_7744,N_6629,N_6778);
or U7745 (N_7745,N_6773,N_6115);
or U7746 (N_7746,N_6569,N_6822);
and U7747 (N_7747,N_6683,N_6546);
and U7748 (N_7748,N_6313,N_6807);
and U7749 (N_7749,N_6539,N_6610);
nor U7750 (N_7750,N_6468,N_6675);
or U7751 (N_7751,N_6833,N_6287);
nor U7752 (N_7752,N_6483,N_6120);
or U7753 (N_7753,N_6463,N_6223);
or U7754 (N_7754,N_6111,N_6537);
nor U7755 (N_7755,N_6552,N_6807);
or U7756 (N_7756,N_6550,N_6276);
and U7757 (N_7757,N_6402,N_6284);
nand U7758 (N_7758,N_6956,N_6034);
nor U7759 (N_7759,N_6178,N_6868);
nand U7760 (N_7760,N_6982,N_6080);
nand U7761 (N_7761,N_6717,N_6924);
nor U7762 (N_7762,N_6567,N_6098);
nand U7763 (N_7763,N_6178,N_6060);
or U7764 (N_7764,N_6699,N_6744);
and U7765 (N_7765,N_6660,N_6743);
nand U7766 (N_7766,N_6321,N_6011);
nor U7767 (N_7767,N_6647,N_6473);
or U7768 (N_7768,N_6193,N_6807);
or U7769 (N_7769,N_6781,N_6146);
nand U7770 (N_7770,N_6338,N_6534);
nand U7771 (N_7771,N_6999,N_6834);
or U7772 (N_7772,N_6505,N_6076);
nor U7773 (N_7773,N_6996,N_6726);
nor U7774 (N_7774,N_6126,N_6934);
or U7775 (N_7775,N_6358,N_6463);
nor U7776 (N_7776,N_6889,N_6920);
or U7777 (N_7777,N_6405,N_6755);
or U7778 (N_7778,N_6047,N_6970);
or U7779 (N_7779,N_6964,N_6685);
or U7780 (N_7780,N_6002,N_6893);
nor U7781 (N_7781,N_6520,N_6629);
nor U7782 (N_7782,N_6488,N_6356);
or U7783 (N_7783,N_6358,N_6466);
or U7784 (N_7784,N_6468,N_6416);
or U7785 (N_7785,N_6736,N_6620);
or U7786 (N_7786,N_6158,N_6411);
nand U7787 (N_7787,N_6834,N_6484);
and U7788 (N_7788,N_6832,N_6990);
nor U7789 (N_7789,N_6755,N_6564);
xor U7790 (N_7790,N_6029,N_6984);
nor U7791 (N_7791,N_6201,N_6279);
or U7792 (N_7792,N_6310,N_6262);
nor U7793 (N_7793,N_6211,N_6207);
nor U7794 (N_7794,N_6600,N_6151);
and U7795 (N_7795,N_6762,N_6122);
and U7796 (N_7796,N_6192,N_6787);
and U7797 (N_7797,N_6287,N_6239);
or U7798 (N_7798,N_6903,N_6432);
or U7799 (N_7799,N_6369,N_6081);
or U7800 (N_7800,N_6811,N_6931);
nor U7801 (N_7801,N_6339,N_6081);
nand U7802 (N_7802,N_6078,N_6827);
nand U7803 (N_7803,N_6096,N_6545);
nand U7804 (N_7804,N_6358,N_6803);
nor U7805 (N_7805,N_6140,N_6022);
nand U7806 (N_7806,N_6253,N_6298);
nand U7807 (N_7807,N_6998,N_6486);
nand U7808 (N_7808,N_6345,N_6168);
nor U7809 (N_7809,N_6850,N_6653);
or U7810 (N_7810,N_6072,N_6891);
and U7811 (N_7811,N_6251,N_6477);
or U7812 (N_7812,N_6062,N_6557);
nand U7813 (N_7813,N_6636,N_6186);
nand U7814 (N_7814,N_6216,N_6046);
and U7815 (N_7815,N_6317,N_6995);
nor U7816 (N_7816,N_6318,N_6194);
nor U7817 (N_7817,N_6804,N_6686);
or U7818 (N_7818,N_6352,N_6240);
nand U7819 (N_7819,N_6030,N_6745);
and U7820 (N_7820,N_6526,N_6898);
or U7821 (N_7821,N_6410,N_6606);
nor U7822 (N_7822,N_6638,N_6106);
or U7823 (N_7823,N_6427,N_6541);
or U7824 (N_7824,N_6299,N_6150);
nor U7825 (N_7825,N_6419,N_6439);
nand U7826 (N_7826,N_6637,N_6540);
nand U7827 (N_7827,N_6216,N_6805);
or U7828 (N_7828,N_6710,N_6791);
and U7829 (N_7829,N_6126,N_6424);
nor U7830 (N_7830,N_6866,N_6702);
and U7831 (N_7831,N_6685,N_6958);
or U7832 (N_7832,N_6638,N_6507);
nor U7833 (N_7833,N_6319,N_6648);
and U7834 (N_7834,N_6254,N_6246);
or U7835 (N_7835,N_6775,N_6122);
or U7836 (N_7836,N_6875,N_6970);
or U7837 (N_7837,N_6871,N_6109);
xor U7838 (N_7838,N_6694,N_6382);
nor U7839 (N_7839,N_6192,N_6735);
and U7840 (N_7840,N_6199,N_6643);
or U7841 (N_7841,N_6174,N_6718);
and U7842 (N_7842,N_6874,N_6292);
and U7843 (N_7843,N_6884,N_6699);
nand U7844 (N_7844,N_6343,N_6223);
nand U7845 (N_7845,N_6186,N_6207);
and U7846 (N_7846,N_6729,N_6848);
nor U7847 (N_7847,N_6717,N_6499);
or U7848 (N_7848,N_6935,N_6827);
nor U7849 (N_7849,N_6618,N_6776);
and U7850 (N_7850,N_6441,N_6401);
nor U7851 (N_7851,N_6924,N_6203);
nand U7852 (N_7852,N_6419,N_6066);
and U7853 (N_7853,N_6724,N_6391);
or U7854 (N_7854,N_6596,N_6438);
nand U7855 (N_7855,N_6598,N_6645);
or U7856 (N_7856,N_6666,N_6143);
or U7857 (N_7857,N_6163,N_6540);
and U7858 (N_7858,N_6062,N_6854);
nor U7859 (N_7859,N_6203,N_6898);
or U7860 (N_7860,N_6092,N_6622);
or U7861 (N_7861,N_6503,N_6360);
nand U7862 (N_7862,N_6429,N_6688);
or U7863 (N_7863,N_6410,N_6236);
nand U7864 (N_7864,N_6751,N_6596);
nor U7865 (N_7865,N_6805,N_6990);
nand U7866 (N_7866,N_6397,N_6244);
or U7867 (N_7867,N_6971,N_6456);
nand U7868 (N_7868,N_6873,N_6034);
nor U7869 (N_7869,N_6971,N_6294);
or U7870 (N_7870,N_6751,N_6732);
or U7871 (N_7871,N_6418,N_6336);
nor U7872 (N_7872,N_6582,N_6600);
or U7873 (N_7873,N_6071,N_6577);
and U7874 (N_7874,N_6076,N_6492);
and U7875 (N_7875,N_6433,N_6800);
or U7876 (N_7876,N_6413,N_6046);
nand U7877 (N_7877,N_6212,N_6300);
nor U7878 (N_7878,N_6759,N_6500);
and U7879 (N_7879,N_6833,N_6118);
nand U7880 (N_7880,N_6345,N_6046);
and U7881 (N_7881,N_6298,N_6072);
or U7882 (N_7882,N_6092,N_6197);
or U7883 (N_7883,N_6806,N_6829);
nand U7884 (N_7884,N_6928,N_6880);
nor U7885 (N_7885,N_6511,N_6283);
and U7886 (N_7886,N_6339,N_6070);
nand U7887 (N_7887,N_6309,N_6121);
or U7888 (N_7888,N_6805,N_6871);
nor U7889 (N_7889,N_6286,N_6547);
or U7890 (N_7890,N_6764,N_6164);
or U7891 (N_7891,N_6287,N_6439);
nand U7892 (N_7892,N_6424,N_6517);
and U7893 (N_7893,N_6840,N_6580);
and U7894 (N_7894,N_6762,N_6321);
nand U7895 (N_7895,N_6766,N_6095);
nor U7896 (N_7896,N_6609,N_6388);
nand U7897 (N_7897,N_6153,N_6529);
and U7898 (N_7898,N_6218,N_6225);
or U7899 (N_7899,N_6488,N_6896);
and U7900 (N_7900,N_6515,N_6321);
nand U7901 (N_7901,N_6379,N_6336);
or U7902 (N_7902,N_6722,N_6323);
nor U7903 (N_7903,N_6656,N_6110);
nand U7904 (N_7904,N_6886,N_6138);
nor U7905 (N_7905,N_6737,N_6736);
nand U7906 (N_7906,N_6418,N_6333);
xnor U7907 (N_7907,N_6078,N_6333);
nor U7908 (N_7908,N_6456,N_6780);
and U7909 (N_7909,N_6528,N_6382);
or U7910 (N_7910,N_6700,N_6393);
nand U7911 (N_7911,N_6488,N_6074);
or U7912 (N_7912,N_6367,N_6612);
and U7913 (N_7913,N_6510,N_6523);
nand U7914 (N_7914,N_6294,N_6962);
nor U7915 (N_7915,N_6592,N_6590);
and U7916 (N_7916,N_6789,N_6651);
nand U7917 (N_7917,N_6323,N_6885);
nor U7918 (N_7918,N_6450,N_6197);
nor U7919 (N_7919,N_6109,N_6786);
nor U7920 (N_7920,N_6230,N_6053);
and U7921 (N_7921,N_6462,N_6658);
xnor U7922 (N_7922,N_6339,N_6148);
or U7923 (N_7923,N_6894,N_6700);
and U7924 (N_7924,N_6001,N_6141);
and U7925 (N_7925,N_6072,N_6753);
and U7926 (N_7926,N_6694,N_6475);
nor U7927 (N_7927,N_6085,N_6359);
nor U7928 (N_7928,N_6651,N_6598);
and U7929 (N_7929,N_6390,N_6340);
nor U7930 (N_7930,N_6030,N_6754);
or U7931 (N_7931,N_6615,N_6899);
nor U7932 (N_7932,N_6432,N_6614);
nand U7933 (N_7933,N_6896,N_6711);
nand U7934 (N_7934,N_6879,N_6102);
nand U7935 (N_7935,N_6072,N_6383);
and U7936 (N_7936,N_6714,N_6227);
nor U7937 (N_7937,N_6456,N_6722);
or U7938 (N_7938,N_6772,N_6521);
and U7939 (N_7939,N_6733,N_6505);
and U7940 (N_7940,N_6369,N_6387);
nor U7941 (N_7941,N_6555,N_6667);
and U7942 (N_7942,N_6820,N_6346);
or U7943 (N_7943,N_6513,N_6588);
nand U7944 (N_7944,N_6481,N_6741);
or U7945 (N_7945,N_6332,N_6597);
nor U7946 (N_7946,N_6706,N_6645);
nor U7947 (N_7947,N_6769,N_6412);
nand U7948 (N_7948,N_6848,N_6858);
nand U7949 (N_7949,N_6026,N_6483);
and U7950 (N_7950,N_6325,N_6093);
or U7951 (N_7951,N_6327,N_6552);
and U7952 (N_7952,N_6435,N_6280);
or U7953 (N_7953,N_6680,N_6218);
and U7954 (N_7954,N_6077,N_6297);
or U7955 (N_7955,N_6191,N_6997);
nand U7956 (N_7956,N_6764,N_6012);
nand U7957 (N_7957,N_6846,N_6953);
and U7958 (N_7958,N_6462,N_6221);
nor U7959 (N_7959,N_6276,N_6163);
nand U7960 (N_7960,N_6540,N_6255);
or U7961 (N_7961,N_6737,N_6934);
nand U7962 (N_7962,N_6365,N_6785);
nand U7963 (N_7963,N_6938,N_6791);
nand U7964 (N_7964,N_6899,N_6371);
nand U7965 (N_7965,N_6434,N_6464);
nor U7966 (N_7966,N_6475,N_6771);
nor U7967 (N_7967,N_6087,N_6339);
nor U7968 (N_7968,N_6418,N_6273);
or U7969 (N_7969,N_6488,N_6834);
and U7970 (N_7970,N_6994,N_6999);
nor U7971 (N_7971,N_6133,N_6627);
nor U7972 (N_7972,N_6836,N_6650);
nand U7973 (N_7973,N_6234,N_6185);
and U7974 (N_7974,N_6194,N_6078);
nor U7975 (N_7975,N_6806,N_6651);
nor U7976 (N_7976,N_6251,N_6827);
nand U7977 (N_7977,N_6267,N_6680);
nor U7978 (N_7978,N_6097,N_6207);
and U7979 (N_7979,N_6263,N_6319);
and U7980 (N_7980,N_6785,N_6305);
or U7981 (N_7981,N_6071,N_6681);
nor U7982 (N_7982,N_6976,N_6624);
nand U7983 (N_7983,N_6300,N_6100);
nor U7984 (N_7984,N_6329,N_6047);
or U7985 (N_7985,N_6075,N_6358);
or U7986 (N_7986,N_6301,N_6360);
or U7987 (N_7987,N_6500,N_6755);
nor U7988 (N_7988,N_6009,N_6498);
nor U7989 (N_7989,N_6489,N_6633);
or U7990 (N_7990,N_6387,N_6386);
and U7991 (N_7991,N_6110,N_6950);
nor U7992 (N_7992,N_6374,N_6387);
or U7993 (N_7993,N_6646,N_6140);
or U7994 (N_7994,N_6219,N_6301);
nand U7995 (N_7995,N_6616,N_6316);
or U7996 (N_7996,N_6501,N_6502);
or U7997 (N_7997,N_6137,N_6715);
nand U7998 (N_7998,N_6983,N_6622);
and U7999 (N_7999,N_6185,N_6563);
nand U8000 (N_8000,N_7195,N_7514);
or U8001 (N_8001,N_7207,N_7430);
and U8002 (N_8002,N_7062,N_7804);
nor U8003 (N_8003,N_7915,N_7972);
nand U8004 (N_8004,N_7864,N_7640);
and U8005 (N_8005,N_7531,N_7180);
nor U8006 (N_8006,N_7811,N_7439);
or U8007 (N_8007,N_7599,N_7923);
and U8008 (N_8008,N_7757,N_7367);
and U8009 (N_8009,N_7803,N_7316);
or U8010 (N_8010,N_7419,N_7620);
nand U8011 (N_8011,N_7097,N_7454);
or U8012 (N_8012,N_7604,N_7641);
and U8013 (N_8013,N_7572,N_7643);
nand U8014 (N_8014,N_7036,N_7224);
and U8015 (N_8015,N_7996,N_7626);
nand U8016 (N_8016,N_7621,N_7472);
nor U8017 (N_8017,N_7593,N_7529);
or U8018 (N_8018,N_7382,N_7606);
and U8019 (N_8019,N_7897,N_7739);
or U8020 (N_8020,N_7326,N_7515);
or U8021 (N_8021,N_7041,N_7007);
or U8022 (N_8022,N_7910,N_7063);
or U8023 (N_8023,N_7901,N_7185);
and U8024 (N_8024,N_7863,N_7563);
or U8025 (N_8025,N_7171,N_7331);
and U8026 (N_8026,N_7278,N_7882);
or U8027 (N_8027,N_7345,N_7952);
nand U8028 (N_8028,N_7833,N_7627);
nand U8029 (N_8029,N_7784,N_7204);
or U8030 (N_8030,N_7905,N_7929);
nand U8031 (N_8031,N_7705,N_7780);
nor U8032 (N_8032,N_7076,N_7302);
nor U8033 (N_8033,N_7000,N_7383);
nand U8034 (N_8034,N_7168,N_7526);
nand U8035 (N_8035,N_7269,N_7501);
nor U8036 (N_8036,N_7338,N_7610);
nand U8037 (N_8037,N_7649,N_7843);
nand U8038 (N_8038,N_7642,N_7675);
nor U8039 (N_8039,N_7039,N_7995);
and U8040 (N_8040,N_7264,N_7979);
nor U8041 (N_8041,N_7286,N_7143);
and U8042 (N_8042,N_7065,N_7712);
or U8043 (N_8043,N_7157,N_7392);
nand U8044 (N_8044,N_7416,N_7552);
nand U8045 (N_8045,N_7442,N_7777);
and U8046 (N_8046,N_7384,N_7032);
nor U8047 (N_8047,N_7744,N_7186);
xor U8048 (N_8048,N_7453,N_7296);
and U8049 (N_8049,N_7589,N_7105);
nor U8050 (N_8050,N_7609,N_7239);
nor U8051 (N_8051,N_7455,N_7769);
or U8052 (N_8052,N_7001,N_7730);
nand U8053 (N_8053,N_7482,N_7216);
nand U8054 (N_8054,N_7436,N_7877);
or U8055 (N_8055,N_7115,N_7376);
and U8056 (N_8056,N_7258,N_7361);
nand U8057 (N_8057,N_7432,N_7054);
nor U8058 (N_8058,N_7665,N_7962);
nand U8059 (N_8059,N_7879,N_7179);
nor U8060 (N_8060,N_7591,N_7373);
and U8061 (N_8061,N_7549,N_7561);
or U8062 (N_8062,N_7834,N_7584);
nand U8063 (N_8063,N_7938,N_7861);
nor U8064 (N_8064,N_7745,N_7406);
and U8065 (N_8065,N_7141,N_7551);
and U8066 (N_8066,N_7029,N_7114);
or U8067 (N_8067,N_7695,N_7876);
nand U8068 (N_8068,N_7789,N_7403);
nor U8069 (N_8069,N_7410,N_7613);
nor U8070 (N_8070,N_7955,N_7071);
or U8071 (N_8071,N_7449,N_7174);
nand U8072 (N_8072,N_7360,N_7639);
nand U8073 (N_8073,N_7450,N_7960);
nand U8074 (N_8074,N_7722,N_7600);
nor U8075 (N_8075,N_7458,N_7898);
or U8076 (N_8076,N_7701,N_7238);
and U8077 (N_8077,N_7451,N_7860);
nor U8078 (N_8078,N_7129,N_7816);
and U8079 (N_8079,N_7194,N_7243);
or U8080 (N_8080,N_7033,N_7577);
or U8081 (N_8081,N_7220,N_7354);
nand U8082 (N_8082,N_7500,N_7127);
or U8083 (N_8083,N_7907,N_7287);
or U8084 (N_8084,N_7902,N_7913);
and U8085 (N_8085,N_7256,N_7528);
nand U8086 (N_8086,N_7149,N_7737);
nand U8087 (N_8087,N_7741,N_7330);
or U8088 (N_8088,N_7104,N_7301);
nand U8089 (N_8089,N_7130,N_7255);
or U8090 (N_8090,N_7058,N_7930);
and U8091 (N_8091,N_7724,N_7344);
or U8092 (N_8092,N_7018,N_7181);
nor U8093 (N_8093,N_7003,N_7377);
nand U8094 (N_8094,N_7132,N_7766);
nand U8095 (N_8095,N_7651,N_7006);
nor U8096 (N_8096,N_7415,N_7874);
or U8097 (N_8097,N_7554,N_7327);
nor U8098 (N_8098,N_7489,N_7478);
and U8099 (N_8099,N_7035,N_7070);
nor U8100 (N_8100,N_7564,N_7959);
nand U8101 (N_8101,N_7203,N_7173);
nand U8102 (N_8102,N_7773,N_7775);
and U8103 (N_8103,N_7004,N_7813);
nor U8104 (N_8104,N_7755,N_7088);
or U8105 (N_8105,N_7809,N_7618);
and U8106 (N_8106,N_7965,N_7854);
and U8107 (N_8107,N_7922,N_7994);
nand U8108 (N_8108,N_7184,N_7867);
xnor U8109 (N_8109,N_7468,N_7349);
nand U8110 (N_8110,N_7120,N_7289);
or U8111 (N_8111,N_7119,N_7556);
and U8112 (N_8112,N_7140,N_7732);
nor U8113 (N_8113,N_7025,N_7365);
or U8114 (N_8114,N_7582,N_7571);
and U8115 (N_8115,N_7051,N_7037);
nand U8116 (N_8116,N_7507,N_7303);
nor U8117 (N_8117,N_7555,N_7534);
nand U8118 (N_8118,N_7425,N_7562);
or U8119 (N_8119,N_7221,N_7026);
and U8120 (N_8120,N_7219,N_7490);
and U8121 (N_8121,N_7064,N_7662);
or U8122 (N_8122,N_7474,N_7652);
and U8123 (N_8123,N_7678,N_7723);
nor U8124 (N_8124,N_7926,N_7801);
or U8125 (N_8125,N_7550,N_7142);
or U8126 (N_8126,N_7683,N_7945);
and U8127 (N_8127,N_7704,N_7259);
or U8128 (N_8128,N_7329,N_7304);
nor U8129 (N_8129,N_7237,N_7366);
and U8130 (N_8130,N_7738,N_7940);
and U8131 (N_8131,N_7570,N_7061);
xor U8132 (N_8132,N_7205,N_7291);
nor U8133 (N_8133,N_7012,N_7399);
nand U8134 (N_8134,N_7873,N_7820);
and U8135 (N_8135,N_7313,N_7791);
nor U8136 (N_8136,N_7282,N_7397);
nor U8137 (N_8137,N_7167,N_7856);
nand U8138 (N_8138,N_7163,N_7423);
and U8139 (N_8139,N_7660,N_7587);
nand U8140 (N_8140,N_7548,N_7608);
or U8141 (N_8141,N_7969,N_7958);
and U8142 (N_8142,N_7146,N_7912);
and U8143 (N_8143,N_7187,N_7761);
or U8144 (N_8144,N_7839,N_7977);
nand U8145 (N_8145,N_7588,N_7160);
and U8146 (N_8146,N_7031,N_7275);
nand U8147 (N_8147,N_7014,N_7395);
nor U8148 (N_8148,N_7385,N_7433);
or U8149 (N_8149,N_7305,N_7916);
or U8150 (N_8150,N_7797,N_7199);
nor U8151 (N_8151,N_7435,N_7772);
and U8152 (N_8152,N_7404,N_7725);
nor U8153 (N_8153,N_7402,N_7583);
nor U8154 (N_8154,N_7829,N_7324);
nand U8155 (N_8155,N_7764,N_7437);
and U8156 (N_8156,N_7073,N_7679);
nor U8157 (N_8157,N_7663,N_7892);
nand U8158 (N_8158,N_7631,N_7246);
or U8159 (N_8159,N_7248,N_7153);
or U8160 (N_8160,N_7218,N_7189);
nand U8161 (N_8161,N_7318,N_7527);
or U8162 (N_8162,N_7310,N_7821);
nand U8163 (N_8163,N_7295,N_7576);
or U8164 (N_8164,N_7636,N_7240);
nand U8165 (N_8165,N_7893,N_7615);
or U8166 (N_8166,N_7699,N_7823);
nor U8167 (N_8167,N_7537,N_7400);
and U8168 (N_8168,N_7447,N_7968);
xnor U8169 (N_8169,N_7920,N_7847);
or U8170 (N_8170,N_7806,N_7147);
nor U8171 (N_8171,N_7352,N_7680);
nor U8172 (N_8172,N_7546,N_7818);
nor U8173 (N_8173,N_7628,N_7111);
and U8174 (N_8174,N_7637,N_7708);
or U8175 (N_8175,N_7710,N_7312);
and U8176 (N_8176,N_7525,N_7340);
or U8177 (N_8177,N_7545,N_7494);
and U8178 (N_8178,N_7081,N_7558);
and U8179 (N_8179,N_7429,N_7573);
and U8180 (N_8180,N_7779,N_7949);
nand U8181 (N_8181,N_7414,N_7428);
nand U8182 (N_8182,N_7050,N_7785);
nor U8183 (N_8183,N_7826,N_7267);
and U8184 (N_8184,N_7096,N_7547);
nand U8185 (N_8185,N_7372,N_7647);
and U8186 (N_8186,N_7603,N_7696);
and U8187 (N_8187,N_7524,N_7578);
or U8188 (N_8188,N_7049,N_7434);
nand U8189 (N_8189,N_7630,N_7850);
nand U8190 (N_8190,N_7445,N_7391);
nor U8191 (N_8191,N_7731,N_7464);
or U8192 (N_8192,N_7060,N_7518);
or U8193 (N_8193,N_7013,N_7164);
nand U8194 (N_8194,N_7162,N_7832);
nor U8195 (N_8195,N_7426,N_7544);
or U8196 (N_8196,N_7894,N_7542);
and U8197 (N_8197,N_7767,N_7093);
and U8198 (N_8198,N_7477,N_7734);
nor U8199 (N_8199,N_7274,N_7212);
or U8200 (N_8200,N_7418,N_7914);
nand U8201 (N_8201,N_7668,N_7904);
nor U8202 (N_8202,N_7565,N_7311);
or U8203 (N_8203,N_7984,N_7686);
nor U8204 (N_8204,N_7814,N_7134);
and U8205 (N_8205,N_7353,N_7133);
or U8206 (N_8206,N_7598,N_7412);
or U8207 (N_8207,N_7188,N_7332);
nand U8208 (N_8208,N_7333,N_7456);
xor U8209 (N_8209,N_7491,N_7232);
and U8210 (N_8210,N_7090,N_7891);
and U8211 (N_8211,N_7646,N_7702);
nor U8212 (N_8212,N_7911,N_7497);
nand U8213 (N_8213,N_7106,N_7198);
nor U8214 (N_8214,N_7431,N_7137);
and U8215 (N_8215,N_7213,N_7844);
and U8216 (N_8216,N_7981,N_7244);
or U8217 (N_8217,N_7749,N_7499);
or U8218 (N_8218,N_7225,N_7231);
and U8219 (N_8219,N_7317,N_7448);
nand U8220 (N_8220,N_7721,N_7250);
nor U8221 (N_8221,N_7091,N_7192);
or U8222 (N_8222,N_7228,N_7590);
nor U8223 (N_8223,N_7299,N_7768);
or U8224 (N_8224,N_7043,N_7175);
or U8225 (N_8225,N_7954,N_7602);
nor U8226 (N_8226,N_7040,N_7953);
nand U8227 (N_8227,N_7211,N_7300);
nand U8228 (N_8228,N_7817,N_7862);
and U8229 (N_8229,N_7698,N_7375);
or U8230 (N_8230,N_7023,N_7424);
or U8231 (N_8231,N_7530,N_7670);
nand U8232 (N_8232,N_7233,N_7476);
nand U8233 (N_8233,N_7417,N_7917);
and U8234 (N_8234,N_7539,N_7123);
nor U8235 (N_8235,N_7144,N_7245);
or U8236 (N_8236,N_7271,N_7511);
and U8237 (N_8237,N_7633,N_7082);
and U8238 (N_8238,N_7463,N_7692);
nand U8239 (N_8239,N_7852,N_7285);
and U8240 (N_8240,N_7151,N_7771);
nand U8241 (N_8241,N_7293,N_7321);
nor U8242 (N_8242,N_7934,N_7294);
nand U8243 (N_8243,N_7002,N_7971);
or U8244 (N_8244,N_7235,N_7292);
or U8245 (N_8245,N_7654,N_7498);
nor U8246 (N_8246,N_7343,N_7650);
and U8247 (N_8247,N_7206,N_7438);
nand U8248 (N_8248,N_7579,N_7394);
nand U8249 (N_8249,N_7249,N_7095);
nor U8250 (N_8250,N_7569,N_7541);
nand U8251 (N_8251,N_7975,N_7276);
or U8252 (N_8252,N_7510,N_7100);
nand U8253 (N_8253,N_7170,N_7196);
and U8254 (N_8254,N_7657,N_7878);
nor U8255 (N_8255,N_7523,N_7900);
and U8256 (N_8256,N_7191,N_7964);
and U8257 (N_8257,N_7348,N_7272);
or U8258 (N_8258,N_7733,N_7297);
nor U8259 (N_8259,N_7655,N_7596);
or U8260 (N_8260,N_7896,N_7728);
or U8261 (N_8261,N_7841,N_7629);
or U8262 (N_8262,N_7568,N_7800);
and U8263 (N_8263,N_7751,N_7208);
nand U8264 (N_8264,N_7812,N_7217);
nor U8265 (N_8265,N_7616,N_7842);
xor U8266 (N_8266,N_7420,N_7674);
and U8267 (N_8267,N_7016,N_7935);
nor U8268 (N_8268,N_7103,N_7931);
or U8269 (N_8269,N_7939,N_7988);
or U8270 (N_8270,N_7488,N_7796);
and U8271 (N_8271,N_7729,N_7786);
and U8272 (N_8272,N_7595,N_7411);
and U8273 (N_8273,N_7347,N_7281);
nand U8274 (N_8274,N_7830,N_7284);
nand U8275 (N_8275,N_7161,N_7697);
and U8276 (N_8276,N_7280,N_7625);
nand U8277 (N_8277,N_7355,N_7156);
and U8278 (N_8278,N_7109,N_7921);
or U8279 (N_8279,N_7906,N_7774);
or U8280 (N_8280,N_7943,N_7009);
nand U8281 (N_8281,N_7325,N_7622);
and U8282 (N_8282,N_7553,N_7866);
nor U8283 (N_8283,N_7740,N_7089);
or U8284 (N_8284,N_7266,N_7941);
nor U8285 (N_8285,N_7201,N_7855);
nand U8286 (N_8286,N_7838,N_7747);
nor U8287 (N_8287,N_7234,N_7822);
nand U8288 (N_8288,N_7516,N_7320);
nor U8289 (N_8289,N_7251,N_7759);
xor U8290 (N_8290,N_7987,N_7241);
nor U8291 (N_8291,N_7015,N_7682);
or U8292 (N_8292,N_7480,N_7306);
nand U8293 (N_8293,N_7193,N_7427);
or U8294 (N_8294,N_7085,N_7351);
nor U8295 (N_8295,N_7807,N_7495);
and U8296 (N_8296,N_7446,N_7750);
and U8297 (N_8297,N_7661,N_7262);
or U8298 (N_8298,N_7986,N_7356);
nand U8299 (N_8299,N_7831,N_7369);
nand U8300 (N_8300,N_7337,N_7145);
nor U8301 (N_8301,N_7967,N_7909);
nor U8302 (N_8302,N_7046,N_7890);
nand U8303 (N_8303,N_7336,N_7288);
nand U8304 (N_8304,N_7452,N_7094);
nor U8305 (N_8305,N_7681,N_7078);
nand U8306 (N_8306,N_7098,N_7635);
or U8307 (N_8307,N_7308,N_7936);
or U8308 (N_8308,N_7273,N_7925);
nor U8309 (N_8309,N_7005,N_7961);
and U8310 (N_8310,N_7440,N_7574);
nor U8311 (N_8311,N_7462,N_7580);
and U8312 (N_8312,N_7357,N_7644);
nand U8313 (N_8313,N_7341,N_7763);
nand U8314 (N_8314,N_7475,N_7172);
and U8315 (N_8315,N_7027,N_7148);
or U8316 (N_8316,N_7080,N_7700);
or U8317 (N_8317,N_7885,N_7887);
nor U8318 (N_8318,N_7042,N_7052);
or U8319 (N_8319,N_7795,N_7837);
nand U8320 (N_8320,N_7077,N_7648);
xor U8321 (N_8321,N_7787,N_7793);
nor U8322 (N_8322,N_7623,N_7719);
or U8323 (N_8323,N_7364,N_7932);
and U8324 (N_8324,N_7017,N_7703);
nand U8325 (N_8325,N_7512,N_7607);
or U8326 (N_8326,N_7790,N_7496);
nand U8327 (N_8327,N_7277,N_7152);
nand U8328 (N_8328,N_7669,N_7517);
and U8329 (N_8329,N_7122,N_7223);
nand U8330 (N_8330,N_7484,N_7976);
or U8331 (N_8331,N_7502,N_7815);
nor U8332 (N_8332,N_7688,N_7942);
and U8333 (N_8333,N_7084,N_7467);
and U8334 (N_8334,N_7726,N_7328);
nor U8335 (N_8335,N_7401,N_7108);
and U8336 (N_8336,N_7533,N_7117);
nor U8337 (N_8337,N_7136,N_7532);
or U8338 (N_8338,N_7835,N_7656);
nand U8339 (N_8339,N_7083,N_7853);
or U8340 (N_8340,N_7808,N_7155);
nor U8341 (N_8341,N_7038,N_7956);
nor U8342 (N_8342,N_7200,N_7851);
and U8343 (N_8343,N_7736,N_7825);
nor U8344 (N_8344,N_7290,N_7581);
or U8345 (N_8345,N_7664,N_7560);
or U8346 (N_8346,N_7727,N_7226);
nand U8347 (N_8347,N_7752,N_7202);
or U8348 (N_8348,N_7802,N_7983);
and U8349 (N_8349,N_7966,N_7858);
xor U8350 (N_8350,N_7503,N_7677);
nor U8351 (N_8351,N_7210,N_7717);
nor U8352 (N_8352,N_7492,N_7638);
and U8353 (N_8353,N_7443,N_7991);
or U8354 (N_8354,N_7504,N_7535);
nor U8355 (N_8355,N_7718,N_7611);
or U8356 (N_8356,N_7706,N_7884);
nor U8357 (N_8357,N_7742,N_7112);
nor U8358 (N_8358,N_7875,N_7386);
and U8359 (N_8359,N_7261,N_7409);
nor U8360 (N_8360,N_7760,N_7614);
nand U8361 (N_8361,N_7982,N_7265);
nor U8362 (N_8362,N_7444,N_7792);
or U8363 (N_8363,N_7849,N_7045);
or U8364 (N_8364,N_7506,N_7810);
or U8365 (N_8365,N_7519,N_7567);
nand U8366 (N_8366,N_7056,N_7177);
and U8367 (N_8367,N_7178,N_7471);
or U8368 (N_8368,N_7260,N_7099);
or U8369 (N_8369,N_7998,N_7086);
and U8370 (N_8370,N_7252,N_7632);
or U8371 (N_8371,N_7165,N_7992);
and U8372 (N_8372,N_7689,N_7840);
nor U8373 (N_8373,N_7575,N_7948);
nand U8374 (N_8374,N_7776,N_7339);
nand U8375 (N_8375,N_7011,N_7557);
nor U8376 (N_8376,N_7393,N_7270);
and U8377 (N_8377,N_7485,N_7634);
nand U8378 (N_8378,N_7176,N_7322);
or U8379 (N_8379,N_7307,N_7126);
and U8380 (N_8380,N_7978,N_7459);
and U8381 (N_8381,N_7460,N_7585);
nand U8382 (N_8382,N_7389,N_7334);
nand U8383 (N_8383,N_7601,N_7951);
and U8384 (N_8384,N_7346,N_7390);
nand U8385 (N_8385,N_7924,N_7693);
or U8386 (N_8386,N_7315,N_7139);
nand U8387 (N_8387,N_7075,N_7946);
or U8388 (N_8388,N_7024,N_7748);
nand U8389 (N_8389,N_7928,N_7888);
nor U8390 (N_8390,N_7169,N_7520);
nand U8391 (N_8391,N_7253,N_7057);
nor U8392 (N_8392,N_7022,N_7672);
and U8393 (N_8393,N_7881,N_7268);
xor U8394 (N_8394,N_7659,N_7685);
nand U8395 (N_8395,N_7413,N_7461);
nand U8396 (N_8396,N_7101,N_7019);
nor U8397 (N_8397,N_7950,N_7113);
nand U8398 (N_8398,N_7690,N_7379);
or U8399 (N_8399,N_7158,N_7368);
nand U8400 (N_8400,N_7128,N_7465);
nor U8401 (N_8401,N_7487,N_7687);
or U8402 (N_8402,N_7788,N_7869);
nor U8403 (N_8403,N_7957,N_7363);
nor U8404 (N_8404,N_7538,N_7388);
or U8405 (N_8405,N_7848,N_7335);
or U8406 (N_8406,N_7597,N_7422);
nand U8407 (N_8407,N_7694,N_7919);
or U8408 (N_8408,N_7483,N_7230);
nand U8409 (N_8409,N_7684,N_7398);
or U8410 (N_8410,N_7008,N_7824);
and U8411 (N_8411,N_7421,N_7215);
and U8412 (N_8412,N_7342,N_7559);
or U8413 (N_8413,N_7985,N_7138);
or U8414 (N_8414,N_7594,N_7937);
nand U8415 (N_8415,N_7716,N_7154);
nand U8416 (N_8416,N_7845,N_7859);
nand U8417 (N_8417,N_7918,N_7380);
nor U8418 (N_8418,N_7713,N_7229);
or U8419 (N_8419,N_7371,N_7805);
nand U8420 (N_8420,N_7479,N_7989);
nor U8421 (N_8421,N_7067,N_7819);
and U8422 (N_8422,N_7799,N_7214);
and U8423 (N_8423,N_7947,N_7666);
or U8424 (N_8424,N_7150,N_7889);
nor U8425 (N_8425,N_7756,N_7254);
or U8426 (N_8426,N_7754,N_7770);
nand U8427 (N_8427,N_7720,N_7466);
or U8428 (N_8428,N_7323,N_7782);
nor U8429 (N_8429,N_7407,N_7586);
nand U8430 (N_8430,N_7624,N_7159);
nor U8431 (N_8431,N_7059,N_7667);
or U8432 (N_8432,N_7197,N_7072);
nor U8433 (N_8433,N_7746,N_7619);
and U8434 (N_8434,N_7509,N_7974);
nor U8435 (N_8435,N_7107,N_7645);
and U8436 (N_8436,N_7798,N_7118);
or U8437 (N_8437,N_7048,N_7047);
nand U8438 (N_8438,N_7309,N_7359);
or U8439 (N_8439,N_7846,N_7944);
or U8440 (N_8440,N_7980,N_7783);
and U8441 (N_8441,N_7707,N_7883);
nand U8442 (N_8442,N_7079,N_7709);
nand U8443 (N_8443,N_7865,N_7183);
or U8444 (N_8444,N_7711,N_7973);
or U8445 (N_8445,N_7381,N_7350);
or U8446 (N_8446,N_7990,N_7970);
and U8447 (N_8447,N_7933,N_7358);
nand U8448 (N_8448,N_7010,N_7899);
and U8449 (N_8449,N_7469,N_7044);
or U8450 (N_8450,N_7020,N_7762);
and U8451 (N_8451,N_7242,N_7209);
nor U8452 (N_8452,N_7868,N_7676);
nor U8453 (N_8453,N_7521,N_7470);
or U8454 (N_8454,N_7021,N_7370);
or U8455 (N_8455,N_7653,N_7714);
nand U8456 (N_8456,N_7870,N_7658);
nor U8457 (N_8457,N_7999,N_7612);
and U8458 (N_8458,N_7135,N_7473);
nor U8459 (N_8459,N_7396,N_7222);
or U8460 (N_8460,N_7074,N_7110);
or U8461 (N_8461,N_7190,N_7121);
or U8462 (N_8462,N_7508,N_7895);
nor U8463 (N_8463,N_7540,N_7493);
and U8464 (N_8464,N_7124,N_7069);
nor U8465 (N_8465,N_7102,N_7927);
and U8466 (N_8466,N_7378,N_7066);
or U8467 (N_8467,N_7055,N_7871);
nor U8468 (N_8468,N_7872,N_7735);
nand U8469 (N_8469,N_7319,N_7125);
nand U8470 (N_8470,N_7087,N_7827);
or U8471 (N_8471,N_7298,N_7481);
nand U8472 (N_8472,N_7405,N_7836);
and U8473 (N_8473,N_7993,N_7068);
or U8474 (N_8474,N_7263,N_7997);
and U8475 (N_8475,N_7753,N_7880);
and U8476 (N_8476,N_7457,N_7227);
nand U8477 (N_8477,N_7828,N_7030);
nor U8478 (N_8478,N_7408,N_7236);
nor U8479 (N_8479,N_7543,N_7781);
and U8480 (N_8480,N_7758,N_7374);
nand U8481 (N_8481,N_7743,N_7028);
nand U8482 (N_8482,N_7513,N_7283);
nand U8483 (N_8483,N_7857,N_7691);
or U8484 (N_8484,N_7362,N_7166);
and U8485 (N_8485,N_7486,N_7963);
and U8486 (N_8486,N_7673,N_7092);
nand U8487 (N_8487,N_7053,N_7182);
nand U8488 (N_8488,N_7257,N_7765);
or U8489 (N_8489,N_7715,N_7536);
nor U8490 (N_8490,N_7131,N_7522);
or U8491 (N_8491,N_7247,N_7794);
or U8492 (N_8492,N_7908,N_7387);
or U8493 (N_8493,N_7903,N_7505);
and U8494 (N_8494,N_7592,N_7778);
nor U8495 (N_8495,N_7314,N_7886);
nor U8496 (N_8496,N_7116,N_7617);
nor U8497 (N_8497,N_7566,N_7441);
nor U8498 (N_8498,N_7605,N_7279);
and U8499 (N_8499,N_7671,N_7034);
or U8500 (N_8500,N_7975,N_7268);
nor U8501 (N_8501,N_7993,N_7372);
nand U8502 (N_8502,N_7941,N_7104);
nand U8503 (N_8503,N_7111,N_7105);
nand U8504 (N_8504,N_7499,N_7794);
or U8505 (N_8505,N_7148,N_7389);
or U8506 (N_8506,N_7771,N_7492);
nor U8507 (N_8507,N_7876,N_7895);
nor U8508 (N_8508,N_7174,N_7706);
and U8509 (N_8509,N_7631,N_7104);
and U8510 (N_8510,N_7400,N_7193);
and U8511 (N_8511,N_7696,N_7310);
xor U8512 (N_8512,N_7830,N_7278);
nand U8513 (N_8513,N_7491,N_7034);
nand U8514 (N_8514,N_7586,N_7059);
and U8515 (N_8515,N_7973,N_7780);
or U8516 (N_8516,N_7748,N_7061);
or U8517 (N_8517,N_7148,N_7295);
or U8518 (N_8518,N_7665,N_7987);
nand U8519 (N_8519,N_7222,N_7403);
or U8520 (N_8520,N_7333,N_7552);
and U8521 (N_8521,N_7170,N_7319);
or U8522 (N_8522,N_7457,N_7635);
nand U8523 (N_8523,N_7570,N_7214);
and U8524 (N_8524,N_7244,N_7636);
nor U8525 (N_8525,N_7920,N_7985);
nor U8526 (N_8526,N_7898,N_7332);
nor U8527 (N_8527,N_7546,N_7796);
nand U8528 (N_8528,N_7602,N_7792);
nand U8529 (N_8529,N_7083,N_7063);
nor U8530 (N_8530,N_7278,N_7641);
and U8531 (N_8531,N_7021,N_7806);
nand U8532 (N_8532,N_7499,N_7123);
nand U8533 (N_8533,N_7323,N_7812);
nand U8534 (N_8534,N_7575,N_7761);
or U8535 (N_8535,N_7349,N_7532);
or U8536 (N_8536,N_7063,N_7633);
and U8537 (N_8537,N_7603,N_7128);
nand U8538 (N_8538,N_7000,N_7790);
and U8539 (N_8539,N_7462,N_7875);
nor U8540 (N_8540,N_7103,N_7447);
or U8541 (N_8541,N_7093,N_7089);
and U8542 (N_8542,N_7926,N_7883);
nand U8543 (N_8543,N_7785,N_7045);
and U8544 (N_8544,N_7626,N_7325);
nor U8545 (N_8545,N_7928,N_7604);
and U8546 (N_8546,N_7922,N_7279);
or U8547 (N_8547,N_7401,N_7842);
or U8548 (N_8548,N_7172,N_7764);
nor U8549 (N_8549,N_7044,N_7536);
and U8550 (N_8550,N_7697,N_7242);
nor U8551 (N_8551,N_7269,N_7149);
or U8552 (N_8552,N_7190,N_7506);
nand U8553 (N_8553,N_7977,N_7176);
nand U8554 (N_8554,N_7280,N_7395);
nand U8555 (N_8555,N_7833,N_7359);
nor U8556 (N_8556,N_7630,N_7345);
nor U8557 (N_8557,N_7523,N_7210);
nand U8558 (N_8558,N_7914,N_7360);
or U8559 (N_8559,N_7342,N_7633);
or U8560 (N_8560,N_7062,N_7881);
nor U8561 (N_8561,N_7411,N_7764);
or U8562 (N_8562,N_7317,N_7773);
nand U8563 (N_8563,N_7448,N_7346);
or U8564 (N_8564,N_7531,N_7755);
or U8565 (N_8565,N_7124,N_7597);
or U8566 (N_8566,N_7028,N_7795);
and U8567 (N_8567,N_7457,N_7601);
or U8568 (N_8568,N_7187,N_7884);
or U8569 (N_8569,N_7397,N_7562);
and U8570 (N_8570,N_7363,N_7483);
or U8571 (N_8571,N_7268,N_7863);
and U8572 (N_8572,N_7903,N_7481);
nand U8573 (N_8573,N_7461,N_7711);
or U8574 (N_8574,N_7967,N_7088);
nor U8575 (N_8575,N_7593,N_7455);
or U8576 (N_8576,N_7620,N_7305);
nor U8577 (N_8577,N_7594,N_7040);
nand U8578 (N_8578,N_7368,N_7977);
and U8579 (N_8579,N_7508,N_7722);
nor U8580 (N_8580,N_7125,N_7389);
and U8581 (N_8581,N_7852,N_7930);
nand U8582 (N_8582,N_7778,N_7089);
nand U8583 (N_8583,N_7687,N_7575);
nand U8584 (N_8584,N_7988,N_7050);
nor U8585 (N_8585,N_7482,N_7297);
nand U8586 (N_8586,N_7192,N_7448);
and U8587 (N_8587,N_7413,N_7822);
and U8588 (N_8588,N_7697,N_7568);
nand U8589 (N_8589,N_7032,N_7944);
xor U8590 (N_8590,N_7528,N_7374);
nor U8591 (N_8591,N_7123,N_7796);
or U8592 (N_8592,N_7001,N_7937);
nand U8593 (N_8593,N_7265,N_7784);
or U8594 (N_8594,N_7283,N_7347);
and U8595 (N_8595,N_7602,N_7228);
xor U8596 (N_8596,N_7667,N_7514);
nor U8597 (N_8597,N_7556,N_7153);
nor U8598 (N_8598,N_7861,N_7578);
nand U8599 (N_8599,N_7532,N_7992);
and U8600 (N_8600,N_7523,N_7864);
or U8601 (N_8601,N_7403,N_7843);
and U8602 (N_8602,N_7136,N_7022);
and U8603 (N_8603,N_7244,N_7284);
or U8604 (N_8604,N_7457,N_7031);
xor U8605 (N_8605,N_7838,N_7018);
and U8606 (N_8606,N_7848,N_7325);
nand U8607 (N_8607,N_7420,N_7814);
or U8608 (N_8608,N_7414,N_7498);
nand U8609 (N_8609,N_7606,N_7153);
or U8610 (N_8610,N_7449,N_7863);
nor U8611 (N_8611,N_7173,N_7599);
or U8612 (N_8612,N_7782,N_7526);
or U8613 (N_8613,N_7902,N_7236);
or U8614 (N_8614,N_7452,N_7817);
and U8615 (N_8615,N_7168,N_7098);
or U8616 (N_8616,N_7687,N_7418);
nor U8617 (N_8617,N_7315,N_7579);
and U8618 (N_8618,N_7483,N_7556);
nand U8619 (N_8619,N_7964,N_7966);
or U8620 (N_8620,N_7832,N_7940);
or U8621 (N_8621,N_7028,N_7345);
xor U8622 (N_8622,N_7183,N_7425);
and U8623 (N_8623,N_7518,N_7792);
or U8624 (N_8624,N_7233,N_7198);
and U8625 (N_8625,N_7195,N_7561);
and U8626 (N_8626,N_7775,N_7244);
or U8627 (N_8627,N_7156,N_7047);
nand U8628 (N_8628,N_7500,N_7662);
and U8629 (N_8629,N_7246,N_7637);
nor U8630 (N_8630,N_7008,N_7406);
or U8631 (N_8631,N_7458,N_7774);
or U8632 (N_8632,N_7553,N_7647);
and U8633 (N_8633,N_7834,N_7778);
and U8634 (N_8634,N_7575,N_7384);
nor U8635 (N_8635,N_7068,N_7923);
nor U8636 (N_8636,N_7902,N_7609);
or U8637 (N_8637,N_7836,N_7664);
nand U8638 (N_8638,N_7550,N_7773);
or U8639 (N_8639,N_7262,N_7111);
nand U8640 (N_8640,N_7282,N_7290);
nor U8641 (N_8641,N_7337,N_7490);
xor U8642 (N_8642,N_7849,N_7982);
xnor U8643 (N_8643,N_7642,N_7671);
nand U8644 (N_8644,N_7665,N_7675);
nand U8645 (N_8645,N_7804,N_7056);
and U8646 (N_8646,N_7448,N_7960);
nor U8647 (N_8647,N_7819,N_7141);
or U8648 (N_8648,N_7147,N_7104);
nand U8649 (N_8649,N_7683,N_7159);
nand U8650 (N_8650,N_7688,N_7436);
nand U8651 (N_8651,N_7551,N_7491);
nor U8652 (N_8652,N_7748,N_7614);
nand U8653 (N_8653,N_7574,N_7378);
and U8654 (N_8654,N_7349,N_7473);
or U8655 (N_8655,N_7170,N_7781);
and U8656 (N_8656,N_7112,N_7375);
nor U8657 (N_8657,N_7157,N_7892);
nor U8658 (N_8658,N_7577,N_7677);
nor U8659 (N_8659,N_7013,N_7377);
and U8660 (N_8660,N_7032,N_7416);
nand U8661 (N_8661,N_7390,N_7745);
and U8662 (N_8662,N_7085,N_7750);
nor U8663 (N_8663,N_7157,N_7797);
nand U8664 (N_8664,N_7737,N_7384);
nand U8665 (N_8665,N_7152,N_7064);
nand U8666 (N_8666,N_7191,N_7975);
nor U8667 (N_8667,N_7679,N_7009);
and U8668 (N_8668,N_7178,N_7642);
xnor U8669 (N_8669,N_7315,N_7016);
nor U8670 (N_8670,N_7291,N_7575);
nor U8671 (N_8671,N_7461,N_7707);
or U8672 (N_8672,N_7844,N_7786);
nand U8673 (N_8673,N_7660,N_7832);
nand U8674 (N_8674,N_7460,N_7851);
nor U8675 (N_8675,N_7408,N_7853);
nor U8676 (N_8676,N_7495,N_7497);
nand U8677 (N_8677,N_7425,N_7373);
nand U8678 (N_8678,N_7909,N_7023);
nor U8679 (N_8679,N_7264,N_7935);
nand U8680 (N_8680,N_7351,N_7334);
nor U8681 (N_8681,N_7534,N_7599);
and U8682 (N_8682,N_7983,N_7121);
nor U8683 (N_8683,N_7843,N_7899);
nand U8684 (N_8684,N_7398,N_7345);
and U8685 (N_8685,N_7599,N_7888);
nor U8686 (N_8686,N_7377,N_7762);
or U8687 (N_8687,N_7903,N_7081);
nand U8688 (N_8688,N_7116,N_7073);
nor U8689 (N_8689,N_7415,N_7124);
or U8690 (N_8690,N_7907,N_7741);
and U8691 (N_8691,N_7652,N_7906);
and U8692 (N_8692,N_7867,N_7761);
or U8693 (N_8693,N_7616,N_7219);
nand U8694 (N_8694,N_7646,N_7156);
nand U8695 (N_8695,N_7235,N_7017);
nand U8696 (N_8696,N_7300,N_7280);
and U8697 (N_8697,N_7067,N_7433);
nor U8698 (N_8698,N_7797,N_7119);
nand U8699 (N_8699,N_7036,N_7348);
nor U8700 (N_8700,N_7485,N_7294);
nor U8701 (N_8701,N_7270,N_7127);
and U8702 (N_8702,N_7241,N_7467);
nand U8703 (N_8703,N_7220,N_7956);
and U8704 (N_8704,N_7568,N_7430);
or U8705 (N_8705,N_7509,N_7999);
and U8706 (N_8706,N_7045,N_7490);
nor U8707 (N_8707,N_7938,N_7088);
and U8708 (N_8708,N_7458,N_7596);
nand U8709 (N_8709,N_7394,N_7140);
nor U8710 (N_8710,N_7229,N_7110);
nand U8711 (N_8711,N_7847,N_7241);
nand U8712 (N_8712,N_7109,N_7045);
or U8713 (N_8713,N_7023,N_7329);
and U8714 (N_8714,N_7139,N_7620);
nor U8715 (N_8715,N_7417,N_7264);
nand U8716 (N_8716,N_7575,N_7429);
or U8717 (N_8717,N_7104,N_7962);
or U8718 (N_8718,N_7317,N_7158);
nor U8719 (N_8719,N_7655,N_7972);
nand U8720 (N_8720,N_7923,N_7146);
or U8721 (N_8721,N_7384,N_7600);
and U8722 (N_8722,N_7289,N_7147);
and U8723 (N_8723,N_7786,N_7816);
nor U8724 (N_8724,N_7733,N_7472);
and U8725 (N_8725,N_7829,N_7860);
nor U8726 (N_8726,N_7163,N_7250);
xnor U8727 (N_8727,N_7015,N_7173);
nand U8728 (N_8728,N_7912,N_7611);
nand U8729 (N_8729,N_7973,N_7250);
nor U8730 (N_8730,N_7143,N_7784);
or U8731 (N_8731,N_7678,N_7484);
and U8732 (N_8732,N_7990,N_7525);
and U8733 (N_8733,N_7611,N_7711);
nor U8734 (N_8734,N_7396,N_7014);
nand U8735 (N_8735,N_7839,N_7215);
nor U8736 (N_8736,N_7755,N_7127);
nor U8737 (N_8737,N_7690,N_7775);
nand U8738 (N_8738,N_7535,N_7526);
nand U8739 (N_8739,N_7817,N_7923);
nor U8740 (N_8740,N_7442,N_7106);
nor U8741 (N_8741,N_7872,N_7264);
nand U8742 (N_8742,N_7571,N_7828);
and U8743 (N_8743,N_7271,N_7935);
and U8744 (N_8744,N_7357,N_7091);
and U8745 (N_8745,N_7023,N_7960);
and U8746 (N_8746,N_7856,N_7379);
nor U8747 (N_8747,N_7070,N_7818);
and U8748 (N_8748,N_7624,N_7433);
and U8749 (N_8749,N_7682,N_7078);
nand U8750 (N_8750,N_7316,N_7426);
or U8751 (N_8751,N_7139,N_7812);
or U8752 (N_8752,N_7952,N_7140);
nand U8753 (N_8753,N_7776,N_7925);
nor U8754 (N_8754,N_7220,N_7988);
or U8755 (N_8755,N_7140,N_7458);
or U8756 (N_8756,N_7871,N_7305);
nor U8757 (N_8757,N_7253,N_7777);
nand U8758 (N_8758,N_7113,N_7482);
nor U8759 (N_8759,N_7864,N_7767);
or U8760 (N_8760,N_7006,N_7870);
nand U8761 (N_8761,N_7886,N_7563);
and U8762 (N_8762,N_7987,N_7538);
nand U8763 (N_8763,N_7034,N_7499);
and U8764 (N_8764,N_7062,N_7662);
nand U8765 (N_8765,N_7947,N_7934);
and U8766 (N_8766,N_7643,N_7599);
or U8767 (N_8767,N_7021,N_7877);
or U8768 (N_8768,N_7245,N_7497);
or U8769 (N_8769,N_7746,N_7692);
nor U8770 (N_8770,N_7665,N_7509);
and U8771 (N_8771,N_7964,N_7553);
and U8772 (N_8772,N_7197,N_7171);
or U8773 (N_8773,N_7300,N_7887);
and U8774 (N_8774,N_7946,N_7210);
and U8775 (N_8775,N_7993,N_7199);
and U8776 (N_8776,N_7111,N_7769);
or U8777 (N_8777,N_7575,N_7295);
nor U8778 (N_8778,N_7679,N_7519);
nor U8779 (N_8779,N_7805,N_7968);
or U8780 (N_8780,N_7137,N_7440);
or U8781 (N_8781,N_7808,N_7674);
and U8782 (N_8782,N_7302,N_7160);
and U8783 (N_8783,N_7360,N_7274);
nor U8784 (N_8784,N_7480,N_7713);
nand U8785 (N_8785,N_7639,N_7781);
nor U8786 (N_8786,N_7058,N_7826);
or U8787 (N_8787,N_7798,N_7218);
nor U8788 (N_8788,N_7076,N_7264);
and U8789 (N_8789,N_7199,N_7242);
nor U8790 (N_8790,N_7687,N_7605);
nand U8791 (N_8791,N_7001,N_7192);
and U8792 (N_8792,N_7740,N_7699);
or U8793 (N_8793,N_7074,N_7187);
and U8794 (N_8794,N_7403,N_7692);
nor U8795 (N_8795,N_7182,N_7762);
or U8796 (N_8796,N_7731,N_7543);
nand U8797 (N_8797,N_7481,N_7755);
nor U8798 (N_8798,N_7407,N_7523);
or U8799 (N_8799,N_7429,N_7812);
and U8800 (N_8800,N_7197,N_7683);
nand U8801 (N_8801,N_7767,N_7271);
and U8802 (N_8802,N_7405,N_7859);
or U8803 (N_8803,N_7249,N_7337);
nor U8804 (N_8804,N_7846,N_7983);
nand U8805 (N_8805,N_7647,N_7873);
or U8806 (N_8806,N_7502,N_7167);
and U8807 (N_8807,N_7729,N_7037);
or U8808 (N_8808,N_7151,N_7928);
nor U8809 (N_8809,N_7492,N_7126);
and U8810 (N_8810,N_7176,N_7151);
nor U8811 (N_8811,N_7250,N_7858);
or U8812 (N_8812,N_7340,N_7934);
nand U8813 (N_8813,N_7921,N_7577);
nand U8814 (N_8814,N_7998,N_7837);
and U8815 (N_8815,N_7758,N_7394);
nor U8816 (N_8816,N_7181,N_7942);
nor U8817 (N_8817,N_7925,N_7007);
or U8818 (N_8818,N_7912,N_7937);
nand U8819 (N_8819,N_7371,N_7557);
or U8820 (N_8820,N_7486,N_7161);
and U8821 (N_8821,N_7649,N_7199);
nand U8822 (N_8822,N_7902,N_7827);
nor U8823 (N_8823,N_7155,N_7697);
nand U8824 (N_8824,N_7273,N_7344);
and U8825 (N_8825,N_7921,N_7257);
and U8826 (N_8826,N_7861,N_7015);
and U8827 (N_8827,N_7668,N_7404);
or U8828 (N_8828,N_7518,N_7089);
and U8829 (N_8829,N_7134,N_7785);
nor U8830 (N_8830,N_7444,N_7635);
nor U8831 (N_8831,N_7849,N_7306);
nor U8832 (N_8832,N_7089,N_7084);
nor U8833 (N_8833,N_7368,N_7481);
or U8834 (N_8834,N_7999,N_7062);
or U8835 (N_8835,N_7761,N_7456);
and U8836 (N_8836,N_7749,N_7564);
nor U8837 (N_8837,N_7794,N_7709);
and U8838 (N_8838,N_7230,N_7330);
nand U8839 (N_8839,N_7199,N_7786);
nand U8840 (N_8840,N_7725,N_7870);
nand U8841 (N_8841,N_7112,N_7874);
nand U8842 (N_8842,N_7821,N_7366);
nor U8843 (N_8843,N_7896,N_7395);
nand U8844 (N_8844,N_7402,N_7093);
nand U8845 (N_8845,N_7906,N_7450);
nand U8846 (N_8846,N_7384,N_7558);
nor U8847 (N_8847,N_7896,N_7636);
nor U8848 (N_8848,N_7606,N_7475);
nor U8849 (N_8849,N_7823,N_7495);
or U8850 (N_8850,N_7149,N_7265);
xor U8851 (N_8851,N_7832,N_7879);
nor U8852 (N_8852,N_7563,N_7392);
or U8853 (N_8853,N_7702,N_7371);
and U8854 (N_8854,N_7769,N_7642);
and U8855 (N_8855,N_7333,N_7421);
or U8856 (N_8856,N_7307,N_7342);
nor U8857 (N_8857,N_7133,N_7041);
or U8858 (N_8858,N_7051,N_7693);
and U8859 (N_8859,N_7713,N_7025);
or U8860 (N_8860,N_7018,N_7418);
or U8861 (N_8861,N_7333,N_7941);
or U8862 (N_8862,N_7989,N_7711);
nor U8863 (N_8863,N_7041,N_7859);
nor U8864 (N_8864,N_7687,N_7401);
and U8865 (N_8865,N_7306,N_7265);
nor U8866 (N_8866,N_7397,N_7101);
nand U8867 (N_8867,N_7151,N_7744);
xor U8868 (N_8868,N_7590,N_7661);
nand U8869 (N_8869,N_7817,N_7744);
nor U8870 (N_8870,N_7642,N_7683);
and U8871 (N_8871,N_7223,N_7830);
nand U8872 (N_8872,N_7788,N_7484);
nor U8873 (N_8873,N_7207,N_7609);
or U8874 (N_8874,N_7313,N_7368);
and U8875 (N_8875,N_7173,N_7087);
or U8876 (N_8876,N_7258,N_7932);
or U8877 (N_8877,N_7524,N_7239);
or U8878 (N_8878,N_7674,N_7732);
and U8879 (N_8879,N_7703,N_7634);
nand U8880 (N_8880,N_7922,N_7372);
and U8881 (N_8881,N_7185,N_7230);
and U8882 (N_8882,N_7495,N_7463);
nor U8883 (N_8883,N_7628,N_7511);
and U8884 (N_8884,N_7184,N_7999);
or U8885 (N_8885,N_7900,N_7360);
nand U8886 (N_8886,N_7935,N_7064);
nand U8887 (N_8887,N_7744,N_7769);
and U8888 (N_8888,N_7639,N_7317);
or U8889 (N_8889,N_7095,N_7467);
nand U8890 (N_8890,N_7897,N_7444);
or U8891 (N_8891,N_7652,N_7804);
nor U8892 (N_8892,N_7401,N_7205);
nor U8893 (N_8893,N_7724,N_7768);
and U8894 (N_8894,N_7435,N_7121);
and U8895 (N_8895,N_7534,N_7450);
nor U8896 (N_8896,N_7439,N_7552);
and U8897 (N_8897,N_7840,N_7043);
nand U8898 (N_8898,N_7957,N_7835);
nand U8899 (N_8899,N_7484,N_7284);
and U8900 (N_8900,N_7961,N_7442);
nand U8901 (N_8901,N_7073,N_7311);
or U8902 (N_8902,N_7036,N_7554);
and U8903 (N_8903,N_7102,N_7210);
xor U8904 (N_8904,N_7507,N_7766);
or U8905 (N_8905,N_7465,N_7890);
or U8906 (N_8906,N_7568,N_7288);
and U8907 (N_8907,N_7528,N_7016);
nand U8908 (N_8908,N_7223,N_7915);
or U8909 (N_8909,N_7902,N_7197);
nor U8910 (N_8910,N_7982,N_7140);
nor U8911 (N_8911,N_7555,N_7013);
or U8912 (N_8912,N_7758,N_7400);
nor U8913 (N_8913,N_7979,N_7391);
nor U8914 (N_8914,N_7902,N_7237);
nor U8915 (N_8915,N_7181,N_7017);
or U8916 (N_8916,N_7885,N_7005);
nor U8917 (N_8917,N_7534,N_7614);
nor U8918 (N_8918,N_7448,N_7587);
or U8919 (N_8919,N_7457,N_7867);
nand U8920 (N_8920,N_7852,N_7194);
and U8921 (N_8921,N_7058,N_7274);
nand U8922 (N_8922,N_7207,N_7291);
nand U8923 (N_8923,N_7802,N_7109);
nand U8924 (N_8924,N_7170,N_7562);
or U8925 (N_8925,N_7852,N_7305);
nand U8926 (N_8926,N_7523,N_7277);
nor U8927 (N_8927,N_7967,N_7139);
nor U8928 (N_8928,N_7633,N_7548);
nand U8929 (N_8929,N_7836,N_7350);
and U8930 (N_8930,N_7868,N_7808);
nand U8931 (N_8931,N_7638,N_7289);
nor U8932 (N_8932,N_7932,N_7526);
nand U8933 (N_8933,N_7778,N_7212);
nand U8934 (N_8934,N_7744,N_7746);
xor U8935 (N_8935,N_7461,N_7339);
and U8936 (N_8936,N_7744,N_7594);
nand U8937 (N_8937,N_7018,N_7934);
or U8938 (N_8938,N_7839,N_7461);
and U8939 (N_8939,N_7020,N_7323);
or U8940 (N_8940,N_7204,N_7289);
nand U8941 (N_8941,N_7712,N_7119);
nand U8942 (N_8942,N_7495,N_7199);
or U8943 (N_8943,N_7743,N_7199);
nand U8944 (N_8944,N_7720,N_7100);
and U8945 (N_8945,N_7377,N_7998);
nor U8946 (N_8946,N_7412,N_7938);
nor U8947 (N_8947,N_7044,N_7132);
or U8948 (N_8948,N_7282,N_7845);
and U8949 (N_8949,N_7087,N_7415);
and U8950 (N_8950,N_7416,N_7578);
and U8951 (N_8951,N_7587,N_7202);
and U8952 (N_8952,N_7644,N_7671);
or U8953 (N_8953,N_7922,N_7109);
or U8954 (N_8954,N_7757,N_7089);
or U8955 (N_8955,N_7054,N_7967);
nor U8956 (N_8956,N_7200,N_7008);
and U8957 (N_8957,N_7448,N_7614);
or U8958 (N_8958,N_7501,N_7393);
xor U8959 (N_8959,N_7912,N_7957);
nand U8960 (N_8960,N_7901,N_7948);
or U8961 (N_8961,N_7680,N_7226);
nand U8962 (N_8962,N_7249,N_7422);
nand U8963 (N_8963,N_7363,N_7752);
or U8964 (N_8964,N_7609,N_7055);
nor U8965 (N_8965,N_7696,N_7346);
and U8966 (N_8966,N_7310,N_7763);
and U8967 (N_8967,N_7411,N_7954);
nor U8968 (N_8968,N_7703,N_7317);
nor U8969 (N_8969,N_7560,N_7649);
nor U8970 (N_8970,N_7575,N_7351);
and U8971 (N_8971,N_7561,N_7221);
or U8972 (N_8972,N_7463,N_7377);
and U8973 (N_8973,N_7373,N_7634);
and U8974 (N_8974,N_7557,N_7226);
nor U8975 (N_8975,N_7995,N_7975);
or U8976 (N_8976,N_7914,N_7293);
or U8977 (N_8977,N_7113,N_7239);
nand U8978 (N_8978,N_7001,N_7214);
and U8979 (N_8979,N_7846,N_7043);
or U8980 (N_8980,N_7432,N_7930);
nor U8981 (N_8981,N_7098,N_7288);
or U8982 (N_8982,N_7194,N_7101);
or U8983 (N_8983,N_7984,N_7503);
nor U8984 (N_8984,N_7827,N_7882);
nand U8985 (N_8985,N_7302,N_7262);
nor U8986 (N_8986,N_7770,N_7627);
or U8987 (N_8987,N_7131,N_7920);
or U8988 (N_8988,N_7176,N_7089);
and U8989 (N_8989,N_7189,N_7828);
and U8990 (N_8990,N_7634,N_7444);
nor U8991 (N_8991,N_7506,N_7842);
nor U8992 (N_8992,N_7863,N_7365);
and U8993 (N_8993,N_7786,N_7572);
nor U8994 (N_8994,N_7366,N_7925);
and U8995 (N_8995,N_7654,N_7980);
or U8996 (N_8996,N_7894,N_7197);
nor U8997 (N_8997,N_7661,N_7368);
nor U8998 (N_8998,N_7588,N_7533);
nand U8999 (N_8999,N_7609,N_7475);
or U9000 (N_9000,N_8361,N_8693);
nand U9001 (N_9001,N_8212,N_8183);
nand U9002 (N_9002,N_8963,N_8200);
and U9003 (N_9003,N_8955,N_8265);
nand U9004 (N_9004,N_8038,N_8329);
or U9005 (N_9005,N_8862,N_8843);
nor U9006 (N_9006,N_8421,N_8445);
and U9007 (N_9007,N_8077,N_8951);
nand U9008 (N_9008,N_8671,N_8112);
or U9009 (N_9009,N_8612,N_8160);
nor U9010 (N_9010,N_8854,N_8100);
nor U9011 (N_9011,N_8455,N_8980);
or U9012 (N_9012,N_8834,N_8477);
nand U9013 (N_9013,N_8378,N_8125);
nor U9014 (N_9014,N_8318,N_8132);
and U9015 (N_9015,N_8607,N_8549);
and U9016 (N_9016,N_8859,N_8882);
nand U9017 (N_9017,N_8878,N_8135);
and U9018 (N_9018,N_8430,N_8780);
nand U9019 (N_9019,N_8102,N_8247);
nor U9020 (N_9020,N_8703,N_8094);
and U9021 (N_9021,N_8023,N_8979);
xnor U9022 (N_9022,N_8062,N_8435);
nor U9023 (N_9023,N_8239,N_8537);
nand U9024 (N_9024,N_8260,N_8974);
or U9025 (N_9025,N_8128,N_8567);
and U9026 (N_9026,N_8064,N_8746);
or U9027 (N_9027,N_8691,N_8641);
nand U9028 (N_9028,N_8017,N_8916);
or U9029 (N_9029,N_8405,N_8444);
nand U9030 (N_9030,N_8093,N_8424);
and U9031 (N_9031,N_8811,N_8787);
or U9032 (N_9032,N_8154,N_8035);
nor U9033 (N_9033,N_8398,N_8485);
nor U9034 (N_9034,N_8753,N_8978);
nor U9035 (N_9035,N_8923,N_8973);
nand U9036 (N_9036,N_8769,N_8947);
and U9037 (N_9037,N_8294,N_8263);
nor U9038 (N_9038,N_8552,N_8512);
nor U9039 (N_9039,N_8039,N_8891);
nor U9040 (N_9040,N_8423,N_8653);
or U9041 (N_9041,N_8729,N_8770);
and U9042 (N_9042,N_8084,N_8598);
or U9043 (N_9043,N_8596,N_8850);
or U9044 (N_9044,N_8801,N_8220);
and U9045 (N_9045,N_8748,N_8033);
and U9046 (N_9046,N_8067,N_8205);
nand U9047 (N_9047,N_8032,N_8600);
nand U9048 (N_9048,N_8027,N_8502);
nand U9049 (N_9049,N_8681,N_8798);
nand U9050 (N_9050,N_8751,N_8050);
nand U9051 (N_9051,N_8351,N_8897);
nand U9052 (N_9052,N_8156,N_8687);
nand U9053 (N_9053,N_8442,N_8108);
or U9054 (N_9054,N_8011,N_8130);
nand U9055 (N_9055,N_8817,N_8254);
nand U9056 (N_9056,N_8383,N_8752);
and U9057 (N_9057,N_8574,N_8180);
and U9058 (N_9058,N_8971,N_8233);
and U9059 (N_9059,N_8056,N_8773);
nor U9060 (N_9060,N_8949,N_8583);
nand U9061 (N_9061,N_8426,N_8219);
nand U9062 (N_9062,N_8203,N_8126);
or U9063 (N_9063,N_8232,N_8704);
or U9064 (N_9064,N_8007,N_8099);
nor U9065 (N_9065,N_8343,N_8287);
nand U9066 (N_9066,N_8396,N_8005);
and U9067 (N_9067,N_8051,N_8117);
nor U9068 (N_9068,N_8909,N_8791);
and U9069 (N_9069,N_8730,N_8532);
xnor U9070 (N_9070,N_8465,N_8985);
and U9071 (N_9071,N_8387,N_8282);
nor U9072 (N_9072,N_8766,N_8347);
and U9073 (N_9073,N_8984,N_8210);
nor U9074 (N_9074,N_8519,N_8257);
or U9075 (N_9075,N_8085,N_8724);
or U9076 (N_9076,N_8790,N_8461);
or U9077 (N_9077,N_8413,N_8699);
or U9078 (N_9078,N_8688,N_8599);
nor U9079 (N_9079,N_8079,N_8745);
nor U9080 (N_9080,N_8358,N_8676);
nor U9081 (N_9081,N_8755,N_8242);
and U9082 (N_9082,N_8914,N_8166);
nand U9083 (N_9083,N_8410,N_8487);
nand U9084 (N_9084,N_8986,N_8606);
nand U9085 (N_9085,N_8412,N_8307);
nand U9086 (N_9086,N_8074,N_8917);
or U9087 (N_9087,N_8721,N_8518);
nand U9088 (N_9088,N_8553,N_8957);
nor U9089 (N_9089,N_8371,N_8913);
or U9090 (N_9090,N_8002,N_8509);
nand U9091 (N_9091,N_8040,N_8860);
and U9092 (N_9092,N_8925,N_8828);
or U9093 (N_9093,N_8514,N_8972);
and U9094 (N_9094,N_8268,N_8261);
nand U9095 (N_9095,N_8929,N_8990);
nor U9096 (N_9096,N_8411,N_8912);
nand U9097 (N_9097,N_8150,N_8161);
nand U9098 (N_9098,N_8975,N_8441);
nand U9099 (N_9099,N_8624,N_8357);
or U9100 (N_9100,N_8407,N_8109);
nand U9101 (N_9101,N_8735,N_8149);
nor U9102 (N_9102,N_8024,N_8018);
or U9103 (N_9103,N_8105,N_8072);
or U9104 (N_9104,N_8523,N_8215);
nand U9105 (N_9105,N_8824,N_8554);
or U9106 (N_9106,N_8896,N_8291);
nor U9107 (N_9107,N_8083,N_8044);
and U9108 (N_9108,N_8422,N_8118);
nand U9109 (N_9109,N_8527,N_8308);
and U9110 (N_9110,N_8388,N_8618);
and U9111 (N_9111,N_8177,N_8175);
nor U9112 (N_9112,N_8259,N_8964);
and U9113 (N_9113,N_8764,N_8999);
or U9114 (N_9114,N_8684,N_8223);
nand U9115 (N_9115,N_8280,N_8097);
nor U9116 (N_9116,N_8370,N_8677);
or U9117 (N_9117,N_8883,N_8073);
nand U9118 (N_9118,N_8070,N_8391);
and U9119 (N_9119,N_8562,N_8868);
or U9120 (N_9120,N_8772,N_8182);
or U9121 (N_9121,N_8471,N_8489);
nand U9122 (N_9122,N_8176,N_8089);
nand U9123 (N_9123,N_8341,N_8826);
nor U9124 (N_9124,N_8248,N_8524);
nor U9125 (N_9125,N_8959,N_8285);
and U9126 (N_9126,N_8473,N_8620);
nand U9127 (N_9127,N_8447,N_8103);
nand U9128 (N_9128,N_8921,N_8068);
nor U9129 (N_9129,N_8706,N_8800);
nand U9130 (N_9130,N_8590,N_8927);
nor U9131 (N_9131,N_8662,N_8720);
nor U9132 (N_9132,N_8181,N_8482);
or U9133 (N_9133,N_8750,N_8838);
nand U9134 (N_9134,N_8216,N_8918);
nand U9135 (N_9135,N_8875,N_8145);
and U9136 (N_9136,N_8174,N_8915);
nor U9137 (N_9137,N_8939,N_8713);
nor U9138 (N_9138,N_8825,N_8781);
nand U9139 (N_9139,N_8414,N_8353);
and U9140 (N_9140,N_8538,N_8907);
and U9141 (N_9141,N_8940,N_8840);
nor U9142 (N_9142,N_8472,N_8744);
nand U9143 (N_9143,N_8484,N_8934);
and U9144 (N_9144,N_8515,N_8983);
or U9145 (N_9145,N_8467,N_8195);
xor U9146 (N_9146,N_8119,N_8451);
and U9147 (N_9147,N_8267,N_8289);
nor U9148 (N_9148,N_8134,N_8303);
and U9149 (N_9149,N_8400,N_8041);
nor U9150 (N_9150,N_8253,N_8580);
or U9151 (N_9151,N_8202,N_8258);
or U9152 (N_9152,N_8301,N_8503);
and U9153 (N_9153,N_8924,N_8363);
and U9154 (N_9154,N_8295,N_8144);
or U9155 (N_9155,N_8292,N_8352);
and U9156 (N_9156,N_8158,N_8698);
nand U9157 (N_9157,N_8799,N_8696);
nand U9158 (N_9158,N_8306,N_8941);
nand U9159 (N_9159,N_8380,N_8082);
and U9160 (N_9160,N_8001,N_8320);
nand U9161 (N_9161,N_8014,N_8667);
nand U9162 (N_9162,N_8457,N_8640);
and U9163 (N_9163,N_8271,N_8053);
nand U9164 (N_9164,N_8446,N_8486);
or U9165 (N_9165,N_8066,N_8340);
or U9166 (N_9166,N_8777,N_8705);
or U9167 (N_9167,N_8581,N_8737);
nor U9168 (N_9168,N_8059,N_8701);
and U9169 (N_9169,N_8855,N_8443);
nand U9170 (N_9170,N_8235,N_8498);
or U9171 (N_9171,N_8305,N_8827);
nor U9172 (N_9172,N_8956,N_8806);
nand U9173 (N_9173,N_8020,N_8015);
or U9174 (N_9174,N_8533,N_8496);
xor U9175 (N_9175,N_8297,N_8165);
and U9176 (N_9176,N_8847,N_8114);
or U9177 (N_9177,N_8448,N_8500);
nor U9178 (N_9178,N_8262,N_8988);
nor U9179 (N_9179,N_8252,N_8829);
and U9180 (N_9180,N_8804,N_8315);
nand U9181 (N_9181,N_8873,N_8568);
or U9182 (N_9182,N_8675,N_8660);
or U9183 (N_9183,N_8768,N_8614);
and U9184 (N_9184,N_8609,N_8708);
or U9185 (N_9185,N_8645,N_8839);
nand U9186 (N_9186,N_8251,N_8522);
or U9187 (N_9187,N_8743,N_8456);
and U9188 (N_9188,N_8364,N_8594);
nor U9189 (N_9189,N_8762,N_8707);
or U9190 (N_9190,N_8098,N_8867);
nor U9191 (N_9191,N_8450,N_8588);
or U9192 (N_9192,N_8187,N_8967);
or U9193 (N_9193,N_8171,N_8576);
nor U9194 (N_9194,N_8314,N_8028);
and U9195 (N_9195,N_8016,N_8564);
nand U9196 (N_9196,N_8841,N_8739);
or U9197 (N_9197,N_8207,N_8619);
nor U9198 (N_9198,N_8731,N_8592);
or U9199 (N_9199,N_8244,N_8278);
or U9200 (N_9200,N_8617,N_8666);
nand U9201 (N_9201,N_8816,N_8481);
nor U9202 (N_9202,N_8655,N_8323);
or U9203 (N_9203,N_8173,N_8765);
or U9204 (N_9204,N_8194,N_8362);
nor U9205 (N_9205,N_8870,N_8530);
nand U9206 (N_9206,N_8389,N_8946);
nand U9207 (N_9207,N_8140,N_8866);
nand U9208 (N_9208,N_8452,N_8511);
nand U9209 (N_9209,N_8399,N_8876);
nor U9210 (N_9210,N_8814,N_8887);
nand U9211 (N_9211,N_8479,N_8366);
nor U9212 (N_9212,N_8243,N_8228);
xnor U9213 (N_9213,N_8899,N_8992);
nor U9214 (N_9214,N_8901,N_8734);
or U9215 (N_9215,N_8784,N_8404);
nor U9216 (N_9216,N_8528,N_8922);
or U9217 (N_9217,N_8153,N_8495);
nand U9218 (N_9218,N_8275,N_8968);
and U9219 (N_9219,N_8309,N_8075);
or U9220 (N_9220,N_8556,N_8204);
nand U9221 (N_9221,N_8492,N_8344);
or U9222 (N_9222,N_8848,N_8629);
xnor U9223 (N_9223,N_8723,N_8636);
nand U9224 (N_9224,N_8147,N_8139);
and U9225 (N_9225,N_8385,N_8402);
or U9226 (N_9226,N_8793,N_8571);
nand U9227 (N_9227,N_8668,N_8143);
or U9228 (N_9228,N_8052,N_8449);
or U9229 (N_9229,N_8326,N_8652);
or U9230 (N_9230,N_8884,N_8335);
and U9231 (N_9231,N_8010,N_8953);
or U9232 (N_9232,N_8822,N_8464);
or U9233 (N_9233,N_8965,N_8328);
and U9234 (N_9234,N_8439,N_8905);
nor U9235 (N_9235,N_8756,N_8792);
or U9236 (N_9236,N_8879,N_8272);
or U9237 (N_9237,N_8663,N_8234);
nor U9238 (N_9238,N_8715,N_8778);
or U9239 (N_9239,N_8551,N_8438);
nand U9240 (N_9240,N_8425,N_8384);
or U9241 (N_9241,N_8279,N_8845);
xor U9242 (N_9242,N_8240,N_8071);
or U9243 (N_9243,N_8127,N_8613);
and U9244 (N_9244,N_8036,N_8683);
nor U9245 (N_9245,N_8397,N_8236);
or U9246 (N_9246,N_8460,N_8987);
nor U9247 (N_9247,N_8131,N_8615);
nand U9248 (N_9248,N_8191,N_8348);
and U9249 (N_9249,N_8851,N_8419);
nor U9250 (N_9250,N_8037,N_8577);
and U9251 (N_9251,N_8434,N_8994);
nand U9252 (N_9252,N_8386,N_8602);
nor U9253 (N_9253,N_8138,N_8319);
nor U9254 (N_9254,N_8547,N_8776);
or U9255 (N_9255,N_8003,N_8217);
nand U9256 (N_9256,N_8749,N_8433);
or U9257 (N_9257,N_8179,N_8497);
nor U9258 (N_9258,N_8904,N_8616);
nand U9259 (N_9259,N_8658,N_8163);
or U9260 (N_9260,N_8944,N_8926);
nand U9261 (N_9261,N_8989,N_8758);
nand U9262 (N_9262,N_8494,N_8585);
nor U9263 (N_9263,N_8360,N_8042);
and U9264 (N_9264,N_8857,N_8638);
and U9265 (N_9265,N_8337,N_8717);
or U9266 (N_9266,N_8898,N_8277);
nand U9267 (N_9267,N_8648,N_8369);
and U9268 (N_9268,N_8356,N_8892);
or U9269 (N_9269,N_8058,N_8453);
nand U9270 (N_9270,N_8719,N_8065);
nand U9271 (N_9271,N_8540,N_8375);
nand U9272 (N_9272,N_8213,N_8754);
or U9273 (N_9273,N_8672,N_8920);
nor U9274 (N_9274,N_8808,N_8632);
nor U9275 (N_9275,N_8786,N_8164);
nand U9276 (N_9276,N_8863,N_8483);
nor U9277 (N_9277,N_8334,N_8785);
nand U9278 (N_9278,N_8810,N_8998);
xnor U9279 (N_9279,N_8539,N_8209);
nor U9280 (N_9280,N_8043,N_8325);
or U9281 (N_9281,N_8470,N_8642);
nand U9282 (N_9282,N_8432,N_8256);
or U9283 (N_9283,N_8055,N_8728);
nor U9284 (N_9284,N_8763,N_8718);
and U9285 (N_9285,N_8649,N_8888);
nand U9286 (N_9286,N_8797,N_8076);
or U9287 (N_9287,N_8637,N_8120);
nand U9288 (N_9288,N_8630,N_8555);
nand U9289 (N_9289,N_8890,N_8508);
nor U9290 (N_9290,N_8833,N_8692);
or U9291 (N_9291,N_8300,N_8650);
nand U9292 (N_9292,N_8429,N_8611);
nor U9293 (N_9293,N_8237,N_8224);
or U9294 (N_9294,N_8513,N_8406);
nor U9295 (N_9295,N_8837,N_8889);
or U9296 (N_9296,N_8088,N_8214);
nand U9297 (N_9297,N_8767,N_8725);
nor U9298 (N_9298,N_8570,N_8111);
or U9299 (N_9299,N_8674,N_8783);
nor U9300 (N_9300,N_8415,N_8871);
nor U9301 (N_9301,N_8293,N_8299);
or U9302 (N_9302,N_8317,N_8678);
and U9303 (N_9303,N_8115,N_8201);
nor U9304 (N_9304,N_8966,N_8910);
nand U9305 (N_9305,N_8991,N_8557);
xor U9306 (N_9306,N_8019,N_8381);
nor U9307 (N_9307,N_8633,N_8022);
or U9308 (N_9308,N_8331,N_8338);
or U9309 (N_9309,N_8782,N_8283);
nor U9310 (N_9310,N_8499,N_8760);
or U9311 (N_9311,N_8893,N_8818);
nor U9312 (N_9312,N_8646,N_8881);
nor U9313 (N_9313,N_8846,N_8566);
or U9314 (N_9314,N_8129,N_8431);
nor U9315 (N_9315,N_8367,N_8643);
nor U9316 (N_9316,N_8995,N_8961);
or U9317 (N_9317,N_8026,N_8006);
xor U9318 (N_9318,N_8936,N_8534);
and U9319 (N_9319,N_8029,N_8218);
and U9320 (N_9320,N_8025,N_8463);
or U9321 (N_9321,N_8342,N_8427);
nand U9322 (N_9322,N_8635,N_8273);
and U9323 (N_9323,N_8198,N_8517);
nor U9324 (N_9324,N_8116,N_8475);
and U9325 (N_9325,N_8466,N_8304);
and U9326 (N_9326,N_8206,N_8536);
nor U9327 (N_9327,N_8241,N_8507);
nor U9328 (N_9328,N_8151,N_8601);
nand U9329 (N_9329,N_8401,N_8542);
nor U9330 (N_9330,N_8759,N_8774);
and U9331 (N_9331,N_8063,N_8480);
nor U9332 (N_9332,N_8008,N_8656);
or U9333 (N_9333,N_8504,N_8659);
nand U9334 (N_9334,N_8416,N_8133);
or U9335 (N_9335,N_8332,N_8565);
or U9336 (N_9336,N_8142,N_8900);
nor U9337 (N_9337,N_8476,N_8208);
nor U9338 (N_9338,N_8771,N_8264);
or U9339 (N_9339,N_8152,N_8679);
nor U9340 (N_9340,N_8420,N_8757);
and U9341 (N_9341,N_8060,N_8061);
nand U9342 (N_9342,N_8324,N_8685);
nand U9343 (N_9343,N_8869,N_8993);
nor U9344 (N_9344,N_8096,N_8950);
or U9345 (N_9345,N_8908,N_8844);
nor U9346 (N_9346,N_8121,N_8546);
nand U9347 (N_9347,N_8584,N_8167);
and U9348 (N_9348,N_8170,N_8579);
or U9349 (N_9349,N_8394,N_8665);
or U9350 (N_9350,N_8977,N_8162);
and U9351 (N_9351,N_8661,N_8911);
or U9352 (N_9352,N_8626,N_8178);
and U9353 (N_9353,N_8428,N_8960);
and U9354 (N_9354,N_8409,N_8976);
nand U9355 (N_9355,N_8852,N_8761);
and U9356 (N_9356,N_8226,N_8591);
nor U9357 (N_9357,N_8469,N_8740);
nor U9358 (N_9358,N_8702,N_8057);
or U9359 (N_9359,N_8933,N_8490);
nand U9360 (N_9360,N_8312,N_8722);
nand U9361 (N_9361,N_8274,N_8578);
and U9362 (N_9362,N_8742,N_8830);
nor U9363 (N_9363,N_8516,N_8726);
or U9364 (N_9364,N_8081,N_8885);
and U9365 (N_9365,N_8937,N_8794);
nand U9366 (N_9366,N_8104,N_8589);
nand U9367 (N_9367,N_8316,N_8390);
and U9368 (N_9368,N_8789,N_8543);
nand U9369 (N_9369,N_8186,N_8238);
nor U9370 (N_9370,N_8747,N_8669);
nor U9371 (N_9371,N_8809,N_8945);
nor U9372 (N_9372,N_8012,N_8709);
nand U9373 (N_9373,N_8004,N_8664);
nand U9374 (N_9374,N_8298,N_8346);
nor U9375 (N_9375,N_8608,N_8694);
nor U9376 (N_9376,N_8284,N_8733);
nor U9377 (N_9377,N_8932,N_8417);
and U9378 (N_9378,N_8820,N_8379);
and U9379 (N_9379,N_8221,N_8313);
nor U9380 (N_9380,N_8886,N_8045);
nor U9381 (N_9381,N_8193,N_8478);
and U9382 (N_9382,N_8711,N_8788);
or U9383 (N_9383,N_8246,N_8894);
and U9384 (N_9384,N_8159,N_8835);
nor U9385 (N_9385,N_8573,N_8561);
nand U9386 (N_9386,N_8831,N_8943);
nor U9387 (N_9387,N_8586,N_8288);
and U9388 (N_9388,N_8141,N_8531);
or U9389 (N_9389,N_8996,N_8714);
and U9390 (N_9390,N_8560,N_8491);
and U9391 (N_9391,N_8529,N_8327);
and U9392 (N_9392,N_8582,N_8505);
nand U9393 (N_9393,N_8069,N_8009);
or U9394 (N_9394,N_8350,N_8697);
or U9395 (N_9395,N_8545,N_8468);
and U9396 (N_9396,N_8550,N_8958);
xor U9397 (N_9397,N_8610,N_8970);
and U9398 (N_9398,N_8354,N_8938);
or U9399 (N_9399,N_8710,N_8031);
nand U9400 (N_9400,N_8330,N_8110);
nand U9401 (N_9401,N_8651,N_8673);
nand U9402 (N_9402,N_8627,N_8872);
nor U9403 (N_9403,N_8842,N_8796);
and U9404 (N_9404,N_8336,N_8510);
or U9405 (N_9405,N_8321,N_8000);
and U9406 (N_9406,N_8593,N_8137);
or U9407 (N_9407,N_8628,N_8322);
nor U9408 (N_9408,N_8107,N_8680);
and U9409 (N_9409,N_8188,N_8185);
and U9410 (N_9410,N_8168,N_8225);
and U9411 (N_9411,N_8270,N_8374);
or U9412 (N_9412,N_8541,N_8245);
nand U9413 (N_9413,N_8928,N_8559);
or U9414 (N_9414,N_8086,N_8962);
or U9415 (N_9415,N_8231,N_8189);
or U9416 (N_9416,N_8080,N_8836);
nor U9417 (N_9417,N_8030,N_8563);
nand U9418 (N_9418,N_8865,N_8544);
and U9419 (N_9419,N_8392,N_8458);
nand U9420 (N_9420,N_8506,N_8395);
nand U9421 (N_9421,N_8190,N_8526);
and U9422 (N_9422,N_8521,N_8136);
nand U9423 (N_9423,N_8372,N_8603);
or U9424 (N_9424,N_8034,N_8874);
nor U9425 (N_9425,N_8172,N_8969);
and U9426 (N_9426,N_8997,N_8169);
and U9427 (N_9427,N_8013,N_8276);
nand U9428 (N_9428,N_8222,N_8775);
nor U9429 (N_9429,N_8339,N_8644);
nand U9430 (N_9430,N_8861,N_8981);
nor U9431 (N_9431,N_8700,N_8712);
and U9432 (N_9432,N_8249,N_8858);
nand U9433 (N_9433,N_8227,N_8310);
or U9434 (N_9434,N_8106,N_8548);
and U9435 (N_9435,N_8113,N_8622);
and U9436 (N_9436,N_8437,N_8286);
nor U9437 (N_9437,N_8365,N_8813);
and U9438 (N_9438,N_8634,N_8695);
nor U9439 (N_9439,N_8047,N_8631);
and U9440 (N_9440,N_8440,N_8501);
nand U9441 (N_9441,N_8952,N_8682);
or U9442 (N_9442,N_8906,N_8230);
and U9443 (N_9443,N_8572,N_8902);
nand U9444 (N_9444,N_8716,N_8123);
nand U9445 (N_9445,N_8393,N_8459);
or U9446 (N_9446,N_8856,N_8368);
and U9447 (N_9447,N_8821,N_8654);
nor U9448 (N_9448,N_8078,N_8657);
nand U9449 (N_9449,N_8625,N_8832);
nand U9450 (N_9450,N_8605,N_8359);
or U9451 (N_9451,N_8408,N_8345);
nand U9452 (N_9452,N_8930,N_8122);
or U9453 (N_9453,N_8880,N_8290);
or U9454 (N_9454,N_8803,N_8101);
nand U9455 (N_9455,N_8157,N_8349);
and U9456 (N_9456,N_8942,N_8812);
or U9457 (N_9457,N_8054,N_8255);
nor U9458 (N_9458,N_8670,N_8587);
or U9459 (N_9459,N_8823,N_8647);
xor U9460 (N_9460,N_8621,N_8802);
nand U9461 (N_9461,N_8376,N_8815);
nand U9462 (N_9462,N_8474,N_8736);
nand U9463 (N_9463,N_8311,N_8795);
or U9464 (N_9464,N_8877,N_8488);
nand U9465 (N_9465,N_8690,N_8197);
nand U9466 (N_9466,N_8184,N_8639);
and U9467 (N_9467,N_8732,N_8373);
or U9468 (N_9468,N_8377,N_8895);
nor U9469 (N_9469,N_8525,N_8575);
nand U9470 (N_9470,N_8807,N_8569);
and U9471 (N_9471,N_8982,N_8948);
nand U9472 (N_9472,N_8046,N_8148);
nand U9473 (N_9473,N_8155,N_8623);
or U9474 (N_9474,N_8436,N_8302);
and U9475 (N_9475,N_8281,N_8124);
nand U9476 (N_9476,N_8090,N_8520);
or U9477 (N_9477,N_8021,N_8211);
or U9478 (N_9478,N_8919,N_8931);
and U9479 (N_9479,N_8535,N_8493);
nand U9480 (N_9480,N_8095,N_8864);
or U9481 (N_9481,N_8196,N_8229);
or U9482 (N_9482,N_8454,N_8333);
and U9483 (N_9483,N_8403,N_8805);
or U9484 (N_9484,N_8738,N_8266);
nor U9485 (N_9485,N_8689,N_8819);
and U9486 (N_9486,N_8087,N_8462);
nand U9487 (N_9487,N_8779,N_8199);
nor U9488 (N_9488,N_8048,N_8146);
or U9489 (N_9489,N_8741,N_8903);
or U9490 (N_9490,N_8382,N_8727);
nand U9491 (N_9491,N_8597,N_8296);
and U9492 (N_9492,N_8092,N_8049);
nand U9493 (N_9493,N_8604,N_8269);
nand U9494 (N_9494,N_8849,N_8192);
nor U9495 (N_9495,N_8355,N_8853);
and U9496 (N_9496,N_8595,N_8250);
or U9497 (N_9497,N_8954,N_8558);
nor U9498 (N_9498,N_8686,N_8091);
and U9499 (N_9499,N_8418,N_8935);
nor U9500 (N_9500,N_8160,N_8700);
and U9501 (N_9501,N_8885,N_8929);
nor U9502 (N_9502,N_8806,N_8572);
nor U9503 (N_9503,N_8956,N_8663);
and U9504 (N_9504,N_8814,N_8647);
nand U9505 (N_9505,N_8779,N_8839);
or U9506 (N_9506,N_8664,N_8877);
nor U9507 (N_9507,N_8088,N_8929);
nor U9508 (N_9508,N_8131,N_8277);
nor U9509 (N_9509,N_8875,N_8179);
nor U9510 (N_9510,N_8111,N_8343);
nor U9511 (N_9511,N_8172,N_8749);
or U9512 (N_9512,N_8475,N_8167);
nand U9513 (N_9513,N_8504,N_8703);
and U9514 (N_9514,N_8614,N_8967);
or U9515 (N_9515,N_8706,N_8505);
or U9516 (N_9516,N_8688,N_8968);
and U9517 (N_9517,N_8237,N_8886);
and U9518 (N_9518,N_8756,N_8908);
nand U9519 (N_9519,N_8180,N_8407);
or U9520 (N_9520,N_8750,N_8112);
nand U9521 (N_9521,N_8501,N_8618);
or U9522 (N_9522,N_8062,N_8144);
nand U9523 (N_9523,N_8080,N_8485);
nand U9524 (N_9524,N_8429,N_8718);
nor U9525 (N_9525,N_8952,N_8361);
nor U9526 (N_9526,N_8598,N_8938);
nor U9527 (N_9527,N_8490,N_8731);
nor U9528 (N_9528,N_8071,N_8551);
nor U9529 (N_9529,N_8542,N_8034);
nor U9530 (N_9530,N_8995,N_8588);
and U9531 (N_9531,N_8970,N_8003);
or U9532 (N_9532,N_8735,N_8501);
or U9533 (N_9533,N_8121,N_8494);
nor U9534 (N_9534,N_8262,N_8551);
and U9535 (N_9535,N_8643,N_8009);
nor U9536 (N_9536,N_8013,N_8815);
nor U9537 (N_9537,N_8935,N_8304);
nor U9538 (N_9538,N_8840,N_8720);
or U9539 (N_9539,N_8090,N_8460);
and U9540 (N_9540,N_8933,N_8790);
or U9541 (N_9541,N_8626,N_8514);
nand U9542 (N_9542,N_8723,N_8985);
nand U9543 (N_9543,N_8012,N_8039);
nor U9544 (N_9544,N_8872,N_8775);
nor U9545 (N_9545,N_8737,N_8797);
nor U9546 (N_9546,N_8614,N_8929);
nor U9547 (N_9547,N_8842,N_8144);
or U9548 (N_9548,N_8916,N_8102);
and U9549 (N_9549,N_8524,N_8900);
and U9550 (N_9550,N_8001,N_8770);
nor U9551 (N_9551,N_8538,N_8172);
or U9552 (N_9552,N_8095,N_8328);
nor U9553 (N_9553,N_8383,N_8368);
nand U9554 (N_9554,N_8143,N_8857);
nor U9555 (N_9555,N_8572,N_8762);
or U9556 (N_9556,N_8625,N_8158);
nor U9557 (N_9557,N_8373,N_8158);
nor U9558 (N_9558,N_8600,N_8043);
nor U9559 (N_9559,N_8626,N_8185);
and U9560 (N_9560,N_8089,N_8249);
nand U9561 (N_9561,N_8484,N_8103);
and U9562 (N_9562,N_8911,N_8203);
nor U9563 (N_9563,N_8857,N_8450);
nor U9564 (N_9564,N_8379,N_8119);
or U9565 (N_9565,N_8427,N_8148);
and U9566 (N_9566,N_8689,N_8355);
or U9567 (N_9567,N_8242,N_8488);
nor U9568 (N_9568,N_8606,N_8165);
nand U9569 (N_9569,N_8157,N_8727);
nor U9570 (N_9570,N_8103,N_8265);
or U9571 (N_9571,N_8725,N_8682);
and U9572 (N_9572,N_8963,N_8248);
nor U9573 (N_9573,N_8321,N_8334);
nand U9574 (N_9574,N_8929,N_8894);
or U9575 (N_9575,N_8734,N_8865);
and U9576 (N_9576,N_8315,N_8646);
nor U9577 (N_9577,N_8855,N_8858);
nor U9578 (N_9578,N_8822,N_8212);
nand U9579 (N_9579,N_8869,N_8566);
and U9580 (N_9580,N_8937,N_8736);
and U9581 (N_9581,N_8494,N_8232);
nor U9582 (N_9582,N_8095,N_8142);
nand U9583 (N_9583,N_8457,N_8817);
nor U9584 (N_9584,N_8154,N_8702);
and U9585 (N_9585,N_8051,N_8617);
nand U9586 (N_9586,N_8161,N_8966);
nor U9587 (N_9587,N_8812,N_8342);
or U9588 (N_9588,N_8163,N_8387);
or U9589 (N_9589,N_8005,N_8128);
nor U9590 (N_9590,N_8926,N_8282);
or U9591 (N_9591,N_8318,N_8665);
nor U9592 (N_9592,N_8209,N_8100);
nand U9593 (N_9593,N_8273,N_8051);
and U9594 (N_9594,N_8315,N_8097);
nand U9595 (N_9595,N_8786,N_8783);
nor U9596 (N_9596,N_8362,N_8356);
or U9597 (N_9597,N_8769,N_8918);
and U9598 (N_9598,N_8247,N_8072);
nand U9599 (N_9599,N_8242,N_8645);
nor U9600 (N_9600,N_8276,N_8564);
nand U9601 (N_9601,N_8835,N_8097);
and U9602 (N_9602,N_8281,N_8718);
or U9603 (N_9603,N_8910,N_8608);
nand U9604 (N_9604,N_8100,N_8845);
nand U9605 (N_9605,N_8314,N_8384);
and U9606 (N_9606,N_8313,N_8381);
nand U9607 (N_9607,N_8316,N_8618);
or U9608 (N_9608,N_8287,N_8221);
xnor U9609 (N_9609,N_8704,N_8393);
nor U9610 (N_9610,N_8650,N_8407);
or U9611 (N_9611,N_8656,N_8159);
and U9612 (N_9612,N_8431,N_8574);
nor U9613 (N_9613,N_8914,N_8489);
nand U9614 (N_9614,N_8412,N_8598);
nand U9615 (N_9615,N_8488,N_8170);
nand U9616 (N_9616,N_8009,N_8107);
or U9617 (N_9617,N_8335,N_8047);
or U9618 (N_9618,N_8459,N_8196);
and U9619 (N_9619,N_8097,N_8531);
and U9620 (N_9620,N_8726,N_8793);
and U9621 (N_9621,N_8476,N_8441);
nor U9622 (N_9622,N_8144,N_8642);
nor U9623 (N_9623,N_8746,N_8012);
xnor U9624 (N_9624,N_8039,N_8629);
or U9625 (N_9625,N_8539,N_8299);
nand U9626 (N_9626,N_8473,N_8750);
nor U9627 (N_9627,N_8337,N_8350);
or U9628 (N_9628,N_8759,N_8549);
or U9629 (N_9629,N_8275,N_8300);
and U9630 (N_9630,N_8934,N_8353);
nand U9631 (N_9631,N_8914,N_8531);
or U9632 (N_9632,N_8538,N_8369);
nand U9633 (N_9633,N_8642,N_8306);
nor U9634 (N_9634,N_8940,N_8560);
or U9635 (N_9635,N_8840,N_8170);
nor U9636 (N_9636,N_8293,N_8552);
or U9637 (N_9637,N_8815,N_8621);
or U9638 (N_9638,N_8510,N_8504);
and U9639 (N_9639,N_8309,N_8791);
nor U9640 (N_9640,N_8404,N_8408);
or U9641 (N_9641,N_8810,N_8013);
nand U9642 (N_9642,N_8720,N_8216);
and U9643 (N_9643,N_8068,N_8030);
nor U9644 (N_9644,N_8460,N_8294);
and U9645 (N_9645,N_8478,N_8601);
and U9646 (N_9646,N_8304,N_8044);
nor U9647 (N_9647,N_8316,N_8069);
or U9648 (N_9648,N_8925,N_8579);
nand U9649 (N_9649,N_8517,N_8446);
nand U9650 (N_9650,N_8125,N_8444);
or U9651 (N_9651,N_8640,N_8320);
and U9652 (N_9652,N_8960,N_8088);
nor U9653 (N_9653,N_8068,N_8165);
and U9654 (N_9654,N_8115,N_8306);
nand U9655 (N_9655,N_8476,N_8807);
and U9656 (N_9656,N_8096,N_8801);
nand U9657 (N_9657,N_8768,N_8112);
nor U9658 (N_9658,N_8173,N_8343);
and U9659 (N_9659,N_8403,N_8705);
nand U9660 (N_9660,N_8275,N_8945);
nand U9661 (N_9661,N_8388,N_8700);
and U9662 (N_9662,N_8156,N_8879);
nand U9663 (N_9663,N_8767,N_8230);
nand U9664 (N_9664,N_8483,N_8132);
and U9665 (N_9665,N_8670,N_8373);
and U9666 (N_9666,N_8905,N_8874);
nor U9667 (N_9667,N_8821,N_8335);
nor U9668 (N_9668,N_8501,N_8328);
and U9669 (N_9669,N_8602,N_8183);
and U9670 (N_9670,N_8569,N_8641);
nor U9671 (N_9671,N_8796,N_8005);
nor U9672 (N_9672,N_8517,N_8166);
or U9673 (N_9673,N_8385,N_8219);
nor U9674 (N_9674,N_8498,N_8070);
and U9675 (N_9675,N_8718,N_8381);
or U9676 (N_9676,N_8696,N_8574);
or U9677 (N_9677,N_8751,N_8341);
nand U9678 (N_9678,N_8373,N_8507);
and U9679 (N_9679,N_8591,N_8876);
and U9680 (N_9680,N_8503,N_8045);
or U9681 (N_9681,N_8018,N_8339);
or U9682 (N_9682,N_8794,N_8684);
nand U9683 (N_9683,N_8267,N_8797);
nand U9684 (N_9684,N_8437,N_8958);
or U9685 (N_9685,N_8996,N_8590);
and U9686 (N_9686,N_8791,N_8441);
or U9687 (N_9687,N_8059,N_8794);
or U9688 (N_9688,N_8799,N_8374);
nor U9689 (N_9689,N_8171,N_8160);
or U9690 (N_9690,N_8708,N_8117);
or U9691 (N_9691,N_8658,N_8778);
or U9692 (N_9692,N_8110,N_8719);
nand U9693 (N_9693,N_8003,N_8654);
nand U9694 (N_9694,N_8036,N_8585);
or U9695 (N_9695,N_8592,N_8985);
nand U9696 (N_9696,N_8251,N_8250);
nand U9697 (N_9697,N_8777,N_8550);
nand U9698 (N_9698,N_8186,N_8671);
nand U9699 (N_9699,N_8204,N_8923);
nor U9700 (N_9700,N_8707,N_8322);
or U9701 (N_9701,N_8952,N_8410);
nand U9702 (N_9702,N_8118,N_8460);
and U9703 (N_9703,N_8926,N_8448);
nand U9704 (N_9704,N_8824,N_8260);
and U9705 (N_9705,N_8091,N_8504);
or U9706 (N_9706,N_8828,N_8819);
nor U9707 (N_9707,N_8323,N_8885);
and U9708 (N_9708,N_8793,N_8357);
nor U9709 (N_9709,N_8211,N_8036);
nand U9710 (N_9710,N_8504,N_8173);
nand U9711 (N_9711,N_8308,N_8554);
and U9712 (N_9712,N_8732,N_8433);
or U9713 (N_9713,N_8789,N_8818);
xnor U9714 (N_9714,N_8293,N_8085);
nor U9715 (N_9715,N_8047,N_8334);
nor U9716 (N_9716,N_8749,N_8842);
or U9717 (N_9717,N_8352,N_8281);
and U9718 (N_9718,N_8559,N_8915);
or U9719 (N_9719,N_8903,N_8960);
and U9720 (N_9720,N_8703,N_8925);
or U9721 (N_9721,N_8426,N_8969);
nand U9722 (N_9722,N_8351,N_8147);
nor U9723 (N_9723,N_8736,N_8001);
nor U9724 (N_9724,N_8183,N_8659);
nand U9725 (N_9725,N_8998,N_8864);
or U9726 (N_9726,N_8372,N_8194);
and U9727 (N_9727,N_8146,N_8001);
nand U9728 (N_9728,N_8063,N_8176);
or U9729 (N_9729,N_8555,N_8575);
and U9730 (N_9730,N_8393,N_8183);
or U9731 (N_9731,N_8425,N_8148);
nand U9732 (N_9732,N_8700,N_8757);
nand U9733 (N_9733,N_8030,N_8394);
and U9734 (N_9734,N_8454,N_8421);
or U9735 (N_9735,N_8157,N_8021);
nand U9736 (N_9736,N_8661,N_8733);
and U9737 (N_9737,N_8617,N_8225);
xnor U9738 (N_9738,N_8757,N_8642);
nand U9739 (N_9739,N_8147,N_8433);
nor U9740 (N_9740,N_8223,N_8351);
or U9741 (N_9741,N_8195,N_8364);
nor U9742 (N_9742,N_8788,N_8720);
and U9743 (N_9743,N_8966,N_8996);
nand U9744 (N_9744,N_8418,N_8716);
or U9745 (N_9745,N_8528,N_8639);
nor U9746 (N_9746,N_8692,N_8204);
nor U9747 (N_9747,N_8347,N_8769);
nor U9748 (N_9748,N_8692,N_8606);
nor U9749 (N_9749,N_8384,N_8524);
or U9750 (N_9750,N_8053,N_8881);
nor U9751 (N_9751,N_8329,N_8242);
nor U9752 (N_9752,N_8173,N_8703);
nand U9753 (N_9753,N_8070,N_8934);
nand U9754 (N_9754,N_8067,N_8846);
nor U9755 (N_9755,N_8791,N_8640);
and U9756 (N_9756,N_8969,N_8601);
nor U9757 (N_9757,N_8112,N_8362);
nand U9758 (N_9758,N_8512,N_8838);
nand U9759 (N_9759,N_8144,N_8923);
and U9760 (N_9760,N_8182,N_8937);
nand U9761 (N_9761,N_8121,N_8373);
nand U9762 (N_9762,N_8643,N_8556);
and U9763 (N_9763,N_8324,N_8561);
nor U9764 (N_9764,N_8033,N_8267);
or U9765 (N_9765,N_8019,N_8205);
or U9766 (N_9766,N_8236,N_8514);
nand U9767 (N_9767,N_8063,N_8625);
nand U9768 (N_9768,N_8018,N_8965);
or U9769 (N_9769,N_8744,N_8669);
nor U9770 (N_9770,N_8541,N_8994);
nor U9771 (N_9771,N_8231,N_8260);
nand U9772 (N_9772,N_8999,N_8783);
and U9773 (N_9773,N_8895,N_8406);
or U9774 (N_9774,N_8116,N_8521);
nor U9775 (N_9775,N_8587,N_8288);
nand U9776 (N_9776,N_8086,N_8141);
nand U9777 (N_9777,N_8974,N_8595);
nor U9778 (N_9778,N_8812,N_8539);
nor U9779 (N_9779,N_8832,N_8090);
nor U9780 (N_9780,N_8047,N_8601);
nor U9781 (N_9781,N_8961,N_8551);
or U9782 (N_9782,N_8903,N_8444);
and U9783 (N_9783,N_8339,N_8290);
nand U9784 (N_9784,N_8715,N_8348);
and U9785 (N_9785,N_8442,N_8520);
nor U9786 (N_9786,N_8994,N_8889);
and U9787 (N_9787,N_8386,N_8892);
nand U9788 (N_9788,N_8928,N_8667);
nand U9789 (N_9789,N_8900,N_8016);
nor U9790 (N_9790,N_8525,N_8053);
nand U9791 (N_9791,N_8485,N_8670);
nor U9792 (N_9792,N_8089,N_8664);
and U9793 (N_9793,N_8065,N_8653);
or U9794 (N_9794,N_8454,N_8527);
nand U9795 (N_9795,N_8778,N_8129);
nand U9796 (N_9796,N_8195,N_8232);
nor U9797 (N_9797,N_8781,N_8583);
nand U9798 (N_9798,N_8290,N_8486);
or U9799 (N_9799,N_8295,N_8386);
nand U9800 (N_9800,N_8570,N_8781);
or U9801 (N_9801,N_8710,N_8285);
and U9802 (N_9802,N_8428,N_8092);
nor U9803 (N_9803,N_8982,N_8827);
or U9804 (N_9804,N_8509,N_8724);
and U9805 (N_9805,N_8672,N_8912);
or U9806 (N_9806,N_8478,N_8661);
nand U9807 (N_9807,N_8132,N_8827);
or U9808 (N_9808,N_8512,N_8848);
nor U9809 (N_9809,N_8847,N_8496);
or U9810 (N_9810,N_8608,N_8866);
nand U9811 (N_9811,N_8708,N_8551);
or U9812 (N_9812,N_8173,N_8860);
nor U9813 (N_9813,N_8957,N_8270);
or U9814 (N_9814,N_8445,N_8425);
nor U9815 (N_9815,N_8846,N_8971);
and U9816 (N_9816,N_8531,N_8887);
or U9817 (N_9817,N_8308,N_8714);
or U9818 (N_9818,N_8862,N_8182);
and U9819 (N_9819,N_8038,N_8582);
or U9820 (N_9820,N_8180,N_8716);
nor U9821 (N_9821,N_8497,N_8649);
and U9822 (N_9822,N_8570,N_8555);
xnor U9823 (N_9823,N_8114,N_8920);
nand U9824 (N_9824,N_8269,N_8229);
nand U9825 (N_9825,N_8658,N_8878);
or U9826 (N_9826,N_8204,N_8614);
nand U9827 (N_9827,N_8839,N_8163);
xor U9828 (N_9828,N_8264,N_8814);
nor U9829 (N_9829,N_8307,N_8645);
nand U9830 (N_9830,N_8972,N_8021);
nand U9831 (N_9831,N_8057,N_8169);
nand U9832 (N_9832,N_8095,N_8064);
or U9833 (N_9833,N_8475,N_8065);
and U9834 (N_9834,N_8501,N_8857);
nand U9835 (N_9835,N_8629,N_8677);
and U9836 (N_9836,N_8124,N_8674);
and U9837 (N_9837,N_8015,N_8891);
xor U9838 (N_9838,N_8878,N_8127);
or U9839 (N_9839,N_8741,N_8415);
or U9840 (N_9840,N_8390,N_8420);
nand U9841 (N_9841,N_8852,N_8115);
and U9842 (N_9842,N_8014,N_8893);
or U9843 (N_9843,N_8634,N_8880);
nor U9844 (N_9844,N_8042,N_8018);
nor U9845 (N_9845,N_8907,N_8988);
or U9846 (N_9846,N_8845,N_8484);
or U9847 (N_9847,N_8409,N_8877);
nor U9848 (N_9848,N_8336,N_8667);
nor U9849 (N_9849,N_8934,N_8446);
nor U9850 (N_9850,N_8578,N_8800);
and U9851 (N_9851,N_8553,N_8350);
or U9852 (N_9852,N_8137,N_8300);
nand U9853 (N_9853,N_8104,N_8747);
and U9854 (N_9854,N_8629,N_8744);
and U9855 (N_9855,N_8250,N_8764);
nor U9856 (N_9856,N_8021,N_8247);
or U9857 (N_9857,N_8662,N_8532);
or U9858 (N_9858,N_8334,N_8500);
nor U9859 (N_9859,N_8302,N_8036);
nor U9860 (N_9860,N_8071,N_8637);
nand U9861 (N_9861,N_8343,N_8989);
or U9862 (N_9862,N_8936,N_8709);
and U9863 (N_9863,N_8260,N_8873);
or U9864 (N_9864,N_8513,N_8526);
nor U9865 (N_9865,N_8332,N_8266);
nor U9866 (N_9866,N_8539,N_8653);
nand U9867 (N_9867,N_8128,N_8253);
and U9868 (N_9868,N_8534,N_8217);
nand U9869 (N_9869,N_8665,N_8422);
nand U9870 (N_9870,N_8150,N_8133);
and U9871 (N_9871,N_8314,N_8317);
or U9872 (N_9872,N_8827,N_8947);
or U9873 (N_9873,N_8291,N_8105);
nor U9874 (N_9874,N_8995,N_8499);
nor U9875 (N_9875,N_8306,N_8126);
and U9876 (N_9876,N_8487,N_8513);
nor U9877 (N_9877,N_8815,N_8193);
nor U9878 (N_9878,N_8135,N_8969);
nor U9879 (N_9879,N_8181,N_8481);
or U9880 (N_9880,N_8597,N_8237);
and U9881 (N_9881,N_8737,N_8002);
nor U9882 (N_9882,N_8933,N_8471);
nand U9883 (N_9883,N_8704,N_8516);
nor U9884 (N_9884,N_8427,N_8848);
or U9885 (N_9885,N_8079,N_8501);
nand U9886 (N_9886,N_8725,N_8127);
or U9887 (N_9887,N_8050,N_8252);
or U9888 (N_9888,N_8055,N_8294);
nand U9889 (N_9889,N_8626,N_8971);
or U9890 (N_9890,N_8370,N_8640);
nor U9891 (N_9891,N_8268,N_8996);
or U9892 (N_9892,N_8489,N_8467);
nand U9893 (N_9893,N_8043,N_8059);
or U9894 (N_9894,N_8224,N_8399);
nand U9895 (N_9895,N_8456,N_8611);
nand U9896 (N_9896,N_8355,N_8690);
nor U9897 (N_9897,N_8951,N_8531);
and U9898 (N_9898,N_8267,N_8606);
nand U9899 (N_9899,N_8919,N_8155);
and U9900 (N_9900,N_8068,N_8937);
or U9901 (N_9901,N_8914,N_8055);
nor U9902 (N_9902,N_8620,N_8109);
or U9903 (N_9903,N_8181,N_8701);
and U9904 (N_9904,N_8176,N_8759);
nor U9905 (N_9905,N_8587,N_8257);
nor U9906 (N_9906,N_8706,N_8248);
nand U9907 (N_9907,N_8198,N_8087);
and U9908 (N_9908,N_8702,N_8976);
or U9909 (N_9909,N_8560,N_8381);
nor U9910 (N_9910,N_8904,N_8432);
nand U9911 (N_9911,N_8901,N_8110);
or U9912 (N_9912,N_8847,N_8231);
and U9913 (N_9913,N_8040,N_8511);
nor U9914 (N_9914,N_8046,N_8709);
or U9915 (N_9915,N_8560,N_8861);
or U9916 (N_9916,N_8089,N_8342);
nor U9917 (N_9917,N_8866,N_8384);
and U9918 (N_9918,N_8134,N_8573);
nand U9919 (N_9919,N_8883,N_8800);
and U9920 (N_9920,N_8912,N_8201);
and U9921 (N_9921,N_8700,N_8038);
nand U9922 (N_9922,N_8852,N_8353);
or U9923 (N_9923,N_8154,N_8468);
nor U9924 (N_9924,N_8508,N_8511);
or U9925 (N_9925,N_8239,N_8189);
or U9926 (N_9926,N_8296,N_8993);
or U9927 (N_9927,N_8888,N_8550);
nand U9928 (N_9928,N_8763,N_8255);
nor U9929 (N_9929,N_8643,N_8750);
nand U9930 (N_9930,N_8472,N_8952);
and U9931 (N_9931,N_8130,N_8990);
nor U9932 (N_9932,N_8745,N_8686);
nor U9933 (N_9933,N_8864,N_8543);
or U9934 (N_9934,N_8785,N_8842);
nand U9935 (N_9935,N_8043,N_8350);
or U9936 (N_9936,N_8259,N_8695);
or U9937 (N_9937,N_8784,N_8043);
and U9938 (N_9938,N_8284,N_8471);
nor U9939 (N_9939,N_8266,N_8655);
nor U9940 (N_9940,N_8176,N_8985);
and U9941 (N_9941,N_8130,N_8968);
or U9942 (N_9942,N_8373,N_8791);
or U9943 (N_9943,N_8888,N_8768);
and U9944 (N_9944,N_8093,N_8283);
nand U9945 (N_9945,N_8579,N_8882);
and U9946 (N_9946,N_8481,N_8103);
and U9947 (N_9947,N_8966,N_8545);
and U9948 (N_9948,N_8369,N_8984);
and U9949 (N_9949,N_8025,N_8144);
nor U9950 (N_9950,N_8434,N_8182);
or U9951 (N_9951,N_8565,N_8228);
nor U9952 (N_9952,N_8893,N_8621);
and U9953 (N_9953,N_8463,N_8866);
or U9954 (N_9954,N_8665,N_8949);
nand U9955 (N_9955,N_8253,N_8164);
or U9956 (N_9956,N_8248,N_8967);
nor U9957 (N_9957,N_8338,N_8354);
and U9958 (N_9958,N_8362,N_8065);
or U9959 (N_9959,N_8897,N_8409);
nand U9960 (N_9960,N_8085,N_8632);
or U9961 (N_9961,N_8106,N_8050);
nand U9962 (N_9962,N_8209,N_8541);
nor U9963 (N_9963,N_8629,N_8887);
nand U9964 (N_9964,N_8319,N_8488);
nor U9965 (N_9965,N_8707,N_8714);
nor U9966 (N_9966,N_8446,N_8716);
nand U9967 (N_9967,N_8547,N_8402);
or U9968 (N_9968,N_8261,N_8402);
and U9969 (N_9969,N_8994,N_8904);
and U9970 (N_9970,N_8034,N_8425);
nor U9971 (N_9971,N_8859,N_8652);
and U9972 (N_9972,N_8522,N_8252);
nor U9973 (N_9973,N_8005,N_8524);
nand U9974 (N_9974,N_8365,N_8822);
or U9975 (N_9975,N_8299,N_8870);
and U9976 (N_9976,N_8891,N_8763);
nand U9977 (N_9977,N_8695,N_8197);
nor U9978 (N_9978,N_8653,N_8749);
nand U9979 (N_9979,N_8189,N_8174);
and U9980 (N_9980,N_8917,N_8631);
and U9981 (N_9981,N_8242,N_8872);
and U9982 (N_9982,N_8044,N_8162);
nand U9983 (N_9983,N_8915,N_8317);
and U9984 (N_9984,N_8094,N_8472);
or U9985 (N_9985,N_8356,N_8620);
or U9986 (N_9986,N_8158,N_8580);
nor U9987 (N_9987,N_8874,N_8386);
or U9988 (N_9988,N_8112,N_8918);
nor U9989 (N_9989,N_8645,N_8959);
or U9990 (N_9990,N_8884,N_8639);
or U9991 (N_9991,N_8161,N_8005);
or U9992 (N_9992,N_8130,N_8864);
and U9993 (N_9993,N_8340,N_8613);
and U9994 (N_9994,N_8172,N_8899);
nor U9995 (N_9995,N_8590,N_8304);
or U9996 (N_9996,N_8166,N_8125);
nand U9997 (N_9997,N_8245,N_8849);
nand U9998 (N_9998,N_8233,N_8099);
nor U9999 (N_9999,N_8180,N_8814);
nor UO_0 (O_0,N_9136,N_9506);
nor UO_1 (O_1,N_9759,N_9826);
or UO_2 (O_2,N_9392,N_9628);
nor UO_3 (O_3,N_9508,N_9089);
nor UO_4 (O_4,N_9597,N_9321);
or UO_5 (O_5,N_9480,N_9630);
and UO_6 (O_6,N_9920,N_9510);
nand UO_7 (O_7,N_9302,N_9256);
nand UO_8 (O_8,N_9808,N_9716);
nand UO_9 (O_9,N_9145,N_9165);
nand UO_10 (O_10,N_9554,N_9365);
or UO_11 (O_11,N_9865,N_9912);
or UO_12 (O_12,N_9450,N_9758);
and UO_13 (O_13,N_9278,N_9542);
nand UO_14 (O_14,N_9440,N_9271);
and UO_15 (O_15,N_9169,N_9578);
nand UO_16 (O_16,N_9997,N_9724);
nand UO_17 (O_17,N_9660,N_9112);
nand UO_18 (O_18,N_9364,N_9613);
or UO_19 (O_19,N_9872,N_9025);
nand UO_20 (O_20,N_9943,N_9174);
or UO_21 (O_21,N_9668,N_9220);
nor UO_22 (O_22,N_9252,N_9176);
or UO_23 (O_23,N_9884,N_9466);
nor UO_24 (O_24,N_9459,N_9074);
and UO_25 (O_25,N_9529,N_9790);
and UO_26 (O_26,N_9345,N_9373);
nand UO_27 (O_27,N_9347,N_9622);
or UO_28 (O_28,N_9532,N_9414);
or UO_29 (O_29,N_9667,N_9471);
nor UO_30 (O_30,N_9188,N_9656);
and UO_31 (O_31,N_9491,N_9571);
or UO_32 (O_32,N_9178,N_9019);
or UO_33 (O_33,N_9574,N_9675);
nand UO_34 (O_34,N_9946,N_9513);
and UO_35 (O_35,N_9703,N_9505);
nand UO_36 (O_36,N_9335,N_9827);
or UO_37 (O_37,N_9251,N_9443);
nand UO_38 (O_38,N_9205,N_9447);
nand UO_39 (O_39,N_9706,N_9867);
and UO_40 (O_40,N_9402,N_9346);
nand UO_41 (O_41,N_9473,N_9782);
and UO_42 (O_42,N_9658,N_9576);
nor UO_43 (O_43,N_9148,N_9989);
xnor UO_44 (O_44,N_9783,N_9289);
or UO_45 (O_45,N_9319,N_9722);
and UO_46 (O_46,N_9767,N_9953);
nor UO_47 (O_47,N_9073,N_9585);
and UO_48 (O_48,N_9963,N_9789);
nand UO_49 (O_49,N_9751,N_9183);
nor UO_50 (O_50,N_9270,N_9031);
and UO_51 (O_51,N_9549,N_9312);
nand UO_52 (O_52,N_9914,N_9893);
nand UO_53 (O_53,N_9299,N_9705);
nor UO_54 (O_54,N_9199,N_9938);
nand UO_55 (O_55,N_9247,N_9113);
nor UO_56 (O_56,N_9540,N_9137);
and UO_57 (O_57,N_9777,N_9330);
and UO_58 (O_58,N_9901,N_9744);
nor UO_59 (O_59,N_9900,N_9971);
nor UO_60 (O_60,N_9479,N_9088);
nor UO_61 (O_61,N_9388,N_9748);
or UO_62 (O_62,N_9063,N_9225);
or UO_63 (O_63,N_9472,N_9755);
nand UO_64 (O_64,N_9526,N_9339);
nand UO_65 (O_65,N_9191,N_9348);
or UO_66 (O_66,N_9184,N_9547);
nor UO_67 (O_67,N_9024,N_9179);
and UO_68 (O_68,N_9951,N_9712);
and UO_69 (O_69,N_9422,N_9700);
and UO_70 (O_70,N_9528,N_9887);
or UO_71 (O_71,N_9754,N_9486);
or UO_72 (O_72,N_9817,N_9014);
or UO_73 (O_73,N_9670,N_9400);
nor UO_74 (O_74,N_9581,N_9367);
nor UO_75 (O_75,N_9389,N_9882);
or UO_76 (O_76,N_9053,N_9322);
and UO_77 (O_77,N_9046,N_9674);
nand UO_78 (O_78,N_9217,N_9383);
nand UO_79 (O_79,N_9854,N_9931);
nand UO_80 (O_80,N_9150,N_9729);
or UO_81 (O_81,N_9430,N_9892);
and UO_82 (O_82,N_9693,N_9678);
nand UO_83 (O_83,N_9267,N_9906);
nand UO_84 (O_84,N_9833,N_9069);
nor UO_85 (O_85,N_9695,N_9066);
nor UO_86 (O_86,N_9370,N_9701);
and UO_87 (O_87,N_9929,N_9657);
nor UO_88 (O_88,N_9326,N_9115);
nand UO_89 (O_89,N_9930,N_9598);
nor UO_90 (O_90,N_9377,N_9149);
and UO_91 (O_91,N_9232,N_9669);
and UO_92 (O_92,N_9993,N_9194);
or UO_93 (O_93,N_9286,N_9504);
or UO_94 (O_94,N_9425,N_9798);
nor UO_95 (O_95,N_9707,N_9041);
or UO_96 (O_96,N_9881,N_9276);
or UO_97 (O_97,N_9093,N_9921);
or UO_98 (O_98,N_9616,N_9406);
or UO_99 (O_99,N_9838,N_9134);
or UO_100 (O_100,N_9792,N_9791);
nand UO_101 (O_101,N_9845,N_9449);
nand UO_102 (O_102,N_9028,N_9825);
nand UO_103 (O_103,N_9720,N_9012);
or UO_104 (O_104,N_9563,N_9966);
and UO_105 (O_105,N_9987,N_9502);
nor UO_106 (O_106,N_9594,N_9280);
and UO_107 (O_107,N_9804,N_9002);
or UO_108 (O_108,N_9683,N_9647);
or UO_109 (O_109,N_9233,N_9124);
nand UO_110 (O_110,N_9340,N_9638);
nand UO_111 (O_111,N_9650,N_9907);
nor UO_112 (O_112,N_9095,N_9342);
nand UO_113 (O_113,N_9062,N_9773);
and UO_114 (O_114,N_9806,N_9379);
nor UO_115 (O_115,N_9454,N_9432);
or UO_116 (O_116,N_9318,N_9663);
nand UO_117 (O_117,N_9990,N_9544);
nand UO_118 (O_118,N_9551,N_9810);
and UO_119 (O_119,N_9283,N_9537);
xor UO_120 (O_120,N_9086,N_9249);
nor UO_121 (O_121,N_9128,N_9435);
nor UO_122 (O_122,N_9005,N_9519);
and UO_123 (O_123,N_9386,N_9204);
nand UO_124 (O_124,N_9468,N_9355);
or UO_125 (O_125,N_9016,N_9009);
nor UO_126 (O_126,N_9814,N_9242);
nand UO_127 (O_127,N_9076,N_9998);
nand UO_128 (O_128,N_9393,N_9306);
and UO_129 (O_129,N_9889,N_9079);
or UO_130 (O_130,N_9250,N_9463);
or UO_131 (O_131,N_9264,N_9610);
nand UO_132 (O_132,N_9894,N_9876);
nor UO_133 (O_133,N_9001,N_9784);
and UO_134 (O_134,N_9467,N_9444);
nor UO_135 (O_135,N_9054,N_9431);
and UO_136 (O_136,N_9317,N_9448);
nor UO_137 (O_137,N_9570,N_9111);
nand UO_138 (O_138,N_9273,N_9637);
nand UO_139 (O_139,N_9118,N_9164);
and UO_140 (O_140,N_9725,N_9438);
and UO_141 (O_141,N_9933,N_9254);
nor UO_142 (O_142,N_9090,N_9763);
or UO_143 (O_143,N_9764,N_9439);
or UO_144 (O_144,N_9044,N_9214);
or UO_145 (O_145,N_9428,N_9607);
or UO_146 (O_146,N_9999,N_9955);
nor UO_147 (O_147,N_9535,N_9923);
and UO_148 (O_148,N_9320,N_9555);
nor UO_149 (O_149,N_9620,N_9851);
nand UO_150 (O_150,N_9853,N_9635);
nor UO_151 (O_151,N_9421,N_9718);
nor UO_152 (O_152,N_9474,N_9499);
nor UO_153 (O_153,N_9922,N_9600);
and UO_154 (O_154,N_9332,N_9794);
and UO_155 (O_155,N_9558,N_9442);
and UO_156 (O_156,N_9941,N_9702);
nor UO_157 (O_157,N_9704,N_9582);
nor UO_158 (O_158,N_9483,N_9646);
nand UO_159 (O_159,N_9268,N_9536);
nor UO_160 (O_160,N_9434,N_9688);
nor UO_161 (O_161,N_9282,N_9445);
nand UO_162 (O_162,N_9307,N_9871);
and UO_163 (O_163,N_9160,N_9200);
nand UO_164 (O_164,N_9116,N_9151);
or UO_165 (O_165,N_9830,N_9836);
nor UO_166 (O_166,N_9885,N_9237);
nand UO_167 (O_167,N_9631,N_9212);
nand UO_168 (O_168,N_9916,N_9553);
nor UO_169 (O_169,N_9114,N_9329);
nand UO_170 (O_170,N_9932,N_9078);
and UO_171 (O_171,N_9296,N_9858);
xor UO_172 (O_172,N_9123,N_9524);
nand UO_173 (O_173,N_9588,N_9691);
nor UO_174 (O_174,N_9511,N_9800);
nand UO_175 (O_175,N_9643,N_9988);
nand UO_176 (O_176,N_9343,N_9244);
or UO_177 (O_177,N_9011,N_9580);
nand UO_178 (O_178,N_9354,N_9316);
or UO_179 (O_179,N_9070,N_9464);
nand UO_180 (O_180,N_9130,N_9618);
and UO_181 (O_181,N_9602,N_9737);
or UO_182 (O_182,N_9498,N_9485);
and UO_183 (O_183,N_9049,N_9301);
nor UO_184 (O_184,N_9293,N_9713);
and UO_185 (O_185,N_9711,N_9223);
nand UO_186 (O_186,N_9862,N_9795);
nand UO_187 (O_187,N_9632,N_9676);
nand UO_188 (O_188,N_9083,N_9786);
nand UO_189 (O_189,N_9008,N_9181);
nor UO_190 (O_190,N_9606,N_9822);
nor UO_191 (O_191,N_9805,N_9275);
nand UO_192 (O_192,N_9038,N_9924);
nor UO_193 (O_193,N_9013,N_9143);
and UO_194 (O_194,N_9153,N_9774);
nand UO_195 (O_195,N_9995,N_9222);
or UO_196 (O_196,N_9304,N_9747);
or UO_197 (O_197,N_9738,N_9935);
and UO_198 (O_198,N_9193,N_9577);
nor UO_199 (O_199,N_9409,N_9741);
or UO_200 (O_200,N_9557,N_9918);
nor UO_201 (O_201,N_9180,N_9021);
and UO_202 (O_202,N_9627,N_9144);
nor UO_203 (O_203,N_9915,N_9840);
or UO_204 (O_204,N_9868,N_9146);
and UO_205 (O_205,N_9664,N_9880);
or UO_206 (O_206,N_9189,N_9689);
nand UO_207 (O_207,N_9832,N_9949);
nor UO_208 (O_208,N_9541,N_9680);
nor UO_209 (O_209,N_9973,N_9352);
nand UO_210 (O_210,N_9040,N_9030);
nor UO_211 (O_211,N_9543,N_9241);
or UO_212 (O_212,N_9465,N_9055);
nor UO_213 (O_213,N_9295,N_9572);
nand UO_214 (O_214,N_9769,N_9801);
or UO_215 (O_215,N_9104,N_9746);
nand UO_216 (O_216,N_9727,N_9757);
and UO_217 (O_217,N_9215,N_9902);
nand UO_218 (O_218,N_9545,N_9441);
nand UO_219 (O_219,N_9015,N_9043);
or UO_220 (O_220,N_9325,N_9477);
or UO_221 (O_221,N_9539,N_9982);
nor UO_222 (O_222,N_9152,N_9719);
or UO_223 (O_223,N_9654,N_9102);
or UO_224 (O_224,N_9481,N_9141);
nor UO_225 (O_225,N_9202,N_9639);
and UO_226 (O_226,N_9775,N_9655);
or UO_227 (O_227,N_9385,N_9977);
and UO_228 (O_228,N_9297,N_9061);
and UO_229 (O_229,N_9484,N_9573);
nand UO_230 (O_230,N_9752,N_9404);
nor UO_231 (O_231,N_9133,N_9171);
nand UO_232 (O_232,N_9824,N_9978);
nand UO_233 (O_233,N_9677,N_9308);
nand UO_234 (O_234,N_9903,N_9257);
nor UO_235 (O_235,N_9029,N_9060);
nand UO_236 (O_236,N_9614,N_9258);
nand UO_237 (O_237,N_9586,N_9382);
nor UO_238 (O_238,N_9723,N_9287);
or UO_239 (O_239,N_9979,N_9904);
nor UO_240 (O_240,N_9899,N_9131);
nor UO_241 (O_241,N_9828,N_9546);
or UO_242 (O_242,N_9839,N_9850);
nor UO_243 (O_243,N_9229,N_9645);
or UO_244 (O_244,N_9624,N_9807);
and UO_245 (O_245,N_9818,N_9391);
nand UO_246 (O_246,N_9168,N_9972);
nor UO_247 (O_247,N_9952,N_9424);
nand UO_248 (O_248,N_9947,N_9652);
nand UO_249 (O_249,N_9636,N_9120);
and UO_250 (O_250,N_9023,N_9412);
and UO_251 (O_251,N_9405,N_9934);
and UO_252 (O_252,N_9052,N_9681);
or UO_253 (O_253,N_9410,N_9496);
nand UO_254 (O_254,N_9333,N_9939);
nand UO_255 (O_255,N_9567,N_9926);
nor UO_256 (O_256,N_9161,N_9714);
nor UO_257 (O_257,N_9453,N_9004);
or UO_258 (O_258,N_9452,N_9662);
and UO_259 (O_259,N_9936,N_9065);
xnor UO_260 (O_260,N_9080,N_9461);
or UO_261 (O_261,N_9026,N_9487);
nor UO_262 (O_262,N_9125,N_9139);
or UO_263 (O_263,N_9359,N_9064);
or UO_264 (O_264,N_9849,N_9905);
and UO_265 (O_265,N_9203,N_9583);
and UO_266 (O_266,N_9556,N_9512);
nor UO_267 (O_267,N_9803,N_9629);
nor UO_268 (O_268,N_9210,N_9960);
nor UO_269 (O_269,N_9928,N_9698);
nor UO_270 (O_270,N_9690,N_9490);
nor UO_271 (O_271,N_9384,N_9206);
nor UO_272 (O_272,N_9619,N_9211);
and UO_273 (O_273,N_9940,N_9132);
or UO_274 (O_274,N_9010,N_9615);
nand UO_275 (O_275,N_9328,N_9238);
nor UO_276 (O_276,N_9686,N_9360);
or UO_277 (O_277,N_9731,N_9173);
and UO_278 (O_278,N_9501,N_9560);
nor UO_279 (O_279,N_9843,N_9020);
and UO_280 (O_280,N_9740,N_9913);
or UO_281 (O_281,N_9240,N_9417);
nand UO_282 (O_282,N_9521,N_9778);
or UO_283 (O_283,N_9185,N_9122);
and UO_284 (O_284,N_9290,N_9277);
or UO_285 (O_285,N_9298,N_9671);
and UO_286 (O_286,N_9523,N_9589);
nor UO_287 (O_287,N_9870,N_9314);
nand UO_288 (O_288,N_9996,N_9397);
and UO_289 (O_289,N_9864,N_9059);
or UO_290 (O_290,N_9942,N_9310);
nand UO_291 (O_291,N_9075,N_9962);
and UO_292 (O_292,N_9592,N_9196);
or UO_293 (O_293,N_9909,N_9035);
or UO_294 (O_294,N_9739,N_9399);
or UO_295 (O_295,N_9208,N_9100);
and UO_296 (O_296,N_9209,N_9495);
and UO_297 (O_297,N_9494,N_9534);
nand UO_298 (O_298,N_9110,N_9927);
nand UO_299 (O_299,N_9155,N_9848);
or UO_300 (O_300,N_9623,N_9037);
and UO_301 (O_301,N_9138,N_9411);
and UO_302 (O_302,N_9047,N_9381);
nand UO_303 (O_303,N_9766,N_9228);
and UO_304 (O_304,N_9983,N_9129);
and UO_305 (O_305,N_9371,N_9599);
nand UO_306 (O_306,N_9891,N_9380);
xor UO_307 (O_307,N_9462,N_9372);
or UO_308 (O_308,N_9022,N_9231);
nand UO_309 (O_309,N_9834,N_9815);
and UO_310 (O_310,N_9538,N_9338);
nor UO_311 (O_311,N_9357,N_9107);
and UO_312 (O_312,N_9324,N_9961);
or UO_313 (O_313,N_9475,N_9919);
nor UO_314 (O_314,N_9263,N_9937);
and UO_315 (O_315,N_9785,N_9793);
nand UO_316 (O_316,N_9964,N_9207);
or UO_317 (O_317,N_9733,N_9245);
or UO_318 (O_318,N_9362,N_9094);
or UO_319 (O_319,N_9750,N_9067);
and UO_320 (O_320,N_9261,N_9562);
nand UO_321 (O_321,N_9696,N_9358);
and UO_322 (O_322,N_9835,N_9500);
or UO_323 (O_323,N_9157,N_9243);
and UO_324 (O_324,N_9423,N_9356);
nand UO_325 (O_325,N_9192,N_9569);
nor UO_326 (O_326,N_9552,N_9837);
nand UO_327 (O_327,N_9687,N_9427);
xor UO_328 (O_328,N_9482,N_9568);
nor UO_329 (O_329,N_9344,N_9732);
nor UO_330 (O_330,N_9559,N_9856);
nor UO_331 (O_331,N_9401,N_9875);
and UO_332 (O_332,N_9366,N_9831);
or UO_333 (O_333,N_9642,N_9768);
and UO_334 (O_334,N_9156,N_9811);
or UO_335 (O_335,N_9957,N_9956);
or UO_336 (O_336,N_9033,N_9072);
and UO_337 (O_337,N_9886,N_9413);
xnor UO_338 (O_338,N_9259,N_9708);
or UO_339 (O_339,N_9036,N_9844);
and UO_340 (O_340,N_9877,N_9561);
nand UO_341 (O_341,N_9959,N_9395);
and UO_342 (O_342,N_9857,N_9260);
nor UO_343 (O_343,N_9641,N_9984);
or UO_344 (O_344,N_9911,N_9699);
nand UO_345 (O_345,N_9895,N_9266);
xnor UO_346 (O_346,N_9077,N_9692);
or UO_347 (O_347,N_9341,N_9787);
or UO_348 (O_348,N_9368,N_9109);
or UO_349 (O_349,N_9595,N_9235);
nor UO_350 (O_350,N_9234,N_9167);
nand UO_351 (O_351,N_9760,N_9315);
or UO_352 (O_352,N_9269,N_9175);
or UO_353 (O_353,N_9458,N_9813);
nor UO_354 (O_354,N_9898,N_9027);
and UO_355 (O_355,N_9084,N_9796);
and UO_356 (O_356,N_9351,N_9292);
or UO_357 (O_357,N_9018,N_9403);
nand UO_358 (O_358,N_9085,N_9349);
or UO_359 (O_359,N_9661,N_9525);
nand UO_360 (O_360,N_9285,N_9633);
nor UO_361 (O_361,N_9520,N_9753);
nor UO_362 (O_362,N_9437,N_9396);
nor UO_363 (O_363,N_9533,N_9159);
nor UO_364 (O_364,N_9416,N_9878);
and UO_365 (O_365,N_9103,N_9866);
or UO_366 (O_366,N_9726,N_9227);
nand UO_367 (O_367,N_9514,N_9305);
or UO_368 (O_368,N_9612,N_9601);
nand UO_369 (O_369,N_9548,N_9954);
and UO_370 (O_370,N_9172,N_9772);
or UO_371 (O_371,N_9198,N_9456);
nor UO_372 (O_372,N_9651,N_9489);
nand UO_373 (O_373,N_9398,N_9994);
nor UO_374 (O_374,N_9756,N_9771);
and UO_375 (O_375,N_9042,N_9226);
nor UO_376 (O_376,N_9608,N_9644);
nor UO_377 (O_377,N_9730,N_9697);
nand UO_378 (O_378,N_9426,N_9742);
nand UO_379 (O_379,N_9334,N_9890);
nand UO_380 (O_380,N_9101,N_9820);
nor UO_381 (O_381,N_9045,N_9219);
nor UO_382 (O_382,N_9099,N_9596);
nand UO_383 (O_383,N_9039,N_9517);
and UO_384 (O_384,N_9378,N_9291);
nor UO_385 (O_385,N_9883,N_9281);
nor UO_386 (O_386,N_9418,N_9842);
nand UO_387 (O_387,N_9779,N_9788);
nor UO_388 (O_388,N_9087,N_9058);
nand UO_389 (O_389,N_9509,N_9313);
nor UO_390 (O_390,N_9311,N_9082);
or UO_391 (O_391,N_9584,N_9709);
nand UO_392 (O_392,N_9455,N_9974);
and UO_393 (O_393,N_9048,N_9390);
or UO_394 (O_394,N_9626,N_9369);
and UO_395 (O_395,N_9071,N_9003);
and UO_396 (O_396,N_9566,N_9518);
and UO_397 (O_397,N_9515,N_9847);
nor UO_398 (O_398,N_9522,N_9809);
nand UO_399 (O_399,N_9121,N_9861);
and UO_400 (O_400,N_9761,N_9694);
nor UO_401 (O_401,N_9050,N_9096);
nand UO_402 (O_402,N_9527,N_9166);
or UO_403 (O_403,N_9303,N_9190);
or UO_404 (O_404,N_9056,N_9488);
nand UO_405 (O_405,N_9991,N_9846);
nor UO_406 (O_406,N_9478,N_9816);
nor UO_407 (O_407,N_9195,N_9640);
nor UO_408 (O_408,N_9965,N_9216);
nor UO_409 (O_409,N_9976,N_9917);
and UO_410 (O_410,N_9309,N_9446);
and UO_411 (O_411,N_9213,N_9460);
nor UO_412 (O_412,N_9006,N_9869);
nor UO_413 (O_413,N_9605,N_9127);
nand UO_414 (O_414,N_9634,N_9253);
nor UO_415 (O_415,N_9743,N_9436);
nand UO_416 (O_416,N_9097,N_9429);
or UO_417 (O_417,N_9565,N_9564);
nand UO_418 (O_418,N_9715,N_9182);
nor UO_419 (O_419,N_9603,N_9140);
nor UO_420 (O_420,N_9162,N_9224);
nor UO_421 (O_421,N_9091,N_9279);
nor UO_422 (O_422,N_9336,N_9665);
and UO_423 (O_423,N_9590,N_9969);
xnor UO_424 (O_424,N_9879,N_9888);
and UO_425 (O_425,N_9717,N_9968);
nor UO_426 (O_426,N_9625,N_9648);
or UO_427 (O_427,N_9457,N_9967);
or UO_428 (O_428,N_9550,N_9821);
nor UO_429 (O_429,N_9980,N_9068);
and UO_430 (O_430,N_9673,N_9781);
or UO_431 (O_431,N_9394,N_9579);
nor UO_432 (O_432,N_9721,N_9530);
and UO_433 (O_433,N_9852,N_9981);
nor UO_434 (O_434,N_9575,N_9908);
or UO_435 (O_435,N_9493,N_9819);
nor UO_436 (O_436,N_9407,N_9142);
and UO_437 (O_437,N_9765,N_9672);
nor UO_438 (O_438,N_9361,N_9363);
or UO_439 (O_439,N_9415,N_9874);
and UO_440 (O_440,N_9007,N_9158);
nand UO_441 (O_441,N_9829,N_9408);
or UO_442 (O_442,N_9531,N_9975);
and UO_443 (O_443,N_9376,N_9469);
or UO_444 (O_444,N_9135,N_9679);
and UO_445 (O_445,N_9236,N_9300);
nor UO_446 (O_446,N_9375,N_9350);
and UO_447 (O_447,N_9736,N_9288);
nor UO_448 (O_448,N_9841,N_9659);
nor UO_449 (O_449,N_9098,N_9119);
and UO_450 (O_450,N_9177,N_9221);
nand UO_451 (O_451,N_9684,N_9925);
and UO_452 (O_452,N_9126,N_9081);
nor UO_453 (O_453,N_9910,N_9106);
and UO_454 (O_454,N_9770,N_9609);
nand UO_455 (O_455,N_9272,N_9780);
or UO_456 (O_456,N_9710,N_9507);
nor UO_457 (O_457,N_9337,N_9163);
and UO_458 (O_458,N_9105,N_9735);
xor UO_459 (O_459,N_9948,N_9776);
and UO_460 (O_460,N_9248,N_9353);
and UO_461 (O_461,N_9516,N_9617);
and UO_462 (O_462,N_9896,N_9218);
and UO_463 (O_463,N_9451,N_9593);
and UO_464 (O_464,N_9117,N_9323);
and UO_465 (O_465,N_9032,N_9470);
nor UO_466 (O_466,N_9653,N_9873);
nor UO_467 (O_467,N_9799,N_9284);
nand UO_468 (O_468,N_9000,N_9503);
or UO_469 (O_469,N_9187,N_9621);
nand UO_470 (O_470,N_9230,N_9945);
nand UO_471 (O_471,N_9108,N_9986);
nand UO_472 (O_472,N_9255,N_9294);
or UO_473 (O_473,N_9201,N_9387);
nor UO_474 (O_474,N_9649,N_9992);
nor UO_475 (O_475,N_9331,N_9327);
or UO_476 (O_476,N_9154,N_9950);
nor UO_477 (O_477,N_9476,N_9017);
or UO_478 (O_478,N_9802,N_9262);
and UO_479 (O_479,N_9985,N_9265);
nor UO_480 (O_480,N_9745,N_9197);
nand UO_481 (O_481,N_9604,N_9970);
and UO_482 (O_482,N_9374,N_9897);
and UO_483 (O_483,N_9433,N_9823);
and UO_484 (O_484,N_9812,N_9419);
nand UO_485 (O_485,N_9863,N_9092);
or UO_486 (O_486,N_9034,N_9944);
and UO_487 (O_487,N_9797,N_9611);
and UO_488 (O_488,N_9728,N_9057);
and UO_489 (O_489,N_9147,N_9587);
nor UO_490 (O_490,N_9682,N_9170);
or UO_491 (O_491,N_9420,N_9246);
and UO_492 (O_492,N_9855,N_9749);
and UO_493 (O_493,N_9685,N_9859);
nand UO_494 (O_494,N_9860,N_9958);
nor UO_495 (O_495,N_9497,N_9274);
nand UO_496 (O_496,N_9186,N_9591);
or UO_497 (O_497,N_9666,N_9762);
or UO_498 (O_498,N_9239,N_9492);
or UO_499 (O_499,N_9734,N_9051);
nand UO_500 (O_500,N_9941,N_9943);
nand UO_501 (O_501,N_9464,N_9912);
nand UO_502 (O_502,N_9184,N_9833);
and UO_503 (O_503,N_9827,N_9558);
nor UO_504 (O_504,N_9611,N_9477);
or UO_505 (O_505,N_9961,N_9768);
nand UO_506 (O_506,N_9081,N_9397);
nand UO_507 (O_507,N_9204,N_9340);
and UO_508 (O_508,N_9731,N_9945);
nor UO_509 (O_509,N_9884,N_9494);
or UO_510 (O_510,N_9868,N_9870);
nand UO_511 (O_511,N_9843,N_9596);
nor UO_512 (O_512,N_9164,N_9855);
nor UO_513 (O_513,N_9373,N_9205);
or UO_514 (O_514,N_9648,N_9165);
nor UO_515 (O_515,N_9126,N_9801);
or UO_516 (O_516,N_9879,N_9426);
nor UO_517 (O_517,N_9358,N_9612);
nand UO_518 (O_518,N_9246,N_9130);
and UO_519 (O_519,N_9035,N_9874);
nand UO_520 (O_520,N_9671,N_9908);
nand UO_521 (O_521,N_9464,N_9492);
nor UO_522 (O_522,N_9691,N_9127);
or UO_523 (O_523,N_9850,N_9777);
and UO_524 (O_524,N_9802,N_9540);
nor UO_525 (O_525,N_9429,N_9953);
nand UO_526 (O_526,N_9243,N_9026);
and UO_527 (O_527,N_9515,N_9647);
and UO_528 (O_528,N_9625,N_9177);
and UO_529 (O_529,N_9522,N_9852);
or UO_530 (O_530,N_9521,N_9353);
and UO_531 (O_531,N_9534,N_9625);
nand UO_532 (O_532,N_9799,N_9003);
nor UO_533 (O_533,N_9562,N_9825);
or UO_534 (O_534,N_9589,N_9996);
and UO_535 (O_535,N_9291,N_9844);
nand UO_536 (O_536,N_9722,N_9056);
nand UO_537 (O_537,N_9286,N_9138);
nor UO_538 (O_538,N_9353,N_9997);
nand UO_539 (O_539,N_9702,N_9447);
or UO_540 (O_540,N_9897,N_9869);
and UO_541 (O_541,N_9454,N_9058);
nand UO_542 (O_542,N_9776,N_9745);
and UO_543 (O_543,N_9055,N_9371);
nor UO_544 (O_544,N_9414,N_9921);
and UO_545 (O_545,N_9754,N_9282);
and UO_546 (O_546,N_9397,N_9022);
nor UO_547 (O_547,N_9328,N_9981);
nor UO_548 (O_548,N_9877,N_9757);
nand UO_549 (O_549,N_9004,N_9241);
nand UO_550 (O_550,N_9838,N_9473);
nor UO_551 (O_551,N_9971,N_9269);
or UO_552 (O_552,N_9107,N_9008);
nand UO_553 (O_553,N_9888,N_9246);
or UO_554 (O_554,N_9732,N_9478);
nand UO_555 (O_555,N_9083,N_9670);
or UO_556 (O_556,N_9376,N_9652);
nand UO_557 (O_557,N_9307,N_9564);
and UO_558 (O_558,N_9553,N_9037);
nor UO_559 (O_559,N_9865,N_9443);
or UO_560 (O_560,N_9936,N_9183);
nor UO_561 (O_561,N_9671,N_9495);
or UO_562 (O_562,N_9981,N_9544);
nand UO_563 (O_563,N_9237,N_9931);
nor UO_564 (O_564,N_9513,N_9319);
or UO_565 (O_565,N_9852,N_9812);
nand UO_566 (O_566,N_9324,N_9936);
nand UO_567 (O_567,N_9235,N_9704);
and UO_568 (O_568,N_9407,N_9613);
nand UO_569 (O_569,N_9074,N_9359);
nor UO_570 (O_570,N_9182,N_9712);
and UO_571 (O_571,N_9925,N_9064);
or UO_572 (O_572,N_9023,N_9582);
nand UO_573 (O_573,N_9087,N_9068);
nand UO_574 (O_574,N_9168,N_9202);
nor UO_575 (O_575,N_9143,N_9860);
and UO_576 (O_576,N_9166,N_9009);
nand UO_577 (O_577,N_9434,N_9634);
and UO_578 (O_578,N_9049,N_9600);
and UO_579 (O_579,N_9547,N_9519);
nand UO_580 (O_580,N_9158,N_9752);
nor UO_581 (O_581,N_9019,N_9812);
nor UO_582 (O_582,N_9570,N_9667);
and UO_583 (O_583,N_9483,N_9580);
and UO_584 (O_584,N_9604,N_9765);
nand UO_585 (O_585,N_9520,N_9184);
and UO_586 (O_586,N_9862,N_9599);
or UO_587 (O_587,N_9228,N_9375);
nor UO_588 (O_588,N_9632,N_9735);
or UO_589 (O_589,N_9307,N_9388);
or UO_590 (O_590,N_9291,N_9213);
xnor UO_591 (O_591,N_9838,N_9107);
and UO_592 (O_592,N_9351,N_9691);
nand UO_593 (O_593,N_9543,N_9070);
xor UO_594 (O_594,N_9021,N_9461);
or UO_595 (O_595,N_9330,N_9088);
nor UO_596 (O_596,N_9923,N_9431);
nor UO_597 (O_597,N_9651,N_9977);
xnor UO_598 (O_598,N_9917,N_9278);
nand UO_599 (O_599,N_9336,N_9754);
nand UO_600 (O_600,N_9806,N_9633);
nand UO_601 (O_601,N_9258,N_9010);
and UO_602 (O_602,N_9049,N_9892);
or UO_603 (O_603,N_9121,N_9452);
nand UO_604 (O_604,N_9845,N_9459);
nand UO_605 (O_605,N_9653,N_9004);
nand UO_606 (O_606,N_9581,N_9083);
or UO_607 (O_607,N_9603,N_9492);
nor UO_608 (O_608,N_9259,N_9129);
or UO_609 (O_609,N_9383,N_9169);
or UO_610 (O_610,N_9673,N_9031);
or UO_611 (O_611,N_9718,N_9386);
nand UO_612 (O_612,N_9596,N_9868);
nor UO_613 (O_613,N_9884,N_9794);
and UO_614 (O_614,N_9045,N_9223);
nand UO_615 (O_615,N_9649,N_9327);
and UO_616 (O_616,N_9725,N_9636);
nor UO_617 (O_617,N_9445,N_9160);
and UO_618 (O_618,N_9528,N_9431);
nor UO_619 (O_619,N_9849,N_9886);
nand UO_620 (O_620,N_9254,N_9596);
and UO_621 (O_621,N_9866,N_9759);
and UO_622 (O_622,N_9756,N_9707);
or UO_623 (O_623,N_9589,N_9965);
nand UO_624 (O_624,N_9454,N_9104);
nand UO_625 (O_625,N_9205,N_9174);
nand UO_626 (O_626,N_9295,N_9254);
or UO_627 (O_627,N_9142,N_9928);
nand UO_628 (O_628,N_9236,N_9563);
or UO_629 (O_629,N_9912,N_9106);
or UO_630 (O_630,N_9380,N_9657);
or UO_631 (O_631,N_9095,N_9413);
and UO_632 (O_632,N_9265,N_9181);
nor UO_633 (O_633,N_9150,N_9938);
or UO_634 (O_634,N_9927,N_9023);
nor UO_635 (O_635,N_9417,N_9885);
or UO_636 (O_636,N_9535,N_9433);
or UO_637 (O_637,N_9711,N_9346);
and UO_638 (O_638,N_9039,N_9443);
and UO_639 (O_639,N_9630,N_9432);
nand UO_640 (O_640,N_9861,N_9606);
nor UO_641 (O_641,N_9977,N_9174);
nor UO_642 (O_642,N_9390,N_9356);
xor UO_643 (O_643,N_9533,N_9628);
and UO_644 (O_644,N_9390,N_9406);
nand UO_645 (O_645,N_9480,N_9396);
or UO_646 (O_646,N_9631,N_9011);
and UO_647 (O_647,N_9357,N_9255);
or UO_648 (O_648,N_9304,N_9843);
and UO_649 (O_649,N_9193,N_9700);
or UO_650 (O_650,N_9646,N_9414);
nand UO_651 (O_651,N_9066,N_9477);
or UO_652 (O_652,N_9492,N_9280);
and UO_653 (O_653,N_9200,N_9493);
or UO_654 (O_654,N_9463,N_9881);
and UO_655 (O_655,N_9870,N_9931);
or UO_656 (O_656,N_9059,N_9105);
nor UO_657 (O_657,N_9708,N_9883);
nor UO_658 (O_658,N_9799,N_9640);
and UO_659 (O_659,N_9770,N_9094);
or UO_660 (O_660,N_9565,N_9636);
nand UO_661 (O_661,N_9529,N_9525);
and UO_662 (O_662,N_9889,N_9847);
nand UO_663 (O_663,N_9814,N_9184);
and UO_664 (O_664,N_9268,N_9881);
xor UO_665 (O_665,N_9990,N_9410);
or UO_666 (O_666,N_9685,N_9318);
nor UO_667 (O_667,N_9987,N_9332);
nor UO_668 (O_668,N_9996,N_9425);
or UO_669 (O_669,N_9732,N_9129);
nor UO_670 (O_670,N_9034,N_9961);
nor UO_671 (O_671,N_9132,N_9535);
and UO_672 (O_672,N_9850,N_9239);
nand UO_673 (O_673,N_9752,N_9078);
or UO_674 (O_674,N_9270,N_9263);
nand UO_675 (O_675,N_9161,N_9409);
and UO_676 (O_676,N_9709,N_9889);
and UO_677 (O_677,N_9915,N_9400);
and UO_678 (O_678,N_9253,N_9760);
or UO_679 (O_679,N_9339,N_9007);
nor UO_680 (O_680,N_9981,N_9125);
nand UO_681 (O_681,N_9141,N_9977);
nor UO_682 (O_682,N_9634,N_9223);
nor UO_683 (O_683,N_9229,N_9821);
nor UO_684 (O_684,N_9268,N_9555);
nand UO_685 (O_685,N_9310,N_9309);
or UO_686 (O_686,N_9594,N_9229);
nor UO_687 (O_687,N_9277,N_9926);
nand UO_688 (O_688,N_9507,N_9790);
nor UO_689 (O_689,N_9922,N_9569);
nor UO_690 (O_690,N_9617,N_9215);
and UO_691 (O_691,N_9763,N_9932);
or UO_692 (O_692,N_9505,N_9133);
nand UO_693 (O_693,N_9656,N_9135);
nor UO_694 (O_694,N_9176,N_9674);
nand UO_695 (O_695,N_9819,N_9616);
nand UO_696 (O_696,N_9137,N_9674);
and UO_697 (O_697,N_9509,N_9225);
and UO_698 (O_698,N_9491,N_9046);
and UO_699 (O_699,N_9986,N_9183);
nand UO_700 (O_700,N_9017,N_9722);
nor UO_701 (O_701,N_9786,N_9829);
and UO_702 (O_702,N_9084,N_9907);
or UO_703 (O_703,N_9219,N_9021);
and UO_704 (O_704,N_9588,N_9866);
nand UO_705 (O_705,N_9252,N_9644);
nand UO_706 (O_706,N_9455,N_9873);
nor UO_707 (O_707,N_9968,N_9554);
and UO_708 (O_708,N_9213,N_9490);
nand UO_709 (O_709,N_9439,N_9920);
nor UO_710 (O_710,N_9962,N_9508);
or UO_711 (O_711,N_9131,N_9652);
nor UO_712 (O_712,N_9983,N_9340);
or UO_713 (O_713,N_9410,N_9571);
and UO_714 (O_714,N_9920,N_9247);
or UO_715 (O_715,N_9476,N_9716);
or UO_716 (O_716,N_9465,N_9618);
or UO_717 (O_717,N_9266,N_9603);
nand UO_718 (O_718,N_9497,N_9151);
nor UO_719 (O_719,N_9142,N_9970);
and UO_720 (O_720,N_9756,N_9687);
nand UO_721 (O_721,N_9542,N_9260);
and UO_722 (O_722,N_9876,N_9900);
nor UO_723 (O_723,N_9189,N_9388);
nor UO_724 (O_724,N_9696,N_9102);
nor UO_725 (O_725,N_9473,N_9152);
nor UO_726 (O_726,N_9207,N_9143);
nor UO_727 (O_727,N_9057,N_9894);
nand UO_728 (O_728,N_9260,N_9818);
and UO_729 (O_729,N_9112,N_9280);
nand UO_730 (O_730,N_9780,N_9003);
nor UO_731 (O_731,N_9135,N_9303);
nor UO_732 (O_732,N_9047,N_9602);
nor UO_733 (O_733,N_9247,N_9222);
or UO_734 (O_734,N_9416,N_9218);
nor UO_735 (O_735,N_9435,N_9446);
and UO_736 (O_736,N_9525,N_9486);
or UO_737 (O_737,N_9787,N_9231);
nor UO_738 (O_738,N_9311,N_9128);
and UO_739 (O_739,N_9517,N_9408);
nor UO_740 (O_740,N_9135,N_9982);
xnor UO_741 (O_741,N_9138,N_9385);
nand UO_742 (O_742,N_9621,N_9740);
or UO_743 (O_743,N_9591,N_9311);
and UO_744 (O_744,N_9847,N_9663);
or UO_745 (O_745,N_9931,N_9327);
nor UO_746 (O_746,N_9678,N_9798);
nand UO_747 (O_747,N_9393,N_9948);
nand UO_748 (O_748,N_9903,N_9302);
and UO_749 (O_749,N_9322,N_9514);
and UO_750 (O_750,N_9711,N_9967);
or UO_751 (O_751,N_9538,N_9447);
nor UO_752 (O_752,N_9030,N_9157);
or UO_753 (O_753,N_9968,N_9321);
and UO_754 (O_754,N_9537,N_9311);
and UO_755 (O_755,N_9354,N_9516);
or UO_756 (O_756,N_9264,N_9531);
nand UO_757 (O_757,N_9360,N_9898);
and UO_758 (O_758,N_9336,N_9627);
or UO_759 (O_759,N_9794,N_9434);
nor UO_760 (O_760,N_9512,N_9374);
nand UO_761 (O_761,N_9128,N_9114);
xnor UO_762 (O_762,N_9718,N_9377);
or UO_763 (O_763,N_9530,N_9892);
or UO_764 (O_764,N_9130,N_9340);
or UO_765 (O_765,N_9308,N_9075);
nand UO_766 (O_766,N_9693,N_9725);
and UO_767 (O_767,N_9131,N_9805);
nor UO_768 (O_768,N_9893,N_9463);
and UO_769 (O_769,N_9617,N_9598);
nor UO_770 (O_770,N_9278,N_9370);
and UO_771 (O_771,N_9458,N_9766);
or UO_772 (O_772,N_9567,N_9253);
nor UO_773 (O_773,N_9192,N_9341);
xor UO_774 (O_774,N_9811,N_9810);
nand UO_775 (O_775,N_9471,N_9330);
nor UO_776 (O_776,N_9754,N_9064);
and UO_777 (O_777,N_9612,N_9950);
and UO_778 (O_778,N_9092,N_9484);
and UO_779 (O_779,N_9003,N_9006);
or UO_780 (O_780,N_9589,N_9654);
or UO_781 (O_781,N_9457,N_9435);
nand UO_782 (O_782,N_9618,N_9300);
nor UO_783 (O_783,N_9547,N_9983);
or UO_784 (O_784,N_9522,N_9979);
and UO_785 (O_785,N_9106,N_9834);
or UO_786 (O_786,N_9470,N_9637);
and UO_787 (O_787,N_9685,N_9204);
or UO_788 (O_788,N_9637,N_9815);
or UO_789 (O_789,N_9642,N_9430);
xnor UO_790 (O_790,N_9507,N_9380);
nand UO_791 (O_791,N_9253,N_9273);
and UO_792 (O_792,N_9734,N_9355);
nor UO_793 (O_793,N_9040,N_9009);
nor UO_794 (O_794,N_9671,N_9356);
nand UO_795 (O_795,N_9616,N_9788);
nor UO_796 (O_796,N_9314,N_9811);
nand UO_797 (O_797,N_9622,N_9367);
nand UO_798 (O_798,N_9708,N_9440);
nand UO_799 (O_799,N_9167,N_9540);
nand UO_800 (O_800,N_9524,N_9113);
nor UO_801 (O_801,N_9582,N_9667);
xnor UO_802 (O_802,N_9438,N_9258);
nor UO_803 (O_803,N_9375,N_9484);
or UO_804 (O_804,N_9998,N_9596);
and UO_805 (O_805,N_9405,N_9233);
nand UO_806 (O_806,N_9409,N_9266);
nand UO_807 (O_807,N_9442,N_9819);
nor UO_808 (O_808,N_9208,N_9410);
or UO_809 (O_809,N_9016,N_9008);
nor UO_810 (O_810,N_9361,N_9209);
and UO_811 (O_811,N_9492,N_9626);
nand UO_812 (O_812,N_9331,N_9599);
and UO_813 (O_813,N_9780,N_9342);
nor UO_814 (O_814,N_9931,N_9583);
nand UO_815 (O_815,N_9590,N_9163);
nor UO_816 (O_816,N_9265,N_9195);
and UO_817 (O_817,N_9386,N_9250);
nor UO_818 (O_818,N_9561,N_9337);
or UO_819 (O_819,N_9575,N_9111);
and UO_820 (O_820,N_9932,N_9128);
nand UO_821 (O_821,N_9767,N_9508);
nand UO_822 (O_822,N_9113,N_9905);
and UO_823 (O_823,N_9155,N_9420);
nor UO_824 (O_824,N_9998,N_9825);
nand UO_825 (O_825,N_9860,N_9253);
nor UO_826 (O_826,N_9356,N_9866);
nor UO_827 (O_827,N_9349,N_9012);
nor UO_828 (O_828,N_9380,N_9207);
or UO_829 (O_829,N_9229,N_9214);
nor UO_830 (O_830,N_9407,N_9670);
nand UO_831 (O_831,N_9520,N_9893);
and UO_832 (O_832,N_9979,N_9930);
nand UO_833 (O_833,N_9752,N_9657);
or UO_834 (O_834,N_9254,N_9321);
and UO_835 (O_835,N_9909,N_9426);
and UO_836 (O_836,N_9614,N_9776);
and UO_837 (O_837,N_9775,N_9587);
nand UO_838 (O_838,N_9281,N_9809);
or UO_839 (O_839,N_9971,N_9835);
nor UO_840 (O_840,N_9413,N_9167);
nor UO_841 (O_841,N_9672,N_9907);
nand UO_842 (O_842,N_9695,N_9954);
and UO_843 (O_843,N_9352,N_9776);
nand UO_844 (O_844,N_9561,N_9451);
nand UO_845 (O_845,N_9034,N_9294);
nand UO_846 (O_846,N_9029,N_9136);
or UO_847 (O_847,N_9763,N_9463);
nor UO_848 (O_848,N_9102,N_9315);
or UO_849 (O_849,N_9304,N_9730);
nor UO_850 (O_850,N_9095,N_9485);
or UO_851 (O_851,N_9857,N_9345);
or UO_852 (O_852,N_9550,N_9218);
nor UO_853 (O_853,N_9700,N_9424);
nand UO_854 (O_854,N_9736,N_9814);
nand UO_855 (O_855,N_9322,N_9165);
and UO_856 (O_856,N_9950,N_9253);
or UO_857 (O_857,N_9299,N_9149);
nor UO_858 (O_858,N_9634,N_9320);
or UO_859 (O_859,N_9980,N_9581);
and UO_860 (O_860,N_9772,N_9800);
and UO_861 (O_861,N_9152,N_9386);
or UO_862 (O_862,N_9626,N_9059);
or UO_863 (O_863,N_9450,N_9127);
or UO_864 (O_864,N_9822,N_9994);
nand UO_865 (O_865,N_9112,N_9250);
nand UO_866 (O_866,N_9546,N_9665);
nand UO_867 (O_867,N_9357,N_9410);
nor UO_868 (O_868,N_9917,N_9458);
nor UO_869 (O_869,N_9481,N_9814);
nand UO_870 (O_870,N_9781,N_9468);
and UO_871 (O_871,N_9685,N_9920);
and UO_872 (O_872,N_9783,N_9250);
nand UO_873 (O_873,N_9219,N_9274);
or UO_874 (O_874,N_9544,N_9487);
or UO_875 (O_875,N_9327,N_9014);
nor UO_876 (O_876,N_9469,N_9268);
or UO_877 (O_877,N_9444,N_9796);
and UO_878 (O_878,N_9398,N_9652);
and UO_879 (O_879,N_9429,N_9157);
or UO_880 (O_880,N_9933,N_9323);
nand UO_881 (O_881,N_9540,N_9231);
nor UO_882 (O_882,N_9459,N_9898);
and UO_883 (O_883,N_9432,N_9910);
and UO_884 (O_884,N_9182,N_9309);
nand UO_885 (O_885,N_9225,N_9042);
nor UO_886 (O_886,N_9758,N_9388);
nand UO_887 (O_887,N_9932,N_9727);
nor UO_888 (O_888,N_9222,N_9621);
or UO_889 (O_889,N_9816,N_9698);
nand UO_890 (O_890,N_9323,N_9271);
nor UO_891 (O_891,N_9942,N_9798);
or UO_892 (O_892,N_9443,N_9193);
nor UO_893 (O_893,N_9785,N_9970);
and UO_894 (O_894,N_9042,N_9308);
nor UO_895 (O_895,N_9707,N_9858);
nand UO_896 (O_896,N_9834,N_9079);
nor UO_897 (O_897,N_9054,N_9767);
nor UO_898 (O_898,N_9714,N_9409);
or UO_899 (O_899,N_9161,N_9969);
and UO_900 (O_900,N_9322,N_9097);
and UO_901 (O_901,N_9466,N_9698);
xnor UO_902 (O_902,N_9960,N_9015);
or UO_903 (O_903,N_9498,N_9930);
or UO_904 (O_904,N_9764,N_9934);
nor UO_905 (O_905,N_9523,N_9117);
and UO_906 (O_906,N_9477,N_9133);
and UO_907 (O_907,N_9833,N_9754);
and UO_908 (O_908,N_9561,N_9253);
nand UO_909 (O_909,N_9660,N_9207);
and UO_910 (O_910,N_9964,N_9362);
nor UO_911 (O_911,N_9965,N_9844);
nand UO_912 (O_912,N_9076,N_9444);
nand UO_913 (O_913,N_9852,N_9616);
and UO_914 (O_914,N_9039,N_9307);
nand UO_915 (O_915,N_9886,N_9049);
nor UO_916 (O_916,N_9207,N_9102);
and UO_917 (O_917,N_9155,N_9852);
xor UO_918 (O_918,N_9559,N_9353);
or UO_919 (O_919,N_9845,N_9227);
nor UO_920 (O_920,N_9896,N_9283);
nand UO_921 (O_921,N_9165,N_9784);
or UO_922 (O_922,N_9157,N_9897);
nor UO_923 (O_923,N_9596,N_9258);
and UO_924 (O_924,N_9340,N_9489);
or UO_925 (O_925,N_9069,N_9949);
nor UO_926 (O_926,N_9396,N_9185);
nor UO_927 (O_927,N_9125,N_9104);
and UO_928 (O_928,N_9367,N_9629);
nand UO_929 (O_929,N_9808,N_9408);
or UO_930 (O_930,N_9393,N_9336);
or UO_931 (O_931,N_9538,N_9547);
nand UO_932 (O_932,N_9098,N_9568);
and UO_933 (O_933,N_9249,N_9927);
nand UO_934 (O_934,N_9171,N_9033);
and UO_935 (O_935,N_9397,N_9487);
or UO_936 (O_936,N_9819,N_9272);
nor UO_937 (O_937,N_9749,N_9097);
or UO_938 (O_938,N_9710,N_9325);
and UO_939 (O_939,N_9309,N_9330);
xnor UO_940 (O_940,N_9008,N_9664);
nand UO_941 (O_941,N_9925,N_9250);
or UO_942 (O_942,N_9603,N_9994);
nand UO_943 (O_943,N_9283,N_9220);
nor UO_944 (O_944,N_9666,N_9483);
nor UO_945 (O_945,N_9590,N_9203);
nor UO_946 (O_946,N_9993,N_9324);
or UO_947 (O_947,N_9977,N_9906);
nor UO_948 (O_948,N_9484,N_9855);
and UO_949 (O_949,N_9071,N_9081);
nand UO_950 (O_950,N_9874,N_9818);
and UO_951 (O_951,N_9615,N_9641);
nor UO_952 (O_952,N_9944,N_9533);
or UO_953 (O_953,N_9194,N_9329);
and UO_954 (O_954,N_9761,N_9551);
nand UO_955 (O_955,N_9149,N_9669);
or UO_956 (O_956,N_9019,N_9701);
nor UO_957 (O_957,N_9477,N_9037);
or UO_958 (O_958,N_9553,N_9235);
and UO_959 (O_959,N_9132,N_9686);
nor UO_960 (O_960,N_9766,N_9189);
nor UO_961 (O_961,N_9082,N_9208);
and UO_962 (O_962,N_9292,N_9960);
nand UO_963 (O_963,N_9493,N_9240);
or UO_964 (O_964,N_9602,N_9787);
nor UO_965 (O_965,N_9381,N_9485);
or UO_966 (O_966,N_9784,N_9128);
and UO_967 (O_967,N_9489,N_9294);
or UO_968 (O_968,N_9663,N_9397);
and UO_969 (O_969,N_9348,N_9880);
nor UO_970 (O_970,N_9065,N_9056);
nand UO_971 (O_971,N_9962,N_9973);
nand UO_972 (O_972,N_9255,N_9920);
and UO_973 (O_973,N_9243,N_9506);
nand UO_974 (O_974,N_9621,N_9612);
nand UO_975 (O_975,N_9585,N_9222);
and UO_976 (O_976,N_9693,N_9407);
nor UO_977 (O_977,N_9864,N_9277);
nor UO_978 (O_978,N_9339,N_9329);
nand UO_979 (O_979,N_9614,N_9100);
or UO_980 (O_980,N_9235,N_9857);
and UO_981 (O_981,N_9866,N_9154);
and UO_982 (O_982,N_9616,N_9761);
nor UO_983 (O_983,N_9126,N_9787);
nor UO_984 (O_984,N_9424,N_9766);
nor UO_985 (O_985,N_9789,N_9827);
and UO_986 (O_986,N_9227,N_9217);
and UO_987 (O_987,N_9689,N_9948);
nor UO_988 (O_988,N_9169,N_9752);
nor UO_989 (O_989,N_9951,N_9482);
nor UO_990 (O_990,N_9886,N_9702);
nor UO_991 (O_991,N_9420,N_9429);
or UO_992 (O_992,N_9703,N_9011);
nor UO_993 (O_993,N_9513,N_9748);
or UO_994 (O_994,N_9494,N_9918);
nand UO_995 (O_995,N_9430,N_9169);
and UO_996 (O_996,N_9144,N_9137);
or UO_997 (O_997,N_9030,N_9847);
nor UO_998 (O_998,N_9014,N_9411);
and UO_999 (O_999,N_9155,N_9601);
or UO_1000 (O_1000,N_9106,N_9460);
nand UO_1001 (O_1001,N_9067,N_9558);
or UO_1002 (O_1002,N_9944,N_9727);
or UO_1003 (O_1003,N_9459,N_9789);
and UO_1004 (O_1004,N_9874,N_9366);
nor UO_1005 (O_1005,N_9005,N_9406);
or UO_1006 (O_1006,N_9160,N_9006);
and UO_1007 (O_1007,N_9582,N_9274);
nor UO_1008 (O_1008,N_9757,N_9573);
nand UO_1009 (O_1009,N_9996,N_9722);
nand UO_1010 (O_1010,N_9907,N_9823);
nand UO_1011 (O_1011,N_9729,N_9891);
or UO_1012 (O_1012,N_9203,N_9810);
nand UO_1013 (O_1013,N_9434,N_9158);
nor UO_1014 (O_1014,N_9380,N_9286);
nand UO_1015 (O_1015,N_9811,N_9019);
or UO_1016 (O_1016,N_9209,N_9782);
or UO_1017 (O_1017,N_9616,N_9158);
and UO_1018 (O_1018,N_9057,N_9948);
and UO_1019 (O_1019,N_9350,N_9971);
and UO_1020 (O_1020,N_9427,N_9851);
or UO_1021 (O_1021,N_9136,N_9893);
or UO_1022 (O_1022,N_9877,N_9334);
nor UO_1023 (O_1023,N_9849,N_9763);
or UO_1024 (O_1024,N_9987,N_9881);
nand UO_1025 (O_1025,N_9412,N_9195);
nor UO_1026 (O_1026,N_9914,N_9848);
nand UO_1027 (O_1027,N_9920,N_9906);
nor UO_1028 (O_1028,N_9665,N_9317);
and UO_1029 (O_1029,N_9756,N_9086);
nand UO_1030 (O_1030,N_9024,N_9359);
and UO_1031 (O_1031,N_9453,N_9144);
or UO_1032 (O_1032,N_9925,N_9714);
or UO_1033 (O_1033,N_9308,N_9945);
nand UO_1034 (O_1034,N_9393,N_9837);
nor UO_1035 (O_1035,N_9730,N_9423);
nor UO_1036 (O_1036,N_9079,N_9202);
nand UO_1037 (O_1037,N_9075,N_9905);
and UO_1038 (O_1038,N_9218,N_9608);
nor UO_1039 (O_1039,N_9551,N_9288);
or UO_1040 (O_1040,N_9195,N_9105);
and UO_1041 (O_1041,N_9623,N_9571);
or UO_1042 (O_1042,N_9118,N_9179);
or UO_1043 (O_1043,N_9433,N_9432);
nand UO_1044 (O_1044,N_9734,N_9494);
nor UO_1045 (O_1045,N_9309,N_9467);
or UO_1046 (O_1046,N_9838,N_9318);
nor UO_1047 (O_1047,N_9581,N_9280);
nand UO_1048 (O_1048,N_9226,N_9045);
or UO_1049 (O_1049,N_9467,N_9990);
nor UO_1050 (O_1050,N_9959,N_9883);
and UO_1051 (O_1051,N_9871,N_9139);
nor UO_1052 (O_1052,N_9778,N_9688);
and UO_1053 (O_1053,N_9540,N_9514);
or UO_1054 (O_1054,N_9029,N_9293);
and UO_1055 (O_1055,N_9588,N_9181);
and UO_1056 (O_1056,N_9034,N_9627);
nand UO_1057 (O_1057,N_9825,N_9560);
or UO_1058 (O_1058,N_9641,N_9601);
nand UO_1059 (O_1059,N_9974,N_9295);
or UO_1060 (O_1060,N_9898,N_9316);
nor UO_1061 (O_1061,N_9959,N_9985);
nand UO_1062 (O_1062,N_9232,N_9327);
nor UO_1063 (O_1063,N_9851,N_9901);
nor UO_1064 (O_1064,N_9561,N_9087);
nand UO_1065 (O_1065,N_9788,N_9359);
nor UO_1066 (O_1066,N_9242,N_9135);
nand UO_1067 (O_1067,N_9509,N_9142);
or UO_1068 (O_1068,N_9686,N_9371);
or UO_1069 (O_1069,N_9284,N_9545);
nand UO_1070 (O_1070,N_9749,N_9447);
xnor UO_1071 (O_1071,N_9382,N_9373);
and UO_1072 (O_1072,N_9784,N_9493);
nor UO_1073 (O_1073,N_9225,N_9671);
nand UO_1074 (O_1074,N_9506,N_9075);
nor UO_1075 (O_1075,N_9003,N_9101);
or UO_1076 (O_1076,N_9997,N_9116);
or UO_1077 (O_1077,N_9440,N_9469);
and UO_1078 (O_1078,N_9684,N_9001);
nand UO_1079 (O_1079,N_9274,N_9981);
nor UO_1080 (O_1080,N_9201,N_9223);
and UO_1081 (O_1081,N_9520,N_9272);
nand UO_1082 (O_1082,N_9643,N_9320);
nand UO_1083 (O_1083,N_9742,N_9781);
or UO_1084 (O_1084,N_9617,N_9489);
or UO_1085 (O_1085,N_9684,N_9885);
nand UO_1086 (O_1086,N_9473,N_9327);
nand UO_1087 (O_1087,N_9617,N_9025);
nand UO_1088 (O_1088,N_9370,N_9584);
nand UO_1089 (O_1089,N_9622,N_9915);
nand UO_1090 (O_1090,N_9961,N_9170);
and UO_1091 (O_1091,N_9619,N_9267);
and UO_1092 (O_1092,N_9366,N_9834);
or UO_1093 (O_1093,N_9104,N_9862);
or UO_1094 (O_1094,N_9991,N_9852);
nor UO_1095 (O_1095,N_9429,N_9050);
and UO_1096 (O_1096,N_9908,N_9244);
or UO_1097 (O_1097,N_9801,N_9500);
xor UO_1098 (O_1098,N_9388,N_9882);
nand UO_1099 (O_1099,N_9273,N_9604);
or UO_1100 (O_1100,N_9950,N_9309);
and UO_1101 (O_1101,N_9025,N_9334);
or UO_1102 (O_1102,N_9691,N_9697);
and UO_1103 (O_1103,N_9788,N_9249);
nor UO_1104 (O_1104,N_9540,N_9292);
and UO_1105 (O_1105,N_9692,N_9807);
and UO_1106 (O_1106,N_9536,N_9780);
nand UO_1107 (O_1107,N_9897,N_9560);
or UO_1108 (O_1108,N_9057,N_9613);
nand UO_1109 (O_1109,N_9298,N_9074);
nand UO_1110 (O_1110,N_9023,N_9430);
nor UO_1111 (O_1111,N_9239,N_9306);
nand UO_1112 (O_1112,N_9135,N_9298);
or UO_1113 (O_1113,N_9074,N_9583);
nand UO_1114 (O_1114,N_9460,N_9787);
nand UO_1115 (O_1115,N_9899,N_9869);
nor UO_1116 (O_1116,N_9720,N_9980);
and UO_1117 (O_1117,N_9922,N_9494);
nor UO_1118 (O_1118,N_9980,N_9604);
or UO_1119 (O_1119,N_9078,N_9781);
and UO_1120 (O_1120,N_9979,N_9603);
or UO_1121 (O_1121,N_9229,N_9121);
nand UO_1122 (O_1122,N_9445,N_9465);
nor UO_1123 (O_1123,N_9499,N_9403);
nand UO_1124 (O_1124,N_9271,N_9179);
nand UO_1125 (O_1125,N_9938,N_9899);
nand UO_1126 (O_1126,N_9100,N_9844);
nand UO_1127 (O_1127,N_9792,N_9913);
and UO_1128 (O_1128,N_9678,N_9447);
or UO_1129 (O_1129,N_9602,N_9794);
nor UO_1130 (O_1130,N_9851,N_9888);
nor UO_1131 (O_1131,N_9914,N_9466);
or UO_1132 (O_1132,N_9298,N_9005);
or UO_1133 (O_1133,N_9657,N_9225);
nor UO_1134 (O_1134,N_9731,N_9794);
or UO_1135 (O_1135,N_9064,N_9538);
nand UO_1136 (O_1136,N_9966,N_9012);
nand UO_1137 (O_1137,N_9737,N_9665);
nor UO_1138 (O_1138,N_9237,N_9536);
and UO_1139 (O_1139,N_9699,N_9567);
and UO_1140 (O_1140,N_9162,N_9998);
and UO_1141 (O_1141,N_9387,N_9606);
or UO_1142 (O_1142,N_9280,N_9337);
nand UO_1143 (O_1143,N_9551,N_9337);
nor UO_1144 (O_1144,N_9261,N_9322);
and UO_1145 (O_1145,N_9593,N_9948);
or UO_1146 (O_1146,N_9833,N_9166);
or UO_1147 (O_1147,N_9583,N_9907);
and UO_1148 (O_1148,N_9149,N_9613);
and UO_1149 (O_1149,N_9361,N_9175);
nor UO_1150 (O_1150,N_9255,N_9435);
and UO_1151 (O_1151,N_9657,N_9125);
nor UO_1152 (O_1152,N_9614,N_9660);
or UO_1153 (O_1153,N_9154,N_9256);
nor UO_1154 (O_1154,N_9811,N_9610);
xor UO_1155 (O_1155,N_9832,N_9668);
and UO_1156 (O_1156,N_9680,N_9118);
and UO_1157 (O_1157,N_9039,N_9880);
nand UO_1158 (O_1158,N_9433,N_9097);
or UO_1159 (O_1159,N_9447,N_9505);
and UO_1160 (O_1160,N_9689,N_9772);
nor UO_1161 (O_1161,N_9660,N_9243);
or UO_1162 (O_1162,N_9379,N_9993);
and UO_1163 (O_1163,N_9188,N_9187);
or UO_1164 (O_1164,N_9908,N_9590);
nor UO_1165 (O_1165,N_9379,N_9671);
nand UO_1166 (O_1166,N_9917,N_9753);
and UO_1167 (O_1167,N_9082,N_9960);
nor UO_1168 (O_1168,N_9351,N_9674);
nor UO_1169 (O_1169,N_9559,N_9855);
or UO_1170 (O_1170,N_9995,N_9607);
and UO_1171 (O_1171,N_9377,N_9908);
nor UO_1172 (O_1172,N_9748,N_9727);
nor UO_1173 (O_1173,N_9528,N_9209);
and UO_1174 (O_1174,N_9290,N_9269);
and UO_1175 (O_1175,N_9281,N_9842);
and UO_1176 (O_1176,N_9190,N_9687);
and UO_1177 (O_1177,N_9067,N_9930);
and UO_1178 (O_1178,N_9835,N_9074);
and UO_1179 (O_1179,N_9918,N_9515);
or UO_1180 (O_1180,N_9261,N_9731);
nand UO_1181 (O_1181,N_9533,N_9897);
nand UO_1182 (O_1182,N_9267,N_9048);
nand UO_1183 (O_1183,N_9549,N_9565);
or UO_1184 (O_1184,N_9150,N_9656);
and UO_1185 (O_1185,N_9880,N_9853);
and UO_1186 (O_1186,N_9235,N_9201);
and UO_1187 (O_1187,N_9133,N_9955);
and UO_1188 (O_1188,N_9043,N_9842);
nand UO_1189 (O_1189,N_9455,N_9832);
nand UO_1190 (O_1190,N_9104,N_9393);
nand UO_1191 (O_1191,N_9296,N_9261);
and UO_1192 (O_1192,N_9547,N_9498);
and UO_1193 (O_1193,N_9568,N_9244);
and UO_1194 (O_1194,N_9942,N_9817);
or UO_1195 (O_1195,N_9468,N_9455);
and UO_1196 (O_1196,N_9831,N_9372);
and UO_1197 (O_1197,N_9931,N_9057);
nand UO_1198 (O_1198,N_9444,N_9877);
nand UO_1199 (O_1199,N_9262,N_9883);
nand UO_1200 (O_1200,N_9905,N_9300);
nand UO_1201 (O_1201,N_9419,N_9937);
and UO_1202 (O_1202,N_9207,N_9448);
or UO_1203 (O_1203,N_9137,N_9789);
and UO_1204 (O_1204,N_9598,N_9729);
and UO_1205 (O_1205,N_9345,N_9205);
nand UO_1206 (O_1206,N_9469,N_9255);
xor UO_1207 (O_1207,N_9079,N_9855);
nor UO_1208 (O_1208,N_9006,N_9873);
nand UO_1209 (O_1209,N_9039,N_9328);
nand UO_1210 (O_1210,N_9939,N_9222);
nor UO_1211 (O_1211,N_9950,N_9090);
nor UO_1212 (O_1212,N_9854,N_9890);
or UO_1213 (O_1213,N_9357,N_9331);
nor UO_1214 (O_1214,N_9380,N_9075);
nor UO_1215 (O_1215,N_9662,N_9220);
nor UO_1216 (O_1216,N_9461,N_9785);
nor UO_1217 (O_1217,N_9716,N_9090);
and UO_1218 (O_1218,N_9198,N_9234);
and UO_1219 (O_1219,N_9705,N_9768);
nand UO_1220 (O_1220,N_9655,N_9399);
nor UO_1221 (O_1221,N_9573,N_9991);
nand UO_1222 (O_1222,N_9862,N_9866);
nand UO_1223 (O_1223,N_9710,N_9458);
nor UO_1224 (O_1224,N_9171,N_9662);
or UO_1225 (O_1225,N_9171,N_9184);
nor UO_1226 (O_1226,N_9910,N_9483);
or UO_1227 (O_1227,N_9100,N_9914);
nand UO_1228 (O_1228,N_9356,N_9167);
and UO_1229 (O_1229,N_9385,N_9563);
and UO_1230 (O_1230,N_9399,N_9268);
nor UO_1231 (O_1231,N_9148,N_9776);
nor UO_1232 (O_1232,N_9171,N_9611);
or UO_1233 (O_1233,N_9341,N_9272);
nand UO_1234 (O_1234,N_9202,N_9508);
or UO_1235 (O_1235,N_9299,N_9914);
and UO_1236 (O_1236,N_9977,N_9525);
nand UO_1237 (O_1237,N_9689,N_9654);
nand UO_1238 (O_1238,N_9908,N_9444);
nor UO_1239 (O_1239,N_9290,N_9042);
nand UO_1240 (O_1240,N_9581,N_9547);
and UO_1241 (O_1241,N_9491,N_9445);
nand UO_1242 (O_1242,N_9534,N_9138);
nand UO_1243 (O_1243,N_9020,N_9612);
xor UO_1244 (O_1244,N_9438,N_9182);
and UO_1245 (O_1245,N_9514,N_9790);
and UO_1246 (O_1246,N_9079,N_9611);
and UO_1247 (O_1247,N_9355,N_9923);
and UO_1248 (O_1248,N_9236,N_9985);
and UO_1249 (O_1249,N_9288,N_9682);
and UO_1250 (O_1250,N_9805,N_9451);
or UO_1251 (O_1251,N_9078,N_9832);
nand UO_1252 (O_1252,N_9808,N_9897);
and UO_1253 (O_1253,N_9385,N_9426);
nor UO_1254 (O_1254,N_9490,N_9635);
and UO_1255 (O_1255,N_9511,N_9287);
or UO_1256 (O_1256,N_9924,N_9876);
nor UO_1257 (O_1257,N_9906,N_9069);
nand UO_1258 (O_1258,N_9696,N_9596);
nand UO_1259 (O_1259,N_9471,N_9420);
nand UO_1260 (O_1260,N_9608,N_9996);
and UO_1261 (O_1261,N_9306,N_9273);
and UO_1262 (O_1262,N_9576,N_9464);
nor UO_1263 (O_1263,N_9146,N_9233);
nand UO_1264 (O_1264,N_9748,N_9930);
nor UO_1265 (O_1265,N_9229,N_9857);
and UO_1266 (O_1266,N_9076,N_9366);
nand UO_1267 (O_1267,N_9993,N_9744);
nor UO_1268 (O_1268,N_9747,N_9521);
nor UO_1269 (O_1269,N_9232,N_9044);
and UO_1270 (O_1270,N_9646,N_9825);
or UO_1271 (O_1271,N_9132,N_9773);
nand UO_1272 (O_1272,N_9479,N_9304);
and UO_1273 (O_1273,N_9497,N_9604);
or UO_1274 (O_1274,N_9966,N_9354);
nor UO_1275 (O_1275,N_9740,N_9618);
and UO_1276 (O_1276,N_9707,N_9940);
or UO_1277 (O_1277,N_9000,N_9098);
or UO_1278 (O_1278,N_9990,N_9873);
or UO_1279 (O_1279,N_9395,N_9763);
and UO_1280 (O_1280,N_9815,N_9102);
nand UO_1281 (O_1281,N_9946,N_9193);
or UO_1282 (O_1282,N_9016,N_9329);
or UO_1283 (O_1283,N_9645,N_9298);
or UO_1284 (O_1284,N_9288,N_9665);
and UO_1285 (O_1285,N_9234,N_9998);
nand UO_1286 (O_1286,N_9796,N_9522);
and UO_1287 (O_1287,N_9732,N_9034);
or UO_1288 (O_1288,N_9276,N_9997);
nand UO_1289 (O_1289,N_9223,N_9549);
or UO_1290 (O_1290,N_9555,N_9745);
nand UO_1291 (O_1291,N_9586,N_9057);
or UO_1292 (O_1292,N_9355,N_9198);
and UO_1293 (O_1293,N_9418,N_9916);
nor UO_1294 (O_1294,N_9364,N_9530);
nand UO_1295 (O_1295,N_9193,N_9799);
or UO_1296 (O_1296,N_9681,N_9262);
nand UO_1297 (O_1297,N_9903,N_9657);
nor UO_1298 (O_1298,N_9790,N_9142);
or UO_1299 (O_1299,N_9291,N_9055);
and UO_1300 (O_1300,N_9791,N_9339);
nand UO_1301 (O_1301,N_9049,N_9154);
nand UO_1302 (O_1302,N_9096,N_9467);
and UO_1303 (O_1303,N_9443,N_9678);
nor UO_1304 (O_1304,N_9237,N_9533);
and UO_1305 (O_1305,N_9006,N_9263);
or UO_1306 (O_1306,N_9419,N_9166);
and UO_1307 (O_1307,N_9259,N_9405);
nand UO_1308 (O_1308,N_9970,N_9164);
nand UO_1309 (O_1309,N_9687,N_9567);
or UO_1310 (O_1310,N_9071,N_9019);
nand UO_1311 (O_1311,N_9923,N_9185);
nand UO_1312 (O_1312,N_9680,N_9621);
or UO_1313 (O_1313,N_9865,N_9223);
nor UO_1314 (O_1314,N_9221,N_9215);
nand UO_1315 (O_1315,N_9828,N_9015);
nor UO_1316 (O_1316,N_9027,N_9004);
and UO_1317 (O_1317,N_9003,N_9017);
and UO_1318 (O_1318,N_9294,N_9044);
or UO_1319 (O_1319,N_9466,N_9284);
or UO_1320 (O_1320,N_9282,N_9610);
or UO_1321 (O_1321,N_9357,N_9007);
nor UO_1322 (O_1322,N_9081,N_9989);
or UO_1323 (O_1323,N_9559,N_9130);
or UO_1324 (O_1324,N_9405,N_9295);
and UO_1325 (O_1325,N_9401,N_9736);
and UO_1326 (O_1326,N_9605,N_9556);
or UO_1327 (O_1327,N_9738,N_9055);
or UO_1328 (O_1328,N_9013,N_9479);
nand UO_1329 (O_1329,N_9597,N_9804);
and UO_1330 (O_1330,N_9320,N_9283);
or UO_1331 (O_1331,N_9027,N_9715);
nand UO_1332 (O_1332,N_9614,N_9287);
nand UO_1333 (O_1333,N_9793,N_9185);
nand UO_1334 (O_1334,N_9614,N_9003);
nor UO_1335 (O_1335,N_9775,N_9608);
nor UO_1336 (O_1336,N_9220,N_9688);
and UO_1337 (O_1337,N_9323,N_9721);
and UO_1338 (O_1338,N_9644,N_9710);
or UO_1339 (O_1339,N_9525,N_9112);
or UO_1340 (O_1340,N_9198,N_9330);
nor UO_1341 (O_1341,N_9773,N_9312);
nor UO_1342 (O_1342,N_9696,N_9006);
or UO_1343 (O_1343,N_9482,N_9682);
nand UO_1344 (O_1344,N_9316,N_9784);
nor UO_1345 (O_1345,N_9916,N_9583);
or UO_1346 (O_1346,N_9490,N_9857);
and UO_1347 (O_1347,N_9467,N_9868);
xnor UO_1348 (O_1348,N_9936,N_9579);
and UO_1349 (O_1349,N_9387,N_9117);
nand UO_1350 (O_1350,N_9965,N_9259);
and UO_1351 (O_1351,N_9546,N_9928);
and UO_1352 (O_1352,N_9999,N_9782);
nor UO_1353 (O_1353,N_9125,N_9182);
and UO_1354 (O_1354,N_9486,N_9687);
and UO_1355 (O_1355,N_9500,N_9856);
nand UO_1356 (O_1356,N_9346,N_9106);
or UO_1357 (O_1357,N_9545,N_9731);
and UO_1358 (O_1358,N_9845,N_9454);
xor UO_1359 (O_1359,N_9626,N_9771);
nor UO_1360 (O_1360,N_9114,N_9181);
or UO_1361 (O_1361,N_9368,N_9733);
or UO_1362 (O_1362,N_9587,N_9966);
or UO_1363 (O_1363,N_9239,N_9923);
and UO_1364 (O_1364,N_9207,N_9671);
nand UO_1365 (O_1365,N_9535,N_9502);
or UO_1366 (O_1366,N_9523,N_9707);
nor UO_1367 (O_1367,N_9350,N_9031);
nor UO_1368 (O_1368,N_9138,N_9773);
nor UO_1369 (O_1369,N_9069,N_9443);
xnor UO_1370 (O_1370,N_9923,N_9836);
nand UO_1371 (O_1371,N_9653,N_9131);
or UO_1372 (O_1372,N_9060,N_9766);
nand UO_1373 (O_1373,N_9069,N_9551);
or UO_1374 (O_1374,N_9205,N_9997);
nor UO_1375 (O_1375,N_9496,N_9786);
nand UO_1376 (O_1376,N_9065,N_9089);
or UO_1377 (O_1377,N_9012,N_9493);
nand UO_1378 (O_1378,N_9993,N_9533);
nand UO_1379 (O_1379,N_9830,N_9048);
and UO_1380 (O_1380,N_9973,N_9637);
or UO_1381 (O_1381,N_9868,N_9890);
and UO_1382 (O_1382,N_9321,N_9414);
nor UO_1383 (O_1383,N_9296,N_9943);
nand UO_1384 (O_1384,N_9470,N_9407);
and UO_1385 (O_1385,N_9861,N_9097);
xnor UO_1386 (O_1386,N_9569,N_9196);
nand UO_1387 (O_1387,N_9372,N_9397);
nor UO_1388 (O_1388,N_9995,N_9745);
nor UO_1389 (O_1389,N_9272,N_9176);
and UO_1390 (O_1390,N_9549,N_9061);
xnor UO_1391 (O_1391,N_9977,N_9928);
and UO_1392 (O_1392,N_9467,N_9106);
and UO_1393 (O_1393,N_9318,N_9308);
and UO_1394 (O_1394,N_9187,N_9082);
and UO_1395 (O_1395,N_9694,N_9365);
or UO_1396 (O_1396,N_9663,N_9518);
nand UO_1397 (O_1397,N_9430,N_9065);
nand UO_1398 (O_1398,N_9846,N_9633);
and UO_1399 (O_1399,N_9264,N_9011);
and UO_1400 (O_1400,N_9644,N_9393);
and UO_1401 (O_1401,N_9531,N_9820);
or UO_1402 (O_1402,N_9874,N_9780);
or UO_1403 (O_1403,N_9313,N_9648);
or UO_1404 (O_1404,N_9309,N_9371);
or UO_1405 (O_1405,N_9397,N_9473);
xor UO_1406 (O_1406,N_9185,N_9970);
nor UO_1407 (O_1407,N_9136,N_9299);
and UO_1408 (O_1408,N_9305,N_9137);
and UO_1409 (O_1409,N_9217,N_9254);
nand UO_1410 (O_1410,N_9262,N_9453);
or UO_1411 (O_1411,N_9880,N_9548);
nor UO_1412 (O_1412,N_9309,N_9733);
nand UO_1413 (O_1413,N_9388,N_9527);
and UO_1414 (O_1414,N_9177,N_9544);
nand UO_1415 (O_1415,N_9920,N_9246);
nor UO_1416 (O_1416,N_9111,N_9237);
nand UO_1417 (O_1417,N_9351,N_9865);
nand UO_1418 (O_1418,N_9716,N_9739);
nand UO_1419 (O_1419,N_9723,N_9825);
nor UO_1420 (O_1420,N_9759,N_9394);
nor UO_1421 (O_1421,N_9726,N_9681);
or UO_1422 (O_1422,N_9509,N_9373);
or UO_1423 (O_1423,N_9002,N_9024);
and UO_1424 (O_1424,N_9706,N_9907);
nor UO_1425 (O_1425,N_9635,N_9452);
or UO_1426 (O_1426,N_9149,N_9576);
nor UO_1427 (O_1427,N_9533,N_9185);
nand UO_1428 (O_1428,N_9039,N_9839);
nor UO_1429 (O_1429,N_9236,N_9910);
nand UO_1430 (O_1430,N_9112,N_9168);
or UO_1431 (O_1431,N_9193,N_9559);
and UO_1432 (O_1432,N_9487,N_9192);
nand UO_1433 (O_1433,N_9648,N_9869);
and UO_1434 (O_1434,N_9819,N_9422);
and UO_1435 (O_1435,N_9862,N_9392);
nor UO_1436 (O_1436,N_9378,N_9537);
nand UO_1437 (O_1437,N_9644,N_9284);
nand UO_1438 (O_1438,N_9455,N_9826);
nor UO_1439 (O_1439,N_9696,N_9476);
or UO_1440 (O_1440,N_9514,N_9912);
or UO_1441 (O_1441,N_9391,N_9030);
nor UO_1442 (O_1442,N_9661,N_9975);
or UO_1443 (O_1443,N_9089,N_9801);
nand UO_1444 (O_1444,N_9706,N_9152);
nor UO_1445 (O_1445,N_9413,N_9504);
and UO_1446 (O_1446,N_9744,N_9638);
nor UO_1447 (O_1447,N_9354,N_9375);
or UO_1448 (O_1448,N_9793,N_9134);
nor UO_1449 (O_1449,N_9436,N_9177);
nand UO_1450 (O_1450,N_9896,N_9579);
nand UO_1451 (O_1451,N_9214,N_9244);
nand UO_1452 (O_1452,N_9644,N_9122);
or UO_1453 (O_1453,N_9641,N_9418);
and UO_1454 (O_1454,N_9930,N_9687);
nor UO_1455 (O_1455,N_9727,N_9097);
or UO_1456 (O_1456,N_9313,N_9600);
nor UO_1457 (O_1457,N_9217,N_9073);
or UO_1458 (O_1458,N_9831,N_9345);
nor UO_1459 (O_1459,N_9397,N_9365);
and UO_1460 (O_1460,N_9037,N_9824);
and UO_1461 (O_1461,N_9076,N_9126);
or UO_1462 (O_1462,N_9555,N_9244);
nand UO_1463 (O_1463,N_9844,N_9927);
nor UO_1464 (O_1464,N_9380,N_9026);
nor UO_1465 (O_1465,N_9029,N_9668);
and UO_1466 (O_1466,N_9803,N_9710);
xnor UO_1467 (O_1467,N_9305,N_9041);
and UO_1468 (O_1468,N_9735,N_9788);
and UO_1469 (O_1469,N_9802,N_9386);
and UO_1470 (O_1470,N_9544,N_9939);
or UO_1471 (O_1471,N_9859,N_9203);
nor UO_1472 (O_1472,N_9153,N_9140);
or UO_1473 (O_1473,N_9394,N_9855);
nand UO_1474 (O_1474,N_9767,N_9305);
nor UO_1475 (O_1475,N_9069,N_9139);
or UO_1476 (O_1476,N_9726,N_9714);
and UO_1477 (O_1477,N_9922,N_9860);
or UO_1478 (O_1478,N_9126,N_9283);
or UO_1479 (O_1479,N_9177,N_9375);
or UO_1480 (O_1480,N_9906,N_9497);
or UO_1481 (O_1481,N_9837,N_9494);
or UO_1482 (O_1482,N_9981,N_9880);
and UO_1483 (O_1483,N_9497,N_9336);
nor UO_1484 (O_1484,N_9025,N_9378);
nor UO_1485 (O_1485,N_9616,N_9824);
nand UO_1486 (O_1486,N_9045,N_9584);
and UO_1487 (O_1487,N_9454,N_9884);
and UO_1488 (O_1488,N_9180,N_9896);
and UO_1489 (O_1489,N_9794,N_9741);
nand UO_1490 (O_1490,N_9294,N_9041);
nor UO_1491 (O_1491,N_9177,N_9927);
or UO_1492 (O_1492,N_9933,N_9265);
nand UO_1493 (O_1493,N_9354,N_9190);
nor UO_1494 (O_1494,N_9906,N_9988);
nand UO_1495 (O_1495,N_9633,N_9258);
and UO_1496 (O_1496,N_9811,N_9926);
or UO_1497 (O_1497,N_9338,N_9293);
nand UO_1498 (O_1498,N_9571,N_9025);
nand UO_1499 (O_1499,N_9361,N_9638);
endmodule