module basic_500_3000_500_3_levels_2xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_484,In_40);
nand U1 (N_1,In_238,In_355);
nor U2 (N_2,In_281,In_30);
and U3 (N_3,In_322,In_331);
nand U4 (N_4,In_323,In_224);
and U5 (N_5,In_488,In_382);
and U6 (N_6,In_92,In_339);
and U7 (N_7,In_466,In_36);
or U8 (N_8,In_402,In_259);
nor U9 (N_9,In_385,In_395);
or U10 (N_10,In_473,In_441);
nor U11 (N_11,In_452,In_279);
or U12 (N_12,In_325,In_405);
and U13 (N_13,In_34,In_438);
or U14 (N_14,In_100,In_164);
or U15 (N_15,In_67,In_13);
nand U16 (N_16,In_18,In_23);
or U17 (N_17,In_123,In_108);
or U18 (N_18,In_449,In_235);
and U19 (N_19,In_494,In_283);
nand U20 (N_20,In_115,In_455);
and U21 (N_21,In_477,In_76);
or U22 (N_22,In_421,In_304);
nor U23 (N_23,In_75,In_432);
xnor U24 (N_24,In_270,In_167);
nand U25 (N_25,In_327,In_109);
xor U26 (N_26,In_51,In_110);
or U27 (N_27,In_362,In_89);
nand U28 (N_28,In_263,In_423);
or U29 (N_29,In_275,In_20);
nand U30 (N_30,In_282,In_239);
and U31 (N_31,In_185,In_15);
nand U32 (N_32,In_461,In_3);
nor U33 (N_33,In_414,In_476);
and U34 (N_34,In_433,In_314);
and U35 (N_35,In_78,In_94);
or U36 (N_36,In_457,In_493);
nand U37 (N_37,In_435,In_284);
or U38 (N_38,In_199,In_212);
and U39 (N_39,In_141,In_374);
or U40 (N_40,In_128,In_230);
nand U41 (N_41,In_243,In_93);
or U42 (N_42,In_286,In_328);
and U43 (N_43,In_17,In_114);
or U44 (N_44,In_448,In_379);
nor U45 (N_45,In_383,In_111);
and U46 (N_46,In_166,In_474);
nand U47 (N_47,In_258,In_136);
nand U48 (N_48,In_104,In_124);
or U49 (N_49,In_27,In_491);
and U50 (N_50,In_344,In_320);
nor U51 (N_51,In_338,In_264);
and U52 (N_52,In_132,In_160);
nand U53 (N_53,In_41,In_209);
and U54 (N_54,In_498,In_143);
nor U55 (N_55,In_139,In_192);
nor U56 (N_56,In_80,In_214);
nor U57 (N_57,In_392,In_145);
nand U58 (N_58,In_483,In_161);
or U59 (N_59,In_496,In_237);
nor U60 (N_60,In_463,In_172);
and U61 (N_61,In_266,In_39);
nor U62 (N_62,In_241,In_408);
nand U63 (N_63,In_45,In_419);
nor U64 (N_64,In_44,In_208);
nand U65 (N_65,In_245,In_1);
nor U66 (N_66,In_31,In_256);
nand U67 (N_67,In_2,In_200);
and U68 (N_68,In_358,In_142);
and U69 (N_69,In_203,In_156);
nor U70 (N_70,In_271,In_194);
nand U71 (N_71,In_404,In_61);
or U72 (N_72,In_380,In_64);
and U73 (N_73,In_240,In_345);
or U74 (N_74,In_425,In_267);
nand U75 (N_75,In_190,In_497);
or U76 (N_76,In_84,In_375);
and U77 (N_77,In_295,In_117);
nor U78 (N_78,In_417,In_310);
or U79 (N_79,In_318,In_9);
and U80 (N_80,In_426,In_356);
and U81 (N_81,In_289,In_377);
nand U82 (N_82,In_430,In_303);
or U83 (N_83,In_407,In_361);
and U84 (N_84,In_149,In_350);
nand U85 (N_85,In_324,In_119);
and U86 (N_86,In_72,In_416);
nand U87 (N_87,In_229,In_255);
nor U88 (N_88,In_305,In_35);
or U89 (N_89,In_265,In_85);
xor U90 (N_90,In_151,In_225);
nor U91 (N_91,In_219,In_446);
nand U92 (N_92,In_301,In_478);
nor U93 (N_93,In_384,In_354);
or U94 (N_94,In_291,In_388);
and U95 (N_95,In_207,In_101);
or U96 (N_96,In_97,In_127);
nor U97 (N_97,In_299,In_113);
or U98 (N_98,In_403,In_312);
nor U99 (N_99,In_376,In_460);
nand U100 (N_100,In_215,In_481);
or U101 (N_101,In_182,In_165);
xor U102 (N_102,In_278,In_471);
nand U103 (N_103,In_492,In_369);
or U104 (N_104,In_216,In_232);
nor U105 (N_105,In_337,In_296);
or U106 (N_106,In_8,In_133);
nand U107 (N_107,In_197,In_46);
xnor U108 (N_108,In_401,In_253);
and U109 (N_109,In_443,In_195);
or U110 (N_110,In_12,In_464);
nand U111 (N_111,In_316,In_251);
nand U112 (N_112,In_334,In_367);
or U113 (N_113,In_418,In_368);
nor U114 (N_114,In_260,In_233);
or U115 (N_115,In_257,In_274);
nand U116 (N_116,In_462,In_24);
nor U117 (N_117,In_198,In_415);
nand U118 (N_118,In_227,In_482);
nor U119 (N_119,In_82,In_87);
nand U120 (N_120,In_411,In_413);
and U121 (N_121,In_321,In_159);
or U122 (N_122,In_188,In_222);
or U123 (N_123,In_174,In_205);
or U124 (N_124,In_7,In_5);
nand U125 (N_125,In_155,In_55);
and U126 (N_126,In_333,In_365);
and U127 (N_127,In_436,In_342);
nor U128 (N_128,In_330,In_183);
nor U129 (N_129,In_276,In_293);
nand U130 (N_130,In_454,In_394);
and U131 (N_131,In_134,In_129);
nor U132 (N_132,In_311,In_479);
and U133 (N_133,In_153,In_158);
or U134 (N_134,In_336,In_68);
and U135 (N_135,In_397,In_187);
or U136 (N_136,In_250,In_366);
and U137 (N_137,In_341,In_352);
and U138 (N_138,In_315,In_178);
or U139 (N_139,In_451,In_437);
nand U140 (N_140,In_191,In_6);
or U141 (N_141,In_247,In_65);
nand U142 (N_142,In_273,In_254);
nor U143 (N_143,In_487,In_81);
and U144 (N_144,In_252,In_154);
or U145 (N_145,In_90,In_43);
nand U146 (N_146,In_79,In_47);
or U147 (N_147,In_292,In_389);
or U148 (N_148,In_300,In_52);
or U149 (N_149,In_399,In_398);
nor U150 (N_150,In_220,In_313);
nor U151 (N_151,In_262,In_175);
nand U152 (N_152,In_363,In_390);
nor U153 (N_153,In_211,In_206);
and U154 (N_154,In_26,In_86);
nor U155 (N_155,In_306,In_201);
nand U156 (N_156,In_246,In_33);
xnor U157 (N_157,In_307,In_290);
or U158 (N_158,In_317,In_288);
nand U159 (N_159,In_410,In_393);
nor U160 (N_160,In_177,In_242);
nor U161 (N_161,In_340,In_456);
or U162 (N_162,In_364,In_202);
nand U163 (N_163,In_346,In_66);
nand U164 (N_164,In_370,In_16);
or U165 (N_165,In_280,In_163);
nor U166 (N_166,In_223,In_450);
or U167 (N_167,In_249,In_131);
and U168 (N_168,In_434,In_122);
and U169 (N_169,In_140,In_373);
nor U170 (N_170,In_217,In_469);
and U171 (N_171,In_126,In_309);
or U172 (N_172,In_32,In_150);
and U173 (N_173,In_70,In_63);
or U174 (N_174,In_261,In_10);
and U175 (N_175,In_59,In_422);
nand U176 (N_176,In_157,In_486);
nor U177 (N_177,In_294,In_357);
nand U178 (N_178,In_360,In_184);
and U179 (N_179,In_14,In_431);
and U180 (N_180,In_147,In_277);
nor U181 (N_181,In_196,In_285);
nor U182 (N_182,In_148,In_269);
xnor U183 (N_183,In_427,In_54);
and U184 (N_184,In_490,In_74);
and U185 (N_185,In_329,In_453);
and U186 (N_186,In_38,In_179);
nor U187 (N_187,In_112,In_189);
or U188 (N_188,In_495,In_121);
and U189 (N_189,In_73,In_347);
and U190 (N_190,In_272,In_475);
nor U191 (N_191,In_442,In_445);
and U192 (N_192,In_99,In_102);
nor U193 (N_193,In_106,In_221);
and U194 (N_194,In_168,In_58);
nand U195 (N_195,In_103,In_428);
or U196 (N_196,In_56,In_302);
or U197 (N_197,In_193,In_459);
nand U198 (N_198,In_396,In_287);
nor U199 (N_199,In_4,In_169);
nor U200 (N_200,In_181,In_95);
and U201 (N_201,In_144,In_218);
or U202 (N_202,In_378,In_424);
nand U203 (N_203,In_391,In_170);
and U204 (N_204,In_332,In_162);
or U205 (N_205,In_28,In_11);
and U206 (N_206,In_236,In_335);
and U207 (N_207,In_387,In_297);
and U208 (N_208,In_234,In_409);
xor U209 (N_209,In_130,In_298);
nor U210 (N_210,In_50,In_359);
or U211 (N_211,In_176,In_37);
and U212 (N_212,In_353,In_372);
nor U213 (N_213,In_146,In_412);
and U214 (N_214,In_120,In_381);
and U215 (N_215,In_351,In_118);
nor U216 (N_216,In_470,In_42);
nor U217 (N_217,In_248,In_231);
nor U218 (N_218,In_420,In_480);
nand U219 (N_219,In_468,In_371);
or U220 (N_220,In_489,In_465);
and U221 (N_221,In_77,In_444);
and U222 (N_222,In_107,In_268);
and U223 (N_223,In_349,In_0);
nor U224 (N_224,In_53,In_499);
nor U225 (N_225,In_19,In_173);
nand U226 (N_226,In_83,In_319);
nand U227 (N_227,In_204,In_440);
nand U228 (N_228,In_472,In_21);
nor U229 (N_229,In_180,In_429);
or U230 (N_230,In_60,In_348);
xor U231 (N_231,In_125,In_138);
nor U232 (N_232,In_62,In_467);
and U233 (N_233,In_326,In_439);
or U234 (N_234,In_186,In_137);
nor U235 (N_235,In_406,In_49);
and U236 (N_236,In_458,In_88);
or U237 (N_237,In_25,In_485);
nand U238 (N_238,In_210,In_152);
and U239 (N_239,In_116,In_135);
nand U240 (N_240,In_171,In_105);
and U241 (N_241,In_69,In_343);
nand U242 (N_242,In_71,In_57);
or U243 (N_243,In_228,In_447);
and U244 (N_244,In_244,In_400);
nor U245 (N_245,In_91,In_226);
or U246 (N_246,In_308,In_96);
and U247 (N_247,In_48,In_386);
nor U248 (N_248,In_22,In_98);
or U249 (N_249,In_29,In_213);
xor U250 (N_250,In_396,In_139);
and U251 (N_251,In_293,In_9);
nand U252 (N_252,In_458,In_82);
or U253 (N_253,In_470,In_243);
and U254 (N_254,In_195,In_326);
or U255 (N_255,In_398,In_61);
or U256 (N_256,In_4,In_178);
nand U257 (N_257,In_233,In_116);
nand U258 (N_258,In_24,In_70);
nand U259 (N_259,In_75,In_103);
or U260 (N_260,In_271,In_285);
nand U261 (N_261,In_420,In_278);
nor U262 (N_262,In_138,In_98);
nor U263 (N_263,In_351,In_55);
nand U264 (N_264,In_403,In_0);
or U265 (N_265,In_21,In_154);
nor U266 (N_266,In_361,In_494);
nor U267 (N_267,In_374,In_237);
nand U268 (N_268,In_403,In_80);
nor U269 (N_269,In_83,In_220);
or U270 (N_270,In_152,In_493);
or U271 (N_271,In_262,In_324);
nor U272 (N_272,In_217,In_395);
nor U273 (N_273,In_385,In_226);
nand U274 (N_274,In_186,In_458);
nor U275 (N_275,In_96,In_238);
or U276 (N_276,In_330,In_69);
or U277 (N_277,In_486,In_136);
and U278 (N_278,In_257,In_27);
or U279 (N_279,In_98,In_31);
or U280 (N_280,In_278,In_105);
nand U281 (N_281,In_54,In_337);
and U282 (N_282,In_170,In_314);
nand U283 (N_283,In_373,In_210);
nor U284 (N_284,In_105,In_62);
or U285 (N_285,In_65,In_337);
nand U286 (N_286,In_283,In_231);
and U287 (N_287,In_141,In_442);
and U288 (N_288,In_397,In_386);
and U289 (N_289,In_18,In_21);
or U290 (N_290,In_136,In_235);
and U291 (N_291,In_152,In_432);
and U292 (N_292,In_272,In_55);
and U293 (N_293,In_473,In_305);
nand U294 (N_294,In_465,In_20);
nor U295 (N_295,In_220,In_165);
nand U296 (N_296,In_76,In_468);
or U297 (N_297,In_195,In_430);
nor U298 (N_298,In_67,In_78);
and U299 (N_299,In_476,In_174);
nor U300 (N_300,In_118,In_384);
xor U301 (N_301,In_77,In_109);
and U302 (N_302,In_432,In_125);
nor U303 (N_303,In_225,In_245);
nand U304 (N_304,In_131,In_212);
or U305 (N_305,In_259,In_66);
nand U306 (N_306,In_276,In_150);
or U307 (N_307,In_142,In_106);
and U308 (N_308,In_336,In_47);
and U309 (N_309,In_36,In_81);
nand U310 (N_310,In_86,In_263);
or U311 (N_311,In_21,In_190);
or U312 (N_312,In_263,In_447);
nand U313 (N_313,In_470,In_382);
nand U314 (N_314,In_180,In_192);
or U315 (N_315,In_126,In_177);
and U316 (N_316,In_78,In_492);
and U317 (N_317,In_55,In_443);
or U318 (N_318,In_248,In_327);
nand U319 (N_319,In_4,In_121);
and U320 (N_320,In_144,In_239);
or U321 (N_321,In_270,In_488);
nor U322 (N_322,In_92,In_416);
and U323 (N_323,In_150,In_79);
nor U324 (N_324,In_422,In_255);
and U325 (N_325,In_244,In_90);
or U326 (N_326,In_244,In_149);
and U327 (N_327,In_221,In_234);
and U328 (N_328,In_56,In_361);
nor U329 (N_329,In_341,In_109);
nor U330 (N_330,In_188,In_413);
nand U331 (N_331,In_84,In_251);
nor U332 (N_332,In_244,In_328);
and U333 (N_333,In_285,In_220);
nand U334 (N_334,In_138,In_104);
and U335 (N_335,In_249,In_330);
and U336 (N_336,In_136,In_412);
and U337 (N_337,In_92,In_175);
nor U338 (N_338,In_76,In_293);
nand U339 (N_339,In_410,In_164);
nand U340 (N_340,In_186,In_272);
nor U341 (N_341,In_228,In_495);
nand U342 (N_342,In_353,In_351);
nand U343 (N_343,In_302,In_47);
or U344 (N_344,In_33,In_359);
nor U345 (N_345,In_353,In_206);
and U346 (N_346,In_84,In_219);
or U347 (N_347,In_5,In_45);
nor U348 (N_348,In_146,In_197);
or U349 (N_349,In_483,In_91);
nor U350 (N_350,In_150,In_105);
and U351 (N_351,In_65,In_482);
nand U352 (N_352,In_324,In_18);
nand U353 (N_353,In_331,In_119);
nand U354 (N_354,In_11,In_84);
or U355 (N_355,In_416,In_167);
or U356 (N_356,In_393,In_254);
nand U357 (N_357,In_397,In_208);
xor U358 (N_358,In_335,In_145);
or U359 (N_359,In_224,In_360);
nor U360 (N_360,In_302,In_81);
nand U361 (N_361,In_485,In_496);
or U362 (N_362,In_58,In_212);
nor U363 (N_363,In_105,In_120);
or U364 (N_364,In_133,In_380);
xnor U365 (N_365,In_431,In_301);
and U366 (N_366,In_310,In_101);
or U367 (N_367,In_307,In_339);
and U368 (N_368,In_354,In_131);
and U369 (N_369,In_15,In_58);
nand U370 (N_370,In_195,In_383);
nor U371 (N_371,In_109,In_285);
or U372 (N_372,In_157,In_81);
and U373 (N_373,In_392,In_476);
or U374 (N_374,In_222,In_257);
and U375 (N_375,In_443,In_155);
nor U376 (N_376,In_201,In_339);
nand U377 (N_377,In_82,In_15);
nor U378 (N_378,In_181,In_29);
nand U379 (N_379,In_207,In_282);
nand U380 (N_380,In_208,In_484);
and U381 (N_381,In_429,In_117);
nor U382 (N_382,In_426,In_146);
nand U383 (N_383,In_97,In_443);
or U384 (N_384,In_31,In_468);
nand U385 (N_385,In_349,In_181);
or U386 (N_386,In_222,In_472);
nand U387 (N_387,In_72,In_401);
and U388 (N_388,In_61,In_380);
and U389 (N_389,In_482,In_201);
nor U390 (N_390,In_377,In_388);
or U391 (N_391,In_9,In_441);
and U392 (N_392,In_406,In_435);
and U393 (N_393,In_275,In_198);
nand U394 (N_394,In_339,In_64);
or U395 (N_395,In_313,In_394);
or U396 (N_396,In_90,In_67);
nor U397 (N_397,In_190,In_279);
and U398 (N_398,In_32,In_441);
or U399 (N_399,In_163,In_61);
nor U400 (N_400,In_330,In_337);
or U401 (N_401,In_431,In_238);
nor U402 (N_402,In_180,In_126);
and U403 (N_403,In_387,In_375);
nand U404 (N_404,In_282,In_397);
or U405 (N_405,In_447,In_173);
or U406 (N_406,In_265,In_423);
nor U407 (N_407,In_231,In_34);
or U408 (N_408,In_423,In_279);
nor U409 (N_409,In_278,In_248);
and U410 (N_410,In_494,In_147);
and U411 (N_411,In_121,In_302);
nor U412 (N_412,In_380,In_73);
nand U413 (N_413,In_228,In_114);
or U414 (N_414,In_304,In_407);
nor U415 (N_415,In_188,In_403);
nor U416 (N_416,In_408,In_342);
and U417 (N_417,In_198,In_130);
and U418 (N_418,In_1,In_244);
nand U419 (N_419,In_200,In_349);
or U420 (N_420,In_372,In_343);
nor U421 (N_421,In_283,In_225);
and U422 (N_422,In_157,In_192);
and U423 (N_423,In_438,In_346);
nand U424 (N_424,In_304,In_399);
or U425 (N_425,In_236,In_153);
and U426 (N_426,In_280,In_474);
or U427 (N_427,In_493,In_210);
nand U428 (N_428,In_462,In_194);
nor U429 (N_429,In_308,In_446);
xor U430 (N_430,In_303,In_39);
nand U431 (N_431,In_433,In_398);
nand U432 (N_432,In_120,In_48);
nor U433 (N_433,In_255,In_175);
nor U434 (N_434,In_109,In_100);
nand U435 (N_435,In_237,In_296);
nor U436 (N_436,In_311,In_97);
nor U437 (N_437,In_498,In_158);
and U438 (N_438,In_320,In_377);
and U439 (N_439,In_441,In_169);
and U440 (N_440,In_485,In_63);
and U441 (N_441,In_105,In_496);
nor U442 (N_442,In_103,In_367);
or U443 (N_443,In_164,In_281);
and U444 (N_444,In_192,In_55);
nand U445 (N_445,In_233,In_361);
and U446 (N_446,In_453,In_153);
nand U447 (N_447,In_258,In_468);
and U448 (N_448,In_353,In_18);
and U449 (N_449,In_343,In_312);
nor U450 (N_450,In_481,In_205);
or U451 (N_451,In_197,In_412);
nor U452 (N_452,In_475,In_450);
or U453 (N_453,In_268,In_181);
nor U454 (N_454,In_316,In_166);
nand U455 (N_455,In_78,In_61);
nor U456 (N_456,In_108,In_404);
or U457 (N_457,In_244,In_144);
and U458 (N_458,In_403,In_208);
and U459 (N_459,In_296,In_449);
nand U460 (N_460,In_232,In_93);
nand U461 (N_461,In_27,In_129);
nand U462 (N_462,In_444,In_360);
or U463 (N_463,In_211,In_481);
nor U464 (N_464,In_202,In_307);
nor U465 (N_465,In_207,In_447);
or U466 (N_466,In_414,In_164);
nor U467 (N_467,In_377,In_489);
nand U468 (N_468,In_10,In_427);
or U469 (N_469,In_441,In_221);
nand U470 (N_470,In_137,In_204);
nand U471 (N_471,In_285,In_167);
or U472 (N_472,In_147,In_210);
nand U473 (N_473,In_185,In_403);
nand U474 (N_474,In_107,In_307);
and U475 (N_475,In_150,In_218);
nor U476 (N_476,In_139,In_437);
or U477 (N_477,In_473,In_483);
nor U478 (N_478,In_307,In_277);
nand U479 (N_479,In_6,In_434);
or U480 (N_480,In_35,In_396);
nand U481 (N_481,In_151,In_290);
nand U482 (N_482,In_417,In_296);
or U483 (N_483,In_58,In_334);
or U484 (N_484,In_368,In_247);
nand U485 (N_485,In_12,In_421);
and U486 (N_486,In_252,In_202);
nor U487 (N_487,In_341,In_404);
nor U488 (N_488,In_208,In_185);
nor U489 (N_489,In_39,In_309);
nand U490 (N_490,In_160,In_6);
and U491 (N_491,In_23,In_423);
nand U492 (N_492,In_474,In_274);
nor U493 (N_493,In_352,In_132);
nor U494 (N_494,In_377,In_493);
and U495 (N_495,In_483,In_432);
or U496 (N_496,In_463,In_79);
nor U497 (N_497,In_99,In_490);
and U498 (N_498,In_167,In_45);
and U499 (N_499,In_296,In_330);
nor U500 (N_500,In_407,In_100);
nor U501 (N_501,In_271,In_6);
xnor U502 (N_502,In_463,In_175);
xor U503 (N_503,In_487,In_3);
and U504 (N_504,In_489,In_25);
or U505 (N_505,In_487,In_324);
or U506 (N_506,In_338,In_30);
nor U507 (N_507,In_274,In_53);
and U508 (N_508,In_347,In_380);
and U509 (N_509,In_186,In_302);
and U510 (N_510,In_82,In_499);
nand U511 (N_511,In_117,In_126);
nor U512 (N_512,In_353,In_196);
nand U513 (N_513,In_116,In_62);
and U514 (N_514,In_263,In_465);
nand U515 (N_515,In_197,In_228);
or U516 (N_516,In_321,In_227);
and U517 (N_517,In_247,In_58);
and U518 (N_518,In_222,In_292);
and U519 (N_519,In_24,In_192);
nor U520 (N_520,In_381,In_56);
nand U521 (N_521,In_349,In_375);
nor U522 (N_522,In_33,In_109);
nand U523 (N_523,In_431,In_73);
and U524 (N_524,In_311,In_420);
and U525 (N_525,In_467,In_4);
nand U526 (N_526,In_402,In_122);
or U527 (N_527,In_64,In_255);
nor U528 (N_528,In_229,In_82);
nor U529 (N_529,In_104,In_232);
and U530 (N_530,In_69,In_156);
nor U531 (N_531,In_271,In_448);
nor U532 (N_532,In_196,In_487);
or U533 (N_533,In_121,In_23);
and U534 (N_534,In_26,In_406);
and U535 (N_535,In_393,In_85);
and U536 (N_536,In_464,In_267);
or U537 (N_537,In_189,In_281);
or U538 (N_538,In_244,In_80);
or U539 (N_539,In_343,In_242);
or U540 (N_540,In_29,In_375);
and U541 (N_541,In_495,In_499);
or U542 (N_542,In_321,In_218);
nand U543 (N_543,In_345,In_421);
nand U544 (N_544,In_5,In_312);
nor U545 (N_545,In_268,In_334);
or U546 (N_546,In_127,In_185);
nor U547 (N_547,In_61,In_152);
nor U548 (N_548,In_483,In_499);
nor U549 (N_549,In_100,In_281);
nand U550 (N_550,In_163,In_388);
nand U551 (N_551,In_134,In_302);
nand U552 (N_552,In_5,In_24);
nor U553 (N_553,In_450,In_332);
nor U554 (N_554,In_333,In_481);
and U555 (N_555,In_32,In_260);
or U556 (N_556,In_111,In_5);
nor U557 (N_557,In_46,In_297);
or U558 (N_558,In_158,In_146);
or U559 (N_559,In_27,In_315);
nand U560 (N_560,In_194,In_321);
or U561 (N_561,In_71,In_489);
and U562 (N_562,In_305,In_281);
and U563 (N_563,In_109,In_355);
and U564 (N_564,In_326,In_55);
nand U565 (N_565,In_151,In_246);
and U566 (N_566,In_78,In_351);
or U567 (N_567,In_448,In_212);
xor U568 (N_568,In_376,In_358);
nand U569 (N_569,In_163,In_154);
or U570 (N_570,In_169,In_55);
and U571 (N_571,In_281,In_456);
and U572 (N_572,In_350,In_343);
nand U573 (N_573,In_458,In_91);
and U574 (N_574,In_385,In_68);
nor U575 (N_575,In_61,In_39);
nand U576 (N_576,In_403,In_283);
nand U577 (N_577,In_212,In_78);
nand U578 (N_578,In_484,In_163);
nand U579 (N_579,In_71,In_47);
or U580 (N_580,In_36,In_165);
and U581 (N_581,In_469,In_488);
nand U582 (N_582,In_267,In_433);
and U583 (N_583,In_66,In_464);
nand U584 (N_584,In_7,In_305);
nand U585 (N_585,In_165,In_407);
or U586 (N_586,In_8,In_117);
or U587 (N_587,In_263,In_201);
or U588 (N_588,In_235,In_38);
nor U589 (N_589,In_188,In_91);
nor U590 (N_590,In_195,In_159);
nand U591 (N_591,In_123,In_26);
nand U592 (N_592,In_347,In_37);
and U593 (N_593,In_34,In_57);
nor U594 (N_594,In_126,In_265);
nand U595 (N_595,In_135,In_180);
nor U596 (N_596,In_16,In_77);
nor U597 (N_597,In_169,In_157);
and U598 (N_598,In_403,In_413);
or U599 (N_599,In_309,In_223);
nand U600 (N_600,In_344,In_446);
and U601 (N_601,In_315,In_338);
or U602 (N_602,In_304,In_344);
nor U603 (N_603,In_95,In_447);
nand U604 (N_604,In_48,In_431);
or U605 (N_605,In_196,In_286);
nand U606 (N_606,In_386,In_442);
nand U607 (N_607,In_197,In_435);
nor U608 (N_608,In_288,In_302);
or U609 (N_609,In_342,In_28);
or U610 (N_610,In_275,In_442);
nor U611 (N_611,In_385,In_223);
nor U612 (N_612,In_416,In_156);
nor U613 (N_613,In_300,In_271);
xor U614 (N_614,In_354,In_78);
nor U615 (N_615,In_256,In_232);
nand U616 (N_616,In_40,In_235);
or U617 (N_617,In_323,In_208);
and U618 (N_618,In_149,In_156);
and U619 (N_619,In_438,In_101);
and U620 (N_620,In_45,In_498);
nor U621 (N_621,In_271,In_34);
nand U622 (N_622,In_373,In_313);
or U623 (N_623,In_368,In_207);
nand U624 (N_624,In_429,In_168);
and U625 (N_625,In_123,In_54);
and U626 (N_626,In_130,In_438);
nand U627 (N_627,In_197,In_362);
nor U628 (N_628,In_236,In_93);
or U629 (N_629,In_79,In_460);
and U630 (N_630,In_236,In_227);
nor U631 (N_631,In_405,In_203);
nand U632 (N_632,In_229,In_436);
nand U633 (N_633,In_283,In_184);
nand U634 (N_634,In_175,In_201);
and U635 (N_635,In_217,In_485);
or U636 (N_636,In_356,In_280);
nor U637 (N_637,In_52,In_87);
or U638 (N_638,In_50,In_258);
nand U639 (N_639,In_185,In_106);
nand U640 (N_640,In_133,In_126);
and U641 (N_641,In_338,In_269);
and U642 (N_642,In_164,In_113);
nor U643 (N_643,In_373,In_76);
nor U644 (N_644,In_173,In_57);
nor U645 (N_645,In_90,In_198);
nand U646 (N_646,In_104,In_89);
and U647 (N_647,In_415,In_370);
and U648 (N_648,In_59,In_78);
nor U649 (N_649,In_352,In_22);
nor U650 (N_650,In_369,In_491);
and U651 (N_651,In_293,In_88);
and U652 (N_652,In_219,In_307);
and U653 (N_653,In_332,In_120);
nor U654 (N_654,In_233,In_210);
nor U655 (N_655,In_371,In_112);
or U656 (N_656,In_267,In_352);
and U657 (N_657,In_468,In_33);
and U658 (N_658,In_445,In_47);
or U659 (N_659,In_135,In_228);
or U660 (N_660,In_114,In_217);
nand U661 (N_661,In_276,In_77);
nor U662 (N_662,In_117,In_13);
nor U663 (N_663,In_471,In_113);
or U664 (N_664,In_288,In_142);
nand U665 (N_665,In_358,In_398);
and U666 (N_666,In_20,In_8);
and U667 (N_667,In_327,In_273);
xnor U668 (N_668,In_209,In_497);
nand U669 (N_669,In_319,In_32);
nor U670 (N_670,In_373,In_434);
or U671 (N_671,In_262,In_22);
nand U672 (N_672,In_112,In_457);
and U673 (N_673,In_281,In_482);
or U674 (N_674,In_309,In_355);
nor U675 (N_675,In_263,In_234);
and U676 (N_676,In_54,In_16);
xnor U677 (N_677,In_54,In_89);
nor U678 (N_678,In_252,In_405);
nor U679 (N_679,In_434,In_282);
or U680 (N_680,In_476,In_460);
nor U681 (N_681,In_258,In_120);
nor U682 (N_682,In_204,In_104);
nor U683 (N_683,In_397,In_296);
nor U684 (N_684,In_259,In_370);
or U685 (N_685,In_243,In_69);
and U686 (N_686,In_490,In_249);
or U687 (N_687,In_365,In_134);
nor U688 (N_688,In_309,In_331);
nand U689 (N_689,In_494,In_199);
nor U690 (N_690,In_487,In_201);
nand U691 (N_691,In_12,In_431);
and U692 (N_692,In_104,In_400);
and U693 (N_693,In_412,In_336);
nand U694 (N_694,In_141,In_289);
and U695 (N_695,In_21,In_102);
and U696 (N_696,In_127,In_199);
xor U697 (N_697,In_290,In_318);
and U698 (N_698,In_1,In_460);
and U699 (N_699,In_459,In_388);
and U700 (N_700,In_105,In_140);
or U701 (N_701,In_281,In_410);
and U702 (N_702,In_418,In_469);
or U703 (N_703,In_498,In_258);
nor U704 (N_704,In_128,In_293);
nor U705 (N_705,In_2,In_265);
nand U706 (N_706,In_303,In_423);
and U707 (N_707,In_123,In_263);
or U708 (N_708,In_90,In_99);
and U709 (N_709,In_327,In_252);
and U710 (N_710,In_306,In_244);
xnor U711 (N_711,In_205,In_438);
nor U712 (N_712,In_322,In_288);
or U713 (N_713,In_11,In_471);
nand U714 (N_714,In_485,In_418);
or U715 (N_715,In_331,In_269);
xor U716 (N_716,In_221,In_118);
nand U717 (N_717,In_444,In_18);
nand U718 (N_718,In_0,In_373);
and U719 (N_719,In_302,In_5);
nand U720 (N_720,In_376,In_150);
nor U721 (N_721,In_75,In_417);
nor U722 (N_722,In_491,In_296);
or U723 (N_723,In_54,In_416);
nor U724 (N_724,In_126,In_317);
nand U725 (N_725,In_280,In_21);
or U726 (N_726,In_241,In_187);
and U727 (N_727,In_431,In_60);
nand U728 (N_728,In_25,In_381);
and U729 (N_729,In_11,In_41);
nand U730 (N_730,In_172,In_464);
nor U731 (N_731,In_302,In_469);
or U732 (N_732,In_356,In_38);
nand U733 (N_733,In_470,In_73);
nor U734 (N_734,In_248,In_194);
or U735 (N_735,In_229,In_372);
nand U736 (N_736,In_202,In_206);
nand U737 (N_737,In_254,In_107);
and U738 (N_738,In_230,In_457);
or U739 (N_739,In_447,In_137);
nor U740 (N_740,In_262,In_334);
and U741 (N_741,In_202,In_415);
nor U742 (N_742,In_36,In_116);
or U743 (N_743,In_29,In_44);
nand U744 (N_744,In_5,In_112);
nor U745 (N_745,In_364,In_428);
and U746 (N_746,In_205,In_470);
xor U747 (N_747,In_45,In_81);
nor U748 (N_748,In_102,In_264);
nand U749 (N_749,In_103,In_479);
nand U750 (N_750,In_138,In_346);
nor U751 (N_751,In_375,In_310);
and U752 (N_752,In_221,In_115);
nor U753 (N_753,In_92,In_24);
or U754 (N_754,In_114,In_391);
nand U755 (N_755,In_101,In_114);
or U756 (N_756,In_380,In_441);
or U757 (N_757,In_222,In_186);
nand U758 (N_758,In_330,In_383);
and U759 (N_759,In_171,In_95);
or U760 (N_760,In_118,In_300);
or U761 (N_761,In_166,In_164);
and U762 (N_762,In_220,In_325);
and U763 (N_763,In_446,In_293);
and U764 (N_764,In_4,In_357);
nand U765 (N_765,In_371,In_485);
or U766 (N_766,In_144,In_174);
and U767 (N_767,In_472,In_376);
and U768 (N_768,In_217,In_37);
and U769 (N_769,In_7,In_296);
or U770 (N_770,In_462,In_18);
or U771 (N_771,In_392,In_44);
and U772 (N_772,In_20,In_175);
nand U773 (N_773,In_154,In_308);
nor U774 (N_774,In_35,In_495);
nand U775 (N_775,In_344,In_325);
nand U776 (N_776,In_176,In_131);
xor U777 (N_777,In_110,In_407);
nand U778 (N_778,In_147,In_489);
and U779 (N_779,In_171,In_123);
nand U780 (N_780,In_112,In_64);
nor U781 (N_781,In_151,In_187);
or U782 (N_782,In_189,In_11);
or U783 (N_783,In_369,In_172);
and U784 (N_784,In_363,In_365);
and U785 (N_785,In_29,In_18);
nor U786 (N_786,In_318,In_194);
nor U787 (N_787,In_286,In_28);
nor U788 (N_788,In_366,In_1);
nor U789 (N_789,In_305,In_347);
and U790 (N_790,In_8,In_131);
or U791 (N_791,In_353,In_187);
or U792 (N_792,In_268,In_231);
nor U793 (N_793,In_24,In_30);
and U794 (N_794,In_166,In_196);
nand U795 (N_795,In_116,In_162);
and U796 (N_796,In_391,In_45);
or U797 (N_797,In_436,In_135);
or U798 (N_798,In_328,In_59);
and U799 (N_799,In_303,In_87);
nand U800 (N_800,In_202,In_170);
nand U801 (N_801,In_88,In_275);
and U802 (N_802,In_286,In_363);
nand U803 (N_803,In_277,In_176);
and U804 (N_804,In_327,In_29);
and U805 (N_805,In_108,In_395);
and U806 (N_806,In_72,In_108);
nand U807 (N_807,In_221,In_86);
nor U808 (N_808,In_453,In_457);
xnor U809 (N_809,In_411,In_225);
and U810 (N_810,In_8,In_386);
nand U811 (N_811,In_417,In_181);
nor U812 (N_812,In_259,In_398);
and U813 (N_813,In_427,In_83);
nor U814 (N_814,In_366,In_152);
nand U815 (N_815,In_239,In_96);
nor U816 (N_816,In_111,In_478);
nand U817 (N_817,In_21,In_113);
nor U818 (N_818,In_228,In_297);
nand U819 (N_819,In_204,In_441);
and U820 (N_820,In_176,In_393);
xor U821 (N_821,In_288,In_117);
nand U822 (N_822,In_75,In_105);
nor U823 (N_823,In_343,In_197);
nor U824 (N_824,In_312,In_142);
nor U825 (N_825,In_478,In_281);
and U826 (N_826,In_245,In_2);
or U827 (N_827,In_182,In_155);
or U828 (N_828,In_95,In_167);
nor U829 (N_829,In_202,In_386);
nand U830 (N_830,In_28,In_496);
nor U831 (N_831,In_293,In_472);
nand U832 (N_832,In_468,In_176);
and U833 (N_833,In_495,In_287);
and U834 (N_834,In_221,In_418);
nand U835 (N_835,In_480,In_242);
or U836 (N_836,In_151,In_308);
and U837 (N_837,In_487,In_142);
and U838 (N_838,In_88,In_419);
and U839 (N_839,In_51,In_140);
and U840 (N_840,In_379,In_297);
or U841 (N_841,In_485,In_109);
and U842 (N_842,In_317,In_121);
nor U843 (N_843,In_6,In_87);
nor U844 (N_844,In_48,In_359);
nor U845 (N_845,In_89,In_460);
or U846 (N_846,In_19,In_297);
xnor U847 (N_847,In_379,In_182);
nor U848 (N_848,In_338,In_44);
or U849 (N_849,In_106,In_388);
or U850 (N_850,In_104,In_355);
nand U851 (N_851,In_467,In_468);
and U852 (N_852,In_224,In_304);
nand U853 (N_853,In_291,In_61);
or U854 (N_854,In_441,In_172);
nor U855 (N_855,In_1,In_314);
or U856 (N_856,In_499,In_497);
nand U857 (N_857,In_74,In_173);
and U858 (N_858,In_340,In_245);
nand U859 (N_859,In_206,In_402);
or U860 (N_860,In_215,In_267);
nand U861 (N_861,In_270,In_421);
and U862 (N_862,In_317,In_87);
and U863 (N_863,In_166,In_258);
or U864 (N_864,In_311,In_0);
nor U865 (N_865,In_254,In_437);
nor U866 (N_866,In_110,In_144);
or U867 (N_867,In_338,In_452);
nor U868 (N_868,In_277,In_88);
or U869 (N_869,In_29,In_456);
or U870 (N_870,In_418,In_476);
and U871 (N_871,In_224,In_227);
or U872 (N_872,In_27,In_376);
nor U873 (N_873,In_334,In_409);
xnor U874 (N_874,In_40,In_211);
nand U875 (N_875,In_462,In_200);
and U876 (N_876,In_107,In_344);
or U877 (N_877,In_241,In_283);
nand U878 (N_878,In_221,In_397);
nor U879 (N_879,In_99,In_497);
nor U880 (N_880,In_487,In_477);
nor U881 (N_881,In_31,In_29);
nor U882 (N_882,In_132,In_15);
nand U883 (N_883,In_71,In_187);
or U884 (N_884,In_412,In_31);
nand U885 (N_885,In_360,In_474);
nor U886 (N_886,In_438,In_203);
nor U887 (N_887,In_367,In_420);
and U888 (N_888,In_434,In_491);
nor U889 (N_889,In_194,In_416);
and U890 (N_890,In_461,In_66);
xor U891 (N_891,In_302,In_262);
nand U892 (N_892,In_301,In_495);
or U893 (N_893,In_91,In_454);
and U894 (N_894,In_330,In_64);
nand U895 (N_895,In_349,In_206);
and U896 (N_896,In_235,In_398);
or U897 (N_897,In_149,In_15);
or U898 (N_898,In_103,In_195);
nor U899 (N_899,In_99,In_341);
nand U900 (N_900,In_481,In_357);
nor U901 (N_901,In_163,In_462);
and U902 (N_902,In_259,In_23);
or U903 (N_903,In_108,In_436);
or U904 (N_904,In_142,In_63);
and U905 (N_905,In_327,In_443);
nor U906 (N_906,In_475,In_215);
and U907 (N_907,In_98,In_96);
nand U908 (N_908,In_217,In_109);
and U909 (N_909,In_352,In_311);
nor U910 (N_910,In_165,In_243);
and U911 (N_911,In_313,In_46);
nor U912 (N_912,In_152,In_427);
and U913 (N_913,In_399,In_450);
or U914 (N_914,In_457,In_298);
or U915 (N_915,In_250,In_382);
nand U916 (N_916,In_264,In_407);
or U917 (N_917,In_142,In_62);
or U918 (N_918,In_440,In_228);
and U919 (N_919,In_383,In_354);
nor U920 (N_920,In_394,In_97);
and U921 (N_921,In_448,In_149);
nand U922 (N_922,In_268,In_323);
and U923 (N_923,In_141,In_60);
or U924 (N_924,In_342,In_238);
nand U925 (N_925,In_396,In_329);
nor U926 (N_926,In_294,In_16);
nand U927 (N_927,In_359,In_430);
or U928 (N_928,In_435,In_238);
or U929 (N_929,In_214,In_491);
and U930 (N_930,In_310,In_336);
and U931 (N_931,In_122,In_467);
and U932 (N_932,In_271,In_265);
nand U933 (N_933,In_108,In_81);
or U934 (N_934,In_374,In_208);
nor U935 (N_935,In_62,In_234);
or U936 (N_936,In_39,In_84);
or U937 (N_937,In_105,In_182);
nand U938 (N_938,In_483,In_334);
or U939 (N_939,In_187,In_91);
nand U940 (N_940,In_165,In_329);
nand U941 (N_941,In_282,In_336);
nor U942 (N_942,In_255,In_139);
and U943 (N_943,In_216,In_62);
and U944 (N_944,In_241,In_489);
nor U945 (N_945,In_358,In_275);
and U946 (N_946,In_188,In_24);
nor U947 (N_947,In_239,In_92);
nand U948 (N_948,In_8,In_114);
and U949 (N_949,In_89,In_377);
xnor U950 (N_950,In_221,In_371);
and U951 (N_951,In_46,In_343);
nand U952 (N_952,In_468,In_336);
and U953 (N_953,In_496,In_277);
and U954 (N_954,In_134,In_126);
and U955 (N_955,In_381,In_217);
or U956 (N_956,In_497,In_438);
or U957 (N_957,In_279,In_278);
or U958 (N_958,In_19,In_216);
xor U959 (N_959,In_124,In_19);
nand U960 (N_960,In_151,In_427);
or U961 (N_961,In_203,In_417);
or U962 (N_962,In_221,In_338);
and U963 (N_963,In_487,In_75);
nor U964 (N_964,In_363,In_105);
and U965 (N_965,In_14,In_79);
and U966 (N_966,In_48,In_280);
and U967 (N_967,In_47,In_223);
or U968 (N_968,In_127,In_59);
nand U969 (N_969,In_466,In_220);
nand U970 (N_970,In_444,In_345);
nor U971 (N_971,In_46,In_245);
xor U972 (N_972,In_38,In_291);
nand U973 (N_973,In_190,In_275);
and U974 (N_974,In_20,In_252);
nor U975 (N_975,In_176,In_403);
nor U976 (N_976,In_315,In_192);
nand U977 (N_977,In_93,In_230);
nand U978 (N_978,In_382,In_1);
nand U979 (N_979,In_499,In_372);
nand U980 (N_980,In_269,In_25);
nor U981 (N_981,In_57,In_466);
nand U982 (N_982,In_430,In_156);
and U983 (N_983,In_472,In_448);
nand U984 (N_984,In_73,In_126);
nor U985 (N_985,In_146,In_372);
nand U986 (N_986,In_243,In_483);
nand U987 (N_987,In_99,In_418);
and U988 (N_988,In_82,In_251);
or U989 (N_989,In_486,In_90);
nor U990 (N_990,In_76,In_146);
or U991 (N_991,In_380,In_95);
nand U992 (N_992,In_155,In_260);
nand U993 (N_993,In_105,In_497);
nor U994 (N_994,In_443,In_16);
nand U995 (N_995,In_5,In_294);
and U996 (N_996,In_11,In_411);
or U997 (N_997,In_74,In_179);
nand U998 (N_998,In_429,In_441);
nand U999 (N_999,In_365,In_420);
nand U1000 (N_1000,N_164,N_87);
nor U1001 (N_1001,N_808,N_48);
xnor U1002 (N_1002,N_274,N_818);
and U1003 (N_1003,N_14,N_157);
nor U1004 (N_1004,N_548,N_773);
or U1005 (N_1005,N_79,N_108);
nor U1006 (N_1006,N_880,N_951);
or U1007 (N_1007,N_500,N_170);
nor U1008 (N_1008,N_696,N_955);
nor U1009 (N_1009,N_94,N_564);
nand U1010 (N_1010,N_238,N_360);
and U1011 (N_1011,N_252,N_332);
and U1012 (N_1012,N_146,N_405);
and U1013 (N_1013,N_900,N_710);
nand U1014 (N_1014,N_557,N_396);
nand U1015 (N_1015,N_546,N_952);
nor U1016 (N_1016,N_203,N_802);
nand U1017 (N_1017,N_188,N_181);
nand U1018 (N_1018,N_941,N_996);
and U1019 (N_1019,N_477,N_39);
nor U1020 (N_1020,N_91,N_662);
and U1021 (N_1021,N_311,N_573);
and U1022 (N_1022,N_531,N_308);
and U1023 (N_1023,N_757,N_118);
nor U1024 (N_1024,N_112,N_836);
nand U1025 (N_1025,N_290,N_226);
nand U1026 (N_1026,N_392,N_465);
nor U1027 (N_1027,N_643,N_798);
nor U1028 (N_1028,N_160,N_421);
and U1029 (N_1029,N_737,N_544);
nor U1030 (N_1030,N_47,N_330);
nor U1031 (N_1031,N_336,N_136);
nor U1032 (N_1032,N_819,N_523);
nor U1033 (N_1033,N_799,N_556);
nand U1034 (N_1034,N_953,N_492);
nand U1035 (N_1035,N_369,N_797);
nand U1036 (N_1036,N_199,N_398);
nand U1037 (N_1037,N_755,N_859);
nand U1038 (N_1038,N_165,N_242);
nand U1039 (N_1039,N_584,N_933);
nor U1040 (N_1040,N_432,N_123);
xor U1041 (N_1041,N_966,N_590);
or U1042 (N_1042,N_293,N_927);
nand U1043 (N_1043,N_302,N_917);
nand U1044 (N_1044,N_697,N_960);
nor U1045 (N_1045,N_763,N_267);
and U1046 (N_1046,N_65,N_762);
nand U1047 (N_1047,N_345,N_152);
or U1048 (N_1048,N_50,N_721);
nor U1049 (N_1049,N_256,N_756);
nand U1050 (N_1050,N_273,N_37);
and U1051 (N_1051,N_230,N_134);
nand U1052 (N_1052,N_17,N_541);
or U1053 (N_1053,N_715,N_71);
and U1054 (N_1054,N_514,N_420);
or U1055 (N_1055,N_816,N_518);
and U1056 (N_1056,N_587,N_645);
nand U1057 (N_1057,N_64,N_839);
nor U1058 (N_1058,N_542,N_881);
nand U1059 (N_1059,N_474,N_426);
nand U1060 (N_1060,N_605,N_980);
or U1061 (N_1061,N_488,N_809);
or U1062 (N_1062,N_942,N_926);
and U1063 (N_1063,N_55,N_22);
nor U1064 (N_1064,N_923,N_574);
nand U1065 (N_1065,N_262,N_61);
xor U1066 (N_1066,N_856,N_716);
nor U1067 (N_1067,N_648,N_578);
nand U1068 (N_1068,N_81,N_462);
nor U1069 (N_1069,N_529,N_476);
nor U1070 (N_1070,N_101,N_359);
or U1071 (N_1071,N_992,N_525);
and U1072 (N_1072,N_785,N_990);
nand U1073 (N_1073,N_860,N_385);
nor U1074 (N_1074,N_51,N_567);
nor U1075 (N_1075,N_822,N_231);
nand U1076 (N_1076,N_604,N_434);
nand U1077 (N_1077,N_389,N_391);
nand U1078 (N_1078,N_347,N_781);
nor U1079 (N_1079,N_335,N_328);
or U1080 (N_1080,N_357,N_814);
or U1081 (N_1081,N_237,N_467);
and U1082 (N_1082,N_764,N_227);
and U1083 (N_1083,N_769,N_639);
and U1084 (N_1084,N_774,N_19);
or U1085 (N_1085,N_495,N_443);
nand U1086 (N_1086,N_982,N_779);
nor U1087 (N_1087,N_34,N_649);
or U1088 (N_1088,N_121,N_104);
and U1089 (N_1089,N_922,N_706);
or U1090 (N_1090,N_276,N_855);
and U1091 (N_1091,N_632,N_868);
and U1092 (N_1092,N_122,N_565);
nand U1093 (N_1093,N_260,N_588);
nor U1094 (N_1094,N_130,N_172);
and U1095 (N_1095,N_343,N_791);
and U1096 (N_1096,N_166,N_538);
or U1097 (N_1097,N_93,N_520);
or U1098 (N_1098,N_246,N_12);
and U1099 (N_1099,N_796,N_449);
nor U1100 (N_1100,N_220,N_837);
or U1101 (N_1101,N_852,N_26);
nor U1102 (N_1102,N_602,N_326);
or U1103 (N_1103,N_218,N_247);
nor U1104 (N_1104,N_793,N_265);
and U1105 (N_1105,N_787,N_853);
and U1106 (N_1106,N_349,N_912);
nand U1107 (N_1107,N_185,N_29);
or U1108 (N_1108,N_315,N_772);
nor U1109 (N_1109,N_88,N_422);
nand U1110 (N_1110,N_279,N_11);
nor U1111 (N_1111,N_981,N_489);
xor U1112 (N_1112,N_415,N_381);
or U1113 (N_1113,N_636,N_968);
nand U1114 (N_1114,N_901,N_760);
nand U1115 (N_1115,N_561,N_599);
or U1116 (N_1116,N_127,N_507);
or U1117 (N_1117,N_191,N_131);
and U1118 (N_1118,N_961,N_299);
nand U1119 (N_1119,N_90,N_743);
or U1120 (N_1120,N_511,N_189);
nor U1121 (N_1121,N_586,N_251);
or U1122 (N_1122,N_195,N_619);
and U1123 (N_1123,N_125,N_817);
or U1124 (N_1124,N_888,N_194);
nand U1125 (N_1125,N_74,N_987);
nand U1126 (N_1126,N_691,N_702);
or U1127 (N_1127,N_496,N_378);
or U1128 (N_1128,N_713,N_254);
and U1129 (N_1129,N_789,N_845);
xor U1130 (N_1130,N_724,N_271);
nand U1131 (N_1131,N_775,N_998);
or U1132 (N_1132,N_733,N_413);
nor U1133 (N_1133,N_228,N_482);
or U1134 (N_1134,N_283,N_698);
and U1135 (N_1135,N_610,N_641);
xnor U1136 (N_1136,N_843,N_92);
and U1137 (N_1137,N_803,N_934);
nand U1138 (N_1138,N_263,N_439);
nor U1139 (N_1139,N_483,N_205);
or U1140 (N_1140,N_659,N_76);
nor U1141 (N_1141,N_402,N_660);
nor U1142 (N_1142,N_569,N_24);
and U1143 (N_1143,N_204,N_686);
nor U1144 (N_1144,N_709,N_921);
nor U1145 (N_1145,N_895,N_431);
or U1146 (N_1146,N_609,N_171);
and U1147 (N_1147,N_493,N_280);
or U1148 (N_1148,N_98,N_635);
and U1149 (N_1149,N_206,N_365);
and U1150 (N_1150,N_616,N_508);
nor U1151 (N_1151,N_806,N_549);
nand U1152 (N_1152,N_284,N_63);
nor U1153 (N_1153,N_509,N_820);
nand U1154 (N_1154,N_295,N_657);
and U1155 (N_1155,N_909,N_794);
nand U1156 (N_1156,N_801,N_846);
and U1157 (N_1157,N_878,N_989);
nor U1158 (N_1158,N_54,N_478);
nand U1159 (N_1159,N_182,N_135);
xnor U1160 (N_1160,N_929,N_249);
or U1161 (N_1161,N_986,N_219);
or U1162 (N_1162,N_240,N_351);
and U1163 (N_1163,N_813,N_133);
and U1164 (N_1164,N_664,N_617);
or U1165 (N_1165,N_628,N_82);
nor U1166 (N_1166,N_43,N_180);
and U1167 (N_1167,N_999,N_902);
and U1168 (N_1168,N_370,N_30);
xnor U1169 (N_1169,N_891,N_253);
and U1170 (N_1170,N_766,N_298);
nand U1171 (N_1171,N_4,N_897);
and U1172 (N_1172,N_811,N_75);
nor U1173 (N_1173,N_212,N_651);
nand U1174 (N_1174,N_908,N_414);
nor U1175 (N_1175,N_368,N_915);
nor U1176 (N_1176,N_409,N_487);
or U1177 (N_1177,N_581,N_233);
or U1178 (N_1178,N_3,N_655);
and U1179 (N_1179,N_364,N_899);
nand U1180 (N_1180,N_670,N_301);
and U1181 (N_1181,N_685,N_903);
nand U1182 (N_1182,N_945,N_503);
and U1183 (N_1183,N_949,N_150);
nor U1184 (N_1184,N_380,N_935);
nor U1185 (N_1185,N_338,N_494);
xnor U1186 (N_1186,N_887,N_403);
or U1187 (N_1187,N_472,N_306);
nand U1188 (N_1188,N_107,N_484);
nor U1189 (N_1189,N_570,N_976);
or U1190 (N_1190,N_235,N_223);
nand U1191 (N_1191,N_23,N_727);
or U1192 (N_1192,N_770,N_20);
nor U1193 (N_1193,N_914,N_857);
nand U1194 (N_1194,N_339,N_292);
or U1195 (N_1195,N_674,N_612);
and U1196 (N_1196,N_278,N_984);
nand U1197 (N_1197,N_348,N_720);
and U1198 (N_1198,N_889,N_374);
nor U1199 (N_1199,N_103,N_867);
or U1200 (N_1200,N_694,N_625);
and U1201 (N_1201,N_501,N_159);
or U1202 (N_1202,N_681,N_675);
or U1203 (N_1203,N_142,N_882);
xnor U1204 (N_1204,N_116,N_754);
nand U1205 (N_1205,N_480,N_871);
or U1206 (N_1206,N_559,N_627);
or U1207 (N_1207,N_416,N_730);
xnor U1208 (N_1208,N_400,N_938);
and U1209 (N_1209,N_601,N_438);
or U1210 (N_1210,N_222,N_245);
nand U1211 (N_1211,N_771,N_318);
nor U1212 (N_1212,N_663,N_861);
and U1213 (N_1213,N_946,N_464);
or U1214 (N_1214,N_163,N_866);
or U1215 (N_1215,N_575,N_49);
nand U1216 (N_1216,N_810,N_446);
or U1217 (N_1217,N_848,N_358);
nand U1218 (N_1218,N_390,N_5);
nor U1219 (N_1219,N_424,N_689);
nor U1220 (N_1220,N_571,N_175);
or U1221 (N_1221,N_27,N_539);
nor U1222 (N_1222,N_849,N_178);
nand U1223 (N_1223,N_393,N_429);
nor U1224 (N_1224,N_0,N_261);
nand U1225 (N_1225,N_739,N_780);
nand U1226 (N_1226,N_688,N_53);
nor U1227 (N_1227,N_115,N_352);
nand U1228 (N_1228,N_807,N_841);
or U1229 (N_1229,N_327,N_863);
xnor U1230 (N_1230,N_873,N_353);
or U1231 (N_1231,N_42,N_905);
or U1232 (N_1232,N_406,N_535);
nor U1233 (N_1233,N_607,N_652);
nand U1234 (N_1234,N_833,N_631);
and U1235 (N_1235,N_551,N_21);
nand U1236 (N_1236,N_350,N_896);
or U1237 (N_1237,N_883,N_408);
and U1238 (N_1238,N_592,N_790);
and U1239 (N_1239,N_25,N_440);
or U1240 (N_1240,N_215,N_303);
nor U1241 (N_1241,N_241,N_579);
and U1242 (N_1242,N_758,N_850);
and U1243 (N_1243,N_582,N_486);
nor U1244 (N_1244,N_453,N_553);
nor U1245 (N_1245,N_777,N_708);
nand U1246 (N_1246,N_840,N_294);
or U1247 (N_1247,N_521,N_309);
and U1248 (N_1248,N_153,N_704);
or U1249 (N_1249,N_624,N_969);
or U1250 (N_1250,N_910,N_532);
or U1251 (N_1251,N_767,N_939);
and U1252 (N_1252,N_40,N_638);
nor U1253 (N_1253,N_57,N_600);
nor U1254 (N_1254,N_6,N_827);
nand U1255 (N_1255,N_38,N_761);
nand U1256 (N_1256,N_591,N_705);
and U1257 (N_1257,N_948,N_786);
xnor U1258 (N_1258,N_944,N_545);
and U1259 (N_1259,N_597,N_211);
nor U1260 (N_1260,N_110,N_16);
or U1261 (N_1261,N_35,N_69);
or U1262 (N_1262,N_872,N_684);
or U1263 (N_1263,N_678,N_892);
and U1264 (N_1264,N_266,N_916);
nor U1265 (N_1265,N_485,N_593);
xor U1266 (N_1266,N_712,N_137);
nand U1267 (N_1267,N_297,N_447);
or U1268 (N_1268,N_44,N_993);
and U1269 (N_1269,N_699,N_46);
nor U1270 (N_1270,N_210,N_826);
or U1271 (N_1271,N_362,N_96);
or U1272 (N_1272,N_490,N_975);
nand U1273 (N_1273,N_964,N_441);
nor U1274 (N_1274,N_322,N_653);
nand U1275 (N_1275,N_615,N_753);
or U1276 (N_1276,N_346,N_626);
and U1277 (N_1277,N_795,N_515);
nor U1278 (N_1278,N_805,N_874);
nor U1279 (N_1279,N_128,N_221);
and U1280 (N_1280,N_355,N_320);
nor U1281 (N_1281,N_979,N_634);
nor U1282 (N_1282,N_864,N_425);
and U1283 (N_1283,N_568,N_457);
nand U1284 (N_1284,N_305,N_451);
and U1285 (N_1285,N_200,N_768);
and U1286 (N_1286,N_158,N_671);
or U1287 (N_1287,N_746,N_154);
and U1288 (N_1288,N_337,N_120);
nand U1289 (N_1289,N_243,N_630);
or U1290 (N_1290,N_621,N_919);
and U1291 (N_1291,N_804,N_275);
nand U1292 (N_1292,N_126,N_419);
nor U1293 (N_1293,N_454,N_77);
nand U1294 (N_1294,N_585,N_458);
nand U1295 (N_1295,N_973,N_931);
or U1296 (N_1296,N_963,N_994);
or U1297 (N_1297,N_875,N_236);
and U1298 (N_1298,N_491,N_461);
and U1299 (N_1299,N_844,N_196);
or U1300 (N_1300,N_264,N_317);
nor U1301 (N_1301,N_886,N_752);
or U1302 (N_1302,N_363,N_516);
nand U1303 (N_1303,N_925,N_66);
nor U1304 (N_1304,N_527,N_959);
nand U1305 (N_1305,N_155,N_456);
nand U1306 (N_1306,N_176,N_455);
nand U1307 (N_1307,N_161,N_732);
or U1308 (N_1308,N_382,N_978);
nand U1309 (N_1309,N_555,N_300);
and U1310 (N_1310,N_576,N_102);
nor U1311 (N_1311,N_714,N_36);
xor U1312 (N_1312,N_765,N_731);
or U1313 (N_1313,N_148,N_383);
and U1314 (N_1314,N_596,N_52);
nor U1315 (N_1315,N_229,N_683);
nor U1316 (N_1316,N_983,N_958);
or U1317 (N_1317,N_445,N_865);
or U1318 (N_1318,N_138,N_847);
nor U1319 (N_1319,N_835,N_404);
nor U1320 (N_1320,N_722,N_473);
and U1321 (N_1321,N_367,N_470);
nor U1322 (N_1322,N_59,N_342);
or U1323 (N_1323,N_736,N_988);
nand U1324 (N_1324,N_985,N_815);
and U1325 (N_1325,N_481,N_504);
nand U1326 (N_1326,N_907,N_726);
or U1327 (N_1327,N_140,N_718);
or U1328 (N_1328,N_418,N_530);
nor U1329 (N_1329,N_524,N_862);
and U1330 (N_1330,N_723,N_748);
and U1331 (N_1331,N_323,N_288);
or U1332 (N_1332,N_537,N_427);
or U1333 (N_1333,N_78,N_310);
and U1334 (N_1334,N_179,N_558);
and U1335 (N_1335,N_991,N_656);
nor U1336 (N_1336,N_307,N_703);
nor U1337 (N_1337,N_10,N_331);
or U1338 (N_1338,N_740,N_735);
nand U1339 (N_1339,N_58,N_208);
xor U1340 (N_1340,N_250,N_312);
or U1341 (N_1341,N_513,N_823);
xnor U1342 (N_1342,N_728,N_669);
or U1343 (N_1343,N_282,N_505);
or U1344 (N_1344,N_407,N_962);
or U1345 (N_1345,N_373,N_838);
and U1346 (N_1346,N_673,N_341);
nand U1347 (N_1347,N_272,N_572);
or U1348 (N_1348,N_313,N_519);
or U1349 (N_1349,N_824,N_930);
and U1350 (N_1350,N_583,N_750);
and U1351 (N_1351,N_316,N_15);
nand U1352 (N_1352,N_654,N_325);
nor U1353 (N_1353,N_388,N_552);
nor U1354 (N_1354,N_598,N_560);
or U1355 (N_1355,N_876,N_543);
nor U1356 (N_1356,N_436,N_729);
and U1357 (N_1357,N_114,N_613);
and U1358 (N_1358,N_324,N_60);
nand U1359 (N_1359,N_45,N_937);
or U1360 (N_1360,N_377,N_672);
and U1361 (N_1361,N_661,N_33);
nand U1362 (N_1362,N_83,N_644);
and U1363 (N_1363,N_717,N_725);
or U1364 (N_1364,N_145,N_614);
or U1365 (N_1365,N_898,N_281);
nand U1366 (N_1366,N_589,N_257);
nand U1367 (N_1367,N_106,N_566);
nand U1368 (N_1368,N_563,N_943);
and U1369 (N_1369,N_526,N_759);
nand U1370 (N_1370,N_2,N_666);
or U1371 (N_1371,N_174,N_700);
and U1372 (N_1372,N_193,N_375);
nand U1373 (N_1373,N_595,N_647);
or U1374 (N_1374,N_974,N_117);
xnor U1375 (N_1375,N_812,N_997);
xor U1376 (N_1376,N_201,N_640);
nand U1377 (N_1377,N_319,N_321);
and U1378 (N_1378,N_448,N_747);
nand U1379 (N_1379,N_97,N_214);
or U1380 (N_1380,N_577,N_73);
nand U1381 (N_1381,N_190,N_858);
nand U1382 (N_1382,N_213,N_8);
or U1383 (N_1383,N_244,N_928);
or U1384 (N_1384,N_622,N_412);
nand U1385 (N_1385,N_784,N_680);
or U1386 (N_1386,N_608,N_749);
or U1387 (N_1387,N_239,N_70);
nand U1388 (N_1388,N_965,N_430);
nand U1389 (N_1389,N_742,N_285);
nand U1390 (N_1390,N_356,N_139);
or U1391 (N_1391,N_85,N_56);
nor U1392 (N_1392,N_450,N_354);
nor U1393 (N_1393,N_745,N_967);
nor U1394 (N_1394,N_894,N_676);
and U1395 (N_1395,N_904,N_950);
nor U1396 (N_1396,N_224,N_554);
nor U1397 (N_1397,N_156,N_851);
nand U1398 (N_1398,N_255,N_842);
nor U1399 (N_1399,N_550,N_437);
nor U1400 (N_1400,N_141,N_920);
or U1401 (N_1401,N_366,N_468);
nand U1402 (N_1402,N_143,N_623);
nor U1403 (N_1403,N_884,N_562);
nor U1404 (N_1404,N_693,N_711);
and U1405 (N_1405,N_778,N_286);
or U1406 (N_1406,N_217,N_258);
nor U1407 (N_1407,N_911,N_417);
or U1408 (N_1408,N_534,N_129);
and U1409 (N_1409,N_738,N_977);
nor U1410 (N_1410,N_89,N_879);
or U1411 (N_1411,N_387,N_62);
nand U1412 (N_1412,N_248,N_751);
xnor U1413 (N_1413,N_970,N_877);
nand U1414 (N_1414,N_401,N_384);
or U1415 (N_1415,N_1,N_506);
and U1416 (N_1416,N_428,N_932);
nand U1417 (N_1417,N_466,N_442);
nand U1418 (N_1418,N_67,N_397);
nor U1419 (N_1419,N_463,N_209);
nor U1420 (N_1420,N_668,N_144);
nand U1421 (N_1421,N_870,N_690);
nor U1422 (N_1422,N_270,N_479);
or U1423 (N_1423,N_192,N_198);
nor U1424 (N_1424,N_162,N_31);
nor U1425 (N_1425,N_776,N_177);
nor U1426 (N_1426,N_633,N_423);
nand U1427 (N_1427,N_695,N_80);
or U1428 (N_1428,N_105,N_854);
and U1429 (N_1429,N_665,N_132);
nor U1430 (N_1430,N_95,N_947);
nor U1431 (N_1431,N_379,N_386);
and U1432 (N_1432,N_376,N_533);
and U1433 (N_1433,N_957,N_679);
and U1434 (N_1434,N_471,N_800);
nand U1435 (N_1435,N_825,N_498);
nor U1436 (N_1436,N_111,N_296);
or U1437 (N_1437,N_893,N_936);
nand U1438 (N_1438,N_314,N_371);
nor U1439 (N_1439,N_821,N_469);
nand U1440 (N_1440,N_832,N_642);
or U1441 (N_1441,N_169,N_940);
and U1442 (N_1442,N_333,N_971);
and U1443 (N_1443,N_834,N_340);
nor U1444 (N_1444,N_828,N_536);
and U1445 (N_1445,N_287,N_637);
and U1446 (N_1446,N_329,N_183);
and U1447 (N_1447,N_618,N_677);
or U1448 (N_1448,N_113,N_399);
nor U1449 (N_1449,N_580,N_831);
or U1450 (N_1450,N_869,N_410);
nand U1451 (N_1451,N_658,N_788);
nand U1452 (N_1452,N_259,N_540);
xor U1453 (N_1453,N_646,N_829);
and U1454 (N_1454,N_701,N_99);
nand U1455 (N_1455,N_510,N_707);
or U1456 (N_1456,N_692,N_913);
and U1457 (N_1457,N_394,N_667);
nor U1458 (N_1458,N_629,N_885);
and U1459 (N_1459,N_603,N_334);
or U1460 (N_1460,N_783,N_277);
nand U1461 (N_1461,N_954,N_18);
xor U1462 (N_1462,N_119,N_100);
nor U1463 (N_1463,N_594,N_956);
or U1464 (N_1464,N_344,N_289);
nand U1465 (N_1465,N_741,N_444);
nor U1466 (N_1466,N_433,N_682);
nand U1467 (N_1467,N_109,N_9);
nand U1468 (N_1468,N_361,N_202);
or U1469 (N_1469,N_32,N_792);
nand U1470 (N_1470,N_167,N_528);
and U1471 (N_1471,N_395,N_620);
or U1472 (N_1472,N_197,N_547);
nor U1473 (N_1473,N_232,N_687);
nor U1474 (N_1474,N_149,N_512);
or U1475 (N_1475,N_147,N_41);
nor U1476 (N_1476,N_68,N_475);
nand U1477 (N_1477,N_522,N_207);
or U1478 (N_1478,N_744,N_225);
or U1479 (N_1479,N_411,N_435);
or U1480 (N_1480,N_497,N_7);
nand U1481 (N_1481,N_268,N_86);
or U1482 (N_1482,N_719,N_924);
and U1483 (N_1483,N_187,N_72);
or U1484 (N_1484,N_499,N_372);
or U1485 (N_1485,N_782,N_611);
nand U1486 (N_1486,N_606,N_502);
xor U1487 (N_1487,N_84,N_168);
and U1488 (N_1488,N_650,N_972);
and U1489 (N_1489,N_186,N_304);
and U1490 (N_1490,N_28,N_918);
nand U1491 (N_1491,N_13,N_124);
and U1492 (N_1492,N_517,N_234);
or U1493 (N_1493,N_151,N_173);
or U1494 (N_1494,N_269,N_452);
or U1495 (N_1495,N_995,N_216);
and U1496 (N_1496,N_890,N_906);
nand U1497 (N_1497,N_459,N_291);
nor U1498 (N_1498,N_830,N_734);
nand U1499 (N_1499,N_460,N_184);
nor U1500 (N_1500,N_2,N_411);
nor U1501 (N_1501,N_733,N_697);
or U1502 (N_1502,N_790,N_529);
nor U1503 (N_1503,N_952,N_931);
or U1504 (N_1504,N_116,N_88);
or U1505 (N_1505,N_826,N_513);
and U1506 (N_1506,N_546,N_358);
or U1507 (N_1507,N_14,N_527);
or U1508 (N_1508,N_986,N_230);
nor U1509 (N_1509,N_475,N_640);
nand U1510 (N_1510,N_946,N_802);
or U1511 (N_1511,N_114,N_876);
or U1512 (N_1512,N_539,N_830);
or U1513 (N_1513,N_1,N_373);
nand U1514 (N_1514,N_528,N_742);
nor U1515 (N_1515,N_232,N_855);
and U1516 (N_1516,N_288,N_642);
nor U1517 (N_1517,N_71,N_363);
or U1518 (N_1518,N_303,N_942);
and U1519 (N_1519,N_684,N_383);
and U1520 (N_1520,N_163,N_578);
or U1521 (N_1521,N_330,N_709);
nor U1522 (N_1522,N_780,N_837);
nand U1523 (N_1523,N_909,N_344);
or U1524 (N_1524,N_585,N_938);
or U1525 (N_1525,N_797,N_577);
nand U1526 (N_1526,N_546,N_562);
and U1527 (N_1527,N_826,N_823);
or U1528 (N_1528,N_426,N_130);
and U1529 (N_1529,N_867,N_522);
nor U1530 (N_1530,N_802,N_957);
or U1531 (N_1531,N_821,N_869);
or U1532 (N_1532,N_506,N_787);
nand U1533 (N_1533,N_46,N_763);
xnor U1534 (N_1534,N_610,N_663);
and U1535 (N_1535,N_872,N_168);
or U1536 (N_1536,N_395,N_830);
and U1537 (N_1537,N_926,N_590);
and U1538 (N_1538,N_499,N_617);
and U1539 (N_1539,N_780,N_999);
and U1540 (N_1540,N_246,N_974);
nand U1541 (N_1541,N_442,N_181);
or U1542 (N_1542,N_959,N_700);
nor U1543 (N_1543,N_981,N_677);
or U1544 (N_1544,N_2,N_393);
and U1545 (N_1545,N_464,N_212);
nand U1546 (N_1546,N_118,N_84);
or U1547 (N_1547,N_541,N_577);
or U1548 (N_1548,N_145,N_764);
or U1549 (N_1549,N_493,N_242);
and U1550 (N_1550,N_138,N_211);
and U1551 (N_1551,N_57,N_256);
nand U1552 (N_1552,N_182,N_220);
and U1553 (N_1553,N_452,N_696);
or U1554 (N_1554,N_510,N_166);
or U1555 (N_1555,N_836,N_849);
or U1556 (N_1556,N_182,N_712);
and U1557 (N_1557,N_919,N_398);
and U1558 (N_1558,N_262,N_68);
or U1559 (N_1559,N_186,N_864);
and U1560 (N_1560,N_521,N_435);
or U1561 (N_1561,N_290,N_991);
nor U1562 (N_1562,N_26,N_208);
or U1563 (N_1563,N_665,N_789);
or U1564 (N_1564,N_336,N_484);
and U1565 (N_1565,N_202,N_981);
or U1566 (N_1566,N_471,N_768);
xnor U1567 (N_1567,N_879,N_979);
nand U1568 (N_1568,N_650,N_342);
nand U1569 (N_1569,N_342,N_684);
nand U1570 (N_1570,N_516,N_255);
or U1571 (N_1571,N_330,N_841);
nor U1572 (N_1572,N_237,N_943);
or U1573 (N_1573,N_385,N_166);
or U1574 (N_1574,N_160,N_545);
or U1575 (N_1575,N_1,N_677);
nand U1576 (N_1576,N_313,N_763);
nor U1577 (N_1577,N_925,N_705);
nand U1578 (N_1578,N_170,N_487);
nand U1579 (N_1579,N_557,N_261);
nand U1580 (N_1580,N_66,N_102);
nand U1581 (N_1581,N_149,N_749);
or U1582 (N_1582,N_4,N_57);
and U1583 (N_1583,N_227,N_783);
or U1584 (N_1584,N_948,N_959);
xnor U1585 (N_1585,N_494,N_988);
and U1586 (N_1586,N_165,N_820);
or U1587 (N_1587,N_599,N_795);
nor U1588 (N_1588,N_246,N_984);
or U1589 (N_1589,N_108,N_409);
and U1590 (N_1590,N_180,N_421);
xor U1591 (N_1591,N_577,N_170);
nand U1592 (N_1592,N_242,N_743);
nor U1593 (N_1593,N_312,N_3);
nor U1594 (N_1594,N_753,N_461);
xnor U1595 (N_1595,N_378,N_614);
and U1596 (N_1596,N_912,N_499);
or U1597 (N_1597,N_707,N_511);
and U1598 (N_1598,N_68,N_461);
or U1599 (N_1599,N_341,N_656);
and U1600 (N_1600,N_454,N_148);
xnor U1601 (N_1601,N_382,N_311);
and U1602 (N_1602,N_821,N_815);
nor U1603 (N_1603,N_272,N_923);
or U1604 (N_1604,N_659,N_60);
nor U1605 (N_1605,N_73,N_484);
or U1606 (N_1606,N_272,N_241);
and U1607 (N_1607,N_829,N_663);
xnor U1608 (N_1608,N_807,N_915);
and U1609 (N_1609,N_695,N_244);
nor U1610 (N_1610,N_942,N_664);
nor U1611 (N_1611,N_401,N_992);
and U1612 (N_1612,N_463,N_319);
nand U1613 (N_1613,N_138,N_478);
and U1614 (N_1614,N_749,N_522);
xor U1615 (N_1615,N_446,N_842);
xnor U1616 (N_1616,N_250,N_39);
nand U1617 (N_1617,N_201,N_185);
nor U1618 (N_1618,N_569,N_639);
and U1619 (N_1619,N_732,N_705);
or U1620 (N_1620,N_815,N_937);
nor U1621 (N_1621,N_677,N_759);
or U1622 (N_1622,N_582,N_621);
nand U1623 (N_1623,N_506,N_12);
and U1624 (N_1624,N_17,N_182);
or U1625 (N_1625,N_265,N_462);
and U1626 (N_1626,N_229,N_56);
and U1627 (N_1627,N_504,N_943);
or U1628 (N_1628,N_16,N_143);
nor U1629 (N_1629,N_554,N_357);
nand U1630 (N_1630,N_485,N_380);
nand U1631 (N_1631,N_56,N_496);
nand U1632 (N_1632,N_14,N_431);
or U1633 (N_1633,N_483,N_198);
nor U1634 (N_1634,N_208,N_287);
and U1635 (N_1635,N_574,N_556);
nor U1636 (N_1636,N_460,N_592);
or U1637 (N_1637,N_220,N_993);
nand U1638 (N_1638,N_303,N_208);
nand U1639 (N_1639,N_460,N_383);
and U1640 (N_1640,N_940,N_762);
or U1641 (N_1641,N_857,N_590);
nand U1642 (N_1642,N_15,N_391);
and U1643 (N_1643,N_785,N_330);
and U1644 (N_1644,N_810,N_297);
or U1645 (N_1645,N_412,N_521);
nor U1646 (N_1646,N_918,N_865);
nor U1647 (N_1647,N_895,N_785);
and U1648 (N_1648,N_433,N_56);
or U1649 (N_1649,N_558,N_296);
nor U1650 (N_1650,N_519,N_30);
nand U1651 (N_1651,N_723,N_944);
xor U1652 (N_1652,N_421,N_709);
nand U1653 (N_1653,N_150,N_143);
or U1654 (N_1654,N_523,N_907);
nor U1655 (N_1655,N_266,N_648);
and U1656 (N_1656,N_385,N_947);
nor U1657 (N_1657,N_124,N_189);
and U1658 (N_1658,N_770,N_593);
xnor U1659 (N_1659,N_258,N_366);
and U1660 (N_1660,N_834,N_344);
nor U1661 (N_1661,N_954,N_352);
and U1662 (N_1662,N_170,N_836);
and U1663 (N_1663,N_984,N_739);
and U1664 (N_1664,N_568,N_928);
xor U1665 (N_1665,N_70,N_698);
nor U1666 (N_1666,N_800,N_94);
or U1667 (N_1667,N_72,N_990);
nand U1668 (N_1668,N_44,N_408);
nor U1669 (N_1669,N_173,N_154);
nand U1670 (N_1670,N_521,N_493);
or U1671 (N_1671,N_496,N_387);
nor U1672 (N_1672,N_723,N_403);
nand U1673 (N_1673,N_965,N_984);
nor U1674 (N_1674,N_154,N_451);
nand U1675 (N_1675,N_214,N_401);
or U1676 (N_1676,N_735,N_244);
nand U1677 (N_1677,N_94,N_134);
and U1678 (N_1678,N_786,N_231);
and U1679 (N_1679,N_347,N_758);
nand U1680 (N_1680,N_728,N_493);
and U1681 (N_1681,N_744,N_147);
nor U1682 (N_1682,N_147,N_870);
nor U1683 (N_1683,N_816,N_933);
and U1684 (N_1684,N_824,N_279);
nor U1685 (N_1685,N_500,N_827);
and U1686 (N_1686,N_549,N_874);
and U1687 (N_1687,N_233,N_938);
and U1688 (N_1688,N_98,N_424);
and U1689 (N_1689,N_210,N_232);
and U1690 (N_1690,N_588,N_923);
and U1691 (N_1691,N_634,N_875);
or U1692 (N_1692,N_178,N_661);
nor U1693 (N_1693,N_646,N_22);
or U1694 (N_1694,N_974,N_127);
or U1695 (N_1695,N_647,N_986);
nand U1696 (N_1696,N_576,N_383);
nand U1697 (N_1697,N_367,N_603);
nor U1698 (N_1698,N_938,N_506);
xnor U1699 (N_1699,N_349,N_325);
or U1700 (N_1700,N_552,N_768);
and U1701 (N_1701,N_905,N_641);
or U1702 (N_1702,N_571,N_357);
nor U1703 (N_1703,N_755,N_668);
and U1704 (N_1704,N_440,N_903);
and U1705 (N_1705,N_876,N_488);
or U1706 (N_1706,N_699,N_166);
and U1707 (N_1707,N_91,N_449);
and U1708 (N_1708,N_924,N_301);
nor U1709 (N_1709,N_727,N_238);
nor U1710 (N_1710,N_30,N_853);
or U1711 (N_1711,N_274,N_339);
nor U1712 (N_1712,N_888,N_32);
nor U1713 (N_1713,N_749,N_19);
nand U1714 (N_1714,N_73,N_611);
and U1715 (N_1715,N_544,N_387);
and U1716 (N_1716,N_837,N_880);
and U1717 (N_1717,N_692,N_881);
and U1718 (N_1718,N_400,N_7);
and U1719 (N_1719,N_203,N_383);
nand U1720 (N_1720,N_101,N_699);
or U1721 (N_1721,N_376,N_839);
and U1722 (N_1722,N_97,N_948);
or U1723 (N_1723,N_308,N_381);
or U1724 (N_1724,N_762,N_867);
or U1725 (N_1725,N_788,N_422);
and U1726 (N_1726,N_555,N_341);
and U1727 (N_1727,N_36,N_145);
nand U1728 (N_1728,N_795,N_826);
nand U1729 (N_1729,N_108,N_669);
or U1730 (N_1730,N_538,N_573);
nor U1731 (N_1731,N_409,N_519);
and U1732 (N_1732,N_608,N_213);
or U1733 (N_1733,N_136,N_276);
nand U1734 (N_1734,N_960,N_791);
and U1735 (N_1735,N_821,N_763);
or U1736 (N_1736,N_760,N_699);
nand U1737 (N_1737,N_779,N_557);
nand U1738 (N_1738,N_787,N_279);
and U1739 (N_1739,N_428,N_802);
nand U1740 (N_1740,N_768,N_450);
nand U1741 (N_1741,N_948,N_365);
xor U1742 (N_1742,N_427,N_681);
or U1743 (N_1743,N_603,N_899);
or U1744 (N_1744,N_853,N_888);
nor U1745 (N_1745,N_947,N_369);
or U1746 (N_1746,N_679,N_652);
and U1747 (N_1747,N_882,N_163);
and U1748 (N_1748,N_347,N_124);
nand U1749 (N_1749,N_374,N_1);
nor U1750 (N_1750,N_460,N_918);
and U1751 (N_1751,N_108,N_428);
nand U1752 (N_1752,N_755,N_474);
and U1753 (N_1753,N_446,N_489);
nor U1754 (N_1754,N_426,N_834);
and U1755 (N_1755,N_534,N_994);
nand U1756 (N_1756,N_443,N_847);
nand U1757 (N_1757,N_271,N_746);
or U1758 (N_1758,N_856,N_157);
and U1759 (N_1759,N_907,N_675);
nand U1760 (N_1760,N_760,N_640);
nor U1761 (N_1761,N_626,N_464);
nand U1762 (N_1762,N_999,N_479);
nand U1763 (N_1763,N_457,N_793);
or U1764 (N_1764,N_657,N_730);
and U1765 (N_1765,N_959,N_955);
nand U1766 (N_1766,N_12,N_435);
or U1767 (N_1767,N_594,N_897);
nor U1768 (N_1768,N_444,N_451);
and U1769 (N_1769,N_901,N_755);
nor U1770 (N_1770,N_459,N_302);
and U1771 (N_1771,N_406,N_542);
and U1772 (N_1772,N_185,N_147);
nand U1773 (N_1773,N_913,N_208);
or U1774 (N_1774,N_189,N_690);
or U1775 (N_1775,N_489,N_228);
nor U1776 (N_1776,N_111,N_249);
and U1777 (N_1777,N_79,N_241);
and U1778 (N_1778,N_969,N_920);
or U1779 (N_1779,N_880,N_532);
or U1780 (N_1780,N_937,N_544);
nor U1781 (N_1781,N_610,N_579);
xnor U1782 (N_1782,N_273,N_478);
or U1783 (N_1783,N_120,N_423);
nor U1784 (N_1784,N_671,N_13);
nor U1785 (N_1785,N_663,N_601);
nor U1786 (N_1786,N_429,N_924);
nor U1787 (N_1787,N_38,N_314);
and U1788 (N_1788,N_106,N_140);
and U1789 (N_1789,N_461,N_103);
and U1790 (N_1790,N_601,N_24);
nand U1791 (N_1791,N_348,N_42);
and U1792 (N_1792,N_345,N_505);
and U1793 (N_1793,N_877,N_309);
nand U1794 (N_1794,N_789,N_479);
nor U1795 (N_1795,N_415,N_183);
or U1796 (N_1796,N_300,N_700);
nor U1797 (N_1797,N_704,N_314);
nor U1798 (N_1798,N_883,N_719);
nor U1799 (N_1799,N_199,N_460);
and U1800 (N_1800,N_574,N_976);
or U1801 (N_1801,N_487,N_594);
and U1802 (N_1802,N_225,N_388);
and U1803 (N_1803,N_667,N_4);
and U1804 (N_1804,N_674,N_290);
nand U1805 (N_1805,N_969,N_808);
nand U1806 (N_1806,N_98,N_126);
xor U1807 (N_1807,N_666,N_148);
nand U1808 (N_1808,N_656,N_273);
xnor U1809 (N_1809,N_746,N_334);
and U1810 (N_1810,N_689,N_591);
nor U1811 (N_1811,N_72,N_461);
nand U1812 (N_1812,N_530,N_372);
or U1813 (N_1813,N_787,N_134);
nand U1814 (N_1814,N_155,N_351);
nor U1815 (N_1815,N_71,N_465);
and U1816 (N_1816,N_207,N_926);
nand U1817 (N_1817,N_54,N_663);
and U1818 (N_1818,N_229,N_933);
and U1819 (N_1819,N_273,N_584);
nand U1820 (N_1820,N_930,N_586);
and U1821 (N_1821,N_373,N_238);
or U1822 (N_1822,N_482,N_551);
nand U1823 (N_1823,N_225,N_330);
or U1824 (N_1824,N_619,N_221);
nand U1825 (N_1825,N_241,N_843);
or U1826 (N_1826,N_806,N_566);
nor U1827 (N_1827,N_617,N_181);
or U1828 (N_1828,N_989,N_350);
or U1829 (N_1829,N_838,N_213);
and U1830 (N_1830,N_995,N_91);
nor U1831 (N_1831,N_381,N_357);
and U1832 (N_1832,N_891,N_817);
or U1833 (N_1833,N_958,N_351);
or U1834 (N_1834,N_448,N_557);
nor U1835 (N_1835,N_62,N_514);
nand U1836 (N_1836,N_269,N_677);
nor U1837 (N_1837,N_291,N_125);
nor U1838 (N_1838,N_82,N_662);
or U1839 (N_1839,N_120,N_473);
nand U1840 (N_1840,N_257,N_325);
nand U1841 (N_1841,N_50,N_100);
nor U1842 (N_1842,N_152,N_120);
nor U1843 (N_1843,N_33,N_663);
or U1844 (N_1844,N_941,N_607);
nor U1845 (N_1845,N_966,N_81);
nor U1846 (N_1846,N_786,N_246);
nand U1847 (N_1847,N_580,N_506);
or U1848 (N_1848,N_288,N_891);
and U1849 (N_1849,N_42,N_431);
or U1850 (N_1850,N_569,N_391);
or U1851 (N_1851,N_250,N_499);
nand U1852 (N_1852,N_938,N_596);
nand U1853 (N_1853,N_308,N_655);
or U1854 (N_1854,N_288,N_570);
nor U1855 (N_1855,N_949,N_703);
nand U1856 (N_1856,N_810,N_62);
and U1857 (N_1857,N_118,N_462);
nor U1858 (N_1858,N_11,N_736);
nand U1859 (N_1859,N_907,N_883);
nand U1860 (N_1860,N_544,N_340);
and U1861 (N_1861,N_347,N_725);
nand U1862 (N_1862,N_579,N_870);
nor U1863 (N_1863,N_161,N_355);
and U1864 (N_1864,N_300,N_494);
nand U1865 (N_1865,N_853,N_504);
nand U1866 (N_1866,N_70,N_68);
nand U1867 (N_1867,N_741,N_365);
and U1868 (N_1868,N_615,N_913);
nor U1869 (N_1869,N_366,N_929);
or U1870 (N_1870,N_346,N_77);
nand U1871 (N_1871,N_329,N_862);
and U1872 (N_1872,N_788,N_642);
and U1873 (N_1873,N_849,N_283);
or U1874 (N_1874,N_345,N_518);
or U1875 (N_1875,N_892,N_297);
nor U1876 (N_1876,N_788,N_54);
or U1877 (N_1877,N_541,N_444);
nand U1878 (N_1878,N_62,N_143);
nand U1879 (N_1879,N_849,N_668);
nor U1880 (N_1880,N_123,N_468);
nor U1881 (N_1881,N_742,N_674);
and U1882 (N_1882,N_72,N_531);
nor U1883 (N_1883,N_949,N_69);
nor U1884 (N_1884,N_685,N_171);
and U1885 (N_1885,N_318,N_283);
and U1886 (N_1886,N_492,N_828);
and U1887 (N_1887,N_935,N_867);
and U1888 (N_1888,N_997,N_774);
and U1889 (N_1889,N_385,N_399);
nand U1890 (N_1890,N_668,N_801);
nand U1891 (N_1891,N_955,N_586);
or U1892 (N_1892,N_195,N_481);
nand U1893 (N_1893,N_287,N_961);
or U1894 (N_1894,N_725,N_901);
nor U1895 (N_1895,N_982,N_402);
and U1896 (N_1896,N_581,N_386);
or U1897 (N_1897,N_0,N_91);
nand U1898 (N_1898,N_874,N_614);
or U1899 (N_1899,N_830,N_332);
or U1900 (N_1900,N_609,N_729);
and U1901 (N_1901,N_947,N_615);
or U1902 (N_1902,N_834,N_685);
nor U1903 (N_1903,N_721,N_89);
nand U1904 (N_1904,N_308,N_931);
nor U1905 (N_1905,N_39,N_936);
and U1906 (N_1906,N_998,N_43);
and U1907 (N_1907,N_537,N_396);
nor U1908 (N_1908,N_731,N_552);
and U1909 (N_1909,N_26,N_373);
or U1910 (N_1910,N_728,N_651);
nand U1911 (N_1911,N_26,N_37);
nand U1912 (N_1912,N_870,N_546);
or U1913 (N_1913,N_694,N_520);
nand U1914 (N_1914,N_238,N_950);
or U1915 (N_1915,N_884,N_525);
nand U1916 (N_1916,N_4,N_382);
or U1917 (N_1917,N_109,N_170);
or U1918 (N_1918,N_724,N_766);
nand U1919 (N_1919,N_708,N_341);
and U1920 (N_1920,N_241,N_330);
nor U1921 (N_1921,N_74,N_488);
nand U1922 (N_1922,N_712,N_971);
nor U1923 (N_1923,N_796,N_342);
nor U1924 (N_1924,N_951,N_156);
nand U1925 (N_1925,N_731,N_668);
and U1926 (N_1926,N_320,N_684);
nand U1927 (N_1927,N_925,N_109);
xor U1928 (N_1928,N_980,N_831);
and U1929 (N_1929,N_137,N_637);
xor U1930 (N_1930,N_713,N_592);
nor U1931 (N_1931,N_434,N_800);
and U1932 (N_1932,N_927,N_941);
nor U1933 (N_1933,N_269,N_363);
nand U1934 (N_1934,N_27,N_33);
nand U1935 (N_1935,N_276,N_257);
nand U1936 (N_1936,N_620,N_171);
nor U1937 (N_1937,N_871,N_325);
or U1938 (N_1938,N_38,N_275);
or U1939 (N_1939,N_676,N_79);
nor U1940 (N_1940,N_805,N_817);
and U1941 (N_1941,N_949,N_495);
and U1942 (N_1942,N_691,N_852);
nor U1943 (N_1943,N_521,N_312);
or U1944 (N_1944,N_321,N_671);
or U1945 (N_1945,N_707,N_553);
and U1946 (N_1946,N_204,N_953);
and U1947 (N_1947,N_781,N_765);
nand U1948 (N_1948,N_99,N_479);
nor U1949 (N_1949,N_614,N_361);
and U1950 (N_1950,N_385,N_515);
nand U1951 (N_1951,N_474,N_21);
nand U1952 (N_1952,N_960,N_465);
nor U1953 (N_1953,N_981,N_214);
nand U1954 (N_1954,N_108,N_95);
xor U1955 (N_1955,N_912,N_132);
and U1956 (N_1956,N_897,N_925);
and U1957 (N_1957,N_324,N_566);
and U1958 (N_1958,N_626,N_412);
or U1959 (N_1959,N_673,N_296);
nor U1960 (N_1960,N_940,N_94);
or U1961 (N_1961,N_200,N_693);
xnor U1962 (N_1962,N_968,N_138);
nand U1963 (N_1963,N_383,N_477);
nor U1964 (N_1964,N_8,N_905);
nand U1965 (N_1965,N_64,N_276);
nor U1966 (N_1966,N_97,N_281);
and U1967 (N_1967,N_498,N_638);
nand U1968 (N_1968,N_313,N_679);
nor U1969 (N_1969,N_142,N_202);
nor U1970 (N_1970,N_714,N_670);
and U1971 (N_1971,N_915,N_299);
nor U1972 (N_1972,N_855,N_879);
and U1973 (N_1973,N_984,N_381);
nor U1974 (N_1974,N_61,N_159);
and U1975 (N_1975,N_726,N_584);
nor U1976 (N_1976,N_208,N_128);
and U1977 (N_1977,N_818,N_202);
nand U1978 (N_1978,N_337,N_286);
and U1979 (N_1979,N_364,N_678);
nand U1980 (N_1980,N_732,N_282);
nor U1981 (N_1981,N_462,N_99);
or U1982 (N_1982,N_836,N_620);
or U1983 (N_1983,N_515,N_637);
nor U1984 (N_1984,N_263,N_534);
and U1985 (N_1985,N_663,N_613);
xor U1986 (N_1986,N_103,N_366);
and U1987 (N_1987,N_412,N_192);
and U1988 (N_1988,N_133,N_926);
and U1989 (N_1989,N_284,N_237);
nand U1990 (N_1990,N_905,N_279);
or U1991 (N_1991,N_256,N_366);
nor U1992 (N_1992,N_1,N_973);
and U1993 (N_1993,N_741,N_230);
nor U1994 (N_1994,N_204,N_610);
nand U1995 (N_1995,N_328,N_906);
and U1996 (N_1996,N_761,N_83);
and U1997 (N_1997,N_815,N_290);
or U1998 (N_1998,N_310,N_751);
nand U1999 (N_1999,N_670,N_876);
nor U2000 (N_2000,N_1081,N_1887);
and U2001 (N_2001,N_1771,N_1387);
nand U2002 (N_2002,N_1686,N_1230);
and U2003 (N_2003,N_1051,N_1216);
and U2004 (N_2004,N_1228,N_1790);
or U2005 (N_2005,N_1429,N_1473);
nor U2006 (N_2006,N_1733,N_1402);
nor U2007 (N_2007,N_1021,N_1439);
or U2008 (N_2008,N_1368,N_1546);
or U2009 (N_2009,N_1743,N_1883);
nor U2010 (N_2010,N_1851,N_1132);
nor U2011 (N_2011,N_1991,N_1122);
nor U2012 (N_2012,N_1826,N_1447);
nor U2013 (N_2013,N_1240,N_1719);
nor U2014 (N_2014,N_1443,N_1938);
or U2015 (N_2015,N_1983,N_1406);
nand U2016 (N_2016,N_1629,N_1695);
or U2017 (N_2017,N_1805,N_1982);
nand U2018 (N_2018,N_1974,N_1811);
xor U2019 (N_2019,N_1188,N_1166);
or U2020 (N_2020,N_1277,N_1403);
nor U2021 (N_2021,N_1264,N_1137);
xnor U2022 (N_2022,N_1547,N_1509);
or U2023 (N_2023,N_1322,N_1298);
nand U2024 (N_2024,N_1342,N_1888);
and U2025 (N_2025,N_1241,N_1693);
and U2026 (N_2026,N_1442,N_1504);
nor U2027 (N_2027,N_1126,N_1287);
nand U2028 (N_2028,N_1049,N_1248);
or U2029 (N_2029,N_1223,N_1857);
and U2030 (N_2030,N_1393,N_1476);
nand U2031 (N_2031,N_1966,N_1191);
nand U2032 (N_2032,N_1142,N_1963);
nand U2033 (N_2033,N_1704,N_1086);
and U2034 (N_2034,N_1478,N_1906);
nor U2035 (N_2035,N_1979,N_1315);
nand U2036 (N_2036,N_1975,N_1925);
or U2037 (N_2037,N_1233,N_1998);
or U2038 (N_2038,N_1073,N_1921);
and U2039 (N_2039,N_1259,N_1506);
or U2040 (N_2040,N_1532,N_1929);
and U2041 (N_2041,N_1076,N_1734);
xor U2042 (N_2042,N_1184,N_1459);
nor U2043 (N_2043,N_1108,N_1808);
xnor U2044 (N_2044,N_1167,N_1822);
nand U2045 (N_2045,N_1356,N_1384);
and U2046 (N_2046,N_1720,N_1499);
or U2047 (N_2047,N_1041,N_1838);
and U2048 (N_2048,N_1551,N_1242);
nor U2049 (N_2049,N_1033,N_1112);
or U2050 (N_2050,N_1934,N_1067);
nor U2051 (N_2051,N_1605,N_1915);
or U2052 (N_2052,N_1467,N_1084);
or U2053 (N_2053,N_1454,N_1872);
and U2054 (N_2054,N_1080,N_1622);
nor U2055 (N_2055,N_1463,N_1903);
nand U2056 (N_2056,N_1489,N_1369);
and U2057 (N_2057,N_1669,N_1363);
nand U2058 (N_2058,N_1200,N_1405);
nor U2059 (N_2059,N_1958,N_1683);
nor U2060 (N_2060,N_1993,N_1741);
and U2061 (N_2061,N_1578,N_1125);
nor U2062 (N_2062,N_1965,N_1378);
or U2063 (N_2063,N_1057,N_1954);
and U2064 (N_2064,N_1528,N_1092);
or U2065 (N_2065,N_1477,N_1799);
or U2066 (N_2066,N_1005,N_1470);
nor U2067 (N_2067,N_1088,N_1381);
or U2068 (N_2068,N_1135,N_1791);
nand U2069 (N_2069,N_1428,N_1379);
nor U2070 (N_2070,N_1948,N_1449);
nand U2071 (N_2071,N_1918,N_1786);
and U2072 (N_2072,N_1770,N_1762);
and U2073 (N_2073,N_1254,N_1004);
or U2074 (N_2074,N_1920,N_1329);
nor U2075 (N_2075,N_1909,N_1845);
nor U2076 (N_2076,N_1019,N_1174);
nand U2077 (N_2077,N_1562,N_1425);
or U2078 (N_2078,N_1859,N_1612);
and U2079 (N_2079,N_1222,N_1272);
nand U2080 (N_2080,N_1468,N_1064);
nor U2081 (N_2081,N_1761,N_1989);
nor U2082 (N_2082,N_1224,N_1995);
nor U2083 (N_2083,N_1904,N_1022);
nor U2084 (N_2084,N_1392,N_1655);
or U2085 (N_2085,N_1816,N_1214);
nor U2086 (N_2086,N_1875,N_1853);
nor U2087 (N_2087,N_1318,N_1246);
nor U2088 (N_2088,N_1830,N_1910);
nand U2089 (N_2089,N_1261,N_1818);
or U2090 (N_2090,N_1139,N_1658);
nand U2091 (N_2091,N_1037,N_1731);
or U2092 (N_2092,N_1180,N_1056);
and U2093 (N_2093,N_1945,N_1210);
or U2094 (N_2094,N_1611,N_1810);
nor U2095 (N_2095,N_1120,N_1623);
nand U2096 (N_2096,N_1131,N_1855);
nand U2097 (N_2097,N_1351,N_1967);
or U2098 (N_2098,N_1335,N_1557);
nand U2099 (N_2099,N_1708,N_1435);
nor U2100 (N_2100,N_1419,N_1821);
and U2101 (N_2101,N_1415,N_1919);
nand U2102 (N_2102,N_1644,N_1880);
or U2103 (N_2103,N_1176,N_1118);
nor U2104 (N_2104,N_1332,N_1577);
nor U2105 (N_2105,N_1520,N_1990);
nor U2106 (N_2106,N_1837,N_1981);
nor U2107 (N_2107,N_1777,N_1508);
nor U2108 (N_2108,N_1692,N_1484);
or U2109 (N_2109,N_1978,N_1048);
nor U2110 (N_2110,N_1186,N_1373);
or U2111 (N_2111,N_1939,N_1098);
nor U2112 (N_2112,N_1573,N_1097);
and U2113 (N_2113,N_1687,N_1788);
or U2114 (N_2114,N_1642,N_1987);
nor U2115 (N_2115,N_1685,N_1533);
nand U2116 (N_2116,N_1712,N_1030);
nor U2117 (N_2117,N_1452,N_1999);
nor U2118 (N_2118,N_1221,N_1566);
and U2119 (N_2119,N_1289,N_1050);
nor U2120 (N_2120,N_1568,N_1581);
nor U2121 (N_2121,N_1785,N_1197);
nand U2122 (N_2122,N_1996,N_1699);
or U2123 (N_2123,N_1119,N_1728);
or U2124 (N_2124,N_1827,N_1388);
or U2125 (N_2125,N_1215,N_1521);
and U2126 (N_2126,N_1279,N_1608);
or U2127 (N_2127,N_1992,N_1794);
or U2128 (N_2128,N_1595,N_1420);
nor U2129 (N_2129,N_1410,N_1867);
nor U2130 (N_2130,N_1278,N_1597);
nand U2131 (N_2131,N_1614,N_1359);
nand U2132 (N_2132,N_1681,N_1072);
nand U2133 (N_2133,N_1040,N_1481);
and U2134 (N_2134,N_1012,N_1198);
or U2135 (N_2135,N_1778,N_1907);
nand U2136 (N_2136,N_1326,N_1361);
nand U2137 (N_2137,N_1567,N_1475);
and U2138 (N_2138,N_1783,N_1205);
and U2139 (N_2139,N_1678,N_1976);
or U2140 (N_2140,N_1294,N_1878);
or U2141 (N_2141,N_1571,N_1398);
or U2142 (N_2142,N_1781,N_1396);
nor U2143 (N_2143,N_1700,N_1601);
nand U2144 (N_2144,N_1657,N_1663);
or U2145 (N_2145,N_1061,N_1864);
and U2146 (N_2146,N_1631,N_1769);
nand U2147 (N_2147,N_1703,N_1923);
nand U2148 (N_2148,N_1090,N_1169);
nand U2149 (N_2149,N_1065,N_1645);
and U2150 (N_2150,N_1480,N_1354);
nand U2151 (N_2151,N_1353,N_1212);
nand U2152 (N_2152,N_1260,N_1150);
or U2153 (N_2153,N_1134,N_1313);
or U2154 (N_2154,N_1082,N_1649);
and U2155 (N_2155,N_1936,N_1209);
nor U2156 (N_2156,N_1213,N_1576);
nor U2157 (N_2157,N_1181,N_1997);
nand U2158 (N_2158,N_1102,N_1660);
nor U2159 (N_2159,N_1165,N_1170);
or U2160 (N_2160,N_1091,N_1764);
or U2161 (N_2161,N_1431,N_1927);
or U2162 (N_2162,N_1585,N_1421);
nand U2163 (N_2163,N_1665,N_1854);
nand U2164 (N_2164,N_1025,N_1691);
nor U2165 (N_2165,N_1549,N_1579);
and U2166 (N_2166,N_1311,N_1063);
nand U2167 (N_2167,N_1324,N_1862);
or U2168 (N_2168,N_1479,N_1148);
and U2169 (N_2169,N_1232,N_1304);
and U2170 (N_2170,N_1413,N_1599);
nor U2171 (N_2171,N_1362,N_1894);
and U2172 (N_2172,N_1843,N_1121);
nor U2173 (N_2173,N_1606,N_1164);
nor U2174 (N_2174,N_1714,N_1423);
or U2175 (N_2175,N_1574,N_1942);
nor U2176 (N_2176,N_1059,N_1775);
nand U2177 (N_2177,N_1806,N_1582);
and U2178 (N_2178,N_1451,N_1625);
or U2179 (N_2179,N_1801,N_1895);
and U2180 (N_2180,N_1675,N_1231);
nor U2181 (N_2181,N_1236,N_1107);
and U2182 (N_2182,N_1093,N_1196);
or U2183 (N_2183,N_1116,N_1671);
nor U2184 (N_2184,N_1530,N_1971);
nand U2185 (N_2185,N_1609,N_1834);
and U2186 (N_2186,N_1793,N_1969);
or U2187 (N_2187,N_1245,N_1548);
nand U2188 (N_2188,N_1662,N_1627);
and U2189 (N_2189,N_1738,N_1905);
nor U2190 (N_2190,N_1094,N_1994);
nor U2191 (N_2191,N_1074,N_1517);
nor U2192 (N_2192,N_1580,N_1271);
nor U2193 (N_2193,N_1512,N_1058);
nor U2194 (N_2194,N_1901,N_1234);
or U2195 (N_2195,N_1346,N_1865);
nor U2196 (N_2196,N_1748,N_1697);
or U2197 (N_2197,N_1679,N_1220);
nor U2198 (N_2198,N_1953,N_1295);
nand U2199 (N_2199,N_1190,N_1676);
nor U2200 (N_2200,N_1427,N_1440);
nor U2201 (N_2201,N_1844,N_1177);
nor U2202 (N_2202,N_1010,N_1922);
and U2203 (N_2203,N_1251,N_1047);
or U2204 (N_2204,N_1607,N_1820);
and U2205 (N_2205,N_1239,N_1143);
nand U2206 (N_2206,N_1465,N_1879);
or U2207 (N_2207,N_1751,N_1485);
nor U2208 (N_2208,N_1858,N_1009);
nand U2209 (N_2209,N_1168,N_1670);
nand U2210 (N_2210,N_1195,N_1682);
or U2211 (N_2211,N_1096,N_1537);
or U2212 (N_2212,N_1270,N_1089);
xor U2213 (N_2213,N_1183,N_1229);
nand U2214 (N_2214,N_1302,N_1510);
and U2215 (N_2215,N_1444,N_1960);
nand U2216 (N_2216,N_1501,N_1062);
or U2217 (N_2217,N_1932,N_1407);
nor U2218 (N_2218,N_1244,N_1689);
nand U2219 (N_2219,N_1068,N_1727);
nand U2220 (N_2220,N_1390,N_1263);
or U2221 (N_2221,N_1587,N_1395);
nor U2222 (N_2222,N_1211,N_1000);
nor U2223 (N_2223,N_1598,N_1717);
and U2224 (N_2224,N_1552,N_1779);
nor U2225 (N_2225,N_1280,N_1747);
or U2226 (N_2226,N_1305,N_1737);
nor U2227 (N_2227,N_1760,N_1266);
or U2228 (N_2228,N_1924,N_1360);
or U2229 (N_2229,N_1060,N_1374);
nand U2230 (N_2230,N_1042,N_1491);
nand U2231 (N_2231,N_1284,N_1202);
nor U2232 (N_2232,N_1634,N_1839);
nor U2233 (N_2233,N_1255,N_1941);
and U2234 (N_2234,N_1647,N_1836);
nand U2235 (N_2235,N_1710,N_1896);
or U2236 (N_2236,N_1192,N_1653);
nand U2237 (N_2237,N_1620,N_1789);
or U2238 (N_2238,N_1952,N_1171);
or U2239 (N_2239,N_1648,N_1893);
nand U2240 (N_2240,N_1928,N_1558);
nand U2241 (N_2241,N_1123,N_1079);
nor U2242 (N_2242,N_1026,N_1028);
nor U2243 (N_2243,N_1153,N_1348);
nor U2244 (N_2244,N_1357,N_1201);
nand U2245 (N_2245,N_1926,N_1956);
and U2246 (N_2246,N_1798,N_1027);
or U2247 (N_2247,N_1460,N_1077);
nor U2248 (N_2248,N_1426,N_1654);
nor U2249 (N_2249,N_1172,N_1204);
nor U2250 (N_2250,N_1610,N_1055);
nor U2251 (N_2251,N_1268,N_1007);
nor U2252 (N_2252,N_1422,N_1561);
nand U2253 (N_2253,N_1591,N_1802);
or U2254 (N_2254,N_1225,N_1386);
nor U2255 (N_2255,N_1780,N_1603);
nand U2256 (N_2256,N_1265,N_1584);
and U2257 (N_2257,N_1039,N_1136);
nor U2258 (N_2258,N_1553,N_1105);
nand U2259 (N_2259,N_1618,N_1430);
xor U2260 (N_2260,N_1688,N_1312);
nor U2261 (N_2261,N_1933,N_1750);
nor U2262 (N_2262,N_1589,N_1564);
and U2263 (N_2263,N_1370,N_1588);
nor U2264 (N_2264,N_1519,N_1319);
nor U2265 (N_2265,N_1085,N_1293);
nand U2266 (N_2266,N_1950,N_1849);
or U2267 (N_2267,N_1711,N_1247);
nand U2268 (N_2268,N_1555,N_1626);
nand U2269 (N_2269,N_1876,N_1913);
nand U2270 (N_2270,N_1892,N_1227);
xnor U2271 (N_2271,N_1046,N_1970);
or U2272 (N_2272,N_1756,N_1029);
or U2273 (N_2273,N_1931,N_1513);
or U2274 (N_2274,N_1505,N_1035);
nand U2275 (N_2275,N_1621,N_1502);
nor U2276 (N_2276,N_1873,N_1514);
and U2277 (N_2277,N_1593,N_1371);
nand U2278 (N_2278,N_1759,N_1038);
or U2279 (N_2279,N_1095,N_1258);
nor U2280 (N_2280,N_1768,N_1943);
nand U2281 (N_2281,N_1382,N_1252);
or U2282 (N_2282,N_1902,N_1490);
and U2283 (N_2283,N_1389,N_1940);
nor U2284 (N_2284,N_1800,N_1643);
and U2285 (N_2285,N_1014,N_1487);
nor U2286 (N_2286,N_1968,N_1414);
or U2287 (N_2287,N_1526,N_1650);
nand U2288 (N_2288,N_1841,N_1848);
nand U2289 (N_2289,N_1453,N_1433);
xnor U2290 (N_2290,N_1787,N_1401);
nand U2291 (N_2291,N_1310,N_1736);
and U2292 (N_2292,N_1297,N_1666);
nor U2293 (N_2293,N_1937,N_1365);
nor U2294 (N_2294,N_1474,N_1347);
nand U2295 (N_2295,N_1912,N_1151);
nand U2296 (N_2296,N_1498,N_1020);
nand U2297 (N_2297,N_1194,N_1957);
nor U2298 (N_2298,N_1256,N_1075);
or U2299 (N_2299,N_1635,N_1897);
and U2300 (N_2300,N_1253,N_1124);
nor U2301 (N_2301,N_1705,N_1099);
and U2302 (N_2302,N_1639,N_1494);
nand U2303 (N_2303,N_1536,N_1540);
or U2304 (N_2304,N_1399,N_1250);
nand U2305 (N_2305,N_1331,N_1630);
and U2306 (N_2306,N_1486,N_1243);
and U2307 (N_2307,N_1018,N_1179);
or U2308 (N_2308,N_1178,N_1182);
or U2309 (N_2309,N_1640,N_1276);
nand U2310 (N_2310,N_1831,N_1110);
nand U2311 (N_2311,N_1586,N_1163);
nor U2312 (N_2312,N_1133,N_1882);
or U2313 (N_2313,N_1409,N_1458);
or U2314 (N_2314,N_1282,N_1636);
and U2315 (N_2315,N_1083,N_1959);
nand U2316 (N_2316,N_1117,N_1217);
nor U2317 (N_2317,N_1742,N_1366);
and U2318 (N_2318,N_1632,N_1377);
or U2319 (N_2319,N_1525,N_1448);
and U2320 (N_2320,N_1814,N_1208);
nand U2321 (N_2321,N_1349,N_1316);
xnor U2322 (N_2322,N_1524,N_1024);
nor U2323 (N_2323,N_1438,N_1193);
nand U2324 (N_2324,N_1031,N_1930);
nand U2325 (N_2325,N_1432,N_1006);
nand U2326 (N_2326,N_1824,N_1604);
and U2327 (N_2327,N_1726,N_1809);
nand U2328 (N_2328,N_1518,N_1337);
or U2329 (N_2329,N_1964,N_1482);
xor U2330 (N_2330,N_1140,N_1492);
or U2331 (N_2331,N_1803,N_1199);
or U2332 (N_2332,N_1900,N_1299);
and U2333 (N_2333,N_1869,N_1462);
nor U2334 (N_2334,N_1267,N_1461);
and U2335 (N_2335,N_1804,N_1596);
and U2336 (N_2336,N_1341,N_1917);
nand U2337 (N_2337,N_1707,N_1773);
xnor U2338 (N_2338,N_1469,N_1702);
or U2339 (N_2339,N_1527,N_1861);
nand U2340 (N_2340,N_1376,N_1721);
or U2341 (N_2341,N_1162,N_1565);
nor U2342 (N_2342,N_1483,N_1291);
or U2343 (N_2343,N_1350,N_1066);
nor U2344 (N_2344,N_1550,N_1559);
or U2345 (N_2345,N_1739,N_1507);
or U2346 (N_2346,N_1890,N_1986);
xnor U2347 (N_2347,N_1283,N_1338);
and U2348 (N_2348,N_1757,N_1103);
or U2349 (N_2349,N_1155,N_1173);
nand U2350 (N_2350,N_1206,N_1624);
nand U2351 (N_2351,N_1149,N_1706);
nand U2352 (N_2352,N_1043,N_1543);
nand U2353 (N_2353,N_1613,N_1397);
nor U2354 (N_2354,N_1516,N_1456);
nor U2355 (N_2355,N_1766,N_1740);
nor U2356 (N_2356,N_1752,N_1497);
and U2357 (N_2357,N_1296,N_1156);
and U2358 (N_2358,N_1735,N_1113);
nand U2359 (N_2359,N_1237,N_1641);
or U2360 (N_2360,N_1765,N_1732);
xor U2361 (N_2361,N_1404,N_1375);
and U2362 (N_2362,N_1411,N_1288);
or U2363 (N_2363,N_1355,N_1087);
or U2364 (N_2364,N_1017,N_1962);
nor U2365 (N_2365,N_1961,N_1380);
and U2366 (N_2366,N_1754,N_1175);
and U2367 (N_2367,N_1916,N_1437);
or U2368 (N_2368,N_1792,N_1146);
nand U2369 (N_2369,N_1301,N_1424);
nor U2370 (N_2370,N_1138,N_1147);
or U2371 (N_2371,N_1796,N_1383);
and U2372 (N_2372,N_1874,N_1819);
or U2373 (N_2373,N_1583,N_1104);
and U2374 (N_2374,N_1908,N_1327);
or U2375 (N_2375,N_1980,N_1914);
nor U2376 (N_2376,N_1617,N_1863);
nand U2377 (N_2377,N_1273,N_1285);
nand U2378 (N_2378,N_1044,N_1493);
nor U2379 (N_2379,N_1825,N_1813);
nand U2380 (N_2380,N_1141,N_1069);
or U2381 (N_2381,N_1496,N_1218);
and U2382 (N_2382,N_1590,N_1701);
nand U2383 (N_2383,N_1889,N_1667);
or U2384 (N_2384,N_1881,N_1145);
or U2385 (N_2385,N_1690,N_1275);
or U2386 (N_2386,N_1344,N_1616);
and U2387 (N_2387,N_1554,N_1729);
nand U2388 (N_2388,N_1320,N_1531);
nor U2389 (N_2389,N_1269,N_1946);
or U2390 (N_2390,N_1951,N_1053);
or U2391 (N_2391,N_1569,N_1127);
nand U2392 (N_2392,N_1730,N_1763);
nand U2393 (N_2393,N_1303,N_1336);
nand U2394 (N_2394,N_1129,N_1772);
or U2395 (N_2395,N_1011,N_1842);
nand U2396 (N_2396,N_1767,N_1441);
xnor U2397 (N_2397,N_1394,N_1840);
or U2398 (N_2398,N_1408,N_1203);
or U2399 (N_2399,N_1651,N_1774);
or U2400 (N_2400,N_1542,N_1828);
and U2401 (N_2401,N_1345,N_1713);
and U2402 (N_2402,N_1955,N_1189);
or U2403 (N_2403,N_1812,N_1071);
and U2404 (N_2404,N_1364,N_1563);
and U2405 (N_2405,N_1755,N_1340);
and U2406 (N_2406,N_1503,N_1886);
nand U2407 (N_2407,N_1947,N_1446);
or U2408 (N_2408,N_1352,N_1130);
nor U2409 (N_2409,N_1417,N_1718);
and U2410 (N_2410,N_1015,N_1317);
or U2411 (N_2411,N_1001,N_1985);
or U2412 (N_2412,N_1972,N_1152);
or U2413 (N_2413,N_1333,N_1776);
or U2414 (N_2414,N_1109,N_1570);
or U2415 (N_2415,N_1973,N_1334);
nand U2416 (N_2416,N_1615,N_1602);
or U2417 (N_2417,N_1758,N_1988);
and U2418 (N_2418,N_1321,N_1450);
or U2419 (N_2419,N_1600,N_1715);
nor U2420 (N_2420,N_1652,N_1877);
and U2421 (N_2421,N_1541,N_1696);
and U2422 (N_2422,N_1157,N_1262);
or U2423 (N_2423,N_1207,N_1725);
nand U2424 (N_2424,N_1013,N_1455);
or U2425 (N_2425,N_1235,N_1833);
nor U2426 (N_2426,N_1308,N_1257);
or U2427 (N_2427,N_1445,N_1846);
or U2428 (N_2428,N_1292,N_1219);
or U2429 (N_2429,N_1339,N_1694);
or U2430 (N_2430,N_1300,N_1935);
or U2431 (N_2431,N_1358,N_1523);
or U2432 (N_2432,N_1003,N_1815);
or U2433 (N_2433,N_1659,N_1898);
nor U2434 (N_2434,N_1782,N_1249);
or U2435 (N_2435,N_1511,N_1238);
or U2436 (N_2436,N_1032,N_1723);
nand U2437 (N_2437,N_1002,N_1870);
nand U2438 (N_2438,N_1400,N_1023);
nand U2439 (N_2439,N_1668,N_1745);
and U2440 (N_2440,N_1817,N_1638);
or U2441 (N_2441,N_1656,N_1034);
nor U2442 (N_2442,N_1753,N_1106);
or U2443 (N_2443,N_1114,N_1367);
nand U2444 (N_2444,N_1944,N_1673);
nor U2445 (N_2445,N_1628,N_1746);
or U2446 (N_2446,N_1307,N_1575);
or U2447 (N_2447,N_1677,N_1797);
nor U2448 (N_2448,N_1418,N_1784);
and U2449 (N_2449,N_1749,N_1646);
nand U2450 (N_2450,N_1471,N_1385);
and U2451 (N_2451,N_1911,N_1416);
nor U2452 (N_2452,N_1538,N_1070);
and U2453 (N_2453,N_1684,N_1852);
nand U2454 (N_2454,N_1343,N_1899);
and U2455 (N_2455,N_1556,N_1466);
nor U2456 (N_2456,N_1515,N_1868);
and U2457 (N_2457,N_1716,N_1328);
nand U2458 (N_2458,N_1619,N_1871);
nor U2459 (N_2459,N_1823,N_1045);
or U2460 (N_2460,N_1464,N_1052);
and U2461 (N_2461,N_1472,N_1674);
nor U2462 (N_2462,N_1160,N_1008);
xor U2463 (N_2463,N_1274,N_1111);
nor U2464 (N_2464,N_1522,N_1860);
nand U2465 (N_2465,N_1835,N_1722);
nand U2466 (N_2466,N_1500,N_1488);
nand U2467 (N_2467,N_1832,N_1698);
nand U2468 (N_2468,N_1187,N_1100);
or U2469 (N_2469,N_1391,N_1560);
and U2470 (N_2470,N_1885,N_1535);
nor U2471 (N_2471,N_1185,N_1545);
and U2472 (N_2472,N_1054,N_1016);
nor U2473 (N_2473,N_1661,N_1847);
and U2474 (N_2474,N_1866,N_1977);
nand U2475 (N_2475,N_1036,N_1323);
nand U2476 (N_2476,N_1078,N_1534);
nor U2477 (N_2477,N_1128,N_1115);
xor U2478 (N_2478,N_1372,N_1161);
or U2479 (N_2479,N_1495,N_1884);
or U2480 (N_2480,N_1795,N_1592);
nand U2481 (N_2481,N_1226,N_1572);
nor U2482 (N_2482,N_1457,N_1101);
nand U2483 (N_2483,N_1637,N_1412);
nor U2484 (N_2484,N_1949,N_1807);
nor U2485 (N_2485,N_1306,N_1891);
or U2486 (N_2486,N_1672,N_1856);
nand U2487 (N_2487,N_1314,N_1529);
or U2488 (N_2488,N_1744,N_1436);
and U2489 (N_2489,N_1850,N_1709);
nor U2490 (N_2490,N_1724,N_1154);
or U2491 (N_2491,N_1633,N_1664);
nor U2492 (N_2492,N_1539,N_1159);
or U2493 (N_2493,N_1984,N_1325);
nand U2494 (N_2494,N_1158,N_1330);
nand U2495 (N_2495,N_1290,N_1829);
or U2496 (N_2496,N_1544,N_1281);
or U2497 (N_2497,N_1144,N_1680);
or U2498 (N_2498,N_1286,N_1434);
and U2499 (N_2499,N_1594,N_1309);
nor U2500 (N_2500,N_1960,N_1153);
nand U2501 (N_2501,N_1212,N_1596);
and U2502 (N_2502,N_1490,N_1432);
nor U2503 (N_2503,N_1805,N_1957);
and U2504 (N_2504,N_1440,N_1302);
and U2505 (N_2505,N_1539,N_1233);
nor U2506 (N_2506,N_1718,N_1723);
and U2507 (N_2507,N_1032,N_1664);
and U2508 (N_2508,N_1368,N_1652);
nand U2509 (N_2509,N_1349,N_1829);
or U2510 (N_2510,N_1131,N_1304);
and U2511 (N_2511,N_1681,N_1361);
or U2512 (N_2512,N_1918,N_1217);
nor U2513 (N_2513,N_1727,N_1514);
and U2514 (N_2514,N_1200,N_1813);
and U2515 (N_2515,N_1516,N_1216);
and U2516 (N_2516,N_1685,N_1188);
nor U2517 (N_2517,N_1625,N_1362);
or U2518 (N_2518,N_1975,N_1760);
nand U2519 (N_2519,N_1449,N_1237);
xor U2520 (N_2520,N_1157,N_1369);
nor U2521 (N_2521,N_1340,N_1039);
nand U2522 (N_2522,N_1446,N_1825);
nand U2523 (N_2523,N_1923,N_1279);
or U2524 (N_2524,N_1285,N_1503);
and U2525 (N_2525,N_1670,N_1312);
and U2526 (N_2526,N_1499,N_1135);
nand U2527 (N_2527,N_1410,N_1238);
and U2528 (N_2528,N_1613,N_1441);
or U2529 (N_2529,N_1377,N_1402);
and U2530 (N_2530,N_1814,N_1344);
or U2531 (N_2531,N_1303,N_1736);
nand U2532 (N_2532,N_1236,N_1135);
nand U2533 (N_2533,N_1276,N_1610);
nand U2534 (N_2534,N_1985,N_1880);
or U2535 (N_2535,N_1728,N_1872);
nand U2536 (N_2536,N_1121,N_1106);
nand U2537 (N_2537,N_1872,N_1957);
nand U2538 (N_2538,N_1834,N_1242);
nor U2539 (N_2539,N_1894,N_1576);
nand U2540 (N_2540,N_1366,N_1825);
or U2541 (N_2541,N_1060,N_1546);
and U2542 (N_2542,N_1944,N_1704);
nand U2543 (N_2543,N_1757,N_1630);
nor U2544 (N_2544,N_1085,N_1809);
nor U2545 (N_2545,N_1749,N_1592);
nor U2546 (N_2546,N_1861,N_1160);
and U2547 (N_2547,N_1910,N_1570);
nand U2548 (N_2548,N_1742,N_1573);
and U2549 (N_2549,N_1401,N_1155);
and U2550 (N_2550,N_1580,N_1556);
or U2551 (N_2551,N_1897,N_1972);
nor U2552 (N_2552,N_1515,N_1432);
nor U2553 (N_2553,N_1241,N_1067);
nor U2554 (N_2554,N_1002,N_1302);
nand U2555 (N_2555,N_1117,N_1335);
xnor U2556 (N_2556,N_1955,N_1404);
and U2557 (N_2557,N_1242,N_1279);
nand U2558 (N_2558,N_1101,N_1973);
nand U2559 (N_2559,N_1932,N_1868);
or U2560 (N_2560,N_1645,N_1112);
and U2561 (N_2561,N_1750,N_1981);
and U2562 (N_2562,N_1125,N_1736);
nand U2563 (N_2563,N_1123,N_1593);
nor U2564 (N_2564,N_1897,N_1167);
nand U2565 (N_2565,N_1751,N_1304);
or U2566 (N_2566,N_1964,N_1051);
and U2567 (N_2567,N_1002,N_1389);
nor U2568 (N_2568,N_1350,N_1112);
nor U2569 (N_2569,N_1140,N_1144);
nor U2570 (N_2570,N_1359,N_1113);
nand U2571 (N_2571,N_1274,N_1871);
or U2572 (N_2572,N_1531,N_1466);
nand U2573 (N_2573,N_1441,N_1300);
nor U2574 (N_2574,N_1333,N_1839);
or U2575 (N_2575,N_1676,N_1821);
and U2576 (N_2576,N_1428,N_1473);
nor U2577 (N_2577,N_1674,N_1250);
or U2578 (N_2578,N_1583,N_1620);
or U2579 (N_2579,N_1336,N_1591);
and U2580 (N_2580,N_1053,N_1526);
nor U2581 (N_2581,N_1541,N_1405);
nand U2582 (N_2582,N_1490,N_1163);
nand U2583 (N_2583,N_1681,N_1421);
nor U2584 (N_2584,N_1307,N_1537);
nor U2585 (N_2585,N_1105,N_1663);
nand U2586 (N_2586,N_1057,N_1245);
nand U2587 (N_2587,N_1704,N_1375);
and U2588 (N_2588,N_1417,N_1071);
and U2589 (N_2589,N_1655,N_1336);
nor U2590 (N_2590,N_1595,N_1986);
and U2591 (N_2591,N_1213,N_1794);
xor U2592 (N_2592,N_1514,N_1939);
or U2593 (N_2593,N_1982,N_1882);
nand U2594 (N_2594,N_1115,N_1858);
xnor U2595 (N_2595,N_1251,N_1291);
nand U2596 (N_2596,N_1495,N_1398);
or U2597 (N_2597,N_1249,N_1964);
and U2598 (N_2598,N_1447,N_1359);
or U2599 (N_2599,N_1613,N_1658);
nand U2600 (N_2600,N_1071,N_1343);
nor U2601 (N_2601,N_1350,N_1273);
and U2602 (N_2602,N_1158,N_1298);
or U2603 (N_2603,N_1815,N_1711);
or U2604 (N_2604,N_1290,N_1166);
or U2605 (N_2605,N_1051,N_1694);
nor U2606 (N_2606,N_1603,N_1190);
or U2607 (N_2607,N_1060,N_1371);
nand U2608 (N_2608,N_1360,N_1959);
or U2609 (N_2609,N_1073,N_1151);
nand U2610 (N_2610,N_1728,N_1402);
nor U2611 (N_2611,N_1156,N_1347);
nand U2612 (N_2612,N_1217,N_1790);
nand U2613 (N_2613,N_1776,N_1355);
or U2614 (N_2614,N_1919,N_1946);
or U2615 (N_2615,N_1186,N_1163);
or U2616 (N_2616,N_1464,N_1134);
and U2617 (N_2617,N_1571,N_1296);
or U2618 (N_2618,N_1429,N_1216);
or U2619 (N_2619,N_1513,N_1679);
nor U2620 (N_2620,N_1760,N_1544);
or U2621 (N_2621,N_1696,N_1415);
nor U2622 (N_2622,N_1910,N_1156);
and U2623 (N_2623,N_1680,N_1615);
nor U2624 (N_2624,N_1384,N_1798);
nor U2625 (N_2625,N_1492,N_1402);
nand U2626 (N_2626,N_1477,N_1341);
and U2627 (N_2627,N_1956,N_1269);
or U2628 (N_2628,N_1695,N_1295);
and U2629 (N_2629,N_1286,N_1334);
and U2630 (N_2630,N_1680,N_1911);
or U2631 (N_2631,N_1721,N_1291);
nor U2632 (N_2632,N_1519,N_1261);
nand U2633 (N_2633,N_1889,N_1351);
nand U2634 (N_2634,N_1646,N_1296);
and U2635 (N_2635,N_1402,N_1893);
xnor U2636 (N_2636,N_1169,N_1072);
nor U2637 (N_2637,N_1894,N_1130);
xnor U2638 (N_2638,N_1038,N_1735);
or U2639 (N_2639,N_1047,N_1521);
nand U2640 (N_2640,N_1486,N_1728);
or U2641 (N_2641,N_1510,N_1281);
and U2642 (N_2642,N_1282,N_1224);
nand U2643 (N_2643,N_1930,N_1543);
and U2644 (N_2644,N_1102,N_1169);
and U2645 (N_2645,N_1789,N_1104);
and U2646 (N_2646,N_1845,N_1559);
and U2647 (N_2647,N_1501,N_1097);
or U2648 (N_2648,N_1297,N_1333);
or U2649 (N_2649,N_1750,N_1874);
nand U2650 (N_2650,N_1518,N_1043);
nand U2651 (N_2651,N_1015,N_1228);
nand U2652 (N_2652,N_1862,N_1352);
nor U2653 (N_2653,N_1542,N_1224);
xnor U2654 (N_2654,N_1258,N_1676);
and U2655 (N_2655,N_1029,N_1305);
nand U2656 (N_2656,N_1351,N_1581);
nand U2657 (N_2657,N_1085,N_1291);
nor U2658 (N_2658,N_1806,N_1889);
nor U2659 (N_2659,N_1602,N_1562);
nor U2660 (N_2660,N_1512,N_1606);
and U2661 (N_2661,N_1163,N_1937);
and U2662 (N_2662,N_1806,N_1679);
nor U2663 (N_2663,N_1650,N_1195);
nor U2664 (N_2664,N_1008,N_1184);
and U2665 (N_2665,N_1314,N_1427);
nor U2666 (N_2666,N_1776,N_1586);
nand U2667 (N_2667,N_1400,N_1931);
nor U2668 (N_2668,N_1183,N_1990);
nand U2669 (N_2669,N_1035,N_1888);
or U2670 (N_2670,N_1601,N_1275);
nand U2671 (N_2671,N_1561,N_1737);
and U2672 (N_2672,N_1960,N_1880);
or U2673 (N_2673,N_1004,N_1021);
nand U2674 (N_2674,N_1878,N_1363);
nand U2675 (N_2675,N_1566,N_1073);
nand U2676 (N_2676,N_1502,N_1610);
xor U2677 (N_2677,N_1828,N_1355);
or U2678 (N_2678,N_1191,N_1390);
or U2679 (N_2679,N_1417,N_1878);
nor U2680 (N_2680,N_1565,N_1539);
and U2681 (N_2681,N_1679,N_1844);
nor U2682 (N_2682,N_1205,N_1151);
nand U2683 (N_2683,N_1871,N_1306);
nand U2684 (N_2684,N_1466,N_1485);
and U2685 (N_2685,N_1177,N_1363);
nor U2686 (N_2686,N_1780,N_1822);
nor U2687 (N_2687,N_1540,N_1777);
and U2688 (N_2688,N_1446,N_1369);
or U2689 (N_2689,N_1032,N_1484);
and U2690 (N_2690,N_1380,N_1520);
xnor U2691 (N_2691,N_1943,N_1581);
nor U2692 (N_2692,N_1215,N_1925);
nor U2693 (N_2693,N_1250,N_1774);
nor U2694 (N_2694,N_1954,N_1305);
and U2695 (N_2695,N_1717,N_1984);
or U2696 (N_2696,N_1049,N_1611);
and U2697 (N_2697,N_1237,N_1373);
or U2698 (N_2698,N_1763,N_1000);
or U2699 (N_2699,N_1338,N_1942);
and U2700 (N_2700,N_1496,N_1828);
nor U2701 (N_2701,N_1094,N_1674);
nand U2702 (N_2702,N_1581,N_1853);
and U2703 (N_2703,N_1279,N_1712);
nand U2704 (N_2704,N_1319,N_1328);
nor U2705 (N_2705,N_1581,N_1254);
and U2706 (N_2706,N_1762,N_1813);
or U2707 (N_2707,N_1429,N_1120);
nand U2708 (N_2708,N_1327,N_1896);
and U2709 (N_2709,N_1504,N_1103);
nand U2710 (N_2710,N_1070,N_1335);
nor U2711 (N_2711,N_1211,N_1692);
or U2712 (N_2712,N_1453,N_1100);
or U2713 (N_2713,N_1868,N_1858);
and U2714 (N_2714,N_1133,N_1502);
nor U2715 (N_2715,N_1521,N_1066);
or U2716 (N_2716,N_1105,N_1399);
nand U2717 (N_2717,N_1000,N_1255);
and U2718 (N_2718,N_1119,N_1821);
nand U2719 (N_2719,N_1847,N_1932);
and U2720 (N_2720,N_1229,N_1980);
nand U2721 (N_2721,N_1040,N_1880);
or U2722 (N_2722,N_1701,N_1659);
and U2723 (N_2723,N_1855,N_1758);
xor U2724 (N_2724,N_1371,N_1641);
or U2725 (N_2725,N_1948,N_1613);
and U2726 (N_2726,N_1483,N_1371);
or U2727 (N_2727,N_1992,N_1132);
nand U2728 (N_2728,N_1570,N_1986);
nand U2729 (N_2729,N_1208,N_1842);
nor U2730 (N_2730,N_1303,N_1500);
nor U2731 (N_2731,N_1559,N_1576);
and U2732 (N_2732,N_1463,N_1445);
or U2733 (N_2733,N_1043,N_1002);
or U2734 (N_2734,N_1114,N_1150);
nor U2735 (N_2735,N_1380,N_1706);
or U2736 (N_2736,N_1360,N_1511);
nand U2737 (N_2737,N_1339,N_1456);
nand U2738 (N_2738,N_1410,N_1686);
and U2739 (N_2739,N_1443,N_1902);
or U2740 (N_2740,N_1415,N_1846);
and U2741 (N_2741,N_1796,N_1604);
and U2742 (N_2742,N_1087,N_1023);
nand U2743 (N_2743,N_1699,N_1184);
xnor U2744 (N_2744,N_1332,N_1267);
and U2745 (N_2745,N_1033,N_1279);
and U2746 (N_2746,N_1660,N_1427);
nor U2747 (N_2747,N_1670,N_1023);
nand U2748 (N_2748,N_1749,N_1147);
or U2749 (N_2749,N_1874,N_1695);
nor U2750 (N_2750,N_1459,N_1971);
and U2751 (N_2751,N_1292,N_1624);
nand U2752 (N_2752,N_1883,N_1960);
or U2753 (N_2753,N_1742,N_1278);
or U2754 (N_2754,N_1505,N_1164);
nor U2755 (N_2755,N_1994,N_1861);
and U2756 (N_2756,N_1845,N_1872);
and U2757 (N_2757,N_1373,N_1074);
and U2758 (N_2758,N_1016,N_1387);
nand U2759 (N_2759,N_1743,N_1680);
and U2760 (N_2760,N_1940,N_1461);
xor U2761 (N_2761,N_1575,N_1703);
and U2762 (N_2762,N_1953,N_1132);
nor U2763 (N_2763,N_1842,N_1439);
nand U2764 (N_2764,N_1732,N_1255);
or U2765 (N_2765,N_1073,N_1138);
nor U2766 (N_2766,N_1583,N_1473);
nor U2767 (N_2767,N_1679,N_1100);
nand U2768 (N_2768,N_1817,N_1011);
nor U2769 (N_2769,N_1798,N_1442);
or U2770 (N_2770,N_1805,N_1792);
nor U2771 (N_2771,N_1222,N_1907);
or U2772 (N_2772,N_1994,N_1409);
nand U2773 (N_2773,N_1629,N_1945);
and U2774 (N_2774,N_1483,N_1696);
nor U2775 (N_2775,N_1388,N_1198);
nand U2776 (N_2776,N_1342,N_1535);
and U2777 (N_2777,N_1927,N_1548);
and U2778 (N_2778,N_1127,N_1647);
nand U2779 (N_2779,N_1974,N_1538);
and U2780 (N_2780,N_1013,N_1368);
and U2781 (N_2781,N_1072,N_1165);
and U2782 (N_2782,N_1902,N_1754);
xnor U2783 (N_2783,N_1992,N_1493);
or U2784 (N_2784,N_1414,N_1022);
xor U2785 (N_2785,N_1054,N_1017);
and U2786 (N_2786,N_1687,N_1061);
nor U2787 (N_2787,N_1027,N_1178);
nand U2788 (N_2788,N_1953,N_1517);
or U2789 (N_2789,N_1720,N_1889);
nor U2790 (N_2790,N_1385,N_1515);
or U2791 (N_2791,N_1703,N_1255);
or U2792 (N_2792,N_1133,N_1383);
or U2793 (N_2793,N_1011,N_1841);
nor U2794 (N_2794,N_1415,N_1630);
nand U2795 (N_2795,N_1922,N_1812);
xnor U2796 (N_2796,N_1055,N_1430);
or U2797 (N_2797,N_1396,N_1336);
nand U2798 (N_2798,N_1364,N_1883);
and U2799 (N_2799,N_1320,N_1493);
xor U2800 (N_2800,N_1600,N_1066);
or U2801 (N_2801,N_1861,N_1139);
and U2802 (N_2802,N_1337,N_1470);
nor U2803 (N_2803,N_1290,N_1540);
nor U2804 (N_2804,N_1899,N_1924);
nand U2805 (N_2805,N_1434,N_1255);
and U2806 (N_2806,N_1228,N_1855);
and U2807 (N_2807,N_1148,N_1448);
nand U2808 (N_2808,N_1531,N_1445);
or U2809 (N_2809,N_1327,N_1215);
nand U2810 (N_2810,N_1283,N_1134);
nor U2811 (N_2811,N_1079,N_1364);
nor U2812 (N_2812,N_1736,N_1011);
nand U2813 (N_2813,N_1357,N_1475);
and U2814 (N_2814,N_1096,N_1600);
nand U2815 (N_2815,N_1079,N_1925);
xnor U2816 (N_2816,N_1347,N_1373);
or U2817 (N_2817,N_1149,N_1959);
and U2818 (N_2818,N_1132,N_1936);
nand U2819 (N_2819,N_1140,N_1775);
or U2820 (N_2820,N_1531,N_1547);
and U2821 (N_2821,N_1752,N_1251);
nand U2822 (N_2822,N_1578,N_1420);
and U2823 (N_2823,N_1141,N_1090);
nand U2824 (N_2824,N_1883,N_1584);
xor U2825 (N_2825,N_1268,N_1553);
or U2826 (N_2826,N_1812,N_1502);
and U2827 (N_2827,N_1743,N_1358);
nand U2828 (N_2828,N_1352,N_1052);
nand U2829 (N_2829,N_1489,N_1827);
nand U2830 (N_2830,N_1977,N_1785);
or U2831 (N_2831,N_1944,N_1607);
nand U2832 (N_2832,N_1828,N_1409);
or U2833 (N_2833,N_1655,N_1628);
and U2834 (N_2834,N_1358,N_1984);
or U2835 (N_2835,N_1047,N_1854);
nand U2836 (N_2836,N_1289,N_1012);
nand U2837 (N_2837,N_1939,N_1888);
nand U2838 (N_2838,N_1606,N_1110);
nand U2839 (N_2839,N_1602,N_1512);
nand U2840 (N_2840,N_1795,N_1677);
and U2841 (N_2841,N_1634,N_1853);
and U2842 (N_2842,N_1984,N_1554);
nand U2843 (N_2843,N_1363,N_1895);
nand U2844 (N_2844,N_1751,N_1095);
and U2845 (N_2845,N_1997,N_1050);
nand U2846 (N_2846,N_1010,N_1356);
xnor U2847 (N_2847,N_1928,N_1738);
or U2848 (N_2848,N_1715,N_1671);
nand U2849 (N_2849,N_1821,N_1906);
and U2850 (N_2850,N_1939,N_1748);
or U2851 (N_2851,N_1898,N_1731);
xor U2852 (N_2852,N_1102,N_1227);
nor U2853 (N_2853,N_1362,N_1802);
and U2854 (N_2854,N_1560,N_1220);
nor U2855 (N_2855,N_1848,N_1437);
nand U2856 (N_2856,N_1105,N_1941);
and U2857 (N_2857,N_1921,N_1748);
or U2858 (N_2858,N_1168,N_1820);
nand U2859 (N_2859,N_1447,N_1080);
nor U2860 (N_2860,N_1458,N_1001);
xor U2861 (N_2861,N_1507,N_1823);
xor U2862 (N_2862,N_1045,N_1768);
nand U2863 (N_2863,N_1272,N_1871);
and U2864 (N_2864,N_1553,N_1341);
or U2865 (N_2865,N_1067,N_1858);
nor U2866 (N_2866,N_1523,N_1884);
nor U2867 (N_2867,N_1194,N_1721);
nand U2868 (N_2868,N_1754,N_1825);
or U2869 (N_2869,N_1932,N_1458);
or U2870 (N_2870,N_1424,N_1767);
nor U2871 (N_2871,N_1184,N_1977);
or U2872 (N_2872,N_1761,N_1833);
nor U2873 (N_2873,N_1399,N_1526);
and U2874 (N_2874,N_1947,N_1514);
and U2875 (N_2875,N_1439,N_1150);
nand U2876 (N_2876,N_1470,N_1456);
and U2877 (N_2877,N_1346,N_1292);
or U2878 (N_2878,N_1419,N_1801);
and U2879 (N_2879,N_1983,N_1407);
nand U2880 (N_2880,N_1211,N_1265);
nand U2881 (N_2881,N_1298,N_1264);
or U2882 (N_2882,N_1939,N_1512);
nor U2883 (N_2883,N_1491,N_1214);
nand U2884 (N_2884,N_1794,N_1747);
and U2885 (N_2885,N_1483,N_1561);
and U2886 (N_2886,N_1043,N_1810);
nor U2887 (N_2887,N_1390,N_1130);
nor U2888 (N_2888,N_1835,N_1782);
and U2889 (N_2889,N_1348,N_1901);
and U2890 (N_2890,N_1949,N_1078);
nor U2891 (N_2891,N_1193,N_1709);
nor U2892 (N_2892,N_1085,N_1314);
or U2893 (N_2893,N_1940,N_1052);
nor U2894 (N_2894,N_1850,N_1420);
nor U2895 (N_2895,N_1730,N_1715);
xor U2896 (N_2896,N_1957,N_1526);
nor U2897 (N_2897,N_1051,N_1068);
and U2898 (N_2898,N_1924,N_1677);
nand U2899 (N_2899,N_1050,N_1978);
xor U2900 (N_2900,N_1946,N_1503);
nor U2901 (N_2901,N_1917,N_1933);
and U2902 (N_2902,N_1248,N_1236);
nand U2903 (N_2903,N_1216,N_1460);
and U2904 (N_2904,N_1518,N_1211);
or U2905 (N_2905,N_1397,N_1391);
nor U2906 (N_2906,N_1507,N_1558);
and U2907 (N_2907,N_1856,N_1834);
and U2908 (N_2908,N_1477,N_1442);
nand U2909 (N_2909,N_1262,N_1123);
nor U2910 (N_2910,N_1153,N_1387);
or U2911 (N_2911,N_1741,N_1345);
xor U2912 (N_2912,N_1163,N_1601);
nor U2913 (N_2913,N_1841,N_1999);
and U2914 (N_2914,N_1906,N_1413);
and U2915 (N_2915,N_1330,N_1730);
or U2916 (N_2916,N_1237,N_1487);
and U2917 (N_2917,N_1110,N_1997);
nand U2918 (N_2918,N_1049,N_1925);
nor U2919 (N_2919,N_1041,N_1283);
nand U2920 (N_2920,N_1121,N_1643);
and U2921 (N_2921,N_1884,N_1700);
or U2922 (N_2922,N_1381,N_1152);
or U2923 (N_2923,N_1156,N_1802);
nor U2924 (N_2924,N_1223,N_1032);
nand U2925 (N_2925,N_1887,N_1502);
nand U2926 (N_2926,N_1332,N_1284);
nor U2927 (N_2927,N_1469,N_1478);
or U2928 (N_2928,N_1425,N_1463);
and U2929 (N_2929,N_1725,N_1047);
or U2930 (N_2930,N_1330,N_1951);
or U2931 (N_2931,N_1069,N_1301);
and U2932 (N_2932,N_1474,N_1456);
nand U2933 (N_2933,N_1841,N_1169);
nand U2934 (N_2934,N_1034,N_1380);
nand U2935 (N_2935,N_1488,N_1783);
and U2936 (N_2936,N_1350,N_1093);
or U2937 (N_2937,N_1672,N_1064);
nor U2938 (N_2938,N_1768,N_1772);
xor U2939 (N_2939,N_1243,N_1271);
xnor U2940 (N_2940,N_1961,N_1220);
nand U2941 (N_2941,N_1384,N_1478);
nor U2942 (N_2942,N_1500,N_1471);
and U2943 (N_2943,N_1589,N_1100);
or U2944 (N_2944,N_1424,N_1036);
nor U2945 (N_2945,N_1752,N_1794);
nor U2946 (N_2946,N_1088,N_1574);
or U2947 (N_2947,N_1990,N_1977);
and U2948 (N_2948,N_1101,N_1293);
and U2949 (N_2949,N_1960,N_1519);
or U2950 (N_2950,N_1150,N_1778);
and U2951 (N_2951,N_1985,N_1744);
and U2952 (N_2952,N_1314,N_1886);
nand U2953 (N_2953,N_1849,N_1445);
or U2954 (N_2954,N_1686,N_1871);
nor U2955 (N_2955,N_1491,N_1106);
and U2956 (N_2956,N_1006,N_1732);
or U2957 (N_2957,N_1126,N_1146);
or U2958 (N_2958,N_1292,N_1691);
nor U2959 (N_2959,N_1975,N_1356);
nor U2960 (N_2960,N_1960,N_1509);
and U2961 (N_2961,N_1075,N_1750);
nor U2962 (N_2962,N_1150,N_1633);
nand U2963 (N_2963,N_1946,N_1959);
or U2964 (N_2964,N_1739,N_1229);
and U2965 (N_2965,N_1306,N_1222);
or U2966 (N_2966,N_1061,N_1847);
and U2967 (N_2967,N_1038,N_1324);
nand U2968 (N_2968,N_1195,N_1550);
and U2969 (N_2969,N_1131,N_1835);
and U2970 (N_2970,N_1896,N_1650);
nor U2971 (N_2971,N_1701,N_1147);
or U2972 (N_2972,N_1897,N_1749);
and U2973 (N_2973,N_1724,N_1803);
or U2974 (N_2974,N_1692,N_1025);
nand U2975 (N_2975,N_1322,N_1618);
and U2976 (N_2976,N_1486,N_1025);
and U2977 (N_2977,N_1260,N_1349);
and U2978 (N_2978,N_1206,N_1082);
and U2979 (N_2979,N_1373,N_1139);
nand U2980 (N_2980,N_1545,N_1473);
nand U2981 (N_2981,N_1761,N_1912);
or U2982 (N_2982,N_1816,N_1752);
and U2983 (N_2983,N_1881,N_1094);
nand U2984 (N_2984,N_1633,N_1453);
nor U2985 (N_2985,N_1218,N_1858);
and U2986 (N_2986,N_1382,N_1322);
and U2987 (N_2987,N_1842,N_1366);
and U2988 (N_2988,N_1001,N_1473);
and U2989 (N_2989,N_1078,N_1365);
or U2990 (N_2990,N_1086,N_1484);
nor U2991 (N_2991,N_1639,N_1625);
and U2992 (N_2992,N_1393,N_1101);
or U2993 (N_2993,N_1347,N_1684);
and U2994 (N_2994,N_1459,N_1390);
and U2995 (N_2995,N_1428,N_1009);
nor U2996 (N_2996,N_1546,N_1725);
or U2997 (N_2997,N_1102,N_1082);
nor U2998 (N_2998,N_1861,N_1099);
and U2999 (N_2999,N_1753,N_1316);
and UO_0 (O_0,N_2180,N_2062);
and UO_1 (O_1,N_2728,N_2580);
and UO_2 (O_2,N_2327,N_2585);
or UO_3 (O_3,N_2702,N_2146);
and UO_4 (O_4,N_2407,N_2615);
and UO_5 (O_5,N_2261,N_2174);
nand UO_6 (O_6,N_2726,N_2276);
and UO_7 (O_7,N_2961,N_2923);
xnor UO_8 (O_8,N_2742,N_2007);
and UO_9 (O_9,N_2222,N_2707);
nor UO_10 (O_10,N_2342,N_2293);
and UO_11 (O_11,N_2470,N_2207);
nor UO_12 (O_12,N_2794,N_2595);
or UO_13 (O_13,N_2769,N_2401);
nand UO_14 (O_14,N_2166,N_2210);
nand UO_15 (O_15,N_2715,N_2879);
or UO_16 (O_16,N_2331,N_2359);
nand UO_17 (O_17,N_2388,N_2937);
nor UO_18 (O_18,N_2861,N_2897);
nor UO_19 (O_19,N_2561,N_2283);
nor UO_20 (O_20,N_2194,N_2380);
and UO_21 (O_21,N_2040,N_2993);
or UO_22 (O_22,N_2853,N_2608);
nand UO_23 (O_23,N_2109,N_2969);
nor UO_24 (O_24,N_2963,N_2968);
or UO_25 (O_25,N_2026,N_2527);
or UO_26 (O_26,N_2893,N_2133);
or UO_27 (O_27,N_2373,N_2243);
xnor UO_28 (O_28,N_2234,N_2217);
and UO_29 (O_29,N_2178,N_2238);
xnor UO_30 (O_30,N_2858,N_2902);
xnor UO_31 (O_31,N_2617,N_2673);
and UO_32 (O_32,N_2928,N_2984);
or UO_33 (O_33,N_2930,N_2036);
or UO_34 (O_34,N_2569,N_2556);
or UO_35 (O_35,N_2254,N_2816);
nand UO_36 (O_36,N_2834,N_2920);
or UO_37 (O_37,N_2572,N_2932);
or UO_38 (O_38,N_2732,N_2131);
or UO_39 (O_39,N_2777,N_2185);
and UO_40 (O_40,N_2637,N_2924);
or UO_41 (O_41,N_2112,N_2960);
and UO_42 (O_42,N_2059,N_2658);
or UO_43 (O_43,N_2134,N_2160);
nor UO_44 (O_44,N_2354,N_2631);
nand UO_45 (O_45,N_2206,N_2111);
nand UO_46 (O_46,N_2657,N_2034);
and UO_47 (O_47,N_2712,N_2095);
xor UO_48 (O_48,N_2457,N_2268);
or UO_49 (O_49,N_2762,N_2357);
nand UO_50 (O_50,N_2278,N_2303);
and UO_51 (O_51,N_2886,N_2014);
nor UO_52 (O_52,N_2730,N_2396);
nand UO_53 (O_53,N_2603,N_2433);
xnor UO_54 (O_54,N_2668,N_2597);
nand UO_55 (O_55,N_2768,N_2314);
nand UO_56 (O_56,N_2934,N_2539);
or UO_57 (O_57,N_2577,N_2517);
nor UO_58 (O_58,N_2905,N_2884);
xor UO_59 (O_59,N_2151,N_2395);
and UO_60 (O_60,N_2624,N_2976);
nor UO_61 (O_61,N_2154,N_2537);
and UO_62 (O_62,N_2697,N_2213);
and UO_63 (O_63,N_2800,N_2127);
and UO_64 (O_64,N_2257,N_2423);
nand UO_65 (O_65,N_2925,N_2320);
xor UO_66 (O_66,N_2656,N_2288);
xor UO_67 (O_67,N_2262,N_2531);
or UO_68 (O_68,N_2755,N_2672);
nand UO_69 (O_69,N_2018,N_2512);
and UO_70 (O_70,N_2247,N_2964);
nand UO_71 (O_71,N_2746,N_2277);
or UO_72 (O_72,N_2236,N_2554);
nor UO_73 (O_73,N_2521,N_2267);
nand UO_74 (O_74,N_2980,N_2460);
and UO_75 (O_75,N_2877,N_2705);
or UO_76 (O_76,N_2872,N_2651);
nor UO_77 (O_77,N_2411,N_2559);
nor UO_78 (O_78,N_2786,N_2016);
and UO_79 (O_79,N_2970,N_2368);
nand UO_80 (O_80,N_2788,N_2035);
or UO_81 (O_81,N_2046,N_2057);
nand UO_82 (O_82,N_2335,N_2749);
nor UO_83 (O_83,N_2900,N_2962);
nand UO_84 (O_84,N_2604,N_2859);
and UO_85 (O_85,N_2004,N_2593);
and UO_86 (O_86,N_2723,N_2116);
or UO_87 (O_87,N_2148,N_2001);
and UO_88 (O_88,N_2379,N_2065);
and UO_89 (O_89,N_2563,N_2850);
and UO_90 (O_90,N_2449,N_2122);
or UO_91 (O_91,N_2224,N_2333);
and UO_92 (O_92,N_2179,N_2391);
nor UO_93 (O_93,N_2558,N_2113);
and UO_94 (O_94,N_2130,N_2764);
or UO_95 (O_95,N_2232,N_2921);
nand UO_96 (O_96,N_2947,N_2197);
and UO_97 (O_97,N_2215,N_2128);
or UO_98 (O_98,N_2802,N_2329);
and UO_99 (O_99,N_2757,N_2434);
or UO_100 (O_100,N_2727,N_2842);
or UO_101 (O_101,N_2248,N_2488);
nand UO_102 (O_102,N_2092,N_2515);
or UO_103 (O_103,N_2621,N_2361);
nor UO_104 (O_104,N_2100,N_2241);
or UO_105 (O_105,N_2177,N_2889);
nand UO_106 (O_106,N_2733,N_2760);
nor UO_107 (O_107,N_2069,N_2143);
and UO_108 (O_108,N_2711,N_2282);
nand UO_109 (O_109,N_2601,N_2381);
nor UO_110 (O_110,N_2880,N_2692);
or UO_111 (O_111,N_2070,N_2562);
nand UO_112 (O_112,N_2084,N_2203);
nor UO_113 (O_113,N_2774,N_2358);
nand UO_114 (O_114,N_2321,N_2010);
nand UO_115 (O_115,N_2867,N_2060);
and UO_116 (O_116,N_2334,N_2101);
nand UO_117 (O_117,N_2633,N_2641);
or UO_118 (O_118,N_2235,N_2856);
nand UO_119 (O_119,N_2804,N_2883);
nand UO_120 (O_120,N_2417,N_2300);
nor UO_121 (O_121,N_2938,N_2287);
and UO_122 (O_122,N_2549,N_2227);
nor UO_123 (O_123,N_2184,N_2564);
nor UO_124 (O_124,N_2781,N_2021);
or UO_125 (O_125,N_2892,N_2497);
and UO_126 (O_126,N_2832,N_2731);
nand UO_127 (O_127,N_2478,N_2110);
and UO_128 (O_128,N_2139,N_2901);
and UO_129 (O_129,N_2170,N_2586);
and UO_130 (O_130,N_2190,N_2191);
nand UO_131 (O_131,N_2119,N_2587);
or UO_132 (O_132,N_2507,N_2522);
nor UO_133 (O_133,N_2458,N_2990);
nand UO_134 (O_134,N_2230,N_2447);
nand UO_135 (O_135,N_2582,N_2799);
and UO_136 (O_136,N_2441,N_2136);
nor UO_137 (O_137,N_2363,N_2374);
and UO_138 (O_138,N_2126,N_2446);
nand UO_139 (O_139,N_2801,N_2894);
nand UO_140 (O_140,N_2041,N_2500);
xnor UO_141 (O_141,N_2703,N_2514);
nand UO_142 (O_142,N_2286,N_2513);
or UO_143 (O_143,N_2677,N_2263);
or UO_144 (O_144,N_2958,N_2294);
and UO_145 (O_145,N_2348,N_2022);
nand UO_146 (O_146,N_2337,N_2750);
nand UO_147 (O_147,N_2653,N_2669);
or UO_148 (O_148,N_2590,N_2156);
nor UO_149 (O_149,N_2941,N_2690);
or UO_150 (O_150,N_2534,N_2142);
and UO_151 (O_151,N_2356,N_2695);
and UO_152 (O_152,N_2685,N_2664);
xor UO_153 (O_153,N_2080,N_2461);
or UO_154 (O_154,N_2017,N_2208);
nand UO_155 (O_155,N_2752,N_2415);
or UO_156 (O_156,N_2408,N_2161);
or UO_157 (O_157,N_2089,N_2281);
nand UO_158 (O_158,N_2273,N_2211);
or UO_159 (O_159,N_2050,N_2214);
nor UO_160 (O_160,N_2548,N_2717);
nor UO_161 (O_161,N_2349,N_2581);
and UO_162 (O_162,N_2484,N_2228);
nand UO_163 (O_163,N_2091,N_2220);
and UO_164 (O_164,N_2384,N_2491);
or UO_165 (O_165,N_2650,N_2706);
nor UO_166 (O_166,N_2583,N_2875);
nand UO_167 (O_167,N_2983,N_2551);
nand UO_168 (O_168,N_2822,N_2412);
nand UO_169 (O_169,N_2318,N_2519);
or UO_170 (O_170,N_2410,N_2860);
or UO_171 (O_171,N_2012,N_2173);
nor UO_172 (O_172,N_2125,N_2868);
nor UO_173 (O_173,N_2103,N_2094);
and UO_174 (O_174,N_2152,N_2871);
or UO_175 (O_175,N_2005,N_2988);
nor UO_176 (O_176,N_2957,N_2767);
and UO_177 (O_177,N_2836,N_2432);
nand UO_178 (O_178,N_2594,N_2175);
and UO_179 (O_179,N_2123,N_2024);
nor UO_180 (O_180,N_2474,N_2828);
or UO_181 (O_181,N_2431,N_2885);
nand UO_182 (O_182,N_2445,N_2301);
nand UO_183 (O_183,N_2629,N_2242);
and UO_184 (O_184,N_2896,N_2870);
nor UO_185 (O_185,N_2782,N_2812);
or UO_186 (O_186,N_2188,N_2847);
nand UO_187 (O_187,N_2444,N_2660);
nor UO_188 (O_188,N_2791,N_2555);
and UO_189 (O_189,N_2663,N_2085);
nor UO_190 (O_190,N_2508,N_2948);
and UO_191 (O_191,N_2443,N_2317);
nor UO_192 (O_192,N_2503,N_2316);
or UO_193 (O_193,N_2223,N_2043);
and UO_194 (O_194,N_2270,N_2102);
or UO_195 (O_195,N_2694,N_2025);
and UO_196 (O_196,N_2611,N_2647);
and UO_197 (O_197,N_2347,N_2124);
nand UO_198 (O_198,N_2783,N_2451);
or UO_199 (O_199,N_2745,N_2216);
nor UO_200 (O_200,N_2231,N_2031);
nand UO_201 (O_201,N_2324,N_2813);
or UO_202 (O_202,N_2201,N_2319);
nor UO_203 (O_203,N_2688,N_2106);
nand UO_204 (O_204,N_2913,N_2833);
or UO_205 (O_205,N_2452,N_2876);
and UO_206 (O_206,N_2542,N_2632);
or UO_207 (O_207,N_2141,N_2667);
nand UO_208 (O_208,N_2399,N_2602);
nand UO_209 (O_209,N_2851,N_2149);
and UO_210 (O_210,N_2066,N_2419);
xnor UO_211 (O_211,N_2121,N_2675);
nand UO_212 (O_212,N_2229,N_2638);
nor UO_213 (O_213,N_2909,N_2392);
nand UO_214 (O_214,N_2761,N_2009);
or UO_215 (O_215,N_2560,N_2074);
nor UO_216 (O_216,N_2353,N_2931);
or UO_217 (O_217,N_2259,N_2492);
nor UO_218 (O_218,N_2129,N_2264);
and UO_219 (O_219,N_2935,N_2489);
nand UO_220 (O_220,N_2082,N_2994);
nor UO_221 (O_221,N_2827,N_2140);
nor UO_222 (O_222,N_2290,N_2953);
or UO_223 (O_223,N_2713,N_2568);
nor UO_224 (O_224,N_2670,N_2328);
or UO_225 (O_225,N_2225,N_2255);
and UO_226 (O_226,N_2516,N_2734);
or UO_227 (O_227,N_2323,N_2051);
nor UO_228 (O_228,N_2943,N_2809);
nand UO_229 (O_229,N_2545,N_2468);
nor UO_230 (O_230,N_2814,N_2400);
nor UO_231 (O_231,N_2792,N_2308);
nand UO_232 (O_232,N_2536,N_2735);
nor UO_233 (O_233,N_2219,N_2553);
or UO_234 (O_234,N_2546,N_2708);
nor UO_235 (O_235,N_2086,N_2779);
and UO_236 (O_236,N_2754,N_2473);
nand UO_237 (O_237,N_2952,N_2493);
nor UO_238 (O_238,N_2540,N_2426);
or UO_239 (O_239,N_2233,N_2793);
or UO_240 (O_240,N_2274,N_2543);
nand UO_241 (O_241,N_2118,N_2033);
and UO_242 (O_242,N_2465,N_2117);
and UO_243 (O_243,N_2682,N_2003);
and UO_244 (O_244,N_2098,N_2592);
or UO_245 (O_245,N_2304,N_2145);
and UO_246 (O_246,N_2296,N_2251);
or UO_247 (O_247,N_2578,N_2881);
xor UO_248 (O_248,N_2710,N_2053);
and UO_249 (O_249,N_2700,N_2153);
or UO_250 (O_250,N_2620,N_2023);
nand UO_251 (O_251,N_2825,N_2639);
nand UO_252 (O_252,N_2138,N_2365);
nand UO_253 (O_253,N_2424,N_2835);
nor UO_254 (O_254,N_2904,N_2908);
and UO_255 (O_255,N_2192,N_2372);
and UO_256 (O_256,N_2698,N_2490);
nand UO_257 (O_257,N_2068,N_2654);
and UO_258 (O_258,N_2075,N_2907);
or UO_259 (O_259,N_2428,N_2830);
or UO_260 (O_260,N_2405,N_2097);
xnor UO_261 (O_261,N_2550,N_2823);
or UO_262 (O_262,N_2917,N_2798);
nand UO_263 (O_263,N_2459,N_2666);
or UO_264 (O_264,N_2951,N_2176);
nand UO_265 (O_265,N_2376,N_2378);
nor UO_266 (O_266,N_2829,N_2849);
nor UO_267 (O_267,N_2996,N_2662);
nand UO_268 (O_268,N_2571,N_2453);
and UO_269 (O_269,N_2093,N_2495);
nor UO_270 (O_270,N_2533,N_2916);
nand UO_271 (O_271,N_2045,N_2502);
nor UO_272 (O_272,N_2476,N_2079);
nor UO_273 (O_273,N_2370,N_2071);
nand UO_274 (O_274,N_2366,N_2462);
nand UO_275 (O_275,N_2427,N_2520);
nand UO_276 (O_276,N_2607,N_2506);
or UO_277 (O_277,N_2403,N_2077);
or UO_278 (O_278,N_2684,N_2808);
nor UO_279 (O_279,N_2387,N_2311);
nand UO_280 (O_280,N_2310,N_2971);
nor UO_281 (O_281,N_2183,N_2250);
nand UO_282 (O_282,N_2162,N_2819);
nor UO_283 (O_283,N_2584,N_2115);
or UO_284 (O_284,N_2529,N_2518);
or UO_285 (O_285,N_2630,N_2440);
and UO_286 (O_286,N_2269,N_2863);
and UO_287 (O_287,N_2891,N_2073);
and UO_288 (O_288,N_2272,N_2439);
nor UO_289 (O_289,N_2628,N_2182);
and UO_290 (O_290,N_2627,N_2414);
nand UO_291 (O_291,N_2911,N_2186);
nor UO_292 (O_292,N_2992,N_2108);
and UO_293 (O_293,N_2168,N_2467);
nor UO_294 (O_294,N_2743,N_2642);
nor UO_295 (O_295,N_2795,N_2736);
and UO_296 (O_296,N_2253,N_2846);
or UO_297 (O_297,N_2946,N_2704);
nor UO_298 (O_298,N_2914,N_2279);
nand UO_299 (O_299,N_2463,N_2390);
nand UO_300 (O_300,N_2817,N_2895);
or UO_301 (O_301,N_2298,N_2854);
nor UO_302 (O_302,N_2693,N_2939);
and UO_303 (O_303,N_2790,N_2864);
and UO_304 (O_304,N_2857,N_2008);
and UO_305 (O_305,N_2701,N_2716);
xnor UO_306 (O_306,N_2865,N_2504);
nor UO_307 (O_307,N_2332,N_2780);
xor UO_308 (O_308,N_2579,N_2634);
and UO_309 (O_309,N_2137,N_2076);
nand UO_310 (O_310,N_2686,N_2785);
nand UO_311 (O_311,N_2944,N_2613);
and UO_312 (O_312,N_2718,N_2049);
nand UO_313 (O_313,N_2888,N_2386);
nand UO_314 (O_314,N_2918,N_2397);
and UO_315 (O_315,N_2343,N_2936);
nor UO_316 (O_316,N_2266,N_2505);
or UO_317 (O_317,N_2037,N_2165);
or UO_318 (O_318,N_2226,N_2691);
and UO_319 (O_319,N_2164,N_2887);
or UO_320 (O_320,N_2326,N_2967);
or UO_321 (O_321,N_2030,N_2525);
or UO_322 (O_322,N_2566,N_2574);
and UO_323 (O_323,N_2966,N_2978);
and UO_324 (O_324,N_2172,N_2501);
or UO_325 (O_325,N_2299,N_2199);
or UO_326 (O_326,N_2605,N_2425);
nor UO_327 (O_327,N_2739,N_2523);
nand UO_328 (O_328,N_2193,N_2949);
nand UO_329 (O_329,N_2028,N_2511);
and UO_330 (O_330,N_2312,N_2635);
nand UO_331 (O_331,N_2275,N_2200);
nor UO_332 (O_332,N_2787,N_2322);
or UO_333 (O_333,N_2776,N_2998);
or UO_334 (O_334,N_2061,N_2150);
and UO_335 (O_335,N_2246,N_2481);
nor UO_336 (O_336,N_2747,N_2438);
nand UO_337 (O_337,N_2950,N_2763);
or UO_338 (O_338,N_2596,N_2430);
nor UO_339 (O_339,N_2524,N_2910);
and UO_340 (O_340,N_2355,N_2088);
nor UO_341 (O_341,N_2011,N_2625);
nand UO_342 (O_342,N_2442,N_2655);
nand UO_343 (O_343,N_2709,N_2078);
or UO_344 (O_344,N_2002,N_2820);
or UO_345 (O_345,N_2413,N_2135);
nor UO_346 (O_346,N_2047,N_2064);
or UO_347 (O_347,N_2464,N_2855);
nand UO_348 (O_348,N_2067,N_2873);
nor UO_349 (O_349,N_2575,N_2671);
or UO_350 (O_350,N_2158,N_2995);
nor UO_351 (O_351,N_2959,N_2541);
nor UO_352 (O_352,N_2090,N_2284);
xor UO_353 (O_353,N_2371,N_2552);
nor UO_354 (O_354,N_2680,N_2659);
and UO_355 (O_355,N_2927,N_2307);
nor UO_356 (O_356,N_2382,N_2991);
or UO_357 (O_357,N_2325,N_2719);
and UO_358 (O_358,N_2058,N_2683);
nor UO_359 (O_359,N_2926,N_2997);
or UO_360 (O_360,N_2422,N_2052);
or UO_361 (O_361,N_2510,N_2899);
and UO_362 (O_362,N_2824,N_2038);
or UO_363 (O_363,N_2072,N_2099);
and UO_364 (O_364,N_2526,N_2985);
or UO_365 (O_365,N_2838,N_2687);
nand UO_366 (O_366,N_2292,N_2942);
nor UO_367 (O_367,N_2039,N_2313);
nand UO_368 (O_368,N_2280,N_2202);
nor UO_369 (O_369,N_2144,N_2239);
and UO_370 (O_370,N_2919,N_2204);
nand UO_371 (O_371,N_2954,N_2929);
nand UO_372 (O_372,N_2773,N_2260);
and UO_373 (O_373,N_2163,N_2104);
nor UO_374 (O_374,N_2351,N_2013);
or UO_375 (O_375,N_2006,N_2418);
nor UO_376 (O_376,N_2171,N_2285);
and UO_377 (O_377,N_2606,N_2610);
nand UO_378 (O_378,N_2645,N_2665);
nand UO_379 (O_379,N_2479,N_2643);
nand UO_380 (O_380,N_2766,N_2544);
and UO_381 (O_381,N_2435,N_2496);
nand UO_382 (O_382,N_2973,N_2999);
nor UO_383 (O_383,N_2981,N_2455);
or UO_384 (O_384,N_2498,N_2797);
nor UO_385 (O_385,N_2898,N_2915);
or UO_386 (O_386,N_2982,N_2448);
nor UO_387 (O_387,N_2565,N_2852);
nand UO_388 (O_388,N_2528,N_2724);
or UO_389 (O_389,N_2362,N_2375);
or UO_390 (O_390,N_2345,N_2421);
nor UO_391 (O_391,N_2722,N_2751);
and UO_392 (O_392,N_2874,N_2912);
and UO_393 (O_393,N_2315,N_2977);
nor UO_394 (O_394,N_2729,N_2840);
nand UO_395 (O_395,N_2297,N_2205);
xnor UO_396 (O_396,N_2483,N_2289);
and UO_397 (O_397,N_2765,N_2056);
nor UO_398 (O_398,N_2081,N_2212);
and UO_399 (O_399,N_2167,N_2107);
nand UO_400 (O_400,N_2922,N_2020);
and UO_401 (O_401,N_2029,N_2841);
and UO_402 (O_402,N_2803,N_2940);
and UO_403 (O_403,N_2393,N_2509);
or UO_404 (O_404,N_2955,N_2420);
or UO_405 (O_405,N_2588,N_2622);
nor UO_406 (O_406,N_2302,N_2600);
and UO_407 (O_407,N_2377,N_2385);
or UO_408 (O_408,N_2573,N_2811);
nand UO_409 (O_409,N_2599,N_2450);
or UO_410 (O_410,N_2394,N_2759);
or UO_411 (O_411,N_2155,N_2339);
or UO_412 (O_412,N_2725,N_2721);
nand UO_413 (O_413,N_2591,N_2689);
nor UO_414 (O_414,N_2352,N_2758);
nand UO_415 (O_415,N_2844,N_2741);
and UO_416 (O_416,N_2187,N_2240);
or UO_417 (O_417,N_2532,N_2044);
nand UO_418 (O_418,N_2619,N_2796);
or UO_419 (O_419,N_2748,N_2878);
and UO_420 (O_420,N_2866,N_2032);
or UO_421 (O_421,N_2696,N_2652);
or UO_422 (O_422,N_2198,N_2636);
and UO_423 (O_423,N_2195,N_2330);
nand UO_424 (O_424,N_2114,N_2810);
nor UO_425 (O_425,N_2530,N_2576);
nor UO_426 (O_426,N_2291,N_2063);
nor UO_427 (O_427,N_2048,N_2956);
nor UO_428 (O_428,N_2972,N_2055);
nand UO_429 (O_429,N_2640,N_2404);
nand UO_430 (O_430,N_2979,N_2494);
or UO_431 (O_431,N_2341,N_2305);
or UO_432 (O_432,N_2648,N_2346);
and UO_433 (O_433,N_2535,N_2890);
or UO_434 (O_434,N_2309,N_2839);
and UO_435 (O_435,N_2649,N_2256);
nand UO_436 (O_436,N_2557,N_2364);
nor UO_437 (O_437,N_2775,N_2054);
xor UO_438 (O_438,N_2678,N_2389);
or UO_439 (O_439,N_2770,N_2805);
nor UO_440 (O_440,N_2598,N_2027);
nand UO_441 (O_441,N_2244,N_2626);
and UO_442 (O_442,N_2087,N_2499);
nand UO_443 (O_443,N_2661,N_2974);
xnor UO_444 (O_444,N_2105,N_2837);
nand UO_445 (O_445,N_2644,N_2265);
nand UO_446 (O_446,N_2986,N_2843);
and UO_447 (O_447,N_2681,N_2096);
xor UO_448 (O_448,N_2845,N_2429);
nand UO_449 (O_449,N_2945,N_2987);
nand UO_450 (O_450,N_2406,N_2567);
nand UO_451 (O_451,N_2570,N_2756);
or UO_452 (O_452,N_2409,N_2609);
and UO_453 (O_453,N_2471,N_2196);
nand UO_454 (O_454,N_2740,N_2295);
nor UO_455 (O_455,N_2245,N_2147);
or UO_456 (O_456,N_2437,N_2000);
nor UO_457 (O_457,N_2538,N_2862);
and UO_458 (O_458,N_2340,N_2042);
or UO_459 (O_459,N_2015,N_2271);
or UO_460 (O_460,N_2367,N_2169);
and UO_461 (O_461,N_2738,N_2882);
and UO_462 (O_462,N_2789,N_2646);
and UO_463 (O_463,N_2674,N_2469);
nor UO_464 (O_464,N_2120,N_2821);
and UO_465 (O_465,N_2258,N_2249);
and UO_466 (O_466,N_2676,N_2189);
and UO_467 (O_467,N_2589,N_2398);
or UO_468 (O_468,N_2618,N_2975);
and UO_469 (O_469,N_2485,N_2784);
nor UO_470 (O_470,N_2714,N_2157);
or UO_471 (O_471,N_2903,N_2132);
or UO_472 (O_472,N_2753,N_2252);
nand UO_473 (O_473,N_2456,N_2778);
or UO_474 (O_474,N_2477,N_2933);
or UO_475 (O_475,N_2612,N_2221);
and UO_476 (O_476,N_2771,N_2869);
and UO_477 (O_477,N_2744,N_2336);
nor UO_478 (O_478,N_2806,N_2209);
or UO_479 (O_479,N_2344,N_2487);
nor UO_480 (O_480,N_2815,N_2482);
or UO_481 (O_481,N_2338,N_2480);
nand UO_482 (O_482,N_2306,N_2218);
or UO_483 (O_483,N_2614,N_2402);
nor UO_484 (O_484,N_2699,N_2679);
and UO_485 (O_485,N_2350,N_2369);
nor UO_486 (O_486,N_2807,N_2616);
and UO_487 (O_487,N_2826,N_2475);
and UO_488 (O_488,N_2472,N_2772);
nor UO_489 (O_489,N_2454,N_2720);
nor UO_490 (O_490,N_2848,N_2416);
nor UO_491 (O_491,N_2486,N_2989);
xor UO_492 (O_492,N_2083,N_2466);
nand UO_493 (O_493,N_2623,N_2906);
xor UO_494 (O_494,N_2383,N_2965);
nor UO_495 (O_495,N_2737,N_2831);
and UO_496 (O_496,N_2436,N_2360);
nor UO_497 (O_497,N_2818,N_2159);
xor UO_498 (O_498,N_2237,N_2019);
or UO_499 (O_499,N_2547,N_2181);
endmodule