module basic_750_5000_1000_25_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_247,In_18);
and U1 (N_1,In_198,In_49);
and U2 (N_2,In_571,In_739);
or U3 (N_3,In_249,In_426);
nand U4 (N_4,In_472,In_686);
or U5 (N_5,In_581,In_604);
and U6 (N_6,In_172,In_524);
or U7 (N_7,In_150,In_241);
or U8 (N_8,In_27,In_430);
nand U9 (N_9,In_421,In_210);
nand U10 (N_10,In_293,In_175);
nor U11 (N_11,In_494,In_577);
or U12 (N_12,In_480,In_443);
and U13 (N_13,In_419,In_567);
nor U14 (N_14,In_559,In_227);
nor U15 (N_15,In_435,In_646);
or U16 (N_16,In_389,In_616);
and U17 (N_17,In_225,In_169);
and U18 (N_18,In_274,In_718);
and U19 (N_19,In_676,In_645);
and U20 (N_20,In_569,In_286);
xnor U21 (N_21,In_254,In_434);
nand U22 (N_22,In_135,In_436);
xor U23 (N_23,In_416,In_107);
nand U24 (N_24,In_272,In_670);
nor U25 (N_25,In_95,In_562);
nand U26 (N_26,In_558,In_582);
nor U27 (N_27,In_4,In_398);
nor U28 (N_28,In_86,In_271);
or U29 (N_29,In_112,In_690);
and U30 (N_30,In_590,In_209);
nor U31 (N_31,In_102,In_193);
and U32 (N_32,In_391,In_136);
or U33 (N_33,In_534,In_712);
nor U34 (N_34,In_194,In_155);
nand U35 (N_35,In_279,In_8);
or U36 (N_36,In_585,In_242);
and U37 (N_37,In_429,In_176);
and U38 (N_38,In_38,In_386);
nand U39 (N_39,In_456,In_723);
nor U40 (N_40,In_99,In_142);
nand U41 (N_41,In_285,In_108);
nand U42 (N_42,In_665,In_10);
and U43 (N_43,In_695,In_167);
nand U44 (N_44,In_470,In_588);
xor U45 (N_45,In_608,In_277);
xnor U46 (N_46,In_121,In_724);
or U47 (N_47,In_168,In_477);
or U48 (N_48,In_230,In_46);
nand U49 (N_49,In_333,In_687);
or U50 (N_50,In_399,In_371);
nor U51 (N_51,In_334,In_433);
nand U52 (N_52,In_613,In_409);
or U53 (N_53,In_586,In_600);
xor U54 (N_54,In_634,In_304);
or U55 (N_55,In_397,In_599);
nand U56 (N_56,In_53,In_404);
and U57 (N_57,In_352,In_415);
nor U58 (N_58,In_189,In_533);
nand U59 (N_59,In_115,In_147);
xnor U60 (N_60,In_614,In_521);
and U61 (N_61,In_266,In_82);
and U62 (N_62,In_405,In_154);
or U63 (N_63,In_342,In_591);
nand U64 (N_64,In_119,In_657);
nand U65 (N_65,In_79,In_734);
and U66 (N_66,In_510,In_693);
nor U67 (N_67,In_64,In_511);
nor U68 (N_68,In_146,In_453);
nor U69 (N_69,In_596,In_417);
and U70 (N_70,In_28,In_680);
nand U71 (N_71,In_654,In_239);
xor U72 (N_72,In_55,In_116);
nand U73 (N_73,In_349,In_207);
nand U74 (N_74,In_716,In_87);
and U75 (N_75,In_41,In_21);
or U76 (N_76,In_183,In_100);
nand U77 (N_77,In_77,In_620);
or U78 (N_78,In_627,In_619);
nor U79 (N_79,In_44,In_156);
xnor U80 (N_80,In_414,In_519);
and U81 (N_81,In_541,In_566);
nand U82 (N_82,In_257,In_265);
nor U83 (N_83,In_216,In_351);
nand U84 (N_84,In_439,In_284);
xnor U85 (N_85,In_308,In_103);
or U86 (N_86,In_466,In_603);
or U87 (N_87,In_451,In_346);
and U88 (N_88,In_626,In_555);
or U89 (N_89,In_644,In_457);
and U90 (N_90,In_393,In_261);
or U91 (N_91,In_326,In_732);
and U92 (N_92,In_675,In_323);
nor U93 (N_93,In_615,In_336);
or U94 (N_94,In_674,In_378);
xnor U95 (N_95,In_89,In_313);
nand U96 (N_96,In_497,In_344);
nor U97 (N_97,In_148,In_388);
nor U98 (N_98,In_493,In_705);
and U99 (N_99,In_500,In_656);
and U100 (N_100,In_671,In_243);
and U101 (N_101,In_425,In_205);
nand U102 (N_102,In_602,In_206);
or U103 (N_103,In_36,In_197);
and U104 (N_104,In_390,In_80);
and U105 (N_105,In_548,In_219);
and U106 (N_106,In_380,In_682);
nor U107 (N_107,In_663,In_660);
nand U108 (N_108,In_158,In_664);
nand U109 (N_109,In_162,In_576);
nand U110 (N_110,In_71,In_637);
nor U111 (N_111,In_338,In_24);
or U112 (N_112,In_502,In_129);
or U113 (N_113,In_594,In_319);
or U114 (N_114,In_413,In_362);
nand U115 (N_115,In_372,In_503);
nand U116 (N_116,In_587,In_631);
nor U117 (N_117,In_655,In_606);
nand U118 (N_118,In_101,In_402);
nand U119 (N_119,In_25,In_746);
and U120 (N_120,In_204,In_294);
nand U121 (N_121,In_505,In_94);
nand U122 (N_122,In_339,In_557);
or U123 (N_123,In_327,In_311);
nor U124 (N_124,In_666,In_552);
nand U125 (N_125,In_273,In_309);
nand U126 (N_126,In_328,In_488);
nor U127 (N_127,In_0,In_228);
and U128 (N_128,In_140,In_161);
or U129 (N_129,In_16,In_343);
and U130 (N_130,In_232,In_618);
and U131 (N_131,In_450,In_706);
xnor U132 (N_132,In_640,In_427);
nand U133 (N_133,In_32,In_727);
nor U134 (N_134,In_650,In_315);
nand U135 (N_135,In_267,In_317);
or U136 (N_136,In_499,In_105);
and U137 (N_137,In_199,In_348);
and U138 (N_138,In_260,In_702);
or U139 (N_139,In_537,In_731);
nand U140 (N_140,In_202,In_479);
or U141 (N_141,In_181,In_486);
and U142 (N_142,In_303,In_341);
and U143 (N_143,In_710,In_517);
nor U144 (N_144,In_395,In_33);
nor U145 (N_145,In_300,In_737);
nor U146 (N_146,In_509,In_258);
and U147 (N_147,In_459,In_489);
and U148 (N_148,In_93,In_120);
nor U149 (N_149,In_195,In_59);
nand U150 (N_150,In_359,In_26);
xor U151 (N_151,In_2,In_446);
nor U152 (N_152,In_691,In_320);
nor U153 (N_153,In_568,In_104);
and U154 (N_154,In_111,In_501);
nor U155 (N_155,In_696,In_551);
nor U156 (N_156,In_471,In_742);
or U157 (N_157,In_68,In_186);
and U158 (N_158,In_275,In_83);
or U159 (N_159,In_356,In_741);
nand U160 (N_160,In_5,In_289);
and U161 (N_161,In_268,In_379);
or U162 (N_162,In_163,In_329);
nor U163 (N_163,In_639,In_353);
and U164 (N_164,In_570,In_628);
and U165 (N_165,In_152,In_495);
or U166 (N_166,In_738,In_392);
nand U167 (N_167,In_612,In_22);
nand U168 (N_168,In_535,In_91);
and U169 (N_169,In_549,In_42);
nor U170 (N_170,In_556,In_74);
or U171 (N_171,In_217,In_423);
and U172 (N_172,In_301,In_234);
nand U173 (N_173,In_445,In_621);
nand U174 (N_174,In_50,In_611);
nor U175 (N_175,In_384,In_238);
or U176 (N_176,In_659,In_444);
xor U177 (N_177,In_29,In_605);
or U178 (N_178,In_667,In_553);
nand U179 (N_179,In_131,In_305);
nor U180 (N_180,In_60,In_647);
nand U181 (N_181,In_78,In_170);
or U182 (N_182,In_632,In_84);
nor U183 (N_183,In_722,In_30);
nor U184 (N_184,In_322,In_244);
or U185 (N_185,In_212,In_48);
nor U186 (N_186,In_231,In_573);
and U187 (N_187,In_730,In_564);
nor U188 (N_188,In_717,In_447);
nor U189 (N_189,In_385,In_708);
and U190 (N_190,In_173,In_295);
or U191 (N_191,In_160,In_331);
xor U192 (N_192,In_482,In_236);
and U193 (N_193,In_282,In_366);
nor U194 (N_194,In_396,In_215);
nor U195 (N_195,In_454,In_629);
nand U196 (N_196,In_504,In_473);
or U197 (N_197,In_307,In_431);
nand U198 (N_198,In_709,In_528);
nand U199 (N_199,In_610,In_364);
nand U200 (N_200,In_350,In_221);
or U201 (N_201,In_491,N_81);
nor U202 (N_202,In_184,In_441);
and U203 (N_203,N_67,N_40);
or U204 (N_204,In_264,N_77);
nor U205 (N_205,In_290,In_31);
nand U206 (N_206,N_92,In_394);
and U207 (N_207,N_20,N_136);
or U208 (N_208,N_110,In_745);
xnor U209 (N_209,N_61,In_332);
nand U210 (N_210,N_123,In_684);
xor U211 (N_211,In_561,In_165);
xor U212 (N_212,In_251,In_250);
xor U213 (N_213,In_642,In_748);
or U214 (N_214,In_547,In_124);
and U215 (N_215,In_291,N_143);
or U216 (N_216,In_428,In_45);
or U217 (N_217,N_104,In_128);
xnor U218 (N_218,In_412,In_259);
nand U219 (N_219,N_169,In_1);
nand U220 (N_220,N_9,In_408);
xor U221 (N_221,In_43,In_468);
and U222 (N_222,In_63,In_375);
and U223 (N_223,N_75,In_635);
or U224 (N_224,N_152,In_66);
nor U225 (N_225,In_410,N_165);
nand U226 (N_226,N_2,In_252);
nand U227 (N_227,In_536,In_522);
nor U228 (N_228,N_195,In_96);
nor U229 (N_229,N_6,N_72);
nor U230 (N_230,N_122,In_114);
nor U231 (N_231,N_121,N_184);
nor U232 (N_232,In_461,N_80);
nor U233 (N_233,In_278,In_192);
and U234 (N_234,N_162,N_177);
nor U235 (N_235,In_335,In_725);
and U236 (N_236,N_173,N_84);
or U237 (N_237,In_514,In_229);
or U238 (N_238,N_54,N_62);
or U239 (N_239,N_48,In_113);
nor U240 (N_240,In_530,In_692);
nand U241 (N_241,In_72,In_546);
nand U242 (N_242,N_172,In_474);
xnor U243 (N_243,N_179,N_85);
nand U244 (N_244,In_40,N_119);
and U245 (N_245,N_22,In_689);
and U246 (N_246,In_166,In_648);
nand U247 (N_247,In_595,In_543);
xnor U248 (N_248,N_111,In_224);
nand U249 (N_249,N_185,N_10);
or U250 (N_250,In_383,N_60);
nand U251 (N_251,In_287,In_88);
or U252 (N_252,In_157,In_719);
nand U253 (N_253,In_132,In_440);
nor U254 (N_254,In_70,In_75);
nand U255 (N_255,In_539,In_593);
nor U256 (N_256,N_197,N_94);
and U257 (N_257,In_525,N_187);
nand U258 (N_258,In_467,N_114);
nand U259 (N_259,N_25,N_91);
nand U260 (N_260,N_132,In_438);
nand U261 (N_261,N_141,In_527);
xor U262 (N_262,In_661,N_58);
and U263 (N_263,N_15,In_669);
or U264 (N_264,N_131,In_733);
nor U265 (N_265,N_151,In_449);
nor U266 (N_266,N_89,In_728);
nor U267 (N_267,In_578,N_101);
or U268 (N_268,In_531,In_248);
nand U269 (N_269,N_55,N_168);
nand U270 (N_270,N_186,N_28);
nor U271 (N_271,N_24,In_297);
or U272 (N_272,N_47,In_73);
and U273 (N_273,N_11,In_117);
nand U274 (N_274,N_97,N_148);
nor U275 (N_275,N_56,In_19);
or U276 (N_276,In_58,In_683);
and U277 (N_277,In_7,N_126);
or U278 (N_278,N_120,In_406);
or U279 (N_279,N_95,N_178);
or U280 (N_280,In_697,In_347);
and U281 (N_281,In_324,N_34);
nor U282 (N_282,In_118,In_592);
and U283 (N_283,N_176,In_462);
nor U284 (N_284,In_143,N_88);
nand U285 (N_285,In_256,In_609);
and U286 (N_286,In_704,In_34);
or U287 (N_287,In_191,N_139);
or U288 (N_288,In_280,In_67);
or U289 (N_289,In_518,In_560);
and U290 (N_290,In_529,In_701);
or U291 (N_291,In_373,In_62);
or U292 (N_292,In_638,In_127);
xnor U293 (N_293,In_544,N_29);
nand U294 (N_294,In_237,In_365);
nor U295 (N_295,In_203,In_677);
nor U296 (N_296,In_312,In_337);
xor U297 (N_297,In_190,N_70);
or U298 (N_298,N_26,In_729);
nand U299 (N_299,In_681,In_658);
nand U300 (N_300,In_233,In_69);
nand U301 (N_301,N_59,In_12);
and U302 (N_302,In_177,In_538);
and U303 (N_303,In_455,In_679);
nand U304 (N_304,In_506,N_157);
nor U305 (N_305,In_51,In_481);
nor U306 (N_306,In_6,In_516);
nor U307 (N_307,In_744,N_18);
nor U308 (N_308,In_263,N_31);
and U309 (N_309,In_448,In_483);
and U310 (N_310,In_139,In_92);
nor U311 (N_311,In_245,In_310);
or U312 (N_312,N_53,In_106);
or U313 (N_313,In_196,N_158);
nand U314 (N_314,In_253,In_330);
and U315 (N_315,In_678,N_189);
or U316 (N_316,N_63,N_30);
nor U317 (N_317,N_149,N_190);
and U318 (N_318,In_688,In_636);
xor U319 (N_319,N_73,In_720);
xor U320 (N_320,In_367,N_191);
and U321 (N_321,In_598,In_721);
nand U322 (N_322,N_198,In_476);
and U323 (N_323,In_65,In_141);
or U324 (N_324,In_711,In_370);
xor U325 (N_325,N_90,In_607);
and U326 (N_326,N_166,N_66);
nor U327 (N_327,In_633,In_355);
or U328 (N_328,In_579,In_218);
or U329 (N_329,N_138,In_246);
nand U330 (N_330,N_1,In_714);
and U331 (N_331,In_381,In_464);
or U332 (N_332,N_112,N_105);
nor U333 (N_333,In_589,In_698);
nand U334 (N_334,In_707,In_185);
or U335 (N_335,In_316,In_475);
and U336 (N_336,In_713,In_283);
nor U337 (N_337,In_179,N_45);
xor U338 (N_338,In_624,In_442);
nand U339 (N_339,N_36,N_130);
xnor U340 (N_340,In_276,In_357);
xor U341 (N_341,In_403,N_156);
or U342 (N_342,In_269,N_137);
or U343 (N_343,In_188,In_694);
or U344 (N_344,In_200,In_630);
xnor U345 (N_345,In_490,In_485);
nor U346 (N_346,In_302,In_735);
and U347 (N_347,In_649,In_382);
nand U348 (N_348,In_743,N_4);
nand U349 (N_349,In_622,In_507);
or U350 (N_350,In_580,In_747);
and U351 (N_351,In_123,In_662);
xor U352 (N_352,N_107,In_358);
or U353 (N_353,In_374,In_532);
or U354 (N_354,In_270,In_512);
nand U355 (N_355,In_15,In_368);
or U356 (N_356,N_32,In_174);
nand U357 (N_357,N_14,In_492);
nor U358 (N_358,N_21,In_90);
nor U359 (N_359,In_144,N_42);
nand U360 (N_360,In_340,N_159);
and U361 (N_361,N_109,N_183);
nand U362 (N_362,In_699,In_496);
or U363 (N_363,N_147,In_597);
and U364 (N_364,In_623,In_159);
nor U365 (N_365,N_79,N_174);
nand U366 (N_366,In_508,In_39);
or U367 (N_367,In_182,In_565);
or U368 (N_368,In_703,In_400);
xnor U369 (N_369,N_106,N_57);
nand U370 (N_370,In_540,In_407);
nor U371 (N_371,N_117,In_3);
nor U372 (N_372,In_515,N_118);
nor U373 (N_373,In_749,N_129);
xnor U374 (N_374,N_160,In_208);
nor U375 (N_375,In_47,N_98);
nor U376 (N_376,In_387,In_201);
nand U377 (N_377,In_240,In_463);
nand U378 (N_378,N_116,In_17);
or U379 (N_379,In_235,In_138);
or U380 (N_380,N_125,In_545);
nand U381 (N_381,In_377,N_43);
nor U382 (N_382,N_134,N_150);
or U383 (N_383,In_369,In_736);
nand U384 (N_384,In_673,In_130);
or U385 (N_385,N_16,In_584);
nand U386 (N_386,In_122,In_422);
nor U387 (N_387,N_181,In_401);
nor U388 (N_388,In_214,In_643);
nand U389 (N_389,In_11,N_23);
nand U390 (N_390,In_550,N_102);
nor U391 (N_391,In_213,In_153);
or U392 (N_392,N_144,In_526);
nor U393 (N_393,In_740,In_554);
xor U394 (N_394,N_17,N_196);
or U395 (N_395,In_126,In_164);
and U396 (N_396,In_432,N_5);
nand U397 (N_397,In_458,In_575);
and U398 (N_398,In_652,N_0);
or U399 (N_399,In_180,In_81);
and U400 (N_400,In_418,N_305);
or U401 (N_401,N_241,In_178);
nor U402 (N_402,In_672,In_360);
and U403 (N_403,N_238,N_291);
nor U404 (N_404,N_3,N_226);
or U405 (N_405,N_248,In_56);
and U406 (N_406,N_373,N_312);
nor U407 (N_407,N_309,In_171);
and U408 (N_408,N_230,N_234);
and U409 (N_409,N_207,In_651);
and U410 (N_410,In_460,In_583);
or U411 (N_411,N_188,N_154);
nor U412 (N_412,N_386,In_57);
and U413 (N_413,In_262,N_385);
nor U414 (N_414,In_487,N_365);
and U415 (N_415,N_311,In_98);
or U416 (N_416,In_321,N_327);
nor U417 (N_417,N_257,N_209);
nor U418 (N_418,N_163,N_299);
nor U419 (N_419,In_133,In_465);
nor U420 (N_420,N_326,In_223);
nor U421 (N_421,N_236,N_124);
xor U422 (N_422,In_520,N_379);
and U423 (N_423,N_351,N_115);
nand U424 (N_424,In_625,N_206);
nor U425 (N_425,In_222,N_100);
or U426 (N_426,N_322,In_411);
or U427 (N_427,In_97,In_617);
or U428 (N_428,N_243,N_357);
xnor U429 (N_429,N_19,In_361);
nor U430 (N_430,N_276,N_382);
or U431 (N_431,N_272,N_282);
nand U432 (N_432,N_389,N_330);
nand U433 (N_433,In_296,N_260);
and U434 (N_434,In_513,N_213);
and U435 (N_435,N_253,N_295);
nor U436 (N_436,N_259,N_356);
nand U437 (N_437,In_685,N_216);
xnor U438 (N_438,N_135,N_358);
and U439 (N_439,N_133,N_142);
and U440 (N_440,N_237,In_37);
or U441 (N_441,N_233,N_7);
or U442 (N_442,N_252,In_211);
or U443 (N_443,N_315,N_210);
or U444 (N_444,N_271,In_13);
and U445 (N_445,N_288,N_249);
or U446 (N_446,N_83,N_310);
nor U447 (N_447,N_333,N_337);
or U448 (N_448,In_149,N_127);
nand U449 (N_449,In_255,N_44);
xnor U450 (N_450,N_231,N_292);
and U451 (N_451,N_283,In_318);
or U452 (N_452,N_346,N_27);
nor U453 (N_453,N_167,N_372);
and U454 (N_454,N_285,N_318);
xnor U455 (N_455,N_355,N_76);
and U456 (N_456,N_203,N_52);
nor U457 (N_457,N_321,N_71);
nand U458 (N_458,N_182,N_323);
and U459 (N_459,N_13,N_201);
nor U460 (N_460,N_275,In_61);
nand U461 (N_461,N_381,N_51);
or U462 (N_462,N_265,N_263);
nand U463 (N_463,N_205,N_258);
and U464 (N_464,N_274,N_270);
and U465 (N_465,N_363,N_300);
nor U466 (N_466,N_87,In_306);
or U467 (N_467,N_342,N_352);
nand U468 (N_468,N_332,In_299);
nor U469 (N_469,N_93,N_223);
and U470 (N_470,In_715,N_281);
and U471 (N_471,In_563,N_307);
nor U472 (N_472,N_329,N_397);
and U473 (N_473,In_363,In_700);
or U474 (N_474,N_286,N_349);
and U475 (N_475,N_74,In_653);
nor U476 (N_476,N_359,N_375);
or U477 (N_477,N_279,In_376);
or U478 (N_478,N_239,In_325);
nor U479 (N_479,In_469,In_14);
nand U480 (N_480,N_217,N_38);
or U481 (N_481,N_103,In_726);
and U482 (N_482,N_214,N_99);
nor U483 (N_483,N_302,N_128);
or U484 (N_484,In_298,N_246);
and U485 (N_485,N_384,N_49);
xor U486 (N_486,N_64,N_254);
and U487 (N_487,N_261,N_278);
or U488 (N_488,N_387,N_399);
nor U489 (N_489,N_145,N_171);
xor U490 (N_490,N_180,In_137);
xnor U491 (N_491,N_350,N_227);
xor U492 (N_492,N_308,N_193);
or U493 (N_493,N_391,N_335);
or U494 (N_494,N_113,N_334);
or U495 (N_495,N_339,N_313);
or U496 (N_496,N_395,In_109);
nand U497 (N_497,N_304,In_601);
or U498 (N_498,In_134,N_398);
or U499 (N_499,N_377,In_314);
or U500 (N_500,In_54,N_362);
nand U501 (N_501,N_328,N_12);
nor U502 (N_502,N_376,N_224);
nor U503 (N_503,In_9,N_244);
and U504 (N_504,N_325,N_370);
or U505 (N_505,In_151,N_86);
and U506 (N_506,In_574,N_164);
and U507 (N_507,N_219,N_390);
or U508 (N_508,N_294,In_187);
or U509 (N_509,N_39,In_23);
nor U510 (N_510,N_245,N_82);
or U511 (N_511,N_65,N_235);
or U512 (N_512,N_394,N_204);
and U513 (N_513,N_303,In_478);
and U514 (N_514,N_37,N_277);
xnor U515 (N_515,N_242,N_262);
nor U516 (N_516,N_348,N_69);
and U517 (N_517,N_33,N_199);
nand U518 (N_518,In_354,N_211);
nor U519 (N_519,N_378,N_371);
or U520 (N_520,N_155,N_218);
xor U521 (N_521,N_343,N_78);
nand U522 (N_522,N_331,In_542);
nand U523 (N_523,N_46,N_320);
nor U524 (N_524,N_267,N_212);
nand U525 (N_525,N_269,N_266);
nand U526 (N_526,N_175,In_35);
and U527 (N_527,N_316,N_347);
or U528 (N_528,N_202,N_341);
nand U529 (N_529,N_353,N_289);
nand U530 (N_530,N_336,In_420);
nand U531 (N_531,N_290,N_369);
and U532 (N_532,N_247,N_301);
nand U533 (N_533,N_222,N_153);
nor U534 (N_534,N_225,N_221);
nand U535 (N_535,N_306,In_125);
nor U536 (N_536,In_498,N_393);
xor U537 (N_537,In_281,N_232);
nand U538 (N_538,N_108,N_361);
nor U539 (N_539,N_287,N_68);
nor U540 (N_540,In_572,N_380);
nor U541 (N_541,N_200,N_354);
nor U542 (N_542,N_240,N_220);
and U543 (N_543,N_344,N_161);
xor U544 (N_544,N_396,N_250);
and U545 (N_545,N_96,N_367);
or U546 (N_546,In_288,N_228);
nor U547 (N_547,In_452,N_140);
nand U548 (N_548,In_220,N_364);
and U549 (N_549,In_85,N_50);
nor U550 (N_550,N_192,In_641);
and U551 (N_551,N_35,N_273);
and U552 (N_552,N_345,In_292);
nor U553 (N_553,N_280,In_668);
nand U554 (N_554,N_215,In_20);
and U555 (N_555,N_293,In_484);
xor U556 (N_556,N_208,N_296);
nand U557 (N_557,N_8,N_324);
nand U558 (N_558,N_251,In_145);
xor U559 (N_559,In_76,N_366);
nand U560 (N_560,N_170,N_284);
or U561 (N_561,N_41,N_374);
or U562 (N_562,N_368,N_264);
and U563 (N_563,In_110,N_255);
or U564 (N_564,In_437,N_319);
xnor U565 (N_565,N_314,N_256);
nor U566 (N_566,N_360,In_345);
nor U567 (N_567,N_146,N_388);
nand U568 (N_568,In_226,N_340);
nand U569 (N_569,N_317,N_338);
and U570 (N_570,N_297,N_298);
nor U571 (N_571,N_383,In_52);
nand U572 (N_572,N_194,In_424);
and U573 (N_573,N_229,N_268);
nand U574 (N_574,In_523,N_392);
nor U575 (N_575,N_33,N_145);
nand U576 (N_576,N_392,N_319);
and U577 (N_577,N_142,In_345);
and U578 (N_578,In_583,In_13);
and U579 (N_579,N_35,N_305);
nand U580 (N_580,N_205,N_188);
and U581 (N_581,In_98,N_304);
nor U582 (N_582,N_113,N_322);
nor U583 (N_583,N_35,In_226);
and U584 (N_584,N_268,N_142);
and U585 (N_585,N_388,N_236);
or U586 (N_586,N_216,N_87);
xor U587 (N_587,N_243,N_49);
nor U588 (N_588,N_209,N_7);
or U589 (N_589,N_238,N_254);
or U590 (N_590,N_241,N_311);
and U591 (N_591,In_487,In_281);
or U592 (N_592,N_325,N_96);
or U593 (N_593,N_230,N_292);
xor U594 (N_594,N_65,N_268);
nor U595 (N_595,N_39,N_364);
nor U596 (N_596,N_333,In_641);
nor U597 (N_597,N_388,N_203);
or U598 (N_598,N_276,In_109);
nand U599 (N_599,N_208,N_124);
xnor U600 (N_600,N_558,N_567);
nand U601 (N_601,N_561,N_410);
nand U602 (N_602,N_463,N_449);
and U603 (N_603,N_547,N_541);
nand U604 (N_604,N_482,N_459);
or U605 (N_605,N_452,N_453);
or U606 (N_606,N_533,N_595);
and U607 (N_607,N_523,N_416);
nor U608 (N_608,N_485,N_401);
nand U609 (N_609,N_503,N_565);
nand U610 (N_610,N_516,N_458);
nand U611 (N_611,N_559,N_478);
and U612 (N_612,N_506,N_446);
and U613 (N_613,N_490,N_405);
nand U614 (N_614,N_487,N_493);
nand U615 (N_615,N_504,N_512);
nand U616 (N_616,N_423,N_414);
xnor U617 (N_617,N_492,N_435);
nor U618 (N_618,N_587,N_467);
or U619 (N_619,N_424,N_545);
nand U620 (N_620,N_593,N_477);
nand U621 (N_621,N_481,N_419);
nand U622 (N_622,N_422,N_454);
nand U623 (N_623,N_542,N_421);
nand U624 (N_624,N_576,N_520);
nand U625 (N_625,N_447,N_577);
nand U626 (N_626,N_497,N_511);
nor U627 (N_627,N_457,N_578);
and U628 (N_628,N_486,N_568);
and U629 (N_629,N_498,N_592);
nor U630 (N_630,N_515,N_584);
nand U631 (N_631,N_473,N_495);
nand U632 (N_632,N_552,N_469);
nor U633 (N_633,N_500,N_427);
or U634 (N_634,N_501,N_536);
and U635 (N_635,N_570,N_403);
and U636 (N_636,N_594,N_466);
and U637 (N_637,N_583,N_589);
and U638 (N_638,N_551,N_445);
and U639 (N_639,N_585,N_433);
nor U640 (N_640,N_409,N_573);
nand U641 (N_641,N_417,N_598);
nand U642 (N_642,N_555,N_451);
and U643 (N_643,N_480,N_455);
and U644 (N_644,N_509,N_596);
xnor U645 (N_645,N_525,N_579);
nand U646 (N_646,N_462,N_513);
nor U647 (N_647,N_425,N_574);
or U648 (N_648,N_468,N_438);
or U649 (N_649,N_441,N_566);
or U650 (N_650,N_434,N_538);
nor U651 (N_651,N_560,N_571);
nand U652 (N_652,N_562,N_460);
and U653 (N_653,N_471,N_586);
or U654 (N_654,N_588,N_575);
or U655 (N_655,N_554,N_564);
or U656 (N_656,N_450,N_510);
xor U657 (N_657,N_428,N_431);
and U658 (N_658,N_444,N_549);
or U659 (N_659,N_507,N_563);
or U660 (N_660,N_443,N_436);
nand U661 (N_661,N_437,N_476);
nand U662 (N_662,N_537,N_569);
nand U663 (N_663,N_475,N_556);
and U664 (N_664,N_429,N_530);
xnor U665 (N_665,N_532,N_521);
nor U666 (N_666,N_517,N_546);
nor U667 (N_667,N_524,N_550);
xnor U668 (N_668,N_580,N_548);
and U669 (N_669,N_599,N_465);
and U670 (N_670,N_432,N_514);
nand U671 (N_671,N_406,N_502);
nor U672 (N_672,N_411,N_543);
nor U673 (N_673,N_420,N_489);
xnor U674 (N_674,N_553,N_519);
nor U675 (N_675,N_582,N_535);
and U676 (N_676,N_400,N_540);
nor U677 (N_677,N_456,N_479);
or U678 (N_678,N_531,N_461);
or U679 (N_679,N_412,N_470);
xnor U680 (N_680,N_442,N_464);
or U681 (N_681,N_408,N_526);
or U682 (N_682,N_539,N_529);
nand U683 (N_683,N_581,N_590);
and U684 (N_684,N_518,N_415);
xor U685 (N_685,N_426,N_557);
or U686 (N_686,N_499,N_528);
or U687 (N_687,N_544,N_488);
and U688 (N_688,N_505,N_430);
or U689 (N_689,N_404,N_591);
nor U690 (N_690,N_534,N_527);
and U691 (N_691,N_484,N_572);
nand U692 (N_692,N_407,N_440);
and U693 (N_693,N_491,N_496);
nand U694 (N_694,N_439,N_494);
and U695 (N_695,N_508,N_413);
xor U696 (N_696,N_472,N_483);
or U697 (N_697,N_522,N_448);
nor U698 (N_698,N_474,N_402);
or U699 (N_699,N_418,N_597);
nand U700 (N_700,N_419,N_431);
or U701 (N_701,N_479,N_536);
nand U702 (N_702,N_539,N_452);
nor U703 (N_703,N_460,N_507);
and U704 (N_704,N_541,N_429);
nor U705 (N_705,N_466,N_533);
or U706 (N_706,N_427,N_560);
nor U707 (N_707,N_419,N_524);
nor U708 (N_708,N_555,N_489);
or U709 (N_709,N_594,N_549);
and U710 (N_710,N_469,N_551);
nor U711 (N_711,N_591,N_415);
xnor U712 (N_712,N_521,N_510);
or U713 (N_713,N_557,N_522);
nand U714 (N_714,N_506,N_550);
nand U715 (N_715,N_409,N_402);
nor U716 (N_716,N_403,N_513);
nand U717 (N_717,N_499,N_491);
nor U718 (N_718,N_495,N_497);
and U719 (N_719,N_571,N_438);
nor U720 (N_720,N_515,N_449);
and U721 (N_721,N_526,N_436);
nor U722 (N_722,N_446,N_460);
nand U723 (N_723,N_581,N_564);
and U724 (N_724,N_491,N_564);
and U725 (N_725,N_544,N_577);
and U726 (N_726,N_418,N_462);
nand U727 (N_727,N_418,N_572);
nor U728 (N_728,N_558,N_591);
and U729 (N_729,N_480,N_458);
and U730 (N_730,N_556,N_575);
xor U731 (N_731,N_447,N_535);
nor U732 (N_732,N_401,N_543);
nand U733 (N_733,N_591,N_486);
xor U734 (N_734,N_482,N_557);
and U735 (N_735,N_515,N_488);
nand U736 (N_736,N_466,N_544);
nor U737 (N_737,N_439,N_459);
or U738 (N_738,N_414,N_528);
nand U739 (N_739,N_407,N_442);
and U740 (N_740,N_590,N_427);
and U741 (N_741,N_411,N_506);
nand U742 (N_742,N_543,N_432);
or U743 (N_743,N_542,N_406);
nand U744 (N_744,N_402,N_523);
and U745 (N_745,N_598,N_570);
and U746 (N_746,N_569,N_416);
and U747 (N_747,N_531,N_494);
and U748 (N_748,N_510,N_597);
nand U749 (N_749,N_583,N_514);
or U750 (N_750,N_472,N_546);
nor U751 (N_751,N_437,N_514);
and U752 (N_752,N_543,N_537);
or U753 (N_753,N_459,N_522);
or U754 (N_754,N_409,N_541);
nand U755 (N_755,N_493,N_525);
or U756 (N_756,N_568,N_426);
nor U757 (N_757,N_520,N_570);
or U758 (N_758,N_403,N_567);
nor U759 (N_759,N_569,N_489);
xnor U760 (N_760,N_546,N_407);
or U761 (N_761,N_439,N_456);
and U762 (N_762,N_436,N_453);
xnor U763 (N_763,N_458,N_540);
or U764 (N_764,N_462,N_533);
xnor U765 (N_765,N_411,N_466);
and U766 (N_766,N_484,N_465);
nor U767 (N_767,N_586,N_503);
xor U768 (N_768,N_582,N_593);
nand U769 (N_769,N_588,N_480);
nand U770 (N_770,N_479,N_537);
or U771 (N_771,N_547,N_475);
and U772 (N_772,N_498,N_469);
and U773 (N_773,N_520,N_519);
nor U774 (N_774,N_424,N_428);
nor U775 (N_775,N_526,N_472);
or U776 (N_776,N_523,N_544);
and U777 (N_777,N_406,N_494);
nand U778 (N_778,N_587,N_522);
or U779 (N_779,N_475,N_483);
nand U780 (N_780,N_440,N_404);
nor U781 (N_781,N_480,N_424);
and U782 (N_782,N_443,N_512);
or U783 (N_783,N_570,N_422);
nand U784 (N_784,N_591,N_581);
and U785 (N_785,N_460,N_406);
nand U786 (N_786,N_549,N_453);
nand U787 (N_787,N_445,N_414);
and U788 (N_788,N_462,N_435);
and U789 (N_789,N_405,N_491);
and U790 (N_790,N_410,N_438);
nor U791 (N_791,N_481,N_517);
nand U792 (N_792,N_570,N_458);
and U793 (N_793,N_449,N_520);
nor U794 (N_794,N_599,N_598);
nor U795 (N_795,N_436,N_570);
nand U796 (N_796,N_488,N_576);
or U797 (N_797,N_457,N_504);
and U798 (N_798,N_551,N_511);
or U799 (N_799,N_595,N_557);
and U800 (N_800,N_745,N_730);
and U801 (N_801,N_659,N_654);
and U802 (N_802,N_667,N_738);
nand U803 (N_803,N_622,N_739);
nor U804 (N_804,N_657,N_767);
xor U805 (N_805,N_630,N_747);
or U806 (N_806,N_719,N_736);
and U807 (N_807,N_639,N_742);
nor U808 (N_808,N_610,N_611);
or U809 (N_809,N_766,N_685);
or U810 (N_810,N_702,N_662);
xor U811 (N_811,N_640,N_712);
nand U812 (N_812,N_614,N_629);
nand U813 (N_813,N_791,N_613);
or U814 (N_814,N_704,N_780);
and U815 (N_815,N_644,N_760);
and U816 (N_816,N_792,N_675);
or U817 (N_817,N_713,N_625);
and U818 (N_818,N_690,N_751);
xor U819 (N_819,N_705,N_627);
or U820 (N_820,N_703,N_683);
and U821 (N_821,N_686,N_774);
xor U822 (N_822,N_664,N_660);
nor U823 (N_823,N_727,N_612);
nand U824 (N_824,N_626,N_600);
nor U825 (N_825,N_618,N_765);
nor U826 (N_826,N_726,N_775);
or U827 (N_827,N_773,N_744);
and U828 (N_828,N_638,N_663);
nor U829 (N_829,N_634,N_688);
xnor U830 (N_830,N_794,N_670);
nand U831 (N_831,N_731,N_759);
and U832 (N_832,N_734,N_674);
nor U833 (N_833,N_620,N_715);
or U834 (N_834,N_782,N_682);
nor U835 (N_835,N_786,N_741);
and U836 (N_836,N_758,N_615);
nor U837 (N_837,N_604,N_680);
nand U838 (N_838,N_743,N_795);
nor U839 (N_839,N_645,N_768);
nor U840 (N_840,N_673,N_684);
nor U841 (N_841,N_710,N_776);
or U842 (N_842,N_716,N_706);
nand U843 (N_843,N_652,N_636);
or U844 (N_844,N_732,N_658);
nand U845 (N_845,N_770,N_616);
xor U846 (N_846,N_756,N_619);
nor U847 (N_847,N_608,N_681);
and U848 (N_848,N_799,N_749);
nor U849 (N_849,N_725,N_717);
nor U850 (N_850,N_602,N_735);
and U851 (N_851,N_790,N_755);
or U852 (N_852,N_781,N_796);
xor U853 (N_853,N_607,N_752);
nand U854 (N_854,N_798,N_707);
and U855 (N_855,N_665,N_623);
xor U856 (N_856,N_723,N_694);
or U857 (N_857,N_721,N_624);
and U858 (N_858,N_720,N_661);
nor U859 (N_859,N_653,N_711);
nor U860 (N_860,N_698,N_646);
and U861 (N_861,N_637,N_648);
nand U862 (N_862,N_763,N_695);
or U863 (N_863,N_650,N_671);
and U864 (N_864,N_693,N_757);
nand U865 (N_865,N_632,N_609);
nor U866 (N_866,N_655,N_679);
or U867 (N_867,N_746,N_606);
and U868 (N_868,N_678,N_687);
nor U869 (N_869,N_777,N_788);
and U870 (N_870,N_651,N_601);
xnor U871 (N_871,N_696,N_697);
nand U872 (N_872,N_691,N_643);
and U873 (N_873,N_722,N_754);
or U874 (N_874,N_787,N_797);
or U875 (N_875,N_793,N_633);
and U876 (N_876,N_631,N_762);
nand U877 (N_877,N_769,N_668);
nand U878 (N_878,N_669,N_605);
or U879 (N_879,N_772,N_709);
nor U880 (N_880,N_701,N_649);
nand U881 (N_881,N_677,N_729);
or U882 (N_882,N_714,N_740);
and U883 (N_883,N_641,N_603);
nor U884 (N_884,N_699,N_617);
nor U885 (N_885,N_750,N_748);
nor U886 (N_886,N_753,N_771);
nor U887 (N_887,N_666,N_764);
nand U888 (N_888,N_761,N_656);
nor U889 (N_889,N_728,N_635);
nand U890 (N_890,N_789,N_784);
and U891 (N_891,N_692,N_778);
nand U892 (N_892,N_737,N_779);
or U893 (N_893,N_708,N_647);
nor U894 (N_894,N_676,N_733);
nand U895 (N_895,N_689,N_642);
or U896 (N_896,N_672,N_783);
xor U897 (N_897,N_724,N_718);
or U898 (N_898,N_628,N_621);
or U899 (N_899,N_700,N_785);
nand U900 (N_900,N_633,N_755);
nand U901 (N_901,N_662,N_634);
and U902 (N_902,N_614,N_613);
and U903 (N_903,N_656,N_650);
xor U904 (N_904,N_635,N_745);
nor U905 (N_905,N_613,N_601);
nand U906 (N_906,N_601,N_656);
xnor U907 (N_907,N_764,N_629);
and U908 (N_908,N_693,N_736);
and U909 (N_909,N_672,N_785);
nor U910 (N_910,N_678,N_683);
xor U911 (N_911,N_624,N_628);
and U912 (N_912,N_600,N_671);
nor U913 (N_913,N_759,N_718);
and U914 (N_914,N_793,N_601);
and U915 (N_915,N_705,N_739);
and U916 (N_916,N_653,N_797);
or U917 (N_917,N_652,N_721);
nor U918 (N_918,N_700,N_779);
or U919 (N_919,N_757,N_604);
nand U920 (N_920,N_706,N_727);
or U921 (N_921,N_767,N_734);
or U922 (N_922,N_762,N_659);
or U923 (N_923,N_780,N_645);
nor U924 (N_924,N_693,N_756);
nand U925 (N_925,N_694,N_734);
and U926 (N_926,N_702,N_749);
nor U927 (N_927,N_773,N_708);
xnor U928 (N_928,N_798,N_726);
nand U929 (N_929,N_648,N_634);
nand U930 (N_930,N_713,N_720);
nand U931 (N_931,N_647,N_788);
nor U932 (N_932,N_793,N_770);
nand U933 (N_933,N_720,N_746);
nand U934 (N_934,N_659,N_691);
or U935 (N_935,N_606,N_773);
or U936 (N_936,N_736,N_723);
and U937 (N_937,N_758,N_764);
or U938 (N_938,N_643,N_796);
nor U939 (N_939,N_709,N_649);
xnor U940 (N_940,N_685,N_756);
and U941 (N_941,N_648,N_684);
or U942 (N_942,N_664,N_768);
xor U943 (N_943,N_734,N_606);
and U944 (N_944,N_737,N_712);
nor U945 (N_945,N_600,N_723);
and U946 (N_946,N_783,N_774);
and U947 (N_947,N_620,N_797);
nor U948 (N_948,N_714,N_631);
nand U949 (N_949,N_702,N_761);
nand U950 (N_950,N_745,N_634);
nor U951 (N_951,N_738,N_791);
or U952 (N_952,N_768,N_612);
and U953 (N_953,N_670,N_667);
and U954 (N_954,N_608,N_774);
nor U955 (N_955,N_685,N_662);
nand U956 (N_956,N_694,N_766);
nand U957 (N_957,N_614,N_790);
nor U958 (N_958,N_733,N_687);
or U959 (N_959,N_705,N_664);
nor U960 (N_960,N_747,N_654);
nor U961 (N_961,N_737,N_610);
or U962 (N_962,N_741,N_766);
nor U963 (N_963,N_762,N_666);
or U964 (N_964,N_767,N_693);
and U965 (N_965,N_724,N_612);
nor U966 (N_966,N_749,N_648);
nand U967 (N_967,N_650,N_773);
nand U968 (N_968,N_758,N_609);
nand U969 (N_969,N_748,N_751);
nor U970 (N_970,N_727,N_616);
or U971 (N_971,N_770,N_780);
nor U972 (N_972,N_638,N_794);
or U973 (N_973,N_724,N_670);
xnor U974 (N_974,N_630,N_637);
or U975 (N_975,N_625,N_745);
and U976 (N_976,N_606,N_626);
or U977 (N_977,N_643,N_697);
or U978 (N_978,N_661,N_674);
nand U979 (N_979,N_678,N_738);
and U980 (N_980,N_771,N_689);
nand U981 (N_981,N_769,N_637);
or U982 (N_982,N_711,N_641);
and U983 (N_983,N_744,N_650);
nor U984 (N_984,N_761,N_651);
nand U985 (N_985,N_664,N_656);
and U986 (N_986,N_778,N_655);
or U987 (N_987,N_621,N_718);
or U988 (N_988,N_703,N_607);
nand U989 (N_989,N_778,N_645);
and U990 (N_990,N_642,N_674);
and U991 (N_991,N_734,N_681);
nand U992 (N_992,N_610,N_717);
or U993 (N_993,N_614,N_745);
or U994 (N_994,N_772,N_741);
and U995 (N_995,N_773,N_672);
nand U996 (N_996,N_697,N_778);
xor U997 (N_997,N_648,N_775);
and U998 (N_998,N_738,N_625);
and U999 (N_999,N_664,N_637);
or U1000 (N_1000,N_923,N_974);
nand U1001 (N_1001,N_946,N_924);
and U1002 (N_1002,N_952,N_840);
and U1003 (N_1003,N_854,N_913);
and U1004 (N_1004,N_837,N_841);
nand U1005 (N_1005,N_908,N_848);
nand U1006 (N_1006,N_811,N_879);
xor U1007 (N_1007,N_806,N_907);
xnor U1008 (N_1008,N_885,N_860);
nand U1009 (N_1009,N_951,N_916);
nor U1010 (N_1010,N_972,N_973);
nand U1011 (N_1011,N_851,N_932);
and U1012 (N_1012,N_877,N_939);
xnor U1013 (N_1013,N_850,N_998);
or U1014 (N_1014,N_993,N_991);
nor U1015 (N_1015,N_988,N_938);
or U1016 (N_1016,N_810,N_893);
or U1017 (N_1017,N_958,N_844);
nand U1018 (N_1018,N_813,N_956);
nor U1019 (N_1019,N_870,N_809);
or U1020 (N_1020,N_803,N_970);
and U1021 (N_1021,N_999,N_947);
and U1022 (N_1022,N_890,N_819);
or U1023 (N_1023,N_839,N_979);
or U1024 (N_1024,N_981,N_836);
or U1025 (N_1025,N_889,N_884);
or U1026 (N_1026,N_928,N_950);
nand U1027 (N_1027,N_962,N_982);
or U1028 (N_1028,N_895,N_849);
and U1029 (N_1029,N_888,N_818);
nor U1030 (N_1030,N_904,N_905);
or U1031 (N_1031,N_978,N_915);
or U1032 (N_1032,N_949,N_825);
nor U1033 (N_1033,N_846,N_968);
nor U1034 (N_1034,N_994,N_874);
xnor U1035 (N_1035,N_808,N_927);
or U1036 (N_1036,N_983,N_990);
nand U1037 (N_1037,N_901,N_826);
xor U1038 (N_1038,N_802,N_801);
and U1039 (N_1039,N_976,N_900);
and U1040 (N_1040,N_896,N_920);
and U1041 (N_1041,N_820,N_912);
or U1042 (N_1042,N_859,N_892);
or U1043 (N_1043,N_984,N_922);
or U1044 (N_1044,N_975,N_882);
nand U1045 (N_1045,N_963,N_891);
or U1046 (N_1046,N_814,N_943);
xnor U1047 (N_1047,N_971,N_842);
and U1048 (N_1048,N_858,N_847);
nand U1049 (N_1049,N_902,N_996);
or U1050 (N_1050,N_873,N_961);
xnor U1051 (N_1051,N_866,N_880);
nor U1052 (N_1052,N_887,N_955);
and U1053 (N_1053,N_987,N_800);
nand U1054 (N_1054,N_948,N_992);
xnor U1055 (N_1055,N_824,N_995);
nor U1056 (N_1056,N_812,N_989);
and U1057 (N_1057,N_899,N_965);
nor U1058 (N_1058,N_934,N_940);
xnor U1059 (N_1059,N_857,N_821);
xnor U1060 (N_1060,N_834,N_898);
or U1061 (N_1061,N_822,N_827);
nand U1062 (N_1062,N_862,N_871);
or U1063 (N_1063,N_816,N_830);
nor U1064 (N_1064,N_852,N_855);
nor U1065 (N_1065,N_967,N_828);
or U1066 (N_1066,N_933,N_966);
or U1067 (N_1067,N_864,N_817);
xnor U1068 (N_1068,N_833,N_917);
or U1069 (N_1069,N_960,N_853);
and U1070 (N_1070,N_845,N_964);
nor U1071 (N_1071,N_823,N_931);
and U1072 (N_1072,N_804,N_881);
xor U1073 (N_1073,N_838,N_835);
nand U1074 (N_1074,N_906,N_897);
nor U1075 (N_1075,N_894,N_930);
or U1076 (N_1076,N_867,N_926);
or U1077 (N_1077,N_883,N_876);
nor U1078 (N_1078,N_959,N_953);
nor U1079 (N_1079,N_986,N_980);
nand U1080 (N_1080,N_868,N_997);
and U1081 (N_1081,N_957,N_969);
and U1082 (N_1082,N_942,N_985);
nor U1083 (N_1083,N_815,N_903);
nor U1084 (N_1084,N_829,N_909);
nand U1085 (N_1085,N_936,N_832);
and U1086 (N_1086,N_911,N_878);
nand U1087 (N_1087,N_869,N_954);
nor U1088 (N_1088,N_807,N_914);
or U1089 (N_1089,N_941,N_919);
nand U1090 (N_1090,N_872,N_843);
nand U1091 (N_1091,N_925,N_875);
nor U1092 (N_1092,N_977,N_856);
or U1093 (N_1093,N_918,N_921);
nand U1094 (N_1094,N_805,N_944);
nor U1095 (N_1095,N_937,N_910);
nor U1096 (N_1096,N_945,N_861);
and U1097 (N_1097,N_865,N_935);
and U1098 (N_1098,N_831,N_863);
or U1099 (N_1099,N_886,N_929);
nor U1100 (N_1100,N_976,N_856);
nor U1101 (N_1101,N_900,N_891);
and U1102 (N_1102,N_831,N_805);
xor U1103 (N_1103,N_975,N_811);
nand U1104 (N_1104,N_946,N_834);
and U1105 (N_1105,N_874,N_854);
nand U1106 (N_1106,N_979,N_826);
xnor U1107 (N_1107,N_941,N_908);
nor U1108 (N_1108,N_829,N_891);
nor U1109 (N_1109,N_975,N_932);
or U1110 (N_1110,N_910,N_853);
nand U1111 (N_1111,N_949,N_943);
nand U1112 (N_1112,N_981,N_864);
or U1113 (N_1113,N_846,N_875);
xnor U1114 (N_1114,N_857,N_854);
nor U1115 (N_1115,N_820,N_963);
nor U1116 (N_1116,N_992,N_962);
nor U1117 (N_1117,N_855,N_806);
xor U1118 (N_1118,N_903,N_832);
nor U1119 (N_1119,N_847,N_840);
nor U1120 (N_1120,N_852,N_885);
nand U1121 (N_1121,N_984,N_935);
and U1122 (N_1122,N_823,N_857);
nor U1123 (N_1123,N_882,N_923);
or U1124 (N_1124,N_915,N_831);
and U1125 (N_1125,N_934,N_868);
nor U1126 (N_1126,N_963,N_920);
nand U1127 (N_1127,N_850,N_944);
or U1128 (N_1128,N_892,N_983);
and U1129 (N_1129,N_922,N_930);
and U1130 (N_1130,N_810,N_924);
or U1131 (N_1131,N_891,N_932);
or U1132 (N_1132,N_974,N_898);
nor U1133 (N_1133,N_887,N_961);
nor U1134 (N_1134,N_935,N_899);
nor U1135 (N_1135,N_910,N_833);
nor U1136 (N_1136,N_924,N_959);
and U1137 (N_1137,N_927,N_948);
nand U1138 (N_1138,N_903,N_845);
and U1139 (N_1139,N_838,N_947);
nand U1140 (N_1140,N_978,N_906);
and U1141 (N_1141,N_810,N_902);
or U1142 (N_1142,N_984,N_954);
and U1143 (N_1143,N_870,N_958);
nor U1144 (N_1144,N_854,N_844);
nor U1145 (N_1145,N_907,N_883);
nand U1146 (N_1146,N_968,N_857);
or U1147 (N_1147,N_988,N_985);
nor U1148 (N_1148,N_861,N_934);
nand U1149 (N_1149,N_842,N_934);
nand U1150 (N_1150,N_906,N_867);
nand U1151 (N_1151,N_882,N_988);
nor U1152 (N_1152,N_886,N_848);
nor U1153 (N_1153,N_918,N_969);
nor U1154 (N_1154,N_917,N_878);
or U1155 (N_1155,N_982,N_949);
nor U1156 (N_1156,N_855,N_897);
xor U1157 (N_1157,N_853,N_859);
and U1158 (N_1158,N_936,N_930);
nand U1159 (N_1159,N_939,N_841);
and U1160 (N_1160,N_874,N_857);
and U1161 (N_1161,N_821,N_995);
or U1162 (N_1162,N_954,N_990);
nor U1163 (N_1163,N_991,N_949);
or U1164 (N_1164,N_953,N_941);
nor U1165 (N_1165,N_912,N_880);
nor U1166 (N_1166,N_951,N_953);
or U1167 (N_1167,N_808,N_973);
nand U1168 (N_1168,N_912,N_803);
xor U1169 (N_1169,N_948,N_981);
xnor U1170 (N_1170,N_956,N_982);
nor U1171 (N_1171,N_891,N_867);
xnor U1172 (N_1172,N_810,N_903);
or U1173 (N_1173,N_835,N_995);
and U1174 (N_1174,N_990,N_902);
and U1175 (N_1175,N_996,N_942);
and U1176 (N_1176,N_861,N_831);
nand U1177 (N_1177,N_901,N_844);
nand U1178 (N_1178,N_930,N_825);
or U1179 (N_1179,N_908,N_955);
nor U1180 (N_1180,N_890,N_944);
or U1181 (N_1181,N_845,N_829);
nand U1182 (N_1182,N_946,N_849);
nor U1183 (N_1183,N_998,N_812);
nand U1184 (N_1184,N_822,N_901);
nor U1185 (N_1185,N_968,N_919);
nand U1186 (N_1186,N_812,N_940);
xor U1187 (N_1187,N_838,N_844);
xor U1188 (N_1188,N_932,N_938);
and U1189 (N_1189,N_817,N_900);
xor U1190 (N_1190,N_857,N_970);
or U1191 (N_1191,N_995,N_817);
nand U1192 (N_1192,N_966,N_858);
and U1193 (N_1193,N_991,N_935);
xor U1194 (N_1194,N_916,N_841);
nor U1195 (N_1195,N_928,N_830);
xor U1196 (N_1196,N_871,N_818);
or U1197 (N_1197,N_874,N_946);
nor U1198 (N_1198,N_938,N_854);
nand U1199 (N_1199,N_915,N_929);
nor U1200 (N_1200,N_1165,N_1067);
and U1201 (N_1201,N_1008,N_1180);
nor U1202 (N_1202,N_1115,N_1184);
or U1203 (N_1203,N_1199,N_1036);
or U1204 (N_1204,N_1113,N_1197);
xor U1205 (N_1205,N_1017,N_1001);
and U1206 (N_1206,N_1040,N_1019);
or U1207 (N_1207,N_1130,N_1049);
nand U1208 (N_1208,N_1077,N_1102);
and U1209 (N_1209,N_1046,N_1093);
and U1210 (N_1210,N_1069,N_1150);
nand U1211 (N_1211,N_1052,N_1138);
xnor U1212 (N_1212,N_1072,N_1182);
nor U1213 (N_1213,N_1034,N_1033);
and U1214 (N_1214,N_1153,N_1122);
and U1215 (N_1215,N_1063,N_1000);
nand U1216 (N_1216,N_1170,N_1148);
or U1217 (N_1217,N_1075,N_1112);
nand U1218 (N_1218,N_1070,N_1065);
nor U1219 (N_1219,N_1198,N_1190);
nand U1220 (N_1220,N_1038,N_1041);
and U1221 (N_1221,N_1010,N_1079);
nor U1222 (N_1222,N_1128,N_1022);
or U1223 (N_1223,N_1045,N_1162);
nand U1224 (N_1224,N_1032,N_1082);
and U1225 (N_1225,N_1014,N_1133);
and U1226 (N_1226,N_1191,N_1071);
xor U1227 (N_1227,N_1178,N_1107);
and U1228 (N_1228,N_1146,N_1193);
and U1229 (N_1229,N_1064,N_1059);
and U1230 (N_1230,N_1066,N_1195);
xor U1231 (N_1231,N_1152,N_1062);
or U1232 (N_1232,N_1140,N_1120);
nand U1233 (N_1233,N_1196,N_1096);
and U1234 (N_1234,N_1157,N_1188);
and U1235 (N_1235,N_1078,N_1176);
xnor U1236 (N_1236,N_1051,N_1137);
nor U1237 (N_1237,N_1095,N_1013);
nor U1238 (N_1238,N_1100,N_1085);
nor U1239 (N_1239,N_1088,N_1117);
and U1240 (N_1240,N_1054,N_1183);
and U1241 (N_1241,N_1101,N_1109);
nor U1242 (N_1242,N_1099,N_1149);
nand U1243 (N_1243,N_1121,N_1098);
xor U1244 (N_1244,N_1159,N_1123);
nor U1245 (N_1245,N_1136,N_1134);
nand U1246 (N_1246,N_1073,N_1015);
or U1247 (N_1247,N_1110,N_1005);
or U1248 (N_1248,N_1158,N_1053);
and U1249 (N_1249,N_1192,N_1141);
or U1250 (N_1250,N_1127,N_1081);
nor U1251 (N_1251,N_1025,N_1104);
and U1252 (N_1252,N_1028,N_1105);
and U1253 (N_1253,N_1163,N_1131);
nor U1254 (N_1254,N_1189,N_1076);
nand U1255 (N_1255,N_1181,N_1090);
nor U1256 (N_1256,N_1151,N_1009);
nand U1257 (N_1257,N_1175,N_1160);
nand U1258 (N_1258,N_1171,N_1023);
nor U1259 (N_1259,N_1166,N_1132);
or U1260 (N_1260,N_1089,N_1068);
nand U1261 (N_1261,N_1050,N_1080);
and U1262 (N_1262,N_1016,N_1021);
nor U1263 (N_1263,N_1057,N_1004);
nand U1264 (N_1264,N_1031,N_1048);
or U1265 (N_1265,N_1111,N_1126);
and U1266 (N_1266,N_1055,N_1020);
xnor U1267 (N_1267,N_1167,N_1083);
and U1268 (N_1268,N_1145,N_1047);
and U1269 (N_1269,N_1035,N_1042);
or U1270 (N_1270,N_1087,N_1177);
nor U1271 (N_1271,N_1125,N_1114);
nand U1272 (N_1272,N_1139,N_1147);
or U1273 (N_1273,N_1161,N_1179);
nand U1274 (N_1274,N_1012,N_1187);
xor U1275 (N_1275,N_1030,N_1044);
nand U1276 (N_1276,N_1164,N_1086);
nor U1277 (N_1277,N_1039,N_1027);
or U1278 (N_1278,N_1097,N_1003);
and U1279 (N_1279,N_1194,N_1058);
or U1280 (N_1280,N_1154,N_1168);
and U1281 (N_1281,N_1007,N_1118);
and U1282 (N_1282,N_1172,N_1106);
and U1283 (N_1283,N_1018,N_1116);
nand U1284 (N_1284,N_1143,N_1142);
xor U1285 (N_1285,N_1119,N_1026);
nor U1286 (N_1286,N_1186,N_1043);
xnor U1287 (N_1287,N_1002,N_1174);
or U1288 (N_1288,N_1173,N_1129);
and U1289 (N_1289,N_1011,N_1084);
or U1290 (N_1290,N_1155,N_1108);
nand U1291 (N_1291,N_1061,N_1135);
and U1292 (N_1292,N_1185,N_1029);
or U1293 (N_1293,N_1091,N_1144);
nor U1294 (N_1294,N_1024,N_1169);
or U1295 (N_1295,N_1124,N_1060);
or U1296 (N_1296,N_1094,N_1103);
nand U1297 (N_1297,N_1074,N_1037);
nor U1298 (N_1298,N_1056,N_1156);
or U1299 (N_1299,N_1006,N_1092);
or U1300 (N_1300,N_1080,N_1101);
nor U1301 (N_1301,N_1093,N_1017);
and U1302 (N_1302,N_1145,N_1019);
xor U1303 (N_1303,N_1000,N_1057);
and U1304 (N_1304,N_1191,N_1027);
or U1305 (N_1305,N_1112,N_1016);
xnor U1306 (N_1306,N_1174,N_1181);
nor U1307 (N_1307,N_1064,N_1066);
and U1308 (N_1308,N_1199,N_1133);
nand U1309 (N_1309,N_1188,N_1149);
nor U1310 (N_1310,N_1190,N_1195);
nor U1311 (N_1311,N_1137,N_1064);
xor U1312 (N_1312,N_1108,N_1164);
or U1313 (N_1313,N_1081,N_1047);
xor U1314 (N_1314,N_1130,N_1171);
nand U1315 (N_1315,N_1000,N_1008);
or U1316 (N_1316,N_1062,N_1012);
and U1317 (N_1317,N_1199,N_1066);
and U1318 (N_1318,N_1013,N_1178);
nor U1319 (N_1319,N_1174,N_1019);
nor U1320 (N_1320,N_1103,N_1098);
and U1321 (N_1321,N_1116,N_1151);
xor U1322 (N_1322,N_1147,N_1001);
and U1323 (N_1323,N_1099,N_1041);
nor U1324 (N_1324,N_1056,N_1006);
or U1325 (N_1325,N_1148,N_1001);
and U1326 (N_1326,N_1080,N_1135);
and U1327 (N_1327,N_1067,N_1080);
nand U1328 (N_1328,N_1067,N_1168);
nor U1329 (N_1329,N_1167,N_1125);
or U1330 (N_1330,N_1110,N_1128);
or U1331 (N_1331,N_1021,N_1077);
or U1332 (N_1332,N_1152,N_1181);
and U1333 (N_1333,N_1099,N_1184);
or U1334 (N_1334,N_1096,N_1192);
and U1335 (N_1335,N_1182,N_1025);
nand U1336 (N_1336,N_1079,N_1124);
nand U1337 (N_1337,N_1061,N_1113);
or U1338 (N_1338,N_1060,N_1090);
nor U1339 (N_1339,N_1006,N_1100);
and U1340 (N_1340,N_1021,N_1136);
nor U1341 (N_1341,N_1073,N_1142);
and U1342 (N_1342,N_1009,N_1007);
nand U1343 (N_1343,N_1069,N_1084);
nand U1344 (N_1344,N_1009,N_1155);
nor U1345 (N_1345,N_1012,N_1027);
or U1346 (N_1346,N_1102,N_1114);
nor U1347 (N_1347,N_1096,N_1121);
nand U1348 (N_1348,N_1179,N_1157);
nor U1349 (N_1349,N_1079,N_1047);
and U1350 (N_1350,N_1186,N_1103);
nor U1351 (N_1351,N_1082,N_1128);
xnor U1352 (N_1352,N_1110,N_1072);
xnor U1353 (N_1353,N_1161,N_1017);
nor U1354 (N_1354,N_1173,N_1104);
nor U1355 (N_1355,N_1165,N_1058);
nor U1356 (N_1356,N_1162,N_1154);
or U1357 (N_1357,N_1186,N_1051);
nand U1358 (N_1358,N_1053,N_1073);
or U1359 (N_1359,N_1161,N_1186);
nand U1360 (N_1360,N_1163,N_1023);
nor U1361 (N_1361,N_1097,N_1181);
nand U1362 (N_1362,N_1080,N_1071);
nor U1363 (N_1363,N_1036,N_1078);
nor U1364 (N_1364,N_1014,N_1092);
nand U1365 (N_1365,N_1008,N_1192);
and U1366 (N_1366,N_1155,N_1016);
and U1367 (N_1367,N_1088,N_1197);
and U1368 (N_1368,N_1151,N_1120);
or U1369 (N_1369,N_1158,N_1168);
and U1370 (N_1370,N_1106,N_1092);
nor U1371 (N_1371,N_1054,N_1198);
nor U1372 (N_1372,N_1091,N_1148);
nand U1373 (N_1373,N_1028,N_1147);
and U1374 (N_1374,N_1035,N_1025);
or U1375 (N_1375,N_1116,N_1021);
nand U1376 (N_1376,N_1009,N_1037);
nor U1377 (N_1377,N_1171,N_1135);
or U1378 (N_1378,N_1049,N_1143);
nand U1379 (N_1379,N_1053,N_1114);
xnor U1380 (N_1380,N_1008,N_1087);
nand U1381 (N_1381,N_1062,N_1046);
and U1382 (N_1382,N_1120,N_1075);
and U1383 (N_1383,N_1129,N_1111);
and U1384 (N_1384,N_1003,N_1111);
xnor U1385 (N_1385,N_1164,N_1160);
xor U1386 (N_1386,N_1044,N_1041);
nand U1387 (N_1387,N_1174,N_1114);
xnor U1388 (N_1388,N_1141,N_1075);
nor U1389 (N_1389,N_1086,N_1052);
and U1390 (N_1390,N_1051,N_1003);
nand U1391 (N_1391,N_1188,N_1190);
or U1392 (N_1392,N_1162,N_1179);
or U1393 (N_1393,N_1110,N_1195);
nor U1394 (N_1394,N_1058,N_1049);
nand U1395 (N_1395,N_1124,N_1062);
xor U1396 (N_1396,N_1198,N_1183);
or U1397 (N_1397,N_1069,N_1095);
nor U1398 (N_1398,N_1034,N_1137);
or U1399 (N_1399,N_1048,N_1034);
xor U1400 (N_1400,N_1387,N_1353);
or U1401 (N_1401,N_1269,N_1334);
nor U1402 (N_1402,N_1378,N_1379);
nor U1403 (N_1403,N_1284,N_1226);
xnor U1404 (N_1404,N_1258,N_1254);
nor U1405 (N_1405,N_1365,N_1299);
or U1406 (N_1406,N_1246,N_1320);
or U1407 (N_1407,N_1229,N_1352);
nor U1408 (N_1408,N_1202,N_1380);
nand U1409 (N_1409,N_1339,N_1250);
or U1410 (N_1410,N_1338,N_1244);
nor U1411 (N_1411,N_1203,N_1393);
or U1412 (N_1412,N_1376,N_1396);
nor U1413 (N_1413,N_1359,N_1397);
nand U1414 (N_1414,N_1364,N_1219);
nand U1415 (N_1415,N_1314,N_1275);
nand U1416 (N_1416,N_1372,N_1337);
or U1417 (N_1417,N_1363,N_1375);
nor U1418 (N_1418,N_1325,N_1398);
nor U1419 (N_1419,N_1266,N_1362);
nand U1420 (N_1420,N_1298,N_1259);
and U1421 (N_1421,N_1241,N_1368);
and U1422 (N_1422,N_1350,N_1377);
nand U1423 (N_1423,N_1370,N_1255);
and U1424 (N_1424,N_1309,N_1336);
nor U1425 (N_1425,N_1331,N_1205);
and U1426 (N_1426,N_1208,N_1392);
nor U1427 (N_1427,N_1347,N_1311);
and U1428 (N_1428,N_1213,N_1328);
xnor U1429 (N_1429,N_1218,N_1214);
nor U1430 (N_1430,N_1300,N_1210);
xnor U1431 (N_1431,N_1312,N_1280);
and U1432 (N_1432,N_1341,N_1316);
and U1433 (N_1433,N_1285,N_1253);
nand U1434 (N_1434,N_1354,N_1342);
or U1435 (N_1435,N_1355,N_1340);
or U1436 (N_1436,N_1228,N_1322);
nand U1437 (N_1437,N_1324,N_1289);
or U1438 (N_1438,N_1385,N_1366);
and U1439 (N_1439,N_1291,N_1274);
and U1440 (N_1440,N_1286,N_1315);
nor U1441 (N_1441,N_1234,N_1327);
or U1442 (N_1442,N_1209,N_1252);
and U1443 (N_1443,N_1304,N_1318);
nor U1444 (N_1444,N_1360,N_1297);
and U1445 (N_1445,N_1367,N_1344);
xor U1446 (N_1446,N_1233,N_1351);
nor U1447 (N_1447,N_1222,N_1382);
xor U1448 (N_1448,N_1217,N_1313);
nor U1449 (N_1449,N_1270,N_1288);
nor U1450 (N_1450,N_1293,N_1395);
and U1451 (N_1451,N_1374,N_1201);
nand U1452 (N_1452,N_1358,N_1207);
xor U1453 (N_1453,N_1333,N_1277);
xor U1454 (N_1454,N_1295,N_1278);
xor U1455 (N_1455,N_1216,N_1230);
and U1456 (N_1456,N_1242,N_1349);
or U1457 (N_1457,N_1256,N_1317);
nand U1458 (N_1458,N_1357,N_1319);
and U1459 (N_1459,N_1248,N_1373);
nand U1460 (N_1460,N_1330,N_1238);
nor U1461 (N_1461,N_1292,N_1281);
and U1462 (N_1462,N_1206,N_1394);
and U1463 (N_1463,N_1240,N_1329);
nand U1464 (N_1464,N_1239,N_1389);
or U1465 (N_1465,N_1303,N_1287);
or U1466 (N_1466,N_1399,N_1371);
nor U1467 (N_1467,N_1227,N_1290);
nor U1468 (N_1468,N_1391,N_1243);
and U1469 (N_1469,N_1326,N_1261);
or U1470 (N_1470,N_1265,N_1308);
and U1471 (N_1471,N_1271,N_1388);
and U1472 (N_1472,N_1305,N_1346);
xor U1473 (N_1473,N_1231,N_1310);
and U1474 (N_1474,N_1267,N_1225);
nand U1475 (N_1475,N_1200,N_1302);
nor U1476 (N_1476,N_1247,N_1361);
and U1477 (N_1477,N_1381,N_1212);
or U1478 (N_1478,N_1235,N_1369);
nor U1479 (N_1479,N_1276,N_1321);
or U1480 (N_1480,N_1223,N_1383);
nor U1481 (N_1481,N_1272,N_1263);
xor U1482 (N_1482,N_1294,N_1356);
or U1483 (N_1483,N_1264,N_1215);
nor U1484 (N_1484,N_1332,N_1282);
nand U1485 (N_1485,N_1296,N_1262);
nand U1486 (N_1486,N_1224,N_1306);
nor U1487 (N_1487,N_1301,N_1257);
xor U1488 (N_1488,N_1260,N_1323);
nand U1489 (N_1489,N_1204,N_1221);
or U1490 (N_1490,N_1268,N_1232);
and U1491 (N_1491,N_1249,N_1220);
or U1492 (N_1492,N_1390,N_1307);
nor U1493 (N_1493,N_1335,N_1245);
nand U1494 (N_1494,N_1348,N_1211);
nor U1495 (N_1495,N_1345,N_1343);
or U1496 (N_1496,N_1386,N_1236);
or U1497 (N_1497,N_1251,N_1279);
nor U1498 (N_1498,N_1273,N_1283);
nor U1499 (N_1499,N_1384,N_1237);
and U1500 (N_1500,N_1271,N_1389);
or U1501 (N_1501,N_1248,N_1276);
nand U1502 (N_1502,N_1239,N_1257);
nand U1503 (N_1503,N_1370,N_1382);
nor U1504 (N_1504,N_1341,N_1333);
xor U1505 (N_1505,N_1330,N_1363);
xor U1506 (N_1506,N_1327,N_1257);
and U1507 (N_1507,N_1345,N_1270);
nand U1508 (N_1508,N_1323,N_1317);
and U1509 (N_1509,N_1378,N_1242);
and U1510 (N_1510,N_1349,N_1389);
nand U1511 (N_1511,N_1344,N_1312);
xor U1512 (N_1512,N_1218,N_1339);
or U1513 (N_1513,N_1332,N_1389);
nor U1514 (N_1514,N_1353,N_1230);
xor U1515 (N_1515,N_1215,N_1345);
xnor U1516 (N_1516,N_1292,N_1245);
nor U1517 (N_1517,N_1354,N_1361);
and U1518 (N_1518,N_1278,N_1391);
and U1519 (N_1519,N_1292,N_1324);
or U1520 (N_1520,N_1384,N_1229);
nor U1521 (N_1521,N_1348,N_1327);
and U1522 (N_1522,N_1231,N_1304);
and U1523 (N_1523,N_1395,N_1343);
nor U1524 (N_1524,N_1360,N_1263);
nor U1525 (N_1525,N_1227,N_1235);
or U1526 (N_1526,N_1266,N_1396);
nand U1527 (N_1527,N_1390,N_1320);
nor U1528 (N_1528,N_1213,N_1289);
and U1529 (N_1529,N_1365,N_1203);
nor U1530 (N_1530,N_1370,N_1332);
or U1531 (N_1531,N_1333,N_1203);
xnor U1532 (N_1532,N_1202,N_1374);
nand U1533 (N_1533,N_1330,N_1381);
or U1534 (N_1534,N_1266,N_1258);
nand U1535 (N_1535,N_1280,N_1286);
nor U1536 (N_1536,N_1369,N_1264);
nor U1537 (N_1537,N_1242,N_1295);
and U1538 (N_1538,N_1354,N_1311);
nand U1539 (N_1539,N_1369,N_1284);
nor U1540 (N_1540,N_1334,N_1267);
nor U1541 (N_1541,N_1319,N_1356);
nor U1542 (N_1542,N_1372,N_1207);
nand U1543 (N_1543,N_1254,N_1375);
and U1544 (N_1544,N_1211,N_1327);
nor U1545 (N_1545,N_1349,N_1365);
nor U1546 (N_1546,N_1295,N_1356);
nor U1547 (N_1547,N_1209,N_1290);
nor U1548 (N_1548,N_1327,N_1201);
and U1549 (N_1549,N_1305,N_1355);
nand U1550 (N_1550,N_1281,N_1383);
or U1551 (N_1551,N_1373,N_1224);
or U1552 (N_1552,N_1232,N_1257);
or U1553 (N_1553,N_1260,N_1395);
and U1554 (N_1554,N_1347,N_1227);
and U1555 (N_1555,N_1235,N_1217);
or U1556 (N_1556,N_1272,N_1357);
or U1557 (N_1557,N_1288,N_1351);
nand U1558 (N_1558,N_1323,N_1244);
nand U1559 (N_1559,N_1249,N_1299);
and U1560 (N_1560,N_1242,N_1320);
and U1561 (N_1561,N_1325,N_1255);
or U1562 (N_1562,N_1228,N_1272);
and U1563 (N_1563,N_1396,N_1243);
nand U1564 (N_1564,N_1200,N_1271);
and U1565 (N_1565,N_1283,N_1229);
and U1566 (N_1566,N_1249,N_1359);
or U1567 (N_1567,N_1394,N_1273);
or U1568 (N_1568,N_1208,N_1203);
nand U1569 (N_1569,N_1236,N_1362);
nand U1570 (N_1570,N_1347,N_1339);
nor U1571 (N_1571,N_1243,N_1393);
or U1572 (N_1572,N_1397,N_1252);
and U1573 (N_1573,N_1329,N_1297);
nor U1574 (N_1574,N_1227,N_1319);
nand U1575 (N_1575,N_1367,N_1314);
nor U1576 (N_1576,N_1389,N_1329);
nand U1577 (N_1577,N_1396,N_1279);
or U1578 (N_1578,N_1264,N_1297);
or U1579 (N_1579,N_1251,N_1315);
and U1580 (N_1580,N_1382,N_1272);
nor U1581 (N_1581,N_1355,N_1227);
nor U1582 (N_1582,N_1288,N_1349);
nor U1583 (N_1583,N_1350,N_1398);
or U1584 (N_1584,N_1377,N_1323);
nand U1585 (N_1585,N_1372,N_1302);
or U1586 (N_1586,N_1340,N_1258);
nor U1587 (N_1587,N_1269,N_1242);
and U1588 (N_1588,N_1207,N_1318);
or U1589 (N_1589,N_1385,N_1301);
xnor U1590 (N_1590,N_1208,N_1233);
nor U1591 (N_1591,N_1233,N_1248);
nand U1592 (N_1592,N_1357,N_1380);
nor U1593 (N_1593,N_1205,N_1271);
nand U1594 (N_1594,N_1393,N_1213);
nor U1595 (N_1595,N_1213,N_1269);
or U1596 (N_1596,N_1334,N_1264);
nor U1597 (N_1597,N_1214,N_1335);
xor U1598 (N_1598,N_1206,N_1244);
or U1599 (N_1599,N_1232,N_1370);
nor U1600 (N_1600,N_1594,N_1478);
or U1601 (N_1601,N_1510,N_1447);
nand U1602 (N_1602,N_1458,N_1502);
and U1603 (N_1603,N_1523,N_1487);
or U1604 (N_1604,N_1521,N_1583);
nand U1605 (N_1605,N_1443,N_1446);
nand U1606 (N_1606,N_1406,N_1522);
and U1607 (N_1607,N_1575,N_1412);
or U1608 (N_1608,N_1483,N_1552);
and U1609 (N_1609,N_1568,N_1449);
and U1610 (N_1610,N_1426,N_1545);
and U1611 (N_1611,N_1414,N_1560);
or U1612 (N_1612,N_1481,N_1581);
nor U1613 (N_1613,N_1513,N_1531);
or U1614 (N_1614,N_1507,N_1473);
nor U1615 (N_1615,N_1579,N_1496);
and U1616 (N_1616,N_1511,N_1469);
or U1617 (N_1617,N_1440,N_1535);
and U1618 (N_1618,N_1453,N_1546);
nor U1619 (N_1619,N_1571,N_1516);
or U1620 (N_1620,N_1574,N_1548);
nor U1621 (N_1621,N_1459,N_1526);
nand U1622 (N_1622,N_1567,N_1556);
nor U1623 (N_1623,N_1451,N_1479);
nor U1624 (N_1624,N_1514,N_1464);
nand U1625 (N_1625,N_1561,N_1551);
or U1626 (N_1626,N_1517,N_1512);
nor U1627 (N_1627,N_1518,N_1407);
nand U1628 (N_1628,N_1591,N_1566);
nor U1629 (N_1629,N_1505,N_1537);
nor U1630 (N_1630,N_1562,N_1588);
xnor U1631 (N_1631,N_1599,N_1405);
nand U1632 (N_1632,N_1422,N_1540);
xnor U1633 (N_1633,N_1532,N_1555);
or U1634 (N_1634,N_1554,N_1564);
or U1635 (N_1635,N_1442,N_1477);
nand U1636 (N_1636,N_1475,N_1441);
nor U1637 (N_1637,N_1509,N_1499);
nor U1638 (N_1638,N_1500,N_1553);
nand U1639 (N_1639,N_1428,N_1456);
nand U1640 (N_1640,N_1462,N_1404);
or U1641 (N_1641,N_1525,N_1429);
nand U1642 (N_1642,N_1558,N_1519);
or U1643 (N_1643,N_1547,N_1401);
nor U1644 (N_1644,N_1520,N_1416);
nor U1645 (N_1645,N_1578,N_1582);
nor U1646 (N_1646,N_1435,N_1415);
or U1647 (N_1647,N_1542,N_1413);
or U1648 (N_1648,N_1592,N_1536);
nor U1649 (N_1649,N_1445,N_1431);
nor U1650 (N_1650,N_1497,N_1533);
nor U1651 (N_1651,N_1529,N_1570);
nor U1652 (N_1652,N_1589,N_1572);
nand U1653 (N_1653,N_1494,N_1490);
or U1654 (N_1654,N_1489,N_1596);
nor U1655 (N_1655,N_1400,N_1504);
nand U1656 (N_1656,N_1450,N_1515);
or U1657 (N_1657,N_1438,N_1538);
and U1658 (N_1658,N_1425,N_1543);
and U1659 (N_1659,N_1430,N_1408);
or U1660 (N_1660,N_1576,N_1423);
xor U1661 (N_1661,N_1508,N_1409);
xnor U1662 (N_1662,N_1433,N_1539);
nor U1663 (N_1663,N_1584,N_1468);
nand U1664 (N_1664,N_1486,N_1418);
or U1665 (N_1665,N_1439,N_1455);
nor U1666 (N_1666,N_1492,N_1527);
xor U1667 (N_1667,N_1586,N_1587);
nand U1668 (N_1668,N_1573,N_1569);
nand U1669 (N_1669,N_1503,N_1463);
xnor U1670 (N_1670,N_1528,N_1436);
or U1671 (N_1671,N_1488,N_1454);
and U1672 (N_1672,N_1472,N_1437);
or U1673 (N_1673,N_1530,N_1544);
or U1674 (N_1674,N_1421,N_1590);
nand U1675 (N_1675,N_1466,N_1585);
and U1676 (N_1676,N_1403,N_1467);
nand U1677 (N_1677,N_1460,N_1550);
nor U1678 (N_1678,N_1595,N_1534);
nor U1679 (N_1679,N_1541,N_1549);
and U1680 (N_1680,N_1597,N_1501);
or U1681 (N_1681,N_1471,N_1557);
and U1682 (N_1682,N_1444,N_1524);
or U1683 (N_1683,N_1465,N_1434);
nor U1684 (N_1684,N_1495,N_1411);
xnor U1685 (N_1685,N_1506,N_1420);
and U1686 (N_1686,N_1498,N_1559);
nor U1687 (N_1687,N_1457,N_1593);
and U1688 (N_1688,N_1577,N_1493);
nor U1689 (N_1689,N_1474,N_1432);
nor U1690 (N_1690,N_1461,N_1419);
nand U1691 (N_1691,N_1598,N_1484);
nor U1692 (N_1692,N_1402,N_1491);
nand U1693 (N_1693,N_1480,N_1563);
and U1694 (N_1694,N_1410,N_1565);
nor U1695 (N_1695,N_1482,N_1485);
and U1696 (N_1696,N_1427,N_1476);
and U1697 (N_1697,N_1452,N_1470);
nor U1698 (N_1698,N_1580,N_1448);
and U1699 (N_1699,N_1424,N_1417);
nand U1700 (N_1700,N_1446,N_1463);
or U1701 (N_1701,N_1436,N_1559);
and U1702 (N_1702,N_1445,N_1403);
and U1703 (N_1703,N_1579,N_1468);
nand U1704 (N_1704,N_1470,N_1565);
xnor U1705 (N_1705,N_1461,N_1505);
xnor U1706 (N_1706,N_1599,N_1425);
nand U1707 (N_1707,N_1448,N_1487);
nand U1708 (N_1708,N_1513,N_1444);
nand U1709 (N_1709,N_1560,N_1402);
or U1710 (N_1710,N_1415,N_1500);
xnor U1711 (N_1711,N_1486,N_1400);
or U1712 (N_1712,N_1446,N_1554);
or U1713 (N_1713,N_1541,N_1511);
nor U1714 (N_1714,N_1498,N_1535);
nor U1715 (N_1715,N_1470,N_1484);
or U1716 (N_1716,N_1500,N_1530);
and U1717 (N_1717,N_1407,N_1553);
or U1718 (N_1718,N_1533,N_1426);
and U1719 (N_1719,N_1486,N_1501);
or U1720 (N_1720,N_1589,N_1474);
or U1721 (N_1721,N_1547,N_1427);
and U1722 (N_1722,N_1572,N_1435);
xnor U1723 (N_1723,N_1557,N_1480);
xnor U1724 (N_1724,N_1563,N_1407);
nor U1725 (N_1725,N_1471,N_1488);
nor U1726 (N_1726,N_1501,N_1490);
and U1727 (N_1727,N_1406,N_1491);
and U1728 (N_1728,N_1579,N_1409);
or U1729 (N_1729,N_1541,N_1571);
or U1730 (N_1730,N_1473,N_1597);
or U1731 (N_1731,N_1475,N_1415);
nor U1732 (N_1732,N_1539,N_1597);
or U1733 (N_1733,N_1544,N_1562);
nor U1734 (N_1734,N_1557,N_1546);
xor U1735 (N_1735,N_1528,N_1578);
or U1736 (N_1736,N_1495,N_1450);
and U1737 (N_1737,N_1432,N_1505);
nand U1738 (N_1738,N_1486,N_1422);
nand U1739 (N_1739,N_1515,N_1581);
and U1740 (N_1740,N_1519,N_1449);
nand U1741 (N_1741,N_1497,N_1550);
nor U1742 (N_1742,N_1488,N_1407);
and U1743 (N_1743,N_1456,N_1417);
and U1744 (N_1744,N_1423,N_1506);
or U1745 (N_1745,N_1509,N_1482);
or U1746 (N_1746,N_1404,N_1523);
xnor U1747 (N_1747,N_1513,N_1489);
nand U1748 (N_1748,N_1412,N_1516);
and U1749 (N_1749,N_1579,N_1472);
nand U1750 (N_1750,N_1529,N_1539);
nor U1751 (N_1751,N_1536,N_1503);
or U1752 (N_1752,N_1431,N_1543);
nor U1753 (N_1753,N_1571,N_1584);
or U1754 (N_1754,N_1427,N_1508);
nor U1755 (N_1755,N_1447,N_1432);
and U1756 (N_1756,N_1408,N_1521);
and U1757 (N_1757,N_1537,N_1534);
nor U1758 (N_1758,N_1407,N_1538);
nand U1759 (N_1759,N_1498,N_1432);
nand U1760 (N_1760,N_1565,N_1525);
or U1761 (N_1761,N_1456,N_1410);
and U1762 (N_1762,N_1428,N_1546);
or U1763 (N_1763,N_1414,N_1407);
nand U1764 (N_1764,N_1513,N_1567);
nand U1765 (N_1765,N_1490,N_1447);
nor U1766 (N_1766,N_1541,N_1578);
xor U1767 (N_1767,N_1582,N_1556);
or U1768 (N_1768,N_1568,N_1439);
nor U1769 (N_1769,N_1429,N_1506);
and U1770 (N_1770,N_1426,N_1586);
or U1771 (N_1771,N_1488,N_1506);
xnor U1772 (N_1772,N_1536,N_1533);
xnor U1773 (N_1773,N_1425,N_1477);
nand U1774 (N_1774,N_1481,N_1539);
or U1775 (N_1775,N_1528,N_1475);
nor U1776 (N_1776,N_1450,N_1594);
xor U1777 (N_1777,N_1529,N_1443);
nor U1778 (N_1778,N_1573,N_1497);
nand U1779 (N_1779,N_1490,N_1561);
or U1780 (N_1780,N_1432,N_1537);
or U1781 (N_1781,N_1455,N_1555);
and U1782 (N_1782,N_1447,N_1401);
nand U1783 (N_1783,N_1438,N_1419);
xnor U1784 (N_1784,N_1550,N_1462);
or U1785 (N_1785,N_1578,N_1418);
nand U1786 (N_1786,N_1501,N_1509);
and U1787 (N_1787,N_1428,N_1413);
or U1788 (N_1788,N_1520,N_1597);
and U1789 (N_1789,N_1466,N_1521);
and U1790 (N_1790,N_1555,N_1559);
and U1791 (N_1791,N_1584,N_1540);
nor U1792 (N_1792,N_1457,N_1444);
and U1793 (N_1793,N_1491,N_1479);
or U1794 (N_1794,N_1401,N_1546);
nand U1795 (N_1795,N_1547,N_1556);
nor U1796 (N_1796,N_1483,N_1410);
nand U1797 (N_1797,N_1415,N_1539);
nand U1798 (N_1798,N_1472,N_1490);
or U1799 (N_1799,N_1525,N_1522);
or U1800 (N_1800,N_1622,N_1670);
or U1801 (N_1801,N_1693,N_1745);
xnor U1802 (N_1802,N_1718,N_1797);
and U1803 (N_1803,N_1686,N_1650);
and U1804 (N_1804,N_1777,N_1760);
and U1805 (N_1805,N_1669,N_1655);
and U1806 (N_1806,N_1742,N_1625);
and U1807 (N_1807,N_1762,N_1657);
and U1808 (N_1808,N_1784,N_1783);
or U1809 (N_1809,N_1609,N_1756);
and U1810 (N_1810,N_1631,N_1724);
or U1811 (N_1811,N_1601,N_1647);
nor U1812 (N_1812,N_1730,N_1785);
xnor U1813 (N_1813,N_1606,N_1674);
nor U1814 (N_1814,N_1640,N_1721);
nor U1815 (N_1815,N_1645,N_1773);
xor U1816 (N_1816,N_1734,N_1683);
and U1817 (N_1817,N_1626,N_1659);
and U1818 (N_1818,N_1664,N_1776);
nor U1819 (N_1819,N_1779,N_1608);
nor U1820 (N_1820,N_1795,N_1714);
xor U1821 (N_1821,N_1663,N_1692);
and U1822 (N_1822,N_1727,N_1765);
nor U1823 (N_1823,N_1636,N_1600);
nand U1824 (N_1824,N_1619,N_1675);
and U1825 (N_1825,N_1708,N_1649);
or U1826 (N_1826,N_1603,N_1732);
xnor U1827 (N_1827,N_1757,N_1658);
nor U1828 (N_1828,N_1768,N_1746);
nor U1829 (N_1829,N_1627,N_1710);
nor U1830 (N_1830,N_1702,N_1643);
and U1831 (N_1831,N_1728,N_1614);
xnor U1832 (N_1832,N_1688,N_1672);
nand U1833 (N_1833,N_1755,N_1753);
nor U1834 (N_1834,N_1646,N_1653);
nand U1835 (N_1835,N_1705,N_1689);
nand U1836 (N_1836,N_1729,N_1671);
xnor U1837 (N_1837,N_1690,N_1673);
nand U1838 (N_1838,N_1759,N_1662);
and U1839 (N_1839,N_1763,N_1656);
xnor U1840 (N_1840,N_1723,N_1667);
or U1841 (N_1841,N_1788,N_1610);
xnor U1842 (N_1842,N_1665,N_1612);
nand U1843 (N_1843,N_1633,N_1735);
nand U1844 (N_1844,N_1651,N_1694);
nor U1845 (N_1845,N_1703,N_1677);
xnor U1846 (N_1846,N_1774,N_1680);
and U1847 (N_1847,N_1628,N_1717);
and U1848 (N_1848,N_1722,N_1715);
or U1849 (N_1849,N_1676,N_1638);
and U1850 (N_1850,N_1615,N_1654);
nand U1851 (N_1851,N_1701,N_1790);
and U1852 (N_1852,N_1697,N_1605);
and U1853 (N_1853,N_1660,N_1704);
nor U1854 (N_1854,N_1764,N_1696);
or U1855 (N_1855,N_1624,N_1700);
nor U1856 (N_1856,N_1639,N_1652);
nand U1857 (N_1857,N_1743,N_1618);
or U1858 (N_1858,N_1720,N_1648);
xnor U1859 (N_1859,N_1786,N_1634);
or U1860 (N_1860,N_1684,N_1716);
nor U1861 (N_1861,N_1616,N_1678);
nand U1862 (N_1862,N_1719,N_1713);
and U1863 (N_1863,N_1733,N_1613);
xor U1864 (N_1864,N_1731,N_1699);
and U1865 (N_1865,N_1794,N_1787);
or U1866 (N_1866,N_1738,N_1754);
and U1867 (N_1867,N_1630,N_1750);
nor U1868 (N_1868,N_1796,N_1668);
xor U1869 (N_1869,N_1681,N_1725);
and U1870 (N_1870,N_1749,N_1644);
nand U1871 (N_1871,N_1637,N_1798);
nand U1872 (N_1872,N_1792,N_1778);
and U1873 (N_1873,N_1747,N_1770);
and U1874 (N_1874,N_1642,N_1739);
or U1875 (N_1875,N_1736,N_1629);
or U1876 (N_1876,N_1691,N_1741);
xnor U1877 (N_1877,N_1782,N_1771);
nand U1878 (N_1878,N_1769,N_1698);
and U1879 (N_1879,N_1758,N_1635);
nor U1880 (N_1880,N_1611,N_1602);
and U1881 (N_1881,N_1789,N_1682);
nor U1882 (N_1882,N_1641,N_1661);
or U1883 (N_1883,N_1766,N_1748);
nand U1884 (N_1884,N_1617,N_1711);
or U1885 (N_1885,N_1666,N_1767);
nor U1886 (N_1886,N_1623,N_1621);
nor U1887 (N_1887,N_1632,N_1709);
and U1888 (N_1888,N_1780,N_1607);
nand U1889 (N_1889,N_1687,N_1775);
xnor U1890 (N_1890,N_1737,N_1712);
or U1891 (N_1891,N_1752,N_1761);
and U1892 (N_1892,N_1604,N_1679);
and U1893 (N_1893,N_1740,N_1726);
or U1894 (N_1894,N_1772,N_1799);
nor U1895 (N_1895,N_1744,N_1707);
nand U1896 (N_1896,N_1791,N_1695);
or U1897 (N_1897,N_1620,N_1751);
and U1898 (N_1898,N_1706,N_1685);
and U1899 (N_1899,N_1793,N_1781);
nor U1900 (N_1900,N_1779,N_1760);
and U1901 (N_1901,N_1673,N_1790);
nor U1902 (N_1902,N_1794,N_1693);
or U1903 (N_1903,N_1674,N_1720);
nor U1904 (N_1904,N_1779,N_1748);
or U1905 (N_1905,N_1691,N_1780);
nor U1906 (N_1906,N_1649,N_1779);
xnor U1907 (N_1907,N_1678,N_1658);
nand U1908 (N_1908,N_1691,N_1602);
and U1909 (N_1909,N_1645,N_1634);
and U1910 (N_1910,N_1714,N_1650);
and U1911 (N_1911,N_1772,N_1689);
nand U1912 (N_1912,N_1788,N_1707);
and U1913 (N_1913,N_1787,N_1662);
nand U1914 (N_1914,N_1632,N_1740);
nand U1915 (N_1915,N_1637,N_1642);
and U1916 (N_1916,N_1729,N_1691);
and U1917 (N_1917,N_1608,N_1775);
and U1918 (N_1918,N_1726,N_1716);
xnor U1919 (N_1919,N_1600,N_1696);
nor U1920 (N_1920,N_1686,N_1632);
or U1921 (N_1921,N_1667,N_1774);
or U1922 (N_1922,N_1629,N_1772);
and U1923 (N_1923,N_1617,N_1758);
or U1924 (N_1924,N_1701,N_1783);
or U1925 (N_1925,N_1689,N_1793);
and U1926 (N_1926,N_1701,N_1799);
nand U1927 (N_1927,N_1712,N_1603);
nand U1928 (N_1928,N_1677,N_1612);
nor U1929 (N_1929,N_1606,N_1671);
and U1930 (N_1930,N_1638,N_1692);
and U1931 (N_1931,N_1648,N_1674);
and U1932 (N_1932,N_1785,N_1796);
nand U1933 (N_1933,N_1623,N_1760);
or U1934 (N_1934,N_1775,N_1780);
or U1935 (N_1935,N_1683,N_1673);
xnor U1936 (N_1936,N_1652,N_1680);
nand U1937 (N_1937,N_1717,N_1785);
nand U1938 (N_1938,N_1755,N_1757);
or U1939 (N_1939,N_1617,N_1788);
or U1940 (N_1940,N_1749,N_1726);
and U1941 (N_1941,N_1717,N_1687);
nand U1942 (N_1942,N_1792,N_1654);
and U1943 (N_1943,N_1715,N_1604);
or U1944 (N_1944,N_1712,N_1689);
and U1945 (N_1945,N_1634,N_1688);
and U1946 (N_1946,N_1641,N_1718);
nand U1947 (N_1947,N_1632,N_1783);
or U1948 (N_1948,N_1649,N_1606);
nor U1949 (N_1949,N_1777,N_1678);
or U1950 (N_1950,N_1769,N_1678);
nor U1951 (N_1951,N_1719,N_1644);
nand U1952 (N_1952,N_1643,N_1764);
nand U1953 (N_1953,N_1755,N_1718);
nand U1954 (N_1954,N_1618,N_1752);
nor U1955 (N_1955,N_1612,N_1642);
nand U1956 (N_1956,N_1657,N_1723);
nand U1957 (N_1957,N_1624,N_1622);
xnor U1958 (N_1958,N_1684,N_1718);
nand U1959 (N_1959,N_1636,N_1682);
xor U1960 (N_1960,N_1654,N_1683);
nand U1961 (N_1961,N_1642,N_1789);
nand U1962 (N_1962,N_1748,N_1621);
and U1963 (N_1963,N_1796,N_1645);
or U1964 (N_1964,N_1795,N_1786);
nor U1965 (N_1965,N_1629,N_1769);
nor U1966 (N_1966,N_1738,N_1631);
nor U1967 (N_1967,N_1616,N_1762);
xnor U1968 (N_1968,N_1795,N_1667);
nand U1969 (N_1969,N_1631,N_1679);
or U1970 (N_1970,N_1749,N_1663);
and U1971 (N_1971,N_1657,N_1769);
or U1972 (N_1972,N_1645,N_1603);
nor U1973 (N_1973,N_1754,N_1676);
xor U1974 (N_1974,N_1670,N_1794);
nand U1975 (N_1975,N_1773,N_1721);
and U1976 (N_1976,N_1686,N_1670);
nor U1977 (N_1977,N_1728,N_1766);
nor U1978 (N_1978,N_1772,N_1665);
nand U1979 (N_1979,N_1636,N_1648);
or U1980 (N_1980,N_1717,N_1732);
and U1981 (N_1981,N_1601,N_1700);
nand U1982 (N_1982,N_1742,N_1794);
nand U1983 (N_1983,N_1707,N_1755);
nand U1984 (N_1984,N_1738,N_1799);
xor U1985 (N_1985,N_1728,N_1781);
nor U1986 (N_1986,N_1630,N_1703);
nor U1987 (N_1987,N_1681,N_1784);
nor U1988 (N_1988,N_1652,N_1722);
nor U1989 (N_1989,N_1736,N_1745);
nor U1990 (N_1990,N_1719,N_1738);
nand U1991 (N_1991,N_1662,N_1655);
and U1992 (N_1992,N_1652,N_1736);
nor U1993 (N_1993,N_1790,N_1716);
nor U1994 (N_1994,N_1716,N_1606);
nor U1995 (N_1995,N_1642,N_1657);
xnor U1996 (N_1996,N_1652,N_1693);
nand U1997 (N_1997,N_1666,N_1777);
or U1998 (N_1998,N_1648,N_1612);
nor U1999 (N_1999,N_1603,N_1796);
or U2000 (N_2000,N_1948,N_1996);
nand U2001 (N_2001,N_1983,N_1963);
nand U2002 (N_2002,N_1962,N_1871);
or U2003 (N_2003,N_1997,N_1842);
or U2004 (N_2004,N_1800,N_1937);
and U2005 (N_2005,N_1801,N_1979);
and U2006 (N_2006,N_1931,N_1816);
and U2007 (N_2007,N_1815,N_1953);
nor U2008 (N_2008,N_1855,N_1819);
or U2009 (N_2009,N_1820,N_1827);
or U2010 (N_2010,N_1951,N_1877);
or U2011 (N_2011,N_1803,N_1821);
and U2012 (N_2012,N_1884,N_1843);
nor U2013 (N_2013,N_1844,N_1859);
nor U2014 (N_2014,N_1916,N_1930);
xnor U2015 (N_2015,N_1894,N_1955);
and U2016 (N_2016,N_1829,N_1926);
nand U2017 (N_2017,N_1857,N_1991);
nand U2018 (N_2018,N_1874,N_1840);
xor U2019 (N_2019,N_1880,N_1858);
nor U2020 (N_2020,N_1920,N_1908);
nand U2021 (N_2021,N_1835,N_1947);
xor U2022 (N_2022,N_1917,N_1866);
or U2023 (N_2023,N_1836,N_1861);
or U2024 (N_2024,N_1817,N_1952);
and U2025 (N_2025,N_1883,N_1886);
or U2026 (N_2026,N_1887,N_1988);
nand U2027 (N_2027,N_1911,N_1933);
xor U2028 (N_2028,N_1964,N_1847);
nor U2029 (N_2029,N_1878,N_1851);
or U2030 (N_2030,N_1876,N_1961);
and U2031 (N_2031,N_1976,N_1927);
and U2032 (N_2032,N_1804,N_1949);
or U2033 (N_2033,N_1832,N_1995);
or U2034 (N_2034,N_1982,N_1823);
nand U2035 (N_2035,N_1939,N_1833);
and U2036 (N_2036,N_1856,N_1872);
nor U2037 (N_2037,N_1936,N_1891);
or U2038 (N_2038,N_1923,N_1987);
nor U2039 (N_2039,N_1919,N_1918);
nand U2040 (N_2040,N_1958,N_1989);
nand U2041 (N_2041,N_1966,N_1845);
nand U2042 (N_2042,N_1882,N_1849);
and U2043 (N_2043,N_1914,N_1915);
or U2044 (N_2044,N_1890,N_1910);
and U2045 (N_2045,N_1826,N_1814);
and U2046 (N_2046,N_1852,N_1959);
nor U2047 (N_2047,N_1934,N_1909);
or U2048 (N_2048,N_1975,N_1970);
nand U2049 (N_2049,N_1839,N_1869);
or U2050 (N_2050,N_1831,N_1881);
and U2051 (N_2051,N_1813,N_1932);
or U2052 (N_2052,N_1818,N_1942);
nand U2053 (N_2053,N_1863,N_1985);
or U2054 (N_2054,N_1913,N_1848);
or U2055 (N_2055,N_1875,N_1957);
nand U2056 (N_2056,N_1921,N_1899);
or U2057 (N_2057,N_1853,N_1954);
and U2058 (N_2058,N_1850,N_1806);
or U2059 (N_2059,N_1834,N_1967);
and U2060 (N_2060,N_1888,N_1893);
and U2061 (N_2061,N_1809,N_1925);
nand U2062 (N_2062,N_1946,N_1825);
and U2063 (N_2063,N_1971,N_1973);
and U2064 (N_2064,N_1960,N_1895);
nand U2065 (N_2065,N_1912,N_1867);
nor U2066 (N_2066,N_1854,N_1900);
or U2067 (N_2067,N_1965,N_1993);
xor U2068 (N_2068,N_1873,N_1922);
and U2069 (N_2069,N_1992,N_1838);
and U2070 (N_2070,N_1812,N_1811);
xnor U2071 (N_2071,N_1805,N_1846);
and U2072 (N_2072,N_1984,N_1892);
or U2073 (N_2073,N_1897,N_1864);
nor U2074 (N_2074,N_1904,N_1860);
xor U2075 (N_2075,N_1924,N_1885);
xor U2076 (N_2076,N_1907,N_1901);
nand U2077 (N_2077,N_1862,N_1974);
nor U2078 (N_2078,N_1990,N_1981);
or U2079 (N_2079,N_1868,N_1994);
and U2080 (N_2080,N_1808,N_1906);
and U2081 (N_2081,N_1810,N_1879);
and U2082 (N_2082,N_1807,N_1828);
or U2083 (N_2083,N_1940,N_1950);
or U2084 (N_2084,N_1802,N_1941);
nor U2085 (N_2085,N_1889,N_1977);
xnor U2086 (N_2086,N_1830,N_1956);
nor U2087 (N_2087,N_1865,N_1824);
and U2088 (N_2088,N_1896,N_1986);
or U2089 (N_2089,N_1945,N_1944);
or U2090 (N_2090,N_1870,N_1980);
and U2091 (N_2091,N_1902,N_1938);
and U2092 (N_2092,N_1998,N_1999);
xnor U2093 (N_2093,N_1943,N_1935);
or U2094 (N_2094,N_1928,N_1969);
nor U2095 (N_2095,N_1978,N_1822);
or U2096 (N_2096,N_1898,N_1929);
nand U2097 (N_2097,N_1841,N_1837);
xor U2098 (N_2098,N_1905,N_1903);
nor U2099 (N_2099,N_1972,N_1968);
or U2100 (N_2100,N_1803,N_1883);
or U2101 (N_2101,N_1946,N_1920);
and U2102 (N_2102,N_1824,N_1866);
and U2103 (N_2103,N_1899,N_1873);
or U2104 (N_2104,N_1857,N_1896);
nor U2105 (N_2105,N_1975,N_1937);
and U2106 (N_2106,N_1981,N_1916);
nor U2107 (N_2107,N_1870,N_1982);
nor U2108 (N_2108,N_1915,N_1904);
or U2109 (N_2109,N_1917,N_1915);
or U2110 (N_2110,N_1802,N_1919);
and U2111 (N_2111,N_1903,N_1937);
and U2112 (N_2112,N_1853,N_1884);
nor U2113 (N_2113,N_1887,N_1871);
nand U2114 (N_2114,N_1862,N_1885);
nor U2115 (N_2115,N_1815,N_1806);
and U2116 (N_2116,N_1987,N_1936);
and U2117 (N_2117,N_1986,N_1974);
and U2118 (N_2118,N_1850,N_1856);
and U2119 (N_2119,N_1927,N_1991);
or U2120 (N_2120,N_1805,N_1908);
nor U2121 (N_2121,N_1871,N_1984);
and U2122 (N_2122,N_1969,N_1944);
nor U2123 (N_2123,N_1843,N_1927);
nor U2124 (N_2124,N_1815,N_1835);
and U2125 (N_2125,N_1965,N_1893);
xnor U2126 (N_2126,N_1818,N_1930);
nor U2127 (N_2127,N_1898,N_1853);
or U2128 (N_2128,N_1867,N_1990);
nor U2129 (N_2129,N_1916,N_1926);
xnor U2130 (N_2130,N_1846,N_1877);
nand U2131 (N_2131,N_1970,N_1996);
nor U2132 (N_2132,N_1926,N_1999);
nor U2133 (N_2133,N_1812,N_1848);
and U2134 (N_2134,N_1971,N_1899);
nand U2135 (N_2135,N_1930,N_1895);
and U2136 (N_2136,N_1862,N_1832);
or U2137 (N_2137,N_1877,N_1847);
and U2138 (N_2138,N_1880,N_1857);
nand U2139 (N_2139,N_1938,N_1848);
and U2140 (N_2140,N_1821,N_1890);
or U2141 (N_2141,N_1910,N_1815);
xnor U2142 (N_2142,N_1857,N_1998);
or U2143 (N_2143,N_1984,N_1947);
and U2144 (N_2144,N_1808,N_1917);
or U2145 (N_2145,N_1941,N_1984);
nor U2146 (N_2146,N_1866,N_1837);
nand U2147 (N_2147,N_1988,N_1973);
nand U2148 (N_2148,N_1884,N_1812);
nand U2149 (N_2149,N_1828,N_1929);
or U2150 (N_2150,N_1898,N_1873);
nor U2151 (N_2151,N_1871,N_1903);
nand U2152 (N_2152,N_1866,N_1924);
nand U2153 (N_2153,N_1869,N_1833);
nor U2154 (N_2154,N_1969,N_1818);
and U2155 (N_2155,N_1925,N_1894);
nand U2156 (N_2156,N_1984,N_1885);
and U2157 (N_2157,N_1861,N_1923);
and U2158 (N_2158,N_1993,N_1985);
and U2159 (N_2159,N_1880,N_1822);
xnor U2160 (N_2160,N_1938,N_1822);
and U2161 (N_2161,N_1803,N_1952);
or U2162 (N_2162,N_1867,N_1869);
and U2163 (N_2163,N_1848,N_1903);
nor U2164 (N_2164,N_1888,N_1848);
nand U2165 (N_2165,N_1837,N_1848);
or U2166 (N_2166,N_1845,N_1847);
or U2167 (N_2167,N_1917,N_1831);
nor U2168 (N_2168,N_1884,N_1958);
nor U2169 (N_2169,N_1907,N_1800);
or U2170 (N_2170,N_1988,N_1960);
nand U2171 (N_2171,N_1908,N_1881);
and U2172 (N_2172,N_1871,N_1963);
or U2173 (N_2173,N_1804,N_1960);
nor U2174 (N_2174,N_1869,N_1996);
nor U2175 (N_2175,N_1900,N_1836);
xnor U2176 (N_2176,N_1935,N_1953);
and U2177 (N_2177,N_1824,N_1973);
xor U2178 (N_2178,N_1839,N_1966);
nand U2179 (N_2179,N_1986,N_1903);
nor U2180 (N_2180,N_1804,N_1828);
or U2181 (N_2181,N_1831,N_1911);
nor U2182 (N_2182,N_1981,N_1827);
nor U2183 (N_2183,N_1922,N_1850);
nand U2184 (N_2184,N_1925,N_1846);
nor U2185 (N_2185,N_1887,N_1836);
nand U2186 (N_2186,N_1816,N_1990);
nand U2187 (N_2187,N_1907,N_1850);
nor U2188 (N_2188,N_1809,N_1958);
nor U2189 (N_2189,N_1827,N_1834);
or U2190 (N_2190,N_1861,N_1855);
or U2191 (N_2191,N_1949,N_1921);
nand U2192 (N_2192,N_1871,N_1826);
or U2193 (N_2193,N_1990,N_1854);
nand U2194 (N_2194,N_1917,N_1804);
nand U2195 (N_2195,N_1840,N_1831);
nand U2196 (N_2196,N_1934,N_1838);
nor U2197 (N_2197,N_1859,N_1954);
or U2198 (N_2198,N_1914,N_1898);
xnor U2199 (N_2199,N_1903,N_1813);
and U2200 (N_2200,N_2114,N_2063);
nand U2201 (N_2201,N_2019,N_2193);
and U2202 (N_2202,N_2059,N_2190);
and U2203 (N_2203,N_2169,N_2108);
nand U2204 (N_2204,N_2198,N_2180);
nor U2205 (N_2205,N_2024,N_2174);
nand U2206 (N_2206,N_2022,N_2181);
or U2207 (N_2207,N_2099,N_2153);
and U2208 (N_2208,N_2138,N_2112);
or U2209 (N_2209,N_2189,N_2034);
nor U2210 (N_2210,N_2003,N_2160);
and U2211 (N_2211,N_2170,N_2026);
or U2212 (N_2212,N_2135,N_2117);
or U2213 (N_2213,N_2044,N_2009);
nand U2214 (N_2214,N_2161,N_2074);
and U2215 (N_2215,N_2113,N_2191);
and U2216 (N_2216,N_2071,N_2076);
and U2217 (N_2217,N_2131,N_2148);
xor U2218 (N_2218,N_2079,N_2168);
xor U2219 (N_2219,N_2029,N_2098);
or U2220 (N_2220,N_2091,N_2163);
nor U2221 (N_2221,N_2109,N_2197);
nor U2222 (N_2222,N_2110,N_2083);
or U2223 (N_2223,N_2152,N_2192);
nor U2224 (N_2224,N_2040,N_2183);
or U2225 (N_2225,N_2142,N_2036);
nand U2226 (N_2226,N_2042,N_2008);
or U2227 (N_2227,N_2014,N_2030);
and U2228 (N_2228,N_2171,N_2082);
nand U2229 (N_2229,N_2066,N_2058);
nand U2230 (N_2230,N_2010,N_2186);
nor U2231 (N_2231,N_2055,N_2086);
xnor U2232 (N_2232,N_2089,N_2027);
nor U2233 (N_2233,N_2023,N_2165);
nor U2234 (N_2234,N_2145,N_2122);
nor U2235 (N_2235,N_2050,N_2007);
nor U2236 (N_2236,N_2123,N_2133);
nand U2237 (N_2237,N_2032,N_2143);
xor U2238 (N_2238,N_2053,N_2105);
and U2239 (N_2239,N_2048,N_2062);
nand U2240 (N_2240,N_2103,N_2031);
xnor U2241 (N_2241,N_2096,N_2176);
nor U2242 (N_2242,N_2144,N_2187);
and U2243 (N_2243,N_2039,N_2139);
nor U2244 (N_2244,N_2017,N_2178);
and U2245 (N_2245,N_2000,N_2068);
and U2246 (N_2246,N_2038,N_2107);
or U2247 (N_2247,N_2167,N_2177);
or U2248 (N_2248,N_2199,N_2094);
xor U2249 (N_2249,N_2060,N_2175);
nor U2250 (N_2250,N_2173,N_2188);
nor U2251 (N_2251,N_2116,N_2052);
nand U2252 (N_2252,N_2021,N_2118);
nand U2253 (N_2253,N_2106,N_2057);
and U2254 (N_2254,N_2157,N_2124);
nand U2255 (N_2255,N_2051,N_2127);
and U2256 (N_2256,N_2047,N_2182);
nor U2257 (N_2257,N_2046,N_2156);
or U2258 (N_2258,N_2061,N_2164);
or U2259 (N_2259,N_2016,N_2125);
nand U2260 (N_2260,N_2100,N_2077);
xnor U2261 (N_2261,N_2101,N_2056);
nand U2262 (N_2262,N_2078,N_2080);
xor U2263 (N_2263,N_2011,N_2088);
nor U2264 (N_2264,N_2025,N_2045);
or U2265 (N_2265,N_2179,N_2041);
or U2266 (N_2266,N_2137,N_2129);
and U2267 (N_2267,N_2097,N_2006);
and U2268 (N_2268,N_2013,N_2162);
or U2269 (N_2269,N_2049,N_2070);
xnor U2270 (N_2270,N_2111,N_2195);
nor U2271 (N_2271,N_2085,N_2035);
and U2272 (N_2272,N_2102,N_2075);
nor U2273 (N_2273,N_2081,N_2194);
and U2274 (N_2274,N_2095,N_2155);
or U2275 (N_2275,N_2064,N_2128);
nand U2276 (N_2276,N_2004,N_2158);
xor U2277 (N_2277,N_2130,N_2149);
and U2278 (N_2278,N_2033,N_2172);
and U2279 (N_2279,N_2012,N_2136);
nand U2280 (N_2280,N_2154,N_2185);
or U2281 (N_2281,N_2015,N_2054);
nor U2282 (N_2282,N_2120,N_2001);
nor U2283 (N_2283,N_2134,N_2147);
or U2284 (N_2284,N_2092,N_2141);
and U2285 (N_2285,N_2132,N_2184);
nand U2286 (N_2286,N_2090,N_2002);
and U2287 (N_2287,N_2073,N_2084);
nor U2288 (N_2288,N_2067,N_2140);
xor U2289 (N_2289,N_2087,N_2043);
and U2290 (N_2290,N_2166,N_2065);
nand U2291 (N_2291,N_2018,N_2196);
nor U2292 (N_2292,N_2151,N_2069);
nor U2293 (N_2293,N_2020,N_2005);
nor U2294 (N_2294,N_2150,N_2119);
and U2295 (N_2295,N_2093,N_2126);
nand U2296 (N_2296,N_2028,N_2121);
xnor U2297 (N_2297,N_2037,N_2146);
or U2298 (N_2298,N_2115,N_2159);
and U2299 (N_2299,N_2104,N_2072);
xor U2300 (N_2300,N_2125,N_2114);
xnor U2301 (N_2301,N_2076,N_2098);
nand U2302 (N_2302,N_2102,N_2099);
nor U2303 (N_2303,N_2038,N_2192);
nor U2304 (N_2304,N_2137,N_2064);
nand U2305 (N_2305,N_2089,N_2021);
nand U2306 (N_2306,N_2066,N_2199);
nand U2307 (N_2307,N_2020,N_2169);
and U2308 (N_2308,N_2187,N_2081);
or U2309 (N_2309,N_2088,N_2055);
nand U2310 (N_2310,N_2171,N_2025);
nand U2311 (N_2311,N_2115,N_2064);
nand U2312 (N_2312,N_2142,N_2188);
and U2313 (N_2313,N_2024,N_2147);
nor U2314 (N_2314,N_2096,N_2069);
or U2315 (N_2315,N_2139,N_2076);
and U2316 (N_2316,N_2198,N_2012);
and U2317 (N_2317,N_2194,N_2100);
and U2318 (N_2318,N_2168,N_2042);
nand U2319 (N_2319,N_2084,N_2013);
or U2320 (N_2320,N_2033,N_2135);
nand U2321 (N_2321,N_2029,N_2051);
and U2322 (N_2322,N_2083,N_2087);
nand U2323 (N_2323,N_2072,N_2089);
and U2324 (N_2324,N_2006,N_2138);
nor U2325 (N_2325,N_2101,N_2010);
nand U2326 (N_2326,N_2123,N_2199);
or U2327 (N_2327,N_2032,N_2000);
or U2328 (N_2328,N_2025,N_2009);
or U2329 (N_2329,N_2031,N_2174);
nand U2330 (N_2330,N_2056,N_2096);
nor U2331 (N_2331,N_2162,N_2186);
or U2332 (N_2332,N_2112,N_2127);
and U2333 (N_2333,N_2012,N_2003);
xor U2334 (N_2334,N_2001,N_2034);
and U2335 (N_2335,N_2123,N_2128);
xnor U2336 (N_2336,N_2017,N_2129);
xnor U2337 (N_2337,N_2156,N_2000);
or U2338 (N_2338,N_2086,N_2164);
nor U2339 (N_2339,N_2118,N_2117);
and U2340 (N_2340,N_2142,N_2110);
and U2341 (N_2341,N_2090,N_2143);
nor U2342 (N_2342,N_2079,N_2036);
nor U2343 (N_2343,N_2040,N_2078);
and U2344 (N_2344,N_2048,N_2034);
xnor U2345 (N_2345,N_2178,N_2123);
or U2346 (N_2346,N_2048,N_2144);
nor U2347 (N_2347,N_2159,N_2156);
nand U2348 (N_2348,N_2150,N_2172);
and U2349 (N_2349,N_2028,N_2175);
or U2350 (N_2350,N_2111,N_2021);
nand U2351 (N_2351,N_2091,N_2021);
or U2352 (N_2352,N_2194,N_2170);
nor U2353 (N_2353,N_2060,N_2170);
nor U2354 (N_2354,N_2178,N_2114);
and U2355 (N_2355,N_2029,N_2078);
and U2356 (N_2356,N_2110,N_2053);
nor U2357 (N_2357,N_2067,N_2058);
nor U2358 (N_2358,N_2184,N_2065);
xor U2359 (N_2359,N_2007,N_2076);
and U2360 (N_2360,N_2117,N_2122);
or U2361 (N_2361,N_2143,N_2075);
nor U2362 (N_2362,N_2070,N_2174);
nand U2363 (N_2363,N_2042,N_2152);
nand U2364 (N_2364,N_2000,N_2062);
nand U2365 (N_2365,N_2034,N_2196);
nand U2366 (N_2366,N_2103,N_2194);
and U2367 (N_2367,N_2136,N_2062);
or U2368 (N_2368,N_2001,N_2085);
xnor U2369 (N_2369,N_2061,N_2063);
and U2370 (N_2370,N_2056,N_2040);
xor U2371 (N_2371,N_2135,N_2122);
nand U2372 (N_2372,N_2149,N_2170);
or U2373 (N_2373,N_2166,N_2051);
nand U2374 (N_2374,N_2039,N_2185);
or U2375 (N_2375,N_2068,N_2166);
nand U2376 (N_2376,N_2108,N_2017);
nand U2377 (N_2377,N_2070,N_2091);
or U2378 (N_2378,N_2049,N_2150);
and U2379 (N_2379,N_2172,N_2013);
and U2380 (N_2380,N_2169,N_2135);
nand U2381 (N_2381,N_2044,N_2185);
nor U2382 (N_2382,N_2054,N_2181);
nor U2383 (N_2383,N_2165,N_2084);
and U2384 (N_2384,N_2170,N_2177);
nor U2385 (N_2385,N_2191,N_2197);
and U2386 (N_2386,N_2061,N_2070);
or U2387 (N_2387,N_2083,N_2115);
nor U2388 (N_2388,N_2089,N_2161);
or U2389 (N_2389,N_2131,N_2087);
or U2390 (N_2390,N_2020,N_2190);
and U2391 (N_2391,N_2052,N_2083);
and U2392 (N_2392,N_2082,N_2097);
nor U2393 (N_2393,N_2143,N_2006);
and U2394 (N_2394,N_2180,N_2169);
or U2395 (N_2395,N_2197,N_2030);
and U2396 (N_2396,N_2003,N_2156);
nand U2397 (N_2397,N_2083,N_2015);
nor U2398 (N_2398,N_2081,N_2011);
nand U2399 (N_2399,N_2024,N_2102);
nor U2400 (N_2400,N_2335,N_2352);
or U2401 (N_2401,N_2289,N_2366);
and U2402 (N_2402,N_2328,N_2355);
nand U2403 (N_2403,N_2395,N_2264);
and U2404 (N_2404,N_2315,N_2287);
and U2405 (N_2405,N_2340,N_2276);
and U2406 (N_2406,N_2344,N_2338);
or U2407 (N_2407,N_2280,N_2269);
xor U2408 (N_2408,N_2250,N_2364);
nand U2409 (N_2409,N_2374,N_2293);
nand U2410 (N_2410,N_2313,N_2390);
nand U2411 (N_2411,N_2296,N_2391);
and U2412 (N_2412,N_2380,N_2388);
nor U2413 (N_2413,N_2238,N_2257);
and U2414 (N_2414,N_2350,N_2327);
or U2415 (N_2415,N_2259,N_2375);
or U2416 (N_2416,N_2399,N_2334);
nand U2417 (N_2417,N_2235,N_2319);
and U2418 (N_2418,N_2249,N_2256);
nor U2419 (N_2419,N_2365,N_2225);
and U2420 (N_2420,N_2255,N_2318);
or U2421 (N_2421,N_2228,N_2201);
nand U2422 (N_2422,N_2370,N_2215);
and U2423 (N_2423,N_2292,N_2302);
and U2424 (N_2424,N_2314,N_2273);
nor U2425 (N_2425,N_2301,N_2279);
nand U2426 (N_2426,N_2231,N_2299);
nor U2427 (N_2427,N_2241,N_2252);
nor U2428 (N_2428,N_2227,N_2378);
and U2429 (N_2429,N_2376,N_2371);
or U2430 (N_2430,N_2271,N_2308);
xnor U2431 (N_2431,N_2382,N_2267);
nand U2432 (N_2432,N_2357,N_2326);
nor U2433 (N_2433,N_2220,N_2331);
or U2434 (N_2434,N_2351,N_2211);
nor U2435 (N_2435,N_2266,N_2345);
or U2436 (N_2436,N_2372,N_2310);
xor U2437 (N_2437,N_2290,N_2222);
and U2438 (N_2438,N_2258,N_2224);
nor U2439 (N_2439,N_2216,N_2284);
nor U2440 (N_2440,N_2393,N_2236);
nand U2441 (N_2441,N_2368,N_2341);
or U2442 (N_2442,N_2226,N_2298);
and U2443 (N_2443,N_2300,N_2398);
and U2444 (N_2444,N_2363,N_2209);
or U2445 (N_2445,N_2200,N_2387);
or U2446 (N_2446,N_2307,N_2281);
and U2447 (N_2447,N_2207,N_2322);
and U2448 (N_2448,N_2294,N_2240);
and U2449 (N_2449,N_2333,N_2362);
xor U2450 (N_2450,N_2246,N_2320);
nor U2451 (N_2451,N_2247,N_2316);
and U2452 (N_2452,N_2379,N_2213);
xor U2453 (N_2453,N_2263,N_2278);
xnor U2454 (N_2454,N_2277,N_2288);
nand U2455 (N_2455,N_2306,N_2237);
nand U2456 (N_2456,N_2384,N_2285);
xnor U2457 (N_2457,N_2274,N_2356);
nor U2458 (N_2458,N_2309,N_2261);
nand U2459 (N_2459,N_2304,N_2212);
nor U2460 (N_2460,N_2381,N_2230);
or U2461 (N_2461,N_2354,N_2223);
nor U2462 (N_2462,N_2324,N_2275);
nor U2463 (N_2463,N_2358,N_2339);
nor U2464 (N_2464,N_2373,N_2330);
and U2465 (N_2465,N_2233,N_2346);
or U2466 (N_2466,N_2234,N_2386);
and U2467 (N_2467,N_2303,N_2253);
nor U2468 (N_2468,N_2360,N_2217);
and U2469 (N_2469,N_2348,N_2396);
xnor U2470 (N_2470,N_2260,N_2336);
and U2471 (N_2471,N_2206,N_2251);
and U2472 (N_2472,N_2337,N_2347);
nor U2473 (N_2473,N_2332,N_2282);
and U2474 (N_2474,N_2286,N_2392);
nor U2475 (N_2475,N_2394,N_2349);
and U2476 (N_2476,N_2218,N_2268);
and U2477 (N_2477,N_2270,N_2219);
nand U2478 (N_2478,N_2353,N_2202);
nand U2479 (N_2479,N_2305,N_2323);
nand U2480 (N_2480,N_2389,N_2208);
or U2481 (N_2481,N_2272,N_2311);
and U2482 (N_2482,N_2245,N_2239);
nand U2483 (N_2483,N_2321,N_2369);
nand U2484 (N_2484,N_2203,N_2221);
nor U2485 (N_2485,N_2329,N_2385);
nand U2486 (N_2486,N_2325,N_2359);
and U2487 (N_2487,N_2214,N_2204);
or U2488 (N_2488,N_2283,N_2229);
or U2489 (N_2489,N_2244,N_2291);
nand U2490 (N_2490,N_2254,N_2383);
and U2491 (N_2491,N_2205,N_2265);
nor U2492 (N_2492,N_2295,N_2297);
xnor U2493 (N_2493,N_2317,N_2343);
xor U2494 (N_2494,N_2248,N_2367);
nand U2495 (N_2495,N_2243,N_2361);
nor U2496 (N_2496,N_2262,N_2312);
nor U2497 (N_2497,N_2232,N_2342);
or U2498 (N_2498,N_2210,N_2397);
nand U2499 (N_2499,N_2377,N_2242);
xnor U2500 (N_2500,N_2372,N_2347);
nor U2501 (N_2501,N_2285,N_2241);
nand U2502 (N_2502,N_2229,N_2303);
and U2503 (N_2503,N_2308,N_2384);
nor U2504 (N_2504,N_2311,N_2202);
xnor U2505 (N_2505,N_2370,N_2348);
nor U2506 (N_2506,N_2205,N_2231);
or U2507 (N_2507,N_2348,N_2367);
nor U2508 (N_2508,N_2220,N_2269);
and U2509 (N_2509,N_2269,N_2318);
nor U2510 (N_2510,N_2265,N_2291);
or U2511 (N_2511,N_2376,N_2244);
nand U2512 (N_2512,N_2388,N_2215);
or U2513 (N_2513,N_2310,N_2276);
nand U2514 (N_2514,N_2202,N_2283);
xnor U2515 (N_2515,N_2342,N_2329);
or U2516 (N_2516,N_2393,N_2279);
nor U2517 (N_2517,N_2361,N_2255);
and U2518 (N_2518,N_2275,N_2359);
and U2519 (N_2519,N_2213,N_2352);
nand U2520 (N_2520,N_2222,N_2251);
and U2521 (N_2521,N_2230,N_2395);
nand U2522 (N_2522,N_2300,N_2307);
and U2523 (N_2523,N_2217,N_2300);
or U2524 (N_2524,N_2282,N_2289);
nor U2525 (N_2525,N_2343,N_2345);
or U2526 (N_2526,N_2316,N_2393);
nor U2527 (N_2527,N_2359,N_2257);
nand U2528 (N_2528,N_2274,N_2328);
and U2529 (N_2529,N_2318,N_2295);
and U2530 (N_2530,N_2230,N_2285);
nor U2531 (N_2531,N_2332,N_2389);
and U2532 (N_2532,N_2363,N_2235);
nand U2533 (N_2533,N_2228,N_2386);
nand U2534 (N_2534,N_2390,N_2354);
xnor U2535 (N_2535,N_2291,N_2325);
or U2536 (N_2536,N_2237,N_2362);
nand U2537 (N_2537,N_2240,N_2238);
and U2538 (N_2538,N_2335,N_2226);
or U2539 (N_2539,N_2399,N_2310);
nor U2540 (N_2540,N_2364,N_2223);
nor U2541 (N_2541,N_2275,N_2218);
and U2542 (N_2542,N_2310,N_2362);
nand U2543 (N_2543,N_2343,N_2251);
and U2544 (N_2544,N_2368,N_2225);
or U2545 (N_2545,N_2291,N_2387);
and U2546 (N_2546,N_2256,N_2312);
and U2547 (N_2547,N_2320,N_2212);
and U2548 (N_2548,N_2243,N_2330);
xor U2549 (N_2549,N_2398,N_2288);
or U2550 (N_2550,N_2308,N_2228);
nor U2551 (N_2551,N_2286,N_2276);
and U2552 (N_2552,N_2338,N_2319);
or U2553 (N_2553,N_2325,N_2395);
and U2554 (N_2554,N_2238,N_2219);
nand U2555 (N_2555,N_2271,N_2231);
and U2556 (N_2556,N_2247,N_2332);
or U2557 (N_2557,N_2288,N_2376);
xor U2558 (N_2558,N_2228,N_2218);
nand U2559 (N_2559,N_2221,N_2379);
and U2560 (N_2560,N_2321,N_2366);
nand U2561 (N_2561,N_2328,N_2352);
and U2562 (N_2562,N_2373,N_2221);
or U2563 (N_2563,N_2371,N_2250);
nor U2564 (N_2564,N_2273,N_2368);
and U2565 (N_2565,N_2313,N_2295);
nand U2566 (N_2566,N_2398,N_2241);
or U2567 (N_2567,N_2292,N_2395);
or U2568 (N_2568,N_2217,N_2398);
nand U2569 (N_2569,N_2302,N_2374);
and U2570 (N_2570,N_2259,N_2266);
nand U2571 (N_2571,N_2228,N_2382);
or U2572 (N_2572,N_2288,N_2221);
or U2573 (N_2573,N_2399,N_2241);
and U2574 (N_2574,N_2279,N_2226);
or U2575 (N_2575,N_2270,N_2260);
nand U2576 (N_2576,N_2255,N_2368);
and U2577 (N_2577,N_2213,N_2251);
and U2578 (N_2578,N_2227,N_2290);
nand U2579 (N_2579,N_2326,N_2261);
and U2580 (N_2580,N_2278,N_2247);
xor U2581 (N_2581,N_2369,N_2305);
nand U2582 (N_2582,N_2347,N_2364);
and U2583 (N_2583,N_2242,N_2277);
and U2584 (N_2584,N_2328,N_2296);
and U2585 (N_2585,N_2258,N_2315);
xnor U2586 (N_2586,N_2259,N_2378);
and U2587 (N_2587,N_2390,N_2318);
and U2588 (N_2588,N_2336,N_2351);
and U2589 (N_2589,N_2243,N_2276);
nor U2590 (N_2590,N_2375,N_2383);
or U2591 (N_2591,N_2226,N_2269);
and U2592 (N_2592,N_2284,N_2339);
nor U2593 (N_2593,N_2320,N_2384);
and U2594 (N_2594,N_2282,N_2219);
nand U2595 (N_2595,N_2245,N_2244);
nand U2596 (N_2596,N_2324,N_2259);
or U2597 (N_2597,N_2300,N_2287);
and U2598 (N_2598,N_2249,N_2301);
nand U2599 (N_2599,N_2345,N_2228);
nor U2600 (N_2600,N_2512,N_2565);
nor U2601 (N_2601,N_2567,N_2453);
nor U2602 (N_2602,N_2548,N_2588);
nand U2603 (N_2603,N_2595,N_2582);
nand U2604 (N_2604,N_2504,N_2463);
nor U2605 (N_2605,N_2473,N_2518);
and U2606 (N_2606,N_2510,N_2415);
nand U2607 (N_2607,N_2498,N_2581);
nor U2608 (N_2608,N_2449,N_2490);
or U2609 (N_2609,N_2487,N_2441);
or U2610 (N_2610,N_2533,N_2444);
or U2611 (N_2611,N_2539,N_2575);
or U2612 (N_2612,N_2553,N_2592);
or U2613 (N_2613,N_2486,N_2438);
xnor U2614 (N_2614,N_2416,N_2437);
or U2615 (N_2615,N_2541,N_2430);
or U2616 (N_2616,N_2400,N_2421);
nand U2617 (N_2617,N_2524,N_2491);
or U2618 (N_2618,N_2420,N_2464);
and U2619 (N_2619,N_2589,N_2440);
nand U2620 (N_2620,N_2591,N_2513);
nand U2621 (N_2621,N_2455,N_2507);
nor U2622 (N_2622,N_2443,N_2471);
or U2623 (N_2623,N_2418,N_2542);
and U2624 (N_2624,N_2561,N_2427);
and U2625 (N_2625,N_2482,N_2563);
nor U2626 (N_2626,N_2517,N_2452);
and U2627 (N_2627,N_2509,N_2496);
nand U2628 (N_2628,N_2599,N_2478);
and U2629 (N_2629,N_2483,N_2521);
nand U2630 (N_2630,N_2404,N_2479);
nor U2631 (N_2631,N_2562,N_2428);
and U2632 (N_2632,N_2474,N_2422);
or U2633 (N_2633,N_2554,N_2556);
and U2634 (N_2634,N_2550,N_2499);
nand U2635 (N_2635,N_2508,N_2451);
nor U2636 (N_2636,N_2450,N_2411);
nand U2637 (N_2637,N_2497,N_2578);
or U2638 (N_2638,N_2472,N_2477);
and U2639 (N_2639,N_2445,N_2585);
nand U2640 (N_2640,N_2405,N_2590);
xor U2641 (N_2641,N_2489,N_2406);
nor U2642 (N_2642,N_2564,N_2429);
nor U2643 (N_2643,N_2460,N_2540);
nor U2644 (N_2644,N_2557,N_2447);
or U2645 (N_2645,N_2537,N_2555);
nand U2646 (N_2646,N_2500,N_2527);
or U2647 (N_2647,N_2596,N_2426);
nor U2648 (N_2648,N_2417,N_2572);
and U2649 (N_2649,N_2543,N_2506);
and U2650 (N_2650,N_2593,N_2401);
or U2651 (N_2651,N_2439,N_2485);
nand U2652 (N_2652,N_2461,N_2546);
xor U2653 (N_2653,N_2403,N_2414);
nor U2654 (N_2654,N_2570,N_2568);
or U2655 (N_2655,N_2419,N_2466);
and U2656 (N_2656,N_2505,N_2494);
nor U2657 (N_2657,N_2462,N_2402);
nand U2658 (N_2658,N_2410,N_2534);
or U2659 (N_2659,N_2523,N_2425);
nand U2660 (N_2660,N_2467,N_2431);
nand U2661 (N_2661,N_2514,N_2434);
nand U2662 (N_2662,N_2424,N_2583);
or U2663 (N_2663,N_2545,N_2488);
nor U2664 (N_2664,N_2480,N_2409);
nor U2665 (N_2665,N_2526,N_2529);
nor U2666 (N_2666,N_2412,N_2502);
nand U2667 (N_2667,N_2525,N_2587);
xnor U2668 (N_2668,N_2530,N_2594);
xnor U2669 (N_2669,N_2566,N_2597);
or U2670 (N_2670,N_2558,N_2551);
and U2671 (N_2671,N_2580,N_2519);
nor U2672 (N_2672,N_2535,N_2468);
and U2673 (N_2673,N_2501,N_2432);
or U2674 (N_2674,N_2436,N_2458);
or U2675 (N_2675,N_2520,N_2569);
nor U2676 (N_2676,N_2538,N_2536);
or U2677 (N_2677,N_2465,N_2469);
and U2678 (N_2678,N_2515,N_2577);
and U2679 (N_2679,N_2407,N_2576);
and U2680 (N_2680,N_2484,N_2586);
or U2681 (N_2681,N_2481,N_2584);
nand U2682 (N_2682,N_2448,N_2459);
and U2683 (N_2683,N_2531,N_2446);
nor U2684 (N_2684,N_2559,N_2532);
and U2685 (N_2685,N_2408,N_2552);
nand U2686 (N_2686,N_2598,N_2470);
nor U2687 (N_2687,N_2573,N_2493);
and U2688 (N_2688,N_2475,N_2423);
nand U2689 (N_2689,N_2457,N_2511);
nor U2690 (N_2690,N_2456,N_2560);
xor U2691 (N_2691,N_2476,N_2544);
and U2692 (N_2692,N_2495,N_2574);
nor U2693 (N_2693,N_2503,N_2579);
or U2694 (N_2694,N_2522,N_2492);
and U2695 (N_2695,N_2442,N_2454);
and U2696 (N_2696,N_2528,N_2571);
or U2697 (N_2697,N_2433,N_2547);
and U2698 (N_2698,N_2549,N_2435);
or U2699 (N_2699,N_2516,N_2413);
nand U2700 (N_2700,N_2547,N_2567);
and U2701 (N_2701,N_2415,N_2507);
nand U2702 (N_2702,N_2401,N_2536);
or U2703 (N_2703,N_2436,N_2574);
or U2704 (N_2704,N_2425,N_2413);
nand U2705 (N_2705,N_2459,N_2537);
and U2706 (N_2706,N_2437,N_2443);
or U2707 (N_2707,N_2480,N_2531);
nor U2708 (N_2708,N_2435,N_2462);
xnor U2709 (N_2709,N_2494,N_2564);
and U2710 (N_2710,N_2520,N_2459);
nor U2711 (N_2711,N_2561,N_2510);
nor U2712 (N_2712,N_2518,N_2442);
or U2713 (N_2713,N_2596,N_2406);
and U2714 (N_2714,N_2413,N_2493);
nand U2715 (N_2715,N_2536,N_2559);
nor U2716 (N_2716,N_2552,N_2452);
nor U2717 (N_2717,N_2553,N_2519);
or U2718 (N_2718,N_2514,N_2588);
and U2719 (N_2719,N_2468,N_2565);
or U2720 (N_2720,N_2491,N_2409);
nand U2721 (N_2721,N_2526,N_2507);
nand U2722 (N_2722,N_2453,N_2416);
nand U2723 (N_2723,N_2557,N_2473);
xnor U2724 (N_2724,N_2578,N_2558);
or U2725 (N_2725,N_2455,N_2478);
nand U2726 (N_2726,N_2487,N_2535);
nor U2727 (N_2727,N_2459,N_2517);
and U2728 (N_2728,N_2473,N_2456);
nand U2729 (N_2729,N_2460,N_2536);
nor U2730 (N_2730,N_2464,N_2438);
or U2731 (N_2731,N_2409,N_2435);
nand U2732 (N_2732,N_2491,N_2481);
or U2733 (N_2733,N_2441,N_2511);
nand U2734 (N_2734,N_2447,N_2598);
xor U2735 (N_2735,N_2442,N_2534);
and U2736 (N_2736,N_2507,N_2508);
and U2737 (N_2737,N_2563,N_2461);
nor U2738 (N_2738,N_2571,N_2494);
nor U2739 (N_2739,N_2434,N_2528);
nand U2740 (N_2740,N_2492,N_2464);
nand U2741 (N_2741,N_2514,N_2595);
nor U2742 (N_2742,N_2546,N_2518);
nand U2743 (N_2743,N_2485,N_2571);
nand U2744 (N_2744,N_2492,N_2469);
or U2745 (N_2745,N_2593,N_2516);
and U2746 (N_2746,N_2579,N_2569);
nand U2747 (N_2747,N_2586,N_2454);
and U2748 (N_2748,N_2477,N_2597);
and U2749 (N_2749,N_2476,N_2487);
xor U2750 (N_2750,N_2538,N_2523);
and U2751 (N_2751,N_2413,N_2597);
or U2752 (N_2752,N_2527,N_2588);
and U2753 (N_2753,N_2487,N_2537);
nand U2754 (N_2754,N_2569,N_2571);
or U2755 (N_2755,N_2419,N_2449);
or U2756 (N_2756,N_2457,N_2525);
or U2757 (N_2757,N_2499,N_2410);
and U2758 (N_2758,N_2403,N_2431);
and U2759 (N_2759,N_2563,N_2448);
nand U2760 (N_2760,N_2418,N_2512);
and U2761 (N_2761,N_2451,N_2463);
nand U2762 (N_2762,N_2508,N_2541);
and U2763 (N_2763,N_2483,N_2543);
and U2764 (N_2764,N_2502,N_2451);
or U2765 (N_2765,N_2529,N_2443);
or U2766 (N_2766,N_2549,N_2525);
nand U2767 (N_2767,N_2591,N_2407);
nand U2768 (N_2768,N_2489,N_2416);
nor U2769 (N_2769,N_2481,N_2423);
and U2770 (N_2770,N_2424,N_2570);
nor U2771 (N_2771,N_2434,N_2575);
and U2772 (N_2772,N_2421,N_2575);
nor U2773 (N_2773,N_2475,N_2469);
nand U2774 (N_2774,N_2572,N_2471);
and U2775 (N_2775,N_2557,N_2458);
nor U2776 (N_2776,N_2425,N_2423);
nor U2777 (N_2777,N_2475,N_2555);
nor U2778 (N_2778,N_2471,N_2431);
and U2779 (N_2779,N_2459,N_2548);
or U2780 (N_2780,N_2527,N_2478);
nor U2781 (N_2781,N_2436,N_2558);
nor U2782 (N_2782,N_2519,N_2482);
nor U2783 (N_2783,N_2485,N_2567);
nor U2784 (N_2784,N_2451,N_2445);
nand U2785 (N_2785,N_2407,N_2493);
nor U2786 (N_2786,N_2509,N_2422);
nand U2787 (N_2787,N_2574,N_2464);
or U2788 (N_2788,N_2518,N_2590);
nor U2789 (N_2789,N_2513,N_2593);
or U2790 (N_2790,N_2464,N_2541);
nand U2791 (N_2791,N_2460,N_2507);
nand U2792 (N_2792,N_2459,N_2585);
nand U2793 (N_2793,N_2539,N_2511);
or U2794 (N_2794,N_2454,N_2536);
nand U2795 (N_2795,N_2460,N_2487);
nor U2796 (N_2796,N_2552,N_2418);
and U2797 (N_2797,N_2464,N_2496);
or U2798 (N_2798,N_2474,N_2492);
and U2799 (N_2799,N_2572,N_2478);
nor U2800 (N_2800,N_2622,N_2689);
nor U2801 (N_2801,N_2798,N_2773);
and U2802 (N_2802,N_2657,N_2619);
xnor U2803 (N_2803,N_2648,N_2610);
and U2804 (N_2804,N_2741,N_2733);
and U2805 (N_2805,N_2656,N_2639);
nor U2806 (N_2806,N_2791,N_2721);
or U2807 (N_2807,N_2718,N_2654);
nand U2808 (N_2808,N_2603,N_2613);
or U2809 (N_2809,N_2694,N_2615);
xor U2810 (N_2810,N_2618,N_2759);
nor U2811 (N_2811,N_2784,N_2680);
or U2812 (N_2812,N_2792,N_2761);
or U2813 (N_2813,N_2658,N_2730);
and U2814 (N_2814,N_2602,N_2663);
or U2815 (N_2815,N_2712,N_2703);
and U2816 (N_2816,N_2769,N_2725);
nand U2817 (N_2817,N_2749,N_2647);
nor U2818 (N_2818,N_2624,N_2644);
xnor U2819 (N_2819,N_2735,N_2767);
nor U2820 (N_2820,N_2632,N_2760);
nor U2821 (N_2821,N_2677,N_2672);
xor U2822 (N_2822,N_2705,N_2756);
or U2823 (N_2823,N_2667,N_2770);
nor U2824 (N_2824,N_2635,N_2780);
nor U2825 (N_2825,N_2740,N_2714);
and U2826 (N_2826,N_2795,N_2734);
and U2827 (N_2827,N_2685,N_2650);
nand U2828 (N_2828,N_2776,N_2628);
xnor U2829 (N_2829,N_2649,N_2777);
xnor U2830 (N_2830,N_2758,N_2607);
nor U2831 (N_2831,N_2660,N_2779);
nand U2832 (N_2832,N_2645,N_2762);
nand U2833 (N_2833,N_2625,N_2768);
or U2834 (N_2834,N_2702,N_2799);
or U2835 (N_2835,N_2742,N_2726);
or U2836 (N_2836,N_2719,N_2745);
nor U2837 (N_2837,N_2690,N_2652);
or U2838 (N_2838,N_2679,N_2605);
nand U2839 (N_2839,N_2642,N_2609);
or U2840 (N_2840,N_2701,N_2637);
or U2841 (N_2841,N_2669,N_2626);
nand U2842 (N_2842,N_2753,N_2699);
or U2843 (N_2843,N_2771,N_2627);
and U2844 (N_2844,N_2772,N_2790);
nor U2845 (N_2845,N_2670,N_2763);
and U2846 (N_2846,N_2692,N_2653);
xnor U2847 (N_2847,N_2629,N_2739);
nand U2848 (N_2848,N_2788,N_2793);
or U2849 (N_2849,N_2783,N_2687);
or U2850 (N_2850,N_2620,N_2708);
nand U2851 (N_2851,N_2722,N_2666);
and U2852 (N_2852,N_2608,N_2698);
xor U2853 (N_2853,N_2766,N_2729);
nand U2854 (N_2854,N_2683,N_2678);
nor U2855 (N_2855,N_2743,N_2785);
nor U2856 (N_2856,N_2674,N_2731);
or U2857 (N_2857,N_2724,N_2736);
nor U2858 (N_2858,N_2693,N_2673);
nor U2859 (N_2859,N_2711,N_2601);
or U2860 (N_2860,N_2728,N_2775);
nor U2861 (N_2861,N_2786,N_2757);
and U2862 (N_2862,N_2655,N_2707);
nand U2863 (N_2863,N_2633,N_2747);
xor U2864 (N_2864,N_2778,N_2746);
nor U2865 (N_2865,N_2676,N_2664);
or U2866 (N_2866,N_2696,N_2782);
and U2867 (N_2867,N_2717,N_2681);
and U2868 (N_2868,N_2755,N_2744);
nor U2869 (N_2869,N_2631,N_2600);
and U2870 (N_2870,N_2641,N_2616);
xor U2871 (N_2871,N_2796,N_2604);
nand U2872 (N_2872,N_2697,N_2715);
nand U2873 (N_2873,N_2710,N_2704);
nor U2874 (N_2874,N_2709,N_2612);
and U2875 (N_2875,N_2727,N_2621);
and U2876 (N_2876,N_2638,N_2695);
and U2877 (N_2877,N_2737,N_2781);
nand U2878 (N_2878,N_2765,N_2668);
nand U2879 (N_2879,N_2732,N_2774);
nor U2880 (N_2880,N_2738,N_2614);
nand U2881 (N_2881,N_2643,N_2682);
or U2882 (N_2882,N_2640,N_2794);
nor U2883 (N_2883,N_2659,N_2691);
nor U2884 (N_2884,N_2662,N_2675);
nor U2885 (N_2885,N_2630,N_2797);
nand U2886 (N_2886,N_2646,N_2764);
nor U2887 (N_2887,N_2623,N_2720);
xor U2888 (N_2888,N_2789,N_2752);
nor U2889 (N_2889,N_2713,N_2606);
xor U2890 (N_2890,N_2754,N_2748);
nand U2891 (N_2891,N_2751,N_2661);
or U2892 (N_2892,N_2671,N_2686);
nor U2893 (N_2893,N_2665,N_2688);
xnor U2894 (N_2894,N_2716,N_2750);
xnor U2895 (N_2895,N_2611,N_2684);
xnor U2896 (N_2896,N_2723,N_2634);
nor U2897 (N_2897,N_2617,N_2700);
or U2898 (N_2898,N_2651,N_2787);
nand U2899 (N_2899,N_2706,N_2636);
xor U2900 (N_2900,N_2624,N_2757);
or U2901 (N_2901,N_2665,N_2773);
xor U2902 (N_2902,N_2630,N_2617);
or U2903 (N_2903,N_2672,N_2685);
and U2904 (N_2904,N_2783,N_2621);
and U2905 (N_2905,N_2725,N_2741);
nor U2906 (N_2906,N_2676,N_2767);
nand U2907 (N_2907,N_2690,N_2780);
or U2908 (N_2908,N_2797,N_2696);
xor U2909 (N_2909,N_2766,N_2701);
nor U2910 (N_2910,N_2656,N_2712);
nor U2911 (N_2911,N_2678,N_2680);
nor U2912 (N_2912,N_2764,N_2777);
nor U2913 (N_2913,N_2742,N_2681);
or U2914 (N_2914,N_2614,N_2751);
nor U2915 (N_2915,N_2726,N_2678);
or U2916 (N_2916,N_2674,N_2676);
nor U2917 (N_2917,N_2713,N_2696);
or U2918 (N_2918,N_2753,N_2686);
nor U2919 (N_2919,N_2774,N_2746);
nor U2920 (N_2920,N_2620,N_2709);
and U2921 (N_2921,N_2732,N_2711);
or U2922 (N_2922,N_2688,N_2731);
nor U2923 (N_2923,N_2628,N_2668);
or U2924 (N_2924,N_2642,N_2703);
nor U2925 (N_2925,N_2753,N_2657);
xnor U2926 (N_2926,N_2715,N_2616);
or U2927 (N_2927,N_2717,N_2642);
xor U2928 (N_2928,N_2606,N_2665);
or U2929 (N_2929,N_2661,N_2750);
and U2930 (N_2930,N_2760,N_2703);
nand U2931 (N_2931,N_2668,N_2694);
and U2932 (N_2932,N_2607,N_2766);
xnor U2933 (N_2933,N_2731,N_2749);
or U2934 (N_2934,N_2764,N_2761);
nand U2935 (N_2935,N_2665,N_2733);
nor U2936 (N_2936,N_2679,N_2693);
or U2937 (N_2937,N_2749,N_2733);
xnor U2938 (N_2938,N_2634,N_2654);
nor U2939 (N_2939,N_2778,N_2779);
nor U2940 (N_2940,N_2771,N_2763);
nand U2941 (N_2941,N_2616,N_2662);
nand U2942 (N_2942,N_2710,N_2644);
nand U2943 (N_2943,N_2772,N_2753);
nand U2944 (N_2944,N_2696,N_2723);
nand U2945 (N_2945,N_2789,N_2673);
and U2946 (N_2946,N_2710,N_2783);
nand U2947 (N_2947,N_2610,N_2759);
nor U2948 (N_2948,N_2735,N_2677);
or U2949 (N_2949,N_2697,N_2616);
nand U2950 (N_2950,N_2622,N_2730);
or U2951 (N_2951,N_2780,N_2694);
nand U2952 (N_2952,N_2654,N_2793);
and U2953 (N_2953,N_2738,N_2653);
nor U2954 (N_2954,N_2725,N_2700);
or U2955 (N_2955,N_2762,N_2750);
xor U2956 (N_2956,N_2676,N_2677);
and U2957 (N_2957,N_2670,N_2632);
nand U2958 (N_2958,N_2681,N_2650);
nor U2959 (N_2959,N_2615,N_2787);
or U2960 (N_2960,N_2626,N_2709);
or U2961 (N_2961,N_2673,N_2686);
or U2962 (N_2962,N_2787,N_2709);
or U2963 (N_2963,N_2760,N_2697);
nor U2964 (N_2964,N_2629,N_2755);
nand U2965 (N_2965,N_2778,N_2627);
nand U2966 (N_2966,N_2672,N_2790);
and U2967 (N_2967,N_2769,N_2644);
nand U2968 (N_2968,N_2624,N_2622);
and U2969 (N_2969,N_2714,N_2708);
nand U2970 (N_2970,N_2745,N_2784);
and U2971 (N_2971,N_2659,N_2750);
nor U2972 (N_2972,N_2738,N_2705);
or U2973 (N_2973,N_2748,N_2670);
or U2974 (N_2974,N_2652,N_2662);
and U2975 (N_2975,N_2754,N_2701);
nor U2976 (N_2976,N_2690,N_2639);
or U2977 (N_2977,N_2686,N_2730);
or U2978 (N_2978,N_2606,N_2661);
xnor U2979 (N_2979,N_2705,N_2706);
nor U2980 (N_2980,N_2726,N_2754);
and U2981 (N_2981,N_2750,N_2648);
nor U2982 (N_2982,N_2757,N_2766);
xnor U2983 (N_2983,N_2779,N_2714);
nor U2984 (N_2984,N_2620,N_2638);
nor U2985 (N_2985,N_2749,N_2672);
nand U2986 (N_2986,N_2658,N_2718);
or U2987 (N_2987,N_2790,N_2638);
and U2988 (N_2988,N_2745,N_2775);
or U2989 (N_2989,N_2736,N_2645);
and U2990 (N_2990,N_2720,N_2604);
or U2991 (N_2991,N_2744,N_2781);
or U2992 (N_2992,N_2787,N_2699);
nor U2993 (N_2993,N_2673,N_2606);
or U2994 (N_2994,N_2705,N_2604);
and U2995 (N_2995,N_2730,N_2716);
nor U2996 (N_2996,N_2780,N_2639);
nor U2997 (N_2997,N_2719,N_2725);
and U2998 (N_2998,N_2643,N_2740);
and U2999 (N_2999,N_2645,N_2666);
xor U3000 (N_3000,N_2886,N_2844);
or U3001 (N_3001,N_2842,N_2976);
nand U3002 (N_3002,N_2907,N_2869);
xnor U3003 (N_3003,N_2892,N_2988);
or U3004 (N_3004,N_2901,N_2876);
and U3005 (N_3005,N_2898,N_2956);
nor U3006 (N_3006,N_2882,N_2867);
nand U3007 (N_3007,N_2905,N_2964);
nor U3008 (N_3008,N_2958,N_2936);
nand U3009 (N_3009,N_2840,N_2879);
or U3010 (N_3010,N_2877,N_2808);
or U3011 (N_3011,N_2946,N_2817);
or U3012 (N_3012,N_2963,N_2991);
or U3013 (N_3013,N_2922,N_2812);
and U3014 (N_3014,N_2954,N_2806);
or U3015 (N_3015,N_2967,N_2854);
or U3016 (N_3016,N_2980,N_2970);
nand U3017 (N_3017,N_2996,N_2997);
xor U3018 (N_3018,N_2872,N_2871);
or U3019 (N_3019,N_2859,N_2982);
nor U3020 (N_3020,N_2951,N_2983);
nand U3021 (N_3021,N_2813,N_2839);
nand U3022 (N_3022,N_2863,N_2800);
nor U3023 (N_3023,N_2929,N_2934);
or U3024 (N_3024,N_2828,N_2957);
nand U3025 (N_3025,N_2841,N_2866);
nor U3026 (N_3026,N_2889,N_2893);
or U3027 (N_3027,N_2947,N_2857);
nand U3028 (N_3028,N_2993,N_2933);
nor U3029 (N_3029,N_2941,N_2815);
or U3030 (N_3030,N_2825,N_2900);
nand U3031 (N_3031,N_2850,N_2918);
nor U3032 (N_3032,N_2920,N_2969);
nand U3033 (N_3033,N_2870,N_2977);
or U3034 (N_3034,N_2834,N_2875);
nor U3035 (N_3035,N_2913,N_2935);
nand U3036 (N_3036,N_2846,N_2939);
and U3037 (N_3037,N_2955,N_2910);
or U3038 (N_3038,N_2942,N_2968);
or U3039 (N_3039,N_2961,N_2899);
nand U3040 (N_3040,N_2928,N_2971);
and U3041 (N_3041,N_2829,N_2809);
or U3042 (N_3042,N_2973,N_2937);
or U3043 (N_3043,N_2916,N_2902);
and U3044 (N_3044,N_2990,N_2995);
or U3045 (N_3045,N_2949,N_2930);
nor U3046 (N_3046,N_2925,N_2822);
or U3047 (N_3047,N_2862,N_2845);
nor U3048 (N_3048,N_2978,N_2975);
and U3049 (N_3049,N_2805,N_2906);
xnor U3050 (N_3050,N_2852,N_2838);
and U3051 (N_3051,N_2880,N_2874);
or U3052 (N_3052,N_2802,N_2940);
nor U3053 (N_3053,N_2959,N_2856);
nand U3054 (N_3054,N_2887,N_2944);
or U3055 (N_3055,N_2921,N_2826);
nand U3056 (N_3056,N_2924,N_2903);
or U3057 (N_3057,N_2803,N_2895);
or U3058 (N_3058,N_2888,N_2897);
nand U3059 (N_3059,N_2965,N_2833);
or U3060 (N_3060,N_2814,N_2926);
nor U3061 (N_3061,N_2927,N_2865);
nor U3062 (N_3062,N_2851,N_2824);
nand U3063 (N_3063,N_2821,N_2868);
and U3064 (N_3064,N_2966,N_2952);
nand U3065 (N_3065,N_2989,N_2938);
xor U3066 (N_3066,N_2915,N_2909);
nor U3067 (N_3067,N_2807,N_2804);
xor U3068 (N_3068,N_2819,N_2823);
nand U3069 (N_3069,N_2960,N_2855);
nand U3070 (N_3070,N_2932,N_2948);
nand U3071 (N_3071,N_2891,N_2998);
nand U3072 (N_3072,N_2953,N_2883);
and U3073 (N_3073,N_2923,N_2873);
or U3074 (N_3074,N_2885,N_2985);
nor U3075 (N_3075,N_2984,N_2853);
and U3076 (N_3076,N_2950,N_2919);
xor U3077 (N_3077,N_2861,N_2847);
xor U3078 (N_3078,N_2972,N_2999);
nor U3079 (N_3079,N_2890,N_2835);
nor U3080 (N_3080,N_2986,N_2884);
nand U3081 (N_3081,N_2837,N_2811);
nand U3082 (N_3082,N_2943,N_2945);
nor U3083 (N_3083,N_2992,N_2830);
nor U3084 (N_3084,N_2914,N_2908);
or U3085 (N_3085,N_2864,N_2858);
nand U3086 (N_3086,N_2981,N_2979);
or U3087 (N_3087,N_2912,N_2974);
nor U3088 (N_3088,N_2878,N_2848);
nand U3089 (N_3089,N_2816,N_2987);
nor U3090 (N_3090,N_2931,N_2827);
xor U3091 (N_3091,N_2818,N_2881);
nor U3092 (N_3092,N_2904,N_2994);
nand U3093 (N_3093,N_2843,N_2831);
nand U3094 (N_3094,N_2820,N_2832);
and U3095 (N_3095,N_2810,N_2917);
and U3096 (N_3096,N_2962,N_2911);
nand U3097 (N_3097,N_2894,N_2801);
nand U3098 (N_3098,N_2849,N_2896);
nor U3099 (N_3099,N_2836,N_2860);
and U3100 (N_3100,N_2820,N_2828);
nor U3101 (N_3101,N_2953,N_2949);
or U3102 (N_3102,N_2822,N_2848);
nand U3103 (N_3103,N_2931,N_2850);
nand U3104 (N_3104,N_2942,N_2943);
and U3105 (N_3105,N_2901,N_2802);
or U3106 (N_3106,N_2936,N_2982);
and U3107 (N_3107,N_2924,N_2887);
nand U3108 (N_3108,N_2979,N_2886);
and U3109 (N_3109,N_2821,N_2917);
nand U3110 (N_3110,N_2910,N_2833);
nor U3111 (N_3111,N_2962,N_2971);
or U3112 (N_3112,N_2900,N_2915);
nor U3113 (N_3113,N_2922,N_2936);
xor U3114 (N_3114,N_2877,N_2822);
and U3115 (N_3115,N_2996,N_2907);
nor U3116 (N_3116,N_2934,N_2862);
xor U3117 (N_3117,N_2955,N_2947);
nor U3118 (N_3118,N_2944,N_2898);
nand U3119 (N_3119,N_2913,N_2883);
and U3120 (N_3120,N_2846,N_2843);
and U3121 (N_3121,N_2884,N_2915);
nand U3122 (N_3122,N_2846,N_2898);
or U3123 (N_3123,N_2862,N_2832);
or U3124 (N_3124,N_2818,N_2912);
xor U3125 (N_3125,N_2959,N_2864);
xnor U3126 (N_3126,N_2859,N_2988);
or U3127 (N_3127,N_2953,N_2817);
nand U3128 (N_3128,N_2898,N_2857);
nor U3129 (N_3129,N_2934,N_2880);
nand U3130 (N_3130,N_2995,N_2802);
xor U3131 (N_3131,N_2998,N_2947);
or U3132 (N_3132,N_2900,N_2801);
nor U3133 (N_3133,N_2895,N_2842);
nand U3134 (N_3134,N_2804,N_2891);
nand U3135 (N_3135,N_2999,N_2827);
xnor U3136 (N_3136,N_2903,N_2986);
and U3137 (N_3137,N_2915,N_2914);
nor U3138 (N_3138,N_2810,N_2949);
nor U3139 (N_3139,N_2960,N_2816);
and U3140 (N_3140,N_2903,N_2839);
and U3141 (N_3141,N_2965,N_2972);
xnor U3142 (N_3142,N_2906,N_2812);
and U3143 (N_3143,N_2800,N_2963);
nand U3144 (N_3144,N_2903,N_2966);
nor U3145 (N_3145,N_2807,N_2847);
and U3146 (N_3146,N_2854,N_2933);
nand U3147 (N_3147,N_2922,N_2917);
or U3148 (N_3148,N_2816,N_2915);
or U3149 (N_3149,N_2869,N_2885);
nand U3150 (N_3150,N_2906,N_2832);
xnor U3151 (N_3151,N_2915,N_2946);
nor U3152 (N_3152,N_2804,N_2962);
and U3153 (N_3153,N_2949,N_2950);
nor U3154 (N_3154,N_2830,N_2879);
nand U3155 (N_3155,N_2823,N_2972);
or U3156 (N_3156,N_2900,N_2834);
and U3157 (N_3157,N_2883,N_2946);
and U3158 (N_3158,N_2951,N_2883);
or U3159 (N_3159,N_2967,N_2871);
and U3160 (N_3160,N_2953,N_2943);
and U3161 (N_3161,N_2830,N_2882);
nor U3162 (N_3162,N_2896,N_2944);
nor U3163 (N_3163,N_2826,N_2963);
nor U3164 (N_3164,N_2829,N_2828);
or U3165 (N_3165,N_2813,N_2898);
or U3166 (N_3166,N_2908,N_2959);
xor U3167 (N_3167,N_2874,N_2901);
and U3168 (N_3168,N_2984,N_2863);
and U3169 (N_3169,N_2822,N_2916);
xor U3170 (N_3170,N_2951,N_2908);
and U3171 (N_3171,N_2947,N_2985);
nand U3172 (N_3172,N_2940,N_2934);
nand U3173 (N_3173,N_2919,N_2810);
nor U3174 (N_3174,N_2988,N_2875);
nand U3175 (N_3175,N_2831,N_2816);
and U3176 (N_3176,N_2911,N_2917);
nor U3177 (N_3177,N_2811,N_2843);
xor U3178 (N_3178,N_2954,N_2996);
and U3179 (N_3179,N_2841,N_2952);
nor U3180 (N_3180,N_2890,N_2910);
nand U3181 (N_3181,N_2978,N_2993);
or U3182 (N_3182,N_2879,N_2872);
nor U3183 (N_3183,N_2966,N_2801);
xor U3184 (N_3184,N_2834,N_2862);
and U3185 (N_3185,N_2849,N_2826);
and U3186 (N_3186,N_2816,N_2935);
or U3187 (N_3187,N_2816,N_2893);
xnor U3188 (N_3188,N_2816,N_2813);
nand U3189 (N_3189,N_2835,N_2951);
nor U3190 (N_3190,N_2928,N_2907);
or U3191 (N_3191,N_2922,N_2860);
nand U3192 (N_3192,N_2852,N_2989);
nor U3193 (N_3193,N_2888,N_2981);
and U3194 (N_3194,N_2974,N_2919);
and U3195 (N_3195,N_2890,N_2940);
and U3196 (N_3196,N_2979,N_2927);
nor U3197 (N_3197,N_2865,N_2803);
and U3198 (N_3198,N_2944,N_2967);
nand U3199 (N_3199,N_2851,N_2951);
nand U3200 (N_3200,N_3093,N_3054);
or U3201 (N_3201,N_3173,N_3053);
nand U3202 (N_3202,N_3117,N_3094);
or U3203 (N_3203,N_3095,N_3147);
and U3204 (N_3204,N_3171,N_3156);
or U3205 (N_3205,N_3049,N_3166);
nand U3206 (N_3206,N_3159,N_3005);
xor U3207 (N_3207,N_3015,N_3006);
or U3208 (N_3208,N_3177,N_3046);
or U3209 (N_3209,N_3103,N_3178);
xnor U3210 (N_3210,N_3089,N_3175);
nor U3211 (N_3211,N_3131,N_3140);
nor U3212 (N_3212,N_3031,N_3190);
xnor U3213 (N_3213,N_3188,N_3198);
nor U3214 (N_3214,N_3116,N_3029);
nand U3215 (N_3215,N_3162,N_3059);
or U3216 (N_3216,N_3084,N_3043);
xor U3217 (N_3217,N_3082,N_3061);
nand U3218 (N_3218,N_3063,N_3060);
and U3219 (N_3219,N_3121,N_3098);
and U3220 (N_3220,N_3144,N_3143);
nand U3221 (N_3221,N_3057,N_3096);
or U3222 (N_3222,N_3042,N_3020);
and U3223 (N_3223,N_3108,N_3045);
or U3224 (N_3224,N_3150,N_3165);
nor U3225 (N_3225,N_3148,N_3114);
nor U3226 (N_3226,N_3182,N_3126);
nand U3227 (N_3227,N_3127,N_3193);
or U3228 (N_3228,N_3081,N_3124);
xnor U3229 (N_3229,N_3163,N_3141);
nor U3230 (N_3230,N_3068,N_3118);
nor U3231 (N_3231,N_3058,N_3047);
nand U3232 (N_3232,N_3184,N_3052);
and U3233 (N_3233,N_3039,N_3038);
xor U3234 (N_3234,N_3123,N_3000);
or U3235 (N_3235,N_3066,N_3050);
and U3236 (N_3236,N_3115,N_3090);
or U3237 (N_3237,N_3062,N_3160);
nor U3238 (N_3238,N_3111,N_3037);
and U3239 (N_3239,N_3197,N_3021);
nor U3240 (N_3240,N_3113,N_3040);
and U3241 (N_3241,N_3137,N_3027);
or U3242 (N_3242,N_3099,N_3088);
nor U3243 (N_3243,N_3036,N_3026);
and U3244 (N_3244,N_3102,N_3086);
or U3245 (N_3245,N_3109,N_3125);
and U3246 (N_3246,N_3051,N_3138);
nor U3247 (N_3247,N_3130,N_3078);
and U3248 (N_3248,N_3009,N_3164);
or U3249 (N_3249,N_3065,N_3191);
nand U3250 (N_3250,N_3196,N_3072);
and U3251 (N_3251,N_3136,N_3167);
nand U3252 (N_3252,N_3157,N_3028);
or U3253 (N_3253,N_3183,N_3018);
nand U3254 (N_3254,N_3187,N_3192);
xnor U3255 (N_3255,N_3002,N_3034);
xnor U3256 (N_3256,N_3149,N_3012);
or U3257 (N_3257,N_3076,N_3186);
nor U3258 (N_3258,N_3080,N_3169);
nand U3259 (N_3259,N_3110,N_3101);
nor U3260 (N_3260,N_3041,N_3001);
nor U3261 (N_3261,N_3142,N_3120);
or U3262 (N_3262,N_3195,N_3172);
and U3263 (N_3263,N_3100,N_3135);
nand U3264 (N_3264,N_3168,N_3181);
and U3265 (N_3265,N_3176,N_3032);
or U3266 (N_3266,N_3154,N_3155);
and U3267 (N_3267,N_3107,N_3074);
nand U3268 (N_3268,N_3122,N_3070);
nand U3269 (N_3269,N_3067,N_3161);
nor U3270 (N_3270,N_3055,N_3016);
nand U3271 (N_3271,N_3199,N_3129);
nand U3272 (N_3272,N_3139,N_3087);
nand U3273 (N_3273,N_3189,N_3019);
nand U3274 (N_3274,N_3025,N_3030);
nor U3275 (N_3275,N_3073,N_3153);
nand U3276 (N_3276,N_3022,N_3075);
nand U3277 (N_3277,N_3151,N_3152);
and U3278 (N_3278,N_3092,N_3105);
nor U3279 (N_3279,N_3069,N_3097);
or U3280 (N_3280,N_3011,N_3180);
nand U3281 (N_3281,N_3014,N_3010);
and U3282 (N_3282,N_3134,N_3003);
or U3283 (N_3283,N_3106,N_3004);
nor U3284 (N_3284,N_3146,N_3071);
nor U3285 (N_3285,N_3083,N_3133);
nor U3286 (N_3286,N_3185,N_3013);
nand U3287 (N_3287,N_3132,N_3119);
and U3288 (N_3288,N_3179,N_3079);
nand U3289 (N_3289,N_3085,N_3158);
and U3290 (N_3290,N_3104,N_3194);
nand U3291 (N_3291,N_3017,N_3145);
and U3292 (N_3292,N_3091,N_3024);
nand U3293 (N_3293,N_3048,N_3035);
and U3294 (N_3294,N_3170,N_3008);
nor U3295 (N_3295,N_3112,N_3056);
nand U3296 (N_3296,N_3077,N_3064);
and U3297 (N_3297,N_3007,N_3128);
and U3298 (N_3298,N_3023,N_3033);
and U3299 (N_3299,N_3044,N_3174);
or U3300 (N_3300,N_3101,N_3175);
xor U3301 (N_3301,N_3007,N_3010);
and U3302 (N_3302,N_3114,N_3119);
nand U3303 (N_3303,N_3031,N_3010);
nor U3304 (N_3304,N_3124,N_3188);
nor U3305 (N_3305,N_3088,N_3159);
or U3306 (N_3306,N_3140,N_3172);
nor U3307 (N_3307,N_3053,N_3085);
or U3308 (N_3308,N_3088,N_3151);
nor U3309 (N_3309,N_3046,N_3019);
or U3310 (N_3310,N_3150,N_3011);
nor U3311 (N_3311,N_3020,N_3190);
or U3312 (N_3312,N_3069,N_3159);
or U3313 (N_3313,N_3174,N_3069);
or U3314 (N_3314,N_3079,N_3070);
nand U3315 (N_3315,N_3079,N_3143);
or U3316 (N_3316,N_3179,N_3043);
nor U3317 (N_3317,N_3031,N_3133);
xor U3318 (N_3318,N_3114,N_3166);
nor U3319 (N_3319,N_3032,N_3130);
nand U3320 (N_3320,N_3020,N_3003);
nor U3321 (N_3321,N_3175,N_3050);
nand U3322 (N_3322,N_3096,N_3086);
nand U3323 (N_3323,N_3033,N_3018);
or U3324 (N_3324,N_3050,N_3194);
nand U3325 (N_3325,N_3173,N_3092);
nand U3326 (N_3326,N_3126,N_3061);
nand U3327 (N_3327,N_3157,N_3193);
nand U3328 (N_3328,N_3153,N_3094);
nor U3329 (N_3329,N_3107,N_3009);
nand U3330 (N_3330,N_3196,N_3193);
or U3331 (N_3331,N_3193,N_3077);
nor U3332 (N_3332,N_3027,N_3161);
nand U3333 (N_3333,N_3082,N_3044);
xnor U3334 (N_3334,N_3040,N_3177);
and U3335 (N_3335,N_3174,N_3179);
or U3336 (N_3336,N_3016,N_3028);
and U3337 (N_3337,N_3171,N_3168);
and U3338 (N_3338,N_3127,N_3083);
and U3339 (N_3339,N_3120,N_3091);
and U3340 (N_3340,N_3112,N_3065);
nor U3341 (N_3341,N_3107,N_3174);
or U3342 (N_3342,N_3178,N_3172);
or U3343 (N_3343,N_3105,N_3024);
or U3344 (N_3344,N_3113,N_3181);
nand U3345 (N_3345,N_3003,N_3034);
nor U3346 (N_3346,N_3130,N_3046);
or U3347 (N_3347,N_3157,N_3062);
nand U3348 (N_3348,N_3026,N_3135);
and U3349 (N_3349,N_3141,N_3144);
or U3350 (N_3350,N_3051,N_3090);
and U3351 (N_3351,N_3179,N_3120);
nor U3352 (N_3352,N_3166,N_3028);
or U3353 (N_3353,N_3153,N_3012);
xnor U3354 (N_3354,N_3099,N_3062);
nand U3355 (N_3355,N_3065,N_3109);
nor U3356 (N_3356,N_3177,N_3174);
nand U3357 (N_3357,N_3193,N_3106);
or U3358 (N_3358,N_3053,N_3062);
nand U3359 (N_3359,N_3149,N_3165);
and U3360 (N_3360,N_3104,N_3161);
and U3361 (N_3361,N_3155,N_3140);
nand U3362 (N_3362,N_3190,N_3060);
and U3363 (N_3363,N_3021,N_3100);
or U3364 (N_3364,N_3158,N_3097);
and U3365 (N_3365,N_3023,N_3062);
nor U3366 (N_3366,N_3038,N_3054);
nor U3367 (N_3367,N_3159,N_3184);
or U3368 (N_3368,N_3141,N_3067);
nor U3369 (N_3369,N_3155,N_3027);
nor U3370 (N_3370,N_3136,N_3005);
nand U3371 (N_3371,N_3164,N_3183);
nor U3372 (N_3372,N_3106,N_3157);
and U3373 (N_3373,N_3190,N_3172);
nor U3374 (N_3374,N_3051,N_3137);
or U3375 (N_3375,N_3119,N_3074);
nor U3376 (N_3376,N_3170,N_3194);
or U3377 (N_3377,N_3035,N_3144);
nand U3378 (N_3378,N_3040,N_3004);
or U3379 (N_3379,N_3163,N_3137);
nand U3380 (N_3380,N_3131,N_3101);
nor U3381 (N_3381,N_3000,N_3032);
or U3382 (N_3382,N_3093,N_3015);
or U3383 (N_3383,N_3062,N_3003);
and U3384 (N_3384,N_3035,N_3141);
xor U3385 (N_3385,N_3102,N_3177);
or U3386 (N_3386,N_3000,N_3079);
nor U3387 (N_3387,N_3026,N_3166);
and U3388 (N_3388,N_3037,N_3056);
xnor U3389 (N_3389,N_3046,N_3173);
or U3390 (N_3390,N_3065,N_3133);
nand U3391 (N_3391,N_3116,N_3178);
nor U3392 (N_3392,N_3042,N_3015);
nand U3393 (N_3393,N_3189,N_3081);
or U3394 (N_3394,N_3079,N_3067);
and U3395 (N_3395,N_3145,N_3181);
nor U3396 (N_3396,N_3057,N_3163);
xor U3397 (N_3397,N_3087,N_3179);
xnor U3398 (N_3398,N_3021,N_3162);
and U3399 (N_3399,N_3110,N_3052);
nand U3400 (N_3400,N_3276,N_3329);
nor U3401 (N_3401,N_3255,N_3335);
nor U3402 (N_3402,N_3399,N_3221);
xor U3403 (N_3403,N_3380,N_3287);
or U3404 (N_3404,N_3397,N_3367);
nor U3405 (N_3405,N_3262,N_3315);
or U3406 (N_3406,N_3272,N_3258);
nor U3407 (N_3407,N_3207,N_3344);
and U3408 (N_3408,N_3271,N_3230);
or U3409 (N_3409,N_3245,N_3268);
nor U3410 (N_3410,N_3267,N_3259);
and U3411 (N_3411,N_3396,N_3390);
nand U3412 (N_3412,N_3204,N_3328);
xnor U3413 (N_3413,N_3235,N_3202);
or U3414 (N_3414,N_3269,N_3281);
nand U3415 (N_3415,N_3282,N_3356);
nand U3416 (N_3416,N_3360,N_3353);
or U3417 (N_3417,N_3270,N_3311);
and U3418 (N_3418,N_3332,N_3351);
nand U3419 (N_3419,N_3296,N_3289);
and U3420 (N_3420,N_3298,N_3244);
or U3421 (N_3421,N_3317,N_3278);
nand U3422 (N_3422,N_3275,N_3265);
xnor U3423 (N_3423,N_3386,N_3212);
nor U3424 (N_3424,N_3337,N_3384);
nand U3425 (N_3425,N_3295,N_3243);
and U3426 (N_3426,N_3261,N_3274);
and U3427 (N_3427,N_3201,N_3361);
and U3428 (N_3428,N_3218,N_3293);
or U3429 (N_3429,N_3266,N_3374);
nor U3430 (N_3430,N_3302,N_3205);
and U3431 (N_3431,N_3220,N_3214);
xor U3432 (N_3432,N_3283,N_3200);
nand U3433 (N_3433,N_3264,N_3333);
xnor U3434 (N_3434,N_3246,N_3294);
nand U3435 (N_3435,N_3217,N_3321);
nor U3436 (N_3436,N_3393,N_3359);
nand U3437 (N_3437,N_3288,N_3395);
or U3438 (N_3438,N_3383,N_3210);
nor U3439 (N_3439,N_3285,N_3290);
nor U3440 (N_3440,N_3372,N_3239);
or U3441 (N_3441,N_3376,N_3325);
nand U3442 (N_3442,N_3224,N_3240);
or U3443 (N_3443,N_3257,N_3382);
and U3444 (N_3444,N_3316,N_3222);
and U3445 (N_3445,N_3352,N_3385);
or U3446 (N_3446,N_3307,N_3377);
nand U3447 (N_3447,N_3324,N_3358);
or U3448 (N_3448,N_3301,N_3343);
or U3449 (N_3449,N_3368,N_3357);
and U3450 (N_3450,N_3347,N_3263);
or U3451 (N_3451,N_3211,N_3319);
nand U3452 (N_3452,N_3330,N_3355);
nand U3453 (N_3453,N_3338,N_3284);
or U3454 (N_3454,N_3387,N_3234);
xnor U3455 (N_3455,N_3241,N_3379);
nand U3456 (N_3456,N_3320,N_3369);
nor U3457 (N_3457,N_3392,N_3312);
and U3458 (N_3458,N_3251,N_3326);
nand U3459 (N_3459,N_3232,N_3350);
nand U3460 (N_3460,N_3226,N_3366);
nor U3461 (N_3461,N_3308,N_3254);
or U3462 (N_3462,N_3306,N_3370);
nor U3463 (N_3463,N_3252,N_3389);
nand U3464 (N_3464,N_3236,N_3229);
nand U3465 (N_3465,N_3247,N_3375);
and U3466 (N_3466,N_3323,N_3314);
and U3467 (N_3467,N_3206,N_3250);
nand U3468 (N_3468,N_3209,N_3341);
nor U3469 (N_3469,N_3345,N_3394);
nand U3470 (N_3470,N_3228,N_3381);
and U3471 (N_3471,N_3363,N_3362);
nand U3472 (N_3472,N_3260,N_3331);
nor U3473 (N_3473,N_3223,N_3208);
and U3474 (N_3474,N_3348,N_3256);
nand U3475 (N_3475,N_3349,N_3340);
nor U3476 (N_3476,N_3215,N_3248);
and U3477 (N_3477,N_3277,N_3310);
nor U3478 (N_3478,N_3322,N_3231);
and U3479 (N_3479,N_3373,N_3354);
or U3480 (N_3480,N_3342,N_3297);
nor U3481 (N_3481,N_3238,N_3305);
nor U3482 (N_3482,N_3313,N_3391);
or U3483 (N_3483,N_3249,N_3334);
xnor U3484 (N_3484,N_3388,N_3216);
or U3485 (N_3485,N_3327,N_3291);
or U3486 (N_3486,N_3365,N_3304);
xor U3487 (N_3487,N_3346,N_3292);
nand U3488 (N_3488,N_3279,N_3398);
xor U3489 (N_3489,N_3300,N_3227);
nand U3490 (N_3490,N_3303,N_3309);
or U3491 (N_3491,N_3339,N_3253);
nor U3492 (N_3492,N_3225,N_3273);
nor U3493 (N_3493,N_3336,N_3203);
nand U3494 (N_3494,N_3237,N_3378);
nor U3495 (N_3495,N_3299,N_3242);
and U3496 (N_3496,N_3371,N_3364);
or U3497 (N_3497,N_3286,N_3213);
and U3498 (N_3498,N_3233,N_3280);
or U3499 (N_3499,N_3318,N_3219);
nand U3500 (N_3500,N_3265,N_3303);
xnor U3501 (N_3501,N_3392,N_3334);
nand U3502 (N_3502,N_3243,N_3207);
nor U3503 (N_3503,N_3394,N_3229);
xor U3504 (N_3504,N_3394,N_3280);
nand U3505 (N_3505,N_3399,N_3241);
nor U3506 (N_3506,N_3310,N_3218);
or U3507 (N_3507,N_3355,N_3398);
and U3508 (N_3508,N_3263,N_3287);
or U3509 (N_3509,N_3215,N_3345);
nand U3510 (N_3510,N_3332,N_3337);
nand U3511 (N_3511,N_3369,N_3206);
nor U3512 (N_3512,N_3246,N_3229);
or U3513 (N_3513,N_3355,N_3258);
or U3514 (N_3514,N_3396,N_3357);
nand U3515 (N_3515,N_3203,N_3308);
nand U3516 (N_3516,N_3236,N_3306);
and U3517 (N_3517,N_3285,N_3369);
or U3518 (N_3518,N_3278,N_3250);
nand U3519 (N_3519,N_3399,N_3254);
xnor U3520 (N_3520,N_3286,N_3262);
and U3521 (N_3521,N_3274,N_3384);
nor U3522 (N_3522,N_3244,N_3312);
nand U3523 (N_3523,N_3288,N_3347);
and U3524 (N_3524,N_3354,N_3347);
or U3525 (N_3525,N_3284,N_3354);
xor U3526 (N_3526,N_3301,N_3235);
nor U3527 (N_3527,N_3365,N_3302);
nor U3528 (N_3528,N_3243,N_3341);
or U3529 (N_3529,N_3250,N_3385);
xor U3530 (N_3530,N_3237,N_3301);
nand U3531 (N_3531,N_3387,N_3383);
and U3532 (N_3532,N_3219,N_3261);
xor U3533 (N_3533,N_3339,N_3343);
xor U3534 (N_3534,N_3239,N_3235);
nor U3535 (N_3535,N_3394,N_3270);
nand U3536 (N_3536,N_3205,N_3376);
nand U3537 (N_3537,N_3219,N_3383);
or U3538 (N_3538,N_3298,N_3346);
nor U3539 (N_3539,N_3298,N_3311);
or U3540 (N_3540,N_3218,N_3281);
nor U3541 (N_3541,N_3238,N_3296);
and U3542 (N_3542,N_3279,N_3235);
xnor U3543 (N_3543,N_3262,N_3260);
or U3544 (N_3544,N_3227,N_3310);
or U3545 (N_3545,N_3374,N_3285);
xnor U3546 (N_3546,N_3306,N_3365);
and U3547 (N_3547,N_3202,N_3317);
xnor U3548 (N_3548,N_3202,N_3201);
or U3549 (N_3549,N_3320,N_3269);
or U3550 (N_3550,N_3218,N_3260);
xor U3551 (N_3551,N_3340,N_3372);
nor U3552 (N_3552,N_3257,N_3256);
and U3553 (N_3553,N_3379,N_3280);
or U3554 (N_3554,N_3363,N_3214);
and U3555 (N_3555,N_3236,N_3379);
or U3556 (N_3556,N_3347,N_3242);
and U3557 (N_3557,N_3399,N_3333);
nor U3558 (N_3558,N_3341,N_3333);
or U3559 (N_3559,N_3284,N_3392);
nor U3560 (N_3560,N_3271,N_3288);
nor U3561 (N_3561,N_3244,N_3236);
nand U3562 (N_3562,N_3347,N_3252);
or U3563 (N_3563,N_3214,N_3372);
and U3564 (N_3564,N_3265,N_3210);
or U3565 (N_3565,N_3358,N_3305);
nor U3566 (N_3566,N_3238,N_3381);
xnor U3567 (N_3567,N_3245,N_3327);
nor U3568 (N_3568,N_3280,N_3289);
nand U3569 (N_3569,N_3233,N_3391);
nand U3570 (N_3570,N_3204,N_3255);
nor U3571 (N_3571,N_3230,N_3375);
nor U3572 (N_3572,N_3376,N_3264);
and U3573 (N_3573,N_3200,N_3212);
nand U3574 (N_3574,N_3255,N_3262);
nand U3575 (N_3575,N_3223,N_3333);
nor U3576 (N_3576,N_3398,N_3345);
nand U3577 (N_3577,N_3314,N_3378);
nor U3578 (N_3578,N_3332,N_3348);
or U3579 (N_3579,N_3226,N_3235);
nor U3580 (N_3580,N_3264,N_3391);
xor U3581 (N_3581,N_3391,N_3339);
nand U3582 (N_3582,N_3333,N_3385);
nor U3583 (N_3583,N_3222,N_3259);
xor U3584 (N_3584,N_3331,N_3240);
or U3585 (N_3585,N_3382,N_3320);
xor U3586 (N_3586,N_3232,N_3356);
and U3587 (N_3587,N_3370,N_3234);
nand U3588 (N_3588,N_3331,N_3203);
or U3589 (N_3589,N_3311,N_3233);
and U3590 (N_3590,N_3363,N_3206);
nor U3591 (N_3591,N_3341,N_3305);
or U3592 (N_3592,N_3205,N_3271);
and U3593 (N_3593,N_3310,N_3246);
nand U3594 (N_3594,N_3264,N_3317);
nand U3595 (N_3595,N_3221,N_3378);
nor U3596 (N_3596,N_3304,N_3214);
nor U3597 (N_3597,N_3394,N_3240);
and U3598 (N_3598,N_3224,N_3309);
or U3599 (N_3599,N_3216,N_3340);
nor U3600 (N_3600,N_3536,N_3489);
or U3601 (N_3601,N_3487,N_3473);
or U3602 (N_3602,N_3406,N_3565);
and U3603 (N_3603,N_3538,N_3527);
or U3604 (N_3604,N_3590,N_3506);
or U3605 (N_3605,N_3583,N_3559);
nor U3606 (N_3606,N_3470,N_3436);
nand U3607 (N_3607,N_3548,N_3566);
nand U3608 (N_3608,N_3481,N_3493);
and U3609 (N_3609,N_3488,N_3495);
or U3610 (N_3610,N_3555,N_3550);
nor U3611 (N_3611,N_3432,N_3558);
and U3612 (N_3612,N_3502,N_3435);
and U3613 (N_3613,N_3476,N_3459);
nor U3614 (N_3614,N_3569,N_3522);
nor U3615 (N_3615,N_3401,N_3517);
or U3616 (N_3616,N_3561,N_3410);
xnor U3617 (N_3617,N_3464,N_3492);
nand U3618 (N_3618,N_3530,N_3532);
nand U3619 (N_3619,N_3462,N_3425);
nand U3620 (N_3620,N_3510,N_3579);
or U3621 (N_3621,N_3466,N_3599);
and U3622 (N_3622,N_3490,N_3444);
nand U3623 (N_3623,N_3526,N_3403);
nor U3624 (N_3624,N_3520,N_3455);
xnor U3625 (N_3625,N_3430,N_3501);
nand U3626 (N_3626,N_3441,N_3428);
and U3627 (N_3627,N_3570,N_3563);
nand U3628 (N_3628,N_3531,N_3547);
xnor U3629 (N_3629,N_3414,N_3443);
and U3630 (N_3630,N_3521,N_3500);
or U3631 (N_3631,N_3504,N_3486);
xor U3632 (N_3632,N_3529,N_3424);
nor U3633 (N_3633,N_3408,N_3453);
nor U3634 (N_3634,N_3440,N_3465);
nand U3635 (N_3635,N_3451,N_3445);
and U3636 (N_3636,N_3588,N_3475);
nand U3637 (N_3637,N_3427,N_3528);
nand U3638 (N_3638,N_3582,N_3420);
nand U3639 (N_3639,N_3519,N_3472);
nand U3640 (N_3640,N_3560,N_3554);
nor U3641 (N_3641,N_3499,N_3498);
and U3642 (N_3642,N_3595,N_3568);
and U3643 (N_3643,N_3457,N_3479);
or U3644 (N_3644,N_3523,N_3442);
and U3645 (N_3645,N_3483,N_3544);
nand U3646 (N_3646,N_3556,N_3447);
nor U3647 (N_3647,N_3407,N_3581);
xnor U3648 (N_3648,N_3450,N_3494);
xor U3649 (N_3649,N_3446,N_3412);
nor U3650 (N_3650,N_3460,N_3598);
xor U3651 (N_3651,N_3404,N_3512);
nand U3652 (N_3652,N_3577,N_3458);
xor U3653 (N_3653,N_3480,N_3478);
nand U3654 (N_3654,N_3454,N_3484);
and U3655 (N_3655,N_3596,N_3589);
nand U3656 (N_3656,N_3497,N_3575);
or U3657 (N_3657,N_3542,N_3433);
and U3658 (N_3658,N_3580,N_3584);
or U3659 (N_3659,N_3594,N_3423);
and U3660 (N_3660,N_3535,N_3562);
xnor U3661 (N_3661,N_3564,N_3503);
and U3662 (N_3662,N_3549,N_3552);
nor U3663 (N_3663,N_3576,N_3400);
and U3664 (N_3664,N_3413,N_3591);
or U3665 (N_3665,N_3438,N_3571);
and U3666 (N_3666,N_3463,N_3417);
nand U3667 (N_3667,N_3448,N_3507);
or U3668 (N_3668,N_3518,N_3511);
nand U3669 (N_3669,N_3482,N_3468);
nand U3670 (N_3670,N_3509,N_3515);
nand U3671 (N_3671,N_3471,N_3553);
or U3672 (N_3672,N_3461,N_3592);
or U3673 (N_3673,N_3437,N_3452);
xor U3674 (N_3674,N_3402,N_3429);
or U3675 (N_3675,N_3467,N_3409);
nand U3676 (N_3676,N_3534,N_3474);
and U3677 (N_3677,N_3586,N_3593);
nor U3678 (N_3678,N_3533,N_3469);
nor U3679 (N_3679,N_3524,N_3419);
nor U3680 (N_3680,N_3587,N_3541);
and U3681 (N_3681,N_3567,N_3426);
and U3682 (N_3682,N_3551,N_3439);
or U3683 (N_3683,N_3514,N_3411);
nand U3684 (N_3684,N_3572,N_3422);
nor U3685 (N_3685,N_3496,N_3421);
or U3686 (N_3686,N_3578,N_3456);
or U3687 (N_3687,N_3585,N_3537);
nand U3688 (N_3688,N_3477,N_3513);
and U3689 (N_3689,N_3573,N_3557);
xnor U3690 (N_3690,N_3516,N_3574);
nor U3691 (N_3691,N_3449,N_3545);
or U3692 (N_3692,N_3508,N_3597);
and U3693 (N_3693,N_3485,N_3415);
xnor U3694 (N_3694,N_3431,N_3525);
nand U3695 (N_3695,N_3418,N_3540);
or U3696 (N_3696,N_3491,N_3434);
nand U3697 (N_3697,N_3405,N_3543);
xor U3698 (N_3698,N_3539,N_3416);
xor U3699 (N_3699,N_3546,N_3505);
nor U3700 (N_3700,N_3459,N_3566);
nor U3701 (N_3701,N_3459,N_3473);
and U3702 (N_3702,N_3539,N_3520);
and U3703 (N_3703,N_3441,N_3596);
nor U3704 (N_3704,N_3460,N_3489);
nand U3705 (N_3705,N_3545,N_3531);
and U3706 (N_3706,N_3461,N_3439);
nand U3707 (N_3707,N_3577,N_3454);
and U3708 (N_3708,N_3517,N_3469);
xor U3709 (N_3709,N_3494,N_3578);
nor U3710 (N_3710,N_3586,N_3521);
and U3711 (N_3711,N_3418,N_3474);
xnor U3712 (N_3712,N_3559,N_3454);
and U3713 (N_3713,N_3444,N_3584);
xor U3714 (N_3714,N_3426,N_3449);
nand U3715 (N_3715,N_3513,N_3553);
and U3716 (N_3716,N_3584,N_3512);
nor U3717 (N_3717,N_3508,N_3404);
nand U3718 (N_3718,N_3464,N_3476);
nor U3719 (N_3719,N_3443,N_3467);
and U3720 (N_3720,N_3520,N_3581);
xor U3721 (N_3721,N_3494,N_3473);
nand U3722 (N_3722,N_3476,N_3577);
and U3723 (N_3723,N_3560,N_3454);
nand U3724 (N_3724,N_3510,N_3599);
nand U3725 (N_3725,N_3548,N_3545);
nand U3726 (N_3726,N_3410,N_3469);
and U3727 (N_3727,N_3460,N_3546);
nand U3728 (N_3728,N_3458,N_3428);
and U3729 (N_3729,N_3557,N_3448);
and U3730 (N_3730,N_3503,N_3501);
xnor U3731 (N_3731,N_3430,N_3419);
nor U3732 (N_3732,N_3579,N_3437);
or U3733 (N_3733,N_3544,N_3503);
nor U3734 (N_3734,N_3568,N_3428);
or U3735 (N_3735,N_3496,N_3411);
nand U3736 (N_3736,N_3541,N_3494);
or U3737 (N_3737,N_3434,N_3525);
or U3738 (N_3738,N_3559,N_3413);
nor U3739 (N_3739,N_3448,N_3431);
and U3740 (N_3740,N_3557,N_3555);
or U3741 (N_3741,N_3528,N_3489);
xor U3742 (N_3742,N_3524,N_3497);
nor U3743 (N_3743,N_3454,N_3506);
nand U3744 (N_3744,N_3481,N_3438);
or U3745 (N_3745,N_3474,N_3475);
and U3746 (N_3746,N_3578,N_3583);
or U3747 (N_3747,N_3525,N_3493);
and U3748 (N_3748,N_3561,N_3575);
nor U3749 (N_3749,N_3418,N_3404);
nand U3750 (N_3750,N_3520,N_3430);
and U3751 (N_3751,N_3520,N_3409);
or U3752 (N_3752,N_3565,N_3537);
nand U3753 (N_3753,N_3497,N_3429);
nor U3754 (N_3754,N_3476,N_3454);
or U3755 (N_3755,N_3448,N_3578);
or U3756 (N_3756,N_3541,N_3418);
nand U3757 (N_3757,N_3556,N_3471);
nor U3758 (N_3758,N_3578,N_3479);
nand U3759 (N_3759,N_3448,N_3465);
and U3760 (N_3760,N_3477,N_3464);
nor U3761 (N_3761,N_3404,N_3449);
nor U3762 (N_3762,N_3405,N_3547);
and U3763 (N_3763,N_3418,N_3499);
and U3764 (N_3764,N_3413,N_3406);
and U3765 (N_3765,N_3550,N_3519);
nor U3766 (N_3766,N_3510,N_3464);
nor U3767 (N_3767,N_3581,N_3503);
nor U3768 (N_3768,N_3446,N_3567);
nand U3769 (N_3769,N_3596,N_3506);
and U3770 (N_3770,N_3417,N_3474);
or U3771 (N_3771,N_3462,N_3529);
or U3772 (N_3772,N_3438,N_3553);
xor U3773 (N_3773,N_3585,N_3583);
and U3774 (N_3774,N_3450,N_3446);
and U3775 (N_3775,N_3479,N_3514);
or U3776 (N_3776,N_3489,N_3527);
nand U3777 (N_3777,N_3443,N_3516);
and U3778 (N_3778,N_3446,N_3541);
and U3779 (N_3779,N_3447,N_3468);
nor U3780 (N_3780,N_3556,N_3403);
nand U3781 (N_3781,N_3574,N_3596);
or U3782 (N_3782,N_3425,N_3429);
xnor U3783 (N_3783,N_3545,N_3572);
and U3784 (N_3784,N_3527,N_3450);
and U3785 (N_3785,N_3460,N_3448);
nor U3786 (N_3786,N_3497,N_3452);
nor U3787 (N_3787,N_3560,N_3599);
nand U3788 (N_3788,N_3556,N_3585);
and U3789 (N_3789,N_3557,N_3584);
nand U3790 (N_3790,N_3410,N_3412);
nor U3791 (N_3791,N_3536,N_3584);
nand U3792 (N_3792,N_3574,N_3501);
nor U3793 (N_3793,N_3440,N_3583);
and U3794 (N_3794,N_3528,N_3567);
or U3795 (N_3795,N_3591,N_3579);
nor U3796 (N_3796,N_3486,N_3477);
nand U3797 (N_3797,N_3492,N_3519);
or U3798 (N_3798,N_3481,N_3536);
and U3799 (N_3799,N_3425,N_3469);
nor U3800 (N_3800,N_3627,N_3630);
and U3801 (N_3801,N_3777,N_3704);
nor U3802 (N_3802,N_3631,N_3647);
nor U3803 (N_3803,N_3635,N_3727);
nor U3804 (N_3804,N_3600,N_3626);
nand U3805 (N_3805,N_3649,N_3609);
nand U3806 (N_3806,N_3786,N_3705);
or U3807 (N_3807,N_3641,N_3767);
nor U3808 (N_3808,N_3654,N_3689);
and U3809 (N_3809,N_3618,N_3646);
and U3810 (N_3810,N_3703,N_3717);
nand U3811 (N_3811,N_3744,N_3690);
nor U3812 (N_3812,N_3745,N_3708);
and U3813 (N_3813,N_3610,N_3663);
or U3814 (N_3814,N_3773,N_3613);
nand U3815 (N_3815,N_3776,N_3664);
or U3816 (N_3816,N_3772,N_3611);
nor U3817 (N_3817,N_3685,N_3707);
nand U3818 (N_3818,N_3608,N_3795);
or U3819 (N_3819,N_3791,N_3742);
nand U3820 (N_3820,N_3665,N_3692);
and U3821 (N_3821,N_3743,N_3667);
and U3822 (N_3822,N_3668,N_3737);
and U3823 (N_3823,N_3721,N_3770);
nor U3824 (N_3824,N_3679,N_3746);
or U3825 (N_3825,N_3758,N_3684);
xor U3826 (N_3826,N_3695,N_3683);
xnor U3827 (N_3827,N_3633,N_3724);
nor U3828 (N_3828,N_3760,N_3785);
or U3829 (N_3829,N_3781,N_3639);
or U3830 (N_3830,N_3660,N_3644);
and U3831 (N_3831,N_3730,N_3702);
or U3832 (N_3832,N_3759,N_3645);
and U3833 (N_3833,N_3797,N_3796);
and U3834 (N_3834,N_3799,N_3761);
xnor U3835 (N_3835,N_3716,N_3748);
nor U3836 (N_3836,N_3619,N_3621);
and U3837 (N_3837,N_3650,N_3655);
nand U3838 (N_3838,N_3775,N_3713);
nand U3839 (N_3839,N_3734,N_3696);
or U3840 (N_3840,N_3782,N_3718);
nand U3841 (N_3841,N_3722,N_3701);
nor U3842 (N_3842,N_3625,N_3669);
nor U3843 (N_3843,N_3728,N_3681);
and U3844 (N_3844,N_3757,N_3687);
nor U3845 (N_3845,N_3714,N_3675);
nand U3846 (N_3846,N_3766,N_3672);
nor U3847 (N_3847,N_3790,N_3726);
and U3848 (N_3848,N_3741,N_3648);
nand U3849 (N_3849,N_3622,N_3688);
xor U3850 (N_3850,N_3674,N_3657);
or U3851 (N_3851,N_3661,N_3620);
nor U3852 (N_3852,N_3798,N_3778);
nand U3853 (N_3853,N_3732,N_3653);
nor U3854 (N_3854,N_3739,N_3753);
xor U3855 (N_3855,N_3623,N_3720);
or U3856 (N_3856,N_3678,N_3751);
nand U3857 (N_3857,N_3700,N_3754);
and U3858 (N_3858,N_3725,N_3694);
and U3859 (N_3859,N_3658,N_3715);
xor U3860 (N_3860,N_3763,N_3711);
nor U3861 (N_3861,N_3762,N_3656);
nand U3862 (N_3862,N_3712,N_3731);
xnor U3863 (N_3863,N_3632,N_3642);
nor U3864 (N_3864,N_3787,N_3768);
nor U3865 (N_3865,N_3607,N_3651);
nand U3866 (N_3866,N_3670,N_3659);
and U3867 (N_3867,N_3752,N_3740);
nand U3868 (N_3868,N_3729,N_3604);
nor U3869 (N_3869,N_3614,N_3765);
xnor U3870 (N_3870,N_3792,N_3699);
nand U3871 (N_3871,N_3636,N_3601);
nand U3872 (N_3872,N_3603,N_3723);
nand U3873 (N_3873,N_3616,N_3774);
or U3874 (N_3874,N_3671,N_3680);
or U3875 (N_3875,N_3682,N_3755);
and U3876 (N_3876,N_3697,N_3750);
or U3877 (N_3877,N_3784,N_3756);
or U3878 (N_3878,N_3733,N_3638);
nor U3879 (N_3879,N_3709,N_3719);
xnor U3880 (N_3880,N_3634,N_3612);
nor U3881 (N_3881,N_3624,N_3602);
nor U3882 (N_3882,N_3788,N_3793);
and U3883 (N_3883,N_3747,N_3698);
or U3884 (N_3884,N_3605,N_3769);
or U3885 (N_3885,N_3794,N_3736);
and U3886 (N_3886,N_3710,N_3643);
or U3887 (N_3887,N_3629,N_3617);
nor U3888 (N_3888,N_3749,N_3693);
nand U3889 (N_3889,N_3783,N_3789);
and U3890 (N_3890,N_3771,N_3735);
and U3891 (N_3891,N_3738,N_3606);
or U3892 (N_3892,N_3662,N_3640);
and U3893 (N_3893,N_3615,N_3686);
nand U3894 (N_3894,N_3666,N_3637);
and U3895 (N_3895,N_3706,N_3764);
nand U3896 (N_3896,N_3691,N_3676);
nand U3897 (N_3897,N_3779,N_3780);
or U3898 (N_3898,N_3673,N_3652);
nand U3899 (N_3899,N_3677,N_3628);
nand U3900 (N_3900,N_3644,N_3775);
nand U3901 (N_3901,N_3762,N_3755);
nand U3902 (N_3902,N_3732,N_3678);
nor U3903 (N_3903,N_3747,N_3613);
or U3904 (N_3904,N_3656,N_3756);
nor U3905 (N_3905,N_3694,N_3792);
and U3906 (N_3906,N_3771,N_3689);
xor U3907 (N_3907,N_3731,N_3638);
or U3908 (N_3908,N_3739,N_3637);
xnor U3909 (N_3909,N_3744,N_3738);
and U3910 (N_3910,N_3777,N_3623);
or U3911 (N_3911,N_3605,N_3663);
xnor U3912 (N_3912,N_3761,N_3678);
xor U3913 (N_3913,N_3664,N_3728);
nand U3914 (N_3914,N_3728,N_3695);
and U3915 (N_3915,N_3692,N_3778);
nand U3916 (N_3916,N_3795,N_3754);
or U3917 (N_3917,N_3796,N_3718);
nand U3918 (N_3918,N_3604,N_3607);
and U3919 (N_3919,N_3613,N_3623);
nand U3920 (N_3920,N_3750,N_3646);
or U3921 (N_3921,N_3671,N_3665);
and U3922 (N_3922,N_3713,N_3654);
and U3923 (N_3923,N_3793,N_3696);
and U3924 (N_3924,N_3702,N_3782);
or U3925 (N_3925,N_3696,N_3673);
or U3926 (N_3926,N_3601,N_3771);
and U3927 (N_3927,N_3652,N_3686);
nor U3928 (N_3928,N_3793,N_3748);
or U3929 (N_3929,N_3706,N_3677);
xor U3930 (N_3930,N_3663,N_3730);
nand U3931 (N_3931,N_3765,N_3773);
nor U3932 (N_3932,N_3765,N_3779);
and U3933 (N_3933,N_3727,N_3620);
and U3934 (N_3934,N_3627,N_3732);
nand U3935 (N_3935,N_3663,N_3722);
or U3936 (N_3936,N_3726,N_3742);
nand U3937 (N_3937,N_3784,N_3738);
and U3938 (N_3938,N_3620,N_3646);
nor U3939 (N_3939,N_3750,N_3675);
nand U3940 (N_3940,N_3669,N_3771);
and U3941 (N_3941,N_3786,N_3798);
and U3942 (N_3942,N_3659,N_3669);
nor U3943 (N_3943,N_3701,N_3796);
nand U3944 (N_3944,N_3640,N_3600);
and U3945 (N_3945,N_3750,N_3678);
nand U3946 (N_3946,N_3630,N_3686);
nand U3947 (N_3947,N_3600,N_3664);
and U3948 (N_3948,N_3632,N_3787);
nor U3949 (N_3949,N_3737,N_3611);
xor U3950 (N_3950,N_3663,N_3674);
xor U3951 (N_3951,N_3783,N_3717);
and U3952 (N_3952,N_3689,N_3718);
xor U3953 (N_3953,N_3778,N_3674);
or U3954 (N_3954,N_3794,N_3703);
or U3955 (N_3955,N_3750,N_3670);
and U3956 (N_3956,N_3742,N_3739);
nor U3957 (N_3957,N_3701,N_3622);
nor U3958 (N_3958,N_3769,N_3606);
and U3959 (N_3959,N_3759,N_3752);
nor U3960 (N_3960,N_3714,N_3666);
nand U3961 (N_3961,N_3722,N_3641);
nand U3962 (N_3962,N_3667,N_3746);
nand U3963 (N_3963,N_3638,N_3796);
and U3964 (N_3964,N_3658,N_3626);
nand U3965 (N_3965,N_3795,N_3766);
nor U3966 (N_3966,N_3753,N_3787);
nand U3967 (N_3967,N_3795,N_3719);
nand U3968 (N_3968,N_3733,N_3702);
nor U3969 (N_3969,N_3689,N_3750);
and U3970 (N_3970,N_3740,N_3768);
or U3971 (N_3971,N_3649,N_3717);
and U3972 (N_3972,N_3727,N_3718);
and U3973 (N_3973,N_3604,N_3663);
nand U3974 (N_3974,N_3796,N_3690);
or U3975 (N_3975,N_3695,N_3747);
or U3976 (N_3976,N_3605,N_3636);
or U3977 (N_3977,N_3708,N_3603);
nand U3978 (N_3978,N_3702,N_3793);
xor U3979 (N_3979,N_3630,N_3744);
nor U3980 (N_3980,N_3615,N_3763);
nand U3981 (N_3981,N_3716,N_3722);
nor U3982 (N_3982,N_3642,N_3732);
or U3983 (N_3983,N_3733,N_3615);
xor U3984 (N_3984,N_3707,N_3694);
or U3985 (N_3985,N_3671,N_3645);
nor U3986 (N_3986,N_3780,N_3794);
xor U3987 (N_3987,N_3788,N_3673);
nor U3988 (N_3988,N_3714,N_3659);
and U3989 (N_3989,N_3680,N_3655);
and U3990 (N_3990,N_3613,N_3641);
nor U3991 (N_3991,N_3647,N_3781);
nand U3992 (N_3992,N_3644,N_3767);
and U3993 (N_3993,N_3636,N_3782);
or U3994 (N_3994,N_3734,N_3660);
or U3995 (N_3995,N_3697,N_3756);
and U3996 (N_3996,N_3793,N_3629);
or U3997 (N_3997,N_3601,N_3659);
nand U3998 (N_3998,N_3777,N_3645);
nor U3999 (N_3999,N_3668,N_3601);
nor U4000 (N_4000,N_3857,N_3893);
nor U4001 (N_4001,N_3880,N_3957);
or U4002 (N_4002,N_3837,N_3997);
or U4003 (N_4003,N_3911,N_3828);
nor U4004 (N_4004,N_3897,N_3803);
or U4005 (N_4005,N_3918,N_3835);
nand U4006 (N_4006,N_3841,N_3962);
or U4007 (N_4007,N_3862,N_3853);
and U4008 (N_4008,N_3882,N_3826);
xor U4009 (N_4009,N_3929,N_3820);
and U4010 (N_4010,N_3941,N_3888);
nor U4011 (N_4011,N_3952,N_3872);
xnor U4012 (N_4012,N_3890,N_3815);
and U4013 (N_4013,N_3833,N_3840);
or U4014 (N_4014,N_3998,N_3933);
nand U4015 (N_4015,N_3969,N_3912);
or U4016 (N_4016,N_3905,N_3894);
xor U4017 (N_4017,N_3855,N_3867);
xor U4018 (N_4018,N_3966,N_3832);
or U4019 (N_4019,N_3866,N_3881);
nor U4020 (N_4020,N_3810,N_3917);
nor U4021 (N_4021,N_3934,N_3825);
and U4022 (N_4022,N_3923,N_3896);
nor U4023 (N_4023,N_3946,N_3886);
xnor U4024 (N_4024,N_3949,N_3987);
and U4025 (N_4025,N_3947,N_3860);
xnor U4026 (N_4026,N_3910,N_3907);
nor U4027 (N_4027,N_3839,N_3807);
xor U4028 (N_4028,N_3895,N_3909);
or U4029 (N_4029,N_3927,N_3887);
nand U4030 (N_4030,N_3816,N_3982);
nand U4031 (N_4031,N_3849,N_3968);
nand U4032 (N_4032,N_3830,N_3842);
xnor U4033 (N_4033,N_3979,N_3956);
xor U4034 (N_4034,N_3906,N_3925);
nand U4035 (N_4035,N_3986,N_3959);
nor U4036 (N_4036,N_3932,N_3821);
or U4037 (N_4037,N_3920,N_3989);
nand U4038 (N_4038,N_3824,N_3964);
and U4039 (N_4039,N_3943,N_3924);
nor U4040 (N_4040,N_3935,N_3983);
or U4041 (N_4041,N_3819,N_3838);
and U4042 (N_4042,N_3990,N_3802);
nand U4043 (N_4043,N_3850,N_3991);
and U4044 (N_4044,N_3811,N_3854);
nand U4045 (N_4045,N_3901,N_3945);
nor U4046 (N_4046,N_3916,N_3831);
nand U4047 (N_4047,N_3926,N_3885);
or U4048 (N_4048,N_3981,N_3823);
nor U4049 (N_4049,N_3873,N_3851);
nor U4050 (N_4050,N_3898,N_3936);
nor U4051 (N_4051,N_3939,N_3861);
or U4052 (N_4052,N_3971,N_3829);
or U4053 (N_4053,N_3868,N_3856);
and U4054 (N_4054,N_3875,N_3836);
and U4055 (N_4055,N_3847,N_3994);
nand U4056 (N_4056,N_3859,N_3974);
or U4057 (N_4057,N_3940,N_3919);
or U4058 (N_4058,N_3852,N_3814);
xnor U4059 (N_4059,N_3812,N_3822);
nor U4060 (N_4060,N_3996,N_3958);
and U4061 (N_4061,N_3928,N_3902);
nor U4062 (N_4062,N_3865,N_3955);
and U4063 (N_4063,N_3953,N_3801);
and U4064 (N_4064,N_3980,N_3874);
and U4065 (N_4065,N_3915,N_3985);
and U4066 (N_4066,N_3995,N_3976);
nand U4067 (N_4067,N_3863,N_3843);
and U4068 (N_4068,N_3848,N_3846);
nand U4069 (N_4069,N_3922,N_3800);
and U4070 (N_4070,N_3883,N_3899);
or U4071 (N_4071,N_3876,N_3977);
or U4072 (N_4072,N_3992,N_3944);
xnor U4073 (N_4073,N_3930,N_3948);
or U4074 (N_4074,N_3931,N_3993);
nor U4075 (N_4075,N_3889,N_3938);
nor U4076 (N_4076,N_3975,N_3978);
nor U4077 (N_4077,N_3805,N_3813);
and U4078 (N_4078,N_3884,N_3864);
and U4079 (N_4079,N_3869,N_3913);
and U4080 (N_4080,N_3965,N_3963);
and U4081 (N_4081,N_3921,N_3973);
and U4082 (N_4082,N_3834,N_3808);
xnor U4083 (N_4083,N_3844,N_3908);
and U4084 (N_4084,N_3914,N_3970);
or U4085 (N_4085,N_3942,N_3967);
and U4086 (N_4086,N_3999,N_3961);
and U4087 (N_4087,N_3892,N_3818);
or U4088 (N_4088,N_3809,N_3870);
xor U4089 (N_4089,N_3817,N_3988);
nor U4090 (N_4090,N_3903,N_3900);
and U4091 (N_4091,N_3904,N_3878);
xor U4092 (N_4092,N_3879,N_3827);
or U4093 (N_4093,N_3960,N_3871);
nor U4094 (N_4094,N_3984,N_3858);
nor U4095 (N_4095,N_3804,N_3951);
or U4096 (N_4096,N_3891,N_3954);
nor U4097 (N_4097,N_3937,N_3806);
nand U4098 (N_4098,N_3972,N_3877);
and U4099 (N_4099,N_3845,N_3950);
or U4100 (N_4100,N_3843,N_3828);
or U4101 (N_4101,N_3962,N_3905);
nor U4102 (N_4102,N_3802,N_3940);
and U4103 (N_4103,N_3869,N_3888);
nor U4104 (N_4104,N_3964,N_3861);
or U4105 (N_4105,N_3810,N_3869);
nand U4106 (N_4106,N_3837,N_3851);
nand U4107 (N_4107,N_3955,N_3964);
and U4108 (N_4108,N_3900,N_3836);
and U4109 (N_4109,N_3934,N_3941);
and U4110 (N_4110,N_3953,N_3967);
nor U4111 (N_4111,N_3862,N_3814);
xor U4112 (N_4112,N_3894,N_3856);
and U4113 (N_4113,N_3834,N_3936);
or U4114 (N_4114,N_3977,N_3809);
xnor U4115 (N_4115,N_3961,N_3918);
and U4116 (N_4116,N_3931,N_3858);
nor U4117 (N_4117,N_3808,N_3868);
and U4118 (N_4118,N_3970,N_3852);
nand U4119 (N_4119,N_3935,N_3851);
or U4120 (N_4120,N_3821,N_3966);
and U4121 (N_4121,N_3997,N_3972);
or U4122 (N_4122,N_3829,N_3962);
or U4123 (N_4123,N_3998,N_3823);
nand U4124 (N_4124,N_3905,N_3909);
nor U4125 (N_4125,N_3999,N_3907);
nor U4126 (N_4126,N_3979,N_3903);
and U4127 (N_4127,N_3934,N_3878);
xnor U4128 (N_4128,N_3857,N_3890);
or U4129 (N_4129,N_3835,N_3858);
nand U4130 (N_4130,N_3997,N_3830);
or U4131 (N_4131,N_3861,N_3869);
xnor U4132 (N_4132,N_3847,N_3978);
xor U4133 (N_4133,N_3969,N_3869);
and U4134 (N_4134,N_3863,N_3857);
and U4135 (N_4135,N_3834,N_3810);
nand U4136 (N_4136,N_3887,N_3934);
or U4137 (N_4137,N_3963,N_3925);
and U4138 (N_4138,N_3823,N_3853);
nand U4139 (N_4139,N_3962,N_3810);
and U4140 (N_4140,N_3870,N_3884);
nand U4141 (N_4141,N_3862,N_3800);
nor U4142 (N_4142,N_3828,N_3831);
nand U4143 (N_4143,N_3822,N_3956);
nor U4144 (N_4144,N_3891,N_3957);
nor U4145 (N_4145,N_3944,N_3848);
nor U4146 (N_4146,N_3878,N_3937);
nand U4147 (N_4147,N_3992,N_3953);
and U4148 (N_4148,N_3962,N_3809);
nand U4149 (N_4149,N_3956,N_3816);
nor U4150 (N_4150,N_3884,N_3899);
nor U4151 (N_4151,N_3832,N_3999);
and U4152 (N_4152,N_3814,N_3870);
or U4153 (N_4153,N_3845,N_3853);
nand U4154 (N_4154,N_3907,N_3849);
and U4155 (N_4155,N_3927,N_3997);
nor U4156 (N_4156,N_3834,N_3880);
and U4157 (N_4157,N_3902,N_3901);
and U4158 (N_4158,N_3978,N_3906);
nand U4159 (N_4159,N_3865,N_3944);
xnor U4160 (N_4160,N_3898,N_3816);
nor U4161 (N_4161,N_3956,N_3817);
nor U4162 (N_4162,N_3951,N_3818);
nor U4163 (N_4163,N_3889,N_3972);
or U4164 (N_4164,N_3850,N_3917);
and U4165 (N_4165,N_3971,N_3947);
or U4166 (N_4166,N_3947,N_3889);
nand U4167 (N_4167,N_3983,N_3948);
and U4168 (N_4168,N_3896,N_3965);
nand U4169 (N_4169,N_3898,N_3979);
xor U4170 (N_4170,N_3884,N_3847);
xor U4171 (N_4171,N_3843,N_3968);
nor U4172 (N_4172,N_3832,N_3876);
nand U4173 (N_4173,N_3878,N_3888);
and U4174 (N_4174,N_3939,N_3921);
nand U4175 (N_4175,N_3939,N_3835);
and U4176 (N_4176,N_3998,N_3961);
and U4177 (N_4177,N_3930,N_3882);
or U4178 (N_4178,N_3821,N_3955);
or U4179 (N_4179,N_3934,N_3868);
or U4180 (N_4180,N_3895,N_3960);
and U4181 (N_4181,N_3988,N_3909);
nand U4182 (N_4182,N_3881,N_3842);
nand U4183 (N_4183,N_3910,N_3852);
and U4184 (N_4184,N_3875,N_3940);
and U4185 (N_4185,N_3872,N_3846);
nand U4186 (N_4186,N_3950,N_3914);
and U4187 (N_4187,N_3951,N_3953);
nor U4188 (N_4188,N_3862,N_3976);
nor U4189 (N_4189,N_3842,N_3812);
nor U4190 (N_4190,N_3905,N_3900);
or U4191 (N_4191,N_3960,N_3920);
and U4192 (N_4192,N_3920,N_3992);
and U4193 (N_4193,N_3828,N_3921);
nand U4194 (N_4194,N_3842,N_3936);
or U4195 (N_4195,N_3993,N_3976);
or U4196 (N_4196,N_3983,N_3993);
nor U4197 (N_4197,N_3897,N_3840);
nor U4198 (N_4198,N_3809,N_3802);
or U4199 (N_4199,N_3939,N_3925);
nor U4200 (N_4200,N_4192,N_4109);
nand U4201 (N_4201,N_4138,N_4014);
or U4202 (N_4202,N_4096,N_4050);
or U4203 (N_4203,N_4193,N_4115);
and U4204 (N_4204,N_4082,N_4052);
and U4205 (N_4205,N_4163,N_4040);
nand U4206 (N_4206,N_4059,N_4048);
nand U4207 (N_4207,N_4039,N_4133);
nand U4208 (N_4208,N_4101,N_4100);
and U4209 (N_4209,N_4197,N_4142);
nand U4210 (N_4210,N_4098,N_4137);
and U4211 (N_4211,N_4134,N_4147);
or U4212 (N_4212,N_4168,N_4081);
nor U4213 (N_4213,N_4186,N_4021);
xnor U4214 (N_4214,N_4057,N_4019);
nand U4215 (N_4215,N_4171,N_4135);
nor U4216 (N_4216,N_4068,N_4055);
nor U4217 (N_4217,N_4003,N_4183);
xnor U4218 (N_4218,N_4159,N_4174);
nor U4219 (N_4219,N_4132,N_4184);
or U4220 (N_4220,N_4090,N_4073);
xor U4221 (N_4221,N_4024,N_4060);
or U4222 (N_4222,N_4111,N_4145);
and U4223 (N_4223,N_4113,N_4185);
and U4224 (N_4224,N_4030,N_4033);
and U4225 (N_4225,N_4141,N_4128);
xor U4226 (N_4226,N_4117,N_4144);
nor U4227 (N_4227,N_4162,N_4054);
and U4228 (N_4228,N_4061,N_4131);
nor U4229 (N_4229,N_4148,N_4175);
and U4230 (N_4230,N_4152,N_4074);
and U4231 (N_4231,N_4170,N_4045);
and U4232 (N_4232,N_4064,N_4124);
and U4233 (N_4233,N_4058,N_4108);
and U4234 (N_4234,N_4002,N_4028);
and U4235 (N_4235,N_4087,N_4049);
or U4236 (N_4236,N_4075,N_4089);
or U4237 (N_4237,N_4027,N_4165);
or U4238 (N_4238,N_4187,N_4072);
xnor U4239 (N_4239,N_4046,N_4023);
nand U4240 (N_4240,N_4155,N_4102);
or U4241 (N_4241,N_4084,N_4047);
and U4242 (N_4242,N_4069,N_4121);
or U4243 (N_4243,N_4161,N_4026);
or U4244 (N_4244,N_4062,N_4078);
or U4245 (N_4245,N_4079,N_4025);
or U4246 (N_4246,N_4169,N_4119);
xnor U4247 (N_4247,N_4116,N_4136);
and U4248 (N_4248,N_4013,N_4146);
nand U4249 (N_4249,N_4035,N_4020);
or U4250 (N_4250,N_4114,N_4157);
or U4251 (N_4251,N_4120,N_4009);
or U4252 (N_4252,N_4151,N_4130);
nor U4253 (N_4253,N_4140,N_4000);
nand U4254 (N_4254,N_4001,N_4189);
and U4255 (N_4255,N_4180,N_4006);
and U4256 (N_4256,N_4066,N_4007);
and U4257 (N_4257,N_4094,N_4037);
or U4258 (N_4258,N_4005,N_4158);
nand U4259 (N_4259,N_4199,N_4143);
nor U4260 (N_4260,N_4092,N_4012);
or U4261 (N_4261,N_4182,N_4016);
or U4262 (N_4262,N_4172,N_4154);
xor U4263 (N_4263,N_4188,N_4125);
or U4264 (N_4264,N_4076,N_4085);
nor U4265 (N_4265,N_4164,N_4106);
nor U4266 (N_4266,N_4160,N_4011);
nand U4267 (N_4267,N_4107,N_4086);
nor U4268 (N_4268,N_4017,N_4008);
nand U4269 (N_4269,N_4194,N_4190);
nor U4270 (N_4270,N_4044,N_4041);
nor U4271 (N_4271,N_4177,N_4112);
or U4272 (N_4272,N_4198,N_4051);
and U4273 (N_4273,N_4127,N_4053);
or U4274 (N_4274,N_4097,N_4126);
nor U4275 (N_4275,N_4043,N_4179);
or U4276 (N_4276,N_4042,N_4156);
nor U4277 (N_4277,N_4010,N_4196);
and U4278 (N_4278,N_4167,N_4015);
nor U4279 (N_4279,N_4022,N_4077);
nor U4280 (N_4280,N_4088,N_4070);
or U4281 (N_4281,N_4139,N_4067);
nor U4282 (N_4282,N_4099,N_4103);
xnor U4283 (N_4283,N_4173,N_4122);
and U4284 (N_4284,N_4181,N_4083);
nor U4285 (N_4285,N_4195,N_4176);
nor U4286 (N_4286,N_4065,N_4166);
xor U4287 (N_4287,N_4036,N_4063);
and U4288 (N_4288,N_4071,N_4029);
and U4289 (N_4289,N_4153,N_4118);
nor U4290 (N_4290,N_4056,N_4150);
nor U4291 (N_4291,N_4105,N_4123);
nand U4292 (N_4292,N_4093,N_4091);
nand U4293 (N_4293,N_4034,N_4080);
and U4294 (N_4294,N_4178,N_4149);
and U4295 (N_4295,N_4191,N_4032);
nor U4296 (N_4296,N_4095,N_4004);
nand U4297 (N_4297,N_4129,N_4031);
or U4298 (N_4298,N_4104,N_4018);
nor U4299 (N_4299,N_4038,N_4110);
nand U4300 (N_4300,N_4188,N_4138);
nand U4301 (N_4301,N_4093,N_4025);
or U4302 (N_4302,N_4000,N_4109);
nor U4303 (N_4303,N_4048,N_4058);
nand U4304 (N_4304,N_4104,N_4143);
and U4305 (N_4305,N_4184,N_4105);
nor U4306 (N_4306,N_4031,N_4160);
and U4307 (N_4307,N_4120,N_4182);
nand U4308 (N_4308,N_4115,N_4025);
nor U4309 (N_4309,N_4016,N_4057);
nand U4310 (N_4310,N_4139,N_4095);
nor U4311 (N_4311,N_4162,N_4177);
nand U4312 (N_4312,N_4049,N_4143);
or U4313 (N_4313,N_4003,N_4158);
or U4314 (N_4314,N_4174,N_4155);
and U4315 (N_4315,N_4171,N_4057);
or U4316 (N_4316,N_4046,N_4089);
and U4317 (N_4317,N_4080,N_4123);
nand U4318 (N_4318,N_4038,N_4147);
nand U4319 (N_4319,N_4003,N_4032);
or U4320 (N_4320,N_4158,N_4133);
or U4321 (N_4321,N_4175,N_4174);
nand U4322 (N_4322,N_4150,N_4167);
nor U4323 (N_4323,N_4078,N_4188);
or U4324 (N_4324,N_4073,N_4158);
nand U4325 (N_4325,N_4154,N_4123);
nand U4326 (N_4326,N_4096,N_4032);
nor U4327 (N_4327,N_4054,N_4091);
xnor U4328 (N_4328,N_4068,N_4106);
nor U4329 (N_4329,N_4176,N_4030);
xnor U4330 (N_4330,N_4176,N_4104);
xnor U4331 (N_4331,N_4080,N_4114);
or U4332 (N_4332,N_4140,N_4036);
nor U4333 (N_4333,N_4015,N_4161);
nand U4334 (N_4334,N_4160,N_4007);
or U4335 (N_4335,N_4098,N_4075);
nor U4336 (N_4336,N_4081,N_4071);
or U4337 (N_4337,N_4032,N_4037);
nor U4338 (N_4338,N_4173,N_4073);
or U4339 (N_4339,N_4114,N_4123);
and U4340 (N_4340,N_4169,N_4095);
and U4341 (N_4341,N_4000,N_4137);
and U4342 (N_4342,N_4162,N_4084);
or U4343 (N_4343,N_4007,N_4182);
and U4344 (N_4344,N_4051,N_4096);
and U4345 (N_4345,N_4159,N_4128);
nor U4346 (N_4346,N_4000,N_4124);
and U4347 (N_4347,N_4068,N_4053);
nor U4348 (N_4348,N_4101,N_4075);
xnor U4349 (N_4349,N_4089,N_4036);
or U4350 (N_4350,N_4146,N_4192);
nand U4351 (N_4351,N_4004,N_4025);
or U4352 (N_4352,N_4098,N_4164);
or U4353 (N_4353,N_4050,N_4156);
xnor U4354 (N_4354,N_4065,N_4160);
and U4355 (N_4355,N_4022,N_4115);
or U4356 (N_4356,N_4172,N_4005);
or U4357 (N_4357,N_4104,N_4199);
nor U4358 (N_4358,N_4160,N_4010);
and U4359 (N_4359,N_4105,N_4025);
or U4360 (N_4360,N_4046,N_4063);
nor U4361 (N_4361,N_4006,N_4176);
xnor U4362 (N_4362,N_4098,N_4113);
and U4363 (N_4363,N_4055,N_4006);
nand U4364 (N_4364,N_4067,N_4173);
nor U4365 (N_4365,N_4143,N_4032);
xor U4366 (N_4366,N_4039,N_4137);
or U4367 (N_4367,N_4145,N_4188);
nor U4368 (N_4368,N_4003,N_4109);
nand U4369 (N_4369,N_4015,N_4139);
nand U4370 (N_4370,N_4029,N_4103);
nor U4371 (N_4371,N_4021,N_4168);
or U4372 (N_4372,N_4164,N_4012);
or U4373 (N_4373,N_4022,N_4144);
xnor U4374 (N_4374,N_4110,N_4154);
nor U4375 (N_4375,N_4074,N_4185);
or U4376 (N_4376,N_4004,N_4100);
and U4377 (N_4377,N_4126,N_4020);
or U4378 (N_4378,N_4042,N_4082);
and U4379 (N_4379,N_4021,N_4049);
nand U4380 (N_4380,N_4022,N_4146);
nand U4381 (N_4381,N_4158,N_4029);
and U4382 (N_4382,N_4186,N_4050);
or U4383 (N_4383,N_4111,N_4135);
nand U4384 (N_4384,N_4024,N_4050);
and U4385 (N_4385,N_4131,N_4013);
and U4386 (N_4386,N_4067,N_4045);
nand U4387 (N_4387,N_4156,N_4045);
or U4388 (N_4388,N_4020,N_4199);
or U4389 (N_4389,N_4177,N_4169);
and U4390 (N_4390,N_4005,N_4081);
and U4391 (N_4391,N_4172,N_4056);
xor U4392 (N_4392,N_4049,N_4122);
nor U4393 (N_4393,N_4099,N_4078);
nor U4394 (N_4394,N_4008,N_4014);
and U4395 (N_4395,N_4108,N_4048);
nand U4396 (N_4396,N_4195,N_4164);
nand U4397 (N_4397,N_4008,N_4043);
nand U4398 (N_4398,N_4043,N_4151);
nand U4399 (N_4399,N_4127,N_4155);
nor U4400 (N_4400,N_4340,N_4305);
and U4401 (N_4401,N_4389,N_4388);
nor U4402 (N_4402,N_4215,N_4283);
nand U4403 (N_4403,N_4297,N_4392);
nor U4404 (N_4404,N_4384,N_4218);
and U4405 (N_4405,N_4375,N_4380);
or U4406 (N_4406,N_4357,N_4238);
or U4407 (N_4407,N_4336,N_4247);
and U4408 (N_4408,N_4367,N_4202);
or U4409 (N_4409,N_4321,N_4379);
nand U4410 (N_4410,N_4311,N_4222);
nand U4411 (N_4411,N_4354,N_4224);
and U4412 (N_4412,N_4217,N_4234);
nand U4413 (N_4413,N_4219,N_4237);
xor U4414 (N_4414,N_4239,N_4214);
or U4415 (N_4415,N_4213,N_4250);
or U4416 (N_4416,N_4211,N_4356);
nor U4417 (N_4417,N_4272,N_4320);
nand U4418 (N_4418,N_4368,N_4240);
nand U4419 (N_4419,N_4361,N_4207);
nand U4420 (N_4420,N_4391,N_4353);
nor U4421 (N_4421,N_4335,N_4270);
nand U4422 (N_4422,N_4387,N_4251);
nand U4423 (N_4423,N_4352,N_4230);
and U4424 (N_4424,N_4294,N_4277);
nand U4425 (N_4425,N_4310,N_4386);
and U4426 (N_4426,N_4268,N_4377);
nand U4427 (N_4427,N_4256,N_4227);
xor U4428 (N_4428,N_4280,N_4314);
nor U4429 (N_4429,N_4249,N_4397);
nor U4430 (N_4430,N_4241,N_4329);
and U4431 (N_4431,N_4366,N_4263);
and U4432 (N_4432,N_4303,N_4350);
nor U4433 (N_4433,N_4383,N_4229);
nand U4434 (N_4434,N_4226,N_4369);
and U4435 (N_4435,N_4206,N_4275);
nand U4436 (N_4436,N_4262,N_4342);
and U4437 (N_4437,N_4209,N_4338);
or U4438 (N_4438,N_4323,N_4278);
or U4439 (N_4439,N_4223,N_4259);
or U4440 (N_4440,N_4279,N_4299);
nor U4441 (N_4441,N_4376,N_4208);
nand U4442 (N_4442,N_4344,N_4390);
nor U4443 (N_4443,N_4243,N_4362);
xor U4444 (N_4444,N_4203,N_4364);
nor U4445 (N_4445,N_4261,N_4260);
nor U4446 (N_4446,N_4381,N_4204);
and U4447 (N_4447,N_4284,N_4317);
xor U4448 (N_4448,N_4269,N_4306);
nand U4449 (N_4449,N_4273,N_4265);
or U4450 (N_4450,N_4205,N_4324);
nand U4451 (N_4451,N_4290,N_4398);
nand U4452 (N_4452,N_4287,N_4395);
or U4453 (N_4453,N_4212,N_4337);
and U4454 (N_4454,N_4292,N_4359);
and U4455 (N_4455,N_4246,N_4348);
nor U4456 (N_4456,N_4382,N_4286);
and U4457 (N_4457,N_4235,N_4231);
xnor U4458 (N_4458,N_4349,N_4347);
or U4459 (N_4459,N_4258,N_4295);
xor U4460 (N_4460,N_4331,N_4300);
nand U4461 (N_4461,N_4319,N_4274);
nand U4462 (N_4462,N_4264,N_4216);
nand U4463 (N_4463,N_4228,N_4365);
or U4464 (N_4464,N_4254,N_4298);
or U4465 (N_4465,N_4225,N_4200);
nor U4466 (N_4466,N_4308,N_4289);
xnor U4467 (N_4467,N_4236,N_4302);
xor U4468 (N_4468,N_4328,N_4355);
and U4469 (N_4469,N_4360,N_4291);
or U4470 (N_4470,N_4339,N_4330);
xor U4471 (N_4471,N_4245,N_4242);
and U4472 (N_4472,N_4307,N_4232);
and U4473 (N_4473,N_4282,N_4201);
or U4474 (N_4474,N_4370,N_4334);
nor U4475 (N_4475,N_4363,N_4276);
or U4476 (N_4476,N_4285,N_4244);
or U4477 (N_4477,N_4316,N_4327);
or U4478 (N_4478,N_4399,N_4393);
and U4479 (N_4479,N_4318,N_4346);
nand U4480 (N_4480,N_4345,N_4293);
nand U4481 (N_4481,N_4332,N_4341);
nand U4482 (N_4482,N_4233,N_4315);
xor U4483 (N_4483,N_4220,N_4296);
nor U4484 (N_4484,N_4221,N_4309);
nor U4485 (N_4485,N_4378,N_4371);
nor U4486 (N_4486,N_4343,N_4333);
xor U4487 (N_4487,N_4325,N_4372);
nor U4488 (N_4488,N_4248,N_4374);
or U4489 (N_4489,N_4266,N_4396);
nand U4490 (N_4490,N_4385,N_4351);
nor U4491 (N_4491,N_4326,N_4255);
and U4492 (N_4492,N_4210,N_4301);
nor U4493 (N_4493,N_4257,N_4253);
or U4494 (N_4494,N_4252,N_4358);
nor U4495 (N_4495,N_4313,N_4267);
nand U4496 (N_4496,N_4288,N_4394);
or U4497 (N_4497,N_4322,N_4271);
or U4498 (N_4498,N_4312,N_4281);
and U4499 (N_4499,N_4304,N_4373);
nand U4500 (N_4500,N_4238,N_4343);
or U4501 (N_4501,N_4264,N_4309);
or U4502 (N_4502,N_4352,N_4310);
or U4503 (N_4503,N_4315,N_4265);
or U4504 (N_4504,N_4280,N_4288);
nor U4505 (N_4505,N_4229,N_4363);
nor U4506 (N_4506,N_4254,N_4288);
nor U4507 (N_4507,N_4254,N_4366);
and U4508 (N_4508,N_4386,N_4294);
nand U4509 (N_4509,N_4365,N_4230);
nor U4510 (N_4510,N_4343,N_4295);
and U4511 (N_4511,N_4297,N_4265);
nor U4512 (N_4512,N_4390,N_4338);
or U4513 (N_4513,N_4269,N_4219);
nand U4514 (N_4514,N_4297,N_4235);
nand U4515 (N_4515,N_4343,N_4304);
and U4516 (N_4516,N_4320,N_4318);
and U4517 (N_4517,N_4257,N_4383);
nand U4518 (N_4518,N_4336,N_4254);
xor U4519 (N_4519,N_4266,N_4208);
xor U4520 (N_4520,N_4268,N_4257);
xnor U4521 (N_4521,N_4244,N_4248);
nor U4522 (N_4522,N_4272,N_4280);
xnor U4523 (N_4523,N_4349,N_4236);
or U4524 (N_4524,N_4379,N_4394);
nor U4525 (N_4525,N_4234,N_4244);
and U4526 (N_4526,N_4323,N_4316);
and U4527 (N_4527,N_4341,N_4253);
nor U4528 (N_4528,N_4312,N_4285);
and U4529 (N_4529,N_4367,N_4232);
or U4530 (N_4530,N_4201,N_4367);
nand U4531 (N_4531,N_4312,N_4349);
nor U4532 (N_4532,N_4224,N_4390);
nor U4533 (N_4533,N_4279,N_4211);
xnor U4534 (N_4534,N_4399,N_4207);
or U4535 (N_4535,N_4210,N_4350);
nor U4536 (N_4536,N_4318,N_4292);
or U4537 (N_4537,N_4208,N_4395);
nor U4538 (N_4538,N_4209,N_4312);
and U4539 (N_4539,N_4242,N_4371);
and U4540 (N_4540,N_4334,N_4213);
and U4541 (N_4541,N_4311,N_4287);
nor U4542 (N_4542,N_4212,N_4243);
xnor U4543 (N_4543,N_4337,N_4257);
or U4544 (N_4544,N_4241,N_4378);
nor U4545 (N_4545,N_4258,N_4304);
and U4546 (N_4546,N_4318,N_4316);
or U4547 (N_4547,N_4367,N_4285);
and U4548 (N_4548,N_4237,N_4310);
nor U4549 (N_4549,N_4308,N_4283);
nand U4550 (N_4550,N_4240,N_4315);
or U4551 (N_4551,N_4395,N_4373);
nor U4552 (N_4552,N_4298,N_4280);
and U4553 (N_4553,N_4284,N_4389);
nor U4554 (N_4554,N_4376,N_4285);
nor U4555 (N_4555,N_4201,N_4371);
and U4556 (N_4556,N_4201,N_4307);
or U4557 (N_4557,N_4265,N_4215);
or U4558 (N_4558,N_4304,N_4215);
nand U4559 (N_4559,N_4206,N_4321);
nand U4560 (N_4560,N_4307,N_4309);
nor U4561 (N_4561,N_4386,N_4255);
and U4562 (N_4562,N_4296,N_4212);
or U4563 (N_4563,N_4332,N_4371);
nor U4564 (N_4564,N_4206,N_4385);
nor U4565 (N_4565,N_4357,N_4216);
nand U4566 (N_4566,N_4299,N_4296);
and U4567 (N_4567,N_4297,N_4375);
and U4568 (N_4568,N_4387,N_4326);
nor U4569 (N_4569,N_4334,N_4397);
or U4570 (N_4570,N_4320,N_4227);
and U4571 (N_4571,N_4293,N_4228);
nand U4572 (N_4572,N_4323,N_4321);
and U4573 (N_4573,N_4344,N_4243);
xor U4574 (N_4574,N_4283,N_4235);
or U4575 (N_4575,N_4204,N_4399);
nand U4576 (N_4576,N_4371,N_4286);
or U4577 (N_4577,N_4257,N_4223);
nand U4578 (N_4578,N_4387,N_4383);
nor U4579 (N_4579,N_4252,N_4385);
nand U4580 (N_4580,N_4371,N_4249);
and U4581 (N_4581,N_4233,N_4322);
or U4582 (N_4582,N_4305,N_4364);
or U4583 (N_4583,N_4366,N_4214);
or U4584 (N_4584,N_4234,N_4304);
nor U4585 (N_4585,N_4385,N_4302);
or U4586 (N_4586,N_4355,N_4235);
nand U4587 (N_4587,N_4273,N_4386);
and U4588 (N_4588,N_4246,N_4210);
or U4589 (N_4589,N_4226,N_4334);
or U4590 (N_4590,N_4394,N_4384);
nor U4591 (N_4591,N_4328,N_4268);
or U4592 (N_4592,N_4336,N_4233);
nand U4593 (N_4593,N_4205,N_4272);
and U4594 (N_4594,N_4286,N_4375);
nand U4595 (N_4595,N_4250,N_4324);
nor U4596 (N_4596,N_4381,N_4284);
and U4597 (N_4597,N_4275,N_4297);
or U4598 (N_4598,N_4291,N_4202);
and U4599 (N_4599,N_4249,N_4292);
xnor U4600 (N_4600,N_4515,N_4436);
and U4601 (N_4601,N_4416,N_4415);
xnor U4602 (N_4602,N_4487,N_4484);
nor U4603 (N_4603,N_4532,N_4439);
nor U4604 (N_4604,N_4521,N_4480);
and U4605 (N_4605,N_4432,N_4522);
nand U4606 (N_4606,N_4543,N_4590);
nor U4607 (N_4607,N_4448,N_4496);
nor U4608 (N_4608,N_4404,N_4508);
nand U4609 (N_4609,N_4463,N_4402);
nand U4610 (N_4610,N_4467,N_4506);
and U4611 (N_4611,N_4425,N_4538);
nor U4612 (N_4612,N_4460,N_4498);
nand U4613 (N_4613,N_4502,N_4580);
or U4614 (N_4614,N_4560,N_4567);
or U4615 (N_4615,N_4566,N_4454);
or U4616 (N_4616,N_4535,N_4469);
nand U4617 (N_4617,N_4572,N_4418);
xnor U4618 (N_4618,N_4514,N_4583);
and U4619 (N_4619,N_4471,N_4458);
nand U4620 (N_4620,N_4599,N_4413);
nor U4621 (N_4621,N_4499,N_4568);
or U4622 (N_4622,N_4529,N_4588);
nand U4623 (N_4623,N_4489,N_4497);
nand U4624 (N_4624,N_4466,N_4513);
nand U4625 (N_4625,N_4531,N_4575);
and U4626 (N_4626,N_4481,N_4527);
nor U4627 (N_4627,N_4452,N_4546);
nor U4628 (N_4628,N_4491,N_4478);
nand U4629 (N_4629,N_4505,N_4435);
or U4630 (N_4630,N_4445,N_4421);
and U4631 (N_4631,N_4406,N_4552);
and U4632 (N_4632,N_4594,N_4537);
and U4633 (N_4633,N_4561,N_4595);
and U4634 (N_4634,N_4585,N_4405);
nand U4635 (N_4635,N_4555,N_4540);
nand U4636 (N_4636,N_4430,N_4455);
xor U4637 (N_4637,N_4541,N_4507);
nor U4638 (N_4638,N_4446,N_4582);
nor U4639 (N_4639,N_4400,N_4420);
and U4640 (N_4640,N_4557,N_4524);
and U4641 (N_4641,N_4441,N_4519);
and U4642 (N_4642,N_4553,N_4509);
nor U4643 (N_4643,N_4417,N_4401);
or U4644 (N_4644,N_4495,N_4556);
xor U4645 (N_4645,N_4477,N_4525);
nor U4646 (N_4646,N_4563,N_4450);
or U4647 (N_4647,N_4479,N_4485);
xnor U4648 (N_4648,N_4438,N_4523);
nor U4649 (N_4649,N_4554,N_4437);
nor U4650 (N_4650,N_4520,N_4596);
or U4651 (N_4651,N_4564,N_4545);
nand U4652 (N_4652,N_4573,N_4407);
nand U4653 (N_4653,N_4449,N_4547);
nand U4654 (N_4654,N_4410,N_4409);
nor U4655 (N_4655,N_4482,N_4592);
and U4656 (N_4656,N_4476,N_4510);
nor U4657 (N_4657,N_4403,N_4411);
or U4658 (N_4658,N_4548,N_4518);
and U4659 (N_4659,N_4549,N_4512);
nor U4660 (N_4660,N_4490,N_4551);
or U4661 (N_4661,N_4593,N_4494);
or U4662 (N_4662,N_4419,N_4465);
or U4663 (N_4663,N_4559,N_4422);
nand U4664 (N_4664,N_4504,N_4483);
nand U4665 (N_4665,N_4459,N_4470);
xnor U4666 (N_4666,N_4558,N_4565);
and U4667 (N_4667,N_4577,N_4571);
nor U4668 (N_4668,N_4501,N_4492);
nand U4669 (N_4669,N_4428,N_4433);
nand U4670 (N_4670,N_4427,N_4550);
and U4671 (N_4671,N_4464,N_4591);
nand U4672 (N_4672,N_4534,N_4536);
xor U4673 (N_4673,N_4586,N_4475);
and U4674 (N_4674,N_4579,N_4424);
nand U4675 (N_4675,N_4472,N_4576);
and U4676 (N_4676,N_4581,N_4451);
nand U4677 (N_4677,N_4493,N_4598);
nor U4678 (N_4678,N_4578,N_4511);
nand U4679 (N_4679,N_4442,N_4569);
xnor U4680 (N_4680,N_4517,N_4503);
nor U4681 (N_4681,N_4408,N_4423);
xnor U4682 (N_4682,N_4434,N_4468);
nand U4683 (N_4683,N_4414,N_4574);
or U4684 (N_4684,N_4533,N_4597);
nor U4685 (N_4685,N_4457,N_4500);
or U4686 (N_4686,N_4447,N_4486);
nor U4687 (N_4687,N_4474,N_4456);
nor U4688 (N_4688,N_4530,N_4444);
xnor U4689 (N_4689,N_4544,N_4473);
nand U4690 (N_4690,N_4453,N_4587);
nor U4691 (N_4691,N_4488,N_4443);
nor U4692 (N_4692,N_4584,N_4440);
nand U4693 (N_4693,N_4426,N_4516);
nor U4694 (N_4694,N_4462,N_4539);
nor U4695 (N_4695,N_4526,N_4570);
nor U4696 (N_4696,N_4528,N_4412);
nor U4697 (N_4697,N_4429,N_4542);
and U4698 (N_4698,N_4562,N_4431);
or U4699 (N_4699,N_4589,N_4461);
or U4700 (N_4700,N_4498,N_4575);
nor U4701 (N_4701,N_4530,N_4544);
xnor U4702 (N_4702,N_4510,N_4473);
or U4703 (N_4703,N_4455,N_4493);
and U4704 (N_4704,N_4467,N_4539);
or U4705 (N_4705,N_4477,N_4597);
or U4706 (N_4706,N_4450,N_4461);
nand U4707 (N_4707,N_4542,N_4496);
or U4708 (N_4708,N_4504,N_4599);
xnor U4709 (N_4709,N_4401,N_4548);
and U4710 (N_4710,N_4552,N_4473);
and U4711 (N_4711,N_4578,N_4494);
nor U4712 (N_4712,N_4598,N_4489);
and U4713 (N_4713,N_4460,N_4506);
or U4714 (N_4714,N_4563,N_4528);
and U4715 (N_4715,N_4457,N_4448);
nor U4716 (N_4716,N_4573,N_4554);
or U4717 (N_4717,N_4450,N_4580);
or U4718 (N_4718,N_4451,N_4554);
xor U4719 (N_4719,N_4514,N_4525);
or U4720 (N_4720,N_4454,N_4493);
and U4721 (N_4721,N_4408,N_4414);
nand U4722 (N_4722,N_4593,N_4465);
nand U4723 (N_4723,N_4573,N_4582);
nor U4724 (N_4724,N_4463,N_4528);
nor U4725 (N_4725,N_4411,N_4544);
xor U4726 (N_4726,N_4486,N_4455);
or U4727 (N_4727,N_4500,N_4409);
nand U4728 (N_4728,N_4562,N_4573);
nor U4729 (N_4729,N_4460,N_4450);
nor U4730 (N_4730,N_4527,N_4582);
or U4731 (N_4731,N_4407,N_4450);
or U4732 (N_4732,N_4419,N_4586);
and U4733 (N_4733,N_4463,N_4438);
or U4734 (N_4734,N_4502,N_4477);
and U4735 (N_4735,N_4592,N_4490);
nor U4736 (N_4736,N_4531,N_4448);
and U4737 (N_4737,N_4423,N_4466);
nand U4738 (N_4738,N_4598,N_4464);
or U4739 (N_4739,N_4437,N_4562);
nor U4740 (N_4740,N_4557,N_4420);
xnor U4741 (N_4741,N_4544,N_4416);
nand U4742 (N_4742,N_4509,N_4558);
xnor U4743 (N_4743,N_4492,N_4536);
and U4744 (N_4744,N_4587,N_4469);
or U4745 (N_4745,N_4454,N_4464);
nand U4746 (N_4746,N_4589,N_4438);
nand U4747 (N_4747,N_4528,N_4534);
nor U4748 (N_4748,N_4513,N_4509);
or U4749 (N_4749,N_4522,N_4570);
nor U4750 (N_4750,N_4536,N_4549);
nor U4751 (N_4751,N_4492,N_4519);
xnor U4752 (N_4752,N_4517,N_4484);
nor U4753 (N_4753,N_4401,N_4572);
and U4754 (N_4754,N_4559,N_4456);
and U4755 (N_4755,N_4467,N_4576);
nand U4756 (N_4756,N_4555,N_4547);
or U4757 (N_4757,N_4543,N_4444);
nor U4758 (N_4758,N_4544,N_4539);
nor U4759 (N_4759,N_4548,N_4449);
xnor U4760 (N_4760,N_4503,N_4509);
or U4761 (N_4761,N_4499,N_4587);
or U4762 (N_4762,N_4535,N_4575);
and U4763 (N_4763,N_4500,N_4599);
and U4764 (N_4764,N_4458,N_4561);
nor U4765 (N_4765,N_4575,N_4492);
or U4766 (N_4766,N_4552,N_4402);
and U4767 (N_4767,N_4515,N_4453);
nand U4768 (N_4768,N_4533,N_4492);
nor U4769 (N_4769,N_4538,N_4581);
and U4770 (N_4770,N_4443,N_4502);
nand U4771 (N_4771,N_4568,N_4593);
or U4772 (N_4772,N_4515,N_4595);
and U4773 (N_4773,N_4423,N_4405);
or U4774 (N_4774,N_4522,N_4502);
and U4775 (N_4775,N_4543,N_4508);
xor U4776 (N_4776,N_4578,N_4411);
xor U4777 (N_4777,N_4584,N_4564);
or U4778 (N_4778,N_4458,N_4532);
and U4779 (N_4779,N_4422,N_4533);
and U4780 (N_4780,N_4585,N_4440);
and U4781 (N_4781,N_4459,N_4553);
nor U4782 (N_4782,N_4556,N_4430);
or U4783 (N_4783,N_4576,N_4406);
nor U4784 (N_4784,N_4561,N_4574);
and U4785 (N_4785,N_4406,N_4416);
or U4786 (N_4786,N_4594,N_4517);
nor U4787 (N_4787,N_4480,N_4575);
nor U4788 (N_4788,N_4474,N_4496);
nand U4789 (N_4789,N_4546,N_4516);
and U4790 (N_4790,N_4403,N_4437);
and U4791 (N_4791,N_4481,N_4577);
xor U4792 (N_4792,N_4408,N_4591);
and U4793 (N_4793,N_4457,N_4545);
nor U4794 (N_4794,N_4435,N_4592);
xnor U4795 (N_4795,N_4563,N_4557);
or U4796 (N_4796,N_4457,N_4585);
and U4797 (N_4797,N_4444,N_4555);
or U4798 (N_4798,N_4504,N_4513);
or U4799 (N_4799,N_4570,N_4533);
and U4800 (N_4800,N_4780,N_4768);
or U4801 (N_4801,N_4799,N_4644);
or U4802 (N_4802,N_4759,N_4600);
and U4803 (N_4803,N_4747,N_4674);
or U4804 (N_4804,N_4648,N_4642);
nand U4805 (N_4805,N_4766,N_4787);
or U4806 (N_4806,N_4686,N_4775);
nand U4807 (N_4807,N_4772,N_4630);
and U4808 (N_4808,N_4779,N_4667);
and U4809 (N_4809,N_4764,N_4632);
xnor U4810 (N_4810,N_4778,N_4774);
nand U4811 (N_4811,N_4635,N_4614);
nand U4812 (N_4812,N_4643,N_4797);
nor U4813 (N_4813,N_4784,N_4697);
nor U4814 (N_4814,N_4703,N_4633);
nand U4815 (N_4815,N_4628,N_4638);
xor U4816 (N_4816,N_4695,N_4657);
xnor U4817 (N_4817,N_4610,N_4711);
xor U4818 (N_4818,N_4704,N_4712);
nor U4819 (N_4819,N_4654,N_4636);
and U4820 (N_4820,N_4691,N_4730);
nand U4821 (N_4821,N_4660,N_4653);
or U4822 (N_4822,N_4692,N_4737);
and U4823 (N_4823,N_4791,N_4786);
or U4824 (N_4824,N_4716,N_4619);
or U4825 (N_4825,N_4662,N_4685);
nand U4826 (N_4826,N_4605,N_4656);
nor U4827 (N_4827,N_4668,N_4626);
xnor U4828 (N_4828,N_4678,N_4721);
and U4829 (N_4829,N_4706,N_4773);
or U4830 (N_4830,N_4677,N_4658);
nor U4831 (N_4831,N_4617,N_4713);
or U4832 (N_4832,N_4618,N_4794);
nor U4833 (N_4833,N_4620,N_4718);
nor U4834 (N_4834,N_4649,N_4680);
nand U4835 (N_4835,N_4696,N_4616);
nand U4836 (N_4836,N_4750,N_4792);
and U4837 (N_4837,N_4751,N_4769);
nor U4838 (N_4838,N_4723,N_4602);
or U4839 (N_4839,N_4702,N_4708);
and U4840 (N_4840,N_4758,N_4663);
or U4841 (N_4841,N_4763,N_4736);
or U4842 (N_4842,N_4623,N_4650);
nand U4843 (N_4843,N_4717,N_4735);
or U4844 (N_4844,N_4631,N_4611);
nand U4845 (N_4845,N_4661,N_4781);
and U4846 (N_4846,N_4762,N_4761);
or U4847 (N_4847,N_4771,N_4714);
and U4848 (N_4848,N_4613,N_4734);
or U4849 (N_4849,N_4744,N_4710);
nand U4850 (N_4850,N_4749,N_4720);
or U4851 (N_4851,N_4752,N_4679);
or U4852 (N_4852,N_4670,N_4690);
and U4853 (N_4853,N_4760,N_4682);
or U4854 (N_4854,N_4743,N_4757);
nand U4855 (N_4855,N_4789,N_4740);
and U4856 (N_4856,N_4637,N_4765);
nand U4857 (N_4857,N_4625,N_4639);
nor U4858 (N_4858,N_4683,N_4615);
or U4859 (N_4859,N_4609,N_4724);
or U4860 (N_4860,N_4673,N_4729);
or U4861 (N_4861,N_4688,N_4700);
nor U4862 (N_4862,N_4782,N_4606);
or U4863 (N_4863,N_4603,N_4627);
nand U4864 (N_4864,N_4742,N_4672);
nor U4865 (N_4865,N_4665,N_4741);
nor U4866 (N_4866,N_4640,N_4604);
xnor U4867 (N_4867,N_4728,N_4693);
xnor U4868 (N_4868,N_4790,N_4681);
and U4869 (N_4869,N_4698,N_4669);
nor U4870 (N_4870,N_4715,N_4755);
nand U4871 (N_4871,N_4659,N_4641);
and U4872 (N_4872,N_4666,N_4793);
nand U4873 (N_4873,N_4785,N_4612);
nor U4874 (N_4874,N_4651,N_4707);
and U4875 (N_4875,N_4745,N_4709);
and U4876 (N_4876,N_4689,N_4795);
or U4877 (N_4877,N_4687,N_4727);
or U4878 (N_4878,N_4607,N_4622);
xor U4879 (N_4879,N_4732,N_4748);
nand U4880 (N_4880,N_4753,N_4647);
xor U4881 (N_4881,N_4646,N_4756);
and U4882 (N_4882,N_4684,N_4731);
or U4883 (N_4883,N_4777,N_4754);
and U4884 (N_4884,N_4676,N_4776);
and U4885 (N_4885,N_4726,N_4699);
nor U4886 (N_4886,N_4621,N_4733);
nor U4887 (N_4887,N_4655,N_4664);
xor U4888 (N_4888,N_4796,N_4634);
or U4889 (N_4889,N_4652,N_4722);
and U4890 (N_4890,N_4645,N_4788);
or U4891 (N_4891,N_4705,N_4671);
or U4892 (N_4892,N_4746,N_4783);
nor U4893 (N_4893,N_4798,N_4767);
nor U4894 (N_4894,N_4738,N_4629);
and U4895 (N_4895,N_4719,N_4739);
nand U4896 (N_4896,N_4608,N_4624);
or U4897 (N_4897,N_4770,N_4701);
or U4898 (N_4898,N_4725,N_4675);
and U4899 (N_4899,N_4601,N_4694);
nor U4900 (N_4900,N_4601,N_4619);
and U4901 (N_4901,N_4791,N_4657);
or U4902 (N_4902,N_4648,N_4697);
or U4903 (N_4903,N_4703,N_4784);
and U4904 (N_4904,N_4722,N_4748);
or U4905 (N_4905,N_4606,N_4772);
xnor U4906 (N_4906,N_4756,N_4630);
nor U4907 (N_4907,N_4646,N_4681);
and U4908 (N_4908,N_4702,N_4733);
and U4909 (N_4909,N_4752,N_4740);
nor U4910 (N_4910,N_4748,N_4642);
and U4911 (N_4911,N_4788,N_4708);
nor U4912 (N_4912,N_4696,N_4613);
nor U4913 (N_4913,N_4740,N_4653);
or U4914 (N_4914,N_4625,N_4709);
nand U4915 (N_4915,N_4634,N_4620);
xnor U4916 (N_4916,N_4664,N_4755);
nand U4917 (N_4917,N_4749,N_4605);
nor U4918 (N_4918,N_4639,N_4736);
nand U4919 (N_4919,N_4701,N_4745);
and U4920 (N_4920,N_4606,N_4779);
nand U4921 (N_4921,N_4722,N_4736);
nand U4922 (N_4922,N_4696,N_4768);
or U4923 (N_4923,N_4691,N_4785);
or U4924 (N_4924,N_4656,N_4771);
xor U4925 (N_4925,N_4759,N_4782);
or U4926 (N_4926,N_4758,N_4605);
and U4927 (N_4927,N_4694,N_4765);
or U4928 (N_4928,N_4730,N_4707);
xor U4929 (N_4929,N_4729,N_4732);
nand U4930 (N_4930,N_4651,N_4645);
or U4931 (N_4931,N_4748,N_4764);
and U4932 (N_4932,N_4792,N_4612);
nand U4933 (N_4933,N_4658,N_4710);
nand U4934 (N_4934,N_4744,N_4645);
nand U4935 (N_4935,N_4632,N_4758);
and U4936 (N_4936,N_4689,N_4785);
nor U4937 (N_4937,N_4607,N_4787);
and U4938 (N_4938,N_4738,N_4693);
nor U4939 (N_4939,N_4736,N_4625);
or U4940 (N_4940,N_4677,N_4671);
nor U4941 (N_4941,N_4780,N_4766);
or U4942 (N_4942,N_4632,N_4607);
or U4943 (N_4943,N_4742,N_4650);
nand U4944 (N_4944,N_4795,N_4608);
or U4945 (N_4945,N_4679,N_4756);
nand U4946 (N_4946,N_4728,N_4611);
nor U4947 (N_4947,N_4602,N_4658);
nand U4948 (N_4948,N_4721,N_4610);
and U4949 (N_4949,N_4792,N_4649);
nor U4950 (N_4950,N_4743,N_4698);
nor U4951 (N_4951,N_4673,N_4638);
and U4952 (N_4952,N_4633,N_4662);
and U4953 (N_4953,N_4712,N_4606);
nor U4954 (N_4954,N_4678,N_4684);
nand U4955 (N_4955,N_4687,N_4735);
or U4956 (N_4956,N_4606,N_4665);
and U4957 (N_4957,N_4749,N_4684);
xnor U4958 (N_4958,N_4785,N_4714);
nor U4959 (N_4959,N_4793,N_4677);
and U4960 (N_4960,N_4769,N_4631);
or U4961 (N_4961,N_4627,N_4716);
nand U4962 (N_4962,N_4735,N_4694);
and U4963 (N_4963,N_4650,N_4695);
or U4964 (N_4964,N_4799,N_4786);
and U4965 (N_4965,N_4628,N_4781);
nand U4966 (N_4966,N_4761,N_4707);
and U4967 (N_4967,N_4688,N_4672);
and U4968 (N_4968,N_4657,N_4750);
nor U4969 (N_4969,N_4747,N_4709);
or U4970 (N_4970,N_4681,N_4771);
nor U4971 (N_4971,N_4766,N_4747);
and U4972 (N_4972,N_4655,N_4611);
nor U4973 (N_4973,N_4667,N_4723);
nand U4974 (N_4974,N_4643,N_4786);
nor U4975 (N_4975,N_4790,N_4794);
and U4976 (N_4976,N_4767,N_4771);
nor U4977 (N_4977,N_4684,N_4630);
nor U4978 (N_4978,N_4788,N_4674);
nand U4979 (N_4979,N_4726,N_4666);
nor U4980 (N_4980,N_4635,N_4609);
and U4981 (N_4981,N_4634,N_4636);
and U4982 (N_4982,N_4710,N_4789);
or U4983 (N_4983,N_4674,N_4704);
nor U4984 (N_4984,N_4663,N_4667);
nand U4985 (N_4985,N_4790,N_4662);
nand U4986 (N_4986,N_4731,N_4683);
nor U4987 (N_4987,N_4695,N_4769);
nor U4988 (N_4988,N_4724,N_4730);
xor U4989 (N_4989,N_4607,N_4698);
nand U4990 (N_4990,N_4641,N_4679);
nand U4991 (N_4991,N_4647,N_4649);
nand U4992 (N_4992,N_4651,N_4740);
nand U4993 (N_4993,N_4663,N_4687);
and U4994 (N_4994,N_4671,N_4757);
or U4995 (N_4995,N_4607,N_4683);
nand U4996 (N_4996,N_4604,N_4790);
nor U4997 (N_4997,N_4778,N_4684);
nand U4998 (N_4998,N_4696,N_4633);
and U4999 (N_4999,N_4673,N_4736);
or UO_0 (O_0,N_4876,N_4984);
nand UO_1 (O_1,N_4900,N_4867);
nand UO_2 (O_2,N_4994,N_4831);
nor UO_3 (O_3,N_4904,N_4998);
xnor UO_4 (O_4,N_4987,N_4850);
nand UO_5 (O_5,N_4883,N_4929);
or UO_6 (O_6,N_4825,N_4974);
or UO_7 (O_7,N_4881,N_4909);
and UO_8 (O_8,N_4912,N_4859);
nor UO_9 (O_9,N_4950,N_4840);
and UO_10 (O_10,N_4873,N_4868);
nor UO_11 (O_11,N_4924,N_4821);
and UO_12 (O_12,N_4939,N_4990);
nor UO_13 (O_13,N_4954,N_4870);
nand UO_14 (O_14,N_4886,N_4852);
nand UO_15 (O_15,N_4996,N_4809);
or UO_16 (O_16,N_4862,N_4969);
nand UO_17 (O_17,N_4874,N_4986);
or UO_18 (O_18,N_4884,N_4894);
or UO_19 (O_19,N_4813,N_4871);
nor UO_20 (O_20,N_4967,N_4846);
or UO_21 (O_21,N_4982,N_4963);
nor UO_22 (O_22,N_4962,N_4952);
and UO_23 (O_23,N_4949,N_4922);
xnor UO_24 (O_24,N_4824,N_4838);
nor UO_25 (O_25,N_4977,N_4810);
nor UO_26 (O_26,N_4842,N_4851);
nor UO_27 (O_27,N_4913,N_4864);
or UO_28 (O_28,N_4923,N_4802);
nor UO_29 (O_29,N_4832,N_4897);
nand UO_30 (O_30,N_4892,N_4828);
or UO_31 (O_31,N_4803,N_4866);
nand UO_32 (O_32,N_4855,N_4889);
nor UO_33 (O_33,N_4878,N_4822);
or UO_34 (O_34,N_4863,N_4818);
nand UO_35 (O_35,N_4845,N_4961);
xnor UO_36 (O_36,N_4826,N_4861);
nand UO_37 (O_37,N_4941,N_4905);
or UO_38 (O_38,N_4916,N_4971);
and UO_39 (O_39,N_4919,N_4808);
or UO_40 (O_40,N_4958,N_4978);
xor UO_41 (O_41,N_4860,N_4956);
xor UO_42 (O_42,N_4898,N_4848);
nand UO_43 (O_43,N_4953,N_4983);
and UO_44 (O_44,N_4937,N_4926);
or UO_45 (O_45,N_4899,N_4968);
nor UO_46 (O_46,N_4921,N_4807);
nand UO_47 (O_47,N_4887,N_4833);
nand UO_48 (O_48,N_4877,N_4829);
xor UO_49 (O_49,N_4975,N_4819);
or UO_50 (O_50,N_4981,N_4865);
or UO_51 (O_51,N_4917,N_4811);
or UO_52 (O_52,N_4928,N_4918);
or UO_53 (O_53,N_4935,N_4925);
xnor UO_54 (O_54,N_4895,N_4903);
and UO_55 (O_55,N_4902,N_4827);
xnor UO_56 (O_56,N_4875,N_4965);
xnor UO_57 (O_57,N_4948,N_4991);
nand UO_58 (O_58,N_4814,N_4801);
or UO_59 (O_59,N_4943,N_4959);
and UO_60 (O_60,N_4988,N_4896);
and UO_61 (O_61,N_4933,N_4955);
and UO_62 (O_62,N_4927,N_4976);
or UO_63 (O_63,N_4907,N_4979);
or UO_64 (O_64,N_4853,N_4880);
or UO_65 (O_65,N_4815,N_4869);
nor UO_66 (O_66,N_4920,N_4938);
nand UO_67 (O_67,N_4957,N_4901);
and UO_68 (O_68,N_4942,N_4970);
or UO_69 (O_69,N_4932,N_4995);
nand UO_70 (O_70,N_4843,N_4985);
nor UO_71 (O_71,N_4966,N_4854);
or UO_72 (O_72,N_4945,N_4817);
or UO_73 (O_73,N_4946,N_4836);
and UO_74 (O_74,N_4890,N_4972);
and UO_75 (O_75,N_4882,N_4804);
nor UO_76 (O_76,N_4891,N_4879);
or UO_77 (O_77,N_4847,N_4888);
or UO_78 (O_78,N_4911,N_4980);
nand UO_79 (O_79,N_4931,N_4857);
nand UO_80 (O_80,N_4858,N_4930);
nor UO_81 (O_81,N_4936,N_4841);
nor UO_82 (O_82,N_4960,N_4837);
and UO_83 (O_83,N_4915,N_4906);
xor UO_84 (O_84,N_4934,N_4835);
and UO_85 (O_85,N_4951,N_4856);
and UO_86 (O_86,N_4820,N_4834);
nand UO_87 (O_87,N_4806,N_4823);
nor UO_88 (O_88,N_4944,N_4908);
nor UO_89 (O_89,N_4844,N_4893);
nand UO_90 (O_90,N_4914,N_4805);
or UO_91 (O_91,N_4992,N_4947);
xnor UO_92 (O_92,N_4973,N_4997);
and UO_93 (O_93,N_4940,N_4993);
nand UO_94 (O_94,N_4910,N_4999);
and UO_95 (O_95,N_4885,N_4830);
or UO_96 (O_96,N_4800,N_4849);
nand UO_97 (O_97,N_4872,N_4816);
nand UO_98 (O_98,N_4839,N_4989);
and UO_99 (O_99,N_4812,N_4964);
or UO_100 (O_100,N_4935,N_4894);
or UO_101 (O_101,N_4835,N_4862);
nand UO_102 (O_102,N_4926,N_4952);
and UO_103 (O_103,N_4939,N_4830);
nand UO_104 (O_104,N_4980,N_4997);
nand UO_105 (O_105,N_4869,N_4832);
nor UO_106 (O_106,N_4839,N_4914);
and UO_107 (O_107,N_4893,N_4919);
or UO_108 (O_108,N_4931,N_4905);
and UO_109 (O_109,N_4924,N_4803);
nor UO_110 (O_110,N_4953,N_4995);
and UO_111 (O_111,N_4812,N_4930);
and UO_112 (O_112,N_4983,N_4986);
nor UO_113 (O_113,N_4872,N_4850);
nand UO_114 (O_114,N_4993,N_4872);
or UO_115 (O_115,N_4874,N_4993);
and UO_116 (O_116,N_4924,N_4903);
nor UO_117 (O_117,N_4886,N_4806);
and UO_118 (O_118,N_4976,N_4937);
or UO_119 (O_119,N_4851,N_4989);
and UO_120 (O_120,N_4827,N_4993);
xor UO_121 (O_121,N_4920,N_4963);
nand UO_122 (O_122,N_4844,N_4915);
nor UO_123 (O_123,N_4991,N_4871);
and UO_124 (O_124,N_4801,N_4963);
nor UO_125 (O_125,N_4823,N_4811);
xor UO_126 (O_126,N_4936,N_4937);
or UO_127 (O_127,N_4857,N_4842);
and UO_128 (O_128,N_4828,N_4929);
nor UO_129 (O_129,N_4900,N_4862);
and UO_130 (O_130,N_4840,N_4831);
and UO_131 (O_131,N_4968,N_4849);
and UO_132 (O_132,N_4824,N_4989);
xor UO_133 (O_133,N_4817,N_4874);
and UO_134 (O_134,N_4922,N_4935);
xor UO_135 (O_135,N_4842,N_4973);
or UO_136 (O_136,N_4845,N_4928);
nor UO_137 (O_137,N_4840,N_4804);
or UO_138 (O_138,N_4980,N_4837);
and UO_139 (O_139,N_4949,N_4873);
and UO_140 (O_140,N_4950,N_4979);
nor UO_141 (O_141,N_4940,N_4936);
and UO_142 (O_142,N_4845,N_4912);
or UO_143 (O_143,N_4921,N_4827);
and UO_144 (O_144,N_4821,N_4945);
and UO_145 (O_145,N_4815,N_4921);
and UO_146 (O_146,N_4933,N_4848);
or UO_147 (O_147,N_4850,N_4978);
nand UO_148 (O_148,N_4803,N_4819);
or UO_149 (O_149,N_4827,N_4879);
nand UO_150 (O_150,N_4807,N_4914);
and UO_151 (O_151,N_4990,N_4846);
and UO_152 (O_152,N_4986,N_4817);
nor UO_153 (O_153,N_4966,N_4881);
or UO_154 (O_154,N_4952,N_4905);
or UO_155 (O_155,N_4938,N_4916);
nor UO_156 (O_156,N_4854,N_4839);
xnor UO_157 (O_157,N_4905,N_4918);
nor UO_158 (O_158,N_4819,N_4943);
xnor UO_159 (O_159,N_4820,N_4939);
nor UO_160 (O_160,N_4815,N_4843);
nor UO_161 (O_161,N_4902,N_4921);
xor UO_162 (O_162,N_4837,N_4842);
and UO_163 (O_163,N_4899,N_4915);
nand UO_164 (O_164,N_4935,N_4999);
nand UO_165 (O_165,N_4981,N_4878);
and UO_166 (O_166,N_4897,N_4902);
nor UO_167 (O_167,N_4869,N_4998);
xnor UO_168 (O_168,N_4824,N_4879);
and UO_169 (O_169,N_4919,N_4951);
nor UO_170 (O_170,N_4831,N_4865);
or UO_171 (O_171,N_4943,N_4956);
or UO_172 (O_172,N_4838,N_4877);
and UO_173 (O_173,N_4989,N_4818);
nand UO_174 (O_174,N_4858,N_4971);
nand UO_175 (O_175,N_4929,N_4990);
and UO_176 (O_176,N_4847,N_4940);
or UO_177 (O_177,N_4929,N_4942);
xnor UO_178 (O_178,N_4939,N_4985);
nor UO_179 (O_179,N_4922,N_4861);
and UO_180 (O_180,N_4964,N_4867);
nand UO_181 (O_181,N_4953,N_4982);
nor UO_182 (O_182,N_4912,N_4880);
or UO_183 (O_183,N_4904,N_4867);
nor UO_184 (O_184,N_4836,N_4952);
xnor UO_185 (O_185,N_4946,N_4892);
or UO_186 (O_186,N_4892,N_4887);
and UO_187 (O_187,N_4978,N_4881);
nand UO_188 (O_188,N_4914,N_4829);
and UO_189 (O_189,N_4959,N_4871);
nand UO_190 (O_190,N_4937,N_4961);
and UO_191 (O_191,N_4826,N_4834);
and UO_192 (O_192,N_4805,N_4930);
nand UO_193 (O_193,N_4984,N_4928);
nor UO_194 (O_194,N_4847,N_4891);
nor UO_195 (O_195,N_4931,N_4871);
nor UO_196 (O_196,N_4963,N_4872);
or UO_197 (O_197,N_4896,N_4901);
or UO_198 (O_198,N_4961,N_4938);
nor UO_199 (O_199,N_4824,N_4930);
xnor UO_200 (O_200,N_4855,N_4877);
nand UO_201 (O_201,N_4872,N_4949);
or UO_202 (O_202,N_4969,N_4922);
nand UO_203 (O_203,N_4876,N_4815);
nor UO_204 (O_204,N_4937,N_4898);
nor UO_205 (O_205,N_4941,N_4901);
nand UO_206 (O_206,N_4896,N_4854);
or UO_207 (O_207,N_4820,N_4969);
and UO_208 (O_208,N_4975,N_4856);
and UO_209 (O_209,N_4844,N_4905);
and UO_210 (O_210,N_4953,N_4822);
and UO_211 (O_211,N_4916,N_4886);
or UO_212 (O_212,N_4878,N_4871);
nor UO_213 (O_213,N_4889,N_4899);
nor UO_214 (O_214,N_4913,N_4917);
nand UO_215 (O_215,N_4973,N_4834);
xor UO_216 (O_216,N_4943,N_4885);
and UO_217 (O_217,N_4951,N_4846);
nor UO_218 (O_218,N_4861,N_4819);
nor UO_219 (O_219,N_4900,N_4803);
or UO_220 (O_220,N_4987,N_4983);
nand UO_221 (O_221,N_4861,N_4894);
xor UO_222 (O_222,N_4826,N_4812);
or UO_223 (O_223,N_4827,N_4806);
nor UO_224 (O_224,N_4970,N_4921);
nand UO_225 (O_225,N_4873,N_4822);
nor UO_226 (O_226,N_4840,N_4877);
nor UO_227 (O_227,N_4981,N_4851);
nand UO_228 (O_228,N_4959,N_4954);
or UO_229 (O_229,N_4983,N_4973);
nor UO_230 (O_230,N_4901,N_4984);
nand UO_231 (O_231,N_4941,N_4870);
nor UO_232 (O_232,N_4872,N_4942);
or UO_233 (O_233,N_4984,N_4872);
nor UO_234 (O_234,N_4969,N_4937);
nand UO_235 (O_235,N_4997,N_4802);
and UO_236 (O_236,N_4855,N_4993);
and UO_237 (O_237,N_4861,N_4803);
xnor UO_238 (O_238,N_4937,N_4995);
or UO_239 (O_239,N_4818,N_4944);
nor UO_240 (O_240,N_4883,N_4845);
xnor UO_241 (O_241,N_4870,N_4835);
and UO_242 (O_242,N_4838,N_4976);
xor UO_243 (O_243,N_4910,N_4873);
nor UO_244 (O_244,N_4968,N_4845);
or UO_245 (O_245,N_4850,N_4956);
or UO_246 (O_246,N_4928,N_4865);
or UO_247 (O_247,N_4820,N_4929);
or UO_248 (O_248,N_4993,N_4913);
or UO_249 (O_249,N_4802,N_4817);
nand UO_250 (O_250,N_4918,N_4992);
nand UO_251 (O_251,N_4839,N_4918);
and UO_252 (O_252,N_4801,N_4897);
or UO_253 (O_253,N_4993,N_4932);
and UO_254 (O_254,N_4982,N_4909);
or UO_255 (O_255,N_4835,N_4816);
nand UO_256 (O_256,N_4832,N_4929);
nor UO_257 (O_257,N_4922,N_4818);
nand UO_258 (O_258,N_4882,N_4957);
and UO_259 (O_259,N_4971,N_4804);
xnor UO_260 (O_260,N_4852,N_4929);
or UO_261 (O_261,N_4824,N_4856);
nor UO_262 (O_262,N_4830,N_4841);
and UO_263 (O_263,N_4881,N_4993);
nand UO_264 (O_264,N_4922,N_4842);
or UO_265 (O_265,N_4904,N_4846);
and UO_266 (O_266,N_4970,N_4909);
nor UO_267 (O_267,N_4800,N_4945);
nor UO_268 (O_268,N_4936,N_4828);
or UO_269 (O_269,N_4906,N_4803);
and UO_270 (O_270,N_4857,N_4863);
or UO_271 (O_271,N_4945,N_4832);
and UO_272 (O_272,N_4957,N_4855);
nand UO_273 (O_273,N_4975,N_4907);
and UO_274 (O_274,N_4936,N_4873);
or UO_275 (O_275,N_4876,N_4987);
xnor UO_276 (O_276,N_4954,N_4935);
nand UO_277 (O_277,N_4961,N_4997);
nand UO_278 (O_278,N_4902,N_4819);
nor UO_279 (O_279,N_4859,N_4926);
nand UO_280 (O_280,N_4816,N_4962);
nand UO_281 (O_281,N_4902,N_4890);
and UO_282 (O_282,N_4931,N_4824);
nand UO_283 (O_283,N_4894,N_4939);
nand UO_284 (O_284,N_4978,N_4892);
or UO_285 (O_285,N_4997,N_4993);
nand UO_286 (O_286,N_4833,N_4938);
or UO_287 (O_287,N_4889,N_4948);
or UO_288 (O_288,N_4811,N_4840);
and UO_289 (O_289,N_4970,N_4889);
and UO_290 (O_290,N_4825,N_4932);
nand UO_291 (O_291,N_4807,N_4901);
or UO_292 (O_292,N_4823,N_4973);
xnor UO_293 (O_293,N_4974,N_4876);
and UO_294 (O_294,N_4800,N_4958);
nor UO_295 (O_295,N_4843,N_4911);
nor UO_296 (O_296,N_4885,N_4871);
or UO_297 (O_297,N_4839,N_4846);
or UO_298 (O_298,N_4815,N_4986);
and UO_299 (O_299,N_4933,N_4954);
and UO_300 (O_300,N_4886,N_4957);
nand UO_301 (O_301,N_4809,N_4995);
or UO_302 (O_302,N_4806,N_4845);
nor UO_303 (O_303,N_4981,N_4913);
nor UO_304 (O_304,N_4839,N_4921);
or UO_305 (O_305,N_4967,N_4944);
or UO_306 (O_306,N_4912,N_4809);
nand UO_307 (O_307,N_4924,N_4920);
nand UO_308 (O_308,N_4998,N_4992);
or UO_309 (O_309,N_4847,N_4968);
nor UO_310 (O_310,N_4823,N_4915);
nand UO_311 (O_311,N_4803,N_4961);
and UO_312 (O_312,N_4962,N_4968);
and UO_313 (O_313,N_4846,N_4968);
nand UO_314 (O_314,N_4978,N_4961);
nor UO_315 (O_315,N_4885,N_4854);
nand UO_316 (O_316,N_4929,N_4928);
or UO_317 (O_317,N_4816,N_4802);
nand UO_318 (O_318,N_4974,N_4827);
and UO_319 (O_319,N_4892,N_4941);
or UO_320 (O_320,N_4903,N_4928);
nor UO_321 (O_321,N_4961,N_4988);
xor UO_322 (O_322,N_4808,N_4823);
nand UO_323 (O_323,N_4988,N_4986);
nand UO_324 (O_324,N_4938,N_4933);
or UO_325 (O_325,N_4892,N_4995);
and UO_326 (O_326,N_4939,N_4973);
nand UO_327 (O_327,N_4853,N_4960);
or UO_328 (O_328,N_4830,N_4917);
or UO_329 (O_329,N_4990,N_4924);
xor UO_330 (O_330,N_4907,N_4984);
nand UO_331 (O_331,N_4993,N_4969);
nand UO_332 (O_332,N_4968,N_4999);
nor UO_333 (O_333,N_4881,N_4945);
and UO_334 (O_334,N_4938,N_4980);
nor UO_335 (O_335,N_4831,N_4898);
and UO_336 (O_336,N_4929,N_4879);
nor UO_337 (O_337,N_4970,N_4926);
and UO_338 (O_338,N_4820,N_4918);
and UO_339 (O_339,N_4958,N_4848);
nand UO_340 (O_340,N_4967,N_4988);
nand UO_341 (O_341,N_4933,N_4835);
nor UO_342 (O_342,N_4802,N_4939);
xor UO_343 (O_343,N_4906,N_4817);
and UO_344 (O_344,N_4805,N_4828);
and UO_345 (O_345,N_4806,N_4818);
nor UO_346 (O_346,N_4980,N_4840);
nand UO_347 (O_347,N_4838,N_4981);
nand UO_348 (O_348,N_4817,N_4882);
xor UO_349 (O_349,N_4907,N_4827);
nand UO_350 (O_350,N_4817,N_4948);
and UO_351 (O_351,N_4881,N_4803);
xor UO_352 (O_352,N_4959,N_4849);
and UO_353 (O_353,N_4932,N_4909);
and UO_354 (O_354,N_4900,N_4958);
or UO_355 (O_355,N_4925,N_4955);
or UO_356 (O_356,N_4811,N_4926);
and UO_357 (O_357,N_4882,N_4849);
or UO_358 (O_358,N_4875,N_4932);
nor UO_359 (O_359,N_4956,N_4893);
xnor UO_360 (O_360,N_4999,N_4878);
xnor UO_361 (O_361,N_4976,N_4969);
nand UO_362 (O_362,N_4833,N_4930);
or UO_363 (O_363,N_4825,N_4976);
or UO_364 (O_364,N_4906,N_4878);
nand UO_365 (O_365,N_4934,N_4851);
xor UO_366 (O_366,N_4836,N_4827);
or UO_367 (O_367,N_4949,N_4939);
xnor UO_368 (O_368,N_4868,N_4995);
nand UO_369 (O_369,N_4883,N_4884);
nand UO_370 (O_370,N_4870,N_4807);
and UO_371 (O_371,N_4913,N_4869);
nand UO_372 (O_372,N_4825,N_4807);
nor UO_373 (O_373,N_4802,N_4958);
nor UO_374 (O_374,N_4893,N_4951);
or UO_375 (O_375,N_4985,N_4965);
nor UO_376 (O_376,N_4933,N_4929);
and UO_377 (O_377,N_4857,N_4925);
nand UO_378 (O_378,N_4970,N_4900);
nand UO_379 (O_379,N_4846,N_4920);
and UO_380 (O_380,N_4967,N_4977);
nand UO_381 (O_381,N_4954,N_4880);
nor UO_382 (O_382,N_4854,N_4871);
nor UO_383 (O_383,N_4823,N_4940);
nand UO_384 (O_384,N_4832,N_4890);
xor UO_385 (O_385,N_4809,N_4993);
and UO_386 (O_386,N_4822,N_4946);
or UO_387 (O_387,N_4953,N_4907);
xor UO_388 (O_388,N_4851,N_4845);
nand UO_389 (O_389,N_4985,N_4966);
and UO_390 (O_390,N_4884,N_4895);
or UO_391 (O_391,N_4991,N_4970);
xnor UO_392 (O_392,N_4985,N_4886);
or UO_393 (O_393,N_4814,N_4865);
or UO_394 (O_394,N_4998,N_4997);
or UO_395 (O_395,N_4866,N_4830);
nor UO_396 (O_396,N_4916,N_4811);
and UO_397 (O_397,N_4910,N_4949);
nor UO_398 (O_398,N_4941,N_4921);
and UO_399 (O_399,N_4924,N_4808);
nand UO_400 (O_400,N_4922,N_4929);
or UO_401 (O_401,N_4986,N_4902);
nor UO_402 (O_402,N_4905,N_4804);
or UO_403 (O_403,N_4801,N_4833);
and UO_404 (O_404,N_4819,N_4989);
or UO_405 (O_405,N_4803,N_4988);
or UO_406 (O_406,N_4849,N_4892);
nor UO_407 (O_407,N_4820,N_4922);
and UO_408 (O_408,N_4950,N_4868);
nand UO_409 (O_409,N_4975,N_4977);
or UO_410 (O_410,N_4844,N_4958);
nor UO_411 (O_411,N_4954,N_4860);
xor UO_412 (O_412,N_4966,N_4901);
or UO_413 (O_413,N_4931,N_4962);
nor UO_414 (O_414,N_4902,N_4860);
nor UO_415 (O_415,N_4954,N_4842);
or UO_416 (O_416,N_4898,N_4882);
xnor UO_417 (O_417,N_4950,N_4814);
nor UO_418 (O_418,N_4966,N_4808);
or UO_419 (O_419,N_4953,N_4824);
nor UO_420 (O_420,N_4999,N_4946);
and UO_421 (O_421,N_4950,N_4931);
or UO_422 (O_422,N_4874,N_4847);
or UO_423 (O_423,N_4852,N_4944);
nor UO_424 (O_424,N_4916,N_4889);
xnor UO_425 (O_425,N_4834,N_4928);
nor UO_426 (O_426,N_4957,N_4946);
and UO_427 (O_427,N_4875,N_4991);
and UO_428 (O_428,N_4938,N_4874);
or UO_429 (O_429,N_4885,N_4941);
nor UO_430 (O_430,N_4956,N_4809);
nor UO_431 (O_431,N_4894,N_4858);
and UO_432 (O_432,N_4965,N_4842);
and UO_433 (O_433,N_4822,N_4875);
or UO_434 (O_434,N_4849,N_4924);
xnor UO_435 (O_435,N_4935,N_4845);
nand UO_436 (O_436,N_4881,N_4916);
nor UO_437 (O_437,N_4894,N_4908);
nor UO_438 (O_438,N_4816,N_4970);
nor UO_439 (O_439,N_4919,N_4894);
nor UO_440 (O_440,N_4914,N_4888);
nor UO_441 (O_441,N_4804,N_4899);
nand UO_442 (O_442,N_4851,N_4920);
nor UO_443 (O_443,N_4874,N_4827);
nor UO_444 (O_444,N_4949,N_4810);
nor UO_445 (O_445,N_4888,N_4861);
nor UO_446 (O_446,N_4931,N_4995);
and UO_447 (O_447,N_4974,N_4886);
and UO_448 (O_448,N_4896,N_4830);
nand UO_449 (O_449,N_4824,N_4832);
or UO_450 (O_450,N_4886,N_4826);
nor UO_451 (O_451,N_4944,N_4928);
or UO_452 (O_452,N_4915,N_4835);
or UO_453 (O_453,N_4828,N_4807);
nor UO_454 (O_454,N_4892,N_4920);
xor UO_455 (O_455,N_4911,N_4936);
and UO_456 (O_456,N_4838,N_4935);
nor UO_457 (O_457,N_4976,N_4857);
xnor UO_458 (O_458,N_4962,N_4882);
xor UO_459 (O_459,N_4838,N_4936);
and UO_460 (O_460,N_4980,N_4993);
or UO_461 (O_461,N_4811,N_4857);
or UO_462 (O_462,N_4908,N_4825);
or UO_463 (O_463,N_4866,N_4919);
xor UO_464 (O_464,N_4992,N_4991);
nor UO_465 (O_465,N_4873,N_4887);
nand UO_466 (O_466,N_4966,N_4821);
xor UO_467 (O_467,N_4816,N_4981);
or UO_468 (O_468,N_4953,N_4949);
or UO_469 (O_469,N_4955,N_4956);
nor UO_470 (O_470,N_4900,N_4804);
or UO_471 (O_471,N_4938,N_4831);
and UO_472 (O_472,N_4847,N_4970);
nand UO_473 (O_473,N_4827,N_4878);
or UO_474 (O_474,N_4887,N_4967);
nor UO_475 (O_475,N_4956,N_4848);
nor UO_476 (O_476,N_4947,N_4955);
nor UO_477 (O_477,N_4926,N_4863);
and UO_478 (O_478,N_4956,N_4916);
and UO_479 (O_479,N_4989,N_4942);
and UO_480 (O_480,N_4860,N_4979);
nor UO_481 (O_481,N_4821,N_4968);
nor UO_482 (O_482,N_4992,N_4980);
nand UO_483 (O_483,N_4890,N_4957);
or UO_484 (O_484,N_4809,N_4806);
or UO_485 (O_485,N_4983,N_4940);
xnor UO_486 (O_486,N_4943,N_4802);
nand UO_487 (O_487,N_4845,N_4856);
nor UO_488 (O_488,N_4827,N_4891);
and UO_489 (O_489,N_4876,N_4962);
and UO_490 (O_490,N_4884,N_4827);
nor UO_491 (O_491,N_4877,N_4979);
and UO_492 (O_492,N_4865,N_4916);
xnor UO_493 (O_493,N_4880,N_4827);
or UO_494 (O_494,N_4914,N_4875);
or UO_495 (O_495,N_4981,N_4899);
or UO_496 (O_496,N_4872,N_4841);
nand UO_497 (O_497,N_4819,N_4999);
and UO_498 (O_498,N_4947,N_4911);
or UO_499 (O_499,N_4867,N_4997);
nand UO_500 (O_500,N_4820,N_4977);
nor UO_501 (O_501,N_4899,N_4898);
and UO_502 (O_502,N_4837,N_4901);
xnor UO_503 (O_503,N_4962,N_4834);
or UO_504 (O_504,N_4968,N_4823);
nor UO_505 (O_505,N_4827,N_4818);
or UO_506 (O_506,N_4992,N_4883);
nor UO_507 (O_507,N_4926,N_4823);
or UO_508 (O_508,N_4876,N_4990);
nand UO_509 (O_509,N_4945,N_4880);
xnor UO_510 (O_510,N_4805,N_4863);
nor UO_511 (O_511,N_4868,N_4837);
nand UO_512 (O_512,N_4926,N_4879);
and UO_513 (O_513,N_4857,N_4898);
nand UO_514 (O_514,N_4889,N_4915);
nor UO_515 (O_515,N_4994,N_4889);
and UO_516 (O_516,N_4911,N_4833);
nor UO_517 (O_517,N_4967,N_4927);
xnor UO_518 (O_518,N_4926,N_4819);
and UO_519 (O_519,N_4926,N_4808);
or UO_520 (O_520,N_4820,N_4961);
or UO_521 (O_521,N_4809,N_4951);
nand UO_522 (O_522,N_4887,N_4931);
nor UO_523 (O_523,N_4980,N_4897);
xor UO_524 (O_524,N_4826,N_4864);
nor UO_525 (O_525,N_4973,N_4844);
nand UO_526 (O_526,N_4918,N_4960);
nand UO_527 (O_527,N_4939,N_4891);
and UO_528 (O_528,N_4842,N_4960);
nor UO_529 (O_529,N_4849,N_4864);
or UO_530 (O_530,N_4948,N_4852);
or UO_531 (O_531,N_4915,N_4969);
and UO_532 (O_532,N_4889,N_4888);
nand UO_533 (O_533,N_4862,N_4846);
or UO_534 (O_534,N_4955,N_4837);
and UO_535 (O_535,N_4884,N_4944);
nand UO_536 (O_536,N_4824,N_4837);
xor UO_537 (O_537,N_4987,N_4813);
xor UO_538 (O_538,N_4962,N_4910);
xnor UO_539 (O_539,N_4910,N_4972);
and UO_540 (O_540,N_4914,N_4854);
or UO_541 (O_541,N_4832,N_4863);
or UO_542 (O_542,N_4927,N_4855);
and UO_543 (O_543,N_4899,N_4905);
nor UO_544 (O_544,N_4859,N_4956);
nand UO_545 (O_545,N_4842,N_4935);
and UO_546 (O_546,N_4966,N_4825);
xor UO_547 (O_547,N_4826,N_4871);
nor UO_548 (O_548,N_4920,N_4935);
and UO_549 (O_549,N_4848,N_4814);
nor UO_550 (O_550,N_4939,N_4991);
xor UO_551 (O_551,N_4811,N_4978);
nand UO_552 (O_552,N_4911,N_4841);
and UO_553 (O_553,N_4901,N_4820);
nand UO_554 (O_554,N_4997,N_4838);
nand UO_555 (O_555,N_4814,N_4843);
nor UO_556 (O_556,N_4904,N_4815);
xnor UO_557 (O_557,N_4945,N_4919);
and UO_558 (O_558,N_4832,N_4875);
and UO_559 (O_559,N_4987,N_4885);
nor UO_560 (O_560,N_4916,N_4914);
nand UO_561 (O_561,N_4871,N_4960);
nand UO_562 (O_562,N_4839,N_4937);
or UO_563 (O_563,N_4898,N_4885);
or UO_564 (O_564,N_4898,N_4809);
nand UO_565 (O_565,N_4896,N_4870);
nor UO_566 (O_566,N_4971,N_4932);
nand UO_567 (O_567,N_4917,N_4989);
xnor UO_568 (O_568,N_4992,N_4898);
and UO_569 (O_569,N_4887,N_4902);
xor UO_570 (O_570,N_4985,N_4837);
xor UO_571 (O_571,N_4854,N_4987);
nor UO_572 (O_572,N_4973,N_4930);
and UO_573 (O_573,N_4859,N_4891);
nor UO_574 (O_574,N_4892,N_4811);
and UO_575 (O_575,N_4982,N_4918);
nand UO_576 (O_576,N_4955,N_4904);
or UO_577 (O_577,N_4913,N_4854);
nor UO_578 (O_578,N_4954,N_4885);
and UO_579 (O_579,N_4996,N_4818);
or UO_580 (O_580,N_4841,N_4955);
nor UO_581 (O_581,N_4983,N_4850);
or UO_582 (O_582,N_4889,N_4911);
or UO_583 (O_583,N_4893,N_4947);
nand UO_584 (O_584,N_4960,N_4846);
or UO_585 (O_585,N_4881,N_4855);
nor UO_586 (O_586,N_4847,N_4832);
and UO_587 (O_587,N_4897,N_4997);
and UO_588 (O_588,N_4823,N_4904);
nand UO_589 (O_589,N_4958,N_4969);
or UO_590 (O_590,N_4938,N_4861);
nand UO_591 (O_591,N_4940,N_4826);
or UO_592 (O_592,N_4919,N_4805);
nor UO_593 (O_593,N_4841,N_4831);
and UO_594 (O_594,N_4886,N_4801);
and UO_595 (O_595,N_4905,N_4935);
xnor UO_596 (O_596,N_4966,N_4852);
nand UO_597 (O_597,N_4870,N_4921);
or UO_598 (O_598,N_4904,N_4810);
or UO_599 (O_599,N_4998,N_4876);
nor UO_600 (O_600,N_4969,N_4806);
and UO_601 (O_601,N_4844,N_4957);
nor UO_602 (O_602,N_4817,N_4864);
nor UO_603 (O_603,N_4990,N_4840);
xnor UO_604 (O_604,N_4922,N_4912);
nand UO_605 (O_605,N_4857,N_4929);
or UO_606 (O_606,N_4883,N_4900);
xnor UO_607 (O_607,N_4960,N_4829);
and UO_608 (O_608,N_4952,N_4935);
xor UO_609 (O_609,N_4839,N_4804);
or UO_610 (O_610,N_4967,N_4830);
and UO_611 (O_611,N_4977,N_4942);
nor UO_612 (O_612,N_4928,N_4810);
xnor UO_613 (O_613,N_4865,N_4920);
nand UO_614 (O_614,N_4834,N_4860);
or UO_615 (O_615,N_4891,N_4923);
nand UO_616 (O_616,N_4912,N_4866);
xnor UO_617 (O_617,N_4803,N_4922);
xor UO_618 (O_618,N_4801,N_4938);
nor UO_619 (O_619,N_4863,N_4821);
nand UO_620 (O_620,N_4888,N_4812);
and UO_621 (O_621,N_4911,N_4977);
xor UO_622 (O_622,N_4814,N_4849);
or UO_623 (O_623,N_4886,N_4810);
nor UO_624 (O_624,N_4973,N_4802);
nand UO_625 (O_625,N_4888,N_4957);
and UO_626 (O_626,N_4858,N_4959);
or UO_627 (O_627,N_4848,N_4895);
and UO_628 (O_628,N_4872,N_4886);
and UO_629 (O_629,N_4912,N_4835);
nor UO_630 (O_630,N_4990,N_4992);
xnor UO_631 (O_631,N_4937,N_4925);
xor UO_632 (O_632,N_4858,N_4900);
and UO_633 (O_633,N_4882,N_4836);
nor UO_634 (O_634,N_4828,N_4837);
and UO_635 (O_635,N_4897,N_4837);
and UO_636 (O_636,N_4820,N_4994);
and UO_637 (O_637,N_4834,N_4873);
nor UO_638 (O_638,N_4817,N_4893);
nor UO_639 (O_639,N_4866,N_4962);
nand UO_640 (O_640,N_4995,N_4923);
and UO_641 (O_641,N_4812,N_4903);
or UO_642 (O_642,N_4845,N_4834);
nor UO_643 (O_643,N_4830,N_4807);
nor UO_644 (O_644,N_4906,N_4997);
nor UO_645 (O_645,N_4902,N_4916);
or UO_646 (O_646,N_4870,N_4979);
and UO_647 (O_647,N_4956,N_4998);
and UO_648 (O_648,N_4919,N_4858);
nor UO_649 (O_649,N_4943,N_4851);
nor UO_650 (O_650,N_4901,N_4976);
xnor UO_651 (O_651,N_4858,N_4842);
or UO_652 (O_652,N_4954,N_4921);
xnor UO_653 (O_653,N_4919,N_4958);
nor UO_654 (O_654,N_4848,N_4975);
and UO_655 (O_655,N_4864,N_4894);
and UO_656 (O_656,N_4978,N_4890);
nand UO_657 (O_657,N_4820,N_4827);
or UO_658 (O_658,N_4862,N_4873);
or UO_659 (O_659,N_4812,N_4939);
nor UO_660 (O_660,N_4840,N_4839);
or UO_661 (O_661,N_4957,N_4929);
nand UO_662 (O_662,N_4855,N_4896);
nand UO_663 (O_663,N_4915,N_4941);
nand UO_664 (O_664,N_4997,N_4851);
or UO_665 (O_665,N_4849,N_4943);
and UO_666 (O_666,N_4997,N_4926);
and UO_667 (O_667,N_4974,N_4903);
and UO_668 (O_668,N_4970,N_4925);
nand UO_669 (O_669,N_4962,N_4891);
nand UO_670 (O_670,N_4836,N_4911);
or UO_671 (O_671,N_4814,N_4800);
nand UO_672 (O_672,N_4963,N_4935);
nor UO_673 (O_673,N_4891,N_4869);
and UO_674 (O_674,N_4933,N_4839);
nor UO_675 (O_675,N_4884,N_4954);
nand UO_676 (O_676,N_4947,N_4995);
nor UO_677 (O_677,N_4888,N_4908);
and UO_678 (O_678,N_4910,N_4924);
nor UO_679 (O_679,N_4932,N_4965);
nor UO_680 (O_680,N_4864,N_4804);
nor UO_681 (O_681,N_4978,N_4923);
or UO_682 (O_682,N_4915,N_4837);
or UO_683 (O_683,N_4834,N_4899);
or UO_684 (O_684,N_4937,N_4921);
and UO_685 (O_685,N_4818,N_4930);
xnor UO_686 (O_686,N_4938,N_4894);
xor UO_687 (O_687,N_4884,N_4836);
and UO_688 (O_688,N_4964,N_4984);
xnor UO_689 (O_689,N_4879,N_4869);
nor UO_690 (O_690,N_4848,N_4821);
or UO_691 (O_691,N_4961,N_4806);
or UO_692 (O_692,N_4878,N_4949);
and UO_693 (O_693,N_4842,N_4951);
nor UO_694 (O_694,N_4975,N_4817);
and UO_695 (O_695,N_4974,N_4897);
nand UO_696 (O_696,N_4811,N_4984);
or UO_697 (O_697,N_4880,N_4843);
nor UO_698 (O_698,N_4996,N_4817);
nor UO_699 (O_699,N_4953,N_4972);
nand UO_700 (O_700,N_4935,N_4981);
nand UO_701 (O_701,N_4954,N_4963);
and UO_702 (O_702,N_4951,N_4977);
or UO_703 (O_703,N_4873,N_4802);
and UO_704 (O_704,N_4912,N_4822);
nand UO_705 (O_705,N_4961,N_4959);
nand UO_706 (O_706,N_4904,N_4866);
or UO_707 (O_707,N_4948,N_4953);
nand UO_708 (O_708,N_4806,N_4994);
and UO_709 (O_709,N_4876,N_4956);
and UO_710 (O_710,N_4971,N_4895);
and UO_711 (O_711,N_4922,N_4821);
nor UO_712 (O_712,N_4935,N_4964);
nand UO_713 (O_713,N_4855,N_4822);
and UO_714 (O_714,N_4995,N_4942);
or UO_715 (O_715,N_4826,N_4896);
and UO_716 (O_716,N_4834,N_4855);
nand UO_717 (O_717,N_4800,N_4937);
or UO_718 (O_718,N_4829,N_4837);
or UO_719 (O_719,N_4973,N_4801);
or UO_720 (O_720,N_4995,N_4864);
nor UO_721 (O_721,N_4995,N_4911);
and UO_722 (O_722,N_4994,N_4938);
nor UO_723 (O_723,N_4811,N_4929);
or UO_724 (O_724,N_4895,N_4862);
and UO_725 (O_725,N_4849,N_4841);
nand UO_726 (O_726,N_4999,N_4867);
and UO_727 (O_727,N_4842,N_4863);
and UO_728 (O_728,N_4907,N_4803);
and UO_729 (O_729,N_4997,N_4987);
or UO_730 (O_730,N_4960,N_4951);
nand UO_731 (O_731,N_4928,N_4964);
and UO_732 (O_732,N_4999,N_4952);
nand UO_733 (O_733,N_4948,N_4886);
or UO_734 (O_734,N_4914,N_4925);
and UO_735 (O_735,N_4910,N_4877);
nor UO_736 (O_736,N_4840,N_4814);
xor UO_737 (O_737,N_4841,N_4944);
or UO_738 (O_738,N_4847,N_4967);
nor UO_739 (O_739,N_4809,N_4826);
and UO_740 (O_740,N_4822,N_4835);
and UO_741 (O_741,N_4813,N_4879);
nand UO_742 (O_742,N_4996,N_4885);
nor UO_743 (O_743,N_4848,N_4962);
and UO_744 (O_744,N_4837,N_4970);
xnor UO_745 (O_745,N_4815,N_4920);
nor UO_746 (O_746,N_4957,N_4872);
nand UO_747 (O_747,N_4998,N_4819);
nand UO_748 (O_748,N_4957,N_4991);
nand UO_749 (O_749,N_4820,N_4863);
nand UO_750 (O_750,N_4835,N_4826);
nor UO_751 (O_751,N_4888,N_4988);
nor UO_752 (O_752,N_4925,N_4997);
and UO_753 (O_753,N_4803,N_4959);
xor UO_754 (O_754,N_4875,N_4926);
and UO_755 (O_755,N_4930,N_4932);
xnor UO_756 (O_756,N_4812,N_4999);
and UO_757 (O_757,N_4884,N_4851);
xor UO_758 (O_758,N_4916,N_4920);
or UO_759 (O_759,N_4970,N_4890);
or UO_760 (O_760,N_4837,N_4999);
and UO_761 (O_761,N_4997,N_4934);
xor UO_762 (O_762,N_4857,N_4894);
and UO_763 (O_763,N_4805,N_4982);
nor UO_764 (O_764,N_4836,N_4925);
and UO_765 (O_765,N_4894,N_4986);
or UO_766 (O_766,N_4957,N_4801);
and UO_767 (O_767,N_4860,N_4827);
and UO_768 (O_768,N_4952,N_4919);
nand UO_769 (O_769,N_4902,N_4992);
nor UO_770 (O_770,N_4924,N_4974);
nand UO_771 (O_771,N_4984,N_4897);
nor UO_772 (O_772,N_4985,N_4920);
and UO_773 (O_773,N_4811,N_4912);
nand UO_774 (O_774,N_4837,N_4802);
nor UO_775 (O_775,N_4990,N_4833);
nand UO_776 (O_776,N_4916,N_4948);
xnor UO_777 (O_777,N_4853,N_4988);
and UO_778 (O_778,N_4812,N_4878);
and UO_779 (O_779,N_4828,N_4836);
and UO_780 (O_780,N_4973,N_4965);
and UO_781 (O_781,N_4930,N_4965);
xor UO_782 (O_782,N_4800,N_4970);
or UO_783 (O_783,N_4989,N_4855);
or UO_784 (O_784,N_4874,N_4888);
nand UO_785 (O_785,N_4818,N_4814);
nand UO_786 (O_786,N_4959,N_4984);
and UO_787 (O_787,N_4980,N_4960);
nand UO_788 (O_788,N_4929,N_4963);
and UO_789 (O_789,N_4993,N_4971);
and UO_790 (O_790,N_4962,N_4983);
nor UO_791 (O_791,N_4805,N_4962);
or UO_792 (O_792,N_4977,N_4988);
xor UO_793 (O_793,N_4918,N_4827);
nor UO_794 (O_794,N_4981,N_4967);
xor UO_795 (O_795,N_4899,N_4888);
nor UO_796 (O_796,N_4928,N_4986);
and UO_797 (O_797,N_4818,N_4903);
nor UO_798 (O_798,N_4885,N_4805);
or UO_799 (O_799,N_4826,N_4897);
nor UO_800 (O_800,N_4843,N_4805);
or UO_801 (O_801,N_4949,N_4807);
nor UO_802 (O_802,N_4954,N_4973);
nor UO_803 (O_803,N_4910,N_4856);
nor UO_804 (O_804,N_4862,N_4979);
nand UO_805 (O_805,N_4891,N_4934);
xor UO_806 (O_806,N_4836,N_4961);
and UO_807 (O_807,N_4883,N_4809);
and UO_808 (O_808,N_4965,N_4979);
nor UO_809 (O_809,N_4913,N_4804);
nand UO_810 (O_810,N_4958,N_4893);
and UO_811 (O_811,N_4986,N_4917);
or UO_812 (O_812,N_4878,N_4804);
nand UO_813 (O_813,N_4996,N_4881);
and UO_814 (O_814,N_4983,N_4878);
nand UO_815 (O_815,N_4843,N_4852);
nor UO_816 (O_816,N_4932,N_4911);
and UO_817 (O_817,N_4915,N_4901);
nand UO_818 (O_818,N_4942,N_4856);
nand UO_819 (O_819,N_4849,N_4949);
nand UO_820 (O_820,N_4928,N_4877);
nor UO_821 (O_821,N_4990,N_4943);
or UO_822 (O_822,N_4809,N_4945);
nor UO_823 (O_823,N_4939,N_4863);
or UO_824 (O_824,N_4920,N_4981);
or UO_825 (O_825,N_4842,N_4801);
xnor UO_826 (O_826,N_4937,N_4959);
nand UO_827 (O_827,N_4862,N_4943);
or UO_828 (O_828,N_4830,N_4879);
nor UO_829 (O_829,N_4816,N_4913);
nor UO_830 (O_830,N_4804,N_4870);
nand UO_831 (O_831,N_4838,N_4960);
or UO_832 (O_832,N_4915,N_4967);
and UO_833 (O_833,N_4998,N_4975);
or UO_834 (O_834,N_4987,N_4895);
or UO_835 (O_835,N_4808,N_4852);
nor UO_836 (O_836,N_4915,N_4866);
and UO_837 (O_837,N_4972,N_4897);
or UO_838 (O_838,N_4841,N_4916);
nor UO_839 (O_839,N_4880,N_4891);
nor UO_840 (O_840,N_4877,N_4817);
and UO_841 (O_841,N_4839,N_4960);
nor UO_842 (O_842,N_4840,N_4879);
xnor UO_843 (O_843,N_4849,N_4938);
and UO_844 (O_844,N_4976,N_4939);
xor UO_845 (O_845,N_4803,N_4983);
or UO_846 (O_846,N_4835,N_4966);
and UO_847 (O_847,N_4918,N_4888);
nor UO_848 (O_848,N_4821,N_4840);
nand UO_849 (O_849,N_4961,N_4928);
nand UO_850 (O_850,N_4957,N_4971);
and UO_851 (O_851,N_4984,N_4906);
or UO_852 (O_852,N_4964,N_4897);
or UO_853 (O_853,N_4837,N_4912);
or UO_854 (O_854,N_4875,N_4994);
nand UO_855 (O_855,N_4975,N_4884);
and UO_856 (O_856,N_4990,N_4914);
or UO_857 (O_857,N_4974,N_4830);
or UO_858 (O_858,N_4997,N_4971);
or UO_859 (O_859,N_4926,N_4868);
xor UO_860 (O_860,N_4905,N_4875);
and UO_861 (O_861,N_4891,N_4815);
and UO_862 (O_862,N_4865,N_4880);
or UO_863 (O_863,N_4909,N_4933);
and UO_864 (O_864,N_4852,N_4862);
nand UO_865 (O_865,N_4926,N_4989);
and UO_866 (O_866,N_4957,N_4988);
and UO_867 (O_867,N_4865,N_4875);
nor UO_868 (O_868,N_4863,N_4812);
and UO_869 (O_869,N_4821,N_4943);
nand UO_870 (O_870,N_4971,N_4921);
nor UO_871 (O_871,N_4928,N_4873);
or UO_872 (O_872,N_4872,N_4989);
nand UO_873 (O_873,N_4955,N_4917);
nand UO_874 (O_874,N_4920,N_4880);
nor UO_875 (O_875,N_4987,N_4815);
and UO_876 (O_876,N_4825,N_4986);
or UO_877 (O_877,N_4858,N_4860);
and UO_878 (O_878,N_4932,N_4984);
nand UO_879 (O_879,N_4952,N_4853);
and UO_880 (O_880,N_4839,N_4871);
xnor UO_881 (O_881,N_4843,N_4894);
xnor UO_882 (O_882,N_4811,N_4817);
nor UO_883 (O_883,N_4823,N_4850);
nor UO_884 (O_884,N_4928,N_4968);
xnor UO_885 (O_885,N_4868,N_4832);
and UO_886 (O_886,N_4945,N_4971);
and UO_887 (O_887,N_4813,N_4889);
nand UO_888 (O_888,N_4934,N_4881);
nor UO_889 (O_889,N_4823,N_4998);
nand UO_890 (O_890,N_4938,N_4860);
nor UO_891 (O_891,N_4998,N_4849);
nor UO_892 (O_892,N_4929,N_4913);
nand UO_893 (O_893,N_4847,N_4861);
xnor UO_894 (O_894,N_4935,N_4846);
nor UO_895 (O_895,N_4985,N_4892);
nor UO_896 (O_896,N_4950,N_4935);
nor UO_897 (O_897,N_4989,N_4945);
xnor UO_898 (O_898,N_4932,N_4991);
and UO_899 (O_899,N_4894,N_4963);
or UO_900 (O_900,N_4928,N_4974);
or UO_901 (O_901,N_4821,N_4950);
xor UO_902 (O_902,N_4874,N_4950);
or UO_903 (O_903,N_4887,N_4972);
or UO_904 (O_904,N_4999,N_4949);
nand UO_905 (O_905,N_4873,N_4913);
and UO_906 (O_906,N_4828,N_4919);
nand UO_907 (O_907,N_4996,N_4900);
or UO_908 (O_908,N_4905,N_4809);
and UO_909 (O_909,N_4877,N_4835);
or UO_910 (O_910,N_4805,N_4945);
nand UO_911 (O_911,N_4854,N_4923);
nand UO_912 (O_912,N_4841,N_4814);
nand UO_913 (O_913,N_4931,N_4921);
and UO_914 (O_914,N_4877,N_4871);
or UO_915 (O_915,N_4811,N_4819);
nand UO_916 (O_916,N_4868,N_4866);
nand UO_917 (O_917,N_4944,N_4961);
and UO_918 (O_918,N_4988,N_4922);
or UO_919 (O_919,N_4934,N_4941);
nor UO_920 (O_920,N_4956,N_4945);
nand UO_921 (O_921,N_4811,N_4971);
or UO_922 (O_922,N_4989,N_4846);
nand UO_923 (O_923,N_4991,N_4894);
or UO_924 (O_924,N_4991,N_4925);
xnor UO_925 (O_925,N_4917,N_4840);
and UO_926 (O_926,N_4807,N_4950);
and UO_927 (O_927,N_4844,N_4839);
or UO_928 (O_928,N_4874,N_4854);
nor UO_929 (O_929,N_4877,N_4867);
and UO_930 (O_930,N_4885,N_4984);
or UO_931 (O_931,N_4822,N_4982);
nand UO_932 (O_932,N_4900,N_4872);
nand UO_933 (O_933,N_4879,N_4817);
and UO_934 (O_934,N_4890,N_4864);
nand UO_935 (O_935,N_4843,N_4876);
nand UO_936 (O_936,N_4997,N_4866);
nand UO_937 (O_937,N_4830,N_4962);
or UO_938 (O_938,N_4944,N_4808);
nand UO_939 (O_939,N_4838,N_4938);
nor UO_940 (O_940,N_4904,N_4826);
and UO_941 (O_941,N_4829,N_4813);
or UO_942 (O_942,N_4873,N_4832);
nor UO_943 (O_943,N_4885,N_4800);
xor UO_944 (O_944,N_4892,N_4857);
or UO_945 (O_945,N_4949,N_4975);
or UO_946 (O_946,N_4868,N_4855);
nand UO_947 (O_947,N_4951,N_4894);
xnor UO_948 (O_948,N_4818,N_4881);
nand UO_949 (O_949,N_4896,N_4983);
nor UO_950 (O_950,N_4931,N_4914);
xnor UO_951 (O_951,N_4880,N_4955);
or UO_952 (O_952,N_4971,N_4806);
or UO_953 (O_953,N_4972,N_4917);
nand UO_954 (O_954,N_4911,N_4804);
nand UO_955 (O_955,N_4849,N_4914);
xnor UO_956 (O_956,N_4877,N_4934);
or UO_957 (O_957,N_4965,N_4944);
xnor UO_958 (O_958,N_4927,N_4979);
nor UO_959 (O_959,N_4855,N_4890);
nor UO_960 (O_960,N_4917,N_4957);
nor UO_961 (O_961,N_4931,N_4801);
or UO_962 (O_962,N_4929,N_4915);
xor UO_963 (O_963,N_4929,N_4819);
nand UO_964 (O_964,N_4834,N_4933);
nand UO_965 (O_965,N_4816,N_4991);
nand UO_966 (O_966,N_4990,N_4820);
nand UO_967 (O_967,N_4958,N_4862);
nor UO_968 (O_968,N_4930,N_4943);
xnor UO_969 (O_969,N_4861,N_4967);
and UO_970 (O_970,N_4879,N_4932);
xor UO_971 (O_971,N_4804,N_4985);
and UO_972 (O_972,N_4999,N_4852);
and UO_973 (O_973,N_4972,N_4961);
and UO_974 (O_974,N_4859,N_4822);
xor UO_975 (O_975,N_4943,N_4994);
or UO_976 (O_976,N_4925,N_4862);
and UO_977 (O_977,N_4959,N_4833);
nand UO_978 (O_978,N_4843,N_4983);
nand UO_979 (O_979,N_4953,N_4861);
nand UO_980 (O_980,N_4972,N_4847);
nor UO_981 (O_981,N_4960,N_4990);
nor UO_982 (O_982,N_4800,N_4815);
xnor UO_983 (O_983,N_4924,N_4870);
or UO_984 (O_984,N_4945,N_4883);
or UO_985 (O_985,N_4890,N_4910);
nand UO_986 (O_986,N_4858,N_4901);
and UO_987 (O_987,N_4922,N_4866);
nor UO_988 (O_988,N_4863,N_4816);
nor UO_989 (O_989,N_4999,N_4917);
and UO_990 (O_990,N_4829,N_4873);
and UO_991 (O_991,N_4911,N_4982);
and UO_992 (O_992,N_4970,N_4853);
nor UO_993 (O_993,N_4862,N_4990);
and UO_994 (O_994,N_4810,N_4958);
and UO_995 (O_995,N_4984,N_4979);
nor UO_996 (O_996,N_4834,N_4857);
or UO_997 (O_997,N_4855,N_4935);
xor UO_998 (O_998,N_4846,N_4822);
nand UO_999 (O_999,N_4894,N_4902);
endmodule