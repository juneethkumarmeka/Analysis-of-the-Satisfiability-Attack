module basic_2500_25000_3000_25_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
and U0 (N_0,In_1655,In_379);
nor U1 (N_1,In_2279,In_1864);
xor U2 (N_2,In_885,In_2413);
nand U3 (N_3,In_453,In_59);
and U4 (N_4,In_1666,In_2034);
or U5 (N_5,In_438,In_892);
and U6 (N_6,In_578,In_2294);
xor U7 (N_7,In_1620,In_406);
and U8 (N_8,In_898,In_1999);
nand U9 (N_9,In_1785,In_447);
and U10 (N_10,In_1578,In_2020);
nor U11 (N_11,In_1483,In_394);
xnor U12 (N_12,In_416,In_2376);
or U13 (N_13,In_2378,In_2400);
nor U14 (N_14,In_1489,In_1735);
and U15 (N_15,In_1567,In_2347);
and U16 (N_16,In_1037,In_2026);
xor U17 (N_17,In_959,In_1584);
nand U18 (N_18,In_642,In_2403);
xor U19 (N_19,In_425,In_997);
and U20 (N_20,In_486,In_1968);
or U21 (N_21,In_585,In_1798);
xnor U22 (N_22,In_1030,In_1733);
nand U23 (N_23,In_1721,In_2252);
xor U24 (N_24,In_1557,In_781);
and U25 (N_25,In_2205,In_2384);
xnor U26 (N_26,In_915,In_2375);
xor U27 (N_27,In_1628,In_1061);
nor U28 (N_28,In_1381,In_2335);
and U29 (N_29,In_2425,In_81);
and U30 (N_30,In_599,In_799);
and U31 (N_31,In_670,In_2043);
or U32 (N_32,In_1141,In_5);
or U33 (N_33,In_161,In_1817);
and U34 (N_34,In_79,In_1335);
or U35 (N_35,In_675,In_780);
and U36 (N_36,In_75,In_2364);
and U37 (N_37,In_2007,In_415);
nand U38 (N_38,In_1123,In_1824);
and U39 (N_39,In_8,In_397);
nand U40 (N_40,In_2325,In_2151);
or U41 (N_41,In_1513,In_407);
or U42 (N_42,In_1209,In_2154);
or U43 (N_43,In_1057,In_1895);
or U44 (N_44,In_882,In_604);
or U45 (N_45,In_1617,In_559);
nor U46 (N_46,In_1741,In_1219);
nor U47 (N_47,In_1164,In_1361);
xnor U48 (N_48,In_1414,In_851);
and U49 (N_49,In_1725,In_1067);
nand U50 (N_50,In_727,In_2157);
or U51 (N_51,In_175,In_134);
nand U52 (N_52,In_146,In_1076);
nor U53 (N_53,In_345,In_1486);
and U54 (N_54,In_2027,In_2048);
and U55 (N_55,In_2153,In_1705);
nand U56 (N_56,In_850,In_2447);
xnor U57 (N_57,In_149,In_1822);
nor U58 (N_58,In_34,In_1972);
xor U59 (N_59,In_1244,In_444);
nand U60 (N_60,In_2396,In_1853);
nor U61 (N_61,In_1920,In_2427);
nor U62 (N_62,In_2052,In_900);
nor U63 (N_63,In_852,In_2306);
or U64 (N_64,In_1607,In_1115);
xor U65 (N_65,In_1826,In_1878);
xor U66 (N_66,In_100,In_1376);
nor U67 (N_67,In_244,In_895);
or U68 (N_68,In_813,In_1954);
nor U69 (N_69,In_726,In_331);
nor U70 (N_70,In_634,In_1544);
nor U71 (N_71,In_23,In_1901);
or U72 (N_72,In_1193,In_2088);
xnor U73 (N_73,In_280,In_1812);
or U74 (N_74,In_1506,In_2074);
or U75 (N_75,In_963,In_2085);
nor U76 (N_76,In_1269,In_1861);
or U77 (N_77,In_63,In_231);
nand U78 (N_78,In_327,In_381);
xnor U79 (N_79,In_360,In_1010);
nor U80 (N_80,In_547,In_2383);
xnor U81 (N_81,In_1162,In_1024);
or U82 (N_82,In_1137,In_1093);
xor U83 (N_83,In_2078,In_1604);
nor U84 (N_84,In_925,In_690);
xnor U85 (N_85,In_1433,In_861);
xnor U86 (N_86,In_1836,In_2408);
xor U87 (N_87,In_340,In_2351);
xnor U88 (N_88,In_1548,In_879);
or U89 (N_89,In_545,In_1151);
and U90 (N_90,In_2231,In_2199);
nand U91 (N_91,In_769,In_907);
or U92 (N_92,In_1158,In_533);
nor U93 (N_93,In_2177,In_249);
xor U94 (N_94,In_405,In_2077);
xnor U95 (N_95,In_56,In_1425);
and U96 (N_96,In_735,In_1202);
or U97 (N_97,In_2286,In_857);
or U98 (N_98,In_1908,In_1247);
nor U99 (N_99,In_1272,In_1637);
nand U100 (N_100,In_370,In_913);
xnor U101 (N_101,In_948,In_1281);
and U102 (N_102,In_1038,In_686);
and U103 (N_103,In_409,In_871);
and U104 (N_104,In_1983,In_470);
and U105 (N_105,In_1399,In_2421);
or U106 (N_106,In_1198,In_229);
and U107 (N_107,In_1287,In_1809);
nor U108 (N_108,In_2476,In_2198);
and U109 (N_109,In_93,In_1386);
or U110 (N_110,In_2387,In_273);
xor U111 (N_111,In_2135,In_884);
nor U112 (N_112,In_1933,In_2379);
nor U113 (N_113,In_1136,In_2099);
xnor U114 (N_114,In_2029,In_2289);
nor U115 (N_115,In_1438,In_1424);
nand U116 (N_116,In_1035,In_776);
xor U117 (N_117,In_1396,In_1215);
nand U118 (N_118,In_877,In_2140);
nor U119 (N_119,In_153,In_2050);
or U120 (N_120,In_2105,In_1967);
xor U121 (N_121,In_2233,In_1251);
nor U122 (N_122,In_1624,In_1978);
and U123 (N_123,In_128,In_133);
xor U124 (N_124,In_1467,In_2467);
xor U125 (N_125,In_514,In_1079);
nand U126 (N_126,In_2158,In_868);
xor U127 (N_127,In_1588,In_999);
xnor U128 (N_128,In_552,In_1563);
xnor U129 (N_129,In_32,In_2036);
and U130 (N_130,In_183,In_2039);
nor U131 (N_131,In_1441,In_433);
xnor U132 (N_132,In_1755,In_402);
xnor U133 (N_133,In_557,In_692);
nand U134 (N_134,In_29,In_1599);
or U135 (N_135,In_355,In_1993);
nand U136 (N_136,In_341,In_1953);
and U137 (N_137,In_304,In_1996);
or U138 (N_138,In_2075,In_1278);
or U139 (N_139,In_795,In_1071);
or U140 (N_140,In_178,In_1600);
or U141 (N_141,In_677,In_2493);
xor U142 (N_142,In_869,In_1085);
nand U143 (N_143,In_946,In_1355);
nand U144 (N_144,In_1815,In_1431);
nand U145 (N_145,In_2272,In_1343);
nor U146 (N_146,In_2355,In_2037);
or U147 (N_147,In_635,In_323);
nand U148 (N_148,In_947,In_181);
nand U149 (N_149,In_1105,In_1777);
xnor U150 (N_150,In_967,In_504);
or U151 (N_151,In_908,In_1491);
and U152 (N_152,In_285,In_234);
or U153 (N_153,In_1195,In_1305);
or U154 (N_154,In_1976,In_176);
xor U155 (N_155,In_1,In_1510);
or U156 (N_156,In_1475,In_1520);
or U157 (N_157,In_794,In_1747);
or U158 (N_158,In_358,In_1442);
and U159 (N_159,In_35,In_203);
nand U160 (N_160,In_1565,In_1044);
nor U161 (N_161,In_2219,In_191);
xor U162 (N_162,In_1471,In_1228);
xor U163 (N_163,In_1683,In_928);
nand U164 (N_164,In_1702,In_2412);
or U165 (N_165,In_673,In_770);
nor U166 (N_166,In_732,In_1060);
or U167 (N_167,In_89,In_1172);
xor U168 (N_168,In_2016,In_154);
xnor U169 (N_169,In_1233,In_1249);
nand U170 (N_170,In_1133,In_827);
nor U171 (N_171,In_91,In_1612);
or U172 (N_172,In_1776,In_344);
nor U173 (N_173,In_1855,In_1333);
and U174 (N_174,In_2280,In_80);
xnor U175 (N_175,In_1937,In_1019);
and U176 (N_176,In_2435,In_1152);
or U177 (N_177,In_1689,In_1793);
or U178 (N_178,In_322,In_1421);
or U179 (N_179,In_839,In_1288);
or U180 (N_180,In_168,In_2430);
or U181 (N_181,In_1778,In_2481);
xor U182 (N_182,In_2262,In_279);
or U183 (N_183,In_1835,In_1979);
xnor U184 (N_184,In_1009,In_1602);
xor U185 (N_185,In_553,In_1282);
nand U186 (N_186,In_970,In_1201);
nand U187 (N_187,In_1810,In_1299);
or U188 (N_188,In_159,In_2066);
nor U189 (N_189,In_1879,In_1256);
nor U190 (N_190,In_1779,In_2118);
nor U191 (N_191,In_1332,In_1615);
nor U192 (N_192,In_198,In_2110);
nor U193 (N_193,In_1929,In_1938);
nand U194 (N_194,In_1488,In_992);
and U195 (N_195,In_1668,In_1827);
or U196 (N_196,In_617,In_945);
nand U197 (N_197,In_202,In_69);
nor U198 (N_198,In_806,In_1517);
nor U199 (N_199,In_2002,In_1562);
and U200 (N_200,In_2031,In_531);
nor U201 (N_201,In_169,In_694);
and U202 (N_202,In_2220,In_2082);
and U203 (N_203,In_87,In_2269);
xor U204 (N_204,In_1610,In_582);
xor U205 (N_205,In_1769,In_237);
nand U206 (N_206,In_520,In_660);
and U207 (N_207,In_853,In_1234);
and U208 (N_208,In_140,In_1239);
and U209 (N_209,In_47,In_1591);
nor U210 (N_210,In_497,In_658);
nor U211 (N_211,In_2474,In_1230);
or U212 (N_212,In_541,In_640);
or U213 (N_213,In_1816,In_307);
or U214 (N_214,In_894,In_1130);
and U215 (N_215,In_576,In_12);
or U216 (N_216,In_1395,In_1865);
nor U217 (N_217,In_812,In_1064);
nor U218 (N_218,In_1698,In_1350);
and U219 (N_219,In_1914,In_25);
or U220 (N_220,In_1950,In_150);
or U221 (N_221,In_1905,In_82);
xnor U222 (N_222,In_1401,In_68);
and U223 (N_223,In_395,In_1648);
nor U224 (N_224,In_2276,In_21);
nand U225 (N_225,In_1728,In_343);
or U226 (N_226,In_2495,In_1519);
nor U227 (N_227,In_1190,In_1238);
and U228 (N_228,In_1558,In_1393);
xnor U229 (N_229,In_1896,In_305);
or U230 (N_230,In_1385,In_589);
or U231 (N_231,In_2482,In_1528);
xnor U232 (N_232,In_99,In_1625);
and U233 (N_233,In_350,In_1882);
nand U234 (N_234,In_890,In_782);
xor U235 (N_235,In_1410,In_1764);
or U236 (N_236,In_1791,In_2166);
nand U237 (N_237,In_2441,In_96);
nor U238 (N_238,In_2455,In_2149);
xnor U239 (N_239,In_2155,In_454);
or U240 (N_240,In_840,In_785);
or U241 (N_241,In_53,In_392);
nand U242 (N_242,In_1984,In_162);
and U243 (N_243,In_1939,In_2247);
xor U244 (N_244,In_1631,In_72);
and U245 (N_245,In_429,In_238);
nor U246 (N_246,In_2139,In_612);
and U247 (N_247,In_2464,In_984);
nand U248 (N_248,In_1383,In_1404);
nand U249 (N_249,In_1677,In_54);
nand U250 (N_250,In_1349,In_940);
nor U251 (N_251,In_2423,In_507);
nor U252 (N_252,In_826,In_2137);
and U253 (N_253,In_2372,In_905);
or U254 (N_254,In_390,In_717);
nor U255 (N_255,In_1459,In_939);
nor U256 (N_256,In_2209,In_27);
and U257 (N_257,In_1831,In_2370);
nand U258 (N_258,In_378,In_2010);
xnor U259 (N_259,In_2101,In_631);
nor U260 (N_260,In_212,In_579);
xnor U261 (N_261,In_84,In_1837);
xnor U262 (N_262,In_1127,In_1461);
nand U263 (N_263,In_1188,In_2117);
or U264 (N_264,In_515,In_382);
nand U265 (N_265,In_1384,In_1918);
nor U266 (N_266,In_2317,In_247);
or U267 (N_267,In_2331,In_2388);
xor U268 (N_268,In_1270,In_1659);
xor U269 (N_269,In_2207,In_808);
or U270 (N_270,In_2449,In_1840);
nor U271 (N_271,In_2256,In_523);
nand U272 (N_272,In_2466,In_297);
or U273 (N_273,In_38,In_957);
and U274 (N_274,In_2361,In_1175);
xnor U275 (N_275,In_1122,In_1113);
and U276 (N_276,In_487,In_1761);
nor U277 (N_277,In_143,In_985);
nand U278 (N_278,In_2263,In_1661);
or U279 (N_279,In_1212,In_1492);
nor U280 (N_280,In_97,In_1267);
xnor U281 (N_281,In_529,In_856);
and U282 (N_282,In_929,In_982);
nand U283 (N_283,In_1416,In_650);
xnor U284 (N_284,In_1797,In_1216);
and U285 (N_285,In_1555,In_2391);
nand U286 (N_286,In_2188,In_7);
nand U287 (N_287,In_156,In_66);
and U288 (N_288,In_434,In_2187);
xor U289 (N_289,In_1751,In_1985);
nand U290 (N_290,In_702,In_1737);
xnor U291 (N_291,In_535,In_1945);
nand U292 (N_292,In_393,In_2015);
and U293 (N_293,In_2073,In_615);
nand U294 (N_294,In_145,In_471);
or U295 (N_295,In_2097,In_2203);
xor U296 (N_296,In_152,In_2454);
nand U297 (N_297,In_1266,In_2485);
xnor U298 (N_298,In_1970,In_2164);
nor U299 (N_299,In_1014,In_28);
xnor U300 (N_300,In_2092,In_330);
or U301 (N_301,In_1499,In_2359);
nand U302 (N_302,In_888,In_2406);
nor U303 (N_303,In_2003,In_995);
xor U304 (N_304,In_2065,In_1371);
or U305 (N_305,In_2393,In_2009);
nand U306 (N_306,In_462,In_1632);
and U307 (N_307,In_2259,In_1833);
nor U308 (N_308,In_1874,In_719);
or U309 (N_309,In_105,In_536);
nor U310 (N_310,In_1360,In_975);
xor U311 (N_311,In_1575,In_728);
nand U312 (N_312,In_1033,In_459);
nor U313 (N_313,In_461,In_1148);
xor U314 (N_314,In_253,In_555);
xor U315 (N_315,In_349,In_2470);
or U316 (N_316,In_2419,In_2319);
nor U317 (N_317,In_1524,In_324);
nor U318 (N_318,In_1946,In_1196);
xor U319 (N_319,In_264,In_1723);
and U320 (N_320,In_1280,In_2273);
nand U321 (N_321,In_1186,In_1790);
and U322 (N_322,In_935,In_137);
nand U323 (N_323,In_432,In_0);
nand U324 (N_324,In_730,In_2450);
xor U325 (N_325,In_2098,In_98);
xnor U326 (N_326,In_362,In_722);
nand U327 (N_327,In_1640,In_2349);
or U328 (N_328,In_1529,In_1549);
nand U329 (N_329,In_2114,In_1095);
nand U330 (N_330,In_952,In_1205);
and U331 (N_331,In_428,In_1375);
and U332 (N_332,In_596,In_22);
nor U333 (N_333,In_991,In_184);
nor U334 (N_334,In_1446,In_1144);
or U335 (N_335,In_116,In_92);
and U336 (N_336,In_309,In_94);
or U337 (N_337,In_2172,In_891);
and U338 (N_338,In_1961,In_15);
or U339 (N_339,In_2463,In_616);
or U340 (N_340,In_512,In_1553);
xnor U341 (N_341,In_2060,In_1448);
nand U342 (N_342,In_1973,In_2056);
xnor U343 (N_343,In_2044,In_1246);
nand U344 (N_344,In_807,In_527);
and U345 (N_345,In_676,In_843);
nand U346 (N_346,In_2080,In_1850);
and U347 (N_347,In_976,In_2439);
nor U348 (N_348,In_1497,In_2251);
xor U349 (N_349,In_2108,In_697);
nand U350 (N_350,In_765,In_1722);
xnor U351 (N_351,In_875,In_1088);
xor U352 (N_352,In_2165,In_798);
xnor U353 (N_353,In_1153,In_463);
nand U354 (N_354,In_1672,In_584);
xor U355 (N_355,In_1873,In_2072);
nor U356 (N_356,In_969,In_2498);
nand U357 (N_357,In_556,In_2196);
nor U358 (N_358,In_2054,In_823);
nor U359 (N_359,In_1400,In_990);
nor U360 (N_360,In_2161,In_1200);
nand U361 (N_361,In_351,In_319);
nand U362 (N_362,In_1956,In_1963);
or U363 (N_363,In_371,In_325);
and U364 (N_364,In_1770,In_902);
xor U365 (N_365,In_1685,In_1104);
xnor U366 (N_366,In_242,In_1058);
xnor U367 (N_367,In_1225,In_365);
xnor U368 (N_368,In_2310,In_740);
xor U369 (N_369,In_1045,In_2235);
xnor U370 (N_370,In_800,In_2488);
nor U371 (N_371,In_318,In_1263);
xor U372 (N_372,In_849,In_464);
or U373 (N_373,In_289,In_2300);
or U374 (N_374,In_125,In_760);
nor U375 (N_375,In_1464,In_1106);
xor U376 (N_376,In_142,In_1684);
xor U377 (N_377,In_1094,In_41);
nor U378 (N_378,In_2225,In_1796);
or U379 (N_379,In_1765,In_865);
and U380 (N_380,In_138,In_1924);
xor U381 (N_381,In_1805,In_130);
nor U382 (N_382,In_398,In_815);
and U383 (N_383,In_1444,In_801);
or U384 (N_384,In_2298,In_46);
xor U385 (N_385,In_588,In_2035);
nor U386 (N_386,In_1081,In_270);
or U387 (N_387,In_1902,In_1884);
nor U388 (N_388,In_2124,In_1883);
and U389 (N_389,In_1587,In_649);
nor U390 (N_390,In_2051,In_1695);
xnor U391 (N_391,In_1843,In_2301);
and U392 (N_392,In_348,In_1596);
nand U393 (N_393,In_2314,In_479);
xnor U394 (N_394,In_1023,In_789);
nor U395 (N_395,In_1825,In_1097);
xor U396 (N_396,In_2451,In_1880);
or U397 (N_397,In_1366,In_9);
nand U398 (N_398,In_2143,In_2171);
nand U399 (N_399,In_2181,In_1931);
or U400 (N_400,In_368,In_2363);
or U401 (N_401,In_1022,In_1654);
nor U402 (N_402,In_2047,In_1813);
and U403 (N_403,In_1821,In_1899);
xnor U404 (N_404,In_216,In_647);
nand U405 (N_405,In_2366,In_1072);
nand U406 (N_406,In_1573,In_2365);
nor U407 (N_407,In_934,In_144);
and U408 (N_408,In_1254,In_1155);
or U409 (N_409,In_2320,In_2264);
nand U410 (N_410,In_2255,In_218);
nor U411 (N_411,In_1353,In_1692);
or U412 (N_412,In_1876,In_2030);
nand U413 (N_413,In_1116,In_70);
nor U414 (N_414,In_1830,In_494);
or U415 (N_415,In_1316,In_2213);
xnor U416 (N_416,In_2302,In_2134);
nand U417 (N_417,In_421,In_448);
nor U418 (N_418,In_951,In_2169);
nor U419 (N_419,In_1616,In_938);
nand U420 (N_420,In_2215,In_276);
nand U421 (N_421,In_1250,In_955);
nor U422 (N_422,In_1566,In_1409);
xnor U423 (N_423,In_753,In_701);
nand U424 (N_424,In_185,In_312);
and U425 (N_425,In_364,In_228);
or U426 (N_426,In_1494,In_236);
and U427 (N_427,In_761,In_1454);
nand U428 (N_428,In_43,In_1619);
nand U429 (N_429,In_980,In_49);
and U430 (N_430,In_1479,In_2443);
and U431 (N_431,In_2023,In_822);
and U432 (N_432,In_958,In_1257);
nor U433 (N_433,In_936,In_1322);
xor U434 (N_434,In_2190,In_546);
xor U435 (N_435,In_2337,In_317);
nand U436 (N_436,In_1647,In_465);
xor U437 (N_437,In_2163,In_1289);
or U438 (N_438,In_20,In_1407);
xnor U439 (N_439,In_713,In_1258);
and U440 (N_440,In_190,In_912);
and U441 (N_441,In_1633,In_2446);
xnor U442 (N_442,In_1759,In_1872);
xor U443 (N_443,In_1975,In_972);
xnor U444 (N_444,In_2227,In_1646);
xor U445 (N_445,In_1580,In_1671);
xnor U446 (N_446,In_1143,In_820);
or U447 (N_447,In_2362,In_44);
xor U448 (N_448,In_1165,In_186);
xor U449 (N_449,In_2316,In_1040);
nor U450 (N_450,In_924,In_2265);
and U451 (N_451,In_2472,In_1049);
and U452 (N_452,In_1521,In_2444);
xor U453 (N_453,In_1688,In_1255);
and U454 (N_454,In_821,In_643);
nor U455 (N_455,In_2241,In_653);
and U456 (N_456,In_906,In_603);
and U457 (N_457,In_1331,In_250);
nor U458 (N_458,In_1626,In_778);
nand U459 (N_459,In_1080,In_499);
nor U460 (N_460,In_564,In_1264);
or U461 (N_461,In_2305,In_771);
xor U462 (N_462,In_2307,In_403);
and U463 (N_463,In_1460,In_286);
and U464 (N_464,In_151,In_227);
or U465 (N_465,In_2250,In_2407);
nand U466 (N_466,In_1069,In_506);
nand U467 (N_467,In_1051,In_1378);
xnor U468 (N_468,In_864,In_988);
and U469 (N_469,In_2128,In_708);
nand U470 (N_470,In_1848,In_422);
nand U471 (N_471,In_2428,In_33);
and U472 (N_472,In_1382,In_430);
and U473 (N_473,In_58,In_1154);
xor U474 (N_474,In_291,In_1284);
and U475 (N_475,In_254,In_1053);
or U476 (N_476,In_1134,In_583);
or U477 (N_477,In_575,In_2017);
nor U478 (N_478,In_1356,In_2288);
nor U479 (N_479,In_1534,In_1504);
or U480 (N_480,In_1303,In_836);
and U481 (N_481,In_2338,In_1713);
or U482 (N_482,In_797,In_2336);
xnor U483 (N_483,In_439,In_1774);
or U484 (N_484,In_662,In_942);
or U485 (N_485,In_918,In_1398);
and U486 (N_486,In_1856,In_554);
nor U487 (N_487,In_1187,In_965);
xor U488 (N_488,In_1098,In_881);
xnor U489 (N_489,In_482,In_1527);
nand U490 (N_490,In_310,In_1394);
nand U491 (N_491,In_2392,In_373);
nand U492 (N_492,In_1174,In_729);
xor U493 (N_493,In_1403,In_347);
nor U494 (N_494,In_505,In_1969);
nor U495 (N_495,In_1101,In_981);
and U496 (N_496,In_1320,In_1161);
xnor U497 (N_497,In_18,In_786);
and U498 (N_498,In_2212,In_1913);
and U499 (N_499,In_290,In_1301);
and U500 (N_500,In_1427,In_628);
and U501 (N_501,In_2332,In_1503);
or U502 (N_502,In_777,In_804);
nor U503 (N_503,In_921,In_2303);
or U504 (N_504,In_141,In_2497);
xnor U505 (N_505,In_2390,In_1227);
nor U506 (N_506,In_171,In_2448);
and U507 (N_507,In_654,In_1339);
xor U508 (N_508,In_1919,In_1845);
xor U509 (N_509,In_1203,In_61);
or U510 (N_510,In_314,In_1804);
nor U511 (N_511,In_391,In_2244);
nand U512 (N_512,In_1430,In_1342);
or U513 (N_513,In_255,In_1468);
nand U514 (N_514,In_1224,In_2465);
xnor U515 (N_515,In_954,In_516);
xnor U516 (N_516,In_2386,In_1315);
nor U517 (N_517,In_95,In_2429);
and U518 (N_518,In_2424,In_1474);
nand U519 (N_519,In_550,In_1715);
or U520 (N_520,In_695,In_1603);
xor U521 (N_521,In_2133,In_2275);
xor U522 (N_522,In_664,In_2452);
or U523 (N_523,In_1470,In_1013);
or U524 (N_524,In_2477,In_1055);
nor U525 (N_525,In_2113,In_1906);
nor U526 (N_526,In_613,In_1163);
nor U527 (N_527,In_863,In_1740);
and U528 (N_528,In_1423,In_1412);
xor U529 (N_529,In_411,In_2120);
xor U530 (N_530,In_1261,In_1718);
xor U531 (N_531,In_1197,In_1710);
xor U532 (N_532,In_1149,In_2290);
and U533 (N_533,In_2218,In_2432);
nor U534 (N_534,In_139,In_2475);
nor U535 (N_535,In_1002,In_1235);
xnor U536 (N_536,In_372,In_566);
nor U537 (N_537,In_1171,In_2479);
or U538 (N_538,In_723,In_271);
nor U539 (N_539,In_870,In_1473);
or U540 (N_540,In_1598,In_1121);
and U541 (N_541,In_277,In_1570);
and U542 (N_542,In_2278,In_1231);
nor U543 (N_543,In_774,In_623);
and U544 (N_544,In_1877,In_114);
xnor U545 (N_545,In_1744,In_2182);
or U546 (N_546,In_1047,In_1732);
nor U547 (N_547,In_591,In_1992);
xnor U548 (N_548,In_189,In_903);
or U549 (N_549,In_2226,In_1749);
nand U550 (N_550,In_225,In_73);
xnor U551 (N_551,In_1437,In_1168);
nor U552 (N_552,In_1241,In_1841);
nand U553 (N_553,In_1008,In_363);
or U554 (N_554,In_845,In_1704);
nor U555 (N_555,In_136,In_1177);
nor U556 (N_556,In_1936,In_1140);
or U557 (N_557,In_1980,In_2156);
and U558 (N_558,In_2234,In_2096);
or U559 (N_559,In_1321,In_1478);
nor U560 (N_560,In_1117,In_1319);
nand U561 (N_561,In_1112,In_2127);
and U562 (N_562,In_467,In_1859);
nand U563 (N_563,In_2090,In_1621);
and U564 (N_564,In_109,In_1229);
nor U565 (N_565,In_488,In_1443);
or U566 (N_566,In_489,In_353);
xnor U567 (N_567,In_744,In_300);
xnor U568 (N_568,In_672,In_2442);
nand U569 (N_569,In_1917,In_1422);
or U570 (N_570,In_899,In_636);
xnor U571 (N_571,In_1476,In_2324);
nor U572 (N_572,In_2360,In_1054);
and U573 (N_573,In_1909,In_517);
or U574 (N_574,In_847,In_222);
and U575 (N_575,In_568,In_910);
nor U576 (N_576,In_177,In_410);
nor U577 (N_577,In_2480,In_356);
or U578 (N_578,In_1028,In_594);
or U579 (N_579,In_2186,In_1886);
xor U580 (N_580,In_949,In_2069);
nand U581 (N_581,In_1243,In_2401);
nor U582 (N_582,In_306,In_1048);
xor U583 (N_583,In_400,In_1703);
xnor U584 (N_584,In_646,In_2191);
xor U585 (N_585,In_2116,In_2445);
nor U586 (N_586,In_1605,In_233);
and U587 (N_587,In_74,In_1370);
xnor U588 (N_588,In_2178,In_1550);
nand U589 (N_589,In_2437,In_607);
nand U590 (N_590,In_275,In_2341);
and U591 (N_591,In_2206,In_498);
nor U592 (N_592,In_721,In_1408);
xor U593 (N_593,In_45,In_876);
nor U594 (N_594,In_1042,In_1189);
nor U595 (N_595,In_1858,In_1569);
and U596 (N_596,In_1276,In_303);
or U597 (N_597,In_920,In_1124);
nand U598 (N_598,In_718,In_256);
and U599 (N_599,In_1531,In_361);
nor U600 (N_600,In_2486,In_36);
nor U601 (N_601,In_1358,In_1629);
xnor U602 (N_602,In_1636,In_745);
and U603 (N_603,In_537,In_2284);
and U604 (N_604,In_1103,In_1611);
nor U605 (N_605,In_1852,In_858);
or U606 (N_606,In_2281,In_1498);
or U607 (N_607,In_1857,In_1700);
nand U608 (N_608,In_1800,In_659);
and U609 (N_609,In_40,In_711);
and U610 (N_610,In_1167,In_226);
nand U611 (N_611,In_1893,In_232);
nand U612 (N_612,In_282,In_1445);
xor U613 (N_613,In_1328,In_1312);
nand U614 (N_614,In_867,In_267);
or U615 (N_615,In_715,In_1743);
and U616 (N_616,In_1087,In_1622);
nor U617 (N_617,In_1971,In_1653);
and U618 (N_618,In_1297,In_2115);
or U619 (N_619,In_292,In_1330);
or U620 (N_620,In_2368,In_10);
nor U621 (N_621,In_1958,In_1223);
and U622 (N_622,In_2274,In_442);
nor U623 (N_623,In_2326,In_809);
and U624 (N_624,In_1965,In_2204);
nor U625 (N_625,In_598,In_1001);
nor U626 (N_626,In_2369,In_1199);
nand U627 (N_627,In_608,In_641);
or U628 (N_628,In_252,In_126);
nand U629 (N_629,In_2285,In_1062);
xnor U630 (N_630,In_1413,In_83);
and U631 (N_631,In_2063,In_1182);
xnor U632 (N_632,In_933,In_413);
or U633 (N_633,In_1015,In_2330);
xor U634 (N_634,In_1540,In_1794);
or U635 (N_635,In_927,In_689);
nor U636 (N_636,In_874,In_1773);
nor U637 (N_637,In_42,In_751);
xor U638 (N_638,In_1389,In_1944);
nor U639 (N_639,In_2142,In_223);
and U640 (N_640,In_243,In_1179);
nor U641 (N_641,In_716,In_1518);
and U642 (N_642,In_102,In_51);
or U643 (N_643,In_669,In_1039);
xnor U644 (N_644,In_1495,In_1334);
xnor U645 (N_645,In_1670,In_2038);
nor U646 (N_646,In_1729,In_2257);
or U647 (N_647,In_490,In_805);
xor U648 (N_648,In_1966,In_614);
xnor U649 (N_649,In_2389,In_1031);
nor U650 (N_650,In_404,In_424);
and U651 (N_651,In_1135,In_1590);
and U652 (N_652,In_197,In_1814);
or U653 (N_653,In_814,In_2076);
nor U654 (N_654,In_1472,In_1726);
nor U655 (N_655,In_2478,In_1948);
nand U656 (N_656,In_2018,In_911);
or U657 (N_657,In_1745,In_1960);
or U658 (N_658,In_831,In_1736);
or U659 (N_659,In_217,In_994);
nand U660 (N_660,In_1799,In_2287);
nand U661 (N_661,In_328,In_1923);
nor U662 (N_662,In_301,In_1808);
and U663 (N_663,In_1453,In_1868);
xnor U664 (N_664,In_2471,In_1579);
xor U665 (N_665,In_1511,In_998);
and U666 (N_666,In_160,In_108);
nand U667 (N_667,In_1897,In_1614);
nor U668 (N_668,In_451,In_1415);
xnor U669 (N_669,In_748,In_790);
xnor U670 (N_670,In_2087,In_2179);
and U671 (N_671,In_944,In_1652);
nand U672 (N_672,In_2440,In_1650);
or U673 (N_673,In_1240,In_2183);
nor U674 (N_674,In_86,In_977);
and U675 (N_675,In_1887,In_742);
nor U676 (N_676,In_260,In_2377);
and U677 (N_677,In_2167,In_2489);
or U678 (N_678,In_1783,In_208);
nor U679 (N_679,In_842,In_1004);
nor U680 (N_680,In_460,In_491);
or U681 (N_681,In_2283,In_200);
and U682 (N_682,In_2112,In_1128);
and U683 (N_683,In_562,In_1428);
or U684 (N_684,In_1667,In_1477);
nand U685 (N_685,In_2395,In_2086);
nor U686 (N_686,In_2297,In_1220);
and U687 (N_687,In_2131,In_163);
or U688 (N_688,In_2339,In_2006);
nand U689 (N_689,In_1568,In_2321);
xor U690 (N_690,In_1708,In_802);
nor U691 (N_691,In_2146,In_272);
xnor U692 (N_692,In_1213,In_110);
or U693 (N_693,In_743,In_1306);
and U694 (N_694,In_2111,In_2024);
or U695 (N_695,In_830,In_6);
or U696 (N_696,In_2356,In_1951);
xnor U697 (N_697,In_158,In_1663);
nor U698 (N_698,In_1782,In_257);
nand U699 (N_699,In_1947,In_2352);
nor U700 (N_700,In_710,In_524);
and U701 (N_701,In_1927,In_2058);
and U702 (N_702,In_64,In_1131);
or U703 (N_703,In_1447,In_375);
nand U704 (N_704,In_586,In_2004);
xor U705 (N_705,In_495,In_2159);
and U706 (N_706,In_1724,In_106);
and U707 (N_707,In_1932,In_132);
or U708 (N_708,In_1206,In_2170);
nand U709 (N_709,In_793,In_860);
nand U710 (N_710,In_2342,In_768);
and U711 (N_711,In_268,In_679);
and U712 (N_712,In_901,In_757);
or U713 (N_713,In_1691,In_2084);
nor U714 (N_714,In_1997,In_883);
nor U715 (N_715,In_762,In_522);
xnor U716 (N_716,In_1977,In_2469);
nor U717 (N_717,In_387,In_1860);
xor U718 (N_718,In_766,In_1678);
nor U719 (N_719,In_179,In_973);
nand U720 (N_720,In_862,In_1012);
and U721 (N_721,In_377,In_1125);
xnor U722 (N_722,In_1086,In_538);
and U723 (N_723,In_824,In_941);
or U724 (N_724,In_2245,In_1419);
and U725 (N_725,In_1184,In_1218);
or U726 (N_726,In_2309,In_214);
or U727 (N_727,In_2490,In_787);
nand U728 (N_728,In_1662,In_848);
xnor U729 (N_729,In_962,In_1046);
xor U730 (N_730,In_561,In_704);
xnor U731 (N_731,In_1390,In_1526);
xor U732 (N_732,In_1731,In_1828);
and U733 (N_733,In_1952,In_811);
or U734 (N_734,In_1434,In_57);
xor U735 (N_735,In_1892,In_2189);
and U736 (N_736,In_386,In_1748);
nand U737 (N_737,In_299,In_2322);
or U738 (N_738,In_746,In_2311);
xnor U739 (N_739,In_1180,In_1940);
and U740 (N_740,In_2014,In_296);
xnor U741 (N_741,In_188,In_2228);
nor U742 (N_742,In_752,In_2200);
xor U743 (N_743,In_1959,In_1807);
or U744 (N_744,In_187,In_1639);
or U745 (N_745,In_103,In_2144);
xnor U746 (N_746,In_315,In_1391);
nor U747 (N_747,In_1537,In_294);
and U748 (N_748,In_1838,In_1716);
and U749 (N_749,In_2242,In_2136);
and U750 (N_750,In_1084,In_887);
xor U751 (N_751,In_1092,In_1114);
or U752 (N_752,In_889,In_2420);
nor U753 (N_753,In_1432,In_1169);
or U754 (N_754,In_1847,In_2046);
nand U755 (N_755,In_1340,In_1806);
nand U756 (N_756,In_657,In_52);
or U757 (N_757,In_1310,In_493);
nor U758 (N_758,In_1368,In_1248);
nor U759 (N_759,In_2238,In_1789);
and U760 (N_760,In_1102,In_1645);
nor U761 (N_761,In_1075,In_119);
and U762 (N_762,In_1222,In_656);
or U763 (N_763,In_592,In_1982);
nor U764 (N_764,In_1253,In_78);
xnor U765 (N_765,In_2160,In_284);
nand U766 (N_766,In_503,In_2145);
nand U767 (N_767,In_979,In_960);
nand U768 (N_768,In_930,In_2346);
and U769 (N_769,In_2221,In_2008);
or U770 (N_770,In_367,In_1236);
nand U771 (N_771,In_2126,In_1642);
or U772 (N_772,In_2208,In_435);
or U773 (N_773,In_455,In_1988);
and U774 (N_774,In_1916,In_1110);
and U775 (N_775,In_1656,In_1679);
xnor U776 (N_776,In_570,In_1585);
xnor U777 (N_777,In_2434,In_1292);
nand U778 (N_778,In_2270,In_2258);
nor U779 (N_779,In_383,In_621);
nor U780 (N_780,In_961,In_1597);
or U781 (N_781,In_1463,In_1074);
xnor U782 (N_782,In_1293,In_60);
and U783 (N_783,In_609,In_1556);
nor U784 (N_784,In_313,In_2348);
and U785 (N_785,In_783,In_2068);
or U786 (N_786,In_1516,In_878);
or U787 (N_787,In_2354,In_693);
nand U788 (N_788,In_90,In_644);
and U789 (N_789,In_1934,In_1634);
nor U790 (N_790,In_1546,In_1942);
and U791 (N_791,In_1304,In_1020);
xor U792 (N_792,In_293,In_1687);
nand U793 (N_793,In_112,In_1922);
nand U794 (N_794,In_1458,In_2001);
xor U795 (N_795,In_691,In_1593);
or U796 (N_796,In_148,In_1160);
nor U797 (N_797,In_2344,In_357);
nor U798 (N_798,In_1943,In_1066);
xnor U799 (N_799,In_55,In_734);
xnor U800 (N_800,In_1065,In_2460);
xnor U801 (N_801,In_2033,In_335);
nor U802 (N_802,In_2249,In_509);
or U803 (N_803,In_2083,In_1449);
xnor U804 (N_804,In_401,In_854);
xor U805 (N_805,In_1456,In_192);
nand U806 (N_806,In_85,In_2094);
nand U807 (N_807,In_1758,In_2104);
or U808 (N_808,In_1000,In_201);
nand U809 (N_809,In_712,In_560);
nor U810 (N_810,In_1834,In_241);
or U811 (N_811,In_1192,In_2130);
nor U812 (N_812,In_477,In_298);
nand U813 (N_813,In_1221,In_246);
nor U814 (N_814,In_1346,In_1623);
nand U815 (N_815,In_2327,In_733);
xnor U816 (N_816,In_909,In_837);
nor U817 (N_817,In_2232,In_2328);
xnor U818 (N_818,In_480,In_24);
xor U819 (N_819,In_1099,In_2418);
and U820 (N_820,In_427,In_419);
nand U821 (N_821,In_182,In_1083);
or U822 (N_822,In_1325,In_329);
xor U823 (N_823,In_1592,In_2210);
nand U824 (N_824,In_1577,In_384);
nand U825 (N_825,In_1739,In_1574);
and U826 (N_826,In_1016,In_2070);
or U827 (N_827,In_1571,In_688);
or U828 (N_828,In_841,In_124);
and U829 (N_829,In_645,In_436);
nand U830 (N_830,In_1420,In_2266);
nand U831 (N_831,In_1354,In_174);
nor U832 (N_832,In_1609,In_2119);
and U833 (N_833,In_687,In_1170);
xor U834 (N_834,In_1763,In_700);
nor U835 (N_835,In_104,In_873);
nand U836 (N_836,In_2385,In_2193);
nor U837 (N_837,In_1337,In_1183);
and U838 (N_838,In_2236,In_1345);
and U839 (N_839,In_829,In_1041);
xor U840 (N_840,In_485,In_207);
nor U841 (N_841,In_1275,In_1362);
and U842 (N_842,In_1307,In_1440);
and U843 (N_843,In_1226,In_2100);
nor U844 (N_844,In_699,In_1658);
nor U845 (N_845,In_235,In_1108);
nand U846 (N_846,In_1981,In_581);
nand U847 (N_847,In_1717,In_567);
or U848 (N_848,In_219,In_209);
and U849 (N_849,In_2064,In_1484);
and U850 (N_850,In_2499,In_996);
nand U851 (N_851,In_1674,In_950);
xor U852 (N_852,In_2185,In_2067);
nand U853 (N_853,In_1508,In_1507);
xnor U854 (N_854,In_964,In_1367);
xnor U855 (N_855,In_2398,In_1987);
or U856 (N_856,In_2243,In_107);
nor U857 (N_857,In_639,In_1618);
and U858 (N_858,In_629,In_525);
nor U859 (N_859,In_1690,In_2103);
and U860 (N_860,In_19,In_1397);
or U861 (N_861,In_551,In_359);
nand U862 (N_862,In_17,In_1651);
nand U863 (N_863,In_2304,In_2223);
or U864 (N_864,In_1753,In_518);
xor U865 (N_865,In_77,In_1986);
or U866 (N_866,In_1138,In_624);
nor U867 (N_867,In_1536,In_1792);
or U868 (N_868,In_338,In_1811);
nand U869 (N_869,In_1829,In_2323);
nor U870 (N_870,In_1754,In_1551);
and U871 (N_871,In_2254,In_597);
nor U872 (N_872,In_431,In_2458);
nor U873 (N_873,In_2409,In_1145);
and U874 (N_874,In_71,In_971);
xor U875 (N_875,In_1455,In_2022);
nor U876 (N_876,In_2436,In_2091);
nor U877 (N_877,In_2315,In_698);
or U878 (N_878,In_846,In_1560);
and U879 (N_879,In_389,In_1296);
and U880 (N_880,In_838,In_426);
nand U881 (N_881,In_1377,In_1373);
nand U882 (N_882,In_1341,In_211);
xnor U883 (N_883,In_2121,In_1730);
or U884 (N_884,In_572,In_714);
nand U885 (N_885,In_2318,In_1514);
xnor U886 (N_886,In_2152,In_627);
and U887 (N_887,In_165,In_1265);
and U888 (N_888,In_164,In_366);
xnor U889 (N_889,In_1502,In_2095);
nand U890 (N_890,In_1576,In_1869);
or U891 (N_891,In_245,In_2483);
xnor U892 (N_892,In_1928,In_989);
xnor U893 (N_893,In_399,In_2012);
nand U894 (N_894,In_937,In_983);
and U895 (N_895,In_65,In_224);
or U896 (N_896,In_1211,In_1129);
nand U897 (N_897,In_2329,In_408);
xor U898 (N_898,In_2416,In_1903);
and U899 (N_899,In_678,In_1760);
nand U900 (N_900,In_308,In_1063);
xor U901 (N_901,In_1935,In_1118);
nand U902 (N_902,In_916,In_195);
and U903 (N_903,In_1581,In_1904);
nor U904 (N_904,In_135,In_113);
or U905 (N_905,In_1649,In_2399);
nor U906 (N_906,In_2494,In_542);
and U907 (N_907,In_2299,In_2197);
nand U908 (N_908,In_855,In_1890);
xnor U909 (N_909,In_1851,In_173);
and U910 (N_910,In_1533,In_1930);
or U911 (N_911,In_1974,In_2055);
and U912 (N_912,In_2260,In_563);
or U913 (N_913,In_2107,In_2484);
nand U914 (N_914,In_2175,In_2367);
and U915 (N_915,In_2248,In_1998);
xnor U916 (N_916,In_2025,In_2106);
and U917 (N_917,In_788,In_1073);
or U918 (N_918,In_1509,In_2013);
nor U919 (N_919,In_2261,In_111);
nand U920 (N_920,In_1146,In_1043);
or U921 (N_921,In_385,In_452);
xor U922 (N_922,In_558,In_2394);
or U923 (N_923,In_1771,In_2333);
or U924 (N_924,In_2487,In_1734);
or U925 (N_925,In_605,In_1682);
xor U926 (N_926,In_321,In_1500);
and U927 (N_927,In_1262,In_194);
or U928 (N_928,In_1364,In_680);
or U929 (N_929,In_2040,In_1784);
nor U930 (N_930,In_1005,In_2230);
nand U931 (N_931,In_2093,In_295);
xnor U932 (N_932,In_2414,In_1819);
or U933 (N_933,In_668,In_1326);
xor U934 (N_934,In_206,In_618);
and U935 (N_935,In_637,In_755);
nor U936 (N_936,In_832,In_458);
nand U937 (N_937,In_167,In_1070);
xnor U938 (N_938,In_1561,In_651);
nor U939 (N_939,In_2081,In_2195);
nand U940 (N_940,In_230,In_414);
and U941 (N_941,In_1552,In_620);
and U942 (N_942,In_240,In_2125);
and U943 (N_943,In_1522,In_1515);
xnor U944 (N_944,In_1271,In_1283);
or U945 (N_945,In_1720,In_611);
nand U946 (N_946,In_2431,In_449);
or U947 (N_947,In_819,In_1352);
xor U948 (N_948,In_2491,In_764);
nand U949 (N_949,In_220,In_897);
and U950 (N_950,In_2041,In_120);
xor U951 (N_951,In_2422,In_101);
nand U952 (N_952,In_1582,In_1572);
or U953 (N_953,In_1036,In_835);
or U954 (N_954,In_496,In_2357);
nor U955 (N_955,In_1595,In_754);
and U956 (N_956,In_288,In_1941);
nand U957 (N_957,In_633,In_1313);
or U958 (N_958,In_2404,In_2201);
nor U959 (N_959,In_1989,In_1379);
and U960 (N_960,In_374,In_573);
nor U961 (N_961,In_526,In_1327);
xor U962 (N_962,In_1026,In_1451);
nor U963 (N_963,In_2334,In_478);
xnor U964 (N_964,In_193,In_1139);
and U965 (N_965,In_1525,In_619);
nand U966 (N_966,In_784,In_1126);
and U967 (N_967,In_2129,In_759);
and U968 (N_968,In_904,In_1900);
xor U969 (N_969,In_334,In_2415);
nand U970 (N_970,In_337,In_1245);
nand U971 (N_971,In_2061,In_1589);
nand U972 (N_972,In_1059,In_2148);
and U973 (N_973,In_1915,In_601);
xnor U974 (N_974,In_1294,In_1242);
nor U975 (N_975,In_26,In_1318);
or U976 (N_976,In_758,In_118);
nor U977 (N_977,In_896,In_1727);
and U978 (N_978,In_590,In_2295);
xor U979 (N_979,In_1606,In_756);
or U980 (N_980,In_519,In_2049);
and U981 (N_981,In_1147,In_1077);
nor U982 (N_982,In_2343,In_953);
nand U983 (N_983,In_1295,In_886);
and U984 (N_984,In_1818,In_2123);
xnor U985 (N_985,In_1564,In_1357);
and U986 (N_986,In_2132,In_251);
and U987 (N_987,In_1324,In_1436);
and U988 (N_988,In_2282,In_2176);
xor U989 (N_989,In_2496,In_1787);
and U990 (N_990,In_1194,In_88);
and U991 (N_991,In_2021,In_1323);
or U992 (N_992,In_2019,In_600);
and U993 (N_993,In_199,In_1387);
xnor U994 (N_994,In_2057,In_828);
or U995 (N_995,In_2296,In_1018);
nand U996 (N_996,In_2217,In_750);
or U997 (N_997,In_67,In_205);
xnor U998 (N_998,In_215,In_987);
and U999 (N_999,In_652,In_1608);
or U1000 (N_1000,N_216,N_168);
xor U1001 (N_1001,In_2042,N_97);
xnor U1002 (N_1002,N_99,In_1995);
xnor U1003 (N_1003,In_2194,In_2380);
nor U1004 (N_1004,In_2059,N_347);
nand U1005 (N_1005,N_475,In_446);
xor U1006 (N_1006,N_290,N_352);
or U1007 (N_1007,In_117,N_632);
nor U1008 (N_1008,N_248,In_510);
nor U1009 (N_1009,N_10,N_678);
xor U1010 (N_1010,N_425,N_780);
and U1011 (N_1011,N_220,N_981);
and U1012 (N_1012,N_696,N_64);
nand U1013 (N_1013,In_1766,N_25);
or U1014 (N_1014,N_584,In_1439);
or U1015 (N_1015,N_138,N_844);
xnor U1016 (N_1016,In_1635,N_122);
nand U1017 (N_1017,N_969,In_336);
xnor U1018 (N_1018,N_803,N_883);
or U1019 (N_1019,N_721,N_51);
and U1020 (N_1020,N_284,N_676);
nand U1021 (N_1021,In_50,N_337);
or U1022 (N_1022,N_386,N_467);
or U1023 (N_1023,N_599,N_809);
or U1024 (N_1024,In_968,In_1686);
nand U1025 (N_1025,In_1991,N_645);
and U1026 (N_1026,N_324,In_893);
or U1027 (N_1027,N_746,N_693);
and U1028 (N_1028,N_956,N_485);
nand U1029 (N_1029,In_1374,N_848);
nor U1030 (N_1030,N_326,N_989);
nand U1031 (N_1031,N_306,N_255);
nand U1032 (N_1032,N_542,N_967);
nor U1033 (N_1033,N_266,In_932);
and U1034 (N_1034,In_1775,N_633);
nor U1035 (N_1035,In_1181,In_528);
or U1036 (N_1036,N_235,N_741);
or U1037 (N_1037,In_1894,N_186);
and U1038 (N_1038,N_373,In_239);
nor U1039 (N_1039,In_473,N_279);
nor U1040 (N_1040,In_931,N_90);
or U1041 (N_1041,N_105,In_724);
xnor U1042 (N_1042,In_1866,In_1871);
nor U1043 (N_1043,N_813,N_655);
or U1044 (N_1044,In_2461,In_418);
nand U1045 (N_1045,In_443,N_217);
nand U1046 (N_1046,In_170,In_1863);
and U1047 (N_1047,N_260,N_995);
nand U1048 (N_1048,In_2,N_408);
or U1049 (N_1049,N_999,N_986);
nor U1050 (N_1050,N_3,N_901);
xor U1051 (N_1051,N_406,N_191);
xor U1052 (N_1052,N_502,In_2350);
xnor U1053 (N_1053,N_582,N_963);
or U1054 (N_1054,In_2291,In_274);
xor U1055 (N_1055,N_32,N_145);
and U1056 (N_1056,N_973,N_635);
and U1057 (N_1057,N_647,N_836);
nand U1058 (N_1058,In_1554,N_244);
nand U1059 (N_1059,In_213,In_655);
or U1060 (N_1060,N_938,N_313);
or U1061 (N_1061,N_81,N_501);
nor U1062 (N_1062,N_157,N_177);
or U1063 (N_1063,N_792,N_155);
and U1064 (N_1064,N_785,N_589);
and U1065 (N_1065,In_1669,N_575);
or U1066 (N_1066,N_144,N_802);
or U1067 (N_1067,In_1003,N_855);
and U1068 (N_1068,In_437,In_1351);
xor U1069 (N_1069,In_1994,In_265);
xor U1070 (N_1070,In_2411,In_1583);
xnor U1071 (N_1071,N_604,N_551);
and U1072 (N_1072,N_513,N_56);
xnor U1073 (N_1073,N_935,N_766);
xor U1074 (N_1074,N_779,In_1132);
xnor U1075 (N_1075,N_682,N_629);
xnor U1076 (N_1076,In_926,N_311);
nor U1077 (N_1077,N_778,In_1898);
nor U1078 (N_1078,N_85,N_865);
and U1079 (N_1079,N_438,N_763);
nor U1080 (N_1080,N_190,In_2312);
nand U1081 (N_1081,N_309,N_98);
nand U1082 (N_1082,N_601,In_469);
nor U1083 (N_1083,N_281,N_600);
nor U1084 (N_1084,In_1862,In_2277);
xor U1085 (N_1085,N_256,N_359);
nand U1086 (N_1086,N_671,In_2433);
xnor U1087 (N_1087,In_1025,N_812);
or U1088 (N_1088,N_932,N_358);
xor U1089 (N_1089,N_821,N_764);
xnor U1090 (N_1090,N_641,N_718);
nand U1091 (N_1091,N_243,N_203);
and U1092 (N_1092,N_499,In_123);
nand U1093 (N_1093,In_326,N_732);
nor U1094 (N_1094,In_2457,In_2473);
nor U1095 (N_1095,In_1709,N_118);
nand U1096 (N_1096,N_623,N_468);
and U1097 (N_1097,In_2271,In_595);
xor U1098 (N_1098,N_831,In_1011);
xnor U1099 (N_1099,N_783,In_1017);
nor U1100 (N_1100,N_903,In_1559);
nand U1101 (N_1101,N_918,N_557);
nor U1102 (N_1102,N_957,N_452);
nor U1103 (N_1103,N_278,N_751);
nor U1104 (N_1104,N_464,N_34);
xnor U1105 (N_1105,N_247,N_919);
and U1106 (N_1106,N_461,In_1846);
or U1107 (N_1107,In_511,In_549);
nand U1108 (N_1108,N_276,In_2028);
and U1109 (N_1109,N_136,N_856);
or U1110 (N_1110,In_796,N_443);
nor U1111 (N_1111,N_885,In_1291);
or U1112 (N_1112,N_710,In_1586);
nand U1113 (N_1113,N_758,N_389);
nand U1114 (N_1114,In_1348,N_677);
nand U1115 (N_1115,N_148,N_941);
nand U1116 (N_1116,In_1302,N_165);
and U1117 (N_1117,N_39,N_598);
xor U1118 (N_1118,N_355,N_992);
nand U1119 (N_1119,In_707,N_556);
xnor U1120 (N_1120,In_1487,N_170);
nor U1121 (N_1121,N_315,N_384);
nor U1122 (N_1122,In_709,N_36);
nor U1123 (N_1123,N_784,N_159);
xnor U1124 (N_1124,N_448,In_2089);
and U1125 (N_1125,N_289,N_158);
nand U1126 (N_1126,In_810,N_178);
xor U1127 (N_1127,N_22,In_476);
or U1128 (N_1128,In_1696,In_587);
and U1129 (N_1129,In_13,N_73);
and U1130 (N_1130,In_76,In_2410);
nand U1131 (N_1131,N_160,N_88);
or U1132 (N_1132,N_454,N_492);
or U1133 (N_1133,N_788,In_866);
and U1134 (N_1134,N_879,In_3);
xor U1135 (N_1135,N_111,In_441);
or U1136 (N_1136,In_2426,N_265);
or U1137 (N_1137,N_429,In_580);
or U1138 (N_1138,In_388,N_712);
nor U1139 (N_1139,N_737,In_1768);
nand U1140 (N_1140,In_706,In_1542);
and U1141 (N_1141,N_924,N_862);
or U1142 (N_1142,N_595,In_685);
nor U1143 (N_1143,N_922,N_53);
nor U1144 (N_1144,In_508,N_724);
nand U1145 (N_1145,N_615,N_307);
xor U1146 (N_1146,N_466,In_258);
nand U1147 (N_1147,N_692,In_2184);
xnor U1148 (N_1148,In_880,In_923);
xor U1149 (N_1149,N_45,N_261);
and U1150 (N_1150,N_297,N_605);
nand U1151 (N_1151,N_330,N_977);
or U1152 (N_1152,N_867,In_763);
nor U1153 (N_1153,N_555,N_670);
nor U1154 (N_1154,N_2,N_790);
nor U1155 (N_1155,N_698,In_1803);
nor U1156 (N_1156,N_344,In_2417);
nand U1157 (N_1157,N_985,N_62);
nor U1158 (N_1158,In_844,N_644);
and U1159 (N_1159,N_701,In_1719);
nand U1160 (N_1160,In_166,N_767);
xnor U1161 (N_1161,N_1,N_562);
and U1162 (N_1162,N_5,In_1493);
and U1163 (N_1163,N_816,N_747);
and U1164 (N_1164,N_121,N_565);
nor U1165 (N_1165,In_1990,In_1676);
nor U1166 (N_1166,N_777,N_907);
and U1167 (N_1167,N_880,In_346);
nor U1168 (N_1168,N_236,In_2237);
xor U1169 (N_1169,N_343,In_1962);
or U1170 (N_1170,In_1697,In_1638);
and U1171 (N_1171,N_317,N_368);
nand U1172 (N_1172,N_868,N_954);
nor U1173 (N_1173,N_338,N_776);
or U1174 (N_1174,N_453,N_881);
nand U1175 (N_1175,N_35,N_46);
and U1176 (N_1176,In_269,In_2180);
and U1177 (N_1177,N_528,N_292);
or U1178 (N_1178,In_1277,N_736);
and U1179 (N_1179,N_752,N_199);
nor U1180 (N_1180,N_971,N_731);
or U1181 (N_1181,N_574,N_87);
xnor U1182 (N_1182,N_818,In_1176);
xnor U1183 (N_1183,N_320,N_583);
nor U1184 (N_1184,N_196,In_571);
nor U1185 (N_1185,In_261,In_1336);
xor U1186 (N_1186,N_639,N_817);
xnor U1187 (N_1187,In_1601,N_876);
nand U1188 (N_1188,In_1411,N_13);
or U1189 (N_1189,In_684,N_411);
nand U1190 (N_1190,N_152,In_196);
xor U1191 (N_1191,In_1780,In_1523);
nor U1192 (N_1192,In_1090,N_327);
xnor U1193 (N_1193,N_852,N_833);
and U1194 (N_1194,N_205,N_651);
and U1195 (N_1195,In_577,N_987);
and U1196 (N_1196,N_192,In_610);
xor U1197 (N_1197,N_195,In_30);
and U1198 (N_1198,In_1844,N_695);
nand U1199 (N_1199,N_472,N_681);
or U1200 (N_1200,N_234,N_318);
or U1201 (N_1201,In_129,N_240);
and U1202 (N_1202,N_331,N_875);
or U1203 (N_1203,In_1082,N_251);
nand U1204 (N_1204,N_913,In_1344);
and U1205 (N_1205,N_937,In_2308);
nand U1206 (N_1206,N_376,N_208);
nand U1207 (N_1207,N_184,N_340);
or U1208 (N_1208,In_352,In_2268);
xor U1209 (N_1209,In_2045,N_805);
or U1210 (N_1210,N_7,N_700);
and U1211 (N_1211,N_274,N_960);
nor U1212 (N_1212,N_864,In_354);
nand U1213 (N_1213,N_976,In_1532);
and U1214 (N_1214,N_891,N_15);
and U1215 (N_1215,In_1450,N_239);
nand U1216 (N_1216,N_460,In_974);
or U1217 (N_1217,N_726,N_462);
and U1218 (N_1218,N_674,N_67);
xnor U1219 (N_1219,N_106,N_378);
and U1220 (N_1220,N_518,N_544);
nand U1221 (N_1221,N_892,N_588);
nand U1222 (N_1222,N_70,N_939);
nand U1223 (N_1223,N_720,N_263);
xnor U1224 (N_1224,In_1481,N_441);
or U1225 (N_1225,N_925,N_154);
xor U1226 (N_1226,In_131,In_825);
nand U1227 (N_1227,In_2150,N_500);
or U1228 (N_1228,In_1309,In_380);
and U1229 (N_1229,N_798,N_760);
and U1230 (N_1230,N_79,N_546);
nor U1231 (N_1231,In_1363,N_893);
and U1232 (N_1232,N_82,N_944);
or U1233 (N_1233,N_611,In_548);
xor U1234 (N_1234,N_962,N_351);
or U1235 (N_1235,In_2224,In_1891);
xor U1236 (N_1236,In_1480,In_534);
nand U1237 (N_1237,N_402,N_447);
and U1238 (N_1238,In_1311,N_275);
xnor U1239 (N_1239,N_863,In_1680);
nor U1240 (N_1240,N_568,N_765);
nor U1241 (N_1241,N_287,N_272);
xnor U1242 (N_1242,N_223,N_364);
nor U1243 (N_1243,N_426,In_1911);
nor U1244 (N_1244,N_38,In_1681);
and U1245 (N_1245,N_446,N_455);
or U1246 (N_1246,N_346,N_839);
xor U1247 (N_1247,N_659,N_543);
nand U1248 (N_1248,N_416,In_1675);
nand U1249 (N_1249,N_808,N_689);
nand U1250 (N_1250,N_725,N_280);
xor U1251 (N_1251,In_917,In_521);
nand U1252 (N_1252,N_249,In_1925);
or U1253 (N_1253,N_666,N_590);
nor U1254 (N_1254,In_1111,In_1173);
or U1255 (N_1255,N_811,N_607);
or U1256 (N_1256,N_908,N_303);
xor U1257 (N_1257,In_1285,N_743);
nor U1258 (N_1258,N_254,N_768);
and U1259 (N_1259,In_302,N_914);
and U1260 (N_1260,N_733,N_224);
nor U1261 (N_1261,N_636,N_702);
or U1262 (N_1262,In_1539,N_484);
nor U1263 (N_1263,In_2239,In_513);
or U1264 (N_1264,In_1955,N_827);
xor U1265 (N_1265,In_450,N_112);
nor U1266 (N_1266,N_807,In_1530);
xor U1267 (N_1267,N_591,N_44);
and U1268 (N_1268,N_614,N_762);
nand U1269 (N_1269,In_1594,N_508);
and U1270 (N_1270,N_124,N_654);
nand U1271 (N_1271,In_741,In_1854);
or U1272 (N_1272,In_1392,In_2381);
or U1273 (N_1273,N_91,N_688);
xnor U1274 (N_1274,N_356,N_246);
and U1275 (N_1275,N_397,In_1701);
nand U1276 (N_1276,In_1426,N_694);
xnor U1277 (N_1277,N_68,N_42);
nor U1278 (N_1278,In_2141,N_873);
and U1279 (N_1279,N_902,In_2222);
xnor U1280 (N_1280,N_434,N_319);
or U1281 (N_1281,In_1541,N_299);
nor U1282 (N_1282,In_966,N_127);
and U1283 (N_1283,In_1772,N_470);
and U1284 (N_1284,N_841,In_311);
nand U1285 (N_1285,N_262,N_755);
nand U1286 (N_1286,N_819,N_396);
xor U1287 (N_1287,N_350,N_237);
and U1288 (N_1288,N_535,N_975);
nand U1289 (N_1289,In_1801,In_1429);
or U1290 (N_1290,N_581,N_179);
or U1291 (N_1291,N_866,In_1644);
nand U1292 (N_1292,N_961,N_212);
or U1293 (N_1293,In_1418,N_314);
or U1294 (N_1294,N_65,N_146);
or U1295 (N_1295,N_577,N_520);
nand U1296 (N_1296,N_722,N_738);
or U1297 (N_1297,N_822,In_481);
nor U1298 (N_1298,In_2246,N_643);
nand U1299 (N_1299,N_321,N_398);
nand U1300 (N_1300,N_395,N_853);
and U1301 (N_1301,In_456,N_167);
and U1302 (N_1302,In_606,N_377);
or U1303 (N_1303,N_569,N_705);
nor U1304 (N_1304,In_502,N_6);
nand U1305 (N_1305,N_305,N_794);
or U1306 (N_1306,N_801,In_1545);
or U1307 (N_1307,N_510,N_909);
xnor U1308 (N_1308,N_672,In_530);
nor U1309 (N_1309,N_310,In_593);
nor U1310 (N_1310,In_2293,N_690);
nand U1311 (N_1311,N_187,In_2358);
and U1312 (N_1312,N_229,N_727);
or U1313 (N_1313,N_89,N_874);
xor U1314 (N_1314,In_420,N_637);
or U1315 (N_1315,N_55,N_4);
or U1316 (N_1316,N_516,In_859);
nand U1317 (N_1317,N_877,N_210);
and U1318 (N_1318,In_287,In_1208);
and U1319 (N_1319,N_950,N_750);
xor U1320 (N_1320,N_537,In_172);
xnor U1321 (N_1321,N_483,In_1178);
nor U1322 (N_1322,In_1142,N_459);
and U1323 (N_1323,N_394,N_990);
nor U1324 (N_1324,N_233,N_172);
nor U1325 (N_1325,In_1359,N_618);
and U1326 (N_1326,N_488,N_498);
nand U1327 (N_1327,In_2162,N_509);
and U1328 (N_1328,In_1150,N_214);
xnor U1329 (N_1329,N_799,N_649);
or U1330 (N_1330,N_421,N_619);
xor U1331 (N_1331,N_800,In_1185);
nor U1332 (N_1332,N_564,In_1885);
nand U1333 (N_1333,N_29,N_380);
and U1334 (N_1334,N_628,In_1823);
or U1335 (N_1335,N_997,N_58);
or U1336 (N_1336,In_474,N_113);
xor U1337 (N_1337,In_1613,N_30);
nor U1338 (N_1338,N_882,N_334);
nand U1339 (N_1339,N_424,N_930);
or U1340 (N_1340,In_2405,In_2353);
or U1341 (N_1341,N_838,N_432);
nor U1342 (N_1342,In_791,In_1365);
and U1343 (N_1343,In_1068,N_753);
xnor U1344 (N_1344,N_849,N_433);
nor U1345 (N_1345,N_409,N_436);
nor U1346 (N_1346,N_795,In_1750);
xnor U1347 (N_1347,In_2079,In_2202);
nand U1348 (N_1348,N_910,In_682);
or U1349 (N_1349,N_156,N_129);
nor U1350 (N_1350,In_316,N_360);
and U1351 (N_1351,N_567,N_285);
nor U1352 (N_1352,N_585,N_739);
xor U1353 (N_1353,N_20,In_919);
nor U1354 (N_1354,In_661,In_818);
and U1355 (N_1355,N_415,N_558);
nor U1356 (N_1356,N_18,In_1466);
nor U1357 (N_1357,In_705,N_563);
xor U1358 (N_1358,N_806,N_664);
xnor U1359 (N_1359,N_295,N_714);
and U1360 (N_1360,N_942,N_829);
nor U1361 (N_1361,N_665,In_1237);
or U1362 (N_1362,N_531,In_1210);
xor U1363 (N_1363,In_1694,N_218);
or U1364 (N_1364,N_850,N_71);
or U1365 (N_1365,N_198,N_328);
nand U1366 (N_1366,N_840,In_1711);
nor U1367 (N_1367,N_414,N_923);
xnor U1368 (N_1368,N_390,N_401);
xnor U1369 (N_1369,N_851,N_456);
nand U1370 (N_1370,N_708,N_781);
xor U1371 (N_1371,In_1380,N_17);
nor U1372 (N_1372,N_222,N_94);
or U1373 (N_1373,N_617,N_114);
or U1374 (N_1374,N_370,N_580);
and U1375 (N_1375,N_391,In_1109);
xor U1376 (N_1376,N_921,N_625);
and U1377 (N_1377,In_278,N_435);
nor U1378 (N_1378,In_1338,N_474);
nor U1379 (N_1379,N_37,N_288);
or U1380 (N_1380,In_720,N_660);
and U1381 (N_1381,N_412,In_2122);
and U1382 (N_1382,N_43,In_1707);
or U1383 (N_1383,N_872,N_616);
or U1384 (N_1384,In_1273,N_592);
or U1385 (N_1385,N_329,N_526);
or U1386 (N_1386,N_169,N_715);
xor U1387 (N_1387,In_2374,In_1078);
nor U1388 (N_1388,N_573,N_23);
nand U1389 (N_1389,In_1664,N_52);
and U1390 (N_1390,N_570,In_674);
nor U1391 (N_1391,In_2053,N_115);
or U1392 (N_1392,N_723,In_472);
and U1393 (N_1393,N_457,N_703);
xor U1394 (N_1394,In_2402,In_914);
and U1395 (N_1395,N_594,In_332);
nor U1396 (N_1396,In_638,In_2382);
and U1397 (N_1397,N_940,In_1738);
xor U1398 (N_1398,In_1867,N_130);
and U1399 (N_1399,N_57,N_140);
nand U1400 (N_1400,N_602,N_860);
or U1401 (N_1401,N_374,In_1096);
nand U1402 (N_1402,N_194,N_163);
and U1403 (N_1403,In_833,In_1888);
or U1404 (N_1404,In_544,N_953);
and U1405 (N_1405,N_787,In_667);
or U1406 (N_1406,In_31,In_543);
nor U1407 (N_1407,N_523,N_810);
or U1408 (N_1408,N_449,N_361);
or U1409 (N_1409,N_984,In_2313);
and U1410 (N_1410,N_587,N_837);
and U1411 (N_1411,N_471,N_161);
xor U1412 (N_1412,In_671,In_1547);
xor U1413 (N_1413,N_171,In_39);
and U1414 (N_1414,In_1490,In_4);
or U1415 (N_1415,N_988,N_182);
nor U1416 (N_1416,In_2138,In_2211);
xnor U1417 (N_1417,In_767,In_342);
or U1418 (N_1418,N_325,N_597);
nand U1419 (N_1419,N_610,N_19);
or U1420 (N_1420,In_1402,N_952);
or U1421 (N_1421,N_173,In_1435);
nor U1422 (N_1422,In_468,N_928);
xnor U1423 (N_1423,N_630,In_1032);
xnor U1424 (N_1424,In_1120,In_772);
and U1425 (N_1425,N_662,N_884);
and U1426 (N_1426,N_333,In_2168);
nand U1427 (N_1427,N_561,In_1752);
nor U1428 (N_1428,In_1329,In_696);
or U1429 (N_1429,In_725,In_540);
or U1430 (N_1430,N_532,N_428);
and U1431 (N_1431,In_1406,In_1693);
or U1432 (N_1432,In_283,N_257);
nand U1433 (N_1433,In_956,In_749);
and U1434 (N_1434,N_545,N_126);
and U1435 (N_1435,N_252,N_400);
nand U1436 (N_1436,N_835,N_540);
or U1437 (N_1437,In_1268,N_354);
nand U1438 (N_1438,N_141,N_209);
and U1439 (N_1439,N_797,N_871);
and U1440 (N_1440,In_501,In_1417);
nor U1441 (N_1441,N_974,N_202);
or U1442 (N_1442,N_119,N_603);
and U1443 (N_1443,N_440,N_189);
or U1444 (N_1444,N_418,N_709);
and U1445 (N_1445,In_1907,N_480);
nand U1446 (N_1446,N_539,N_661);
nor U1447 (N_1447,In_1217,N_994);
and U1448 (N_1448,In_834,N_175);
or U1449 (N_1449,In_1388,N_832);
and U1450 (N_1450,In_2005,N_21);
or U1451 (N_1451,N_745,N_711);
xor U1452 (N_1452,In_266,N_153);
or U1453 (N_1453,N_646,N_72);
or U1454 (N_1454,In_1964,In_978);
xnor U1455 (N_1455,N_282,N_296);
xnor U1456 (N_1456,In_1786,N_686);
xnor U1457 (N_1457,In_2229,N_342);
nand U1458 (N_1458,In_1469,In_483);
nand U1459 (N_1459,In_773,N_291);
nand U1460 (N_1460,In_2456,N_147);
or U1461 (N_1461,N_519,In_736);
and U1462 (N_1462,In_281,In_1300);
nand U1463 (N_1463,N_900,N_497);
nand U1464 (N_1464,N_365,In_2438);
nor U1465 (N_1465,N_770,N_897);
or U1466 (N_1466,N_270,N_571);
nor U1467 (N_1467,In_1643,N_385);
or U1468 (N_1468,N_522,In_115);
and U1469 (N_1469,N_300,N_123);
nand U1470 (N_1470,In_986,N_238);
or U1471 (N_1471,N_357,N_135);
xnor U1472 (N_1472,N_773,In_2109);
nor U1473 (N_1473,N_566,N_9);
nand U1474 (N_1474,N_463,N_652);
xor U1475 (N_1475,In_2253,N_505);
nor U1476 (N_1476,N_59,N_669);
xor U1477 (N_1477,N_185,In_475);
and U1478 (N_1478,N_366,N_744);
or U1479 (N_1479,N_620,N_0);
xnor U1480 (N_1480,In_2147,N_174);
and U1481 (N_1481,In_779,In_1485);
xor U1482 (N_1482,N_399,In_1029);
xnor U1483 (N_1483,In_1274,In_2240);
and U1484 (N_1484,In_259,N_66);
or U1485 (N_1485,In_1298,N_204);
and U1486 (N_1486,N_525,N_176);
nor U1487 (N_1487,In_1627,N_658);
nand U1488 (N_1488,In_2062,N_477);
xnor U1489 (N_1489,N_60,N_323);
and U1490 (N_1490,N_609,N_993);
nor U1491 (N_1491,N_572,In_396);
nand U1492 (N_1492,In_1100,In_2371);
and U1493 (N_1493,N_381,N_998);
or U1494 (N_1494,N_857,N_54);
nand U1495 (N_1495,N_363,N_26);
xnor U1496 (N_1496,In_2032,N_107);
nor U1497 (N_1497,In_2174,N_943);
and U1498 (N_1498,In_1191,In_2173);
or U1499 (N_1499,In_1214,N_886);
and U1500 (N_1500,N_142,N_920);
xnor U1501 (N_1501,N_14,N_393);
nor U1502 (N_1502,N_707,In_2216);
nor U1503 (N_1503,In_2459,N_634);
nand U1504 (N_1504,N_527,N_201);
nand U1505 (N_1505,In_1027,In_1207);
xnor U1506 (N_1506,N_84,N_815);
nand U1507 (N_1507,N_521,N_286);
and U1508 (N_1508,N_912,In_2102);
or U1509 (N_1509,N_367,In_1279);
or U1510 (N_1510,N_858,N_151);
and U1511 (N_1511,In_630,In_1372);
xnor U1512 (N_1512,N_524,In_993);
nand U1513 (N_1513,N_756,N_859);
or U1514 (N_1514,In_37,N_627);
xor U1515 (N_1515,In_1457,N_258);
nand U1516 (N_1516,In_666,N_996);
nand U1517 (N_1517,N_972,In_155);
and U1518 (N_1518,N_916,N_225);
nand U1519 (N_1519,In_2462,N_231);
nor U1520 (N_1520,N_444,In_1762);
and U1521 (N_1521,N_245,N_469);
xnor U1522 (N_1522,N_308,N_259);
xnor U1523 (N_1523,N_814,In_2292);
nor U1524 (N_1524,N_869,In_1820);
nor U1525 (N_1525,In_1881,N_417);
xnor U1526 (N_1526,N_775,In_569);
xor U1527 (N_1527,In_1496,N_298);
nor U1528 (N_1528,N_946,N_890);
and U1529 (N_1529,N_951,In_369);
xor U1530 (N_1530,N_109,N_339);
nand U1531 (N_1531,N_250,In_1006);
nand U1532 (N_1532,In_1756,N_697);
nor U1533 (N_1533,N_423,In_1091);
nand U1534 (N_1534,N_133,N_656);
xor U1535 (N_1535,N_547,In_1159);
nor U1536 (N_1536,N_28,N_131);
nand U1537 (N_1537,In_2000,In_440);
and U1538 (N_1538,In_2468,In_2192);
and U1539 (N_1539,N_979,N_489);
or U1540 (N_1540,N_451,N_895);
and U1541 (N_1541,N_959,N_541);
nand U1542 (N_1542,In_1875,In_1921);
xnor U1543 (N_1543,N_716,In_1543);
or U1544 (N_1544,N_679,N_422);
and U1545 (N_1545,In_262,In_1795);
and U1546 (N_1546,N_887,N_302);
xor U1547 (N_1547,N_241,N_622);
nor U1548 (N_1548,N_104,N_215);
nor U1549 (N_1549,N_668,In_663);
nor U1550 (N_1550,N_754,N_495);
and U1551 (N_1551,N_948,N_899);
or U1552 (N_1552,N_640,In_1767);
or U1553 (N_1553,N_180,In_16);
or U1554 (N_1554,N_947,In_739);
or U1555 (N_1555,N_847,N_442);
xnor U1556 (N_1556,N_271,N_143);
and U1557 (N_1557,In_1746,N_917);
xor U1558 (N_1558,N_650,In_2397);
or U1559 (N_1559,N_102,In_622);
nand U1560 (N_1560,N_12,In_1842);
and U1561 (N_1561,N_137,N_786);
or U1562 (N_1562,N_47,N_369);
or U1563 (N_1563,N_734,N_188);
nor U1564 (N_1564,In_1889,N_823);
or U1565 (N_1565,In_48,In_1452);
and U1566 (N_1566,N_949,N_529);
and U1567 (N_1567,In_180,N_536);
nor U1568 (N_1568,In_1260,N_405);
or U1569 (N_1569,N_478,N_970);
nand U1570 (N_1570,N_117,N_40);
and U1571 (N_1571,N_904,N_162);
and U1572 (N_1572,N_578,N_503);
nand U1573 (N_1573,N_232,N_978);
and U1574 (N_1574,N_704,In_602);
and U1575 (N_1575,N_684,N_404);
xnor U1576 (N_1576,In_1252,N_663);
or U1577 (N_1577,N_789,N_253);
and U1578 (N_1578,N_322,In_1505);
xnor U1579 (N_1579,N_403,N_530);
nand U1580 (N_1580,N_889,In_320);
and U1581 (N_1581,N_61,In_1926);
or U1582 (N_1582,N_101,N_86);
nand U1583 (N_1583,In_1156,In_1119);
and U1584 (N_1584,N_379,N_538);
or U1585 (N_1585,N_268,In_539);
xor U1586 (N_1586,N_490,N_514);
nor U1587 (N_1587,N_496,N_473);
and U1588 (N_1588,N_683,In_2453);
nand U1589 (N_1589,In_872,In_263);
nand U1590 (N_1590,In_2071,N_699);
or U1591 (N_1591,N_273,N_894);
nand U1592 (N_1592,N_507,N_820);
nand U1593 (N_1593,In_1788,N_120);
or U1594 (N_1594,In_1050,In_1673);
nand U1595 (N_1595,N_830,N_332);
or U1596 (N_1596,N_16,In_1802);
xnor U1597 (N_1597,N_491,In_1757);
and U1598 (N_1598,N_667,N_878);
xnor U1599 (N_1599,In_683,In_943);
xnor U1600 (N_1600,N_828,In_1657);
xnor U1601 (N_1601,N_181,In_500);
nor U1602 (N_1602,In_1706,N_653);
nand U1603 (N_1603,In_2267,N_958);
and U1604 (N_1604,N_606,N_933);
or U1605 (N_1605,N_934,N_729);
nand U1606 (N_1606,In_1912,N_430);
or U1607 (N_1607,In_1347,N_965);
nand U1608 (N_1608,In_1910,N_312);
and U1609 (N_1609,N_69,N_929);
xnor U1610 (N_1610,N_458,N_139);
xnor U1611 (N_1611,N_277,N_166);
xnor U1612 (N_1612,N_533,N_431);
nand U1613 (N_1613,In_121,N_713);
nand U1614 (N_1614,In_2214,N_730);
and U1615 (N_1615,N_294,N_772);
nor U1616 (N_1616,N_769,In_339);
and U1617 (N_1617,N_193,N_896);
or U1618 (N_1618,N_226,N_372);
xnor U1619 (N_1619,In_2373,In_625);
or U1620 (N_1620,N_675,N_685);
xnor U1621 (N_1621,N_548,In_14);
or U1622 (N_1622,N_24,N_132);
and U1623 (N_1623,N_116,N_771);
and U1624 (N_1624,N_931,N_479);
nand U1625 (N_1625,N_748,In_731);
and U1626 (N_1626,N_517,In_147);
nor U1627 (N_1627,N_96,N_717);
and U1628 (N_1628,In_2492,In_1308);
or U1629 (N_1629,N_83,N_631);
nand U1630 (N_1630,N_427,In_1089);
nand U1631 (N_1631,N_906,N_966);
and U1632 (N_1632,In_1781,N_382);
xnor U1633 (N_1633,N_74,N_657);
nor U1634 (N_1634,N_576,In_1405);
xor U1635 (N_1635,N_596,N_11);
nor U1636 (N_1636,N_345,N_63);
or U1637 (N_1637,N_854,In_1204);
and U1638 (N_1638,N_608,N_392);
nand U1639 (N_1639,In_817,N_774);
and U1640 (N_1640,In_1290,N_846);
nand U1641 (N_1641,N_197,N_75);
nand U1642 (N_1642,N_719,In_574);
or U1643 (N_1643,In_665,N_964);
nor U1644 (N_1644,In_445,N_183);
and U1645 (N_1645,In_703,N_48);
nor U1646 (N_1646,N_735,N_200);
nand U1647 (N_1647,In_1034,N_861);
and U1648 (N_1648,N_559,N_945);
xnor U1649 (N_1649,N_335,N_553);
or U1650 (N_1650,In_1286,N_230);
or U1651 (N_1651,In_248,N_41);
nor U1652 (N_1652,In_2011,N_349);
and U1653 (N_1653,In_417,In_492);
nand U1654 (N_1654,N_487,N_341);
and U1655 (N_1655,In_1107,In_1665);
xnor U1656 (N_1656,N_826,In_1314);
or U1657 (N_1657,N_164,In_1512);
xor U1658 (N_1658,N_437,In_1839);
or U1659 (N_1659,In_803,N_982);
nor U1660 (N_1660,In_1157,N_968);
or U1661 (N_1661,N_482,In_1259);
xnor U1662 (N_1662,N_825,In_626);
nand U1663 (N_1663,N_486,N_749);
nand U1664 (N_1664,N_465,N_387);
nand U1665 (N_1665,N_804,N_445);
xor U1666 (N_1666,In_1232,N_742);
nand U1667 (N_1667,N_936,In_792);
and U1668 (N_1668,N_80,N_560);
or U1669 (N_1669,N_77,In_457);
nor U1670 (N_1670,N_845,N_450);
nor U1671 (N_1671,N_413,In_1870);
nor U1672 (N_1672,N_31,N_125);
and U1673 (N_1673,N_991,In_210);
xor U1674 (N_1674,In_648,N_691);
and U1675 (N_1675,N_301,N_304);
xnor U1676 (N_1676,N_481,N_980);
or U1677 (N_1677,N_793,N_50);
and U1678 (N_1678,N_375,In_1482);
nand U1679 (N_1679,N_316,N_293);
and U1680 (N_1680,In_816,In_333);
nor U1681 (N_1681,In_221,In_1462);
xor U1682 (N_1682,In_1832,N_283);
and U1683 (N_1683,N_782,N_336);
and U1684 (N_1684,In_1056,In_747);
nand U1685 (N_1685,N_228,N_843);
xnor U1686 (N_1686,N_100,In_738);
nand U1687 (N_1687,N_410,In_1538);
xor U1688 (N_1688,N_27,In_122);
or U1689 (N_1689,N_706,In_1714);
and U1690 (N_1690,N_213,N_579);
and U1691 (N_1691,In_1007,In_737);
nand U1692 (N_1692,In_11,N_504);
or U1693 (N_1693,N_439,In_412);
xor U1694 (N_1694,N_150,In_1166);
nand U1695 (N_1695,In_1021,N_728);
nor U1696 (N_1696,N_586,N_898);
nor U1697 (N_1697,In_1317,N_353);
xnor U1698 (N_1698,In_775,N_796);
nor U1699 (N_1699,N_870,In_1465);
nand U1700 (N_1700,N_108,N_134);
or U1701 (N_1701,In_2340,N_506);
nor U1702 (N_1702,In_1660,In_1535);
nand U1703 (N_1703,N_219,N_550);
and U1704 (N_1704,N_8,N_549);
or U1705 (N_1705,N_511,In_1630);
nor U1706 (N_1706,N_824,In_1949);
or U1707 (N_1707,In_376,N_642);
xnor U1708 (N_1708,N_242,N_687);
and U1709 (N_1709,N_348,N_149);
or U1710 (N_1710,N_419,N_638);
nor U1711 (N_1711,N_593,N_621);
and U1712 (N_1712,N_92,In_632);
nand U1713 (N_1713,N_227,N_362);
xor U1714 (N_1714,N_269,N_206);
or U1715 (N_1715,N_371,N_926);
or U1716 (N_1716,N_211,N_267);
and U1717 (N_1717,N_626,In_922);
xnor U1718 (N_1718,N_78,N_915);
and U1719 (N_1719,N_388,N_673);
and U1720 (N_1720,In_157,N_264);
and U1721 (N_1721,N_983,N_512);
nand U1722 (N_1722,N_221,In_1742);
nor U1723 (N_1723,N_407,N_740);
nand U1724 (N_1724,In_681,N_761);
or U1725 (N_1725,In_62,N_842);
xnor U1726 (N_1726,In_1957,N_420);
nor U1727 (N_1727,N_905,In_484);
nor U1728 (N_1728,N_648,N_515);
xnor U1729 (N_1729,N_911,N_757);
nor U1730 (N_1730,N_624,N_494);
nand U1731 (N_1731,N_680,N_552);
and U1732 (N_1732,N_95,N_33);
xor U1733 (N_1733,In_466,N_759);
nor U1734 (N_1734,In_2345,In_532);
xor U1735 (N_1735,N_554,In_1369);
or U1736 (N_1736,In_1641,N_955);
nand U1737 (N_1737,In_1849,In_204);
and U1738 (N_1738,In_1699,N_476);
or U1739 (N_1739,N_103,N_49);
nor U1740 (N_1740,N_493,N_534);
or U1741 (N_1741,N_888,N_612);
nor U1742 (N_1742,N_834,In_423);
xnor U1743 (N_1743,N_93,In_127);
and U1744 (N_1744,N_207,In_1712);
or U1745 (N_1745,N_110,N_791);
nor U1746 (N_1746,N_76,N_128);
nand U1747 (N_1747,In_565,N_927);
or U1748 (N_1748,In_1052,In_1501);
or U1749 (N_1749,N_613,N_383);
nor U1750 (N_1750,N_706,N_613);
nand U1751 (N_1751,N_367,In_1142);
nor U1752 (N_1752,N_962,N_794);
or U1753 (N_1753,N_284,N_281);
nand U1754 (N_1754,N_437,N_136);
and U1755 (N_1755,N_174,N_799);
or U1756 (N_1756,N_783,N_745);
or U1757 (N_1757,N_357,N_951);
or U1758 (N_1758,N_884,In_1780);
or U1759 (N_1759,N_309,In_2005);
or U1760 (N_1760,N_164,N_171);
nand U1761 (N_1761,N_153,N_366);
nor U1762 (N_1762,In_1643,N_359);
and U1763 (N_1763,In_968,In_1056);
xnor U1764 (N_1764,N_74,N_242);
xnor U1765 (N_1765,In_1482,N_64);
nand U1766 (N_1766,N_625,N_561);
and U1767 (N_1767,In_2059,In_1539);
and U1768 (N_1768,N_526,N_959);
xnor U1769 (N_1769,N_363,N_37);
xor U1770 (N_1770,N_514,N_847);
or U1771 (N_1771,In_1351,N_270);
xor U1772 (N_1772,N_532,N_618);
nand U1773 (N_1773,N_807,In_287);
and U1774 (N_1774,In_1314,N_906);
xnor U1775 (N_1775,N_987,N_884);
and U1776 (N_1776,In_261,N_994);
xnor U1777 (N_1777,N_446,N_903);
and U1778 (N_1778,N_498,N_863);
xnor U1779 (N_1779,N_174,N_711);
or U1780 (N_1780,N_353,In_931);
xnor U1781 (N_1781,In_1601,N_167);
or U1782 (N_1782,N_376,N_971);
nand U1783 (N_1783,In_2162,N_368);
nor U1784 (N_1784,N_443,N_605);
and U1785 (N_1785,N_400,N_741);
or U1786 (N_1786,N_422,N_303);
xnor U1787 (N_1787,In_622,N_927);
nor U1788 (N_1788,N_30,N_987);
nor U1789 (N_1789,In_500,N_815);
or U1790 (N_1790,N_849,N_658);
nor U1791 (N_1791,N_131,N_840);
nand U1792 (N_1792,N_936,In_336);
xor U1793 (N_1793,N_121,In_655);
xnor U1794 (N_1794,N_914,In_2268);
and U1795 (N_1795,In_472,N_131);
xor U1796 (N_1796,In_1962,In_1680);
or U1797 (N_1797,N_234,N_401);
and U1798 (N_1798,N_220,In_587);
xor U1799 (N_1799,In_1757,In_117);
and U1800 (N_1800,N_415,N_755);
or U1801 (N_1801,In_2358,N_883);
nand U1802 (N_1802,N_144,N_967);
and U1803 (N_1803,N_242,N_240);
nand U1804 (N_1804,N_804,N_728);
xor U1805 (N_1805,N_154,N_935);
xor U1806 (N_1806,N_287,In_1052);
or U1807 (N_1807,N_845,In_1694);
nand U1808 (N_1808,N_755,N_939);
nor U1809 (N_1809,N_156,N_368);
nor U1810 (N_1810,N_982,N_877);
nand U1811 (N_1811,N_917,N_965);
and U1812 (N_1812,N_463,N_258);
nor U1813 (N_1813,In_530,N_988);
nand U1814 (N_1814,N_990,N_550);
nand U1815 (N_1815,In_1429,N_823);
nand U1816 (N_1816,N_727,N_768);
xnor U1817 (N_1817,N_301,N_120);
xnor U1818 (N_1818,N_904,N_620);
nor U1819 (N_1819,In_500,In_376);
or U1820 (N_1820,N_951,N_805);
nor U1821 (N_1821,N_756,In_736);
nand U1822 (N_1822,N_320,N_809);
nor U1823 (N_1823,N_299,N_785);
or U1824 (N_1824,In_767,N_65);
xnor U1825 (N_1825,N_339,In_2433);
nand U1826 (N_1826,In_1185,In_1707);
xor U1827 (N_1827,In_1832,N_197);
and U1828 (N_1828,N_295,In_210);
nand U1829 (N_1829,In_626,In_131);
xor U1830 (N_1830,N_496,N_159);
and U1831 (N_1831,N_47,N_286);
nand U1832 (N_1832,N_108,N_468);
nor U1833 (N_1833,N_477,N_335);
or U1834 (N_1834,N_173,N_378);
nor U1835 (N_1835,N_915,N_692);
or U1836 (N_1836,N_48,In_1641);
nand U1837 (N_1837,N_213,In_1738);
xor U1838 (N_1838,N_701,In_1711);
nor U1839 (N_1839,N_809,In_919);
nand U1840 (N_1840,N_904,N_330);
xnor U1841 (N_1841,N_142,In_3);
xnor U1842 (N_1842,In_1021,N_329);
nor U1843 (N_1843,In_1693,N_201);
xnor U1844 (N_1844,N_532,In_333);
nand U1845 (N_1845,N_914,N_960);
nand U1846 (N_1846,N_685,In_705);
xor U1847 (N_1847,N_187,N_345);
or U1848 (N_1848,In_1554,N_765);
and U1849 (N_1849,N_963,N_943);
nor U1850 (N_1850,N_812,N_467);
nor U1851 (N_1851,N_731,In_880);
xor U1852 (N_1852,N_801,N_80);
xor U1853 (N_1853,N_654,N_123);
xnor U1854 (N_1854,N_681,In_626);
nor U1855 (N_1855,N_566,In_1003);
nand U1856 (N_1856,N_583,In_2192);
xor U1857 (N_1857,N_399,N_123);
or U1858 (N_1858,N_555,In_2071);
nor U1859 (N_1859,N_46,In_1870);
nand U1860 (N_1860,In_2380,N_805);
or U1861 (N_1861,In_540,In_792);
or U1862 (N_1862,In_2492,N_246);
xor U1863 (N_1863,N_468,In_2045);
xnor U1864 (N_1864,N_10,N_73);
xnor U1865 (N_1865,N_727,N_78);
nor U1866 (N_1866,N_294,N_705);
and U1867 (N_1867,N_66,N_115);
nand U1868 (N_1868,In_157,In_665);
nand U1869 (N_1869,N_336,N_925);
xnor U1870 (N_1870,In_263,N_54);
xnor U1871 (N_1871,N_579,N_439);
nand U1872 (N_1872,N_252,N_179);
or U1873 (N_1873,N_43,N_975);
nor U1874 (N_1874,N_915,N_33);
or U1875 (N_1875,N_956,In_1259);
and U1876 (N_1876,In_2162,N_62);
nor U1877 (N_1877,In_1363,In_1870);
or U1878 (N_1878,N_122,N_680);
nor U1879 (N_1879,In_1891,N_605);
or U1880 (N_1880,In_775,In_1090);
nand U1881 (N_1881,In_1844,In_1380);
nor U1882 (N_1882,N_9,N_11);
and U1883 (N_1883,N_723,In_2492);
xnor U1884 (N_1884,N_919,In_508);
or U1885 (N_1885,N_606,In_1709);
nor U1886 (N_1886,N_524,N_936);
and U1887 (N_1887,In_1156,N_592);
nor U1888 (N_1888,N_872,N_684);
and U1889 (N_1889,In_1964,In_50);
nor U1890 (N_1890,In_978,N_163);
and U1891 (N_1891,In_2433,N_780);
or U1892 (N_1892,N_119,N_391);
and U1893 (N_1893,N_508,N_451);
xnor U1894 (N_1894,In_1757,In_1056);
and U1895 (N_1895,In_565,N_950);
or U1896 (N_1896,N_16,N_921);
and U1897 (N_1897,N_212,N_378);
xor U1898 (N_1898,In_1314,N_913);
xor U1899 (N_1899,N_895,N_222);
xor U1900 (N_1900,N_609,In_731);
and U1901 (N_1901,N_441,In_1738);
nor U1902 (N_1902,In_1210,N_239);
or U1903 (N_1903,N_979,N_379);
nand U1904 (N_1904,In_481,N_343);
xor U1905 (N_1905,In_2358,N_346);
or U1906 (N_1906,In_1329,In_1676);
nor U1907 (N_1907,In_917,N_657);
nor U1908 (N_1908,In_1406,N_478);
and U1909 (N_1909,In_922,N_403);
or U1910 (N_1910,N_554,N_320);
nor U1911 (N_1911,N_989,N_150);
and U1912 (N_1912,N_146,N_477);
nor U1913 (N_1913,N_340,N_195);
and U1914 (N_1914,N_288,N_505);
and U1915 (N_1915,N_20,In_2374);
and U1916 (N_1916,N_547,In_336);
nand U1917 (N_1917,N_29,In_380);
or U1918 (N_1918,N_488,N_416);
nor U1919 (N_1919,N_203,N_477);
nor U1920 (N_1920,In_287,In_1021);
nand U1921 (N_1921,N_914,N_679);
xor U1922 (N_1922,N_341,N_872);
nor U1923 (N_1923,N_477,N_143);
nand U1924 (N_1924,N_592,N_256);
or U1925 (N_1925,In_450,N_530);
nand U1926 (N_1926,N_678,N_824);
xor U1927 (N_1927,N_532,In_369);
and U1928 (N_1928,In_248,N_352);
nor U1929 (N_1929,In_587,In_1388);
or U1930 (N_1930,N_402,N_553);
or U1931 (N_1931,N_609,In_810);
xnor U1932 (N_1932,N_9,N_972);
nand U1933 (N_1933,N_806,N_514);
nor U1934 (N_1934,In_259,In_1308);
xnor U1935 (N_1935,In_737,N_730);
xor U1936 (N_1936,N_466,In_738);
and U1937 (N_1937,N_354,N_820);
xnor U1938 (N_1938,N_816,In_1469);
nand U1939 (N_1939,In_446,N_644);
nand U1940 (N_1940,N_84,In_1586);
and U1941 (N_1941,In_606,In_1025);
nor U1942 (N_1942,N_81,In_2312);
nor U1943 (N_1943,In_1912,N_573);
and U1944 (N_1944,In_166,N_205);
or U1945 (N_1945,In_475,N_418);
and U1946 (N_1946,N_481,N_688);
or U1947 (N_1947,N_992,N_296);
or U1948 (N_1948,In_1119,N_748);
nand U1949 (N_1949,In_1532,N_890);
nand U1950 (N_1950,N_535,In_859);
or U1951 (N_1951,N_268,In_1273);
and U1952 (N_1952,N_738,N_258);
nand U1953 (N_1953,N_725,In_1844);
nor U1954 (N_1954,In_258,N_629);
or U1955 (N_1955,In_738,N_758);
xnor U1956 (N_1956,N_747,N_644);
nor U1957 (N_1957,In_1714,N_203);
nor U1958 (N_1958,N_141,N_891);
nor U1959 (N_1959,N_582,N_136);
xor U1960 (N_1960,N_632,In_2042);
or U1961 (N_1961,In_2373,In_2224);
xnor U1962 (N_1962,In_2011,N_864);
or U1963 (N_1963,N_55,In_2473);
xor U1964 (N_1964,In_450,In_1925);
nor U1965 (N_1965,N_297,N_191);
nor U1966 (N_1966,N_37,In_1490);
and U1967 (N_1967,In_2174,N_934);
or U1968 (N_1968,N_34,N_455);
or U1969 (N_1969,In_1132,N_216);
xnor U1970 (N_1970,N_382,N_613);
and U1971 (N_1971,In_720,N_771);
or U1972 (N_1972,N_0,N_929);
nor U1973 (N_1973,N_472,N_662);
or U1974 (N_1974,N_621,In_775);
nand U1975 (N_1975,N_70,N_706);
nand U1976 (N_1976,In_703,In_76);
nor U1977 (N_1977,In_1309,N_362);
xnor U1978 (N_1978,N_970,N_59);
xor U1979 (N_1979,In_2168,N_985);
and U1980 (N_1980,In_1870,N_206);
xor U1981 (N_1981,N_708,N_174);
or U1982 (N_1982,In_1232,In_1957);
or U1983 (N_1983,N_88,N_410);
nor U1984 (N_1984,N_268,In_48);
xor U1985 (N_1985,N_120,N_678);
nor U1986 (N_1986,N_903,N_115);
nand U1987 (N_1987,N_599,N_29);
or U1988 (N_1988,In_833,N_90);
and U1989 (N_1989,In_326,In_2410);
and U1990 (N_1990,N_560,N_625);
and U1991 (N_1991,N_223,N_216);
and U1992 (N_1992,N_286,N_238);
or U1993 (N_1993,In_1369,In_1482);
nand U1994 (N_1994,N_349,N_35);
or U1995 (N_1995,N_246,In_1021);
xor U1996 (N_1996,N_383,In_354);
or U1997 (N_1997,N_700,In_2216);
nand U1998 (N_1998,In_1100,In_48);
nand U1999 (N_1999,N_338,N_976);
xor U2000 (N_2000,N_1602,N_1880);
xor U2001 (N_2001,N_1504,N_1596);
nand U2002 (N_2002,N_1384,N_1426);
xor U2003 (N_2003,N_1538,N_1148);
nand U2004 (N_2004,N_1065,N_1410);
nand U2005 (N_2005,N_1976,N_1645);
xor U2006 (N_2006,N_1516,N_1280);
nor U2007 (N_2007,N_1002,N_1531);
or U2008 (N_2008,N_1197,N_1887);
nor U2009 (N_2009,N_1147,N_1279);
and U2010 (N_2010,N_1144,N_1106);
xnor U2011 (N_2011,N_1671,N_1035);
xnor U2012 (N_2012,N_1510,N_1096);
or U2013 (N_2013,N_1665,N_1822);
or U2014 (N_2014,N_1211,N_1508);
and U2015 (N_2015,N_1001,N_1398);
and U2016 (N_2016,N_1291,N_1678);
or U2017 (N_2017,N_1313,N_1448);
and U2018 (N_2018,N_1404,N_1111);
or U2019 (N_2019,N_1618,N_1885);
nor U2020 (N_2020,N_1092,N_1394);
and U2021 (N_2021,N_1753,N_1859);
xor U2022 (N_2022,N_1617,N_1764);
xnor U2023 (N_2023,N_1662,N_1659);
nand U2024 (N_2024,N_1483,N_1988);
xnor U2025 (N_2025,N_1803,N_1331);
or U2026 (N_2026,N_1808,N_1995);
nor U2027 (N_2027,N_1315,N_1863);
nor U2028 (N_2028,N_1858,N_1079);
and U2029 (N_2029,N_1402,N_1977);
or U2030 (N_2030,N_1798,N_1725);
xnor U2031 (N_2031,N_1588,N_1867);
nand U2032 (N_2032,N_1775,N_1584);
and U2033 (N_2033,N_1129,N_1806);
or U2034 (N_2034,N_1233,N_1193);
or U2035 (N_2035,N_1467,N_1639);
and U2036 (N_2036,N_1955,N_1889);
nand U2037 (N_2037,N_1325,N_1706);
nor U2038 (N_2038,N_1541,N_1982);
and U2039 (N_2039,N_1535,N_1991);
or U2040 (N_2040,N_1968,N_1554);
xnor U2041 (N_2041,N_1260,N_1396);
or U2042 (N_2042,N_1479,N_1375);
nand U2043 (N_2043,N_1607,N_1821);
nor U2044 (N_2044,N_1388,N_1024);
and U2045 (N_2045,N_1393,N_1075);
nand U2046 (N_2046,N_1500,N_1012);
or U2047 (N_2047,N_1540,N_1062);
and U2048 (N_2048,N_1589,N_1274);
nor U2049 (N_2049,N_1297,N_1761);
nand U2050 (N_2050,N_1462,N_1542);
nand U2051 (N_2051,N_1293,N_1557);
nand U2052 (N_2052,N_1401,N_1055);
nor U2053 (N_2053,N_1149,N_1351);
xnor U2054 (N_2054,N_1027,N_1695);
and U2055 (N_2055,N_1537,N_1314);
or U2056 (N_2056,N_1304,N_1009);
and U2057 (N_2057,N_1757,N_1031);
xor U2058 (N_2058,N_1872,N_1511);
nand U2059 (N_2059,N_1369,N_1308);
nand U2060 (N_2060,N_1344,N_1568);
and U2061 (N_2061,N_1956,N_1974);
or U2062 (N_2062,N_1321,N_1323);
nand U2063 (N_2063,N_1524,N_1747);
or U2064 (N_2064,N_1654,N_1492);
and U2065 (N_2065,N_1383,N_1132);
nor U2066 (N_2066,N_1135,N_1326);
and U2067 (N_2067,N_1506,N_1916);
or U2068 (N_2068,N_1340,N_1622);
or U2069 (N_2069,N_1102,N_1305);
nor U2070 (N_2070,N_1324,N_1360);
nor U2071 (N_2071,N_1998,N_1239);
nor U2072 (N_2072,N_1629,N_1306);
or U2073 (N_2073,N_1637,N_1390);
or U2074 (N_2074,N_1153,N_1558);
nor U2075 (N_2075,N_1781,N_1407);
nand U2076 (N_2076,N_1660,N_1406);
or U2077 (N_2077,N_1041,N_1578);
and U2078 (N_2078,N_1533,N_1472);
nand U2079 (N_2079,N_1905,N_1018);
nor U2080 (N_2080,N_1139,N_1947);
or U2081 (N_2081,N_1235,N_1037);
or U2082 (N_2082,N_1507,N_1784);
or U2083 (N_2083,N_1985,N_1796);
nor U2084 (N_2084,N_1019,N_1150);
xnor U2085 (N_2085,N_1021,N_1690);
or U2086 (N_2086,N_1631,N_1854);
xnor U2087 (N_2087,N_1845,N_1620);
nor U2088 (N_2088,N_1015,N_1437);
or U2089 (N_2089,N_1846,N_1301);
or U2090 (N_2090,N_1316,N_1336);
or U2091 (N_2091,N_1105,N_1376);
and U2092 (N_2092,N_1115,N_1994);
nor U2093 (N_2093,N_1302,N_1932);
and U2094 (N_2094,N_1057,N_1054);
nor U2095 (N_2095,N_1721,N_1941);
nor U2096 (N_2096,N_1641,N_1726);
nand U2097 (N_2097,N_1493,N_1922);
nand U2098 (N_2098,N_1480,N_1957);
and U2099 (N_2099,N_1552,N_1934);
or U2100 (N_2100,N_1777,N_1627);
and U2101 (N_2101,N_1759,N_1320);
nor U2102 (N_2102,N_1429,N_1299);
nor U2103 (N_2103,N_1431,N_1458);
nand U2104 (N_2104,N_1460,N_1563);
or U2105 (N_2105,N_1415,N_1952);
nand U2106 (N_2106,N_1623,N_1186);
or U2107 (N_2107,N_1137,N_1285);
xnor U2108 (N_2108,N_1481,N_1230);
nor U2109 (N_2109,N_1244,N_1087);
and U2110 (N_2110,N_1553,N_1489);
xor U2111 (N_2111,N_1463,N_1779);
nand U2112 (N_2112,N_1261,N_1714);
nor U2113 (N_2113,N_1748,N_1095);
nand U2114 (N_2114,N_1549,N_1457);
nand U2115 (N_2115,N_1679,N_1612);
or U2116 (N_2116,N_1090,N_1848);
and U2117 (N_2117,N_1071,N_1920);
xor U2118 (N_2118,N_1194,N_1283);
xnor U2119 (N_2119,N_1760,N_1249);
nand U2120 (N_2120,N_1082,N_1337);
xor U2121 (N_2121,N_1339,N_1456);
nand U2122 (N_2122,N_1767,N_1736);
nand U2123 (N_2123,N_1074,N_1091);
xor U2124 (N_2124,N_1754,N_1616);
or U2125 (N_2125,N_1517,N_1518);
nor U2126 (N_2126,N_1635,N_1583);
nand U2127 (N_2127,N_1704,N_1007);
nand U2128 (N_2128,N_1182,N_1569);
nor U2129 (N_2129,N_1694,N_1983);
nor U2130 (N_2130,N_1048,N_1923);
nor U2131 (N_2131,N_1909,N_1547);
and U2132 (N_2132,N_1005,N_1898);
xnor U2133 (N_2133,N_1046,N_1644);
or U2134 (N_2134,N_1051,N_1405);
nor U2135 (N_2135,N_1373,N_1113);
nor U2136 (N_2136,N_1972,N_1318);
or U2137 (N_2137,N_1029,N_1902);
or U2138 (N_2138,N_1495,N_1167);
nand U2139 (N_2139,N_1927,N_1403);
and U2140 (N_2140,N_1136,N_1829);
nor U2141 (N_2141,N_1591,N_1795);
nand U2142 (N_2142,N_1750,N_1544);
or U2143 (N_2143,N_1443,N_1159);
and U2144 (N_2144,N_1935,N_1545);
and U2145 (N_2145,N_1897,N_1418);
xor U2146 (N_2146,N_1119,N_1298);
nor U2147 (N_2147,N_1990,N_1422);
and U2148 (N_2148,N_1441,N_1669);
xor U2149 (N_2149,N_1514,N_1461);
nand U2150 (N_2150,N_1815,N_1901);
xnor U2151 (N_2151,N_1276,N_1411);
and U2152 (N_2152,N_1951,N_1653);
and U2153 (N_2153,N_1765,N_1603);
nor U2154 (N_2154,N_1469,N_1294);
and U2155 (N_2155,N_1424,N_1890);
nand U2156 (N_2156,N_1329,N_1427);
xor U2157 (N_2157,N_1894,N_1685);
nor U2158 (N_2158,N_1487,N_1392);
xor U2159 (N_2159,N_1361,N_1494);
or U2160 (N_2160,N_1442,N_1131);
nor U2161 (N_2161,N_1000,N_1278);
nand U2162 (N_2162,N_1053,N_1190);
nand U2163 (N_2163,N_1900,N_1787);
nand U2164 (N_2164,N_1817,N_1502);
or U2165 (N_2165,N_1327,N_1770);
xor U2166 (N_2166,N_1272,N_1634);
and U2167 (N_2167,N_1248,N_1959);
and U2168 (N_2168,N_1640,N_1925);
and U2169 (N_2169,N_1751,N_1794);
nor U2170 (N_2170,N_1921,N_1610);
or U2171 (N_2171,N_1058,N_1226);
and U2172 (N_2172,N_1838,N_1961);
nor U2173 (N_2173,N_1946,N_1070);
and U2174 (N_2174,N_1512,N_1275);
or U2175 (N_2175,N_1891,N_1824);
nand U2176 (N_2176,N_1245,N_1643);
nand U2177 (N_2177,N_1341,N_1939);
or U2178 (N_2178,N_1421,N_1056);
or U2179 (N_2179,N_1723,N_1258);
nand U2180 (N_2180,N_1451,N_1828);
nand U2181 (N_2181,N_1300,N_1399);
xnor U2182 (N_2182,N_1371,N_1040);
or U2183 (N_2183,N_1937,N_1948);
or U2184 (N_2184,N_1270,N_1256);
and U2185 (N_2185,N_1162,N_1104);
nand U2186 (N_2186,N_1997,N_1744);
nor U2187 (N_2187,N_1417,N_1598);
nand U2188 (N_2188,N_1866,N_1606);
xnor U2189 (N_2189,N_1818,N_1906);
nand U2190 (N_2190,N_1212,N_1713);
nor U2191 (N_2191,N_1912,N_1797);
nand U2192 (N_2192,N_1061,N_1509);
nor U2193 (N_2193,N_1594,N_1154);
or U2194 (N_2194,N_1960,N_1400);
nand U2195 (N_2195,N_1525,N_1677);
nor U2196 (N_2196,N_1930,N_1161);
nand U2197 (N_2197,N_1731,N_1222);
nor U2198 (N_2198,N_1391,N_1560);
and U2199 (N_2199,N_1919,N_1852);
and U2200 (N_2200,N_1221,N_1895);
nand U2201 (N_2201,N_1830,N_1447);
or U2202 (N_2202,N_1661,N_1003);
or U2203 (N_2203,N_1878,N_1564);
and U2204 (N_2204,N_1730,N_1166);
nand U2205 (N_2205,N_1819,N_1561);
or U2206 (N_2206,N_1409,N_1605);
or U2207 (N_2207,N_1163,N_1993);
or U2208 (N_2208,N_1452,N_1883);
or U2209 (N_2209,N_1851,N_1084);
and U2210 (N_2210,N_1380,N_1364);
and U2211 (N_2211,N_1236,N_1551);
nand U2212 (N_2212,N_1292,N_1374);
nand U2213 (N_2213,N_1028,N_1936);
xor U2214 (N_2214,N_1680,N_1042);
or U2215 (N_2215,N_1101,N_1387);
and U2216 (N_2216,N_1146,N_1367);
and U2217 (N_2217,N_1804,N_1672);
nand U2218 (N_2218,N_1739,N_1876);
and U2219 (N_2219,N_1773,N_1098);
nor U2220 (N_2220,N_1227,N_1756);
nor U2221 (N_2221,N_1624,N_1832);
or U2222 (N_2222,N_1984,N_1853);
and U2223 (N_2223,N_1045,N_1567);
or U2224 (N_2224,N_1008,N_1171);
xor U2225 (N_2225,N_1379,N_1783);
nand U2226 (N_2226,N_1468,N_1099);
xor U2227 (N_2227,N_1185,N_1017);
nor U2228 (N_2228,N_1626,N_1097);
or U2229 (N_2229,N_1791,N_1121);
nor U2230 (N_2230,N_1143,N_1666);
nand U2231 (N_2231,N_1196,N_1928);
xor U2232 (N_2232,N_1204,N_1250);
xor U2233 (N_2233,N_1440,N_1733);
nand U2234 (N_2234,N_1559,N_1856);
or U2235 (N_2235,N_1523,N_1078);
nand U2236 (N_2236,N_1953,N_1216);
or U2237 (N_2237,N_1215,N_1032);
xor U2238 (N_2238,N_1884,N_1122);
nor U2239 (N_2239,N_1837,N_1816);
or U2240 (N_2240,N_1217,N_1214);
or U2241 (N_2241,N_1039,N_1944);
nand U2242 (N_2242,N_1899,N_1788);
nor U2243 (N_2243,N_1195,N_1157);
xor U2244 (N_2244,N_1004,N_1491);
or U2245 (N_2245,N_1580,N_1484);
and U2246 (N_2246,N_1420,N_1419);
nor U2247 (N_2247,N_1439,N_1334);
and U2248 (N_2248,N_1833,N_1289);
nor U2249 (N_2249,N_1727,N_1698);
nor U2250 (N_2250,N_1152,N_1962);
xor U2251 (N_2251,N_1158,N_1273);
nand U2252 (N_2252,N_1813,N_1823);
nand U2253 (N_2253,N_1613,N_1430);
or U2254 (N_2254,N_1772,N_1486);
nand U2255 (N_2255,N_1573,N_1353);
nor U2256 (N_2256,N_1218,N_1942);
or U2257 (N_2257,N_1188,N_1971);
nor U2258 (N_2258,N_1413,N_1436);
xor U2259 (N_2259,N_1582,N_1220);
and U2260 (N_2260,N_1908,N_1776);
nor U2261 (N_2261,N_1342,N_1475);
and U2262 (N_2262,N_1565,N_1160);
or U2263 (N_2263,N_1911,N_1574);
nand U2264 (N_2264,N_1740,N_1742);
xnor U2265 (N_2265,N_1670,N_1842);
or U2266 (N_2266,N_1886,N_1156);
xnor U2267 (N_2267,N_1903,N_1368);
and U2268 (N_2268,N_1904,N_1649);
xor U2269 (N_2269,N_1711,N_1766);
nor U2270 (N_2270,N_1438,N_1827);
or U2271 (N_2271,N_1362,N_1673);
nand U2272 (N_2272,N_1478,N_1938);
xnor U2273 (N_2273,N_1126,N_1423);
nor U2274 (N_2274,N_1253,N_1072);
and U2275 (N_2275,N_1724,N_1917);
xor U2276 (N_2276,N_1433,N_1338);
xnor U2277 (N_2277,N_1141,N_1333);
or U2278 (N_2278,N_1628,N_1309);
xor U2279 (N_2279,N_1026,N_1599);
xor U2280 (N_2280,N_1970,N_1052);
or U2281 (N_2281,N_1348,N_1496);
and U2282 (N_2282,N_1782,N_1043);
xnor U2283 (N_2283,N_1940,N_1625);
nand U2284 (N_2284,N_1130,N_1522);
nand U2285 (N_2285,N_1109,N_1702);
nor U2286 (N_2286,N_1701,N_1246);
xnor U2287 (N_2287,N_1805,N_1534);
nand U2288 (N_2288,N_1208,N_1023);
or U2289 (N_2289,N_1521,N_1519);
nor U2290 (N_2290,N_1288,N_1192);
or U2291 (N_2291,N_1020,N_1682);
or U2292 (N_2292,N_1083,N_1597);
and U2293 (N_2293,N_1785,N_1254);
and U2294 (N_2294,N_1973,N_1155);
nand U2295 (N_2295,N_1989,N_1501);
and U2296 (N_2296,N_1255,N_1172);
nor U2297 (N_2297,N_1202,N_1763);
or U2298 (N_2298,N_1322,N_1556);
nor U2299 (N_2299,N_1175,N_1191);
nor U2300 (N_2300,N_1893,N_1992);
and U2301 (N_2301,N_1950,N_1151);
and U2302 (N_2302,N_1145,N_1869);
nand U2303 (N_2303,N_1650,N_1737);
nor U2304 (N_2304,N_1600,N_1619);
nor U2305 (N_2305,N_1550,N_1967);
nand U2306 (N_2306,N_1435,N_1926);
and U2307 (N_2307,N_1868,N_1059);
nor U2308 (N_2308,N_1862,N_1127);
xnor U2309 (N_2309,N_1474,N_1710);
nand U2310 (N_2310,N_1428,N_1389);
xor U2311 (N_2311,N_1980,N_1864);
nand U2312 (N_2312,N_1257,N_1814);
and U2313 (N_2313,N_1238,N_1080);
nor U2314 (N_2314,N_1527,N_1482);
nor U2315 (N_2315,N_1466,N_1014);
nor U2316 (N_2316,N_1692,N_1780);
nor U2317 (N_2317,N_1476,N_1664);
nand U2318 (N_2318,N_1453,N_1709);
xor U2319 (N_2319,N_1271,N_1943);
nand U2320 (N_2320,N_1125,N_1356);
nand U2321 (N_2321,N_1570,N_1366);
xnor U2322 (N_2322,N_1687,N_1703);
nand U2323 (N_2323,N_1432,N_1609);
nand U2324 (N_2324,N_1181,N_1312);
and U2325 (N_2325,N_1357,N_1729);
nor U2326 (N_2326,N_1498,N_1614);
nor U2327 (N_2327,N_1601,N_1232);
nor U2328 (N_2328,N_1543,N_1810);
xor U2329 (N_2329,N_1807,N_1945);
or U2330 (N_2330,N_1178,N_1663);
nor U2331 (N_2331,N_1134,N_1718);
nor U2332 (N_2332,N_1686,N_1958);
xnor U2333 (N_2333,N_1888,N_1963);
or U2334 (N_2334,N_1789,N_1310);
or U2335 (N_2335,N_1343,N_1259);
nand U2336 (N_2336,N_1656,N_1874);
or U2337 (N_2337,N_1077,N_1228);
and U2338 (N_2338,N_1473,N_1128);
nor U2339 (N_2339,N_1385,N_1231);
and U2340 (N_2340,N_1268,N_1116);
xor U2341 (N_2341,N_1987,N_1611);
and U2342 (N_2342,N_1571,N_1877);
or U2343 (N_2343,N_1450,N_1831);
xor U2344 (N_2344,N_1657,N_1728);
and U2345 (N_2345,N_1286,N_1319);
nand U2346 (N_2346,N_1749,N_1219);
nand U2347 (N_2347,N_1290,N_1719);
nand U2348 (N_2348,N_1395,N_1240);
nor U2349 (N_2349,N_1790,N_1386);
or U2350 (N_2350,N_1022,N_1464);
nand U2351 (N_2351,N_1370,N_1434);
and U2352 (N_2352,N_1068,N_1536);
nor U2353 (N_2353,N_1277,N_1873);
or U2354 (N_2354,N_1840,N_1755);
nor U2355 (N_2355,N_1016,N_1425);
nor U2356 (N_2356,N_1683,N_1865);
or U2357 (N_2357,N_1229,N_1455);
and U2358 (N_2358,N_1834,N_1741);
nor U2359 (N_2359,N_1849,N_1615);
or U2360 (N_2360,N_1459,N_1913);
or U2361 (N_2361,N_1529,N_1505);
and U2362 (N_2362,N_1575,N_1247);
nand U2363 (N_2363,N_1604,N_1281);
or U2364 (N_2364,N_1855,N_1546);
nor U2365 (N_2365,N_1732,N_1363);
and U2366 (N_2366,N_1203,N_1608);
nor U2367 (N_2367,N_1110,N_1882);
or U2368 (N_2368,N_1734,N_1520);
and U2369 (N_2369,N_1799,N_1592);
nor U2370 (N_2370,N_1595,N_1949);
nor U2371 (N_2371,N_1267,N_1843);
nand U2372 (N_2372,N_1223,N_1875);
nand U2373 (N_2373,N_1802,N_1445);
and U2374 (N_2374,N_1497,N_1847);
or U2375 (N_2375,N_1896,N_1047);
and U2376 (N_2376,N_1700,N_1081);
nand U2377 (N_2377,N_1655,N_1586);
nor U2378 (N_2378,N_1209,N_1577);
xnor U2379 (N_2379,N_1225,N_1964);
and U2380 (N_2380,N_1006,N_1213);
or U2381 (N_2381,N_1881,N_1720);
nand U2382 (N_2382,N_1572,N_1381);
and U2383 (N_2383,N_1237,N_1735);
and U2384 (N_2384,N_1470,N_1555);
nor U2385 (N_2385,N_1978,N_1176);
nor U2386 (N_2386,N_1969,N_1689);
nor U2387 (N_2387,N_1712,N_1630);
and U2388 (N_2388,N_1296,N_1397);
or U2389 (N_2389,N_1786,N_1762);
nor U2390 (N_2390,N_1528,N_1243);
nand U2391 (N_2391,N_1579,N_1076);
nor U2392 (N_2392,N_1861,N_1086);
xor U2393 (N_2393,N_1752,N_1030);
nand U2394 (N_2394,N_1117,N_1485);
or U2395 (N_2395,N_1165,N_1490);
and U2396 (N_2396,N_1372,N_1722);
or U2397 (N_2397,N_1716,N_1044);
xor U2398 (N_2398,N_1382,N_1870);
nand U2399 (N_2399,N_1841,N_1581);
nor U2400 (N_2400,N_1089,N_1515);
and U2401 (N_2401,N_1668,N_1647);
nor U2402 (N_2402,N_1063,N_1771);
nand U2403 (N_2403,N_1860,N_1871);
or U2404 (N_2404,N_1996,N_1346);
nor U2405 (N_2405,N_1252,N_1187);
nand U2406 (N_2406,N_1778,N_1262);
and U2407 (N_2407,N_1060,N_1264);
and U2408 (N_2408,N_1064,N_1133);
and U2409 (N_2409,N_1120,N_1835);
nand U2410 (N_2410,N_1915,N_1705);
or U2411 (N_2411,N_1743,N_1295);
or U2412 (N_2412,N_1688,N_1566);
nor U2413 (N_2413,N_1929,N_1981);
nor U2414 (N_2414,N_1774,N_1532);
or U2415 (N_2415,N_1038,N_1801);
or U2416 (N_2416,N_1715,N_1931);
xor U2417 (N_2417,N_1446,N_1242);
nor U2418 (N_2418,N_1812,N_1234);
nor U2419 (N_2419,N_1954,N_1352);
xor U2420 (N_2420,N_1738,N_1085);
nand U2421 (N_2421,N_1358,N_1093);
and U2422 (N_2422,N_1684,N_1966);
xor U2423 (N_2423,N_1266,N_1562);
nor U2424 (N_2424,N_1693,N_1768);
or U2425 (N_2425,N_1050,N_1349);
and U2426 (N_2426,N_1345,N_1590);
nor U2427 (N_2427,N_1124,N_1658);
or U2428 (N_2428,N_1174,N_1844);
xnor U2429 (N_2429,N_1180,N_1793);
and U2430 (N_2430,N_1034,N_1576);
xnor U2431 (N_2431,N_1114,N_1699);
or U2432 (N_2432,N_1696,N_1667);
nand U2433 (N_2433,N_1924,N_1697);
nor U2434 (N_2434,N_1013,N_1593);
nor U2435 (N_2435,N_1317,N_1033);
nor U2436 (N_2436,N_1335,N_1621);
nand U2437 (N_2437,N_1168,N_1287);
xor U2438 (N_2438,N_1269,N_1408);
and U2439 (N_2439,N_1642,N_1914);
xor U2440 (N_2440,N_1173,N_1675);
and U2441 (N_2441,N_1284,N_1108);
nor U2442 (N_2442,N_1359,N_1025);
nand U2443 (N_2443,N_1758,N_1347);
nor U2444 (N_2444,N_1539,N_1189);
or U2445 (N_2445,N_1811,N_1010);
xor U2446 (N_2446,N_1036,N_1454);
or U2447 (N_2447,N_1307,N_1850);
or U2448 (N_2448,N_1330,N_1488);
nor U2449 (N_2449,N_1975,N_1303);
nand U2450 (N_2450,N_1587,N_1179);
or U2451 (N_2451,N_1892,N_1999);
or U2452 (N_2452,N_1839,N_1365);
xnor U2453 (N_2453,N_1530,N_1328);
nor U2454 (N_2454,N_1412,N_1350);
nand U2455 (N_2455,N_1826,N_1513);
nand U2456 (N_2456,N_1332,N_1107);
nand U2457 (N_2457,N_1674,N_1088);
and U2458 (N_2458,N_1651,N_1465);
and U2459 (N_2459,N_1707,N_1499);
nand U2460 (N_2460,N_1676,N_1708);
or U2461 (N_2461,N_1164,N_1548);
nand U2462 (N_2462,N_1449,N_1251);
nor U2463 (N_2463,N_1652,N_1918);
nand U2464 (N_2464,N_1184,N_1681);
xnor U2465 (N_2465,N_1224,N_1857);
nand U2466 (N_2466,N_1444,N_1311);
and U2467 (N_2467,N_1067,N_1414);
or U2468 (N_2468,N_1636,N_1103);
or U2469 (N_2469,N_1207,N_1879);
or U2470 (N_2470,N_1112,N_1073);
xor U2471 (N_2471,N_1416,N_1825);
or U2472 (N_2472,N_1138,N_1206);
and U2473 (N_2473,N_1646,N_1069);
nand U2474 (N_2474,N_1378,N_1263);
xnor U2475 (N_2475,N_1282,N_1965);
xnor U2476 (N_2476,N_1066,N_1377);
and U2477 (N_2477,N_1907,N_1201);
nor U2478 (N_2478,N_1769,N_1355);
nand U2479 (N_2479,N_1100,N_1265);
nor U2480 (N_2480,N_1836,N_1638);
nor U2481 (N_2481,N_1910,N_1933);
or U2482 (N_2482,N_1169,N_1986);
or U2483 (N_2483,N_1199,N_1049);
nand U2484 (N_2484,N_1094,N_1717);
or U2485 (N_2485,N_1979,N_1170);
xor U2486 (N_2486,N_1800,N_1633);
xor U2487 (N_2487,N_1746,N_1792);
and U2488 (N_2488,N_1820,N_1177);
and U2489 (N_2489,N_1477,N_1205);
nor U2490 (N_2490,N_1210,N_1123);
nand U2491 (N_2491,N_1503,N_1241);
or U2492 (N_2492,N_1198,N_1526);
nand U2493 (N_2493,N_1809,N_1745);
or U2494 (N_2494,N_1691,N_1118);
or U2495 (N_2495,N_1142,N_1648);
and U2496 (N_2496,N_1471,N_1585);
and U2497 (N_2497,N_1140,N_1183);
nor U2498 (N_2498,N_1354,N_1011);
or U2499 (N_2499,N_1200,N_1632);
or U2500 (N_2500,N_1654,N_1313);
nand U2501 (N_2501,N_1066,N_1524);
xor U2502 (N_2502,N_1482,N_1123);
nand U2503 (N_2503,N_1120,N_1813);
nor U2504 (N_2504,N_1591,N_1229);
nor U2505 (N_2505,N_1187,N_1650);
nor U2506 (N_2506,N_1479,N_1666);
and U2507 (N_2507,N_1409,N_1629);
nor U2508 (N_2508,N_1561,N_1173);
nor U2509 (N_2509,N_1591,N_1628);
and U2510 (N_2510,N_1382,N_1420);
and U2511 (N_2511,N_1147,N_1671);
and U2512 (N_2512,N_1655,N_1043);
nor U2513 (N_2513,N_1945,N_1726);
or U2514 (N_2514,N_1687,N_1255);
nor U2515 (N_2515,N_1932,N_1004);
xor U2516 (N_2516,N_1987,N_1457);
nand U2517 (N_2517,N_1141,N_1652);
xnor U2518 (N_2518,N_1236,N_1643);
or U2519 (N_2519,N_1741,N_1253);
or U2520 (N_2520,N_1874,N_1679);
and U2521 (N_2521,N_1923,N_1958);
nand U2522 (N_2522,N_1000,N_1990);
nor U2523 (N_2523,N_1618,N_1723);
and U2524 (N_2524,N_1968,N_1427);
nor U2525 (N_2525,N_1691,N_1143);
and U2526 (N_2526,N_1669,N_1568);
or U2527 (N_2527,N_1398,N_1767);
or U2528 (N_2528,N_1339,N_1669);
nand U2529 (N_2529,N_1714,N_1505);
nor U2530 (N_2530,N_1436,N_1440);
nand U2531 (N_2531,N_1688,N_1428);
or U2532 (N_2532,N_1775,N_1334);
or U2533 (N_2533,N_1950,N_1552);
nand U2534 (N_2534,N_1454,N_1489);
nor U2535 (N_2535,N_1133,N_1375);
and U2536 (N_2536,N_1652,N_1823);
xnor U2537 (N_2537,N_1190,N_1986);
nor U2538 (N_2538,N_1399,N_1648);
nand U2539 (N_2539,N_1237,N_1729);
or U2540 (N_2540,N_1023,N_1570);
xor U2541 (N_2541,N_1148,N_1699);
nor U2542 (N_2542,N_1609,N_1718);
and U2543 (N_2543,N_1772,N_1078);
or U2544 (N_2544,N_1347,N_1029);
or U2545 (N_2545,N_1896,N_1315);
xor U2546 (N_2546,N_1022,N_1333);
and U2547 (N_2547,N_1451,N_1670);
and U2548 (N_2548,N_1013,N_1112);
xnor U2549 (N_2549,N_1001,N_1653);
xor U2550 (N_2550,N_1325,N_1825);
xor U2551 (N_2551,N_1615,N_1446);
and U2552 (N_2552,N_1731,N_1419);
xor U2553 (N_2553,N_1334,N_1403);
and U2554 (N_2554,N_1821,N_1257);
nand U2555 (N_2555,N_1021,N_1495);
xor U2556 (N_2556,N_1608,N_1505);
xor U2557 (N_2557,N_1588,N_1678);
nor U2558 (N_2558,N_1273,N_1015);
or U2559 (N_2559,N_1056,N_1212);
or U2560 (N_2560,N_1913,N_1620);
xnor U2561 (N_2561,N_1854,N_1081);
or U2562 (N_2562,N_1893,N_1875);
nor U2563 (N_2563,N_1862,N_1794);
and U2564 (N_2564,N_1903,N_1848);
nor U2565 (N_2565,N_1717,N_1012);
nor U2566 (N_2566,N_1024,N_1869);
nor U2567 (N_2567,N_1369,N_1484);
xnor U2568 (N_2568,N_1491,N_1656);
nor U2569 (N_2569,N_1140,N_1974);
or U2570 (N_2570,N_1440,N_1256);
xor U2571 (N_2571,N_1603,N_1746);
or U2572 (N_2572,N_1914,N_1945);
and U2573 (N_2573,N_1995,N_1828);
nor U2574 (N_2574,N_1565,N_1094);
and U2575 (N_2575,N_1721,N_1607);
nand U2576 (N_2576,N_1626,N_1954);
xor U2577 (N_2577,N_1429,N_1857);
xor U2578 (N_2578,N_1753,N_1023);
and U2579 (N_2579,N_1189,N_1783);
and U2580 (N_2580,N_1215,N_1305);
nor U2581 (N_2581,N_1489,N_1755);
or U2582 (N_2582,N_1008,N_1523);
or U2583 (N_2583,N_1479,N_1247);
or U2584 (N_2584,N_1391,N_1104);
xor U2585 (N_2585,N_1904,N_1339);
or U2586 (N_2586,N_1114,N_1112);
and U2587 (N_2587,N_1477,N_1152);
xnor U2588 (N_2588,N_1122,N_1803);
xnor U2589 (N_2589,N_1950,N_1714);
and U2590 (N_2590,N_1708,N_1834);
nor U2591 (N_2591,N_1767,N_1689);
or U2592 (N_2592,N_1419,N_1340);
nand U2593 (N_2593,N_1544,N_1756);
xor U2594 (N_2594,N_1155,N_1950);
nor U2595 (N_2595,N_1649,N_1451);
or U2596 (N_2596,N_1644,N_1700);
nand U2597 (N_2597,N_1393,N_1823);
or U2598 (N_2598,N_1365,N_1913);
nand U2599 (N_2599,N_1120,N_1628);
xor U2600 (N_2600,N_1811,N_1222);
xnor U2601 (N_2601,N_1229,N_1458);
nor U2602 (N_2602,N_1031,N_1485);
and U2603 (N_2603,N_1248,N_1810);
and U2604 (N_2604,N_1124,N_1056);
nor U2605 (N_2605,N_1677,N_1449);
nor U2606 (N_2606,N_1813,N_1418);
xor U2607 (N_2607,N_1724,N_1199);
or U2608 (N_2608,N_1497,N_1328);
or U2609 (N_2609,N_1939,N_1667);
and U2610 (N_2610,N_1999,N_1130);
and U2611 (N_2611,N_1843,N_1948);
or U2612 (N_2612,N_1685,N_1152);
nor U2613 (N_2613,N_1037,N_1717);
or U2614 (N_2614,N_1464,N_1661);
xnor U2615 (N_2615,N_1743,N_1814);
and U2616 (N_2616,N_1133,N_1541);
xor U2617 (N_2617,N_1958,N_1865);
xnor U2618 (N_2618,N_1258,N_1515);
nor U2619 (N_2619,N_1341,N_1684);
and U2620 (N_2620,N_1544,N_1643);
and U2621 (N_2621,N_1032,N_1549);
and U2622 (N_2622,N_1597,N_1315);
nand U2623 (N_2623,N_1636,N_1431);
nand U2624 (N_2624,N_1223,N_1848);
or U2625 (N_2625,N_1815,N_1354);
xnor U2626 (N_2626,N_1732,N_1687);
nand U2627 (N_2627,N_1870,N_1903);
nor U2628 (N_2628,N_1581,N_1814);
nor U2629 (N_2629,N_1601,N_1043);
xor U2630 (N_2630,N_1448,N_1022);
xnor U2631 (N_2631,N_1418,N_1367);
nor U2632 (N_2632,N_1882,N_1629);
xnor U2633 (N_2633,N_1740,N_1371);
or U2634 (N_2634,N_1102,N_1429);
or U2635 (N_2635,N_1944,N_1446);
or U2636 (N_2636,N_1430,N_1340);
xor U2637 (N_2637,N_1468,N_1601);
xnor U2638 (N_2638,N_1053,N_1188);
or U2639 (N_2639,N_1986,N_1284);
nor U2640 (N_2640,N_1614,N_1779);
xnor U2641 (N_2641,N_1151,N_1411);
xnor U2642 (N_2642,N_1852,N_1897);
or U2643 (N_2643,N_1442,N_1454);
and U2644 (N_2644,N_1355,N_1738);
xnor U2645 (N_2645,N_1074,N_1446);
xnor U2646 (N_2646,N_1800,N_1328);
and U2647 (N_2647,N_1594,N_1762);
nand U2648 (N_2648,N_1519,N_1568);
and U2649 (N_2649,N_1796,N_1354);
xnor U2650 (N_2650,N_1608,N_1171);
nand U2651 (N_2651,N_1027,N_1351);
and U2652 (N_2652,N_1753,N_1739);
or U2653 (N_2653,N_1337,N_1384);
nor U2654 (N_2654,N_1236,N_1099);
nand U2655 (N_2655,N_1865,N_1675);
nand U2656 (N_2656,N_1817,N_1765);
nor U2657 (N_2657,N_1066,N_1492);
nand U2658 (N_2658,N_1963,N_1730);
or U2659 (N_2659,N_1776,N_1816);
nand U2660 (N_2660,N_1728,N_1549);
nor U2661 (N_2661,N_1814,N_1061);
nor U2662 (N_2662,N_1633,N_1054);
xor U2663 (N_2663,N_1952,N_1912);
nor U2664 (N_2664,N_1726,N_1432);
and U2665 (N_2665,N_1938,N_1403);
or U2666 (N_2666,N_1107,N_1621);
nor U2667 (N_2667,N_1343,N_1229);
and U2668 (N_2668,N_1582,N_1084);
nand U2669 (N_2669,N_1630,N_1467);
nand U2670 (N_2670,N_1100,N_1606);
nor U2671 (N_2671,N_1398,N_1075);
nor U2672 (N_2672,N_1536,N_1264);
and U2673 (N_2673,N_1464,N_1657);
and U2674 (N_2674,N_1736,N_1061);
and U2675 (N_2675,N_1710,N_1583);
and U2676 (N_2676,N_1483,N_1345);
or U2677 (N_2677,N_1477,N_1530);
nor U2678 (N_2678,N_1007,N_1881);
and U2679 (N_2679,N_1911,N_1303);
xnor U2680 (N_2680,N_1677,N_1057);
xor U2681 (N_2681,N_1007,N_1321);
nand U2682 (N_2682,N_1094,N_1327);
or U2683 (N_2683,N_1542,N_1518);
nor U2684 (N_2684,N_1502,N_1304);
nand U2685 (N_2685,N_1566,N_1400);
and U2686 (N_2686,N_1055,N_1526);
nor U2687 (N_2687,N_1791,N_1665);
or U2688 (N_2688,N_1503,N_1139);
nor U2689 (N_2689,N_1893,N_1884);
xnor U2690 (N_2690,N_1005,N_1446);
nor U2691 (N_2691,N_1205,N_1286);
xor U2692 (N_2692,N_1718,N_1699);
nand U2693 (N_2693,N_1358,N_1001);
nor U2694 (N_2694,N_1587,N_1318);
and U2695 (N_2695,N_1618,N_1958);
xnor U2696 (N_2696,N_1526,N_1223);
nand U2697 (N_2697,N_1973,N_1587);
xnor U2698 (N_2698,N_1999,N_1807);
nor U2699 (N_2699,N_1192,N_1713);
nor U2700 (N_2700,N_1469,N_1215);
or U2701 (N_2701,N_1940,N_1399);
or U2702 (N_2702,N_1458,N_1808);
nand U2703 (N_2703,N_1290,N_1275);
or U2704 (N_2704,N_1013,N_1426);
nand U2705 (N_2705,N_1988,N_1653);
nand U2706 (N_2706,N_1927,N_1773);
xnor U2707 (N_2707,N_1420,N_1403);
and U2708 (N_2708,N_1045,N_1617);
nand U2709 (N_2709,N_1150,N_1932);
nand U2710 (N_2710,N_1522,N_1507);
or U2711 (N_2711,N_1387,N_1494);
xor U2712 (N_2712,N_1990,N_1025);
nand U2713 (N_2713,N_1937,N_1790);
and U2714 (N_2714,N_1196,N_1881);
or U2715 (N_2715,N_1257,N_1483);
nand U2716 (N_2716,N_1394,N_1669);
nor U2717 (N_2717,N_1555,N_1030);
nor U2718 (N_2718,N_1887,N_1759);
and U2719 (N_2719,N_1692,N_1701);
and U2720 (N_2720,N_1709,N_1569);
nand U2721 (N_2721,N_1432,N_1931);
xor U2722 (N_2722,N_1946,N_1573);
and U2723 (N_2723,N_1422,N_1959);
nor U2724 (N_2724,N_1964,N_1858);
nor U2725 (N_2725,N_1865,N_1476);
and U2726 (N_2726,N_1929,N_1582);
xnor U2727 (N_2727,N_1768,N_1338);
or U2728 (N_2728,N_1229,N_1698);
or U2729 (N_2729,N_1904,N_1496);
or U2730 (N_2730,N_1295,N_1574);
or U2731 (N_2731,N_1253,N_1162);
and U2732 (N_2732,N_1292,N_1637);
or U2733 (N_2733,N_1383,N_1575);
and U2734 (N_2734,N_1074,N_1639);
or U2735 (N_2735,N_1562,N_1620);
or U2736 (N_2736,N_1186,N_1465);
and U2737 (N_2737,N_1290,N_1276);
and U2738 (N_2738,N_1885,N_1765);
xor U2739 (N_2739,N_1405,N_1572);
nor U2740 (N_2740,N_1246,N_1556);
nor U2741 (N_2741,N_1314,N_1831);
and U2742 (N_2742,N_1287,N_1189);
and U2743 (N_2743,N_1374,N_1388);
nand U2744 (N_2744,N_1839,N_1076);
nand U2745 (N_2745,N_1791,N_1138);
nand U2746 (N_2746,N_1460,N_1497);
and U2747 (N_2747,N_1874,N_1348);
xor U2748 (N_2748,N_1314,N_1765);
nor U2749 (N_2749,N_1373,N_1743);
xnor U2750 (N_2750,N_1771,N_1193);
xor U2751 (N_2751,N_1574,N_1388);
and U2752 (N_2752,N_1911,N_1561);
nand U2753 (N_2753,N_1091,N_1710);
nand U2754 (N_2754,N_1146,N_1788);
xor U2755 (N_2755,N_1429,N_1927);
or U2756 (N_2756,N_1820,N_1860);
nor U2757 (N_2757,N_1089,N_1343);
xnor U2758 (N_2758,N_1742,N_1305);
or U2759 (N_2759,N_1034,N_1314);
xnor U2760 (N_2760,N_1118,N_1715);
and U2761 (N_2761,N_1021,N_1906);
nand U2762 (N_2762,N_1709,N_1146);
nand U2763 (N_2763,N_1236,N_1433);
or U2764 (N_2764,N_1694,N_1636);
nand U2765 (N_2765,N_1394,N_1854);
or U2766 (N_2766,N_1527,N_1767);
nand U2767 (N_2767,N_1710,N_1842);
nor U2768 (N_2768,N_1168,N_1905);
nand U2769 (N_2769,N_1725,N_1175);
xor U2770 (N_2770,N_1634,N_1957);
nand U2771 (N_2771,N_1874,N_1962);
or U2772 (N_2772,N_1170,N_1866);
xnor U2773 (N_2773,N_1000,N_1355);
xor U2774 (N_2774,N_1336,N_1303);
and U2775 (N_2775,N_1783,N_1827);
nand U2776 (N_2776,N_1636,N_1010);
xor U2777 (N_2777,N_1854,N_1023);
nand U2778 (N_2778,N_1049,N_1197);
nor U2779 (N_2779,N_1100,N_1990);
and U2780 (N_2780,N_1353,N_1359);
and U2781 (N_2781,N_1840,N_1611);
nor U2782 (N_2782,N_1365,N_1476);
or U2783 (N_2783,N_1754,N_1530);
and U2784 (N_2784,N_1490,N_1188);
nor U2785 (N_2785,N_1775,N_1055);
or U2786 (N_2786,N_1505,N_1917);
nand U2787 (N_2787,N_1055,N_1114);
or U2788 (N_2788,N_1931,N_1503);
xor U2789 (N_2789,N_1869,N_1581);
nor U2790 (N_2790,N_1952,N_1598);
xnor U2791 (N_2791,N_1731,N_1570);
and U2792 (N_2792,N_1047,N_1364);
nand U2793 (N_2793,N_1605,N_1234);
or U2794 (N_2794,N_1590,N_1115);
xor U2795 (N_2795,N_1545,N_1567);
xor U2796 (N_2796,N_1266,N_1901);
nand U2797 (N_2797,N_1207,N_1283);
xor U2798 (N_2798,N_1864,N_1804);
nor U2799 (N_2799,N_1171,N_1970);
nor U2800 (N_2800,N_1064,N_1822);
xnor U2801 (N_2801,N_1795,N_1168);
xor U2802 (N_2802,N_1895,N_1746);
or U2803 (N_2803,N_1399,N_1995);
nor U2804 (N_2804,N_1635,N_1370);
or U2805 (N_2805,N_1277,N_1946);
xnor U2806 (N_2806,N_1759,N_1956);
nor U2807 (N_2807,N_1724,N_1310);
and U2808 (N_2808,N_1010,N_1679);
nand U2809 (N_2809,N_1554,N_1152);
nand U2810 (N_2810,N_1462,N_1008);
xnor U2811 (N_2811,N_1421,N_1686);
xor U2812 (N_2812,N_1377,N_1535);
and U2813 (N_2813,N_1927,N_1581);
nor U2814 (N_2814,N_1550,N_1411);
xor U2815 (N_2815,N_1503,N_1781);
or U2816 (N_2816,N_1903,N_1417);
nor U2817 (N_2817,N_1890,N_1054);
xnor U2818 (N_2818,N_1015,N_1851);
or U2819 (N_2819,N_1943,N_1894);
nor U2820 (N_2820,N_1453,N_1123);
or U2821 (N_2821,N_1228,N_1124);
nor U2822 (N_2822,N_1331,N_1020);
xor U2823 (N_2823,N_1141,N_1444);
xnor U2824 (N_2824,N_1867,N_1308);
nor U2825 (N_2825,N_1728,N_1913);
xor U2826 (N_2826,N_1592,N_1366);
nor U2827 (N_2827,N_1419,N_1869);
nor U2828 (N_2828,N_1943,N_1374);
or U2829 (N_2829,N_1557,N_1816);
nand U2830 (N_2830,N_1525,N_1038);
nor U2831 (N_2831,N_1708,N_1384);
and U2832 (N_2832,N_1005,N_1091);
or U2833 (N_2833,N_1924,N_1829);
nand U2834 (N_2834,N_1199,N_1334);
nor U2835 (N_2835,N_1990,N_1269);
nor U2836 (N_2836,N_1756,N_1343);
or U2837 (N_2837,N_1135,N_1205);
or U2838 (N_2838,N_1808,N_1419);
nor U2839 (N_2839,N_1197,N_1813);
xor U2840 (N_2840,N_1435,N_1746);
nor U2841 (N_2841,N_1963,N_1345);
xor U2842 (N_2842,N_1782,N_1274);
nand U2843 (N_2843,N_1046,N_1365);
xor U2844 (N_2844,N_1182,N_1915);
and U2845 (N_2845,N_1857,N_1183);
or U2846 (N_2846,N_1862,N_1376);
and U2847 (N_2847,N_1705,N_1719);
or U2848 (N_2848,N_1649,N_1155);
nand U2849 (N_2849,N_1625,N_1084);
and U2850 (N_2850,N_1739,N_1012);
xor U2851 (N_2851,N_1025,N_1800);
and U2852 (N_2852,N_1216,N_1322);
nand U2853 (N_2853,N_1030,N_1412);
or U2854 (N_2854,N_1603,N_1348);
or U2855 (N_2855,N_1720,N_1199);
or U2856 (N_2856,N_1400,N_1227);
nor U2857 (N_2857,N_1278,N_1983);
nand U2858 (N_2858,N_1479,N_1328);
xnor U2859 (N_2859,N_1011,N_1341);
and U2860 (N_2860,N_1409,N_1600);
xor U2861 (N_2861,N_1246,N_1546);
or U2862 (N_2862,N_1212,N_1741);
or U2863 (N_2863,N_1336,N_1677);
and U2864 (N_2864,N_1708,N_1316);
nand U2865 (N_2865,N_1456,N_1215);
nand U2866 (N_2866,N_1154,N_1847);
and U2867 (N_2867,N_1741,N_1833);
nor U2868 (N_2868,N_1222,N_1286);
and U2869 (N_2869,N_1327,N_1771);
and U2870 (N_2870,N_1096,N_1386);
nor U2871 (N_2871,N_1876,N_1042);
or U2872 (N_2872,N_1236,N_1730);
and U2873 (N_2873,N_1102,N_1110);
xnor U2874 (N_2874,N_1437,N_1636);
nor U2875 (N_2875,N_1250,N_1921);
nand U2876 (N_2876,N_1213,N_1192);
xor U2877 (N_2877,N_1657,N_1233);
and U2878 (N_2878,N_1445,N_1936);
or U2879 (N_2879,N_1080,N_1100);
or U2880 (N_2880,N_1999,N_1162);
or U2881 (N_2881,N_1638,N_1082);
nor U2882 (N_2882,N_1132,N_1599);
xnor U2883 (N_2883,N_1012,N_1760);
or U2884 (N_2884,N_1745,N_1380);
nand U2885 (N_2885,N_1571,N_1198);
nand U2886 (N_2886,N_1309,N_1830);
xor U2887 (N_2887,N_1227,N_1127);
and U2888 (N_2888,N_1248,N_1317);
nor U2889 (N_2889,N_1769,N_1072);
and U2890 (N_2890,N_1824,N_1906);
or U2891 (N_2891,N_1548,N_1049);
or U2892 (N_2892,N_1004,N_1933);
and U2893 (N_2893,N_1520,N_1334);
nor U2894 (N_2894,N_1714,N_1663);
and U2895 (N_2895,N_1801,N_1247);
nand U2896 (N_2896,N_1485,N_1771);
or U2897 (N_2897,N_1663,N_1762);
or U2898 (N_2898,N_1448,N_1976);
nor U2899 (N_2899,N_1351,N_1215);
xnor U2900 (N_2900,N_1709,N_1212);
nand U2901 (N_2901,N_1240,N_1799);
xor U2902 (N_2902,N_1836,N_1980);
and U2903 (N_2903,N_1089,N_1912);
or U2904 (N_2904,N_1425,N_1744);
xnor U2905 (N_2905,N_1279,N_1831);
xor U2906 (N_2906,N_1826,N_1938);
nand U2907 (N_2907,N_1958,N_1597);
xor U2908 (N_2908,N_1223,N_1215);
xnor U2909 (N_2909,N_1825,N_1646);
and U2910 (N_2910,N_1298,N_1674);
nor U2911 (N_2911,N_1427,N_1036);
or U2912 (N_2912,N_1328,N_1447);
and U2913 (N_2913,N_1457,N_1284);
nand U2914 (N_2914,N_1973,N_1533);
xor U2915 (N_2915,N_1686,N_1860);
or U2916 (N_2916,N_1006,N_1891);
nand U2917 (N_2917,N_1753,N_1582);
nor U2918 (N_2918,N_1362,N_1497);
nand U2919 (N_2919,N_1541,N_1542);
and U2920 (N_2920,N_1247,N_1061);
nor U2921 (N_2921,N_1414,N_1361);
and U2922 (N_2922,N_1704,N_1776);
and U2923 (N_2923,N_1330,N_1795);
or U2924 (N_2924,N_1833,N_1321);
nor U2925 (N_2925,N_1331,N_1144);
or U2926 (N_2926,N_1867,N_1824);
or U2927 (N_2927,N_1081,N_1715);
nor U2928 (N_2928,N_1390,N_1424);
or U2929 (N_2929,N_1395,N_1718);
nand U2930 (N_2930,N_1738,N_1943);
nand U2931 (N_2931,N_1080,N_1739);
or U2932 (N_2932,N_1566,N_1980);
and U2933 (N_2933,N_1264,N_1963);
nand U2934 (N_2934,N_1790,N_1588);
and U2935 (N_2935,N_1433,N_1948);
or U2936 (N_2936,N_1064,N_1767);
nand U2937 (N_2937,N_1864,N_1800);
or U2938 (N_2938,N_1740,N_1242);
nor U2939 (N_2939,N_1664,N_1411);
nand U2940 (N_2940,N_1259,N_1619);
nand U2941 (N_2941,N_1971,N_1115);
or U2942 (N_2942,N_1813,N_1072);
xor U2943 (N_2943,N_1976,N_1168);
nor U2944 (N_2944,N_1548,N_1733);
xnor U2945 (N_2945,N_1603,N_1439);
nand U2946 (N_2946,N_1324,N_1378);
or U2947 (N_2947,N_1497,N_1581);
nand U2948 (N_2948,N_1126,N_1863);
nor U2949 (N_2949,N_1954,N_1562);
nor U2950 (N_2950,N_1183,N_1489);
and U2951 (N_2951,N_1425,N_1006);
and U2952 (N_2952,N_1898,N_1876);
xnor U2953 (N_2953,N_1059,N_1922);
nor U2954 (N_2954,N_1901,N_1650);
nor U2955 (N_2955,N_1755,N_1406);
nor U2956 (N_2956,N_1304,N_1719);
and U2957 (N_2957,N_1780,N_1504);
and U2958 (N_2958,N_1585,N_1036);
and U2959 (N_2959,N_1256,N_1943);
or U2960 (N_2960,N_1678,N_1692);
nor U2961 (N_2961,N_1100,N_1646);
nand U2962 (N_2962,N_1389,N_1234);
xor U2963 (N_2963,N_1024,N_1107);
or U2964 (N_2964,N_1591,N_1081);
and U2965 (N_2965,N_1487,N_1529);
nor U2966 (N_2966,N_1703,N_1180);
xor U2967 (N_2967,N_1032,N_1577);
and U2968 (N_2968,N_1380,N_1419);
and U2969 (N_2969,N_1117,N_1672);
or U2970 (N_2970,N_1657,N_1125);
or U2971 (N_2971,N_1992,N_1237);
or U2972 (N_2972,N_1259,N_1744);
nand U2973 (N_2973,N_1999,N_1470);
nor U2974 (N_2974,N_1821,N_1582);
xor U2975 (N_2975,N_1534,N_1162);
or U2976 (N_2976,N_1651,N_1233);
or U2977 (N_2977,N_1802,N_1211);
xor U2978 (N_2978,N_1246,N_1369);
and U2979 (N_2979,N_1934,N_1619);
xnor U2980 (N_2980,N_1325,N_1383);
and U2981 (N_2981,N_1274,N_1349);
and U2982 (N_2982,N_1168,N_1945);
nor U2983 (N_2983,N_1274,N_1183);
or U2984 (N_2984,N_1808,N_1321);
xor U2985 (N_2985,N_1576,N_1527);
and U2986 (N_2986,N_1035,N_1813);
nand U2987 (N_2987,N_1710,N_1355);
nand U2988 (N_2988,N_1148,N_1806);
or U2989 (N_2989,N_1468,N_1013);
nand U2990 (N_2990,N_1565,N_1513);
xor U2991 (N_2991,N_1007,N_1609);
nand U2992 (N_2992,N_1207,N_1905);
nand U2993 (N_2993,N_1956,N_1962);
nor U2994 (N_2994,N_1286,N_1831);
and U2995 (N_2995,N_1879,N_1559);
and U2996 (N_2996,N_1988,N_1610);
nor U2997 (N_2997,N_1516,N_1112);
xnor U2998 (N_2998,N_1981,N_1392);
nand U2999 (N_2999,N_1467,N_1693);
nor U3000 (N_3000,N_2401,N_2311);
or U3001 (N_3001,N_2623,N_2417);
nor U3002 (N_3002,N_2461,N_2420);
nor U3003 (N_3003,N_2439,N_2016);
nor U3004 (N_3004,N_2823,N_2127);
and U3005 (N_3005,N_2858,N_2494);
nor U3006 (N_3006,N_2866,N_2309);
or U3007 (N_3007,N_2380,N_2470);
or U3008 (N_3008,N_2937,N_2749);
or U3009 (N_3009,N_2410,N_2226);
nand U3010 (N_3010,N_2617,N_2353);
and U3011 (N_3011,N_2169,N_2750);
xnor U3012 (N_3012,N_2041,N_2221);
and U3013 (N_3013,N_2554,N_2973);
nor U3014 (N_3014,N_2595,N_2718);
or U3015 (N_3015,N_2341,N_2174);
nor U3016 (N_3016,N_2443,N_2317);
or U3017 (N_3017,N_2789,N_2658);
nand U3018 (N_3018,N_2359,N_2728);
nand U3019 (N_3019,N_2824,N_2519);
xnor U3020 (N_3020,N_2388,N_2037);
and U3021 (N_3021,N_2030,N_2611);
or U3022 (N_3022,N_2576,N_2490);
xnor U3023 (N_3023,N_2269,N_2668);
and U3024 (N_3024,N_2477,N_2746);
and U3025 (N_3025,N_2367,N_2516);
xor U3026 (N_3026,N_2638,N_2276);
nand U3027 (N_3027,N_2508,N_2548);
or U3028 (N_3028,N_2721,N_2608);
xnor U3029 (N_3029,N_2830,N_2241);
nor U3030 (N_3030,N_2959,N_2000);
or U3031 (N_3031,N_2346,N_2374);
or U3032 (N_3032,N_2084,N_2408);
xor U3033 (N_3033,N_2072,N_2774);
nor U3034 (N_3034,N_2020,N_2334);
and U3035 (N_3035,N_2292,N_2969);
nand U3036 (N_3036,N_2135,N_2946);
or U3037 (N_3037,N_2647,N_2085);
or U3038 (N_3038,N_2115,N_2021);
and U3039 (N_3039,N_2726,N_2633);
or U3040 (N_3040,N_2808,N_2524);
nand U3041 (N_3041,N_2351,N_2087);
and U3042 (N_3042,N_2143,N_2971);
and U3043 (N_3043,N_2500,N_2216);
nand U3044 (N_3044,N_2887,N_2450);
or U3045 (N_3045,N_2755,N_2680);
and U3046 (N_3046,N_2395,N_2596);
xor U3047 (N_3047,N_2160,N_2600);
and U3048 (N_3048,N_2202,N_2869);
or U3049 (N_3049,N_2626,N_2274);
or U3050 (N_3050,N_2422,N_2104);
or U3051 (N_3051,N_2916,N_2511);
nand U3052 (N_3052,N_2102,N_2674);
nor U3053 (N_3053,N_2863,N_2393);
and U3054 (N_3054,N_2308,N_2144);
nor U3055 (N_3055,N_2938,N_2207);
xor U3056 (N_3056,N_2203,N_2448);
xor U3057 (N_3057,N_2200,N_2473);
and U3058 (N_3058,N_2909,N_2571);
nor U3059 (N_3059,N_2871,N_2430);
nand U3060 (N_3060,N_2224,N_2953);
or U3061 (N_3061,N_2319,N_2635);
xnor U3062 (N_3062,N_2483,N_2826);
nand U3063 (N_3063,N_2318,N_2819);
nand U3064 (N_3064,N_2418,N_2372);
nor U3065 (N_3065,N_2132,N_2167);
nand U3066 (N_3066,N_2384,N_2445);
nand U3067 (N_3067,N_2897,N_2933);
nand U3068 (N_3068,N_2504,N_2788);
or U3069 (N_3069,N_2109,N_2591);
or U3070 (N_3070,N_2099,N_2559);
xor U3071 (N_3071,N_2835,N_2485);
nand U3072 (N_3072,N_2773,N_2503);
xor U3073 (N_3073,N_2066,N_2427);
and U3074 (N_3074,N_2236,N_2431);
nand U3075 (N_3075,N_2853,N_2392);
xnor U3076 (N_3076,N_2211,N_2632);
nand U3077 (N_3077,N_2277,N_2995);
xor U3078 (N_3078,N_2634,N_2931);
nor U3079 (N_3079,N_2533,N_2337);
and U3080 (N_3080,N_2165,N_2088);
or U3081 (N_3081,N_2235,N_2506);
or U3082 (N_3082,N_2760,N_2197);
and U3083 (N_3083,N_2349,N_2093);
xor U3084 (N_3084,N_2272,N_2779);
xor U3085 (N_3085,N_2090,N_2042);
nand U3086 (N_3086,N_2368,N_2011);
nand U3087 (N_3087,N_2669,N_2809);
and U3088 (N_3088,N_2446,N_2238);
nor U3089 (N_3089,N_2345,N_2405);
nor U3090 (N_3090,N_2022,N_2950);
and U3091 (N_3091,N_2205,N_2312);
nor U3092 (N_3092,N_2720,N_2283);
nor U3093 (N_3093,N_2861,N_2191);
nor U3094 (N_3094,N_2284,N_2355);
nor U3095 (N_3095,N_2710,N_2057);
xor U3096 (N_3096,N_2570,N_2105);
or U3097 (N_3097,N_2291,N_2547);
xnor U3098 (N_3098,N_2204,N_2002);
nand U3099 (N_3099,N_2474,N_2754);
or U3100 (N_3100,N_2502,N_2069);
and U3101 (N_3101,N_2761,N_2336);
nor U3102 (N_3102,N_2872,N_2980);
nand U3103 (N_3103,N_2992,N_2537);
nand U3104 (N_3104,N_2817,N_2389);
nor U3105 (N_3105,N_2646,N_2192);
nand U3106 (N_3106,N_2925,N_2096);
or U3107 (N_3107,N_2112,N_2440);
nor U3108 (N_3108,N_2257,N_2320);
xnor U3109 (N_3109,N_2149,N_2364);
and U3110 (N_3110,N_2521,N_2219);
nand U3111 (N_3111,N_2074,N_2162);
nor U3112 (N_3112,N_2376,N_2326);
nor U3113 (N_3113,N_2759,N_2910);
xnor U3114 (N_3114,N_2766,N_2601);
nor U3115 (N_3115,N_2068,N_2052);
nor U3116 (N_3116,N_2438,N_2930);
nand U3117 (N_3117,N_2557,N_2715);
or U3118 (N_3118,N_2469,N_2286);
and U3119 (N_3119,N_2912,N_2048);
and U3120 (N_3120,N_2542,N_2703);
xnor U3121 (N_3121,N_2531,N_2199);
or U3122 (N_3122,N_2017,N_2491);
nor U3123 (N_3123,N_2731,N_2400);
nor U3124 (N_3124,N_2517,N_2498);
or U3125 (N_3125,N_2369,N_2957);
or U3126 (N_3126,N_2214,N_2907);
nand U3127 (N_3127,N_2509,N_2051);
and U3128 (N_3128,N_2541,N_2118);
nor U3129 (N_3129,N_2390,N_2184);
xor U3130 (N_3130,N_2700,N_2386);
or U3131 (N_3131,N_2613,N_2796);
and U3132 (N_3132,N_2151,N_2932);
xnor U3133 (N_3133,N_2990,N_2854);
or U3134 (N_3134,N_2860,N_2083);
or U3135 (N_3135,N_2295,N_2593);
and U3136 (N_3136,N_2639,N_2018);
nor U3137 (N_3137,N_2706,N_2044);
or U3138 (N_3138,N_2077,N_2507);
nor U3139 (N_3139,N_2232,N_2315);
and U3140 (N_3140,N_2078,N_2046);
nor U3141 (N_3141,N_2222,N_2810);
or U3142 (N_3142,N_2873,N_2194);
xor U3143 (N_3143,N_2765,N_2242);
nand U3144 (N_3144,N_2362,N_2103);
or U3145 (N_3145,N_2625,N_2347);
and U3146 (N_3146,N_2492,N_2421);
and U3147 (N_3147,N_2223,N_2079);
nor U3148 (N_3148,N_2486,N_2929);
nor U3149 (N_3149,N_2606,N_2574);
nor U3150 (N_3150,N_2956,N_2790);
nor U3151 (N_3151,N_2947,N_2268);
xor U3152 (N_3152,N_2629,N_2979);
nor U3153 (N_3153,N_2905,N_2831);
and U3154 (N_3154,N_2560,N_2894);
nor U3155 (N_3155,N_2131,N_2350);
nand U3156 (N_3156,N_2654,N_2913);
xor U3157 (N_3157,N_2514,N_2845);
nand U3158 (N_3158,N_2862,N_2186);
or U3159 (N_3159,N_2839,N_2949);
nor U3160 (N_3160,N_2164,N_2076);
nand U3161 (N_3161,N_2785,N_2058);
nand U3162 (N_3162,N_2073,N_2178);
xor U3163 (N_3163,N_2126,N_2966);
nand U3164 (N_3164,N_2459,N_2125);
nor U3165 (N_3165,N_2964,N_2177);
or U3166 (N_3166,N_2803,N_2451);
or U3167 (N_3167,N_2857,N_2049);
nor U3168 (N_3168,N_2140,N_2884);
nor U3169 (N_3169,N_2424,N_2665);
xnor U3170 (N_3170,N_2447,N_2371);
or U3171 (N_3171,N_2101,N_2047);
nand U3172 (N_3172,N_2651,N_2592);
nor U3173 (N_3173,N_2004,N_2114);
or U3174 (N_3174,N_2153,N_2195);
or U3175 (N_3175,N_2532,N_2702);
or U3176 (N_3176,N_2807,N_2024);
nor U3177 (N_3177,N_2977,N_2227);
and U3178 (N_3178,N_2050,N_2951);
xnor U3179 (N_3179,N_2425,N_2279);
nor U3180 (N_3180,N_2649,N_2888);
or U3181 (N_3181,N_2799,N_2482);
nand U3182 (N_3182,N_2928,N_2527);
nor U3183 (N_3183,N_2305,N_2027);
nand U3184 (N_3184,N_2786,N_2138);
and U3185 (N_3185,N_2842,N_2442);
or U3186 (N_3186,N_2480,N_2433);
nand U3187 (N_3187,N_2742,N_2847);
or U3188 (N_3188,N_2008,N_2610);
nor U3189 (N_3189,N_2210,N_2113);
and U3190 (N_3190,N_2373,N_2919);
and U3191 (N_3191,N_2762,N_2801);
or U3192 (N_3192,N_2339,N_2675);
xnor U3193 (N_3193,N_2997,N_2663);
nand U3194 (N_3194,N_2121,N_2695);
nor U3195 (N_3195,N_2147,N_2944);
nand U3196 (N_3196,N_2612,N_2399);
or U3197 (N_3197,N_2696,N_2117);
and U3198 (N_3198,N_2974,N_2539);
nor U3199 (N_3199,N_2730,N_2954);
xnor U3200 (N_3200,N_2978,N_2522);
nor U3201 (N_3201,N_2940,N_2895);
nor U3202 (N_3202,N_2465,N_2265);
or U3203 (N_3203,N_2429,N_2802);
nor U3204 (N_3204,N_2201,N_2917);
and U3205 (N_3205,N_2852,N_2218);
and U3206 (N_3206,N_2015,N_2397);
and U3207 (N_3207,N_2619,N_2264);
xnor U3208 (N_3208,N_2411,N_2948);
or U3209 (N_3209,N_2701,N_2587);
xor U3210 (N_3210,N_2678,N_2414);
nor U3211 (N_3211,N_2544,N_2379);
or U3212 (N_3212,N_2820,N_2900);
nor U3213 (N_3213,N_2206,N_2182);
nand U3214 (N_3214,N_2540,N_2981);
nor U3215 (N_3215,N_2994,N_2495);
nor U3216 (N_3216,N_2889,N_2825);
and U3217 (N_3217,N_2325,N_2436);
xor U3218 (N_3218,N_2775,N_2636);
xnor U3219 (N_3219,N_2816,N_2901);
or U3220 (N_3220,N_2868,N_2363);
and U3221 (N_3221,N_2179,N_2562);
nand U3222 (N_3222,N_2432,N_2784);
or U3223 (N_3223,N_2903,N_2130);
nand U3224 (N_3224,N_2588,N_2768);
xnor U3225 (N_3225,N_2941,N_2091);
or U3226 (N_3226,N_2984,N_2428);
and U3227 (N_3227,N_2187,N_2630);
nand U3228 (N_3228,N_2229,N_2882);
nor U3229 (N_3229,N_2920,N_2190);
nor U3230 (N_3230,N_2230,N_2094);
nand U3231 (N_3231,N_2444,N_2594);
xnor U3232 (N_3232,N_2158,N_2449);
nand U3233 (N_3233,N_2288,N_2829);
and U3234 (N_3234,N_2879,N_2965);
xor U3235 (N_3235,N_2770,N_2366);
and U3236 (N_3236,N_2124,N_2457);
nor U3237 (N_3237,N_2505,N_2468);
or U3238 (N_3238,N_2378,N_2526);
nand U3239 (N_3239,N_2566,N_2679);
or U3240 (N_3240,N_2855,N_2716);
and U3241 (N_3241,N_2725,N_2262);
and U3242 (N_3242,N_2426,N_2692);
nand U3243 (N_3243,N_2906,N_2189);
and U3244 (N_3244,N_2097,N_2381);
nor U3245 (N_3245,N_2253,N_2690);
nor U3246 (N_3246,N_2307,N_2342);
nor U3247 (N_3247,N_2813,N_2551);
and U3248 (N_3248,N_2840,N_2324);
or U3249 (N_3249,N_2166,N_2181);
or U3250 (N_3250,N_2510,N_2982);
xor U3251 (N_3251,N_2234,N_2038);
nor U3252 (N_3252,N_2299,N_2119);
and U3253 (N_3253,N_2106,N_2452);
nor U3254 (N_3254,N_2943,N_2838);
nand U3255 (N_3255,N_2719,N_2332);
and U3256 (N_3256,N_2806,N_2361);
nand U3257 (N_3257,N_2699,N_2598);
nand U3258 (N_3258,N_2565,N_2233);
nand U3259 (N_3259,N_2877,N_2159);
and U3260 (N_3260,N_2472,N_2063);
nand U3261 (N_3261,N_2846,N_2727);
or U3262 (N_3262,N_2603,N_2578);
xor U3263 (N_3263,N_2609,N_2689);
nor U3264 (N_3264,N_2120,N_2313);
nand U3265 (N_3265,N_2848,N_2331);
or U3266 (N_3266,N_2543,N_2275);
nor U3267 (N_3267,N_2215,N_2142);
nor U3268 (N_3268,N_2377,N_2797);
xnor U3269 (N_3269,N_2843,N_2059);
nand U3270 (N_3270,N_2391,N_2530);
or U3271 (N_3271,N_2653,N_2009);
xnor U3272 (N_3272,N_2743,N_2631);
and U3273 (N_3273,N_2758,N_2794);
xor U3274 (N_3274,N_2060,N_2375);
nor U3275 (N_3275,N_2403,N_2487);
nand U3276 (N_3276,N_2128,N_2248);
or U3277 (N_3277,N_2306,N_2735);
nand U3278 (N_3278,N_2952,N_2175);
xor U3279 (N_3279,N_2958,N_2180);
and U3280 (N_3280,N_2382,N_2012);
or U3281 (N_3281,N_2404,N_2471);
and U3282 (N_3282,N_2739,N_2423);
nor U3283 (N_3283,N_2891,N_2352);
and U3284 (N_3284,N_2267,N_2693);
xor U3285 (N_3285,N_2586,N_2890);
xor U3286 (N_3286,N_2314,N_2327);
or U3287 (N_3287,N_2316,N_2185);
nor U3288 (N_3288,N_2239,N_2585);
nor U3289 (N_3289,N_2805,N_2915);
and U3290 (N_3290,N_2053,N_2628);
and U3291 (N_3291,N_2518,N_2019);
or U3292 (N_3292,N_2407,N_2564);
nand U3293 (N_3293,N_2911,N_2589);
nor U3294 (N_3294,N_2732,N_2171);
nor U3295 (N_3295,N_2642,N_2927);
nor U3296 (N_3296,N_2338,N_2029);
xor U3297 (N_3297,N_2662,N_2737);
nor U3298 (N_3298,N_2798,N_2045);
nand U3299 (N_3299,N_2303,N_2864);
and U3300 (N_3300,N_2168,N_2258);
nor U3301 (N_3301,N_2032,N_2385);
nor U3302 (N_3302,N_2043,N_2462);
nor U3303 (N_3303,N_2714,N_2064);
xnor U3304 (N_3304,N_2875,N_2481);
nor U3305 (N_3305,N_2767,N_2605);
nand U3306 (N_3306,N_2294,N_2659);
xnor U3307 (N_3307,N_2014,N_2682);
nand U3308 (N_3308,N_2252,N_2455);
or U3309 (N_3309,N_2479,N_2967);
nand U3310 (N_3310,N_2095,N_2552);
or U3311 (N_3311,N_2133,N_2358);
xnor U3312 (N_3312,N_2081,N_2070);
or U3313 (N_3313,N_2985,N_2246);
xor U3314 (N_3314,N_2599,N_2323);
and U3315 (N_3315,N_2413,N_2711);
and U3316 (N_3316,N_2523,N_2225);
nor U3317 (N_3317,N_2828,N_2260);
or U3318 (N_3318,N_2643,N_2661);
and U3319 (N_3319,N_2056,N_2496);
nor U3320 (N_3320,N_2525,N_2415);
nor U3321 (N_3321,N_2529,N_2939);
xnor U3322 (N_3322,N_2263,N_2736);
or U3323 (N_3323,N_2163,N_2859);
nand U3324 (N_3324,N_2991,N_2899);
nand U3325 (N_3325,N_2034,N_2209);
and U3326 (N_3326,N_2033,N_2466);
xnor U3327 (N_3327,N_2614,N_2188);
xnor U3328 (N_3328,N_2827,N_2281);
nor U3329 (N_3329,N_2025,N_2934);
and U3330 (N_3330,N_2987,N_2579);
and U3331 (N_3331,N_2387,N_2712);
nor U3332 (N_3332,N_2244,N_2963);
and U3333 (N_3333,N_2467,N_2935);
or U3334 (N_3334,N_2989,N_2818);
or U3335 (N_3335,N_2792,N_2183);
nand U3336 (N_3336,N_2691,N_2893);
xnor U3337 (N_3337,N_2580,N_2454);
or U3338 (N_3338,N_2584,N_2620);
or U3339 (N_3339,N_2329,N_2146);
nand U3340 (N_3340,N_2285,N_2412);
and U3341 (N_3341,N_2741,N_2793);
nand U3342 (N_3342,N_2247,N_2771);
nor U3343 (N_3343,N_2534,N_2968);
nor U3344 (N_3344,N_2561,N_2441);
and U3345 (N_3345,N_2667,N_2322);
xor U3346 (N_3346,N_2804,N_2627);
or U3347 (N_3347,N_2370,N_2110);
or U3348 (N_3348,N_2256,N_2815);
nor U3349 (N_3349,N_2228,N_2220);
nand U3350 (N_3350,N_2249,N_2139);
xnor U3351 (N_3351,N_2898,N_2394);
nand U3352 (N_3352,N_2409,N_2867);
or U3353 (N_3353,N_2856,N_2876);
xnor U3354 (N_3354,N_2217,N_2333);
xor U3355 (N_3355,N_2962,N_2621);
and U3356 (N_3356,N_2681,N_2670);
xor U3357 (N_3357,N_2787,N_2499);
and U3358 (N_3358,N_2812,N_2243);
or U3359 (N_3359,N_2035,N_2713);
xor U3360 (N_3360,N_2535,N_2054);
nor U3361 (N_3361,N_2092,N_2883);
nor U3362 (N_3362,N_2708,N_2777);
xor U3363 (N_3363,N_2513,N_2624);
nor U3364 (N_3364,N_2672,N_2955);
xnor U3365 (N_3365,N_2137,N_2604);
xor U3366 (N_3366,N_2040,N_2172);
or U3367 (N_3367,N_2098,N_2640);
or U3368 (N_3368,N_2908,N_2023);
xnor U3369 (N_3369,N_2841,N_2729);
xnor U3370 (N_3370,N_2763,N_2237);
nor U3371 (N_3371,N_2145,N_2273);
nand U3372 (N_3372,N_2751,N_2581);
and U3373 (N_3373,N_2833,N_2383);
xor U3374 (N_3374,N_2936,N_2772);
nand U3375 (N_3375,N_2563,N_2549);
nor U3376 (N_3376,N_2707,N_2902);
xor U3377 (N_3377,N_2822,N_2055);
nand U3378 (N_3378,N_2301,N_2031);
and U3379 (N_3379,N_2402,N_2880);
nor U3380 (N_3380,N_2924,N_2321);
xor U3381 (N_3381,N_2489,N_2512);
nor U3382 (N_3382,N_2709,N_2278);
nand U3383 (N_3383,N_2302,N_2289);
nand U3384 (N_3384,N_2255,N_2501);
or U3385 (N_3385,N_2811,N_2136);
nor U3386 (N_3386,N_2983,N_2365);
or U3387 (N_3387,N_2849,N_2569);
and U3388 (N_3388,N_2999,N_2271);
and U3389 (N_3389,N_2006,N_2615);
and U3390 (N_3390,N_2434,N_2607);
nor U3391 (N_3391,N_2567,N_2821);
or U3392 (N_3392,N_2546,N_2697);
nor U3393 (N_3393,N_2622,N_2800);
nor U3394 (N_3394,N_2300,N_2769);
nor U3395 (N_3395,N_2885,N_2155);
nand U3396 (N_3396,N_2998,N_2280);
or U3397 (N_3397,N_2437,N_2922);
xnor U3398 (N_3398,N_2001,N_2780);
and U3399 (N_3399,N_2553,N_2666);
nand U3400 (N_3400,N_2173,N_2791);
or U3401 (N_3401,N_2976,N_2213);
nand U3402 (N_3402,N_2705,N_2003);
or U3403 (N_3403,N_2328,N_2590);
or U3404 (N_3404,N_2484,N_2538);
and U3405 (N_3405,N_2007,N_2193);
and U3406 (N_3406,N_2597,N_2488);
xnor U3407 (N_3407,N_2161,N_2704);
nor U3408 (N_3408,N_2684,N_2671);
nand U3409 (N_3409,N_2677,N_2686);
nor U3410 (N_3410,N_2343,N_2129);
nor U3411 (N_3411,N_2111,N_2988);
nor U3412 (N_3412,N_2896,N_2497);
xor U3413 (N_3413,N_2108,N_2918);
nand U3414 (N_3414,N_2198,N_2694);
and U3415 (N_3415,N_2722,N_2290);
nand U3416 (N_3416,N_2536,N_2348);
xor U3417 (N_3417,N_2745,N_2287);
nand U3418 (N_3418,N_2583,N_2028);
and U3419 (N_3419,N_2254,N_2738);
or U3420 (N_3420,N_2107,N_2764);
nor U3421 (N_3421,N_2116,N_2558);
nand U3422 (N_3422,N_2396,N_2556);
xor U3423 (N_3423,N_2354,N_2756);
nand U3424 (N_3424,N_2656,N_2170);
and U3425 (N_3425,N_2753,N_2075);
xor U3426 (N_3426,N_2575,N_2357);
or U3427 (N_3427,N_2961,N_2356);
nand U3428 (N_3428,N_2850,N_2795);
nor U3429 (N_3429,N_2086,N_2717);
and U3430 (N_3430,N_2881,N_2259);
nor U3431 (N_3431,N_2212,N_2698);
nor U3432 (N_3432,N_2344,N_2993);
xor U3433 (N_3433,N_2250,N_2089);
xor U3434 (N_3434,N_2945,N_2520);
and U3435 (N_3435,N_2655,N_2062);
or U3436 (N_3436,N_2005,N_2456);
nor U3437 (N_3437,N_2757,N_2834);
or U3438 (N_3438,N_2748,N_2435);
xnor U3439 (N_3439,N_2419,N_2865);
nor U3440 (N_3440,N_2781,N_2026);
nor U3441 (N_3441,N_2196,N_2874);
nand U3442 (N_3442,N_2261,N_2723);
xnor U3443 (N_3443,N_2878,N_2996);
or U3444 (N_3444,N_2776,N_2618);
and U3445 (N_3445,N_2778,N_2747);
and U3446 (N_3446,N_2645,N_2270);
or U3447 (N_3447,N_2602,N_2231);
xor U3448 (N_3448,N_2061,N_2039);
nor U3449 (N_3449,N_2687,N_2582);
or U3450 (N_3450,N_2475,N_2464);
nand U3451 (N_3451,N_2036,N_2648);
nor U3452 (N_3452,N_2340,N_2071);
and U3453 (N_3453,N_2572,N_2975);
and U3454 (N_3454,N_2152,N_2515);
or U3455 (N_3455,N_2870,N_2310);
and U3456 (N_3456,N_2904,N_2360);
and U3457 (N_3457,N_2245,N_2463);
xor U3458 (N_3458,N_2154,N_2157);
or U3459 (N_3459,N_2555,N_2100);
nor U3460 (N_3460,N_2676,N_2914);
nor U3461 (N_3461,N_2067,N_2851);
nor U3462 (N_3462,N_2550,N_2065);
and U3463 (N_3463,N_2782,N_2493);
and U3464 (N_3464,N_2685,N_2148);
or U3465 (N_3465,N_2740,N_2733);
nand U3466 (N_3466,N_2573,N_2960);
nor U3467 (N_3467,N_2293,N_2082);
nand U3468 (N_3468,N_2123,N_2296);
nor U3469 (N_3469,N_2568,N_2783);
nor U3470 (N_3470,N_2832,N_2266);
nor U3471 (N_3471,N_2970,N_2837);
nor U3472 (N_3472,N_2010,N_2458);
xor U3473 (N_3473,N_2298,N_2013);
nor U3474 (N_3474,N_2986,N_2886);
or U3475 (N_3475,N_2923,N_2644);
and U3476 (N_3476,N_2416,N_2453);
xnor U3477 (N_3477,N_2080,N_2673);
nand U3478 (N_3478,N_2282,N_2926);
and U3479 (N_3479,N_2921,N_2688);
nor U3480 (N_3480,N_2657,N_2134);
or U3481 (N_3481,N_2724,N_2297);
and U3482 (N_3482,N_2616,N_2330);
or U3483 (N_3483,N_2528,N_2122);
nand U3484 (N_3484,N_2476,N_2844);
and U3485 (N_3485,N_2150,N_2942);
and U3486 (N_3486,N_2251,N_2972);
and U3487 (N_3487,N_2460,N_2156);
nor U3488 (N_3488,N_2141,N_2545);
or U3489 (N_3489,N_2398,N_2652);
xnor U3490 (N_3490,N_2577,N_2660);
nand U3491 (N_3491,N_2176,N_2892);
nand U3492 (N_3492,N_2752,N_2836);
nor U3493 (N_3493,N_2683,N_2744);
xnor U3494 (N_3494,N_2814,N_2304);
nand U3495 (N_3495,N_2637,N_2641);
xnor U3496 (N_3496,N_2406,N_2664);
and U3497 (N_3497,N_2208,N_2478);
xnor U3498 (N_3498,N_2240,N_2335);
or U3499 (N_3499,N_2650,N_2734);
nand U3500 (N_3500,N_2840,N_2687);
or U3501 (N_3501,N_2587,N_2973);
xnor U3502 (N_3502,N_2304,N_2733);
nor U3503 (N_3503,N_2597,N_2319);
nor U3504 (N_3504,N_2740,N_2797);
and U3505 (N_3505,N_2862,N_2458);
nor U3506 (N_3506,N_2744,N_2160);
nor U3507 (N_3507,N_2780,N_2174);
xnor U3508 (N_3508,N_2714,N_2229);
nor U3509 (N_3509,N_2984,N_2728);
nand U3510 (N_3510,N_2214,N_2635);
nand U3511 (N_3511,N_2397,N_2109);
and U3512 (N_3512,N_2197,N_2927);
nand U3513 (N_3513,N_2641,N_2108);
xor U3514 (N_3514,N_2649,N_2107);
and U3515 (N_3515,N_2927,N_2834);
nor U3516 (N_3516,N_2974,N_2394);
and U3517 (N_3517,N_2175,N_2794);
xnor U3518 (N_3518,N_2327,N_2723);
xnor U3519 (N_3519,N_2212,N_2352);
xor U3520 (N_3520,N_2193,N_2413);
xnor U3521 (N_3521,N_2663,N_2468);
xnor U3522 (N_3522,N_2831,N_2333);
xnor U3523 (N_3523,N_2103,N_2981);
and U3524 (N_3524,N_2969,N_2525);
xnor U3525 (N_3525,N_2039,N_2128);
or U3526 (N_3526,N_2390,N_2693);
xor U3527 (N_3527,N_2885,N_2664);
nand U3528 (N_3528,N_2992,N_2737);
xor U3529 (N_3529,N_2723,N_2822);
xor U3530 (N_3530,N_2444,N_2550);
and U3531 (N_3531,N_2159,N_2944);
xor U3532 (N_3532,N_2097,N_2216);
nand U3533 (N_3533,N_2635,N_2231);
or U3534 (N_3534,N_2289,N_2474);
nor U3535 (N_3535,N_2189,N_2186);
nor U3536 (N_3536,N_2127,N_2554);
or U3537 (N_3537,N_2722,N_2332);
and U3538 (N_3538,N_2876,N_2543);
nor U3539 (N_3539,N_2363,N_2057);
nor U3540 (N_3540,N_2846,N_2852);
and U3541 (N_3541,N_2267,N_2894);
and U3542 (N_3542,N_2276,N_2862);
or U3543 (N_3543,N_2045,N_2800);
xor U3544 (N_3544,N_2721,N_2370);
nand U3545 (N_3545,N_2462,N_2795);
xor U3546 (N_3546,N_2301,N_2868);
nand U3547 (N_3547,N_2857,N_2319);
nand U3548 (N_3548,N_2883,N_2120);
nor U3549 (N_3549,N_2099,N_2749);
nand U3550 (N_3550,N_2945,N_2309);
or U3551 (N_3551,N_2223,N_2393);
nand U3552 (N_3552,N_2376,N_2897);
and U3553 (N_3553,N_2290,N_2664);
and U3554 (N_3554,N_2576,N_2005);
nand U3555 (N_3555,N_2699,N_2032);
or U3556 (N_3556,N_2147,N_2263);
xnor U3557 (N_3557,N_2875,N_2126);
nor U3558 (N_3558,N_2454,N_2286);
or U3559 (N_3559,N_2614,N_2036);
xor U3560 (N_3560,N_2952,N_2505);
xnor U3561 (N_3561,N_2366,N_2231);
nor U3562 (N_3562,N_2449,N_2386);
nand U3563 (N_3563,N_2256,N_2700);
or U3564 (N_3564,N_2993,N_2551);
nand U3565 (N_3565,N_2384,N_2191);
xor U3566 (N_3566,N_2069,N_2178);
and U3567 (N_3567,N_2353,N_2345);
or U3568 (N_3568,N_2899,N_2058);
xor U3569 (N_3569,N_2290,N_2556);
and U3570 (N_3570,N_2793,N_2014);
or U3571 (N_3571,N_2889,N_2139);
nor U3572 (N_3572,N_2191,N_2455);
and U3573 (N_3573,N_2436,N_2235);
nor U3574 (N_3574,N_2920,N_2384);
or U3575 (N_3575,N_2967,N_2136);
nor U3576 (N_3576,N_2885,N_2666);
nand U3577 (N_3577,N_2128,N_2981);
and U3578 (N_3578,N_2936,N_2344);
xor U3579 (N_3579,N_2879,N_2074);
nor U3580 (N_3580,N_2932,N_2573);
or U3581 (N_3581,N_2722,N_2936);
nand U3582 (N_3582,N_2513,N_2809);
or U3583 (N_3583,N_2539,N_2940);
nand U3584 (N_3584,N_2484,N_2980);
xnor U3585 (N_3585,N_2340,N_2625);
nor U3586 (N_3586,N_2673,N_2340);
and U3587 (N_3587,N_2951,N_2453);
and U3588 (N_3588,N_2202,N_2169);
and U3589 (N_3589,N_2257,N_2346);
and U3590 (N_3590,N_2493,N_2980);
nand U3591 (N_3591,N_2290,N_2076);
or U3592 (N_3592,N_2382,N_2281);
nor U3593 (N_3593,N_2419,N_2372);
nor U3594 (N_3594,N_2380,N_2820);
and U3595 (N_3595,N_2417,N_2331);
or U3596 (N_3596,N_2779,N_2337);
nand U3597 (N_3597,N_2866,N_2775);
nand U3598 (N_3598,N_2930,N_2994);
xnor U3599 (N_3599,N_2057,N_2568);
xnor U3600 (N_3600,N_2037,N_2561);
or U3601 (N_3601,N_2324,N_2235);
xnor U3602 (N_3602,N_2745,N_2636);
or U3603 (N_3603,N_2109,N_2214);
or U3604 (N_3604,N_2748,N_2659);
nor U3605 (N_3605,N_2295,N_2699);
and U3606 (N_3606,N_2811,N_2675);
nor U3607 (N_3607,N_2847,N_2836);
and U3608 (N_3608,N_2059,N_2985);
xor U3609 (N_3609,N_2662,N_2198);
xor U3610 (N_3610,N_2296,N_2535);
xor U3611 (N_3611,N_2339,N_2798);
nand U3612 (N_3612,N_2760,N_2209);
nand U3613 (N_3613,N_2016,N_2187);
and U3614 (N_3614,N_2128,N_2669);
and U3615 (N_3615,N_2279,N_2471);
and U3616 (N_3616,N_2077,N_2818);
or U3617 (N_3617,N_2446,N_2722);
xor U3618 (N_3618,N_2051,N_2467);
nand U3619 (N_3619,N_2961,N_2497);
and U3620 (N_3620,N_2895,N_2137);
or U3621 (N_3621,N_2521,N_2642);
xor U3622 (N_3622,N_2269,N_2962);
nand U3623 (N_3623,N_2170,N_2069);
xnor U3624 (N_3624,N_2643,N_2578);
nor U3625 (N_3625,N_2090,N_2939);
and U3626 (N_3626,N_2094,N_2398);
nand U3627 (N_3627,N_2963,N_2199);
xnor U3628 (N_3628,N_2863,N_2570);
nand U3629 (N_3629,N_2064,N_2711);
or U3630 (N_3630,N_2781,N_2796);
and U3631 (N_3631,N_2439,N_2039);
nand U3632 (N_3632,N_2401,N_2235);
and U3633 (N_3633,N_2543,N_2463);
nand U3634 (N_3634,N_2849,N_2684);
xor U3635 (N_3635,N_2543,N_2420);
xnor U3636 (N_3636,N_2858,N_2435);
nor U3637 (N_3637,N_2054,N_2511);
and U3638 (N_3638,N_2605,N_2733);
nor U3639 (N_3639,N_2689,N_2091);
xor U3640 (N_3640,N_2302,N_2725);
nand U3641 (N_3641,N_2419,N_2509);
nor U3642 (N_3642,N_2880,N_2719);
or U3643 (N_3643,N_2893,N_2586);
and U3644 (N_3644,N_2076,N_2051);
and U3645 (N_3645,N_2400,N_2399);
xnor U3646 (N_3646,N_2172,N_2383);
nand U3647 (N_3647,N_2311,N_2885);
and U3648 (N_3648,N_2581,N_2578);
xor U3649 (N_3649,N_2565,N_2933);
and U3650 (N_3650,N_2818,N_2613);
nor U3651 (N_3651,N_2516,N_2394);
nor U3652 (N_3652,N_2978,N_2594);
xnor U3653 (N_3653,N_2299,N_2841);
nand U3654 (N_3654,N_2073,N_2433);
nand U3655 (N_3655,N_2969,N_2512);
xor U3656 (N_3656,N_2172,N_2887);
xor U3657 (N_3657,N_2387,N_2257);
and U3658 (N_3658,N_2641,N_2377);
and U3659 (N_3659,N_2865,N_2478);
and U3660 (N_3660,N_2805,N_2907);
nand U3661 (N_3661,N_2815,N_2886);
nor U3662 (N_3662,N_2539,N_2102);
and U3663 (N_3663,N_2410,N_2807);
and U3664 (N_3664,N_2729,N_2700);
nand U3665 (N_3665,N_2865,N_2670);
nor U3666 (N_3666,N_2340,N_2055);
xor U3667 (N_3667,N_2927,N_2890);
and U3668 (N_3668,N_2834,N_2058);
nor U3669 (N_3669,N_2572,N_2783);
and U3670 (N_3670,N_2118,N_2273);
nor U3671 (N_3671,N_2756,N_2161);
nand U3672 (N_3672,N_2993,N_2140);
nor U3673 (N_3673,N_2828,N_2079);
nor U3674 (N_3674,N_2917,N_2850);
and U3675 (N_3675,N_2836,N_2026);
and U3676 (N_3676,N_2394,N_2733);
nand U3677 (N_3677,N_2746,N_2785);
and U3678 (N_3678,N_2093,N_2428);
nand U3679 (N_3679,N_2397,N_2114);
or U3680 (N_3680,N_2736,N_2599);
nor U3681 (N_3681,N_2403,N_2885);
nor U3682 (N_3682,N_2559,N_2124);
or U3683 (N_3683,N_2661,N_2452);
or U3684 (N_3684,N_2568,N_2127);
nor U3685 (N_3685,N_2123,N_2605);
and U3686 (N_3686,N_2562,N_2046);
and U3687 (N_3687,N_2955,N_2153);
or U3688 (N_3688,N_2511,N_2436);
nor U3689 (N_3689,N_2193,N_2526);
nor U3690 (N_3690,N_2286,N_2236);
or U3691 (N_3691,N_2938,N_2540);
xnor U3692 (N_3692,N_2402,N_2109);
nand U3693 (N_3693,N_2111,N_2136);
nor U3694 (N_3694,N_2838,N_2029);
nor U3695 (N_3695,N_2588,N_2532);
nor U3696 (N_3696,N_2556,N_2227);
nand U3697 (N_3697,N_2569,N_2039);
nand U3698 (N_3698,N_2366,N_2759);
xor U3699 (N_3699,N_2365,N_2497);
and U3700 (N_3700,N_2406,N_2603);
or U3701 (N_3701,N_2657,N_2851);
nor U3702 (N_3702,N_2560,N_2721);
and U3703 (N_3703,N_2400,N_2872);
nand U3704 (N_3704,N_2988,N_2243);
nand U3705 (N_3705,N_2570,N_2910);
and U3706 (N_3706,N_2428,N_2925);
and U3707 (N_3707,N_2149,N_2676);
nor U3708 (N_3708,N_2914,N_2915);
xnor U3709 (N_3709,N_2639,N_2158);
nor U3710 (N_3710,N_2891,N_2026);
nor U3711 (N_3711,N_2327,N_2384);
and U3712 (N_3712,N_2348,N_2312);
or U3713 (N_3713,N_2275,N_2307);
nand U3714 (N_3714,N_2476,N_2313);
xnor U3715 (N_3715,N_2684,N_2745);
and U3716 (N_3716,N_2606,N_2190);
nor U3717 (N_3717,N_2703,N_2581);
nor U3718 (N_3718,N_2447,N_2482);
or U3719 (N_3719,N_2510,N_2314);
or U3720 (N_3720,N_2768,N_2730);
and U3721 (N_3721,N_2385,N_2779);
xnor U3722 (N_3722,N_2428,N_2653);
or U3723 (N_3723,N_2276,N_2440);
and U3724 (N_3724,N_2836,N_2098);
nand U3725 (N_3725,N_2498,N_2474);
nor U3726 (N_3726,N_2813,N_2300);
or U3727 (N_3727,N_2495,N_2932);
and U3728 (N_3728,N_2553,N_2530);
nor U3729 (N_3729,N_2674,N_2301);
nand U3730 (N_3730,N_2615,N_2223);
nand U3731 (N_3731,N_2171,N_2194);
nor U3732 (N_3732,N_2962,N_2822);
or U3733 (N_3733,N_2911,N_2016);
nand U3734 (N_3734,N_2743,N_2519);
and U3735 (N_3735,N_2862,N_2356);
or U3736 (N_3736,N_2596,N_2564);
and U3737 (N_3737,N_2014,N_2605);
nand U3738 (N_3738,N_2850,N_2623);
nand U3739 (N_3739,N_2483,N_2119);
nand U3740 (N_3740,N_2102,N_2476);
xnor U3741 (N_3741,N_2945,N_2721);
and U3742 (N_3742,N_2421,N_2945);
or U3743 (N_3743,N_2650,N_2822);
nand U3744 (N_3744,N_2388,N_2050);
and U3745 (N_3745,N_2864,N_2847);
and U3746 (N_3746,N_2658,N_2311);
xnor U3747 (N_3747,N_2374,N_2465);
and U3748 (N_3748,N_2595,N_2707);
or U3749 (N_3749,N_2195,N_2905);
xnor U3750 (N_3750,N_2746,N_2963);
nand U3751 (N_3751,N_2439,N_2554);
nor U3752 (N_3752,N_2505,N_2243);
or U3753 (N_3753,N_2499,N_2443);
xnor U3754 (N_3754,N_2157,N_2217);
xor U3755 (N_3755,N_2268,N_2979);
nand U3756 (N_3756,N_2690,N_2380);
and U3757 (N_3757,N_2330,N_2792);
nor U3758 (N_3758,N_2323,N_2531);
or U3759 (N_3759,N_2393,N_2674);
xor U3760 (N_3760,N_2487,N_2964);
xor U3761 (N_3761,N_2140,N_2658);
or U3762 (N_3762,N_2790,N_2767);
nor U3763 (N_3763,N_2729,N_2842);
and U3764 (N_3764,N_2845,N_2759);
nand U3765 (N_3765,N_2002,N_2005);
nand U3766 (N_3766,N_2053,N_2200);
nor U3767 (N_3767,N_2835,N_2933);
xnor U3768 (N_3768,N_2661,N_2741);
nand U3769 (N_3769,N_2629,N_2438);
or U3770 (N_3770,N_2468,N_2267);
and U3771 (N_3771,N_2403,N_2038);
or U3772 (N_3772,N_2868,N_2186);
nor U3773 (N_3773,N_2626,N_2221);
nand U3774 (N_3774,N_2826,N_2536);
and U3775 (N_3775,N_2744,N_2786);
nor U3776 (N_3776,N_2477,N_2591);
and U3777 (N_3777,N_2621,N_2728);
nand U3778 (N_3778,N_2566,N_2200);
nand U3779 (N_3779,N_2364,N_2233);
or U3780 (N_3780,N_2537,N_2012);
nand U3781 (N_3781,N_2613,N_2825);
and U3782 (N_3782,N_2793,N_2752);
xnor U3783 (N_3783,N_2723,N_2403);
xnor U3784 (N_3784,N_2464,N_2752);
and U3785 (N_3785,N_2313,N_2391);
and U3786 (N_3786,N_2369,N_2571);
xor U3787 (N_3787,N_2968,N_2897);
nand U3788 (N_3788,N_2268,N_2975);
nor U3789 (N_3789,N_2063,N_2058);
and U3790 (N_3790,N_2890,N_2648);
nor U3791 (N_3791,N_2701,N_2728);
nand U3792 (N_3792,N_2812,N_2245);
xnor U3793 (N_3793,N_2466,N_2629);
or U3794 (N_3794,N_2904,N_2756);
nor U3795 (N_3795,N_2177,N_2332);
xnor U3796 (N_3796,N_2087,N_2884);
or U3797 (N_3797,N_2688,N_2322);
nor U3798 (N_3798,N_2254,N_2069);
and U3799 (N_3799,N_2461,N_2576);
xnor U3800 (N_3800,N_2923,N_2320);
nor U3801 (N_3801,N_2694,N_2032);
nand U3802 (N_3802,N_2367,N_2976);
nand U3803 (N_3803,N_2704,N_2019);
nand U3804 (N_3804,N_2726,N_2942);
nand U3805 (N_3805,N_2636,N_2525);
xnor U3806 (N_3806,N_2858,N_2649);
and U3807 (N_3807,N_2797,N_2458);
nor U3808 (N_3808,N_2862,N_2763);
nor U3809 (N_3809,N_2763,N_2086);
or U3810 (N_3810,N_2445,N_2948);
or U3811 (N_3811,N_2770,N_2198);
and U3812 (N_3812,N_2347,N_2388);
nor U3813 (N_3813,N_2964,N_2156);
nor U3814 (N_3814,N_2633,N_2606);
nor U3815 (N_3815,N_2119,N_2225);
or U3816 (N_3816,N_2416,N_2465);
xnor U3817 (N_3817,N_2473,N_2752);
xor U3818 (N_3818,N_2243,N_2919);
or U3819 (N_3819,N_2662,N_2034);
xnor U3820 (N_3820,N_2394,N_2249);
and U3821 (N_3821,N_2754,N_2496);
or U3822 (N_3822,N_2134,N_2103);
and U3823 (N_3823,N_2670,N_2095);
nor U3824 (N_3824,N_2392,N_2698);
or U3825 (N_3825,N_2018,N_2535);
and U3826 (N_3826,N_2300,N_2698);
xnor U3827 (N_3827,N_2151,N_2510);
nor U3828 (N_3828,N_2325,N_2817);
nand U3829 (N_3829,N_2319,N_2009);
or U3830 (N_3830,N_2798,N_2817);
xnor U3831 (N_3831,N_2804,N_2245);
and U3832 (N_3832,N_2505,N_2022);
nor U3833 (N_3833,N_2429,N_2086);
nor U3834 (N_3834,N_2901,N_2894);
or U3835 (N_3835,N_2807,N_2920);
xor U3836 (N_3836,N_2635,N_2661);
or U3837 (N_3837,N_2612,N_2253);
nand U3838 (N_3838,N_2142,N_2431);
nor U3839 (N_3839,N_2470,N_2149);
and U3840 (N_3840,N_2107,N_2682);
and U3841 (N_3841,N_2761,N_2518);
nand U3842 (N_3842,N_2811,N_2321);
xor U3843 (N_3843,N_2729,N_2719);
and U3844 (N_3844,N_2616,N_2785);
nor U3845 (N_3845,N_2107,N_2566);
nor U3846 (N_3846,N_2655,N_2735);
and U3847 (N_3847,N_2659,N_2357);
nor U3848 (N_3848,N_2614,N_2217);
and U3849 (N_3849,N_2402,N_2986);
and U3850 (N_3850,N_2240,N_2647);
nand U3851 (N_3851,N_2896,N_2562);
and U3852 (N_3852,N_2364,N_2164);
and U3853 (N_3853,N_2245,N_2476);
xor U3854 (N_3854,N_2636,N_2583);
and U3855 (N_3855,N_2545,N_2521);
nand U3856 (N_3856,N_2075,N_2746);
nand U3857 (N_3857,N_2300,N_2096);
or U3858 (N_3858,N_2487,N_2842);
xor U3859 (N_3859,N_2099,N_2772);
nor U3860 (N_3860,N_2460,N_2358);
and U3861 (N_3861,N_2870,N_2752);
nand U3862 (N_3862,N_2974,N_2864);
nand U3863 (N_3863,N_2842,N_2546);
or U3864 (N_3864,N_2832,N_2440);
and U3865 (N_3865,N_2233,N_2744);
nor U3866 (N_3866,N_2272,N_2618);
and U3867 (N_3867,N_2315,N_2600);
nand U3868 (N_3868,N_2529,N_2739);
and U3869 (N_3869,N_2697,N_2067);
and U3870 (N_3870,N_2335,N_2469);
nor U3871 (N_3871,N_2700,N_2298);
and U3872 (N_3872,N_2211,N_2767);
nor U3873 (N_3873,N_2906,N_2849);
nand U3874 (N_3874,N_2014,N_2267);
nor U3875 (N_3875,N_2542,N_2085);
xor U3876 (N_3876,N_2461,N_2784);
xor U3877 (N_3877,N_2080,N_2982);
nor U3878 (N_3878,N_2618,N_2175);
and U3879 (N_3879,N_2929,N_2238);
or U3880 (N_3880,N_2115,N_2742);
xor U3881 (N_3881,N_2227,N_2936);
nor U3882 (N_3882,N_2293,N_2579);
nor U3883 (N_3883,N_2074,N_2070);
or U3884 (N_3884,N_2573,N_2832);
xnor U3885 (N_3885,N_2193,N_2148);
xnor U3886 (N_3886,N_2629,N_2546);
or U3887 (N_3887,N_2434,N_2569);
nor U3888 (N_3888,N_2348,N_2478);
and U3889 (N_3889,N_2201,N_2143);
and U3890 (N_3890,N_2131,N_2561);
xor U3891 (N_3891,N_2578,N_2488);
and U3892 (N_3892,N_2161,N_2571);
or U3893 (N_3893,N_2580,N_2271);
and U3894 (N_3894,N_2403,N_2647);
nand U3895 (N_3895,N_2510,N_2443);
xnor U3896 (N_3896,N_2589,N_2406);
nor U3897 (N_3897,N_2940,N_2833);
nand U3898 (N_3898,N_2354,N_2657);
nand U3899 (N_3899,N_2832,N_2891);
and U3900 (N_3900,N_2010,N_2994);
xor U3901 (N_3901,N_2112,N_2294);
nor U3902 (N_3902,N_2383,N_2028);
and U3903 (N_3903,N_2450,N_2386);
xor U3904 (N_3904,N_2007,N_2516);
nor U3905 (N_3905,N_2798,N_2907);
nor U3906 (N_3906,N_2541,N_2995);
and U3907 (N_3907,N_2614,N_2867);
nand U3908 (N_3908,N_2236,N_2735);
or U3909 (N_3909,N_2905,N_2020);
or U3910 (N_3910,N_2762,N_2245);
or U3911 (N_3911,N_2578,N_2522);
or U3912 (N_3912,N_2569,N_2523);
and U3913 (N_3913,N_2138,N_2967);
or U3914 (N_3914,N_2997,N_2961);
xor U3915 (N_3915,N_2447,N_2759);
xor U3916 (N_3916,N_2359,N_2889);
xnor U3917 (N_3917,N_2877,N_2249);
nand U3918 (N_3918,N_2912,N_2949);
xnor U3919 (N_3919,N_2469,N_2265);
nor U3920 (N_3920,N_2617,N_2163);
nor U3921 (N_3921,N_2702,N_2467);
or U3922 (N_3922,N_2581,N_2437);
nand U3923 (N_3923,N_2313,N_2447);
xor U3924 (N_3924,N_2701,N_2400);
xnor U3925 (N_3925,N_2800,N_2610);
and U3926 (N_3926,N_2373,N_2742);
nand U3927 (N_3927,N_2508,N_2426);
and U3928 (N_3928,N_2208,N_2212);
and U3929 (N_3929,N_2912,N_2515);
nand U3930 (N_3930,N_2175,N_2908);
nor U3931 (N_3931,N_2517,N_2574);
xor U3932 (N_3932,N_2111,N_2986);
or U3933 (N_3933,N_2089,N_2650);
xor U3934 (N_3934,N_2708,N_2291);
nor U3935 (N_3935,N_2525,N_2973);
nor U3936 (N_3936,N_2903,N_2637);
xor U3937 (N_3937,N_2926,N_2242);
nor U3938 (N_3938,N_2256,N_2236);
nand U3939 (N_3939,N_2194,N_2080);
xor U3940 (N_3940,N_2792,N_2655);
nor U3941 (N_3941,N_2416,N_2002);
nand U3942 (N_3942,N_2235,N_2751);
or U3943 (N_3943,N_2490,N_2671);
nor U3944 (N_3944,N_2281,N_2511);
nand U3945 (N_3945,N_2363,N_2913);
and U3946 (N_3946,N_2239,N_2748);
nand U3947 (N_3947,N_2176,N_2193);
or U3948 (N_3948,N_2221,N_2049);
xor U3949 (N_3949,N_2065,N_2244);
or U3950 (N_3950,N_2814,N_2664);
xnor U3951 (N_3951,N_2848,N_2829);
xnor U3952 (N_3952,N_2948,N_2420);
nand U3953 (N_3953,N_2686,N_2785);
nand U3954 (N_3954,N_2268,N_2135);
nor U3955 (N_3955,N_2932,N_2479);
and U3956 (N_3956,N_2439,N_2247);
nand U3957 (N_3957,N_2849,N_2334);
or U3958 (N_3958,N_2903,N_2748);
nor U3959 (N_3959,N_2753,N_2370);
or U3960 (N_3960,N_2557,N_2062);
xnor U3961 (N_3961,N_2900,N_2401);
nand U3962 (N_3962,N_2950,N_2000);
nor U3963 (N_3963,N_2724,N_2557);
xor U3964 (N_3964,N_2209,N_2661);
xnor U3965 (N_3965,N_2177,N_2019);
xor U3966 (N_3966,N_2344,N_2963);
nor U3967 (N_3967,N_2866,N_2853);
or U3968 (N_3968,N_2871,N_2850);
and U3969 (N_3969,N_2901,N_2696);
nand U3970 (N_3970,N_2948,N_2813);
or U3971 (N_3971,N_2657,N_2820);
nand U3972 (N_3972,N_2477,N_2204);
xnor U3973 (N_3973,N_2493,N_2700);
or U3974 (N_3974,N_2761,N_2251);
and U3975 (N_3975,N_2927,N_2450);
and U3976 (N_3976,N_2479,N_2514);
nor U3977 (N_3977,N_2563,N_2339);
and U3978 (N_3978,N_2442,N_2902);
xnor U3979 (N_3979,N_2607,N_2133);
xnor U3980 (N_3980,N_2565,N_2802);
or U3981 (N_3981,N_2303,N_2962);
nor U3982 (N_3982,N_2363,N_2492);
xor U3983 (N_3983,N_2938,N_2222);
xnor U3984 (N_3984,N_2054,N_2228);
nor U3985 (N_3985,N_2092,N_2161);
or U3986 (N_3986,N_2463,N_2166);
nand U3987 (N_3987,N_2922,N_2310);
xnor U3988 (N_3988,N_2748,N_2039);
nor U3989 (N_3989,N_2723,N_2984);
and U3990 (N_3990,N_2442,N_2192);
nand U3991 (N_3991,N_2197,N_2650);
and U3992 (N_3992,N_2950,N_2572);
nand U3993 (N_3993,N_2622,N_2991);
and U3994 (N_3994,N_2525,N_2020);
or U3995 (N_3995,N_2773,N_2559);
nand U3996 (N_3996,N_2000,N_2294);
nand U3997 (N_3997,N_2397,N_2310);
nor U3998 (N_3998,N_2263,N_2157);
xor U3999 (N_3999,N_2340,N_2446);
nand U4000 (N_4000,N_3012,N_3923);
nand U4001 (N_4001,N_3645,N_3649);
nor U4002 (N_4002,N_3078,N_3793);
nor U4003 (N_4003,N_3032,N_3456);
or U4004 (N_4004,N_3668,N_3701);
nor U4005 (N_4005,N_3410,N_3756);
and U4006 (N_4006,N_3089,N_3884);
and U4007 (N_4007,N_3841,N_3204);
xor U4008 (N_4008,N_3058,N_3936);
nand U4009 (N_4009,N_3026,N_3974);
and U4010 (N_4010,N_3972,N_3886);
nor U4011 (N_4011,N_3951,N_3201);
nand U4012 (N_4012,N_3132,N_3134);
or U4013 (N_4013,N_3270,N_3890);
or U4014 (N_4014,N_3784,N_3937);
nand U4015 (N_4015,N_3573,N_3938);
nand U4016 (N_4016,N_3583,N_3188);
nand U4017 (N_4017,N_3397,N_3712);
and U4018 (N_4018,N_3006,N_3077);
nand U4019 (N_4019,N_3084,N_3116);
nand U4020 (N_4020,N_3344,N_3167);
and U4021 (N_4021,N_3297,N_3404);
or U4022 (N_4022,N_3355,N_3378);
xor U4023 (N_4023,N_3422,N_3342);
or U4024 (N_4024,N_3955,N_3045);
nand U4025 (N_4025,N_3778,N_3950);
and U4026 (N_4026,N_3284,N_3449);
xor U4027 (N_4027,N_3105,N_3265);
nand U4028 (N_4028,N_3008,N_3389);
nor U4029 (N_4029,N_3692,N_3716);
nand U4030 (N_4030,N_3862,N_3585);
or U4031 (N_4031,N_3138,N_3211);
xor U4032 (N_4032,N_3027,N_3803);
nand U4033 (N_4033,N_3327,N_3602);
nand U4034 (N_4034,N_3703,N_3436);
nand U4035 (N_4035,N_3306,N_3907);
nand U4036 (N_4036,N_3213,N_3177);
nand U4037 (N_4037,N_3964,N_3372);
nand U4038 (N_4038,N_3751,N_3215);
or U4039 (N_4039,N_3471,N_3905);
nand U4040 (N_4040,N_3067,N_3179);
nor U4041 (N_4041,N_3894,N_3816);
xnor U4042 (N_4042,N_3450,N_3021);
nand U4043 (N_4043,N_3652,N_3486);
and U4044 (N_4044,N_3693,N_3352);
and U4045 (N_4045,N_3070,N_3186);
nor U4046 (N_4046,N_3853,N_3590);
nor U4047 (N_4047,N_3060,N_3570);
nor U4048 (N_4048,N_3219,N_3588);
nand U4049 (N_4049,N_3965,N_3453);
or U4050 (N_4050,N_3738,N_3343);
nand U4051 (N_4051,N_3603,N_3085);
xnor U4052 (N_4052,N_3561,N_3673);
xor U4053 (N_4053,N_3596,N_3749);
nand U4054 (N_4054,N_3128,N_3662);
nand U4055 (N_4055,N_3592,N_3648);
nor U4056 (N_4056,N_3051,N_3987);
and U4057 (N_4057,N_3903,N_3710);
nand U4058 (N_4058,N_3249,N_3996);
nor U4059 (N_4059,N_3586,N_3001);
or U4060 (N_4060,N_3605,N_3216);
nor U4061 (N_4061,N_3178,N_3010);
or U4062 (N_4062,N_3727,N_3137);
or U4063 (N_4063,N_3121,N_3148);
nand U4064 (N_4064,N_3665,N_3824);
and U4065 (N_4065,N_3607,N_3124);
xor U4066 (N_4066,N_3229,N_3799);
nand U4067 (N_4067,N_3904,N_3455);
or U4068 (N_4068,N_3960,N_3830);
xor U4069 (N_4069,N_3019,N_3809);
nand U4070 (N_4070,N_3625,N_3767);
nor U4071 (N_4071,N_3675,N_3777);
nand U4072 (N_4072,N_3879,N_3090);
nor U4073 (N_4073,N_3258,N_3944);
or U4074 (N_4074,N_3567,N_3413);
or U4075 (N_4075,N_3971,N_3543);
or U4076 (N_4076,N_3104,N_3736);
or U4077 (N_4077,N_3677,N_3542);
xor U4078 (N_4078,N_3446,N_3826);
xnor U4079 (N_4079,N_3264,N_3755);
or U4080 (N_4080,N_3250,N_3334);
and U4081 (N_4081,N_3241,N_3516);
or U4082 (N_4082,N_3139,N_3745);
and U4083 (N_4083,N_3472,N_3156);
and U4084 (N_4084,N_3521,N_3792);
nand U4085 (N_4085,N_3383,N_3339);
xnor U4086 (N_4086,N_3257,N_3035);
nand U4087 (N_4087,N_3639,N_3055);
or U4088 (N_4088,N_3240,N_3642);
nor U4089 (N_4089,N_3071,N_3052);
nand U4090 (N_4090,N_3034,N_3844);
and U4091 (N_4091,N_3761,N_3544);
nand U4092 (N_4092,N_3330,N_3308);
or U4093 (N_4093,N_3949,N_3096);
and U4094 (N_4094,N_3406,N_3108);
and U4095 (N_4095,N_3385,N_3395);
or U4096 (N_4096,N_3735,N_3539);
nand U4097 (N_4097,N_3806,N_3222);
nand U4098 (N_4098,N_3817,N_3847);
xnor U4099 (N_4099,N_3838,N_3787);
and U4100 (N_4100,N_3380,N_3910);
and U4101 (N_4101,N_3582,N_3225);
and U4102 (N_4102,N_3367,N_3564);
nor U4103 (N_4103,N_3985,N_3202);
nand U4104 (N_4104,N_3261,N_3888);
and U4105 (N_4105,N_3260,N_3644);
nor U4106 (N_4106,N_3968,N_3811);
and U4107 (N_4107,N_3580,N_3037);
or U4108 (N_4108,N_3362,N_3289);
xor U4109 (N_4109,N_3454,N_3946);
or U4110 (N_4110,N_3109,N_3232);
xor U4111 (N_4111,N_3236,N_3114);
xor U4112 (N_4112,N_3520,N_3502);
nand U4113 (N_4113,N_3214,N_3717);
xor U4114 (N_4114,N_3152,N_3758);
nor U4115 (N_4115,N_3220,N_3402);
or U4116 (N_4116,N_3933,N_3233);
nor U4117 (N_4117,N_3237,N_3640);
xor U4118 (N_4118,N_3063,N_3865);
or U4119 (N_4119,N_3018,N_3895);
and U4120 (N_4120,N_3919,N_3613);
or U4121 (N_4121,N_3863,N_3628);
xor U4122 (N_4122,N_3978,N_3254);
xor U4123 (N_4123,N_3111,N_3812);
nand U4124 (N_4124,N_3650,N_3932);
xor U4125 (N_4125,N_3617,N_3655);
xor U4126 (N_4126,N_3268,N_3195);
xnor U4127 (N_4127,N_3427,N_3529);
or U4128 (N_4128,N_3540,N_3118);
and U4129 (N_4129,N_3506,N_3780);
and U4130 (N_4130,N_3206,N_3331);
and U4131 (N_4131,N_3341,N_3381);
nand U4132 (N_4132,N_3474,N_3072);
nor U4133 (N_4133,N_3880,N_3878);
nor U4134 (N_4134,N_3493,N_3347);
or U4135 (N_4135,N_3171,N_3252);
nor U4136 (N_4136,N_3468,N_3476);
nand U4137 (N_4137,N_3351,N_3439);
nor U4138 (N_4138,N_3646,N_3141);
or U4139 (N_4139,N_3255,N_3672);
and U4140 (N_4140,N_3414,N_3050);
and U4141 (N_4141,N_3804,N_3666);
nand U4142 (N_4142,N_3015,N_3357);
xor U4143 (N_4143,N_3688,N_3835);
nor U4144 (N_4144,N_3365,N_3979);
and U4145 (N_4145,N_3747,N_3958);
and U4146 (N_4146,N_3193,N_3901);
or U4147 (N_4147,N_3143,N_3684);
nor U4148 (N_4148,N_3740,N_3431);
nand U4149 (N_4149,N_3752,N_3320);
xor U4150 (N_4150,N_3388,N_3300);
or U4151 (N_4151,N_3718,N_3970);
and U4152 (N_4152,N_3401,N_3842);
or U4153 (N_4153,N_3638,N_3952);
and U4154 (N_4154,N_3151,N_3384);
nor U4155 (N_4155,N_3174,N_3783);
and U4156 (N_4156,N_3595,N_3527);
nor U4157 (N_4157,N_3925,N_3897);
nand U4158 (N_4158,N_3463,N_3366);
and U4159 (N_4159,N_3855,N_3130);
nand U4160 (N_4160,N_3360,N_3230);
nor U4161 (N_4161,N_3243,N_3510);
or U4162 (N_4162,N_3656,N_3739);
and U4163 (N_4163,N_3391,N_3191);
xnor U4164 (N_4164,N_3073,N_3429);
nand U4165 (N_4165,N_3094,N_3545);
nand U4166 (N_4166,N_3658,N_3262);
xnor U4167 (N_4167,N_3864,N_3800);
nor U4168 (N_4168,N_3851,N_3190);
nand U4169 (N_4169,N_3930,N_3281);
or U4170 (N_4170,N_3578,N_3408);
or U4171 (N_4171,N_3368,N_3575);
xnor U4172 (N_4172,N_3212,N_3166);
nor U4173 (N_4173,N_3560,N_3228);
xor U4174 (N_4174,N_3871,N_3869);
xor U4175 (N_4175,N_3843,N_3850);
or U4176 (N_4176,N_3197,N_3538);
and U4177 (N_4177,N_3957,N_3962);
or U4178 (N_4178,N_3092,N_3305);
and U4179 (N_4179,N_3523,N_3664);
nand U4180 (N_4180,N_3594,N_3165);
and U4181 (N_4181,N_3282,N_3119);
nand U4182 (N_4182,N_3597,N_3392);
nand U4183 (N_4183,N_3379,N_3122);
nand U4184 (N_4184,N_3318,N_3273);
or U4185 (N_4185,N_3068,N_3789);
and U4186 (N_4186,N_3013,N_3867);
or U4187 (N_4187,N_3834,N_3891);
or U4188 (N_4188,N_3786,N_3988);
and U4189 (N_4189,N_3428,N_3437);
or U4190 (N_4190,N_3478,N_3140);
and U4191 (N_4191,N_3609,N_3481);
and U4192 (N_4192,N_3568,N_3671);
or U4193 (N_4193,N_3555,N_3981);
or U4194 (N_4194,N_3200,N_3432);
and U4195 (N_4195,N_3998,N_3292);
nor U4196 (N_4196,N_3822,N_3420);
xor U4197 (N_4197,N_3490,N_3993);
xnor U4198 (N_4198,N_3153,N_3390);
nand U4199 (N_4199,N_3421,N_3795);
and U4200 (N_4200,N_3698,N_3947);
or U4201 (N_4201,N_3661,N_3541);
or U4202 (N_4202,N_3043,N_3031);
or U4203 (N_4203,N_3857,N_3976);
and U4204 (N_4204,N_3505,N_3659);
or U4205 (N_4205,N_3808,N_3694);
and U4206 (N_4206,N_3967,N_3517);
nand U4207 (N_4207,N_3883,N_3393);
nor U4208 (N_4208,N_3742,N_3566);
and U4209 (N_4209,N_3537,N_3346);
or U4210 (N_4210,N_3107,N_3364);
nor U4211 (N_4211,N_3906,N_3088);
nor U4212 (N_4212,N_3409,N_3820);
and U4213 (N_4213,N_3093,N_3504);
nor U4214 (N_4214,N_3374,N_3482);
xor U4215 (N_4215,N_3163,N_3730);
nor U4216 (N_4216,N_3791,N_3160);
or U4217 (N_4217,N_3172,N_3417);
xnor U4218 (N_4218,N_3917,N_3158);
and U4219 (N_4219,N_3556,N_3729);
xor U4220 (N_4220,N_3584,N_3775);
or U4221 (N_4221,N_3059,N_3721);
and U4222 (N_4222,N_3227,N_3324);
nand U4223 (N_4223,N_3732,N_3685);
xnor U4224 (N_4224,N_3161,N_3245);
or U4225 (N_4225,N_3833,N_3038);
nand U4226 (N_4226,N_3303,N_3579);
nand U4227 (N_4227,N_3036,N_3087);
nor U4228 (N_4228,N_3915,N_3501);
nand U4229 (N_4229,N_3435,N_3312);
xor U4230 (N_4230,N_3647,N_3902);
and U4231 (N_4231,N_3748,N_3768);
or U4232 (N_4232,N_3176,N_3136);
xnor U4233 (N_4233,N_3479,N_3709);
nor U4234 (N_4234,N_3494,N_3358);
xnor U4235 (N_4235,N_3011,N_3242);
nand U4236 (N_4236,N_3610,N_3608);
xor U4237 (N_4237,N_3304,N_3440);
nand U4238 (N_4238,N_3674,N_3489);
nor U4239 (N_4239,N_3335,N_3969);
nor U4240 (N_4240,N_3881,N_3899);
xor U4241 (N_4241,N_3928,N_3198);
and U4242 (N_4242,N_3629,N_3029);
nor U4243 (N_4243,N_3612,N_3005);
xor U4244 (N_4244,N_3587,N_3144);
and U4245 (N_4245,N_3689,N_3291);
xor U4246 (N_4246,N_3407,N_3209);
or U4247 (N_4247,N_3491,N_3434);
nor U4248 (N_4248,N_3248,N_3877);
or U4249 (N_4249,N_3983,N_3829);
nor U4250 (N_4250,N_3123,N_3375);
nand U4251 (N_4251,N_3512,N_3507);
or U4252 (N_4252,N_3218,N_3086);
nor U4253 (N_4253,N_3553,N_3091);
nor U4254 (N_4254,N_3794,N_3256);
nand U4255 (N_4255,N_3999,N_3276);
nand U4256 (N_4256,N_3142,N_3991);
nor U4257 (N_4257,N_3591,N_3196);
nand U4258 (N_4258,N_3790,N_3492);
nor U4259 (N_4259,N_3513,N_3657);
nand U4260 (N_4260,N_3854,N_3889);
nand U4261 (N_4261,N_3102,N_3117);
nor U4262 (N_4262,N_3048,N_3623);
or U4263 (N_4263,N_3317,N_3173);
or U4264 (N_4264,N_3531,N_3313);
and U4265 (N_4265,N_3253,N_3425);
and U4266 (N_4266,N_3737,N_3430);
or U4267 (N_4267,N_3461,N_3373);
and U4268 (N_4268,N_3619,N_3080);
or U4269 (N_4269,N_3876,N_3338);
nand U4270 (N_4270,N_3547,N_3667);
nand U4271 (N_4271,N_3269,N_3574);
nand U4272 (N_4272,N_3785,N_3340);
nor U4273 (N_4273,N_3187,N_3175);
or U4274 (N_4274,N_3700,N_3075);
nor U4275 (N_4275,N_3849,N_3945);
xor U4276 (N_4276,N_3887,N_3133);
or U4277 (N_4277,N_3975,N_3781);
and U4278 (N_4278,N_3299,N_3146);
or U4279 (N_4279,N_3845,N_3707);
nand U4280 (N_4280,N_3852,N_3097);
or U4281 (N_4281,N_3654,N_3741);
nand U4282 (N_4282,N_3286,N_3120);
or U4283 (N_4283,N_3959,N_3444);
or U4284 (N_4284,N_3182,N_3274);
and U4285 (N_4285,N_3495,N_3589);
xnor U4286 (N_4286,N_3802,N_3563);
nor U4287 (N_4287,N_3251,N_3115);
nor U4288 (N_4288,N_3924,N_3247);
and U4289 (N_4289,N_3469,N_3065);
or U4290 (N_4290,N_3020,N_3484);
xnor U4291 (N_4291,N_3451,N_3480);
and U4292 (N_4292,N_3931,N_3095);
nand U4293 (N_4293,N_3956,N_3558);
xnor U4294 (N_4294,N_3690,N_3832);
nor U4295 (N_4295,N_3713,N_3641);
or U4296 (N_4296,N_3315,N_3942);
and U4297 (N_4297,N_3294,N_3418);
nand U4298 (N_4298,N_3874,N_3181);
and U4299 (N_4299,N_3234,N_3620);
nand U4300 (N_4300,N_3714,N_3776);
and U4301 (N_4301,N_3016,N_3990);
and U4302 (N_4302,N_3370,N_3731);
nand U4303 (N_4303,N_3686,N_3488);
and U4304 (N_4304,N_3125,N_3840);
xnor U4305 (N_4305,N_3056,N_3861);
xor U4306 (N_4306,N_3185,N_3473);
nor U4307 (N_4307,N_3680,N_3514);
nor U4308 (N_4308,N_3278,N_3509);
nand U4309 (N_4309,N_3550,N_3669);
nand U4310 (N_4310,N_3183,N_3994);
or U4311 (N_4311,N_3235,N_3162);
and U4312 (N_4312,N_3475,N_3135);
and U4313 (N_4313,N_3022,N_3062);
and U4314 (N_4314,N_3356,N_3462);
nand U4315 (N_4315,N_3546,N_3929);
nand U4316 (N_4316,N_3989,N_3064);
nand U4317 (N_4317,N_3192,N_3394);
and U4318 (N_4318,N_3918,N_3728);
and U4319 (N_4319,N_3184,N_3061);
nand U4320 (N_4320,N_3326,N_3023);
nand U4321 (N_4321,N_3565,N_3239);
nor U4322 (N_4322,N_3810,N_3333);
or U4323 (N_4323,N_3601,N_3042);
and U4324 (N_4324,N_3131,N_3290);
xor U4325 (N_4325,N_3155,N_3773);
nand U4326 (N_4326,N_3287,N_3328);
and U4327 (N_4327,N_3637,N_3499);
and U4328 (N_4328,N_3189,N_3017);
nand U4329 (N_4329,N_3599,N_3549);
and U4330 (N_4330,N_3321,N_3726);
xor U4331 (N_4331,N_3986,N_3708);
nor U4332 (N_4332,N_3244,N_3277);
nand U4333 (N_4333,N_3581,N_3870);
nand U4334 (N_4334,N_3154,N_3839);
and U4335 (N_4335,N_3415,N_3129);
xnor U4336 (N_4336,N_3697,N_3298);
and U4337 (N_4337,N_3359,N_3757);
nand U4338 (N_4338,N_3280,N_3720);
or U4339 (N_4339,N_3653,N_3103);
nor U4340 (N_4340,N_3875,N_3487);
nor U4341 (N_4341,N_3569,N_3283);
nand U4342 (N_4342,N_3866,N_3076);
and U4343 (N_4343,N_3515,N_3528);
nand U4344 (N_4344,N_3912,N_3846);
nand U4345 (N_4345,N_3632,N_3961);
nand U4346 (N_4346,N_3054,N_3765);
nand U4347 (N_4347,N_3069,N_3941);
and U4348 (N_4348,N_3412,N_3293);
nand U4349 (N_4349,N_3459,N_3746);
nor U4350 (N_4350,N_3231,N_3705);
nand U4351 (N_4351,N_3725,N_3633);
nand U4352 (N_4352,N_3796,N_3426);
nand U4353 (N_4353,N_3263,N_3606);
nand U4354 (N_4354,N_3940,N_3369);
or U4355 (N_4355,N_3953,N_3033);
and U4356 (N_4356,N_3896,N_3980);
nor U4357 (N_4357,N_3503,N_3150);
nor U4358 (N_4358,N_3691,N_3470);
nand U4359 (N_4359,N_3467,N_3621);
xor U4360 (N_4360,N_3309,N_3868);
nor U4361 (N_4361,N_3438,N_3788);
and U4362 (N_4362,N_3643,N_3681);
and U4363 (N_4363,N_3682,N_3534);
and U4364 (N_4364,N_3763,N_3966);
nor U4365 (N_4365,N_3577,N_3423);
or U4366 (N_4366,N_3948,N_3525);
xnor U4367 (N_4367,N_3651,N_3954);
or U4368 (N_4368,N_3719,N_3836);
nand U4369 (N_4369,N_3624,N_3224);
nor U4370 (N_4370,N_3079,N_3464);
or U4371 (N_4371,N_3296,N_3660);
nand U4372 (N_4372,N_3801,N_3205);
or U4373 (N_4373,N_3618,N_3458);
and U4374 (N_4374,N_3272,N_3530);
xnor U4375 (N_4375,N_3002,N_3722);
nand U4376 (N_4376,N_3419,N_3935);
and U4377 (N_4377,N_3635,N_3535);
nor U4378 (N_4378,N_3110,N_3814);
nor U4379 (N_4379,N_3246,N_3337);
and U4380 (N_4380,N_3083,N_3350);
and U4381 (N_4381,N_3101,N_3518);
nand U4382 (N_4382,N_3387,N_3536);
xor U4383 (N_4383,N_3199,N_3047);
nor U4384 (N_4384,N_3927,N_3611);
and U4385 (N_4385,N_3500,N_3798);
and U4386 (N_4386,N_3302,N_3074);
nor U4387 (N_4387,N_3433,N_3319);
and U4388 (N_4388,N_3267,N_3552);
nor U4389 (N_4389,N_3771,N_3898);
nand U4390 (N_4390,N_3279,N_3670);
and U4391 (N_4391,N_3403,N_3551);
and U4392 (N_4392,N_3443,N_3399);
or U4393 (N_4393,N_3100,N_3711);
nor U4394 (N_4394,N_3992,N_3485);
nor U4395 (N_4395,N_3593,N_3828);
xnor U4396 (N_4396,N_3963,N_3872);
xor U4397 (N_4397,N_3003,N_3926);
and U4398 (N_4398,N_3893,N_3572);
nand U4399 (N_4399,N_3465,N_3098);
nand U4400 (N_4400,N_3081,N_3702);
and U4401 (N_4401,N_3024,N_3914);
nor U4402 (N_4402,N_3683,N_3827);
or U4403 (N_4403,N_3149,N_3025);
and U4404 (N_4404,N_3044,N_3977);
xnor U4405 (N_4405,N_3511,N_3445);
xor U4406 (N_4406,N_3679,N_3706);
nor U4407 (N_4407,N_3626,N_3754);
nor U4408 (N_4408,N_3532,N_3028);
or U4409 (N_4409,N_3049,N_3921);
nor U4410 (N_4410,N_3571,N_3604);
nor U4411 (N_4411,N_3180,N_3909);
and U4412 (N_4412,N_3557,N_3769);
nor U4413 (N_4413,N_3782,N_3271);
or U4414 (N_4414,N_3634,N_3457);
xor U4415 (N_4415,N_3398,N_3554);
or U4416 (N_4416,N_3424,N_3477);
nor U4417 (N_4417,N_3934,N_3126);
and U4418 (N_4418,N_3325,N_3900);
or U4419 (N_4419,N_3396,N_3329);
or U4420 (N_4420,N_3562,N_3112);
nand U4421 (N_4421,N_3805,N_3837);
xor U4422 (N_4422,N_3039,N_3377);
nor U4423 (N_4423,N_3524,N_3483);
or U4424 (N_4424,N_3452,N_3759);
or U4425 (N_4425,N_3715,N_3772);
or U4426 (N_4426,N_3519,N_3332);
or U4427 (N_4427,N_3275,N_3818);
or U4428 (N_4428,N_3223,N_3695);
and U4429 (N_4429,N_3363,N_3295);
nand U4430 (N_4430,N_3676,N_3466);
nand U4431 (N_4431,N_3939,N_3526);
or U4432 (N_4432,N_3442,N_3856);
or U4433 (N_4433,N_3997,N_3724);
and U4434 (N_4434,N_3170,N_3882);
or U4435 (N_4435,N_3386,N_3766);
or U4436 (N_4436,N_3311,N_3441);
xor U4437 (N_4437,N_3920,N_3014);
or U4438 (N_4438,N_3371,N_3885);
xor U4439 (N_4439,N_3663,N_3508);
and U4440 (N_4440,N_3807,N_3743);
nand U4441 (N_4441,N_3723,N_3522);
or U4442 (N_4442,N_3687,N_3908);
and U4443 (N_4443,N_3345,N_3744);
or U4444 (N_4444,N_3113,N_3226);
xor U4445 (N_4445,N_3873,N_3825);
or U4446 (N_4446,N_3310,N_3943);
nor U4447 (N_4447,N_3911,N_3400);
and U4448 (N_4448,N_3217,N_3498);
nor U4449 (N_4449,N_3349,N_3627);
xor U4450 (N_4450,N_3622,N_3460);
xnor U4451 (N_4451,N_3099,N_3982);
or U4452 (N_4452,N_3040,N_3760);
nor U4453 (N_4453,N_3066,N_3823);
or U4454 (N_4454,N_3616,N_3764);
xnor U4455 (N_4455,N_3405,N_3009);
and U4456 (N_4456,N_3448,N_3630);
nand U4457 (N_4457,N_3314,N_3208);
nor U4458 (N_4458,N_3750,N_3753);
nor U4459 (N_4459,N_3147,N_3770);
xnor U4460 (N_4460,N_3984,N_3210);
nand U4461 (N_4461,N_3615,N_3636);
or U4462 (N_4462,N_3007,N_3382);
xor U4463 (N_4463,N_3678,N_3819);
nand U4464 (N_4464,N_3361,N_3922);
xnor U4465 (N_4465,N_3533,N_3779);
or U4466 (N_4466,N_3266,N_3916);
xor U4467 (N_4467,N_3041,N_3631);
or U4468 (N_4468,N_3157,N_3762);
or U4469 (N_4469,N_3733,N_3598);
or U4470 (N_4470,N_3813,N_3348);
and U4471 (N_4471,N_3548,N_3030);
xor U4472 (N_4472,N_3576,N_3559);
nor U4473 (N_4473,N_3203,N_3336);
xnor U4474 (N_4474,N_3285,N_3316);
and U4475 (N_4475,N_3164,N_3995);
nor U4476 (N_4476,N_3145,N_3973);
nor U4477 (N_4477,N_3696,N_3057);
nor U4478 (N_4478,N_3704,N_3322);
xor U4479 (N_4479,N_3238,N_3082);
and U4480 (N_4480,N_3734,N_3821);
or U4481 (N_4481,N_3600,N_3323);
and U4482 (N_4482,N_3699,N_3411);
and U4483 (N_4483,N_3447,N_3000);
nor U4484 (N_4484,N_3354,N_3858);
xnor U4485 (N_4485,N_3797,N_3860);
xor U4486 (N_4486,N_3416,N_3376);
and U4487 (N_4487,N_3831,N_3207);
and U4488 (N_4488,N_3159,N_3046);
and U4489 (N_4489,N_3774,N_3288);
xor U4490 (N_4490,N_3127,N_3106);
nor U4491 (N_4491,N_3307,N_3859);
and U4492 (N_4492,N_3004,N_3497);
nand U4493 (N_4493,N_3848,N_3194);
nand U4494 (N_4494,N_3892,N_3496);
or U4495 (N_4495,N_3614,N_3353);
nor U4496 (N_4496,N_3221,N_3913);
xnor U4497 (N_4497,N_3259,N_3168);
nand U4498 (N_4498,N_3053,N_3301);
xor U4499 (N_4499,N_3815,N_3169);
and U4500 (N_4500,N_3660,N_3550);
nor U4501 (N_4501,N_3035,N_3102);
nand U4502 (N_4502,N_3694,N_3380);
nand U4503 (N_4503,N_3070,N_3767);
and U4504 (N_4504,N_3341,N_3147);
nor U4505 (N_4505,N_3211,N_3087);
or U4506 (N_4506,N_3658,N_3195);
nand U4507 (N_4507,N_3773,N_3839);
nor U4508 (N_4508,N_3961,N_3605);
nand U4509 (N_4509,N_3350,N_3556);
xnor U4510 (N_4510,N_3347,N_3668);
nor U4511 (N_4511,N_3636,N_3684);
nor U4512 (N_4512,N_3126,N_3167);
nand U4513 (N_4513,N_3088,N_3180);
or U4514 (N_4514,N_3426,N_3105);
xnor U4515 (N_4515,N_3219,N_3001);
nand U4516 (N_4516,N_3024,N_3097);
or U4517 (N_4517,N_3059,N_3742);
or U4518 (N_4518,N_3409,N_3711);
nor U4519 (N_4519,N_3144,N_3523);
xor U4520 (N_4520,N_3085,N_3807);
nor U4521 (N_4521,N_3489,N_3095);
nor U4522 (N_4522,N_3434,N_3667);
nor U4523 (N_4523,N_3132,N_3550);
nor U4524 (N_4524,N_3843,N_3301);
or U4525 (N_4525,N_3367,N_3099);
nand U4526 (N_4526,N_3729,N_3915);
nor U4527 (N_4527,N_3279,N_3693);
or U4528 (N_4528,N_3702,N_3602);
nand U4529 (N_4529,N_3668,N_3609);
and U4530 (N_4530,N_3603,N_3568);
and U4531 (N_4531,N_3309,N_3079);
or U4532 (N_4532,N_3934,N_3424);
or U4533 (N_4533,N_3178,N_3298);
xnor U4534 (N_4534,N_3364,N_3337);
xnor U4535 (N_4535,N_3084,N_3732);
nand U4536 (N_4536,N_3217,N_3831);
xnor U4537 (N_4537,N_3547,N_3563);
and U4538 (N_4538,N_3426,N_3549);
and U4539 (N_4539,N_3243,N_3263);
or U4540 (N_4540,N_3322,N_3376);
xnor U4541 (N_4541,N_3628,N_3459);
nor U4542 (N_4542,N_3393,N_3816);
and U4543 (N_4543,N_3546,N_3346);
nand U4544 (N_4544,N_3179,N_3427);
and U4545 (N_4545,N_3746,N_3165);
nand U4546 (N_4546,N_3317,N_3275);
or U4547 (N_4547,N_3748,N_3824);
and U4548 (N_4548,N_3721,N_3225);
xor U4549 (N_4549,N_3228,N_3819);
and U4550 (N_4550,N_3926,N_3930);
or U4551 (N_4551,N_3166,N_3695);
or U4552 (N_4552,N_3645,N_3243);
nand U4553 (N_4553,N_3887,N_3402);
or U4554 (N_4554,N_3321,N_3072);
or U4555 (N_4555,N_3371,N_3188);
and U4556 (N_4556,N_3440,N_3705);
or U4557 (N_4557,N_3696,N_3591);
xnor U4558 (N_4558,N_3767,N_3910);
nor U4559 (N_4559,N_3930,N_3839);
or U4560 (N_4560,N_3820,N_3100);
or U4561 (N_4561,N_3675,N_3438);
or U4562 (N_4562,N_3845,N_3474);
nand U4563 (N_4563,N_3997,N_3466);
nor U4564 (N_4564,N_3968,N_3204);
and U4565 (N_4565,N_3509,N_3430);
xor U4566 (N_4566,N_3439,N_3919);
and U4567 (N_4567,N_3559,N_3880);
or U4568 (N_4568,N_3296,N_3580);
or U4569 (N_4569,N_3160,N_3782);
nor U4570 (N_4570,N_3130,N_3362);
nand U4571 (N_4571,N_3542,N_3300);
or U4572 (N_4572,N_3325,N_3947);
or U4573 (N_4573,N_3817,N_3652);
xnor U4574 (N_4574,N_3570,N_3421);
xor U4575 (N_4575,N_3634,N_3249);
xnor U4576 (N_4576,N_3737,N_3275);
nor U4577 (N_4577,N_3611,N_3732);
xnor U4578 (N_4578,N_3059,N_3403);
nor U4579 (N_4579,N_3996,N_3311);
nand U4580 (N_4580,N_3553,N_3738);
xnor U4581 (N_4581,N_3831,N_3295);
xnor U4582 (N_4582,N_3157,N_3326);
nand U4583 (N_4583,N_3460,N_3062);
and U4584 (N_4584,N_3833,N_3044);
nand U4585 (N_4585,N_3517,N_3820);
nor U4586 (N_4586,N_3830,N_3520);
and U4587 (N_4587,N_3616,N_3410);
and U4588 (N_4588,N_3272,N_3270);
nand U4589 (N_4589,N_3642,N_3629);
and U4590 (N_4590,N_3219,N_3623);
or U4591 (N_4591,N_3184,N_3010);
and U4592 (N_4592,N_3708,N_3042);
or U4593 (N_4593,N_3444,N_3353);
nor U4594 (N_4594,N_3844,N_3872);
and U4595 (N_4595,N_3596,N_3857);
nand U4596 (N_4596,N_3947,N_3597);
or U4597 (N_4597,N_3603,N_3675);
nor U4598 (N_4598,N_3892,N_3025);
nor U4599 (N_4599,N_3510,N_3891);
xnor U4600 (N_4600,N_3828,N_3596);
nor U4601 (N_4601,N_3227,N_3966);
nor U4602 (N_4602,N_3612,N_3400);
or U4603 (N_4603,N_3728,N_3388);
or U4604 (N_4604,N_3080,N_3284);
nand U4605 (N_4605,N_3981,N_3287);
nand U4606 (N_4606,N_3428,N_3268);
or U4607 (N_4607,N_3449,N_3243);
nor U4608 (N_4608,N_3550,N_3069);
or U4609 (N_4609,N_3202,N_3236);
nand U4610 (N_4610,N_3760,N_3736);
or U4611 (N_4611,N_3113,N_3027);
or U4612 (N_4612,N_3802,N_3794);
xor U4613 (N_4613,N_3299,N_3761);
or U4614 (N_4614,N_3813,N_3589);
nand U4615 (N_4615,N_3162,N_3051);
nor U4616 (N_4616,N_3058,N_3444);
nand U4617 (N_4617,N_3058,N_3012);
nand U4618 (N_4618,N_3878,N_3959);
nor U4619 (N_4619,N_3807,N_3689);
xor U4620 (N_4620,N_3524,N_3875);
xnor U4621 (N_4621,N_3547,N_3662);
and U4622 (N_4622,N_3985,N_3105);
nand U4623 (N_4623,N_3703,N_3641);
xor U4624 (N_4624,N_3211,N_3862);
nor U4625 (N_4625,N_3034,N_3662);
nand U4626 (N_4626,N_3346,N_3463);
nor U4627 (N_4627,N_3418,N_3083);
xnor U4628 (N_4628,N_3551,N_3358);
nor U4629 (N_4629,N_3809,N_3661);
nand U4630 (N_4630,N_3295,N_3696);
nor U4631 (N_4631,N_3399,N_3934);
nor U4632 (N_4632,N_3237,N_3582);
nand U4633 (N_4633,N_3752,N_3430);
xor U4634 (N_4634,N_3207,N_3984);
xnor U4635 (N_4635,N_3869,N_3507);
xor U4636 (N_4636,N_3056,N_3593);
or U4637 (N_4637,N_3289,N_3270);
and U4638 (N_4638,N_3204,N_3569);
nand U4639 (N_4639,N_3473,N_3376);
nand U4640 (N_4640,N_3312,N_3407);
nor U4641 (N_4641,N_3423,N_3750);
and U4642 (N_4642,N_3412,N_3655);
or U4643 (N_4643,N_3946,N_3219);
and U4644 (N_4644,N_3117,N_3047);
nand U4645 (N_4645,N_3820,N_3371);
nand U4646 (N_4646,N_3468,N_3924);
or U4647 (N_4647,N_3913,N_3256);
nand U4648 (N_4648,N_3152,N_3894);
nand U4649 (N_4649,N_3383,N_3483);
nor U4650 (N_4650,N_3088,N_3398);
nand U4651 (N_4651,N_3496,N_3038);
nand U4652 (N_4652,N_3439,N_3431);
nand U4653 (N_4653,N_3375,N_3342);
xor U4654 (N_4654,N_3859,N_3544);
or U4655 (N_4655,N_3763,N_3179);
xor U4656 (N_4656,N_3119,N_3539);
xor U4657 (N_4657,N_3992,N_3209);
xor U4658 (N_4658,N_3060,N_3301);
and U4659 (N_4659,N_3515,N_3988);
nor U4660 (N_4660,N_3508,N_3898);
nand U4661 (N_4661,N_3232,N_3337);
or U4662 (N_4662,N_3803,N_3990);
and U4663 (N_4663,N_3521,N_3772);
or U4664 (N_4664,N_3438,N_3907);
nor U4665 (N_4665,N_3074,N_3770);
nand U4666 (N_4666,N_3982,N_3815);
nor U4667 (N_4667,N_3702,N_3371);
or U4668 (N_4668,N_3052,N_3011);
nand U4669 (N_4669,N_3859,N_3813);
nor U4670 (N_4670,N_3375,N_3511);
nand U4671 (N_4671,N_3592,N_3249);
xnor U4672 (N_4672,N_3759,N_3556);
xnor U4673 (N_4673,N_3914,N_3425);
or U4674 (N_4674,N_3137,N_3710);
or U4675 (N_4675,N_3348,N_3931);
xnor U4676 (N_4676,N_3916,N_3697);
nand U4677 (N_4677,N_3493,N_3365);
xor U4678 (N_4678,N_3841,N_3766);
nand U4679 (N_4679,N_3289,N_3495);
or U4680 (N_4680,N_3799,N_3497);
nor U4681 (N_4681,N_3323,N_3020);
xnor U4682 (N_4682,N_3640,N_3378);
and U4683 (N_4683,N_3738,N_3294);
nor U4684 (N_4684,N_3582,N_3242);
xor U4685 (N_4685,N_3033,N_3400);
nor U4686 (N_4686,N_3650,N_3904);
xor U4687 (N_4687,N_3042,N_3195);
and U4688 (N_4688,N_3332,N_3577);
and U4689 (N_4689,N_3420,N_3390);
nor U4690 (N_4690,N_3562,N_3881);
xor U4691 (N_4691,N_3551,N_3350);
or U4692 (N_4692,N_3537,N_3543);
xor U4693 (N_4693,N_3304,N_3483);
and U4694 (N_4694,N_3091,N_3110);
nand U4695 (N_4695,N_3801,N_3445);
nand U4696 (N_4696,N_3278,N_3809);
xor U4697 (N_4697,N_3662,N_3829);
or U4698 (N_4698,N_3137,N_3697);
and U4699 (N_4699,N_3685,N_3331);
or U4700 (N_4700,N_3132,N_3087);
xor U4701 (N_4701,N_3464,N_3125);
or U4702 (N_4702,N_3742,N_3388);
or U4703 (N_4703,N_3940,N_3012);
xor U4704 (N_4704,N_3716,N_3484);
and U4705 (N_4705,N_3738,N_3230);
xor U4706 (N_4706,N_3860,N_3646);
nand U4707 (N_4707,N_3830,N_3730);
and U4708 (N_4708,N_3538,N_3742);
nor U4709 (N_4709,N_3981,N_3579);
nor U4710 (N_4710,N_3411,N_3671);
and U4711 (N_4711,N_3709,N_3172);
nand U4712 (N_4712,N_3652,N_3367);
or U4713 (N_4713,N_3539,N_3063);
xnor U4714 (N_4714,N_3573,N_3619);
xor U4715 (N_4715,N_3634,N_3921);
nor U4716 (N_4716,N_3313,N_3786);
nor U4717 (N_4717,N_3540,N_3202);
nor U4718 (N_4718,N_3173,N_3291);
nor U4719 (N_4719,N_3846,N_3461);
xnor U4720 (N_4720,N_3846,N_3093);
and U4721 (N_4721,N_3965,N_3231);
nor U4722 (N_4722,N_3253,N_3273);
nand U4723 (N_4723,N_3348,N_3183);
nor U4724 (N_4724,N_3173,N_3959);
and U4725 (N_4725,N_3763,N_3592);
nand U4726 (N_4726,N_3952,N_3064);
or U4727 (N_4727,N_3064,N_3162);
nor U4728 (N_4728,N_3234,N_3828);
nor U4729 (N_4729,N_3100,N_3309);
and U4730 (N_4730,N_3427,N_3325);
xnor U4731 (N_4731,N_3828,N_3004);
or U4732 (N_4732,N_3956,N_3939);
or U4733 (N_4733,N_3356,N_3299);
xor U4734 (N_4734,N_3463,N_3760);
nor U4735 (N_4735,N_3527,N_3593);
or U4736 (N_4736,N_3835,N_3428);
and U4737 (N_4737,N_3658,N_3575);
or U4738 (N_4738,N_3130,N_3728);
or U4739 (N_4739,N_3226,N_3699);
and U4740 (N_4740,N_3641,N_3124);
xor U4741 (N_4741,N_3706,N_3764);
nand U4742 (N_4742,N_3327,N_3852);
nand U4743 (N_4743,N_3563,N_3989);
nand U4744 (N_4744,N_3793,N_3211);
and U4745 (N_4745,N_3737,N_3928);
or U4746 (N_4746,N_3558,N_3419);
nor U4747 (N_4747,N_3335,N_3200);
nor U4748 (N_4748,N_3789,N_3630);
and U4749 (N_4749,N_3903,N_3690);
xor U4750 (N_4750,N_3046,N_3308);
or U4751 (N_4751,N_3841,N_3750);
nand U4752 (N_4752,N_3194,N_3252);
and U4753 (N_4753,N_3042,N_3617);
and U4754 (N_4754,N_3488,N_3675);
and U4755 (N_4755,N_3771,N_3377);
and U4756 (N_4756,N_3302,N_3099);
nor U4757 (N_4757,N_3876,N_3610);
and U4758 (N_4758,N_3380,N_3757);
xnor U4759 (N_4759,N_3212,N_3741);
and U4760 (N_4760,N_3547,N_3129);
and U4761 (N_4761,N_3035,N_3262);
nand U4762 (N_4762,N_3916,N_3165);
and U4763 (N_4763,N_3184,N_3927);
or U4764 (N_4764,N_3201,N_3261);
nor U4765 (N_4765,N_3759,N_3957);
xor U4766 (N_4766,N_3821,N_3596);
xor U4767 (N_4767,N_3283,N_3238);
xnor U4768 (N_4768,N_3294,N_3140);
xor U4769 (N_4769,N_3937,N_3896);
nand U4770 (N_4770,N_3652,N_3731);
xor U4771 (N_4771,N_3887,N_3950);
xnor U4772 (N_4772,N_3108,N_3616);
nand U4773 (N_4773,N_3432,N_3928);
nor U4774 (N_4774,N_3462,N_3743);
nor U4775 (N_4775,N_3390,N_3848);
nor U4776 (N_4776,N_3627,N_3817);
xnor U4777 (N_4777,N_3964,N_3579);
and U4778 (N_4778,N_3861,N_3007);
xor U4779 (N_4779,N_3995,N_3614);
or U4780 (N_4780,N_3911,N_3207);
nand U4781 (N_4781,N_3846,N_3500);
nand U4782 (N_4782,N_3290,N_3874);
nand U4783 (N_4783,N_3822,N_3610);
xnor U4784 (N_4784,N_3109,N_3468);
xnor U4785 (N_4785,N_3332,N_3318);
xnor U4786 (N_4786,N_3499,N_3314);
nor U4787 (N_4787,N_3801,N_3011);
and U4788 (N_4788,N_3992,N_3603);
xnor U4789 (N_4789,N_3879,N_3025);
and U4790 (N_4790,N_3342,N_3085);
nor U4791 (N_4791,N_3492,N_3600);
xor U4792 (N_4792,N_3218,N_3574);
nand U4793 (N_4793,N_3330,N_3307);
and U4794 (N_4794,N_3349,N_3261);
nor U4795 (N_4795,N_3950,N_3242);
nand U4796 (N_4796,N_3582,N_3688);
and U4797 (N_4797,N_3700,N_3146);
nand U4798 (N_4798,N_3995,N_3770);
nor U4799 (N_4799,N_3809,N_3830);
nor U4800 (N_4800,N_3013,N_3159);
nand U4801 (N_4801,N_3542,N_3152);
nor U4802 (N_4802,N_3900,N_3352);
xor U4803 (N_4803,N_3984,N_3533);
nor U4804 (N_4804,N_3437,N_3959);
nand U4805 (N_4805,N_3000,N_3901);
xnor U4806 (N_4806,N_3520,N_3711);
or U4807 (N_4807,N_3383,N_3818);
or U4808 (N_4808,N_3773,N_3104);
or U4809 (N_4809,N_3632,N_3038);
nor U4810 (N_4810,N_3373,N_3992);
or U4811 (N_4811,N_3745,N_3082);
and U4812 (N_4812,N_3862,N_3919);
or U4813 (N_4813,N_3752,N_3191);
or U4814 (N_4814,N_3698,N_3284);
or U4815 (N_4815,N_3876,N_3238);
nand U4816 (N_4816,N_3414,N_3452);
or U4817 (N_4817,N_3616,N_3419);
nor U4818 (N_4818,N_3268,N_3345);
xor U4819 (N_4819,N_3283,N_3666);
xor U4820 (N_4820,N_3630,N_3002);
xnor U4821 (N_4821,N_3860,N_3239);
xor U4822 (N_4822,N_3536,N_3641);
or U4823 (N_4823,N_3665,N_3548);
nor U4824 (N_4824,N_3470,N_3511);
or U4825 (N_4825,N_3879,N_3754);
and U4826 (N_4826,N_3317,N_3371);
xor U4827 (N_4827,N_3576,N_3888);
nand U4828 (N_4828,N_3363,N_3019);
and U4829 (N_4829,N_3436,N_3061);
and U4830 (N_4830,N_3152,N_3300);
xor U4831 (N_4831,N_3824,N_3240);
and U4832 (N_4832,N_3615,N_3625);
nor U4833 (N_4833,N_3860,N_3472);
xor U4834 (N_4834,N_3633,N_3204);
or U4835 (N_4835,N_3115,N_3702);
nor U4836 (N_4836,N_3501,N_3947);
nand U4837 (N_4837,N_3275,N_3538);
nor U4838 (N_4838,N_3549,N_3736);
xor U4839 (N_4839,N_3918,N_3761);
nand U4840 (N_4840,N_3528,N_3090);
xnor U4841 (N_4841,N_3728,N_3155);
xnor U4842 (N_4842,N_3540,N_3635);
or U4843 (N_4843,N_3367,N_3261);
nand U4844 (N_4844,N_3195,N_3233);
and U4845 (N_4845,N_3486,N_3662);
and U4846 (N_4846,N_3478,N_3679);
or U4847 (N_4847,N_3111,N_3312);
nor U4848 (N_4848,N_3715,N_3788);
nor U4849 (N_4849,N_3837,N_3224);
or U4850 (N_4850,N_3796,N_3572);
or U4851 (N_4851,N_3122,N_3427);
nor U4852 (N_4852,N_3723,N_3714);
xor U4853 (N_4853,N_3414,N_3954);
and U4854 (N_4854,N_3143,N_3978);
and U4855 (N_4855,N_3416,N_3616);
or U4856 (N_4856,N_3204,N_3386);
xnor U4857 (N_4857,N_3715,N_3950);
nor U4858 (N_4858,N_3878,N_3299);
nor U4859 (N_4859,N_3083,N_3396);
or U4860 (N_4860,N_3636,N_3724);
and U4861 (N_4861,N_3380,N_3666);
nand U4862 (N_4862,N_3441,N_3029);
nor U4863 (N_4863,N_3710,N_3097);
xnor U4864 (N_4864,N_3607,N_3487);
nor U4865 (N_4865,N_3162,N_3613);
xnor U4866 (N_4866,N_3831,N_3986);
xor U4867 (N_4867,N_3916,N_3419);
nand U4868 (N_4868,N_3308,N_3092);
and U4869 (N_4869,N_3221,N_3900);
and U4870 (N_4870,N_3892,N_3467);
xnor U4871 (N_4871,N_3644,N_3412);
nor U4872 (N_4872,N_3018,N_3325);
and U4873 (N_4873,N_3378,N_3673);
xnor U4874 (N_4874,N_3178,N_3908);
nor U4875 (N_4875,N_3880,N_3507);
xnor U4876 (N_4876,N_3832,N_3176);
or U4877 (N_4877,N_3140,N_3121);
nor U4878 (N_4878,N_3046,N_3351);
nand U4879 (N_4879,N_3930,N_3363);
xor U4880 (N_4880,N_3344,N_3751);
or U4881 (N_4881,N_3140,N_3773);
and U4882 (N_4882,N_3890,N_3970);
xor U4883 (N_4883,N_3065,N_3348);
xor U4884 (N_4884,N_3960,N_3917);
nor U4885 (N_4885,N_3906,N_3520);
and U4886 (N_4886,N_3429,N_3987);
or U4887 (N_4887,N_3276,N_3916);
xor U4888 (N_4888,N_3911,N_3053);
or U4889 (N_4889,N_3070,N_3273);
or U4890 (N_4890,N_3701,N_3859);
nor U4891 (N_4891,N_3456,N_3143);
or U4892 (N_4892,N_3427,N_3538);
or U4893 (N_4893,N_3680,N_3845);
nand U4894 (N_4894,N_3478,N_3563);
xnor U4895 (N_4895,N_3690,N_3430);
xor U4896 (N_4896,N_3177,N_3154);
or U4897 (N_4897,N_3268,N_3711);
and U4898 (N_4898,N_3223,N_3400);
or U4899 (N_4899,N_3204,N_3848);
and U4900 (N_4900,N_3055,N_3455);
and U4901 (N_4901,N_3886,N_3228);
and U4902 (N_4902,N_3112,N_3733);
xnor U4903 (N_4903,N_3841,N_3635);
or U4904 (N_4904,N_3029,N_3289);
xnor U4905 (N_4905,N_3160,N_3677);
and U4906 (N_4906,N_3933,N_3329);
nor U4907 (N_4907,N_3765,N_3100);
and U4908 (N_4908,N_3170,N_3039);
nor U4909 (N_4909,N_3010,N_3832);
or U4910 (N_4910,N_3949,N_3786);
or U4911 (N_4911,N_3374,N_3666);
nand U4912 (N_4912,N_3220,N_3522);
nor U4913 (N_4913,N_3976,N_3536);
or U4914 (N_4914,N_3687,N_3995);
xor U4915 (N_4915,N_3766,N_3219);
nor U4916 (N_4916,N_3791,N_3774);
nor U4917 (N_4917,N_3179,N_3884);
or U4918 (N_4918,N_3554,N_3325);
and U4919 (N_4919,N_3829,N_3683);
and U4920 (N_4920,N_3779,N_3954);
nand U4921 (N_4921,N_3719,N_3117);
and U4922 (N_4922,N_3307,N_3097);
nor U4923 (N_4923,N_3457,N_3598);
or U4924 (N_4924,N_3879,N_3933);
and U4925 (N_4925,N_3446,N_3557);
nand U4926 (N_4926,N_3910,N_3344);
nand U4927 (N_4927,N_3052,N_3121);
nor U4928 (N_4928,N_3777,N_3952);
nand U4929 (N_4929,N_3071,N_3145);
or U4930 (N_4930,N_3174,N_3676);
nor U4931 (N_4931,N_3263,N_3760);
or U4932 (N_4932,N_3386,N_3329);
or U4933 (N_4933,N_3627,N_3753);
nor U4934 (N_4934,N_3590,N_3120);
nand U4935 (N_4935,N_3812,N_3854);
or U4936 (N_4936,N_3015,N_3211);
and U4937 (N_4937,N_3360,N_3678);
nor U4938 (N_4938,N_3758,N_3062);
nor U4939 (N_4939,N_3476,N_3016);
xor U4940 (N_4940,N_3209,N_3931);
or U4941 (N_4941,N_3907,N_3387);
and U4942 (N_4942,N_3169,N_3381);
and U4943 (N_4943,N_3956,N_3476);
nor U4944 (N_4944,N_3545,N_3689);
and U4945 (N_4945,N_3794,N_3180);
xnor U4946 (N_4946,N_3180,N_3695);
xnor U4947 (N_4947,N_3208,N_3515);
nand U4948 (N_4948,N_3972,N_3617);
nor U4949 (N_4949,N_3011,N_3574);
xor U4950 (N_4950,N_3360,N_3187);
nand U4951 (N_4951,N_3809,N_3820);
and U4952 (N_4952,N_3613,N_3708);
and U4953 (N_4953,N_3843,N_3065);
xnor U4954 (N_4954,N_3007,N_3541);
nand U4955 (N_4955,N_3361,N_3479);
nor U4956 (N_4956,N_3864,N_3807);
nor U4957 (N_4957,N_3779,N_3708);
or U4958 (N_4958,N_3846,N_3750);
xor U4959 (N_4959,N_3193,N_3821);
and U4960 (N_4960,N_3090,N_3239);
nand U4961 (N_4961,N_3293,N_3061);
xnor U4962 (N_4962,N_3045,N_3805);
xor U4963 (N_4963,N_3430,N_3713);
and U4964 (N_4964,N_3746,N_3048);
xnor U4965 (N_4965,N_3646,N_3718);
and U4966 (N_4966,N_3970,N_3358);
nor U4967 (N_4967,N_3961,N_3962);
nor U4968 (N_4968,N_3154,N_3628);
nand U4969 (N_4969,N_3252,N_3584);
and U4970 (N_4970,N_3663,N_3119);
xnor U4971 (N_4971,N_3563,N_3551);
or U4972 (N_4972,N_3097,N_3968);
xor U4973 (N_4973,N_3147,N_3261);
nor U4974 (N_4974,N_3904,N_3675);
nand U4975 (N_4975,N_3047,N_3604);
nor U4976 (N_4976,N_3667,N_3968);
and U4977 (N_4977,N_3834,N_3296);
nor U4978 (N_4978,N_3627,N_3042);
or U4979 (N_4979,N_3672,N_3624);
xor U4980 (N_4980,N_3804,N_3049);
nor U4981 (N_4981,N_3491,N_3131);
nand U4982 (N_4982,N_3898,N_3661);
nor U4983 (N_4983,N_3099,N_3935);
nor U4984 (N_4984,N_3182,N_3443);
and U4985 (N_4985,N_3879,N_3479);
and U4986 (N_4986,N_3897,N_3089);
or U4987 (N_4987,N_3168,N_3011);
xor U4988 (N_4988,N_3323,N_3140);
xnor U4989 (N_4989,N_3366,N_3988);
and U4990 (N_4990,N_3469,N_3137);
xnor U4991 (N_4991,N_3569,N_3416);
nor U4992 (N_4992,N_3357,N_3692);
xnor U4993 (N_4993,N_3258,N_3871);
nand U4994 (N_4994,N_3238,N_3118);
or U4995 (N_4995,N_3605,N_3190);
nand U4996 (N_4996,N_3498,N_3062);
or U4997 (N_4997,N_3118,N_3312);
xor U4998 (N_4998,N_3812,N_3122);
or U4999 (N_4999,N_3093,N_3771);
nor U5000 (N_5000,N_4471,N_4262);
nand U5001 (N_5001,N_4584,N_4160);
nand U5002 (N_5002,N_4637,N_4945);
or U5003 (N_5003,N_4914,N_4545);
or U5004 (N_5004,N_4589,N_4339);
nand U5005 (N_5005,N_4394,N_4617);
or U5006 (N_5006,N_4614,N_4532);
and U5007 (N_5007,N_4598,N_4707);
xnor U5008 (N_5008,N_4890,N_4655);
xor U5009 (N_5009,N_4091,N_4196);
nor U5010 (N_5010,N_4712,N_4088);
or U5011 (N_5011,N_4951,N_4922);
nand U5012 (N_5012,N_4536,N_4549);
xnor U5013 (N_5013,N_4029,N_4492);
nor U5014 (N_5014,N_4576,N_4984);
and U5015 (N_5015,N_4155,N_4817);
xor U5016 (N_5016,N_4008,N_4554);
and U5017 (N_5017,N_4408,N_4791);
xor U5018 (N_5018,N_4104,N_4676);
nor U5019 (N_5019,N_4907,N_4487);
nand U5020 (N_5020,N_4470,N_4601);
nand U5021 (N_5021,N_4942,N_4926);
and U5022 (N_5022,N_4904,N_4916);
and U5023 (N_5023,N_4322,N_4131);
nor U5024 (N_5024,N_4099,N_4895);
or U5025 (N_5025,N_4047,N_4546);
or U5026 (N_5026,N_4948,N_4181);
nor U5027 (N_5027,N_4575,N_4176);
or U5028 (N_5028,N_4718,N_4445);
nand U5029 (N_5029,N_4423,N_4743);
or U5030 (N_5030,N_4499,N_4596);
or U5031 (N_5031,N_4043,N_4038);
xor U5032 (N_5032,N_4253,N_4792);
and U5033 (N_5033,N_4337,N_4336);
xnor U5034 (N_5034,N_4971,N_4952);
or U5035 (N_5035,N_4870,N_4986);
nand U5036 (N_5036,N_4095,N_4831);
xnor U5037 (N_5037,N_4422,N_4703);
xnor U5038 (N_5038,N_4530,N_4562);
nand U5039 (N_5039,N_4608,N_4180);
nor U5040 (N_5040,N_4663,N_4863);
and U5041 (N_5041,N_4194,N_4868);
or U5042 (N_5042,N_4212,N_4654);
and U5043 (N_5043,N_4526,N_4117);
and U5044 (N_5044,N_4508,N_4533);
and U5045 (N_5045,N_4889,N_4325);
nand U5046 (N_5046,N_4192,N_4938);
nor U5047 (N_5047,N_4275,N_4885);
or U5048 (N_5048,N_4209,N_4820);
nand U5049 (N_5049,N_4615,N_4051);
or U5050 (N_5050,N_4740,N_4515);
nor U5051 (N_5051,N_4041,N_4841);
nand U5052 (N_5052,N_4271,N_4704);
or U5053 (N_5053,N_4719,N_4344);
xnor U5054 (N_5054,N_4130,N_4363);
nand U5055 (N_5055,N_4741,N_4141);
xor U5056 (N_5056,N_4026,N_4071);
nor U5057 (N_5057,N_4396,N_4065);
or U5058 (N_5058,N_4233,N_4427);
xor U5059 (N_5059,N_4923,N_4933);
xnor U5060 (N_5060,N_4972,N_4757);
or U5061 (N_5061,N_4812,N_4714);
nor U5062 (N_5062,N_4222,N_4643);
nand U5063 (N_5063,N_4382,N_4838);
xnor U5064 (N_5064,N_4320,N_4200);
or U5065 (N_5065,N_4268,N_4767);
xnor U5066 (N_5066,N_4717,N_4659);
nor U5067 (N_5067,N_4444,N_4847);
or U5068 (N_5068,N_4054,N_4298);
nor U5069 (N_5069,N_4686,N_4706);
xor U5070 (N_5070,N_4779,N_4512);
nor U5071 (N_5071,N_4775,N_4855);
xor U5072 (N_5072,N_4033,N_4207);
nand U5073 (N_5073,N_4888,N_4928);
xor U5074 (N_5074,N_4254,N_4014);
or U5075 (N_5075,N_4144,N_4699);
and U5076 (N_5076,N_4488,N_4429);
xnor U5077 (N_5077,N_4030,N_4806);
xnor U5078 (N_5078,N_4467,N_4896);
and U5079 (N_5079,N_4446,N_4786);
nand U5080 (N_5080,N_4419,N_4833);
nand U5081 (N_5081,N_4188,N_4224);
and U5082 (N_5082,N_4208,N_4688);
and U5083 (N_5083,N_4352,N_4119);
nand U5084 (N_5084,N_4813,N_4929);
or U5085 (N_5085,N_4992,N_4609);
xor U5086 (N_5086,N_4366,N_4527);
and U5087 (N_5087,N_4050,N_4101);
and U5088 (N_5088,N_4883,N_4338);
xnor U5089 (N_5089,N_4510,N_4305);
or U5090 (N_5090,N_4872,N_4357);
or U5091 (N_5091,N_4257,N_4435);
or U5092 (N_5092,N_4874,N_4912);
nand U5093 (N_5093,N_4878,N_4146);
nor U5094 (N_5094,N_4534,N_4186);
or U5095 (N_5095,N_4826,N_4226);
nand U5096 (N_5096,N_4607,N_4441);
nand U5097 (N_5097,N_4997,N_4129);
nand U5098 (N_5098,N_4594,N_4206);
nand U5099 (N_5099,N_4183,N_4683);
nor U5100 (N_5100,N_4436,N_4134);
or U5101 (N_5101,N_4279,N_4987);
nand U5102 (N_5102,N_4836,N_4317);
nand U5103 (N_5103,N_4892,N_4684);
nand U5104 (N_5104,N_4877,N_4003);
or U5105 (N_5105,N_4004,N_4383);
xor U5106 (N_5106,N_4705,N_4649);
nand U5107 (N_5107,N_4613,N_4165);
nand U5108 (N_5108,N_4407,N_4780);
nor U5109 (N_5109,N_4314,N_4873);
or U5110 (N_5110,N_4140,N_4177);
nand U5111 (N_5111,N_4302,N_4135);
nor U5112 (N_5112,N_4893,N_4284);
nand U5113 (N_5113,N_4572,N_4620);
xnor U5114 (N_5114,N_4341,N_4650);
or U5115 (N_5115,N_4789,N_4159);
xnor U5116 (N_5116,N_4588,N_4976);
nand U5117 (N_5117,N_4236,N_4090);
and U5118 (N_5118,N_4542,N_4642);
and U5119 (N_5119,N_4681,N_4956);
nor U5120 (N_5120,N_4694,N_4535);
xor U5121 (N_5121,N_4720,N_4970);
nand U5122 (N_5122,N_4934,N_4055);
and U5123 (N_5123,N_4387,N_4677);
nor U5124 (N_5124,N_4031,N_4981);
nor U5125 (N_5125,N_4269,N_4485);
nand U5126 (N_5126,N_4519,N_4678);
nor U5127 (N_5127,N_4425,N_4784);
or U5128 (N_5128,N_4447,N_4328);
xor U5129 (N_5129,N_4231,N_4539);
nand U5130 (N_5130,N_4368,N_4056);
and U5131 (N_5131,N_4932,N_4538);
xor U5132 (N_5132,N_4968,N_4799);
nor U5133 (N_5133,N_4518,N_4709);
nand U5134 (N_5134,N_4566,N_4203);
or U5135 (N_5135,N_4244,N_4045);
and U5136 (N_5136,N_4288,N_4067);
or U5137 (N_5137,N_4964,N_4392);
or U5138 (N_5138,N_4816,N_4927);
or U5139 (N_5139,N_4115,N_4658);
xnor U5140 (N_5140,N_4046,N_4547);
and U5141 (N_5141,N_4397,N_4738);
nand U5142 (N_5142,N_4410,N_4733);
and U5143 (N_5143,N_4591,N_4028);
or U5144 (N_5144,N_4763,N_4310);
and U5145 (N_5145,N_4500,N_4327);
xnor U5146 (N_5146,N_4721,N_4876);
nor U5147 (N_5147,N_4808,N_4901);
or U5148 (N_5148,N_4283,N_4145);
xor U5149 (N_5149,N_4248,N_4568);
and U5150 (N_5150,N_4991,N_4225);
and U5151 (N_5151,N_4675,N_4316);
xnor U5152 (N_5152,N_4300,N_4502);
or U5153 (N_5153,N_4440,N_4100);
or U5154 (N_5154,N_4960,N_4079);
xor U5155 (N_5155,N_4053,N_4304);
or U5156 (N_5156,N_4857,N_4162);
or U5157 (N_5157,N_4449,N_4918);
or U5158 (N_5158,N_4012,N_4552);
xor U5159 (N_5159,N_4370,N_4085);
or U5160 (N_5160,N_4521,N_4076);
and U5161 (N_5161,N_4377,N_4689);
and U5162 (N_5162,N_4967,N_4274);
nor U5163 (N_5163,N_4651,N_4980);
and U5164 (N_5164,N_4661,N_4834);
xnor U5165 (N_5165,N_4749,N_4798);
nor U5166 (N_5166,N_4680,N_4815);
nor U5167 (N_5167,N_4742,N_4656);
and U5168 (N_5168,N_4173,N_4944);
xnor U5169 (N_5169,N_4021,N_4010);
and U5170 (N_5170,N_4124,N_4151);
nand U5171 (N_5171,N_4998,N_4715);
xnor U5172 (N_5172,N_4416,N_4865);
xnor U5173 (N_5173,N_4850,N_4286);
nor U5174 (N_5174,N_4781,N_4120);
and U5175 (N_5175,N_4657,N_4406);
nand U5176 (N_5176,N_4541,N_4195);
and U5177 (N_5177,N_4511,N_4567);
or U5178 (N_5178,N_4957,N_4946);
and U5179 (N_5179,N_4007,N_4632);
or U5180 (N_5180,N_4861,N_4975);
xnor U5181 (N_5181,N_4999,N_4641);
or U5182 (N_5182,N_4788,N_4579);
or U5183 (N_5183,N_4765,N_4285);
or U5184 (N_5184,N_4402,N_4674);
nand U5185 (N_5185,N_4832,N_4062);
nor U5186 (N_5186,N_4520,N_4548);
xnor U5187 (N_5187,N_4747,N_4645);
nand U5188 (N_5188,N_4947,N_4334);
and U5189 (N_5189,N_4830,N_4580);
nor U5190 (N_5190,N_4710,N_4218);
nand U5191 (N_5191,N_4306,N_4531);
nand U5192 (N_5192,N_4060,N_4586);
nor U5193 (N_5193,N_4480,N_4561);
or U5194 (N_5194,N_4154,N_4727);
nor U5195 (N_5195,N_4204,N_4513);
nor U5196 (N_5196,N_4260,N_4428);
xnor U5197 (N_5197,N_4197,N_4070);
and U5198 (N_5198,N_4000,N_4941);
xor U5199 (N_5199,N_4910,N_4624);
xnor U5200 (N_5200,N_4287,N_4246);
nand U5201 (N_5201,N_4551,N_4315);
nor U5202 (N_5202,N_4295,N_4389);
nand U5203 (N_5203,N_4193,N_4221);
or U5204 (N_5204,N_4125,N_4768);
and U5205 (N_5205,N_4149,N_4219);
nand U5206 (N_5206,N_4662,N_4309);
and U5207 (N_5207,N_4002,N_4171);
and U5208 (N_5208,N_4034,N_4015);
and U5209 (N_5209,N_4042,N_4793);
nor U5210 (N_5210,N_4856,N_4109);
xnor U5211 (N_5211,N_4438,N_4454);
or U5212 (N_5212,N_4503,N_4859);
nor U5213 (N_5213,N_4629,N_4107);
and U5214 (N_5214,N_4582,N_4577);
or U5215 (N_5215,N_4189,N_4092);
and U5216 (N_5216,N_4434,N_4032);
and U5217 (N_5217,N_4573,N_4354);
and U5218 (N_5218,N_4824,N_4736);
nand U5219 (N_5219,N_4665,N_4342);
and U5220 (N_5220,N_4294,N_4660);
xnor U5221 (N_5221,N_4773,N_4278);
xor U5222 (N_5222,N_4073,N_4756);
nor U5223 (N_5223,N_4698,N_4350);
or U5224 (N_5224,N_4989,N_4086);
xnor U5225 (N_5225,N_4058,N_4565);
xnor U5226 (N_5226,N_4769,N_4600);
or U5227 (N_5227,N_4023,N_4909);
nor U5228 (N_5228,N_4475,N_4735);
nor U5229 (N_5229,N_4668,N_4498);
and U5230 (N_5230,N_4908,N_4163);
or U5231 (N_5231,N_4619,N_4112);
xnor U5232 (N_5232,N_4333,N_4628);
nor U5233 (N_5233,N_4977,N_4574);
nor U5234 (N_5234,N_4994,N_4955);
and U5235 (N_5235,N_4583,N_4569);
and U5236 (N_5236,N_4880,N_4361);
xor U5237 (N_5237,N_4887,N_4852);
or U5238 (N_5238,N_4190,N_4522);
or U5239 (N_5239,N_4481,N_4018);
and U5240 (N_5240,N_4148,N_4867);
nor U5241 (N_5241,N_4473,N_4647);
and U5242 (N_5242,N_4412,N_4858);
nand U5243 (N_5243,N_4770,N_4057);
xor U5244 (N_5244,N_4814,N_4525);
xor U5245 (N_5245,N_4965,N_4232);
xnor U5246 (N_5246,N_4543,N_4068);
xnor U5247 (N_5247,N_4172,N_4372);
or U5248 (N_5248,N_4039,N_4006);
and U5249 (N_5249,N_4182,N_4954);
and U5250 (N_5250,N_4343,N_4962);
and U5251 (N_5251,N_4009,N_4161);
or U5252 (N_5252,N_4752,N_4842);
xor U5253 (N_5253,N_4087,N_4332);
and U5254 (N_5254,N_4708,N_4762);
nand U5255 (N_5255,N_4556,N_4638);
nand U5256 (N_5256,N_4292,N_4381);
and U5257 (N_5257,N_4673,N_4102);
nor U5258 (N_5258,N_4474,N_4760);
and U5259 (N_5259,N_4256,N_4465);
or U5260 (N_5260,N_4001,N_4585);
nor U5261 (N_5261,N_4745,N_4157);
and U5262 (N_5262,N_4881,N_4595);
or U5263 (N_5263,N_4138,N_4078);
xor U5264 (N_5264,N_4979,N_4367);
xor U5265 (N_5265,N_4170,N_4958);
and U5266 (N_5266,N_4346,N_4199);
nand U5267 (N_5267,N_4599,N_4150);
xnor U5268 (N_5268,N_4995,N_4625);
or U5269 (N_5269,N_4633,N_4516);
xor U5270 (N_5270,N_4722,N_4634);
nor U5271 (N_5271,N_4137,N_4022);
nor U5272 (N_5272,N_4251,N_4216);
nand U5273 (N_5273,N_4737,N_4025);
or U5274 (N_5274,N_4646,N_4882);
or U5275 (N_5275,N_4239,N_4621);
xor U5276 (N_5276,N_4924,N_4729);
nor U5277 (N_5277,N_4682,N_4731);
and U5278 (N_5278,N_4631,N_4825);
xnor U5279 (N_5279,N_4853,N_4671);
and U5280 (N_5280,N_4730,N_4234);
and U5281 (N_5281,N_4755,N_4744);
xnor U5282 (N_5282,N_4917,N_4851);
and U5283 (N_5283,N_4461,N_4027);
nand U5284 (N_5284,N_4395,N_4460);
or U5285 (N_5285,N_4884,N_4349);
nand U5286 (N_5286,N_4862,N_4795);
nor U5287 (N_5287,N_4456,N_4311);
nand U5288 (N_5288,N_4996,N_4153);
xnor U5289 (N_5289,N_4803,N_4243);
nor U5290 (N_5290,N_4894,N_4228);
nor U5291 (N_5291,N_4261,N_4017);
and U5292 (N_5292,N_4403,N_4122);
and U5293 (N_5293,N_4761,N_4011);
xor U5294 (N_5294,N_4774,N_4993);
and U5295 (N_5295,N_4493,N_4409);
nand U5296 (N_5296,N_4811,N_4871);
and U5297 (N_5297,N_4345,N_4961);
nand U5298 (N_5298,N_4420,N_4670);
nand U5299 (N_5299,N_4564,N_4364);
nor U5300 (N_5300,N_4509,N_4167);
xnor U5301 (N_5301,N_4804,N_4466);
xor U5302 (N_5302,N_4477,N_4691);
nor U5303 (N_5303,N_4754,N_4590);
or U5304 (N_5304,N_4690,N_4431);
nor U5305 (N_5305,N_4950,N_4911);
and U5306 (N_5306,N_4476,N_4953);
and U5307 (N_5307,N_4772,N_4277);
xnor U5308 (N_5308,N_4201,N_4297);
nor U5309 (N_5309,N_4846,N_4483);
or U5310 (N_5310,N_4990,N_4255);
or U5311 (N_5311,N_4351,N_4906);
or U5312 (N_5312,N_4083,N_4829);
nand U5313 (N_5313,N_4644,N_4652);
xor U5314 (N_5314,N_4365,N_4616);
nor U5315 (N_5315,N_4184,N_4164);
or U5316 (N_5316,N_4818,N_4238);
nand U5317 (N_5317,N_4358,N_4840);
xnor U5318 (N_5318,N_4211,N_4347);
nand U5319 (N_5319,N_4093,N_4462);
xnor U5320 (N_5320,N_4005,N_4430);
nor U5321 (N_5321,N_4782,N_4214);
or U5322 (N_5322,N_4692,N_4237);
or U5323 (N_5323,N_4400,N_4711);
or U5324 (N_5324,N_4270,N_4902);
nand U5325 (N_5325,N_4866,N_4915);
nor U5326 (N_5326,N_4726,N_4081);
xnor U5327 (N_5327,N_4442,N_4728);
or U5328 (N_5328,N_4507,N_4899);
or U5329 (N_5329,N_4685,N_4903);
nand U5330 (N_5330,N_4399,N_4303);
or U5331 (N_5331,N_4724,N_4390);
xor U5332 (N_5332,N_4725,N_4578);
nor U5333 (N_5333,N_4291,N_4605);
xor U5334 (N_5334,N_4052,N_4307);
nand U5335 (N_5335,N_4653,N_4105);
or U5336 (N_5336,N_4417,N_4759);
nand U5337 (N_5337,N_4404,N_4766);
nor U5338 (N_5338,N_4080,N_4355);
nor U5339 (N_5339,N_4603,N_4864);
xor U5340 (N_5340,N_4020,N_4191);
xor U5341 (N_5341,N_4827,N_4179);
nand U5342 (N_5342,N_4937,N_4697);
nand U5343 (N_5343,N_4356,N_4802);
and U5344 (N_5344,N_4949,N_4453);
or U5345 (N_5345,N_4110,N_4514);
nand U5346 (N_5346,N_4069,N_4432);
and U5347 (N_5347,N_4024,N_4178);
and U5348 (N_5348,N_4540,N_4648);
xor U5349 (N_5349,N_4463,N_4597);
xor U5350 (N_5350,N_4920,N_4116);
or U5351 (N_5351,N_4464,N_4869);
xnor U5352 (N_5352,N_4822,N_4426);
xor U5353 (N_5353,N_4571,N_4044);
and U5354 (N_5354,N_4391,N_4785);
nor U5355 (N_5355,N_4592,N_4494);
and U5356 (N_5356,N_4626,N_4169);
nand U5357 (N_5357,N_4983,N_4443);
nand U5358 (N_5358,N_4142,N_4611);
nand U5359 (N_5359,N_4544,N_4205);
xor U5360 (N_5360,N_4898,N_4348);
or U5361 (N_5361,N_4240,N_4281);
or U5362 (N_5362,N_4258,N_4790);
nor U5363 (N_5363,N_4734,N_4469);
nor U5364 (N_5364,N_4959,N_4839);
and U5365 (N_5365,N_4235,N_4259);
xor U5366 (N_5366,N_4837,N_4771);
or U5367 (N_5367,N_4136,N_4973);
xor U5368 (N_5368,N_4411,N_4319);
nor U5369 (N_5369,N_4293,N_4969);
nor U5370 (N_5370,N_4560,N_4249);
and U5371 (N_5371,N_4335,N_4921);
nor U5372 (N_5372,N_4123,N_4220);
xnor U5373 (N_5373,N_4468,N_4491);
nand U5374 (N_5374,N_4787,N_4340);
or U5375 (N_5375,N_4451,N_4776);
xor U5376 (N_5376,N_4604,N_4982);
nand U5377 (N_5377,N_4210,N_4750);
or U5378 (N_5378,N_4247,N_4482);
xnor U5379 (N_5379,N_4373,N_4794);
nor U5380 (N_5380,N_4418,N_4523);
nand U5381 (N_5381,N_4398,N_4074);
or U5382 (N_5382,N_4764,N_4623);
nor U5383 (N_5383,N_4299,N_4939);
nor U5384 (N_5384,N_4702,N_4700);
nand U5385 (N_5385,N_4848,N_4168);
xor U5386 (N_5386,N_4801,N_4324);
nand U5387 (N_5387,N_4809,N_4943);
or U5388 (N_5388,N_4679,N_4486);
or U5389 (N_5389,N_4405,N_4424);
nor U5390 (N_5390,N_4301,N_4985);
or U5391 (N_5391,N_4312,N_4393);
and U5392 (N_5392,N_4040,N_4529);
xor U5393 (N_5393,N_4223,N_4879);
xnor U5394 (N_5394,N_4187,N_4267);
nor U5395 (N_5395,N_4118,N_4369);
xnor U5396 (N_5396,N_4783,N_4886);
nand U5397 (N_5397,N_4797,N_4931);
nand U5398 (N_5398,N_4553,N_4266);
or U5399 (N_5399,N_4121,N_4413);
nor U5400 (N_5400,N_4753,N_4640);
nand U5401 (N_5401,N_4618,N_4158);
xor U5402 (N_5402,N_4059,N_4126);
nor U5403 (N_5403,N_4061,N_4835);
or U5404 (N_5404,N_4630,N_4359);
xor U5405 (N_5405,N_4152,N_4810);
or U5406 (N_5406,N_4940,N_4156);
or U5407 (N_5407,N_4988,N_4495);
nand U5408 (N_5408,N_4897,N_4290);
xor U5409 (N_5409,N_4935,N_4805);
nor U5410 (N_5410,N_4606,N_4064);
nand U5411 (N_5411,N_4353,N_4245);
nor U5412 (N_5412,N_4748,N_4376);
and U5413 (N_5413,N_4555,N_4384);
nand U5414 (N_5414,N_4213,N_4252);
xor U5415 (N_5415,N_4570,N_4635);
and U5416 (N_5416,N_4739,N_4506);
xnor U5417 (N_5417,N_4414,N_4891);
xor U5418 (N_5418,N_4103,N_4035);
nand U5419 (N_5419,N_4166,N_4746);
and U5420 (N_5420,N_4378,N_4280);
or U5421 (N_5421,N_4558,N_4106);
and U5422 (N_5422,N_4289,N_4693);
and U5423 (N_5423,N_4557,N_4321);
nand U5424 (N_5424,N_4437,N_4672);
or U5425 (N_5425,N_4496,N_4386);
or U5426 (N_5426,N_4296,N_4272);
xor U5427 (N_5427,N_4777,N_4501);
or U5428 (N_5428,N_4550,N_4821);
xor U5429 (N_5429,N_4127,N_4593);
nand U5430 (N_5430,N_4687,N_4505);
nand U5431 (N_5431,N_4978,N_4097);
or U5432 (N_5432,N_4075,N_4385);
nand U5433 (N_5433,N_4913,N_4843);
and U5434 (N_5434,N_4013,N_4936);
xor U5435 (N_5435,N_4497,N_4326);
xnor U5436 (N_5436,N_4174,N_4215);
or U5437 (N_5437,N_4823,N_4066);
xor U5438 (N_5438,N_4537,N_4147);
or U5439 (N_5439,N_4854,N_4919);
or U5440 (N_5440,N_4133,N_4612);
and U5441 (N_5441,N_4610,N_4844);
nand U5442 (N_5442,N_4966,N_4930);
nand U5443 (N_5443,N_4925,N_4563);
nor U5444 (N_5444,N_4669,N_4380);
xnor U5445 (N_5445,N_4667,N_4371);
xnor U5446 (N_5446,N_4900,N_4559);
nor U5447 (N_5447,N_4128,N_4263);
or U5448 (N_5448,N_4143,N_4751);
nor U5449 (N_5449,N_4063,N_4388);
or U5450 (N_5450,N_4330,N_4250);
nand U5451 (N_5451,N_4113,N_4323);
or U5452 (N_5452,N_4450,N_4094);
nor U5453 (N_5453,N_4528,N_4108);
nor U5454 (N_5454,N_4963,N_4375);
xor U5455 (N_5455,N_4489,N_4360);
nand U5456 (N_5456,N_4265,N_4448);
or U5457 (N_5457,N_4778,N_4082);
or U5458 (N_5458,N_4308,N_4227);
nand U5459 (N_5459,N_4627,N_4723);
and U5460 (N_5460,N_4401,N_4484);
or U5461 (N_5461,N_4273,N_4587);
nand U5462 (N_5462,N_4504,N_4807);
and U5463 (N_5463,N_4077,N_4282);
or U5464 (N_5464,N_4472,N_4490);
nor U5465 (N_5465,N_4202,N_4132);
nor U5466 (N_5466,N_4049,N_4229);
and U5467 (N_5467,N_4701,N_4517);
or U5468 (N_5468,N_4318,N_4139);
or U5469 (N_5469,N_4636,N_4098);
and U5470 (N_5470,N_4379,N_4374);
and U5471 (N_5471,N_4800,N_4732);
or U5472 (N_5472,N_4114,N_4622);
xor U5473 (N_5473,N_4230,N_4602);
and U5474 (N_5474,N_4048,N_4037);
or U5475 (N_5475,N_4185,N_4713);
or U5476 (N_5476,N_4524,N_4276);
and U5477 (N_5477,N_4452,N_4845);
nor U5478 (N_5478,N_4217,N_4019);
xnor U5479 (N_5479,N_4581,N_4479);
nand U5480 (N_5480,N_4875,N_4796);
xnor U5481 (N_5481,N_4415,N_4455);
or U5482 (N_5482,N_4695,N_4758);
xor U5483 (N_5483,N_4849,N_4860);
xnor U5484 (N_5484,N_4457,N_4458);
nor U5485 (N_5485,N_4313,N_4459);
or U5486 (N_5486,N_4439,N_4696);
nand U5487 (N_5487,N_4639,N_4089);
nand U5488 (N_5488,N_4819,N_4974);
nor U5489 (N_5489,N_4329,N_4716);
xor U5490 (N_5490,N_4242,N_4664);
or U5491 (N_5491,N_4666,N_4421);
and U5492 (N_5492,N_4036,N_4828);
nand U5493 (N_5493,N_4433,N_4331);
nor U5494 (N_5494,N_4096,N_4084);
nand U5495 (N_5495,N_4111,N_4241);
and U5496 (N_5496,N_4198,N_4016);
nor U5497 (N_5497,N_4478,N_4264);
nand U5498 (N_5498,N_4072,N_4175);
xor U5499 (N_5499,N_4362,N_4905);
and U5500 (N_5500,N_4724,N_4944);
and U5501 (N_5501,N_4783,N_4022);
or U5502 (N_5502,N_4911,N_4303);
and U5503 (N_5503,N_4465,N_4300);
or U5504 (N_5504,N_4262,N_4006);
nand U5505 (N_5505,N_4120,N_4171);
nand U5506 (N_5506,N_4640,N_4080);
or U5507 (N_5507,N_4030,N_4467);
and U5508 (N_5508,N_4236,N_4600);
xor U5509 (N_5509,N_4784,N_4526);
nand U5510 (N_5510,N_4287,N_4915);
nand U5511 (N_5511,N_4967,N_4199);
and U5512 (N_5512,N_4301,N_4556);
nor U5513 (N_5513,N_4731,N_4492);
nand U5514 (N_5514,N_4621,N_4614);
and U5515 (N_5515,N_4002,N_4348);
nor U5516 (N_5516,N_4367,N_4677);
nand U5517 (N_5517,N_4243,N_4590);
xor U5518 (N_5518,N_4666,N_4966);
xnor U5519 (N_5519,N_4897,N_4089);
nor U5520 (N_5520,N_4340,N_4474);
and U5521 (N_5521,N_4903,N_4911);
nor U5522 (N_5522,N_4134,N_4621);
and U5523 (N_5523,N_4575,N_4134);
and U5524 (N_5524,N_4076,N_4425);
and U5525 (N_5525,N_4070,N_4608);
xor U5526 (N_5526,N_4395,N_4123);
nand U5527 (N_5527,N_4308,N_4453);
nor U5528 (N_5528,N_4793,N_4210);
nor U5529 (N_5529,N_4777,N_4403);
xor U5530 (N_5530,N_4613,N_4117);
or U5531 (N_5531,N_4879,N_4018);
and U5532 (N_5532,N_4044,N_4935);
and U5533 (N_5533,N_4260,N_4104);
nor U5534 (N_5534,N_4574,N_4135);
and U5535 (N_5535,N_4192,N_4880);
xnor U5536 (N_5536,N_4572,N_4422);
or U5537 (N_5537,N_4372,N_4743);
nor U5538 (N_5538,N_4395,N_4011);
xnor U5539 (N_5539,N_4508,N_4014);
or U5540 (N_5540,N_4041,N_4441);
nand U5541 (N_5541,N_4439,N_4011);
nor U5542 (N_5542,N_4119,N_4633);
and U5543 (N_5543,N_4573,N_4266);
or U5544 (N_5544,N_4073,N_4490);
or U5545 (N_5545,N_4560,N_4776);
and U5546 (N_5546,N_4309,N_4934);
nand U5547 (N_5547,N_4684,N_4075);
xnor U5548 (N_5548,N_4603,N_4735);
and U5549 (N_5549,N_4379,N_4676);
nor U5550 (N_5550,N_4689,N_4000);
or U5551 (N_5551,N_4552,N_4495);
or U5552 (N_5552,N_4171,N_4858);
or U5553 (N_5553,N_4787,N_4850);
nand U5554 (N_5554,N_4468,N_4932);
and U5555 (N_5555,N_4603,N_4032);
nand U5556 (N_5556,N_4157,N_4812);
xnor U5557 (N_5557,N_4715,N_4548);
and U5558 (N_5558,N_4236,N_4696);
xor U5559 (N_5559,N_4666,N_4826);
xnor U5560 (N_5560,N_4600,N_4220);
xor U5561 (N_5561,N_4701,N_4803);
nand U5562 (N_5562,N_4052,N_4173);
or U5563 (N_5563,N_4740,N_4039);
or U5564 (N_5564,N_4035,N_4045);
xor U5565 (N_5565,N_4482,N_4619);
xnor U5566 (N_5566,N_4625,N_4571);
and U5567 (N_5567,N_4654,N_4426);
or U5568 (N_5568,N_4495,N_4035);
or U5569 (N_5569,N_4288,N_4304);
xor U5570 (N_5570,N_4659,N_4586);
xnor U5571 (N_5571,N_4962,N_4586);
nand U5572 (N_5572,N_4054,N_4947);
xnor U5573 (N_5573,N_4718,N_4758);
nor U5574 (N_5574,N_4581,N_4908);
xnor U5575 (N_5575,N_4689,N_4928);
nor U5576 (N_5576,N_4918,N_4558);
nor U5577 (N_5577,N_4680,N_4836);
xnor U5578 (N_5578,N_4031,N_4386);
xor U5579 (N_5579,N_4667,N_4381);
and U5580 (N_5580,N_4173,N_4410);
nand U5581 (N_5581,N_4259,N_4696);
and U5582 (N_5582,N_4584,N_4164);
xnor U5583 (N_5583,N_4982,N_4190);
nor U5584 (N_5584,N_4097,N_4371);
nand U5585 (N_5585,N_4597,N_4462);
nand U5586 (N_5586,N_4820,N_4165);
xnor U5587 (N_5587,N_4375,N_4047);
and U5588 (N_5588,N_4343,N_4640);
nor U5589 (N_5589,N_4179,N_4670);
and U5590 (N_5590,N_4177,N_4841);
nor U5591 (N_5591,N_4821,N_4098);
and U5592 (N_5592,N_4870,N_4589);
nand U5593 (N_5593,N_4598,N_4988);
xor U5594 (N_5594,N_4540,N_4789);
or U5595 (N_5595,N_4748,N_4342);
xor U5596 (N_5596,N_4853,N_4849);
or U5597 (N_5597,N_4782,N_4663);
nand U5598 (N_5598,N_4061,N_4468);
or U5599 (N_5599,N_4274,N_4462);
and U5600 (N_5600,N_4797,N_4531);
and U5601 (N_5601,N_4890,N_4505);
nand U5602 (N_5602,N_4971,N_4978);
or U5603 (N_5603,N_4145,N_4485);
or U5604 (N_5604,N_4378,N_4271);
nor U5605 (N_5605,N_4066,N_4908);
nor U5606 (N_5606,N_4680,N_4909);
and U5607 (N_5607,N_4140,N_4272);
nand U5608 (N_5608,N_4376,N_4541);
and U5609 (N_5609,N_4100,N_4835);
or U5610 (N_5610,N_4269,N_4496);
nand U5611 (N_5611,N_4205,N_4384);
or U5612 (N_5612,N_4888,N_4169);
nand U5613 (N_5613,N_4078,N_4906);
and U5614 (N_5614,N_4508,N_4910);
nand U5615 (N_5615,N_4504,N_4765);
nor U5616 (N_5616,N_4716,N_4772);
xor U5617 (N_5617,N_4250,N_4810);
nand U5618 (N_5618,N_4459,N_4285);
or U5619 (N_5619,N_4142,N_4294);
nor U5620 (N_5620,N_4672,N_4793);
nor U5621 (N_5621,N_4114,N_4921);
xnor U5622 (N_5622,N_4516,N_4675);
and U5623 (N_5623,N_4998,N_4124);
nand U5624 (N_5624,N_4878,N_4378);
or U5625 (N_5625,N_4261,N_4500);
nor U5626 (N_5626,N_4903,N_4524);
nand U5627 (N_5627,N_4978,N_4497);
xor U5628 (N_5628,N_4157,N_4728);
nand U5629 (N_5629,N_4665,N_4953);
xor U5630 (N_5630,N_4646,N_4656);
nand U5631 (N_5631,N_4570,N_4685);
nand U5632 (N_5632,N_4033,N_4741);
nor U5633 (N_5633,N_4181,N_4139);
or U5634 (N_5634,N_4376,N_4868);
or U5635 (N_5635,N_4090,N_4770);
xnor U5636 (N_5636,N_4031,N_4546);
or U5637 (N_5637,N_4029,N_4926);
or U5638 (N_5638,N_4227,N_4700);
or U5639 (N_5639,N_4084,N_4171);
and U5640 (N_5640,N_4268,N_4265);
or U5641 (N_5641,N_4464,N_4772);
or U5642 (N_5642,N_4074,N_4007);
xor U5643 (N_5643,N_4968,N_4319);
xor U5644 (N_5644,N_4953,N_4371);
and U5645 (N_5645,N_4512,N_4171);
nor U5646 (N_5646,N_4307,N_4638);
nor U5647 (N_5647,N_4063,N_4784);
and U5648 (N_5648,N_4308,N_4977);
or U5649 (N_5649,N_4161,N_4163);
xnor U5650 (N_5650,N_4064,N_4979);
and U5651 (N_5651,N_4990,N_4329);
nor U5652 (N_5652,N_4478,N_4128);
nor U5653 (N_5653,N_4799,N_4094);
xor U5654 (N_5654,N_4535,N_4965);
nor U5655 (N_5655,N_4792,N_4285);
and U5656 (N_5656,N_4669,N_4490);
xor U5657 (N_5657,N_4636,N_4614);
nand U5658 (N_5658,N_4088,N_4192);
nor U5659 (N_5659,N_4673,N_4141);
nand U5660 (N_5660,N_4111,N_4207);
nand U5661 (N_5661,N_4987,N_4957);
nand U5662 (N_5662,N_4704,N_4746);
xnor U5663 (N_5663,N_4482,N_4935);
nor U5664 (N_5664,N_4989,N_4508);
or U5665 (N_5665,N_4221,N_4804);
or U5666 (N_5666,N_4230,N_4894);
nor U5667 (N_5667,N_4298,N_4861);
or U5668 (N_5668,N_4968,N_4419);
and U5669 (N_5669,N_4671,N_4805);
or U5670 (N_5670,N_4272,N_4929);
nand U5671 (N_5671,N_4406,N_4318);
xnor U5672 (N_5672,N_4595,N_4096);
xnor U5673 (N_5673,N_4018,N_4718);
xnor U5674 (N_5674,N_4176,N_4422);
nand U5675 (N_5675,N_4503,N_4225);
xor U5676 (N_5676,N_4139,N_4437);
and U5677 (N_5677,N_4191,N_4498);
xor U5678 (N_5678,N_4700,N_4129);
xor U5679 (N_5679,N_4844,N_4720);
and U5680 (N_5680,N_4662,N_4900);
xor U5681 (N_5681,N_4690,N_4025);
xor U5682 (N_5682,N_4548,N_4839);
or U5683 (N_5683,N_4989,N_4479);
nand U5684 (N_5684,N_4393,N_4558);
or U5685 (N_5685,N_4979,N_4384);
nor U5686 (N_5686,N_4474,N_4071);
nor U5687 (N_5687,N_4684,N_4776);
xor U5688 (N_5688,N_4286,N_4349);
nor U5689 (N_5689,N_4201,N_4446);
and U5690 (N_5690,N_4186,N_4387);
nand U5691 (N_5691,N_4944,N_4166);
and U5692 (N_5692,N_4268,N_4422);
and U5693 (N_5693,N_4938,N_4684);
or U5694 (N_5694,N_4445,N_4466);
nor U5695 (N_5695,N_4914,N_4088);
nor U5696 (N_5696,N_4693,N_4174);
xor U5697 (N_5697,N_4475,N_4048);
nand U5698 (N_5698,N_4522,N_4267);
xnor U5699 (N_5699,N_4619,N_4137);
and U5700 (N_5700,N_4257,N_4926);
or U5701 (N_5701,N_4320,N_4411);
and U5702 (N_5702,N_4208,N_4094);
xor U5703 (N_5703,N_4135,N_4077);
nor U5704 (N_5704,N_4515,N_4315);
or U5705 (N_5705,N_4277,N_4073);
xnor U5706 (N_5706,N_4641,N_4001);
and U5707 (N_5707,N_4331,N_4656);
nor U5708 (N_5708,N_4934,N_4547);
xnor U5709 (N_5709,N_4882,N_4956);
and U5710 (N_5710,N_4261,N_4707);
and U5711 (N_5711,N_4791,N_4464);
and U5712 (N_5712,N_4043,N_4261);
or U5713 (N_5713,N_4401,N_4831);
or U5714 (N_5714,N_4812,N_4702);
nor U5715 (N_5715,N_4511,N_4196);
or U5716 (N_5716,N_4801,N_4251);
or U5717 (N_5717,N_4153,N_4208);
nand U5718 (N_5718,N_4581,N_4114);
nor U5719 (N_5719,N_4403,N_4802);
nor U5720 (N_5720,N_4258,N_4627);
xnor U5721 (N_5721,N_4388,N_4877);
or U5722 (N_5722,N_4155,N_4266);
or U5723 (N_5723,N_4576,N_4539);
and U5724 (N_5724,N_4767,N_4191);
nor U5725 (N_5725,N_4671,N_4722);
xnor U5726 (N_5726,N_4798,N_4815);
and U5727 (N_5727,N_4787,N_4250);
nor U5728 (N_5728,N_4470,N_4294);
nor U5729 (N_5729,N_4533,N_4009);
xnor U5730 (N_5730,N_4038,N_4217);
and U5731 (N_5731,N_4735,N_4848);
nand U5732 (N_5732,N_4117,N_4407);
nand U5733 (N_5733,N_4482,N_4503);
nor U5734 (N_5734,N_4248,N_4334);
nor U5735 (N_5735,N_4836,N_4133);
nor U5736 (N_5736,N_4418,N_4073);
and U5737 (N_5737,N_4095,N_4953);
nor U5738 (N_5738,N_4406,N_4887);
xnor U5739 (N_5739,N_4434,N_4184);
nor U5740 (N_5740,N_4910,N_4312);
nor U5741 (N_5741,N_4546,N_4553);
xor U5742 (N_5742,N_4252,N_4539);
and U5743 (N_5743,N_4129,N_4942);
xor U5744 (N_5744,N_4444,N_4834);
nor U5745 (N_5745,N_4634,N_4560);
nand U5746 (N_5746,N_4648,N_4546);
nor U5747 (N_5747,N_4869,N_4089);
and U5748 (N_5748,N_4300,N_4603);
nand U5749 (N_5749,N_4001,N_4276);
xor U5750 (N_5750,N_4587,N_4108);
and U5751 (N_5751,N_4901,N_4502);
and U5752 (N_5752,N_4941,N_4536);
nand U5753 (N_5753,N_4045,N_4203);
or U5754 (N_5754,N_4957,N_4913);
nand U5755 (N_5755,N_4792,N_4281);
or U5756 (N_5756,N_4002,N_4828);
nor U5757 (N_5757,N_4428,N_4693);
nor U5758 (N_5758,N_4742,N_4216);
and U5759 (N_5759,N_4083,N_4891);
nand U5760 (N_5760,N_4568,N_4987);
nand U5761 (N_5761,N_4659,N_4523);
nand U5762 (N_5762,N_4515,N_4557);
nand U5763 (N_5763,N_4896,N_4605);
nor U5764 (N_5764,N_4307,N_4806);
and U5765 (N_5765,N_4955,N_4369);
xnor U5766 (N_5766,N_4590,N_4435);
nor U5767 (N_5767,N_4288,N_4401);
and U5768 (N_5768,N_4034,N_4785);
and U5769 (N_5769,N_4994,N_4937);
xnor U5770 (N_5770,N_4536,N_4251);
nand U5771 (N_5771,N_4257,N_4806);
and U5772 (N_5772,N_4372,N_4496);
xor U5773 (N_5773,N_4325,N_4700);
or U5774 (N_5774,N_4678,N_4253);
nor U5775 (N_5775,N_4493,N_4538);
nand U5776 (N_5776,N_4683,N_4507);
or U5777 (N_5777,N_4431,N_4861);
xnor U5778 (N_5778,N_4376,N_4749);
xnor U5779 (N_5779,N_4025,N_4887);
nand U5780 (N_5780,N_4040,N_4641);
nand U5781 (N_5781,N_4307,N_4634);
or U5782 (N_5782,N_4721,N_4825);
xor U5783 (N_5783,N_4979,N_4296);
nor U5784 (N_5784,N_4818,N_4480);
nand U5785 (N_5785,N_4016,N_4665);
and U5786 (N_5786,N_4687,N_4708);
nor U5787 (N_5787,N_4702,N_4626);
nand U5788 (N_5788,N_4265,N_4356);
nand U5789 (N_5789,N_4621,N_4595);
or U5790 (N_5790,N_4134,N_4953);
xnor U5791 (N_5791,N_4131,N_4090);
or U5792 (N_5792,N_4202,N_4907);
xor U5793 (N_5793,N_4131,N_4993);
xnor U5794 (N_5794,N_4365,N_4238);
or U5795 (N_5795,N_4994,N_4946);
and U5796 (N_5796,N_4088,N_4559);
nand U5797 (N_5797,N_4007,N_4302);
or U5798 (N_5798,N_4871,N_4065);
xnor U5799 (N_5799,N_4859,N_4164);
or U5800 (N_5800,N_4290,N_4906);
nand U5801 (N_5801,N_4174,N_4578);
nor U5802 (N_5802,N_4280,N_4129);
nor U5803 (N_5803,N_4310,N_4433);
nor U5804 (N_5804,N_4086,N_4287);
nor U5805 (N_5805,N_4581,N_4625);
nor U5806 (N_5806,N_4836,N_4937);
xnor U5807 (N_5807,N_4589,N_4170);
xnor U5808 (N_5808,N_4226,N_4613);
or U5809 (N_5809,N_4242,N_4080);
nand U5810 (N_5810,N_4510,N_4896);
or U5811 (N_5811,N_4826,N_4539);
nor U5812 (N_5812,N_4154,N_4871);
and U5813 (N_5813,N_4113,N_4102);
nor U5814 (N_5814,N_4970,N_4288);
nand U5815 (N_5815,N_4163,N_4832);
nand U5816 (N_5816,N_4954,N_4596);
or U5817 (N_5817,N_4258,N_4248);
xor U5818 (N_5818,N_4183,N_4315);
or U5819 (N_5819,N_4866,N_4751);
nor U5820 (N_5820,N_4583,N_4257);
nand U5821 (N_5821,N_4547,N_4214);
nor U5822 (N_5822,N_4526,N_4828);
nor U5823 (N_5823,N_4535,N_4817);
xnor U5824 (N_5824,N_4692,N_4299);
xor U5825 (N_5825,N_4686,N_4549);
or U5826 (N_5826,N_4882,N_4508);
nand U5827 (N_5827,N_4295,N_4910);
nor U5828 (N_5828,N_4105,N_4767);
xnor U5829 (N_5829,N_4169,N_4496);
xor U5830 (N_5830,N_4161,N_4549);
or U5831 (N_5831,N_4550,N_4875);
or U5832 (N_5832,N_4951,N_4433);
xnor U5833 (N_5833,N_4249,N_4552);
nand U5834 (N_5834,N_4960,N_4316);
xor U5835 (N_5835,N_4301,N_4733);
and U5836 (N_5836,N_4815,N_4417);
xor U5837 (N_5837,N_4218,N_4701);
nor U5838 (N_5838,N_4202,N_4774);
and U5839 (N_5839,N_4973,N_4316);
nand U5840 (N_5840,N_4816,N_4166);
xor U5841 (N_5841,N_4457,N_4289);
nor U5842 (N_5842,N_4913,N_4721);
nor U5843 (N_5843,N_4099,N_4936);
nor U5844 (N_5844,N_4344,N_4201);
and U5845 (N_5845,N_4344,N_4642);
nand U5846 (N_5846,N_4058,N_4614);
and U5847 (N_5847,N_4707,N_4811);
nand U5848 (N_5848,N_4937,N_4412);
nand U5849 (N_5849,N_4879,N_4260);
and U5850 (N_5850,N_4034,N_4342);
nand U5851 (N_5851,N_4766,N_4813);
and U5852 (N_5852,N_4806,N_4310);
nor U5853 (N_5853,N_4478,N_4977);
nor U5854 (N_5854,N_4657,N_4786);
or U5855 (N_5855,N_4678,N_4160);
or U5856 (N_5856,N_4094,N_4087);
and U5857 (N_5857,N_4102,N_4876);
and U5858 (N_5858,N_4585,N_4464);
and U5859 (N_5859,N_4348,N_4792);
xor U5860 (N_5860,N_4376,N_4045);
nand U5861 (N_5861,N_4884,N_4865);
xnor U5862 (N_5862,N_4589,N_4463);
nor U5863 (N_5863,N_4714,N_4676);
or U5864 (N_5864,N_4254,N_4815);
xnor U5865 (N_5865,N_4541,N_4971);
or U5866 (N_5866,N_4753,N_4517);
nor U5867 (N_5867,N_4455,N_4929);
nor U5868 (N_5868,N_4443,N_4562);
or U5869 (N_5869,N_4062,N_4683);
nor U5870 (N_5870,N_4152,N_4520);
nor U5871 (N_5871,N_4337,N_4771);
or U5872 (N_5872,N_4310,N_4187);
nand U5873 (N_5873,N_4944,N_4874);
nor U5874 (N_5874,N_4296,N_4072);
or U5875 (N_5875,N_4623,N_4153);
nor U5876 (N_5876,N_4279,N_4473);
and U5877 (N_5877,N_4123,N_4485);
or U5878 (N_5878,N_4548,N_4846);
nor U5879 (N_5879,N_4040,N_4979);
xor U5880 (N_5880,N_4443,N_4031);
and U5881 (N_5881,N_4425,N_4017);
nand U5882 (N_5882,N_4719,N_4992);
nor U5883 (N_5883,N_4087,N_4953);
or U5884 (N_5884,N_4361,N_4784);
or U5885 (N_5885,N_4327,N_4628);
xnor U5886 (N_5886,N_4880,N_4963);
and U5887 (N_5887,N_4557,N_4101);
nor U5888 (N_5888,N_4781,N_4683);
nand U5889 (N_5889,N_4384,N_4482);
xnor U5890 (N_5890,N_4841,N_4871);
and U5891 (N_5891,N_4339,N_4073);
or U5892 (N_5892,N_4819,N_4087);
nand U5893 (N_5893,N_4186,N_4965);
nand U5894 (N_5894,N_4012,N_4694);
nand U5895 (N_5895,N_4741,N_4745);
nor U5896 (N_5896,N_4160,N_4266);
nor U5897 (N_5897,N_4821,N_4119);
nand U5898 (N_5898,N_4147,N_4078);
nand U5899 (N_5899,N_4021,N_4465);
and U5900 (N_5900,N_4746,N_4440);
or U5901 (N_5901,N_4542,N_4297);
nor U5902 (N_5902,N_4061,N_4802);
nand U5903 (N_5903,N_4681,N_4995);
and U5904 (N_5904,N_4596,N_4552);
and U5905 (N_5905,N_4010,N_4577);
nand U5906 (N_5906,N_4810,N_4245);
or U5907 (N_5907,N_4927,N_4598);
or U5908 (N_5908,N_4860,N_4742);
xor U5909 (N_5909,N_4153,N_4211);
or U5910 (N_5910,N_4163,N_4805);
and U5911 (N_5911,N_4184,N_4098);
nor U5912 (N_5912,N_4872,N_4962);
and U5913 (N_5913,N_4321,N_4746);
xnor U5914 (N_5914,N_4378,N_4517);
nor U5915 (N_5915,N_4670,N_4875);
nand U5916 (N_5916,N_4569,N_4214);
nor U5917 (N_5917,N_4094,N_4870);
or U5918 (N_5918,N_4761,N_4464);
or U5919 (N_5919,N_4046,N_4579);
and U5920 (N_5920,N_4412,N_4706);
and U5921 (N_5921,N_4680,N_4819);
xnor U5922 (N_5922,N_4499,N_4111);
nor U5923 (N_5923,N_4700,N_4230);
nand U5924 (N_5924,N_4554,N_4494);
and U5925 (N_5925,N_4858,N_4961);
and U5926 (N_5926,N_4134,N_4714);
and U5927 (N_5927,N_4782,N_4781);
and U5928 (N_5928,N_4945,N_4562);
nor U5929 (N_5929,N_4596,N_4745);
xor U5930 (N_5930,N_4537,N_4157);
xnor U5931 (N_5931,N_4033,N_4069);
and U5932 (N_5932,N_4144,N_4102);
and U5933 (N_5933,N_4635,N_4206);
or U5934 (N_5934,N_4950,N_4358);
nand U5935 (N_5935,N_4495,N_4289);
or U5936 (N_5936,N_4374,N_4209);
nand U5937 (N_5937,N_4197,N_4789);
or U5938 (N_5938,N_4104,N_4502);
and U5939 (N_5939,N_4491,N_4583);
nand U5940 (N_5940,N_4818,N_4690);
nor U5941 (N_5941,N_4609,N_4349);
nand U5942 (N_5942,N_4631,N_4724);
xor U5943 (N_5943,N_4570,N_4259);
or U5944 (N_5944,N_4766,N_4769);
or U5945 (N_5945,N_4854,N_4541);
nand U5946 (N_5946,N_4466,N_4555);
nand U5947 (N_5947,N_4628,N_4392);
nand U5948 (N_5948,N_4471,N_4723);
nand U5949 (N_5949,N_4017,N_4343);
xor U5950 (N_5950,N_4182,N_4666);
or U5951 (N_5951,N_4036,N_4261);
xnor U5952 (N_5952,N_4172,N_4443);
and U5953 (N_5953,N_4718,N_4186);
or U5954 (N_5954,N_4669,N_4726);
xor U5955 (N_5955,N_4800,N_4853);
xor U5956 (N_5956,N_4875,N_4552);
and U5957 (N_5957,N_4937,N_4517);
xnor U5958 (N_5958,N_4361,N_4630);
and U5959 (N_5959,N_4820,N_4014);
nand U5960 (N_5960,N_4627,N_4222);
nand U5961 (N_5961,N_4853,N_4597);
nor U5962 (N_5962,N_4531,N_4242);
nor U5963 (N_5963,N_4291,N_4601);
and U5964 (N_5964,N_4987,N_4210);
and U5965 (N_5965,N_4627,N_4415);
nor U5966 (N_5966,N_4517,N_4117);
or U5967 (N_5967,N_4822,N_4349);
and U5968 (N_5968,N_4796,N_4776);
nand U5969 (N_5969,N_4941,N_4703);
nor U5970 (N_5970,N_4183,N_4253);
or U5971 (N_5971,N_4598,N_4423);
and U5972 (N_5972,N_4046,N_4146);
nor U5973 (N_5973,N_4013,N_4905);
and U5974 (N_5974,N_4880,N_4506);
or U5975 (N_5975,N_4715,N_4328);
nand U5976 (N_5976,N_4653,N_4401);
nor U5977 (N_5977,N_4610,N_4845);
xor U5978 (N_5978,N_4848,N_4182);
xnor U5979 (N_5979,N_4110,N_4552);
or U5980 (N_5980,N_4024,N_4283);
or U5981 (N_5981,N_4671,N_4581);
xor U5982 (N_5982,N_4936,N_4391);
nor U5983 (N_5983,N_4970,N_4233);
xnor U5984 (N_5984,N_4024,N_4046);
nor U5985 (N_5985,N_4730,N_4362);
nor U5986 (N_5986,N_4916,N_4795);
or U5987 (N_5987,N_4570,N_4819);
nand U5988 (N_5988,N_4990,N_4849);
nor U5989 (N_5989,N_4367,N_4023);
xor U5990 (N_5990,N_4994,N_4329);
and U5991 (N_5991,N_4074,N_4223);
nand U5992 (N_5992,N_4593,N_4453);
or U5993 (N_5993,N_4763,N_4717);
nand U5994 (N_5994,N_4375,N_4069);
nand U5995 (N_5995,N_4800,N_4303);
nor U5996 (N_5996,N_4429,N_4986);
and U5997 (N_5997,N_4424,N_4324);
xnor U5998 (N_5998,N_4928,N_4642);
or U5999 (N_5999,N_4119,N_4280);
nor U6000 (N_6000,N_5331,N_5481);
or U6001 (N_6001,N_5667,N_5322);
nor U6002 (N_6002,N_5855,N_5191);
and U6003 (N_6003,N_5278,N_5611);
and U6004 (N_6004,N_5868,N_5026);
nor U6005 (N_6005,N_5090,N_5174);
xor U6006 (N_6006,N_5081,N_5066);
xor U6007 (N_6007,N_5860,N_5872);
and U6008 (N_6008,N_5824,N_5939);
nor U6009 (N_6009,N_5114,N_5375);
nor U6010 (N_6010,N_5429,N_5753);
xnor U6011 (N_6011,N_5008,N_5875);
or U6012 (N_6012,N_5943,N_5615);
or U6013 (N_6013,N_5166,N_5165);
nand U6014 (N_6014,N_5188,N_5249);
nand U6015 (N_6015,N_5691,N_5258);
or U6016 (N_6016,N_5480,N_5305);
nor U6017 (N_6017,N_5313,N_5538);
nand U6018 (N_6018,N_5403,N_5514);
and U6019 (N_6019,N_5347,N_5612);
nand U6020 (N_6020,N_5454,N_5969);
nor U6021 (N_6021,N_5492,N_5862);
xnor U6022 (N_6022,N_5512,N_5938);
xor U6023 (N_6023,N_5948,N_5228);
nand U6024 (N_6024,N_5282,N_5326);
or U6025 (N_6025,N_5241,N_5685);
or U6026 (N_6026,N_5518,N_5925);
nand U6027 (N_6027,N_5646,N_5863);
nand U6028 (N_6028,N_5636,N_5741);
xor U6029 (N_6029,N_5884,N_5426);
and U6030 (N_6030,N_5537,N_5186);
xnor U6031 (N_6031,N_5441,N_5353);
and U6032 (N_6032,N_5694,N_5418);
or U6033 (N_6033,N_5276,N_5149);
nand U6034 (N_6034,N_5421,N_5910);
or U6035 (N_6035,N_5142,N_5742);
xor U6036 (N_6036,N_5665,N_5034);
xnor U6037 (N_6037,N_5124,N_5298);
nor U6038 (N_6038,N_5084,N_5865);
nor U6039 (N_6039,N_5401,N_5467);
or U6040 (N_6040,N_5195,N_5409);
nor U6041 (N_6041,N_5766,N_5462);
and U6042 (N_6042,N_5369,N_5787);
xor U6043 (N_6043,N_5912,N_5772);
or U6044 (N_6044,N_5755,N_5058);
nand U6045 (N_6045,N_5333,N_5083);
xnor U6046 (N_6046,N_5593,N_5745);
or U6047 (N_6047,N_5847,N_5926);
nand U6048 (N_6048,N_5966,N_5318);
nor U6049 (N_6049,N_5849,N_5352);
or U6050 (N_6050,N_5580,N_5343);
or U6051 (N_6051,N_5113,N_5569);
nor U6052 (N_6052,N_5754,N_5054);
and U6053 (N_6053,N_5351,N_5416);
or U6054 (N_6054,N_5128,N_5112);
and U6055 (N_6055,N_5460,N_5025);
xnor U6056 (N_6056,N_5103,N_5048);
or U6057 (N_6057,N_5233,N_5229);
nor U6058 (N_6058,N_5055,N_5422);
nand U6059 (N_6059,N_5820,N_5961);
and U6060 (N_6060,N_5695,N_5052);
xor U6061 (N_6061,N_5931,N_5744);
xnor U6062 (N_6062,N_5749,N_5704);
nor U6063 (N_6063,N_5159,N_5509);
nand U6064 (N_6064,N_5620,N_5002);
xor U6065 (N_6065,N_5334,N_5639);
or U6066 (N_6066,N_5899,N_5701);
or U6067 (N_6067,N_5486,N_5871);
or U6068 (N_6068,N_5136,N_5781);
and U6069 (N_6069,N_5041,N_5516);
xnor U6070 (N_6070,N_5354,N_5858);
xor U6071 (N_6071,N_5303,N_5271);
or U6072 (N_6072,N_5221,N_5402);
or U6073 (N_6073,N_5891,N_5212);
nor U6074 (N_6074,N_5545,N_5823);
or U6075 (N_6075,N_5914,N_5247);
and U6076 (N_6076,N_5867,N_5069);
xor U6077 (N_6077,N_5019,N_5153);
nand U6078 (N_6078,N_5385,N_5762);
xor U6079 (N_6079,N_5958,N_5094);
xor U6080 (N_6080,N_5707,N_5503);
nor U6081 (N_6081,N_5944,N_5976);
nor U6082 (N_6082,N_5987,N_5692);
nand U6083 (N_6083,N_5873,N_5489);
nor U6084 (N_6084,N_5582,N_5187);
nand U6085 (N_6085,N_5208,N_5295);
nor U6086 (N_6086,N_5556,N_5380);
and U6087 (N_6087,N_5184,N_5599);
or U6088 (N_6088,N_5382,N_5785);
and U6089 (N_6089,N_5164,N_5200);
nor U6090 (N_6090,N_5673,N_5606);
or U6091 (N_6091,N_5118,N_5534);
xnor U6092 (N_6092,N_5696,N_5363);
nand U6093 (N_6093,N_5230,N_5449);
nor U6094 (N_6094,N_5361,N_5622);
and U6095 (N_6095,N_5963,N_5199);
or U6096 (N_6096,N_5829,N_5493);
nor U6097 (N_6097,N_5260,N_5774);
nor U6098 (N_6098,N_5979,N_5138);
or U6099 (N_6099,N_5653,N_5381);
or U6100 (N_6100,N_5324,N_5728);
nand U6101 (N_6101,N_5876,N_5285);
xnor U6102 (N_6102,N_5670,N_5339);
and U6103 (N_6103,N_5491,N_5359);
and U6104 (N_6104,N_5548,N_5275);
and U6105 (N_6105,N_5951,N_5145);
or U6106 (N_6106,N_5777,N_5444);
nand U6107 (N_6107,N_5553,N_5714);
or U6108 (N_6108,N_5917,N_5344);
nand U6109 (N_6109,N_5049,N_5497);
or U6110 (N_6110,N_5367,N_5407);
xor U6111 (N_6111,N_5915,N_5879);
nand U6112 (N_6112,N_5342,N_5220);
and U6113 (N_6113,N_5908,N_5971);
xor U6114 (N_6114,N_5430,N_5869);
and U6115 (N_6115,N_5960,N_5182);
nor U6116 (N_6116,N_5818,N_5500);
nor U6117 (N_6117,N_5909,N_5368);
and U6118 (N_6118,N_5709,N_5924);
nand U6119 (N_6119,N_5323,N_5686);
and U6120 (N_6120,N_5137,N_5870);
or U6121 (N_6121,N_5716,N_5970);
xor U6122 (N_6122,N_5946,N_5307);
nor U6123 (N_6123,N_5732,N_5237);
nor U6124 (N_6124,N_5030,N_5340);
nand U6125 (N_6125,N_5294,N_5798);
nor U6126 (N_6126,N_5940,N_5074);
nand U6127 (N_6127,N_5115,N_5127);
xor U6128 (N_6128,N_5698,N_5578);
nor U6129 (N_6129,N_5614,N_5097);
or U6130 (N_6130,N_5110,N_5861);
nor U6131 (N_6131,N_5389,N_5736);
and U6132 (N_6132,N_5243,N_5280);
xnor U6133 (N_6133,N_5045,N_5125);
or U6134 (N_6134,N_5029,N_5794);
nor U6135 (N_6135,N_5757,N_5102);
nand U6136 (N_6136,N_5886,N_5256);
and U6137 (N_6137,N_5255,N_5445);
xor U6138 (N_6138,N_5618,N_5535);
nand U6139 (N_6139,N_5064,N_5994);
nand U6140 (N_6140,N_5597,N_5629);
xnor U6141 (N_6141,N_5116,N_5201);
or U6142 (N_6142,N_5037,N_5038);
nor U6143 (N_6143,N_5690,N_5522);
and U6144 (N_6144,N_5494,N_5532);
xnor U6145 (N_6145,N_5455,N_5120);
nor U6146 (N_6146,N_5495,N_5091);
nand U6147 (N_6147,N_5327,N_5645);
or U6148 (N_6148,N_5675,N_5998);
xor U6149 (N_6149,N_5895,N_5790);
xor U6150 (N_6150,N_5121,N_5376);
xnor U6151 (N_6151,N_5496,N_5205);
nor U6152 (N_6152,N_5050,N_5250);
nor U6153 (N_6153,N_5042,N_5404);
xor U6154 (N_6154,N_5773,N_5374);
and U6155 (N_6155,N_5711,N_5238);
or U6156 (N_6156,N_5185,N_5180);
and U6157 (N_6157,N_5160,N_5983);
nor U6158 (N_6158,N_5544,N_5498);
nand U6159 (N_6159,N_5217,N_5133);
and U6160 (N_6160,N_5688,N_5279);
xor U6161 (N_6161,N_5433,N_5542);
nor U6162 (N_6162,N_5130,N_5296);
xnor U6163 (N_6163,N_5651,N_5078);
xnor U6164 (N_6164,N_5077,N_5778);
and U6165 (N_6165,N_5490,N_5655);
xor U6166 (N_6166,N_5656,N_5851);
nand U6167 (N_6167,N_5056,N_5134);
nand U6168 (N_6168,N_5251,N_5316);
or U6169 (N_6169,N_5902,N_5458);
xor U6170 (N_6170,N_5517,N_5981);
xor U6171 (N_6171,N_5779,N_5477);
and U6172 (N_6172,N_5579,N_5093);
or U6173 (N_6173,N_5431,N_5436);
nand U6174 (N_6174,N_5274,N_5715);
nand U6175 (N_6175,N_5028,N_5650);
or U6176 (N_6176,N_5016,N_5395);
or U6177 (N_6177,N_5293,N_5482);
nand U6178 (N_6178,N_5668,N_5011);
and U6179 (N_6179,N_5239,N_5394);
and U6180 (N_6180,N_5904,N_5504);
or U6181 (N_6181,N_5747,N_5405);
xor U6182 (N_6182,N_5519,N_5759);
nand U6183 (N_6183,N_5272,N_5617);
nor U6184 (N_6184,N_5047,N_5649);
nand U6185 (N_6185,N_5758,N_5572);
nand U6186 (N_6186,N_5771,N_5007);
and U6187 (N_6187,N_5521,N_5219);
nand U6188 (N_6188,N_5246,N_5549);
nor U6189 (N_6189,N_5213,N_5834);
nand U6190 (N_6190,N_5240,N_5555);
xnor U6191 (N_6191,N_5515,N_5529);
or U6192 (N_6192,N_5877,N_5788);
nand U6193 (N_6193,N_5268,N_5725);
or U6194 (N_6194,N_5364,N_5738);
nor U6195 (N_6195,N_5562,N_5878);
or U6196 (N_6196,N_5459,N_5986);
nor U6197 (N_6197,N_5586,N_5892);
xnor U6198 (N_6198,N_5883,N_5306);
or U6199 (N_6199,N_5378,N_5658);
xnor U6200 (N_6200,N_5447,N_5852);
xor U6201 (N_6201,N_5839,N_5320);
xnor U6202 (N_6202,N_5513,N_5528);
and U6203 (N_6203,N_5793,N_5705);
nor U6204 (N_6204,N_5721,N_5487);
and U6205 (N_6205,N_5581,N_5393);
nor U6206 (N_6206,N_5400,N_5756);
xor U6207 (N_6207,N_5576,N_5536);
and U6208 (N_6208,N_5044,N_5977);
nor U6209 (N_6209,N_5065,N_5697);
and U6210 (N_6210,N_5484,N_5428);
and U6211 (N_6211,N_5842,N_5355);
or U6212 (N_6212,N_5710,N_5062);
xnor U6213 (N_6213,N_5464,N_5223);
xor U6214 (N_6214,N_5857,N_5760);
xnor U6215 (N_6215,N_5216,N_5499);
nor U6216 (N_6216,N_5634,N_5952);
or U6217 (N_6217,N_5501,N_5060);
or U6218 (N_6218,N_5328,N_5408);
nand U6219 (N_6219,N_5575,N_5973);
nand U6220 (N_6220,N_5630,N_5589);
nand U6221 (N_6221,N_5141,N_5360);
nor U6222 (N_6222,N_5901,N_5526);
nand U6223 (N_6223,N_5642,N_5613);
and U6224 (N_6224,N_5088,N_5123);
xor U6225 (N_6225,N_5392,N_5992);
or U6226 (N_6226,N_5261,N_5985);
xor U6227 (N_6227,N_5254,N_5154);
nor U6228 (N_6228,N_5903,N_5348);
xnor U6229 (N_6229,N_5804,N_5674);
xnor U6230 (N_6230,N_5232,N_5928);
nor U6231 (N_6231,N_5453,N_5432);
or U6232 (N_6232,N_5227,N_5706);
or U6233 (N_6233,N_5485,N_5263);
and U6234 (N_6234,N_5671,N_5505);
or U6235 (N_6235,N_5085,N_5267);
xnor U6236 (N_6236,N_5962,N_5846);
xor U6237 (N_6237,N_5662,N_5726);
xor U6238 (N_6238,N_5746,N_5838);
nand U6239 (N_6239,N_5168,N_5978);
nor U6240 (N_6240,N_5189,N_5853);
or U6241 (N_6241,N_5057,N_5967);
nor U6242 (N_6242,N_5737,N_5761);
and U6243 (N_6243,N_5812,N_5330);
xor U6244 (N_6244,N_5292,N_5748);
or U6245 (N_6245,N_5752,N_5601);
nand U6246 (N_6246,N_5291,N_5638);
xnor U6247 (N_6247,N_5273,N_5805);
and U6248 (N_6248,N_5730,N_5299);
nor U6249 (N_6249,N_5178,N_5033);
nand U6250 (N_6250,N_5425,N_5446);
or U6251 (N_6251,N_5616,N_5531);
nor U6252 (N_6252,N_5552,N_5561);
and U6253 (N_6253,N_5577,N_5996);
and U6254 (N_6254,N_5063,N_5071);
or U6255 (N_6255,N_5072,N_5724);
xnor U6256 (N_6256,N_5310,N_5682);
and U6257 (N_6257,N_5807,N_5396);
or U6258 (N_6258,N_5982,N_5397);
nand U6259 (N_6259,N_5043,N_5573);
or U6260 (N_6260,N_5419,N_5666);
nand U6261 (N_6261,N_5699,N_5218);
nand U6262 (N_6262,N_5678,N_5933);
xnor U6263 (N_6263,N_5564,N_5265);
and U6264 (N_6264,N_5897,N_5335);
and U6265 (N_6265,N_5073,N_5792);
nor U6266 (N_6266,N_5520,N_5635);
and U6267 (N_6267,N_5681,N_5006);
nand U6268 (N_6268,N_5739,N_5362);
xnor U6269 (N_6269,N_5676,N_5988);
nand U6270 (N_6270,N_5059,N_5632);
nand U6271 (N_6271,N_5702,N_5181);
nor U6272 (N_6272,N_5075,N_5286);
nand U6273 (N_6273,N_5743,N_5720);
and U6274 (N_6274,N_5470,N_5633);
nor U6275 (N_6275,N_5923,N_5341);
nor U6276 (N_6276,N_5816,N_5995);
xor U6277 (N_6277,N_5209,N_5874);
xor U6278 (N_6278,N_5398,N_5889);
nor U6279 (N_6279,N_5584,N_5448);
nand U6280 (N_6280,N_5104,N_5173);
or U6281 (N_6281,N_5196,N_5106);
or U6282 (N_6282,N_5111,N_5828);
or U6283 (N_6283,N_5974,N_5864);
nor U6284 (N_6284,N_5881,N_5587);
or U6285 (N_6285,N_5916,N_5021);
or U6286 (N_6286,N_5010,N_5559);
nor U6287 (N_6287,N_5770,N_5117);
or U6288 (N_6288,N_5171,N_5379);
xnor U6289 (N_6289,N_5595,N_5964);
or U6290 (N_6290,N_5972,N_5511);
nor U6291 (N_6291,N_5214,N_5070);
and U6292 (N_6292,N_5769,N_5604);
nor U6293 (N_6293,N_5859,N_5930);
or U6294 (N_6294,N_5197,N_5383);
and U6295 (N_6295,N_5882,N_5399);
xor U6296 (N_6296,N_5927,N_5162);
and U6297 (N_6297,N_5848,N_5169);
nor U6298 (N_6298,N_5051,N_5370);
nand U6299 (N_6299,N_5336,N_5894);
nor U6300 (N_6300,N_5596,N_5605);
xnor U6301 (N_6301,N_5621,N_5791);
nor U6302 (N_6302,N_5797,N_5092);
nor U6303 (N_6303,N_5411,N_5022);
nand U6304 (N_6304,N_5713,N_5896);
nand U6305 (N_6305,N_5032,N_5679);
nor U6306 (N_6306,N_5479,N_5570);
nor U6307 (N_6307,N_5936,N_5061);
xor U6308 (N_6308,N_5827,N_5795);
and U6309 (N_6309,N_5350,N_5955);
and U6310 (N_6310,N_5456,N_5819);
xnor U6311 (N_6311,N_5947,N_5833);
or U6312 (N_6312,N_5796,N_5101);
nor U6313 (N_6313,N_5937,N_5391);
nor U6314 (N_6314,N_5800,N_5959);
xor U6315 (N_6315,N_5832,N_5808);
nand U6316 (N_6316,N_5202,N_5954);
or U6317 (N_6317,N_5427,N_5161);
nor U6318 (N_6318,N_5317,N_5751);
nor U6319 (N_6319,N_5471,N_5566);
xor U6320 (N_6320,N_5727,N_5684);
or U6321 (N_6321,N_5680,N_5731);
nand U6322 (N_6322,N_5100,N_5990);
or U6323 (N_6323,N_5356,N_5004);
xnor U6324 (N_6324,N_5468,N_5235);
and U6325 (N_6325,N_5096,N_5358);
or U6326 (N_6326,N_5035,N_5371);
nand U6327 (N_6327,N_5508,N_5949);
and U6328 (N_6328,N_5139,N_5919);
nand U6329 (N_6329,N_5012,N_5300);
and U6330 (N_6330,N_5719,N_5469);
nand U6331 (N_6331,N_5211,N_5281);
and U6332 (N_6332,N_5906,N_5365);
nor U6333 (N_6333,N_5163,N_5693);
nand U6334 (N_6334,N_5890,N_5898);
xnor U6335 (N_6335,N_5424,N_5451);
or U6336 (N_6336,N_5473,N_5763);
and U6337 (N_6337,N_5068,N_5089);
xnor U6338 (N_6338,N_5015,N_5321);
xnor U6339 (N_6339,N_5373,N_5053);
and U6340 (N_6340,N_5266,N_5527);
nand U6341 (N_6341,N_5129,N_5836);
nand U6342 (N_6342,N_5929,N_5677);
nand U6343 (N_6343,N_5913,N_5193);
xor U6344 (N_6344,N_5588,N_5225);
nand U6345 (N_6345,N_5700,N_5108);
or U6346 (N_6346,N_5119,N_5357);
xor U6347 (N_6347,N_5099,N_5253);
and U6348 (N_6348,N_5231,N_5813);
nand U6349 (N_6349,N_5712,N_5703);
and U6350 (N_6350,N_5014,N_5502);
nor U6351 (N_6351,N_5603,N_5640);
nor U6352 (N_6352,N_5524,N_5297);
and U6353 (N_6353,N_5172,N_5269);
nand U6354 (N_6354,N_5277,N_5020);
nor U6355 (N_6355,N_5067,N_5417);
nor U6356 (N_6356,N_5017,N_5786);
and U6357 (N_6357,N_5594,N_5289);
nand U6358 (N_6358,N_5845,N_5483);
nor U6359 (N_6359,N_5717,N_5920);
and U6360 (N_6360,N_5844,N_5003);
and U6361 (N_6361,N_5264,N_5461);
or U6362 (N_6362,N_5372,N_5406);
nor U6363 (N_6363,N_5325,N_5236);
xnor U6364 (N_6364,N_5087,N_5013);
nand U6365 (N_6365,N_5510,N_5539);
and U6366 (N_6366,N_5175,N_5183);
nand U6367 (N_6367,N_5387,N_5377);
and U6368 (N_6368,N_5784,N_5132);
and U6369 (N_6369,N_5095,N_5652);
xor U6370 (N_6370,N_5854,N_5583);
and U6371 (N_6371,N_5571,N_5301);
nor U6372 (N_6372,N_5148,N_5563);
xnor U6373 (N_6373,N_5957,N_5776);
nor U6374 (N_6374,N_5222,N_5574);
and U6375 (N_6375,N_5598,N_5474);
and U6376 (N_6376,N_5866,N_5507);
nor U6377 (N_6377,N_5567,N_5911);
xnor U6378 (N_6378,N_5143,N_5657);
and U6379 (N_6379,N_5435,N_5329);
xnor U6380 (N_6380,N_5669,N_5031);
and U6381 (N_6381,N_5105,N_5506);
nor U6382 (N_6382,N_5304,N_5244);
or U6383 (N_6383,N_5830,N_5659);
or U6384 (N_6384,N_5607,N_5591);
nor U6385 (N_6385,N_5144,N_5600);
xnor U6386 (N_6386,N_5346,N_5345);
nand U6387 (N_6387,N_5809,N_5131);
and U6388 (N_6388,N_5107,N_5672);
xor U6389 (N_6389,N_5609,N_5158);
and U6390 (N_6390,N_5475,N_5687);
xor U6391 (N_6391,N_5437,N_5547);
nand U6392 (N_6392,N_5953,N_5817);
nand U6393 (N_6393,N_5815,N_5980);
nor U6394 (N_6394,N_5440,N_5643);
nor U6395 (N_6395,N_5729,N_5789);
and U6396 (N_6396,N_5525,N_5146);
or U6397 (N_6397,N_5177,N_5005);
nor U6398 (N_6398,N_5245,N_5631);
xnor U6399 (N_6399,N_5999,N_5624);
nand U6400 (N_6400,N_5248,N_5689);
and U6401 (N_6401,N_5541,N_5989);
or U6402 (N_6402,N_5592,N_5893);
nor U6403 (N_6403,N_5626,N_5001);
xnor U6404 (N_6404,N_5991,N_5628);
or U6405 (N_6405,N_5558,N_5488);
or U6406 (N_6406,N_5109,N_5557);
nand U6407 (N_6407,N_5024,N_5811);
xnor U6408 (N_6408,N_5841,N_5550);
nand U6409 (N_6409,N_5434,N_5147);
nand U6410 (N_6410,N_5523,N_5224);
or U6411 (N_6411,N_5637,N_5465);
or U6412 (N_6412,N_5450,N_5801);
nand U6413 (N_6413,N_5625,N_5887);
xnor U6414 (N_6414,N_5956,N_5152);
nand U6415 (N_6415,N_5082,N_5009);
or U6416 (N_6416,N_5036,N_5079);
and U6417 (N_6417,N_5206,N_5466);
xor U6418 (N_6418,N_5288,N_5386);
and U6419 (N_6419,N_5767,N_5905);
nor U6420 (N_6420,N_5565,N_5540);
nand U6421 (N_6421,N_5315,N_5941);
xnor U6422 (N_6422,N_5270,N_5803);
or U6423 (N_6423,N_5443,N_5661);
xor U6424 (N_6424,N_5332,N_5080);
nor U6425 (N_6425,N_5027,N_5900);
nand U6426 (N_6426,N_5806,N_5740);
nor U6427 (N_6427,N_5412,N_5568);
and U6428 (N_6428,N_5155,N_5627);
and U6429 (N_6429,N_5438,N_5610);
and U6430 (N_6430,N_5735,N_5623);
xor U6431 (N_6431,N_5683,N_5478);
xnor U6432 (N_6432,N_5945,N_5423);
or U6433 (N_6433,N_5856,N_5780);
or U6434 (N_6434,N_5608,N_5319);
xor U6435 (N_6435,N_5420,N_5039);
nor U6436 (N_6436,N_5157,N_5907);
nor U6437 (N_6437,N_5338,N_5156);
and U6438 (N_6438,N_5170,N_5198);
nor U6439 (N_6439,N_5259,N_5718);
xnor U6440 (N_6440,N_5918,N_5257);
nor U6441 (N_6441,N_5210,N_5641);
or U6442 (N_6442,N_5086,N_5993);
and U6443 (N_6443,N_5837,N_5708);
and U6444 (N_6444,N_5647,N_5843);
nor U6445 (N_6445,N_5533,N_5337);
xor U6446 (N_6446,N_5442,N_5850);
nor U6447 (N_6447,N_5975,N_5302);
xnor U6448 (N_6448,N_5921,N_5457);
nand U6449 (N_6449,N_5413,N_5194);
xor U6450 (N_6450,N_5734,N_5190);
nor U6451 (N_6451,N_5040,N_5046);
nand U6452 (N_6452,N_5775,N_5826);
xor U6453 (N_6453,N_5414,N_5415);
nand U6454 (N_6454,N_5965,N_5176);
xor U6455 (N_6455,N_5309,N_5722);
xor U6456 (N_6456,N_5590,N_5822);
nor U6457 (N_6457,N_5215,N_5750);
and U6458 (N_6458,N_5135,N_5452);
nand U6459 (N_6459,N_5410,N_5619);
nand U6460 (N_6460,N_5950,N_5076);
nor U6461 (N_6461,N_5551,N_5314);
nor U6462 (N_6462,N_5207,N_5098);
xnor U6463 (N_6463,N_5648,N_5840);
and U6464 (N_6464,N_5799,N_5810);
or U6465 (N_6465,N_5126,N_5723);
and U6466 (N_6466,N_5234,N_5765);
or U6467 (N_6467,N_5782,N_5167);
nor U6468 (N_6468,N_5825,N_5984);
or U6469 (N_6469,N_5935,N_5283);
and U6470 (N_6470,N_5140,N_5733);
and U6471 (N_6471,N_5151,N_5888);
and U6472 (N_6472,N_5814,N_5942);
xnor U6473 (N_6473,N_5543,N_5476);
and U6474 (N_6474,N_5602,N_5831);
nand U6475 (N_6475,N_5554,N_5663);
xor U6476 (N_6476,N_5122,N_5000);
and U6477 (N_6477,N_5366,N_5934);
xnor U6478 (N_6478,N_5472,N_5997);
xnor U6479 (N_6479,N_5546,N_5880);
nor U6480 (N_6480,N_5585,N_5644);
and U6481 (N_6481,N_5764,N_5179);
nor U6482 (N_6482,N_5018,N_5932);
xnor U6483 (N_6483,N_5192,N_5654);
nand U6484 (N_6484,N_5311,N_5242);
and U6485 (N_6485,N_5390,N_5262);
xor U6486 (N_6486,N_5388,N_5349);
or U6487 (N_6487,N_5821,N_5287);
nor U6488 (N_6488,N_5660,N_5226);
nor U6489 (N_6489,N_5768,N_5968);
and U6490 (N_6490,N_5203,N_5802);
xnor U6491 (N_6491,N_5252,N_5150);
and U6492 (N_6492,N_5308,N_5783);
or U6493 (N_6493,N_5384,N_5530);
nand U6494 (N_6494,N_5922,N_5284);
or U6495 (N_6495,N_5463,N_5023);
nand U6496 (N_6496,N_5664,N_5312);
nor U6497 (N_6497,N_5204,N_5439);
nor U6498 (N_6498,N_5290,N_5885);
xor U6499 (N_6499,N_5560,N_5835);
and U6500 (N_6500,N_5882,N_5590);
xor U6501 (N_6501,N_5198,N_5219);
and U6502 (N_6502,N_5002,N_5382);
and U6503 (N_6503,N_5664,N_5816);
xor U6504 (N_6504,N_5257,N_5818);
nand U6505 (N_6505,N_5359,N_5523);
nand U6506 (N_6506,N_5948,N_5853);
xnor U6507 (N_6507,N_5909,N_5102);
or U6508 (N_6508,N_5317,N_5932);
or U6509 (N_6509,N_5957,N_5601);
xnor U6510 (N_6510,N_5487,N_5912);
nor U6511 (N_6511,N_5126,N_5714);
xnor U6512 (N_6512,N_5039,N_5271);
xnor U6513 (N_6513,N_5767,N_5364);
and U6514 (N_6514,N_5887,N_5175);
nor U6515 (N_6515,N_5364,N_5034);
nand U6516 (N_6516,N_5121,N_5064);
nand U6517 (N_6517,N_5552,N_5613);
nand U6518 (N_6518,N_5512,N_5421);
nor U6519 (N_6519,N_5444,N_5074);
nand U6520 (N_6520,N_5700,N_5930);
nand U6521 (N_6521,N_5328,N_5025);
nor U6522 (N_6522,N_5726,N_5660);
nor U6523 (N_6523,N_5204,N_5247);
nand U6524 (N_6524,N_5281,N_5543);
or U6525 (N_6525,N_5002,N_5139);
nand U6526 (N_6526,N_5404,N_5088);
and U6527 (N_6527,N_5848,N_5342);
xnor U6528 (N_6528,N_5544,N_5384);
nor U6529 (N_6529,N_5296,N_5256);
xor U6530 (N_6530,N_5335,N_5359);
nand U6531 (N_6531,N_5636,N_5798);
and U6532 (N_6532,N_5715,N_5306);
or U6533 (N_6533,N_5829,N_5861);
nor U6534 (N_6534,N_5389,N_5096);
or U6535 (N_6535,N_5647,N_5017);
nand U6536 (N_6536,N_5747,N_5422);
nand U6537 (N_6537,N_5681,N_5588);
or U6538 (N_6538,N_5284,N_5511);
and U6539 (N_6539,N_5410,N_5590);
nand U6540 (N_6540,N_5577,N_5372);
nand U6541 (N_6541,N_5705,N_5455);
nor U6542 (N_6542,N_5873,N_5290);
and U6543 (N_6543,N_5463,N_5735);
xnor U6544 (N_6544,N_5699,N_5470);
nand U6545 (N_6545,N_5760,N_5853);
and U6546 (N_6546,N_5991,N_5091);
xor U6547 (N_6547,N_5084,N_5794);
xnor U6548 (N_6548,N_5567,N_5518);
nand U6549 (N_6549,N_5922,N_5262);
nor U6550 (N_6550,N_5519,N_5377);
nand U6551 (N_6551,N_5977,N_5184);
and U6552 (N_6552,N_5974,N_5593);
xnor U6553 (N_6553,N_5593,N_5151);
nand U6554 (N_6554,N_5289,N_5605);
xor U6555 (N_6555,N_5991,N_5672);
or U6556 (N_6556,N_5562,N_5213);
xnor U6557 (N_6557,N_5797,N_5485);
or U6558 (N_6558,N_5386,N_5074);
or U6559 (N_6559,N_5320,N_5292);
or U6560 (N_6560,N_5416,N_5192);
and U6561 (N_6561,N_5401,N_5082);
nand U6562 (N_6562,N_5042,N_5616);
and U6563 (N_6563,N_5319,N_5137);
nand U6564 (N_6564,N_5536,N_5093);
nand U6565 (N_6565,N_5246,N_5515);
xor U6566 (N_6566,N_5512,N_5172);
nor U6567 (N_6567,N_5189,N_5726);
nand U6568 (N_6568,N_5985,N_5417);
nor U6569 (N_6569,N_5041,N_5313);
nor U6570 (N_6570,N_5749,N_5813);
xnor U6571 (N_6571,N_5385,N_5145);
or U6572 (N_6572,N_5228,N_5741);
nand U6573 (N_6573,N_5594,N_5322);
nor U6574 (N_6574,N_5236,N_5423);
or U6575 (N_6575,N_5103,N_5675);
and U6576 (N_6576,N_5050,N_5186);
nor U6577 (N_6577,N_5256,N_5236);
xnor U6578 (N_6578,N_5238,N_5854);
xor U6579 (N_6579,N_5521,N_5826);
xnor U6580 (N_6580,N_5113,N_5141);
nand U6581 (N_6581,N_5551,N_5505);
nor U6582 (N_6582,N_5868,N_5967);
nor U6583 (N_6583,N_5087,N_5793);
and U6584 (N_6584,N_5762,N_5284);
nand U6585 (N_6585,N_5694,N_5662);
or U6586 (N_6586,N_5251,N_5859);
nor U6587 (N_6587,N_5379,N_5226);
nand U6588 (N_6588,N_5227,N_5399);
nor U6589 (N_6589,N_5943,N_5053);
nand U6590 (N_6590,N_5745,N_5515);
and U6591 (N_6591,N_5978,N_5820);
or U6592 (N_6592,N_5424,N_5368);
or U6593 (N_6593,N_5164,N_5564);
and U6594 (N_6594,N_5181,N_5212);
or U6595 (N_6595,N_5462,N_5370);
xor U6596 (N_6596,N_5682,N_5417);
nor U6597 (N_6597,N_5218,N_5059);
xor U6598 (N_6598,N_5311,N_5393);
and U6599 (N_6599,N_5993,N_5474);
or U6600 (N_6600,N_5029,N_5289);
and U6601 (N_6601,N_5258,N_5505);
and U6602 (N_6602,N_5241,N_5861);
xor U6603 (N_6603,N_5631,N_5421);
and U6604 (N_6604,N_5238,N_5990);
nand U6605 (N_6605,N_5065,N_5245);
nand U6606 (N_6606,N_5537,N_5826);
or U6607 (N_6607,N_5868,N_5962);
nand U6608 (N_6608,N_5382,N_5693);
or U6609 (N_6609,N_5640,N_5323);
nor U6610 (N_6610,N_5817,N_5226);
xor U6611 (N_6611,N_5050,N_5404);
nor U6612 (N_6612,N_5430,N_5590);
nor U6613 (N_6613,N_5744,N_5789);
or U6614 (N_6614,N_5508,N_5879);
xor U6615 (N_6615,N_5742,N_5199);
xor U6616 (N_6616,N_5521,N_5801);
xnor U6617 (N_6617,N_5758,N_5977);
xor U6618 (N_6618,N_5391,N_5583);
xor U6619 (N_6619,N_5984,N_5596);
nor U6620 (N_6620,N_5566,N_5480);
or U6621 (N_6621,N_5112,N_5481);
nor U6622 (N_6622,N_5535,N_5613);
xnor U6623 (N_6623,N_5687,N_5612);
xor U6624 (N_6624,N_5633,N_5709);
nand U6625 (N_6625,N_5958,N_5919);
nand U6626 (N_6626,N_5969,N_5079);
xor U6627 (N_6627,N_5101,N_5768);
and U6628 (N_6628,N_5647,N_5130);
nor U6629 (N_6629,N_5386,N_5867);
or U6630 (N_6630,N_5795,N_5480);
xor U6631 (N_6631,N_5317,N_5992);
xor U6632 (N_6632,N_5151,N_5670);
or U6633 (N_6633,N_5821,N_5920);
nor U6634 (N_6634,N_5777,N_5653);
xnor U6635 (N_6635,N_5934,N_5030);
and U6636 (N_6636,N_5892,N_5533);
nand U6637 (N_6637,N_5067,N_5880);
nand U6638 (N_6638,N_5771,N_5043);
nor U6639 (N_6639,N_5495,N_5875);
nand U6640 (N_6640,N_5839,N_5341);
nand U6641 (N_6641,N_5635,N_5026);
and U6642 (N_6642,N_5826,N_5907);
and U6643 (N_6643,N_5816,N_5321);
or U6644 (N_6644,N_5191,N_5033);
nor U6645 (N_6645,N_5624,N_5168);
and U6646 (N_6646,N_5557,N_5239);
xor U6647 (N_6647,N_5840,N_5308);
xor U6648 (N_6648,N_5265,N_5252);
nor U6649 (N_6649,N_5211,N_5755);
nor U6650 (N_6650,N_5292,N_5418);
nand U6651 (N_6651,N_5270,N_5962);
and U6652 (N_6652,N_5109,N_5449);
nor U6653 (N_6653,N_5131,N_5584);
nor U6654 (N_6654,N_5691,N_5151);
or U6655 (N_6655,N_5636,N_5155);
or U6656 (N_6656,N_5937,N_5593);
and U6657 (N_6657,N_5674,N_5715);
or U6658 (N_6658,N_5178,N_5281);
nand U6659 (N_6659,N_5674,N_5208);
nor U6660 (N_6660,N_5644,N_5611);
nand U6661 (N_6661,N_5192,N_5297);
or U6662 (N_6662,N_5222,N_5296);
and U6663 (N_6663,N_5131,N_5555);
and U6664 (N_6664,N_5807,N_5260);
or U6665 (N_6665,N_5856,N_5384);
nand U6666 (N_6666,N_5509,N_5980);
nor U6667 (N_6667,N_5232,N_5756);
xnor U6668 (N_6668,N_5844,N_5445);
xnor U6669 (N_6669,N_5213,N_5700);
or U6670 (N_6670,N_5760,N_5318);
or U6671 (N_6671,N_5347,N_5084);
nand U6672 (N_6672,N_5157,N_5890);
nand U6673 (N_6673,N_5085,N_5887);
and U6674 (N_6674,N_5442,N_5853);
nor U6675 (N_6675,N_5741,N_5429);
and U6676 (N_6676,N_5566,N_5784);
and U6677 (N_6677,N_5183,N_5304);
and U6678 (N_6678,N_5327,N_5509);
xnor U6679 (N_6679,N_5760,N_5200);
xor U6680 (N_6680,N_5694,N_5777);
or U6681 (N_6681,N_5523,N_5936);
xnor U6682 (N_6682,N_5712,N_5394);
xnor U6683 (N_6683,N_5537,N_5086);
xor U6684 (N_6684,N_5881,N_5751);
nor U6685 (N_6685,N_5276,N_5417);
nand U6686 (N_6686,N_5445,N_5873);
nor U6687 (N_6687,N_5100,N_5858);
and U6688 (N_6688,N_5179,N_5066);
or U6689 (N_6689,N_5438,N_5007);
xnor U6690 (N_6690,N_5681,N_5906);
xnor U6691 (N_6691,N_5602,N_5078);
xor U6692 (N_6692,N_5875,N_5634);
nor U6693 (N_6693,N_5305,N_5676);
xor U6694 (N_6694,N_5330,N_5550);
nand U6695 (N_6695,N_5510,N_5043);
nand U6696 (N_6696,N_5598,N_5928);
nor U6697 (N_6697,N_5180,N_5685);
nand U6698 (N_6698,N_5435,N_5636);
or U6699 (N_6699,N_5030,N_5297);
xor U6700 (N_6700,N_5582,N_5451);
and U6701 (N_6701,N_5266,N_5959);
or U6702 (N_6702,N_5565,N_5652);
or U6703 (N_6703,N_5832,N_5804);
or U6704 (N_6704,N_5230,N_5002);
nor U6705 (N_6705,N_5514,N_5305);
nor U6706 (N_6706,N_5753,N_5778);
nor U6707 (N_6707,N_5436,N_5443);
and U6708 (N_6708,N_5414,N_5375);
or U6709 (N_6709,N_5190,N_5214);
and U6710 (N_6710,N_5133,N_5331);
or U6711 (N_6711,N_5329,N_5832);
nand U6712 (N_6712,N_5659,N_5389);
or U6713 (N_6713,N_5118,N_5970);
nor U6714 (N_6714,N_5019,N_5626);
or U6715 (N_6715,N_5002,N_5649);
or U6716 (N_6716,N_5627,N_5033);
xor U6717 (N_6717,N_5246,N_5431);
nand U6718 (N_6718,N_5123,N_5213);
xor U6719 (N_6719,N_5682,N_5505);
nor U6720 (N_6720,N_5942,N_5849);
and U6721 (N_6721,N_5182,N_5267);
nand U6722 (N_6722,N_5392,N_5566);
or U6723 (N_6723,N_5403,N_5894);
nor U6724 (N_6724,N_5144,N_5626);
xor U6725 (N_6725,N_5554,N_5776);
nor U6726 (N_6726,N_5425,N_5324);
nand U6727 (N_6727,N_5230,N_5317);
or U6728 (N_6728,N_5982,N_5583);
xor U6729 (N_6729,N_5982,N_5657);
or U6730 (N_6730,N_5313,N_5508);
xor U6731 (N_6731,N_5196,N_5897);
or U6732 (N_6732,N_5780,N_5942);
nand U6733 (N_6733,N_5517,N_5513);
nand U6734 (N_6734,N_5691,N_5731);
and U6735 (N_6735,N_5502,N_5683);
nand U6736 (N_6736,N_5759,N_5855);
and U6737 (N_6737,N_5999,N_5200);
xor U6738 (N_6738,N_5269,N_5136);
or U6739 (N_6739,N_5128,N_5334);
nor U6740 (N_6740,N_5030,N_5866);
nand U6741 (N_6741,N_5990,N_5651);
or U6742 (N_6742,N_5470,N_5065);
xor U6743 (N_6743,N_5126,N_5838);
or U6744 (N_6744,N_5725,N_5710);
or U6745 (N_6745,N_5791,N_5294);
and U6746 (N_6746,N_5720,N_5845);
nor U6747 (N_6747,N_5887,N_5113);
nor U6748 (N_6748,N_5027,N_5012);
or U6749 (N_6749,N_5447,N_5500);
nor U6750 (N_6750,N_5005,N_5651);
or U6751 (N_6751,N_5367,N_5440);
xor U6752 (N_6752,N_5638,N_5600);
xnor U6753 (N_6753,N_5129,N_5477);
nor U6754 (N_6754,N_5485,N_5123);
nand U6755 (N_6755,N_5321,N_5499);
and U6756 (N_6756,N_5175,N_5774);
and U6757 (N_6757,N_5251,N_5420);
or U6758 (N_6758,N_5096,N_5069);
nor U6759 (N_6759,N_5661,N_5608);
xor U6760 (N_6760,N_5841,N_5289);
xor U6761 (N_6761,N_5017,N_5212);
nor U6762 (N_6762,N_5675,N_5640);
nand U6763 (N_6763,N_5996,N_5249);
and U6764 (N_6764,N_5659,N_5861);
nor U6765 (N_6765,N_5008,N_5211);
or U6766 (N_6766,N_5717,N_5489);
nor U6767 (N_6767,N_5638,N_5075);
nand U6768 (N_6768,N_5202,N_5164);
nor U6769 (N_6769,N_5859,N_5799);
nand U6770 (N_6770,N_5868,N_5635);
nor U6771 (N_6771,N_5062,N_5564);
or U6772 (N_6772,N_5658,N_5063);
nand U6773 (N_6773,N_5123,N_5802);
nor U6774 (N_6774,N_5896,N_5383);
nor U6775 (N_6775,N_5709,N_5676);
xor U6776 (N_6776,N_5048,N_5030);
and U6777 (N_6777,N_5777,N_5229);
nor U6778 (N_6778,N_5755,N_5268);
and U6779 (N_6779,N_5113,N_5977);
nand U6780 (N_6780,N_5706,N_5299);
and U6781 (N_6781,N_5982,N_5149);
nor U6782 (N_6782,N_5585,N_5093);
nor U6783 (N_6783,N_5962,N_5182);
or U6784 (N_6784,N_5501,N_5837);
nor U6785 (N_6785,N_5970,N_5896);
xor U6786 (N_6786,N_5848,N_5019);
and U6787 (N_6787,N_5741,N_5651);
xor U6788 (N_6788,N_5133,N_5883);
and U6789 (N_6789,N_5621,N_5883);
nor U6790 (N_6790,N_5957,N_5613);
or U6791 (N_6791,N_5369,N_5424);
or U6792 (N_6792,N_5562,N_5048);
xor U6793 (N_6793,N_5195,N_5041);
and U6794 (N_6794,N_5827,N_5754);
nor U6795 (N_6795,N_5721,N_5809);
and U6796 (N_6796,N_5716,N_5598);
and U6797 (N_6797,N_5773,N_5329);
nor U6798 (N_6798,N_5604,N_5075);
xor U6799 (N_6799,N_5213,N_5324);
xnor U6800 (N_6800,N_5210,N_5082);
and U6801 (N_6801,N_5026,N_5439);
nand U6802 (N_6802,N_5987,N_5210);
or U6803 (N_6803,N_5933,N_5379);
and U6804 (N_6804,N_5609,N_5809);
and U6805 (N_6805,N_5457,N_5275);
or U6806 (N_6806,N_5941,N_5891);
nand U6807 (N_6807,N_5378,N_5818);
and U6808 (N_6808,N_5893,N_5743);
nand U6809 (N_6809,N_5600,N_5022);
nand U6810 (N_6810,N_5657,N_5226);
xnor U6811 (N_6811,N_5239,N_5249);
nor U6812 (N_6812,N_5158,N_5522);
and U6813 (N_6813,N_5734,N_5840);
nand U6814 (N_6814,N_5052,N_5899);
nand U6815 (N_6815,N_5656,N_5462);
or U6816 (N_6816,N_5330,N_5800);
xnor U6817 (N_6817,N_5500,N_5961);
nand U6818 (N_6818,N_5683,N_5729);
and U6819 (N_6819,N_5128,N_5589);
nor U6820 (N_6820,N_5265,N_5109);
or U6821 (N_6821,N_5276,N_5931);
xnor U6822 (N_6822,N_5563,N_5748);
nand U6823 (N_6823,N_5032,N_5151);
nand U6824 (N_6824,N_5453,N_5922);
nor U6825 (N_6825,N_5042,N_5409);
or U6826 (N_6826,N_5889,N_5753);
nand U6827 (N_6827,N_5646,N_5099);
xor U6828 (N_6828,N_5489,N_5274);
nor U6829 (N_6829,N_5582,N_5548);
or U6830 (N_6830,N_5602,N_5717);
nand U6831 (N_6831,N_5166,N_5754);
or U6832 (N_6832,N_5477,N_5365);
or U6833 (N_6833,N_5678,N_5400);
and U6834 (N_6834,N_5036,N_5785);
xor U6835 (N_6835,N_5298,N_5688);
or U6836 (N_6836,N_5385,N_5099);
or U6837 (N_6837,N_5087,N_5547);
nor U6838 (N_6838,N_5633,N_5817);
nand U6839 (N_6839,N_5993,N_5556);
or U6840 (N_6840,N_5766,N_5814);
nand U6841 (N_6841,N_5634,N_5944);
and U6842 (N_6842,N_5830,N_5988);
xor U6843 (N_6843,N_5723,N_5065);
or U6844 (N_6844,N_5105,N_5280);
and U6845 (N_6845,N_5727,N_5118);
and U6846 (N_6846,N_5396,N_5794);
nand U6847 (N_6847,N_5866,N_5050);
and U6848 (N_6848,N_5041,N_5631);
nand U6849 (N_6849,N_5877,N_5807);
nand U6850 (N_6850,N_5211,N_5920);
xnor U6851 (N_6851,N_5195,N_5189);
nor U6852 (N_6852,N_5105,N_5552);
nand U6853 (N_6853,N_5074,N_5425);
nor U6854 (N_6854,N_5694,N_5165);
nor U6855 (N_6855,N_5106,N_5153);
nor U6856 (N_6856,N_5898,N_5793);
xor U6857 (N_6857,N_5732,N_5833);
or U6858 (N_6858,N_5719,N_5007);
or U6859 (N_6859,N_5029,N_5689);
nor U6860 (N_6860,N_5691,N_5747);
and U6861 (N_6861,N_5302,N_5644);
nand U6862 (N_6862,N_5812,N_5514);
nand U6863 (N_6863,N_5405,N_5287);
and U6864 (N_6864,N_5640,N_5535);
and U6865 (N_6865,N_5787,N_5545);
or U6866 (N_6866,N_5682,N_5099);
or U6867 (N_6867,N_5467,N_5275);
nand U6868 (N_6868,N_5908,N_5473);
nand U6869 (N_6869,N_5141,N_5827);
or U6870 (N_6870,N_5368,N_5717);
xnor U6871 (N_6871,N_5607,N_5756);
nor U6872 (N_6872,N_5332,N_5457);
xnor U6873 (N_6873,N_5672,N_5634);
and U6874 (N_6874,N_5657,N_5449);
and U6875 (N_6875,N_5952,N_5658);
and U6876 (N_6876,N_5126,N_5929);
nand U6877 (N_6877,N_5374,N_5020);
or U6878 (N_6878,N_5714,N_5768);
and U6879 (N_6879,N_5126,N_5942);
or U6880 (N_6880,N_5908,N_5723);
nand U6881 (N_6881,N_5445,N_5932);
nand U6882 (N_6882,N_5596,N_5597);
and U6883 (N_6883,N_5598,N_5042);
and U6884 (N_6884,N_5284,N_5643);
or U6885 (N_6885,N_5220,N_5633);
and U6886 (N_6886,N_5132,N_5518);
xor U6887 (N_6887,N_5618,N_5769);
or U6888 (N_6888,N_5705,N_5411);
and U6889 (N_6889,N_5549,N_5510);
or U6890 (N_6890,N_5173,N_5364);
and U6891 (N_6891,N_5861,N_5571);
nor U6892 (N_6892,N_5665,N_5412);
xor U6893 (N_6893,N_5264,N_5094);
nand U6894 (N_6894,N_5594,N_5820);
and U6895 (N_6895,N_5736,N_5162);
nand U6896 (N_6896,N_5614,N_5713);
and U6897 (N_6897,N_5543,N_5519);
xnor U6898 (N_6898,N_5344,N_5188);
and U6899 (N_6899,N_5162,N_5918);
nor U6900 (N_6900,N_5964,N_5120);
nor U6901 (N_6901,N_5519,N_5522);
nor U6902 (N_6902,N_5115,N_5254);
and U6903 (N_6903,N_5906,N_5761);
xnor U6904 (N_6904,N_5562,N_5887);
nor U6905 (N_6905,N_5068,N_5551);
xnor U6906 (N_6906,N_5431,N_5770);
xor U6907 (N_6907,N_5190,N_5974);
xnor U6908 (N_6908,N_5069,N_5041);
xnor U6909 (N_6909,N_5477,N_5011);
or U6910 (N_6910,N_5169,N_5628);
and U6911 (N_6911,N_5232,N_5446);
xor U6912 (N_6912,N_5793,N_5506);
nand U6913 (N_6913,N_5185,N_5081);
nor U6914 (N_6914,N_5480,N_5051);
nand U6915 (N_6915,N_5095,N_5689);
nor U6916 (N_6916,N_5699,N_5501);
nor U6917 (N_6917,N_5087,N_5721);
and U6918 (N_6918,N_5059,N_5344);
and U6919 (N_6919,N_5065,N_5269);
xnor U6920 (N_6920,N_5155,N_5194);
and U6921 (N_6921,N_5695,N_5767);
xnor U6922 (N_6922,N_5687,N_5322);
xnor U6923 (N_6923,N_5375,N_5760);
or U6924 (N_6924,N_5780,N_5141);
and U6925 (N_6925,N_5156,N_5239);
nor U6926 (N_6926,N_5374,N_5510);
and U6927 (N_6927,N_5871,N_5576);
and U6928 (N_6928,N_5293,N_5474);
or U6929 (N_6929,N_5565,N_5401);
and U6930 (N_6930,N_5700,N_5620);
and U6931 (N_6931,N_5563,N_5431);
or U6932 (N_6932,N_5737,N_5109);
nor U6933 (N_6933,N_5954,N_5190);
xnor U6934 (N_6934,N_5925,N_5607);
and U6935 (N_6935,N_5567,N_5892);
nand U6936 (N_6936,N_5638,N_5296);
and U6937 (N_6937,N_5315,N_5530);
nor U6938 (N_6938,N_5998,N_5608);
nand U6939 (N_6939,N_5711,N_5584);
nor U6940 (N_6940,N_5500,N_5345);
nand U6941 (N_6941,N_5103,N_5098);
xnor U6942 (N_6942,N_5557,N_5488);
xor U6943 (N_6943,N_5216,N_5190);
xor U6944 (N_6944,N_5108,N_5948);
xnor U6945 (N_6945,N_5321,N_5360);
or U6946 (N_6946,N_5733,N_5324);
or U6947 (N_6947,N_5315,N_5556);
and U6948 (N_6948,N_5380,N_5976);
xnor U6949 (N_6949,N_5425,N_5461);
nor U6950 (N_6950,N_5913,N_5677);
xor U6951 (N_6951,N_5516,N_5548);
xor U6952 (N_6952,N_5890,N_5421);
and U6953 (N_6953,N_5534,N_5930);
or U6954 (N_6954,N_5193,N_5532);
nand U6955 (N_6955,N_5677,N_5037);
and U6956 (N_6956,N_5508,N_5944);
xor U6957 (N_6957,N_5158,N_5976);
xnor U6958 (N_6958,N_5598,N_5437);
nor U6959 (N_6959,N_5809,N_5379);
or U6960 (N_6960,N_5426,N_5258);
nor U6961 (N_6961,N_5854,N_5053);
xnor U6962 (N_6962,N_5177,N_5562);
nor U6963 (N_6963,N_5547,N_5872);
nor U6964 (N_6964,N_5405,N_5052);
and U6965 (N_6965,N_5491,N_5940);
nor U6966 (N_6966,N_5922,N_5921);
and U6967 (N_6967,N_5792,N_5212);
xor U6968 (N_6968,N_5195,N_5010);
xor U6969 (N_6969,N_5724,N_5044);
nand U6970 (N_6970,N_5660,N_5570);
or U6971 (N_6971,N_5649,N_5478);
and U6972 (N_6972,N_5353,N_5935);
nor U6973 (N_6973,N_5304,N_5983);
xor U6974 (N_6974,N_5307,N_5111);
or U6975 (N_6975,N_5256,N_5252);
xnor U6976 (N_6976,N_5927,N_5675);
xor U6977 (N_6977,N_5651,N_5530);
xnor U6978 (N_6978,N_5134,N_5916);
nor U6979 (N_6979,N_5095,N_5063);
xnor U6980 (N_6980,N_5128,N_5805);
and U6981 (N_6981,N_5869,N_5293);
nor U6982 (N_6982,N_5319,N_5218);
nor U6983 (N_6983,N_5997,N_5030);
and U6984 (N_6984,N_5768,N_5370);
xor U6985 (N_6985,N_5748,N_5879);
and U6986 (N_6986,N_5984,N_5767);
nand U6987 (N_6987,N_5632,N_5261);
nand U6988 (N_6988,N_5598,N_5776);
xor U6989 (N_6989,N_5857,N_5270);
nor U6990 (N_6990,N_5815,N_5160);
nand U6991 (N_6991,N_5775,N_5662);
and U6992 (N_6992,N_5057,N_5623);
nand U6993 (N_6993,N_5914,N_5597);
xor U6994 (N_6994,N_5183,N_5639);
or U6995 (N_6995,N_5148,N_5803);
and U6996 (N_6996,N_5620,N_5652);
nor U6997 (N_6997,N_5939,N_5523);
nor U6998 (N_6998,N_5262,N_5751);
nand U6999 (N_6999,N_5037,N_5763);
xnor U7000 (N_7000,N_6456,N_6263);
and U7001 (N_7001,N_6151,N_6753);
xor U7002 (N_7002,N_6642,N_6204);
xnor U7003 (N_7003,N_6691,N_6484);
nor U7004 (N_7004,N_6964,N_6703);
or U7005 (N_7005,N_6757,N_6390);
nand U7006 (N_7006,N_6354,N_6621);
nand U7007 (N_7007,N_6450,N_6277);
nor U7008 (N_7008,N_6178,N_6735);
nor U7009 (N_7009,N_6461,N_6377);
nand U7010 (N_7010,N_6304,N_6818);
nand U7011 (N_7011,N_6882,N_6474);
nand U7012 (N_7012,N_6466,N_6025);
nand U7013 (N_7013,N_6696,N_6939);
nor U7014 (N_7014,N_6519,N_6965);
nor U7015 (N_7015,N_6530,N_6901);
or U7016 (N_7016,N_6117,N_6660);
xnor U7017 (N_7017,N_6617,N_6306);
nand U7018 (N_7018,N_6294,N_6969);
nor U7019 (N_7019,N_6083,N_6813);
or U7020 (N_7020,N_6472,N_6995);
xnor U7021 (N_7021,N_6459,N_6315);
or U7022 (N_7022,N_6548,N_6942);
and U7023 (N_7023,N_6575,N_6047);
nand U7024 (N_7024,N_6455,N_6708);
or U7025 (N_7025,N_6234,N_6003);
and U7026 (N_7026,N_6400,N_6168);
nand U7027 (N_7027,N_6623,N_6994);
or U7028 (N_7028,N_6150,N_6787);
nor U7029 (N_7029,N_6470,N_6602);
nor U7030 (N_7030,N_6807,N_6038);
nand U7031 (N_7031,N_6560,N_6355);
or U7032 (N_7032,N_6092,N_6610);
or U7033 (N_7033,N_6608,N_6481);
xnor U7034 (N_7034,N_6944,N_6903);
or U7035 (N_7035,N_6358,N_6546);
nand U7036 (N_7036,N_6556,N_6177);
xor U7037 (N_7037,N_6430,N_6570);
nand U7038 (N_7038,N_6700,N_6926);
nor U7039 (N_7039,N_6588,N_6115);
nor U7040 (N_7040,N_6501,N_6085);
xor U7041 (N_7041,N_6561,N_6899);
or U7042 (N_7042,N_6462,N_6288);
nand U7043 (N_7043,N_6783,N_6884);
nand U7044 (N_7044,N_6376,N_6385);
nor U7045 (N_7045,N_6603,N_6246);
nand U7046 (N_7046,N_6191,N_6075);
and U7047 (N_7047,N_6488,N_6477);
and U7048 (N_7048,N_6834,N_6279);
or U7049 (N_7049,N_6322,N_6791);
nor U7050 (N_7050,N_6004,N_6070);
nor U7051 (N_7051,N_6058,N_6250);
xnor U7052 (N_7052,N_6665,N_6129);
nor U7053 (N_7053,N_6754,N_6479);
and U7054 (N_7054,N_6962,N_6482);
or U7055 (N_7055,N_6175,N_6051);
xnor U7056 (N_7056,N_6679,N_6024);
xor U7057 (N_7057,N_6021,N_6976);
nand U7058 (N_7058,N_6883,N_6521);
nor U7059 (N_7059,N_6821,N_6001);
nor U7060 (N_7060,N_6580,N_6532);
nand U7061 (N_7061,N_6871,N_6592);
and U7062 (N_7062,N_6208,N_6644);
nor U7063 (N_7063,N_6285,N_6291);
or U7064 (N_7064,N_6084,N_6153);
nor U7065 (N_7065,N_6956,N_6720);
nor U7066 (N_7066,N_6292,N_6030);
nor U7067 (N_7067,N_6724,N_6612);
or U7068 (N_7068,N_6431,N_6977);
or U7069 (N_7069,N_6205,N_6106);
nand U7070 (N_7070,N_6314,N_6303);
nor U7071 (N_7071,N_6138,N_6137);
nand U7072 (N_7072,N_6636,N_6081);
and U7073 (N_7073,N_6631,N_6023);
or U7074 (N_7074,N_6752,N_6067);
nor U7075 (N_7075,N_6607,N_6209);
xnor U7076 (N_7076,N_6054,N_6493);
xnor U7077 (N_7077,N_6173,N_6321);
and U7078 (N_7078,N_6330,N_6225);
nor U7079 (N_7079,N_6566,N_6310);
nand U7080 (N_7080,N_6780,N_6674);
and U7081 (N_7081,N_6991,N_6830);
xnor U7082 (N_7082,N_6522,N_6252);
and U7083 (N_7083,N_6931,N_6750);
or U7084 (N_7084,N_6904,N_6073);
xnor U7085 (N_7085,N_6859,N_6254);
nand U7086 (N_7086,N_6567,N_6378);
or U7087 (N_7087,N_6946,N_6971);
nor U7088 (N_7088,N_6542,N_6823);
nor U7089 (N_7089,N_6940,N_6874);
xor U7090 (N_7090,N_6202,N_6562);
nand U7091 (N_7091,N_6077,N_6917);
nor U7092 (N_7092,N_6244,N_6978);
and U7093 (N_7093,N_6436,N_6412);
xnor U7094 (N_7094,N_6258,N_6844);
and U7095 (N_7095,N_6913,N_6534);
nand U7096 (N_7096,N_6214,N_6076);
or U7097 (N_7097,N_6465,N_6808);
xor U7098 (N_7098,N_6798,N_6448);
and U7099 (N_7099,N_6606,N_6241);
nand U7100 (N_7100,N_6121,N_6941);
and U7101 (N_7101,N_6020,N_6900);
xor U7102 (N_7102,N_6949,N_6107);
xor U7103 (N_7103,N_6555,N_6184);
nand U7104 (N_7104,N_6505,N_6410);
or U7105 (N_7105,N_6549,N_6706);
nor U7106 (N_7106,N_6260,N_6773);
and U7107 (N_7107,N_6265,N_6007);
and U7108 (N_7108,N_6825,N_6654);
and U7109 (N_7109,N_6511,N_6622);
nor U7110 (N_7110,N_6719,N_6282);
and U7111 (N_7111,N_6272,N_6257);
or U7112 (N_7112,N_6768,N_6427);
or U7113 (N_7113,N_6704,N_6396);
nand U7114 (N_7114,N_6036,N_6537);
and U7115 (N_7115,N_6576,N_6332);
nor U7116 (N_7116,N_6953,N_6167);
and U7117 (N_7117,N_6335,N_6865);
xnor U7118 (N_7118,N_6127,N_6181);
or U7119 (N_7119,N_6498,N_6447);
or U7120 (N_7120,N_6952,N_6143);
nor U7121 (N_7121,N_6095,N_6919);
nor U7122 (N_7122,N_6895,N_6563);
xnor U7123 (N_7123,N_6437,N_6583);
nand U7124 (N_7124,N_6155,N_6223);
and U7125 (N_7125,N_6711,N_6341);
nor U7126 (N_7126,N_6990,N_6658);
xnor U7127 (N_7127,N_6048,N_6096);
or U7128 (N_7128,N_6347,N_6035);
xnor U7129 (N_7129,N_6433,N_6630);
xnor U7130 (N_7130,N_6662,N_6331);
and U7131 (N_7131,N_6170,N_6135);
and U7132 (N_7132,N_6782,N_6156);
nor U7133 (N_7133,N_6625,N_6862);
xor U7134 (N_7134,N_6579,N_6718);
xnor U7135 (N_7135,N_6774,N_6487);
xnor U7136 (N_7136,N_6682,N_6937);
and U7137 (N_7137,N_6795,N_6118);
and U7138 (N_7138,N_6984,N_6295);
nand U7139 (N_7139,N_6329,N_6681);
nor U7140 (N_7140,N_6515,N_6595);
or U7141 (N_7141,N_6896,N_6451);
or U7142 (N_7142,N_6283,N_6849);
and U7143 (N_7143,N_6478,N_6394);
nor U7144 (N_7144,N_6399,N_6226);
or U7145 (N_7145,N_6230,N_6827);
and U7146 (N_7146,N_6045,N_6222);
and U7147 (N_7147,N_6967,N_6756);
nand U7148 (N_7148,N_6163,N_6099);
nand U7149 (N_7149,N_6614,N_6317);
xnor U7150 (N_7150,N_6417,N_6559);
and U7151 (N_7151,N_6641,N_6728);
xor U7152 (N_7152,N_6227,N_6837);
xnor U7153 (N_7153,N_6235,N_6543);
nand U7154 (N_7154,N_6591,N_6932);
and U7155 (N_7155,N_6206,N_6116);
xnor U7156 (N_7156,N_6529,N_6471);
xnor U7157 (N_7157,N_6707,N_6078);
nand U7158 (N_7158,N_6790,N_6668);
nand U7159 (N_7159,N_6444,N_6594);
xor U7160 (N_7160,N_6912,N_6684);
and U7161 (N_7161,N_6908,N_6187);
nor U7162 (N_7162,N_6945,N_6819);
nand U7163 (N_7163,N_6368,N_6535);
nand U7164 (N_7164,N_6979,N_6179);
or U7165 (N_7165,N_6973,N_6388);
and U7166 (N_7166,N_6716,N_6403);
nor U7167 (N_7167,N_6460,N_6664);
nand U7168 (N_7168,N_6924,N_6892);
nor U7169 (N_7169,N_6087,N_6373);
nand U7170 (N_7170,N_6935,N_6613);
or U7171 (N_7171,N_6069,N_6350);
or U7172 (N_7172,N_6360,N_6936);
nor U7173 (N_7173,N_6928,N_6667);
or U7174 (N_7174,N_6144,N_6705);
nand U7175 (N_7175,N_6506,N_6278);
and U7176 (N_7176,N_6647,N_6564);
and U7177 (N_7177,N_6639,N_6723);
or U7178 (N_7178,N_6043,N_6324);
and U7179 (N_7179,N_6046,N_6822);
xor U7180 (N_7180,N_6996,N_6800);
or U7181 (N_7181,N_6041,N_6852);
nor U7182 (N_7182,N_6238,N_6133);
xor U7183 (N_7183,N_6803,N_6476);
xnor U7184 (N_7184,N_6503,N_6231);
or U7185 (N_7185,N_6497,N_6139);
xor U7186 (N_7186,N_6902,N_6446);
xor U7187 (N_7187,N_6270,N_6961);
nand U7188 (N_7188,N_6183,N_6652);
and U7189 (N_7189,N_6199,N_6290);
xor U7190 (N_7190,N_6981,N_6361);
or U7191 (N_7191,N_6404,N_6374);
or U7192 (N_7192,N_6551,N_6382);
nand U7193 (N_7193,N_6338,N_6611);
nand U7194 (N_7194,N_6366,N_6645);
nor U7195 (N_7195,N_6312,N_6055);
xor U7196 (N_7196,N_6197,N_6925);
or U7197 (N_7197,N_6655,N_6565);
and U7198 (N_7198,N_6624,N_6861);
nor U7199 (N_7199,N_6885,N_6228);
nand U7200 (N_7200,N_6469,N_6997);
nand U7201 (N_7201,N_6948,N_6810);
nor U7202 (N_7202,N_6022,N_6587);
nand U7203 (N_7203,N_6596,N_6261);
xor U7204 (N_7204,N_6186,N_6876);
and U7205 (N_7205,N_6300,N_6082);
or U7206 (N_7206,N_6142,N_6552);
xor U7207 (N_7207,N_6766,N_6402);
nor U7208 (N_7208,N_6445,N_6066);
and U7209 (N_7209,N_6453,N_6159);
nand U7210 (N_7210,N_6855,N_6112);
or U7211 (N_7211,N_6702,N_6605);
or U7212 (N_7212,N_6289,N_6425);
and U7213 (N_7213,N_6218,N_6353);
or U7214 (N_7214,N_6966,N_6216);
xnor U7215 (N_7215,N_6510,N_6590);
xor U7216 (N_7216,N_6856,N_6034);
nand U7217 (N_7217,N_6789,N_6369);
nor U7218 (N_7218,N_6989,N_6011);
nor U7219 (N_7219,N_6262,N_6348);
nor U7220 (N_7220,N_6547,N_6119);
or U7221 (N_7221,N_6898,N_6334);
and U7222 (N_7222,N_6748,N_6792);
or U7223 (N_7223,N_6864,N_6105);
or U7224 (N_7224,N_6922,N_6824);
xnor U7225 (N_7225,N_6166,N_6414);
or U7226 (N_7226,N_6713,N_6520);
xnor U7227 (N_7227,N_6508,N_6777);
xnor U7228 (N_7228,N_6835,N_6029);
or U7229 (N_7229,N_6710,N_6620);
and U7230 (N_7230,N_6909,N_6585);
or U7231 (N_7231,N_6749,N_6879);
and U7232 (N_7232,N_6714,N_6140);
and U7233 (N_7233,N_6751,N_6313);
nand U7234 (N_7234,N_6762,N_6485);
or U7235 (N_7235,N_6316,N_6598);
and U7236 (N_7236,N_6923,N_6027);
or U7237 (N_7237,N_6694,N_6632);
nor U7238 (N_7238,N_6514,N_6490);
xor U7239 (N_7239,N_6804,N_6089);
or U7240 (N_7240,N_6581,N_6097);
nor U7241 (N_7241,N_6379,N_6866);
or U7242 (N_7242,N_6729,N_6761);
or U7243 (N_7243,N_6820,N_6811);
and U7244 (N_7244,N_6242,N_6528);
or U7245 (N_7245,N_6554,N_6464);
or U7246 (N_7246,N_6851,N_6880);
nor U7247 (N_7247,N_6154,N_6165);
nor U7248 (N_7248,N_6217,N_6688);
xnor U7249 (N_7249,N_6806,N_6391);
xnor U7250 (N_7250,N_6421,N_6829);
nand U7251 (N_7251,N_6028,N_6088);
nor U7252 (N_7252,N_6286,N_6201);
nor U7253 (N_7253,N_6873,N_6571);
nor U7254 (N_7254,N_6409,N_6346);
and U7255 (N_7255,N_6068,N_6420);
nor U7256 (N_7256,N_6259,N_6693);
nand U7257 (N_7257,N_6669,N_6463);
xor U7258 (N_7258,N_6722,N_6299);
nor U7259 (N_7259,N_6816,N_6287);
nand U7260 (N_7260,N_6677,N_6149);
and U7261 (N_7261,N_6318,N_6527);
and U7262 (N_7262,N_6578,N_6675);
nor U7263 (N_7263,N_6507,N_6059);
and U7264 (N_7264,N_6429,N_6771);
and U7265 (N_7265,N_6267,N_6424);
xnor U7266 (N_7266,N_6185,N_6005);
or U7267 (N_7267,N_6999,N_6531);
xnor U7268 (N_7268,N_6843,N_6715);
nand U7269 (N_7269,N_6509,N_6525);
nand U7270 (N_7270,N_6232,N_6957);
nor U7271 (N_7271,N_6577,N_6943);
xor U7272 (N_7272,N_6114,N_6128);
nand U7273 (N_7273,N_6858,N_6040);
nor U7274 (N_7274,N_6689,N_6094);
nor U7275 (N_7275,N_6203,N_6363);
nor U7276 (N_7276,N_6039,N_6086);
xnor U7277 (N_7277,N_6890,N_6176);
xnor U7278 (N_7278,N_6817,N_6224);
or U7279 (N_7279,N_6921,N_6698);
xnor U7280 (N_7280,N_6877,N_6418);
nand U7281 (N_7281,N_6838,N_6502);
nand U7282 (N_7282,N_6545,N_6311);
and U7283 (N_7283,N_6635,N_6213);
and U7284 (N_7284,N_6008,N_6000);
or U7285 (N_7285,N_6916,N_6435);
nand U7286 (N_7286,N_6033,N_6247);
or U7287 (N_7287,N_6333,N_6695);
and U7288 (N_7288,N_6649,N_6539);
nand U7289 (N_7289,N_6933,N_6002);
nor U7290 (N_7290,N_6062,N_6255);
and U7291 (N_7291,N_6071,N_6572);
xnor U7292 (N_7292,N_6010,N_6875);
nor U7293 (N_7293,N_6440,N_6491);
nor U7294 (N_7294,N_6785,N_6383);
xor U7295 (N_7295,N_6918,N_6536);
or U7296 (N_7296,N_6443,N_6125);
nor U7297 (N_7297,N_6422,N_6275);
xor U7298 (N_7298,N_6124,N_6998);
nand U7299 (N_7299,N_6389,N_6986);
nand U7300 (N_7300,N_6738,N_6670);
and U7301 (N_7301,N_6721,N_6309);
xnor U7302 (N_7302,N_6626,N_6467);
nor U7303 (N_7303,N_6604,N_6018);
nand U7304 (N_7304,N_6557,N_6169);
nand U7305 (N_7305,N_6929,N_6074);
and U7306 (N_7306,N_6357,N_6584);
and U7307 (N_7307,N_6930,N_6646);
xor U7308 (N_7308,N_6192,N_6887);
or U7309 (N_7309,N_6573,N_6320);
xnor U7310 (N_7310,N_6256,N_6065);
and U7311 (N_7311,N_6663,N_6405);
nor U7312 (N_7312,N_6836,N_6057);
nor U7313 (N_7313,N_6015,N_6148);
or U7314 (N_7314,N_6914,N_6867);
nand U7315 (N_7315,N_6158,N_6273);
and U7316 (N_7316,N_6079,N_6362);
or U7317 (N_7317,N_6832,N_6019);
xor U7318 (N_7318,N_6372,N_6518);
xnor U7319 (N_7319,N_6031,N_6236);
nor U7320 (N_7320,N_6954,N_6486);
nor U7321 (N_7321,N_6589,N_6841);
nand U7322 (N_7322,N_6731,N_6266);
and U7323 (N_7323,N_6123,N_6709);
and U7324 (N_7324,N_6056,N_6784);
xor U7325 (N_7325,N_6134,N_6758);
nor U7326 (N_7326,N_6305,N_6200);
or U7327 (N_7327,N_6906,N_6993);
and U7328 (N_7328,N_6108,N_6064);
nor U7329 (N_7329,N_6540,N_6744);
nand U7330 (N_7330,N_6538,N_6365);
xor U7331 (N_7331,N_6764,N_6982);
xor U7332 (N_7332,N_6210,N_6745);
and U7333 (N_7333,N_6245,N_6947);
nor U7334 (N_7334,N_6893,N_6136);
and U7335 (N_7335,N_6586,N_6653);
nor U7336 (N_7336,N_6833,N_6523);
xnor U7337 (N_7337,N_6325,N_6182);
or U7338 (N_7338,N_6326,N_6174);
or U7339 (N_7339,N_6869,N_6006);
nand U7340 (N_7340,N_6190,N_6683);
and U7341 (N_7341,N_6725,N_6513);
and U7342 (N_7342,N_6416,N_6794);
xor U7343 (N_7343,N_6426,N_6344);
or U7344 (N_7344,N_6815,N_6381);
nand U7345 (N_7345,N_6276,N_6516);
and U7346 (N_7346,N_6863,N_6407);
or U7347 (N_7347,N_6860,N_6298);
or U7348 (N_7348,N_6072,N_6162);
xnor U7349 (N_7349,N_6233,N_6568);
xor U7350 (N_7350,N_6061,N_6145);
xor U7351 (N_7351,N_6375,N_6911);
nor U7352 (N_7352,N_6517,N_6685);
nand U7353 (N_7353,N_6016,N_6680);
nor U7354 (N_7354,N_6401,N_6323);
xnor U7355 (N_7355,N_6558,N_6499);
nor U7356 (N_7356,N_6013,N_6220);
nand U7357 (N_7357,N_6458,N_6413);
nand U7358 (N_7358,N_6959,N_6746);
and U7359 (N_7359,N_6452,N_6141);
xor U7360 (N_7360,N_6364,N_6249);
xnor U7361 (N_7361,N_6779,N_6915);
and U7362 (N_7362,N_6661,N_6593);
or U7363 (N_7363,N_6975,N_6297);
and U7364 (N_7364,N_6248,N_6889);
xnor U7365 (N_7365,N_6219,N_6500);
and U7366 (N_7366,N_6666,N_6193);
nor U7367 (N_7367,N_6386,N_6739);
xor U7368 (N_7368,N_6012,N_6340);
nand U7369 (N_7369,N_6483,N_6293);
xor U7370 (N_7370,N_6619,N_6442);
nor U7371 (N_7371,N_6793,N_6747);
and U7372 (N_7372,N_6831,N_6659);
and U7373 (N_7373,N_6524,N_6734);
nand U7374 (N_7374,N_6207,N_6687);
nor U7375 (N_7375,N_6737,N_6473);
or U7376 (N_7376,N_6958,N_6643);
nand U7377 (N_7377,N_6699,N_6343);
nor U7378 (N_7378,N_6809,N_6131);
or U7379 (N_7379,N_6093,N_6146);
nand U7380 (N_7380,N_6868,N_6968);
or U7381 (N_7381,N_6846,N_6198);
nor U7382 (N_7382,N_6042,N_6098);
nor U7383 (N_7383,N_6988,N_6101);
nand U7384 (N_7384,N_6161,N_6104);
xor U7385 (N_7385,N_6627,N_6296);
and U7386 (N_7386,N_6897,N_6733);
and U7387 (N_7387,N_6157,N_6950);
nor U7388 (N_7388,N_6727,N_6618);
or U7389 (N_7389,N_6406,N_6411);
nand U7390 (N_7390,N_6934,N_6063);
xnor U7391 (N_7391,N_6495,N_6457);
and U7392 (N_7392,N_6171,N_6438);
or U7393 (N_7393,N_6398,N_6251);
and U7394 (N_7394,N_6049,N_6983);
or U7395 (N_7395,N_6980,N_6671);
nand U7396 (N_7396,N_6215,N_6100);
nand U7397 (N_7397,N_6533,N_6423);
xnor U7398 (N_7398,N_6480,N_6845);
xor U7399 (N_7399,N_6814,N_6392);
and U7400 (N_7400,N_6441,N_6113);
nor U7401 (N_7401,N_6351,N_6188);
nor U7402 (N_7402,N_6726,N_6775);
or U7403 (N_7403,N_6319,N_6102);
or U7404 (N_7404,N_6090,N_6504);
and U7405 (N_7405,N_6648,N_6308);
and U7406 (N_7406,N_6195,N_6044);
xor U7407 (N_7407,N_6797,N_6972);
and U7408 (N_7408,N_6052,N_6629);
and U7409 (N_7409,N_6640,N_6468);
and U7410 (N_7410,N_6280,N_6781);
or U7411 (N_7411,N_6327,N_6686);
xor U7412 (N_7412,N_6434,N_6951);
or U7413 (N_7413,N_6609,N_6269);
xor U7414 (N_7414,N_6512,N_6927);
xor U7415 (N_7415,N_6164,N_6111);
and U7416 (N_7416,N_6872,N_6886);
nand U7417 (N_7417,N_6229,N_6454);
or U7418 (N_7418,N_6328,N_6740);
xor U7419 (N_7419,N_6690,N_6786);
and U7420 (N_7420,N_6359,N_6032);
nor U7421 (N_7421,N_6211,N_6582);
nor U7422 (N_7422,N_6840,N_6281);
and U7423 (N_7423,N_6408,N_6541);
or U7424 (N_7424,N_6337,N_6307);
nor U7425 (N_7425,N_6014,N_6553);
or U7426 (N_7426,N_6475,N_6920);
nand U7427 (N_7427,N_6237,N_6352);
and U7428 (N_7428,N_6050,N_6599);
nor U7429 (N_7429,N_6743,N_6770);
nor U7430 (N_7430,N_6132,N_6905);
nor U7431 (N_7431,N_6616,N_6302);
and U7432 (N_7432,N_6776,N_6060);
and U7433 (N_7433,N_6240,N_6569);
or U7434 (N_7434,N_6415,N_6439);
and U7435 (N_7435,N_6544,N_6349);
and U7436 (N_7436,N_6712,N_6697);
nor U7437 (N_7437,N_6763,N_6345);
nor U7438 (N_7438,N_6628,N_6130);
nor U7439 (N_7439,N_6799,N_6839);
xor U7440 (N_7440,N_6633,N_6615);
nand U7441 (N_7441,N_6676,N_6026);
xnor U7442 (N_7442,N_6253,N_6126);
nor U7443 (N_7443,N_6650,N_6271);
nor U7444 (N_7444,N_6189,N_6387);
xnor U7445 (N_7445,N_6494,N_6356);
and U7446 (N_7446,N_6891,N_6772);
xnor U7447 (N_7447,N_6080,N_6857);
nand U7448 (N_7448,N_6651,N_6730);
nor U7449 (N_7449,N_6853,N_6881);
or U7450 (N_7450,N_6180,N_6393);
nor U7451 (N_7451,N_6212,N_6842);
xnor U7452 (N_7452,N_6878,N_6147);
or U7453 (N_7453,N_6963,N_6938);
nand U7454 (N_7454,N_6395,N_6701);
nor U7455 (N_7455,N_6339,N_6239);
and U7456 (N_7456,N_6634,N_6432);
nor U7457 (N_7457,N_6760,N_6370);
xor U7458 (N_7458,N_6769,N_6910);
xnor U7459 (N_7459,N_6801,N_6091);
nand U7460 (N_7460,N_6759,N_6742);
xnor U7461 (N_7461,N_6673,N_6597);
or U7462 (N_7462,N_6656,N_6657);
nand U7463 (N_7463,N_6987,N_6301);
and U7464 (N_7464,N_6371,N_6601);
and U7465 (N_7465,N_6672,N_6870);
xnor U7466 (N_7466,N_6053,N_6828);
and U7467 (N_7467,N_6678,N_6692);
xnor U7468 (N_7468,N_6384,N_6152);
nand U7469 (N_7469,N_6600,N_6888);
and U7470 (N_7470,N_6243,N_6017);
xor U7471 (N_7471,N_6109,N_6492);
or U7472 (N_7472,N_6221,N_6848);
xor U7473 (N_7473,N_6741,N_6037);
or U7474 (N_7474,N_6550,N_6196);
or U7475 (N_7475,N_6974,N_6732);
nor U7476 (N_7476,N_6489,N_6717);
and U7477 (N_7477,N_6960,N_6110);
nand U7478 (N_7478,N_6574,N_6284);
or U7479 (N_7479,N_6637,N_6992);
xor U7480 (N_7480,N_6765,N_6496);
xor U7481 (N_7481,N_6955,N_6802);
or U7482 (N_7482,N_6638,N_6274);
nand U7483 (N_7483,N_6847,N_6120);
and U7484 (N_7484,N_6788,N_6907);
or U7485 (N_7485,N_6160,N_6419);
nor U7486 (N_7486,N_6778,N_6755);
xor U7487 (N_7487,N_6342,N_6428);
nor U7488 (N_7488,N_6736,N_6526);
xnor U7489 (N_7489,N_6894,N_6826);
or U7490 (N_7490,N_6449,N_6397);
xnor U7491 (N_7491,N_6103,N_6122);
xnor U7492 (N_7492,N_6336,N_6854);
nand U7493 (N_7493,N_6985,N_6812);
xor U7494 (N_7494,N_6367,N_6009);
nor U7495 (N_7495,N_6970,N_6805);
or U7496 (N_7496,N_6767,N_6380);
nor U7497 (N_7497,N_6850,N_6172);
nor U7498 (N_7498,N_6264,N_6194);
nor U7499 (N_7499,N_6268,N_6796);
nor U7500 (N_7500,N_6629,N_6203);
and U7501 (N_7501,N_6090,N_6062);
or U7502 (N_7502,N_6272,N_6983);
nand U7503 (N_7503,N_6359,N_6357);
nor U7504 (N_7504,N_6234,N_6889);
xor U7505 (N_7505,N_6501,N_6394);
and U7506 (N_7506,N_6493,N_6637);
or U7507 (N_7507,N_6741,N_6995);
xor U7508 (N_7508,N_6834,N_6683);
xnor U7509 (N_7509,N_6363,N_6025);
nor U7510 (N_7510,N_6441,N_6922);
nand U7511 (N_7511,N_6108,N_6349);
xor U7512 (N_7512,N_6945,N_6814);
and U7513 (N_7513,N_6798,N_6508);
xor U7514 (N_7514,N_6670,N_6473);
xor U7515 (N_7515,N_6166,N_6192);
nor U7516 (N_7516,N_6882,N_6745);
and U7517 (N_7517,N_6619,N_6693);
or U7518 (N_7518,N_6970,N_6527);
or U7519 (N_7519,N_6669,N_6714);
or U7520 (N_7520,N_6290,N_6703);
nand U7521 (N_7521,N_6595,N_6288);
xnor U7522 (N_7522,N_6261,N_6614);
nand U7523 (N_7523,N_6269,N_6920);
and U7524 (N_7524,N_6511,N_6387);
xnor U7525 (N_7525,N_6268,N_6793);
nand U7526 (N_7526,N_6861,N_6655);
or U7527 (N_7527,N_6711,N_6191);
nor U7528 (N_7528,N_6285,N_6833);
xor U7529 (N_7529,N_6806,N_6120);
nand U7530 (N_7530,N_6432,N_6512);
and U7531 (N_7531,N_6341,N_6537);
nand U7532 (N_7532,N_6805,N_6425);
or U7533 (N_7533,N_6077,N_6592);
nand U7534 (N_7534,N_6534,N_6765);
and U7535 (N_7535,N_6281,N_6004);
or U7536 (N_7536,N_6650,N_6029);
xnor U7537 (N_7537,N_6255,N_6526);
nand U7538 (N_7538,N_6771,N_6482);
and U7539 (N_7539,N_6310,N_6859);
or U7540 (N_7540,N_6826,N_6758);
nand U7541 (N_7541,N_6873,N_6840);
nor U7542 (N_7542,N_6433,N_6921);
or U7543 (N_7543,N_6710,N_6571);
and U7544 (N_7544,N_6347,N_6435);
and U7545 (N_7545,N_6963,N_6830);
nor U7546 (N_7546,N_6357,N_6415);
and U7547 (N_7547,N_6110,N_6527);
nor U7548 (N_7548,N_6801,N_6803);
and U7549 (N_7549,N_6540,N_6855);
nand U7550 (N_7550,N_6605,N_6519);
xnor U7551 (N_7551,N_6675,N_6604);
nand U7552 (N_7552,N_6733,N_6006);
nand U7553 (N_7553,N_6886,N_6750);
nand U7554 (N_7554,N_6398,N_6911);
nor U7555 (N_7555,N_6282,N_6946);
nor U7556 (N_7556,N_6461,N_6228);
or U7557 (N_7557,N_6657,N_6081);
and U7558 (N_7558,N_6715,N_6544);
xnor U7559 (N_7559,N_6392,N_6829);
xor U7560 (N_7560,N_6928,N_6735);
nand U7561 (N_7561,N_6129,N_6332);
xor U7562 (N_7562,N_6560,N_6550);
xnor U7563 (N_7563,N_6129,N_6786);
nand U7564 (N_7564,N_6306,N_6045);
and U7565 (N_7565,N_6875,N_6123);
or U7566 (N_7566,N_6961,N_6177);
xnor U7567 (N_7567,N_6631,N_6989);
or U7568 (N_7568,N_6415,N_6404);
xnor U7569 (N_7569,N_6271,N_6321);
nor U7570 (N_7570,N_6166,N_6535);
and U7571 (N_7571,N_6629,N_6375);
nand U7572 (N_7572,N_6871,N_6012);
nand U7573 (N_7573,N_6605,N_6359);
and U7574 (N_7574,N_6819,N_6852);
or U7575 (N_7575,N_6733,N_6544);
nand U7576 (N_7576,N_6404,N_6105);
nor U7577 (N_7577,N_6884,N_6878);
and U7578 (N_7578,N_6006,N_6122);
nand U7579 (N_7579,N_6699,N_6646);
nand U7580 (N_7580,N_6202,N_6510);
and U7581 (N_7581,N_6548,N_6962);
or U7582 (N_7582,N_6084,N_6452);
nand U7583 (N_7583,N_6552,N_6051);
or U7584 (N_7584,N_6533,N_6032);
xor U7585 (N_7585,N_6871,N_6654);
nand U7586 (N_7586,N_6787,N_6509);
nor U7587 (N_7587,N_6047,N_6894);
nand U7588 (N_7588,N_6183,N_6636);
nor U7589 (N_7589,N_6074,N_6451);
and U7590 (N_7590,N_6714,N_6452);
nor U7591 (N_7591,N_6243,N_6413);
xor U7592 (N_7592,N_6818,N_6598);
xor U7593 (N_7593,N_6710,N_6384);
nand U7594 (N_7594,N_6323,N_6387);
nand U7595 (N_7595,N_6877,N_6301);
and U7596 (N_7596,N_6156,N_6518);
nor U7597 (N_7597,N_6033,N_6922);
and U7598 (N_7598,N_6227,N_6828);
and U7599 (N_7599,N_6602,N_6862);
nand U7600 (N_7600,N_6081,N_6297);
or U7601 (N_7601,N_6185,N_6262);
nor U7602 (N_7602,N_6184,N_6644);
nand U7603 (N_7603,N_6069,N_6838);
or U7604 (N_7604,N_6445,N_6148);
nor U7605 (N_7605,N_6747,N_6858);
or U7606 (N_7606,N_6279,N_6071);
or U7607 (N_7607,N_6268,N_6252);
nor U7608 (N_7608,N_6252,N_6102);
xor U7609 (N_7609,N_6270,N_6456);
xnor U7610 (N_7610,N_6663,N_6777);
nor U7611 (N_7611,N_6347,N_6390);
and U7612 (N_7612,N_6349,N_6822);
xor U7613 (N_7613,N_6866,N_6925);
nand U7614 (N_7614,N_6303,N_6716);
and U7615 (N_7615,N_6968,N_6214);
xor U7616 (N_7616,N_6486,N_6284);
or U7617 (N_7617,N_6388,N_6754);
xor U7618 (N_7618,N_6295,N_6642);
nor U7619 (N_7619,N_6083,N_6229);
xor U7620 (N_7620,N_6126,N_6863);
xnor U7621 (N_7621,N_6346,N_6771);
and U7622 (N_7622,N_6321,N_6698);
xor U7623 (N_7623,N_6916,N_6372);
xor U7624 (N_7624,N_6996,N_6963);
nor U7625 (N_7625,N_6763,N_6505);
nor U7626 (N_7626,N_6208,N_6688);
and U7627 (N_7627,N_6065,N_6999);
nor U7628 (N_7628,N_6481,N_6496);
xnor U7629 (N_7629,N_6251,N_6026);
or U7630 (N_7630,N_6941,N_6620);
nand U7631 (N_7631,N_6018,N_6689);
or U7632 (N_7632,N_6761,N_6549);
nand U7633 (N_7633,N_6480,N_6595);
and U7634 (N_7634,N_6358,N_6841);
nand U7635 (N_7635,N_6366,N_6154);
and U7636 (N_7636,N_6937,N_6880);
or U7637 (N_7637,N_6869,N_6043);
and U7638 (N_7638,N_6157,N_6976);
nand U7639 (N_7639,N_6178,N_6454);
nor U7640 (N_7640,N_6881,N_6442);
or U7641 (N_7641,N_6234,N_6680);
nand U7642 (N_7642,N_6253,N_6735);
or U7643 (N_7643,N_6530,N_6072);
and U7644 (N_7644,N_6501,N_6409);
nor U7645 (N_7645,N_6183,N_6233);
or U7646 (N_7646,N_6706,N_6422);
or U7647 (N_7647,N_6608,N_6701);
xor U7648 (N_7648,N_6370,N_6222);
nand U7649 (N_7649,N_6650,N_6571);
and U7650 (N_7650,N_6165,N_6279);
nand U7651 (N_7651,N_6917,N_6245);
xnor U7652 (N_7652,N_6310,N_6779);
xnor U7653 (N_7653,N_6225,N_6689);
nor U7654 (N_7654,N_6327,N_6793);
nand U7655 (N_7655,N_6867,N_6365);
nand U7656 (N_7656,N_6238,N_6771);
nand U7657 (N_7657,N_6931,N_6722);
or U7658 (N_7658,N_6520,N_6447);
xnor U7659 (N_7659,N_6641,N_6618);
xnor U7660 (N_7660,N_6543,N_6480);
nor U7661 (N_7661,N_6882,N_6075);
xor U7662 (N_7662,N_6989,N_6656);
nand U7663 (N_7663,N_6890,N_6524);
nand U7664 (N_7664,N_6490,N_6765);
or U7665 (N_7665,N_6178,N_6044);
nand U7666 (N_7666,N_6126,N_6449);
nand U7667 (N_7667,N_6640,N_6840);
xnor U7668 (N_7668,N_6794,N_6435);
and U7669 (N_7669,N_6923,N_6841);
nand U7670 (N_7670,N_6536,N_6090);
nor U7671 (N_7671,N_6307,N_6338);
or U7672 (N_7672,N_6414,N_6221);
nor U7673 (N_7673,N_6637,N_6870);
xor U7674 (N_7674,N_6439,N_6189);
xnor U7675 (N_7675,N_6901,N_6379);
nor U7676 (N_7676,N_6196,N_6702);
nor U7677 (N_7677,N_6193,N_6562);
nand U7678 (N_7678,N_6163,N_6382);
xnor U7679 (N_7679,N_6054,N_6628);
nand U7680 (N_7680,N_6898,N_6631);
nor U7681 (N_7681,N_6784,N_6529);
or U7682 (N_7682,N_6400,N_6847);
or U7683 (N_7683,N_6646,N_6282);
xor U7684 (N_7684,N_6060,N_6361);
and U7685 (N_7685,N_6752,N_6194);
and U7686 (N_7686,N_6066,N_6378);
or U7687 (N_7687,N_6013,N_6542);
nand U7688 (N_7688,N_6236,N_6761);
nor U7689 (N_7689,N_6061,N_6813);
xor U7690 (N_7690,N_6920,N_6506);
nand U7691 (N_7691,N_6973,N_6902);
or U7692 (N_7692,N_6523,N_6607);
or U7693 (N_7693,N_6047,N_6145);
or U7694 (N_7694,N_6945,N_6115);
nor U7695 (N_7695,N_6455,N_6809);
nor U7696 (N_7696,N_6707,N_6949);
nor U7697 (N_7697,N_6088,N_6308);
or U7698 (N_7698,N_6113,N_6866);
xor U7699 (N_7699,N_6579,N_6164);
and U7700 (N_7700,N_6305,N_6302);
or U7701 (N_7701,N_6733,N_6489);
nand U7702 (N_7702,N_6742,N_6492);
xor U7703 (N_7703,N_6176,N_6880);
xor U7704 (N_7704,N_6413,N_6497);
nand U7705 (N_7705,N_6885,N_6334);
nor U7706 (N_7706,N_6550,N_6055);
and U7707 (N_7707,N_6458,N_6351);
or U7708 (N_7708,N_6326,N_6340);
and U7709 (N_7709,N_6114,N_6269);
nand U7710 (N_7710,N_6923,N_6623);
nand U7711 (N_7711,N_6222,N_6098);
xnor U7712 (N_7712,N_6680,N_6522);
or U7713 (N_7713,N_6107,N_6950);
xor U7714 (N_7714,N_6338,N_6843);
xor U7715 (N_7715,N_6484,N_6788);
and U7716 (N_7716,N_6606,N_6268);
or U7717 (N_7717,N_6530,N_6438);
nand U7718 (N_7718,N_6923,N_6322);
or U7719 (N_7719,N_6625,N_6068);
or U7720 (N_7720,N_6677,N_6040);
xor U7721 (N_7721,N_6788,N_6868);
nor U7722 (N_7722,N_6976,N_6080);
and U7723 (N_7723,N_6988,N_6064);
or U7724 (N_7724,N_6416,N_6284);
xor U7725 (N_7725,N_6662,N_6127);
xnor U7726 (N_7726,N_6700,N_6548);
and U7727 (N_7727,N_6368,N_6044);
nor U7728 (N_7728,N_6105,N_6398);
or U7729 (N_7729,N_6941,N_6524);
xnor U7730 (N_7730,N_6512,N_6804);
or U7731 (N_7731,N_6003,N_6768);
or U7732 (N_7732,N_6895,N_6571);
or U7733 (N_7733,N_6633,N_6089);
nand U7734 (N_7734,N_6865,N_6349);
or U7735 (N_7735,N_6015,N_6282);
xor U7736 (N_7736,N_6456,N_6412);
nand U7737 (N_7737,N_6338,N_6166);
nor U7738 (N_7738,N_6686,N_6482);
and U7739 (N_7739,N_6917,N_6516);
and U7740 (N_7740,N_6416,N_6805);
nor U7741 (N_7741,N_6002,N_6264);
xor U7742 (N_7742,N_6646,N_6805);
nand U7743 (N_7743,N_6171,N_6115);
nor U7744 (N_7744,N_6416,N_6662);
or U7745 (N_7745,N_6937,N_6062);
xnor U7746 (N_7746,N_6653,N_6720);
nor U7747 (N_7747,N_6780,N_6270);
xor U7748 (N_7748,N_6028,N_6879);
or U7749 (N_7749,N_6711,N_6375);
xor U7750 (N_7750,N_6735,N_6966);
and U7751 (N_7751,N_6538,N_6273);
and U7752 (N_7752,N_6582,N_6643);
xnor U7753 (N_7753,N_6752,N_6944);
nand U7754 (N_7754,N_6490,N_6618);
nand U7755 (N_7755,N_6864,N_6219);
nand U7756 (N_7756,N_6172,N_6238);
nor U7757 (N_7757,N_6665,N_6358);
xnor U7758 (N_7758,N_6126,N_6149);
xor U7759 (N_7759,N_6302,N_6374);
or U7760 (N_7760,N_6054,N_6845);
and U7761 (N_7761,N_6900,N_6135);
or U7762 (N_7762,N_6892,N_6399);
nand U7763 (N_7763,N_6001,N_6345);
and U7764 (N_7764,N_6161,N_6011);
and U7765 (N_7765,N_6506,N_6430);
xor U7766 (N_7766,N_6184,N_6079);
nand U7767 (N_7767,N_6233,N_6562);
or U7768 (N_7768,N_6070,N_6630);
and U7769 (N_7769,N_6987,N_6512);
and U7770 (N_7770,N_6354,N_6666);
nand U7771 (N_7771,N_6584,N_6287);
xnor U7772 (N_7772,N_6856,N_6897);
or U7773 (N_7773,N_6001,N_6269);
nor U7774 (N_7774,N_6554,N_6898);
and U7775 (N_7775,N_6352,N_6810);
and U7776 (N_7776,N_6545,N_6309);
nor U7777 (N_7777,N_6805,N_6147);
nor U7778 (N_7778,N_6688,N_6118);
xor U7779 (N_7779,N_6045,N_6948);
nor U7780 (N_7780,N_6380,N_6457);
nand U7781 (N_7781,N_6485,N_6220);
and U7782 (N_7782,N_6963,N_6785);
nand U7783 (N_7783,N_6344,N_6020);
nor U7784 (N_7784,N_6872,N_6520);
and U7785 (N_7785,N_6618,N_6229);
nand U7786 (N_7786,N_6006,N_6448);
or U7787 (N_7787,N_6592,N_6261);
or U7788 (N_7788,N_6427,N_6033);
xnor U7789 (N_7789,N_6037,N_6250);
and U7790 (N_7790,N_6867,N_6595);
nor U7791 (N_7791,N_6174,N_6657);
and U7792 (N_7792,N_6975,N_6889);
and U7793 (N_7793,N_6307,N_6280);
or U7794 (N_7794,N_6202,N_6032);
xnor U7795 (N_7795,N_6387,N_6060);
xnor U7796 (N_7796,N_6349,N_6720);
or U7797 (N_7797,N_6541,N_6440);
and U7798 (N_7798,N_6652,N_6656);
nor U7799 (N_7799,N_6454,N_6222);
nor U7800 (N_7800,N_6263,N_6041);
or U7801 (N_7801,N_6962,N_6792);
nand U7802 (N_7802,N_6964,N_6791);
nor U7803 (N_7803,N_6838,N_6689);
nand U7804 (N_7804,N_6186,N_6147);
xnor U7805 (N_7805,N_6647,N_6814);
nand U7806 (N_7806,N_6721,N_6254);
nor U7807 (N_7807,N_6183,N_6663);
xnor U7808 (N_7808,N_6837,N_6085);
and U7809 (N_7809,N_6643,N_6874);
xor U7810 (N_7810,N_6954,N_6894);
nor U7811 (N_7811,N_6189,N_6348);
and U7812 (N_7812,N_6642,N_6918);
and U7813 (N_7813,N_6681,N_6255);
xnor U7814 (N_7814,N_6965,N_6800);
or U7815 (N_7815,N_6236,N_6149);
xor U7816 (N_7816,N_6741,N_6144);
xnor U7817 (N_7817,N_6881,N_6572);
or U7818 (N_7818,N_6265,N_6318);
nor U7819 (N_7819,N_6236,N_6604);
and U7820 (N_7820,N_6508,N_6447);
nand U7821 (N_7821,N_6509,N_6077);
xnor U7822 (N_7822,N_6849,N_6165);
xor U7823 (N_7823,N_6494,N_6374);
xor U7824 (N_7824,N_6477,N_6542);
xnor U7825 (N_7825,N_6177,N_6268);
nor U7826 (N_7826,N_6651,N_6501);
nand U7827 (N_7827,N_6822,N_6851);
nor U7828 (N_7828,N_6465,N_6182);
nand U7829 (N_7829,N_6691,N_6222);
and U7830 (N_7830,N_6021,N_6352);
nor U7831 (N_7831,N_6440,N_6666);
xor U7832 (N_7832,N_6335,N_6251);
nand U7833 (N_7833,N_6423,N_6525);
nor U7834 (N_7834,N_6787,N_6536);
xnor U7835 (N_7835,N_6609,N_6215);
xor U7836 (N_7836,N_6770,N_6537);
nor U7837 (N_7837,N_6782,N_6439);
and U7838 (N_7838,N_6893,N_6333);
nand U7839 (N_7839,N_6910,N_6959);
nand U7840 (N_7840,N_6563,N_6189);
nor U7841 (N_7841,N_6956,N_6766);
xnor U7842 (N_7842,N_6240,N_6720);
and U7843 (N_7843,N_6164,N_6341);
nor U7844 (N_7844,N_6205,N_6311);
nor U7845 (N_7845,N_6267,N_6232);
or U7846 (N_7846,N_6187,N_6365);
and U7847 (N_7847,N_6348,N_6486);
nor U7848 (N_7848,N_6322,N_6149);
xnor U7849 (N_7849,N_6514,N_6364);
xor U7850 (N_7850,N_6163,N_6936);
xor U7851 (N_7851,N_6946,N_6141);
xnor U7852 (N_7852,N_6603,N_6068);
xnor U7853 (N_7853,N_6284,N_6280);
nor U7854 (N_7854,N_6625,N_6143);
or U7855 (N_7855,N_6683,N_6489);
or U7856 (N_7856,N_6839,N_6289);
nand U7857 (N_7857,N_6628,N_6156);
xnor U7858 (N_7858,N_6163,N_6362);
or U7859 (N_7859,N_6567,N_6060);
and U7860 (N_7860,N_6420,N_6348);
xor U7861 (N_7861,N_6509,N_6686);
nor U7862 (N_7862,N_6255,N_6676);
nand U7863 (N_7863,N_6848,N_6207);
nor U7864 (N_7864,N_6369,N_6255);
xnor U7865 (N_7865,N_6080,N_6151);
or U7866 (N_7866,N_6977,N_6810);
or U7867 (N_7867,N_6427,N_6291);
nor U7868 (N_7868,N_6024,N_6615);
xnor U7869 (N_7869,N_6387,N_6237);
nor U7870 (N_7870,N_6721,N_6549);
or U7871 (N_7871,N_6507,N_6185);
and U7872 (N_7872,N_6905,N_6509);
or U7873 (N_7873,N_6701,N_6744);
xnor U7874 (N_7874,N_6053,N_6370);
nand U7875 (N_7875,N_6901,N_6376);
nor U7876 (N_7876,N_6877,N_6935);
or U7877 (N_7877,N_6146,N_6500);
nor U7878 (N_7878,N_6390,N_6497);
nand U7879 (N_7879,N_6812,N_6080);
and U7880 (N_7880,N_6004,N_6722);
nand U7881 (N_7881,N_6086,N_6498);
and U7882 (N_7882,N_6571,N_6267);
nor U7883 (N_7883,N_6304,N_6044);
and U7884 (N_7884,N_6533,N_6410);
or U7885 (N_7885,N_6923,N_6814);
or U7886 (N_7886,N_6703,N_6566);
and U7887 (N_7887,N_6388,N_6887);
or U7888 (N_7888,N_6294,N_6574);
nor U7889 (N_7889,N_6100,N_6306);
nor U7890 (N_7890,N_6025,N_6223);
nor U7891 (N_7891,N_6608,N_6651);
nor U7892 (N_7892,N_6857,N_6467);
nand U7893 (N_7893,N_6186,N_6822);
and U7894 (N_7894,N_6134,N_6346);
nor U7895 (N_7895,N_6034,N_6802);
xor U7896 (N_7896,N_6821,N_6206);
nor U7897 (N_7897,N_6911,N_6504);
or U7898 (N_7898,N_6503,N_6327);
xor U7899 (N_7899,N_6803,N_6292);
xor U7900 (N_7900,N_6828,N_6835);
xnor U7901 (N_7901,N_6022,N_6592);
or U7902 (N_7902,N_6089,N_6462);
and U7903 (N_7903,N_6240,N_6037);
or U7904 (N_7904,N_6168,N_6724);
xor U7905 (N_7905,N_6696,N_6096);
nor U7906 (N_7906,N_6096,N_6409);
or U7907 (N_7907,N_6683,N_6732);
and U7908 (N_7908,N_6385,N_6926);
nor U7909 (N_7909,N_6919,N_6904);
nand U7910 (N_7910,N_6835,N_6730);
and U7911 (N_7911,N_6289,N_6614);
or U7912 (N_7912,N_6809,N_6658);
xnor U7913 (N_7913,N_6295,N_6800);
xor U7914 (N_7914,N_6850,N_6973);
nor U7915 (N_7915,N_6425,N_6095);
or U7916 (N_7916,N_6513,N_6873);
and U7917 (N_7917,N_6249,N_6862);
and U7918 (N_7918,N_6129,N_6657);
nand U7919 (N_7919,N_6768,N_6582);
nor U7920 (N_7920,N_6063,N_6581);
nand U7921 (N_7921,N_6434,N_6162);
or U7922 (N_7922,N_6861,N_6625);
nand U7923 (N_7923,N_6517,N_6931);
nor U7924 (N_7924,N_6760,N_6851);
nand U7925 (N_7925,N_6157,N_6521);
nand U7926 (N_7926,N_6275,N_6722);
or U7927 (N_7927,N_6044,N_6296);
nand U7928 (N_7928,N_6099,N_6027);
or U7929 (N_7929,N_6152,N_6091);
and U7930 (N_7930,N_6724,N_6114);
or U7931 (N_7931,N_6241,N_6505);
nand U7932 (N_7932,N_6366,N_6978);
xnor U7933 (N_7933,N_6022,N_6609);
nor U7934 (N_7934,N_6396,N_6238);
nor U7935 (N_7935,N_6373,N_6138);
nand U7936 (N_7936,N_6780,N_6842);
nand U7937 (N_7937,N_6965,N_6130);
nor U7938 (N_7938,N_6853,N_6341);
xnor U7939 (N_7939,N_6657,N_6690);
and U7940 (N_7940,N_6162,N_6666);
nor U7941 (N_7941,N_6379,N_6024);
nand U7942 (N_7942,N_6696,N_6709);
nor U7943 (N_7943,N_6036,N_6238);
nand U7944 (N_7944,N_6795,N_6739);
and U7945 (N_7945,N_6593,N_6134);
and U7946 (N_7946,N_6597,N_6267);
nor U7947 (N_7947,N_6400,N_6275);
and U7948 (N_7948,N_6033,N_6843);
xnor U7949 (N_7949,N_6099,N_6539);
xor U7950 (N_7950,N_6801,N_6153);
nor U7951 (N_7951,N_6070,N_6751);
or U7952 (N_7952,N_6546,N_6669);
and U7953 (N_7953,N_6922,N_6192);
nand U7954 (N_7954,N_6536,N_6514);
and U7955 (N_7955,N_6369,N_6473);
xnor U7956 (N_7956,N_6258,N_6719);
or U7957 (N_7957,N_6706,N_6400);
xor U7958 (N_7958,N_6505,N_6322);
xnor U7959 (N_7959,N_6943,N_6129);
nand U7960 (N_7960,N_6147,N_6282);
nor U7961 (N_7961,N_6089,N_6063);
and U7962 (N_7962,N_6747,N_6953);
and U7963 (N_7963,N_6293,N_6129);
nor U7964 (N_7964,N_6993,N_6408);
and U7965 (N_7965,N_6119,N_6574);
xor U7966 (N_7966,N_6971,N_6531);
or U7967 (N_7967,N_6644,N_6450);
and U7968 (N_7968,N_6124,N_6609);
and U7969 (N_7969,N_6188,N_6244);
and U7970 (N_7970,N_6371,N_6741);
nor U7971 (N_7971,N_6237,N_6976);
nand U7972 (N_7972,N_6257,N_6304);
nor U7973 (N_7973,N_6830,N_6954);
or U7974 (N_7974,N_6486,N_6823);
or U7975 (N_7975,N_6368,N_6838);
and U7976 (N_7976,N_6407,N_6488);
nand U7977 (N_7977,N_6730,N_6913);
nand U7978 (N_7978,N_6953,N_6071);
nor U7979 (N_7979,N_6692,N_6388);
nor U7980 (N_7980,N_6168,N_6481);
and U7981 (N_7981,N_6576,N_6514);
nand U7982 (N_7982,N_6319,N_6330);
nor U7983 (N_7983,N_6974,N_6896);
and U7984 (N_7984,N_6904,N_6345);
nand U7985 (N_7985,N_6338,N_6892);
nand U7986 (N_7986,N_6600,N_6990);
nor U7987 (N_7987,N_6437,N_6466);
and U7988 (N_7988,N_6854,N_6566);
xnor U7989 (N_7989,N_6890,N_6793);
or U7990 (N_7990,N_6062,N_6853);
nor U7991 (N_7991,N_6424,N_6134);
and U7992 (N_7992,N_6926,N_6003);
and U7993 (N_7993,N_6940,N_6626);
or U7994 (N_7994,N_6844,N_6583);
nor U7995 (N_7995,N_6713,N_6582);
and U7996 (N_7996,N_6195,N_6183);
nor U7997 (N_7997,N_6722,N_6562);
xor U7998 (N_7998,N_6651,N_6219);
or U7999 (N_7999,N_6137,N_6563);
and U8000 (N_8000,N_7906,N_7136);
nand U8001 (N_8001,N_7152,N_7976);
or U8002 (N_8002,N_7553,N_7446);
nand U8003 (N_8003,N_7192,N_7880);
nand U8004 (N_8004,N_7320,N_7038);
xor U8005 (N_8005,N_7035,N_7308);
and U8006 (N_8006,N_7934,N_7274);
and U8007 (N_8007,N_7220,N_7262);
nor U8008 (N_8008,N_7734,N_7706);
nand U8009 (N_8009,N_7813,N_7070);
nand U8010 (N_8010,N_7882,N_7673);
or U8011 (N_8011,N_7771,N_7477);
or U8012 (N_8012,N_7503,N_7504);
nor U8013 (N_8013,N_7143,N_7228);
nor U8014 (N_8014,N_7573,N_7806);
nand U8015 (N_8015,N_7025,N_7109);
nand U8016 (N_8016,N_7049,N_7453);
or U8017 (N_8017,N_7582,N_7926);
nor U8018 (N_8018,N_7326,N_7467);
nor U8019 (N_8019,N_7655,N_7741);
and U8020 (N_8020,N_7956,N_7726);
nor U8021 (N_8021,N_7384,N_7554);
nor U8022 (N_8022,N_7358,N_7563);
and U8023 (N_8023,N_7762,N_7279);
nor U8024 (N_8024,N_7885,N_7822);
or U8025 (N_8025,N_7509,N_7249);
nor U8026 (N_8026,N_7912,N_7046);
xnor U8027 (N_8027,N_7953,N_7597);
nand U8028 (N_8028,N_7742,N_7286);
xor U8029 (N_8029,N_7469,N_7260);
nor U8030 (N_8030,N_7856,N_7349);
nand U8031 (N_8031,N_7105,N_7300);
or U8032 (N_8032,N_7481,N_7548);
or U8033 (N_8033,N_7555,N_7993);
xor U8034 (N_8034,N_7017,N_7492);
and U8035 (N_8035,N_7275,N_7016);
or U8036 (N_8036,N_7996,N_7617);
nor U8037 (N_8037,N_7518,N_7858);
or U8038 (N_8038,N_7306,N_7499);
or U8039 (N_8039,N_7416,N_7658);
xor U8040 (N_8040,N_7718,N_7204);
or U8041 (N_8041,N_7559,N_7955);
nand U8042 (N_8042,N_7997,N_7857);
or U8043 (N_8043,N_7244,N_7276);
nand U8044 (N_8044,N_7412,N_7685);
nand U8045 (N_8045,N_7310,N_7799);
nor U8046 (N_8046,N_7913,N_7432);
nand U8047 (N_8047,N_7950,N_7414);
xnor U8048 (N_8048,N_7805,N_7480);
or U8049 (N_8049,N_7929,N_7606);
xnor U8050 (N_8050,N_7870,N_7705);
or U8051 (N_8051,N_7425,N_7285);
nor U8052 (N_8052,N_7680,N_7634);
or U8053 (N_8053,N_7712,N_7397);
xnor U8054 (N_8054,N_7466,N_7268);
and U8055 (N_8055,N_7500,N_7359);
or U8056 (N_8056,N_7866,N_7602);
nand U8057 (N_8057,N_7002,N_7339);
nor U8058 (N_8058,N_7508,N_7398);
nand U8059 (N_8059,N_7487,N_7059);
nor U8060 (N_8060,N_7238,N_7878);
and U8061 (N_8061,N_7795,N_7200);
xnor U8062 (N_8062,N_7945,N_7507);
xnor U8063 (N_8063,N_7153,N_7482);
or U8064 (N_8064,N_7264,N_7635);
or U8065 (N_8065,N_7571,N_7701);
nor U8066 (N_8066,N_7526,N_7015);
or U8067 (N_8067,N_7226,N_7041);
and U8068 (N_8068,N_7545,N_7170);
and U8069 (N_8069,N_7447,N_7373);
xor U8070 (N_8070,N_7861,N_7883);
xor U8071 (N_8071,N_7061,N_7445);
and U8072 (N_8072,N_7840,N_7340);
nand U8073 (N_8073,N_7135,N_7291);
and U8074 (N_8074,N_7263,N_7158);
or U8075 (N_8075,N_7045,N_7778);
or U8076 (N_8076,N_7328,N_7325);
nor U8077 (N_8077,N_7909,N_7527);
and U8078 (N_8078,N_7704,N_7368);
or U8079 (N_8079,N_7639,N_7483);
xor U8080 (N_8080,N_7042,N_7405);
or U8081 (N_8081,N_7937,N_7128);
nor U8082 (N_8082,N_7221,N_7892);
xor U8083 (N_8083,N_7255,N_7441);
nor U8084 (N_8084,N_7583,N_7399);
nor U8085 (N_8085,N_7756,N_7242);
and U8086 (N_8086,N_7970,N_7120);
nand U8087 (N_8087,N_7863,N_7572);
and U8088 (N_8088,N_7738,N_7211);
xor U8089 (N_8089,N_7438,N_7356);
xor U8090 (N_8090,N_7694,N_7000);
nor U8091 (N_8091,N_7295,N_7853);
or U8092 (N_8092,N_7251,N_7519);
nand U8093 (N_8093,N_7486,N_7385);
xor U8094 (N_8094,N_7184,N_7951);
or U8095 (N_8095,N_7243,N_7345);
nand U8096 (N_8096,N_7029,N_7598);
and U8097 (N_8097,N_7093,N_7779);
or U8098 (N_8098,N_7832,N_7815);
nand U8099 (N_8099,N_7921,N_7064);
nand U8100 (N_8100,N_7936,N_7944);
or U8101 (N_8101,N_7139,N_7828);
and U8102 (N_8102,N_7485,N_7194);
nand U8103 (N_8103,N_7952,N_7835);
xnor U8104 (N_8104,N_7969,N_7644);
nor U8105 (N_8105,N_7550,N_7721);
nor U8106 (N_8106,N_7925,N_7475);
or U8107 (N_8107,N_7430,N_7390);
nor U8108 (N_8108,N_7411,N_7068);
nand U8109 (N_8109,N_7071,N_7013);
nand U8110 (N_8110,N_7730,N_7422);
xor U8111 (N_8111,N_7531,N_7148);
or U8112 (N_8112,N_7773,N_7253);
nor U8113 (N_8113,N_7871,N_7100);
xor U8114 (N_8114,N_7556,N_7116);
nand U8115 (N_8115,N_7651,N_7740);
nor U8116 (N_8116,N_7981,N_7624);
or U8117 (N_8117,N_7387,N_7661);
or U8118 (N_8118,N_7175,N_7660);
nand U8119 (N_8119,N_7776,N_7298);
and U8120 (N_8120,N_7337,N_7169);
xnor U8121 (N_8121,N_7722,N_7056);
xor U8122 (N_8122,N_7393,N_7094);
or U8123 (N_8123,N_7267,N_7625);
nand U8124 (N_8124,N_7178,N_7428);
nand U8125 (N_8125,N_7665,N_7501);
nand U8126 (N_8126,N_7307,N_7725);
or U8127 (N_8127,N_7463,N_7332);
or U8128 (N_8128,N_7719,N_7363);
nand U8129 (N_8129,N_7887,N_7587);
nor U8130 (N_8130,N_7766,N_7731);
and U8131 (N_8131,N_7163,N_7055);
nand U8132 (N_8132,N_7090,N_7096);
nand U8133 (N_8133,N_7561,N_7189);
nor U8134 (N_8134,N_7562,N_7331);
xor U8135 (N_8135,N_7099,N_7551);
and U8136 (N_8136,N_7123,N_7218);
or U8137 (N_8137,N_7581,N_7686);
nand U8138 (N_8138,N_7942,N_7511);
and U8139 (N_8139,N_7232,N_7736);
nand U8140 (N_8140,N_7770,N_7727);
xor U8141 (N_8141,N_7588,N_7374);
and U8142 (N_8142,N_7205,N_7697);
xnor U8143 (N_8143,N_7314,N_7614);
and U8144 (N_8144,N_7065,N_7372);
or U8145 (N_8145,N_7724,N_7304);
or U8146 (N_8146,N_7278,N_7860);
nor U8147 (N_8147,N_7353,N_7058);
nor U8148 (N_8148,N_7210,N_7968);
and U8149 (N_8149,N_7842,N_7137);
nor U8150 (N_8150,N_7224,N_7073);
nor U8151 (N_8151,N_7437,N_7034);
or U8152 (N_8152,N_7987,N_7979);
and U8153 (N_8153,N_7810,N_7132);
xnor U8154 (N_8154,N_7846,N_7348);
and U8155 (N_8155,N_7746,N_7973);
and U8156 (N_8156,N_7418,N_7819);
and U8157 (N_8157,N_7580,N_7708);
xor U8158 (N_8158,N_7149,N_7789);
xnor U8159 (N_8159,N_7185,N_7141);
and U8160 (N_8160,N_7535,N_7663);
and U8161 (N_8161,N_7947,N_7765);
nor U8162 (N_8162,N_7855,N_7943);
and U8163 (N_8163,N_7388,N_7395);
and U8164 (N_8164,N_7008,N_7893);
xor U8165 (N_8165,N_7958,N_7851);
or U8166 (N_8166,N_7547,N_7436);
nand U8167 (N_8167,N_7330,N_7591);
nor U8168 (N_8168,N_7316,N_7329);
or U8169 (N_8169,N_7579,N_7922);
nand U8170 (N_8170,N_7821,N_7191);
and U8171 (N_8171,N_7261,N_7400);
or U8172 (N_8172,N_7837,N_7693);
nand U8173 (N_8173,N_7811,N_7684);
and U8174 (N_8174,N_7462,N_7653);
nor U8175 (N_8175,N_7824,N_7723);
xnor U8176 (N_8176,N_7424,N_7360);
and U8177 (N_8177,N_7596,N_7364);
nor U8178 (N_8178,N_7510,N_7747);
and U8179 (N_8179,N_7010,N_7516);
nand U8180 (N_8180,N_7523,N_7054);
or U8181 (N_8181,N_7812,N_7172);
or U8182 (N_8182,N_7303,N_7146);
and U8183 (N_8183,N_7538,N_7769);
xnor U8184 (N_8184,N_7933,N_7830);
nor U8185 (N_8185,N_7084,N_7471);
and U8186 (N_8186,N_7378,N_7402);
and U8187 (N_8187,N_7122,N_7618);
nor U8188 (N_8188,N_7103,N_7833);
or U8189 (N_8189,N_7592,N_7667);
and U8190 (N_8190,N_7566,N_7609);
or U8191 (N_8191,N_7020,N_7062);
or U8192 (N_8192,N_7688,N_7108);
nor U8193 (N_8193,N_7315,N_7560);
and U8194 (N_8194,N_7003,N_7959);
nand U8195 (N_8195,N_7623,N_7273);
or U8196 (N_8196,N_7282,N_7759);
or U8197 (N_8197,N_7850,N_7567);
and U8198 (N_8198,N_7362,N_7377);
nor U8199 (N_8199,N_7604,N_7423);
nor U8200 (N_8200,N_7967,N_7739);
nand U8201 (N_8201,N_7230,N_7793);
or U8202 (N_8202,N_7459,N_7394);
xor U8203 (N_8203,N_7001,N_7656);
and U8204 (N_8204,N_7903,N_7245);
nand U8205 (N_8205,N_7338,N_7490);
nand U8206 (N_8206,N_7197,N_7751);
nand U8207 (N_8207,N_7048,N_7069);
and U8208 (N_8208,N_7534,N_7294);
and U8209 (N_8209,N_7415,N_7729);
nand U8210 (N_8210,N_7111,N_7130);
nor U8211 (N_8211,N_7841,N_7608);
nand U8212 (N_8212,N_7112,N_7803);
nor U8213 (N_8213,N_7974,N_7764);
nand U8214 (N_8214,N_7156,N_7030);
xnor U8215 (N_8215,N_7343,N_7067);
xor U8216 (N_8216,N_7344,N_7124);
or U8217 (N_8217,N_7995,N_7027);
and U8218 (N_8218,N_7570,N_7082);
nor U8219 (N_8219,N_7804,N_7732);
or U8220 (N_8220,N_7413,N_7834);
nor U8221 (N_8221,N_7376,N_7992);
nand U8222 (N_8222,N_7988,N_7578);
and U8223 (N_8223,N_7964,N_7826);
xnor U8224 (N_8224,N_7365,N_7820);
nor U8225 (N_8225,N_7502,N_7528);
xor U8226 (N_8226,N_7616,N_7297);
xor U8227 (N_8227,N_7788,N_7775);
nand U8228 (N_8228,N_7790,N_7539);
nand U8229 (N_8229,N_7986,N_7451);
xnor U8230 (N_8230,N_7134,N_7886);
and U8231 (N_8231,N_7900,N_7650);
and U8232 (N_8232,N_7464,N_7050);
xor U8233 (N_8233,N_7435,N_7918);
and U8234 (N_8234,N_7391,N_7076);
or U8235 (N_8235,N_7816,N_7575);
or U8236 (N_8236,N_7229,N_7406);
nor U8237 (N_8237,N_7468,N_7470);
nand U8238 (N_8238,N_7537,N_7881);
nand U8239 (N_8239,N_7915,N_7089);
nand U8240 (N_8240,N_7195,N_7293);
nand U8241 (N_8241,N_7875,N_7493);
or U8242 (N_8242,N_7317,N_7101);
xor U8243 (N_8243,N_7755,N_7199);
nor U8244 (N_8244,N_7808,N_7642);
or U8245 (N_8245,N_7410,N_7777);
or U8246 (N_8246,N_7198,N_7075);
xor U8247 (N_8247,N_7088,N_7202);
nor U8248 (N_8248,N_7322,N_7506);
nand U8249 (N_8249,N_7182,N_7434);
nor U8250 (N_8250,N_7823,N_7495);
xnor U8251 (N_8251,N_7289,N_7839);
xor U8252 (N_8252,N_7234,N_7845);
and U8253 (N_8253,N_7714,N_7515);
nand U8254 (N_8254,N_7744,N_7443);
or U8255 (N_8255,N_7864,N_7085);
nand U8256 (N_8256,N_7737,N_7774);
xnor U8257 (N_8257,N_7521,N_7709);
and U8258 (N_8258,N_7350,N_7215);
nand U8259 (N_8259,N_7159,N_7664);
nor U8260 (N_8260,N_7862,N_7381);
and U8261 (N_8261,N_7342,N_7346);
nand U8262 (N_8262,N_7525,N_7250);
nand U8263 (N_8263,N_7066,N_7629);
nor U8264 (N_8264,N_7142,N_7319);
nand U8265 (N_8265,N_7847,N_7902);
or U8266 (N_8266,N_7849,N_7817);
xor U8267 (N_8267,N_7290,N_7626);
xnor U8268 (N_8268,N_7802,N_7520);
nand U8269 (N_8269,N_7392,N_7540);
xnor U8270 (N_8270,N_7814,N_7077);
nor U8271 (N_8271,N_7999,N_7352);
nand U8272 (N_8272,N_7031,N_7183);
or U8273 (N_8273,N_7208,N_7807);
and U8274 (N_8274,N_7375,N_7831);
or U8275 (N_8275,N_7961,N_7455);
or U8276 (N_8276,N_7063,N_7948);
and U8277 (N_8277,N_7404,N_7167);
xor U8278 (N_8278,N_7081,N_7074);
nor U8279 (N_8279,N_7783,N_7569);
and U8280 (N_8280,N_7825,N_7233);
nor U8281 (N_8281,N_7876,N_7043);
nor U8282 (N_8282,N_7772,N_7098);
xor U8283 (N_8283,N_7919,N_7780);
nor U8284 (N_8284,N_7179,N_7636);
nor U8285 (N_8285,N_7690,N_7897);
xor U8286 (N_8286,N_7785,N_7894);
or U8287 (N_8287,N_7333,N_7036);
nor U8288 (N_8288,N_7728,N_7219);
or U8289 (N_8289,N_7440,N_7594);
nand U8290 (N_8290,N_7461,N_7646);
nor U8291 (N_8291,N_7786,N_7473);
xnor U8292 (N_8292,N_7087,N_7652);
or U8293 (N_8293,N_7239,N_7032);
nor U8294 (N_8294,N_7630,N_7932);
or U8295 (N_8295,N_7852,N_7254);
nor U8296 (N_8296,N_7843,N_7186);
nand U8297 (N_8297,N_7427,N_7888);
nand U8298 (N_8298,N_7641,N_7014);
or U8299 (N_8299,N_7662,N_7484);
or U8300 (N_8300,N_7657,N_7749);
nor U8301 (N_8301,N_7798,N_7426);
nor U8302 (N_8302,N_7072,N_7246);
and U8303 (N_8303,N_7299,N_7166);
or U8304 (N_8304,N_7750,N_7674);
and U8305 (N_8305,N_7227,N_7313);
or U8306 (N_8306,N_7905,N_7079);
nand U8307 (N_8307,N_7542,N_7867);
nor U8308 (N_8308,N_7683,N_7160);
or U8309 (N_8309,N_7498,N_7884);
and U8310 (N_8310,N_7287,N_7341);
and U8311 (N_8311,N_7458,N_7106);
nand U8312 (N_8312,N_7713,N_7114);
nor U8313 (N_8313,N_7396,N_7118);
xnor U8314 (N_8314,N_7336,N_7335);
xnor U8315 (N_8315,N_7627,N_7433);
or U8316 (N_8316,N_7465,N_7366);
xnor U8317 (N_8317,N_7006,N_7666);
xor U8318 (N_8318,N_7868,N_7162);
or U8319 (N_8319,N_7154,N_7370);
or U8320 (N_8320,N_7557,N_7612);
nand U8321 (N_8321,N_7615,N_7083);
and U8322 (N_8322,N_7647,N_7829);
xor U8323 (N_8323,N_7910,N_7768);
or U8324 (N_8324,N_7188,N_7354);
xor U8325 (N_8325,N_7407,N_7181);
xnor U8326 (N_8326,N_7421,N_7827);
or U8327 (N_8327,N_7599,N_7442);
xor U8328 (N_8328,N_7060,N_7125);
nor U8329 (N_8329,N_7691,N_7164);
xnor U8330 (N_8330,N_7367,N_7576);
xor U8331 (N_8331,N_7018,N_7379);
nand U8332 (N_8332,N_7628,N_7654);
nand U8333 (N_8333,N_7758,N_7984);
nand U8334 (N_8334,N_7613,N_7859);
xnor U8335 (N_8335,N_7532,N_7873);
xor U8336 (N_8336,N_7659,N_7311);
nor U8337 (N_8337,N_7488,N_7126);
xor U8338 (N_8338,N_7865,N_7552);
and U8339 (N_8339,N_7217,N_7632);
nand U8340 (N_8340,N_7110,N_7678);
or U8341 (N_8341,N_7403,N_7257);
nor U8342 (N_8342,N_7140,N_7874);
and U8343 (N_8343,N_7895,N_7104);
xor U8344 (N_8344,N_7223,N_7983);
or U8345 (N_8345,N_7904,N_7095);
and U8346 (N_8346,N_7190,N_7097);
and U8347 (N_8347,N_7675,N_7703);
nand U8348 (N_8348,N_7165,N_7147);
or U8349 (N_8349,N_7935,N_7752);
and U8350 (N_8350,N_7222,N_7931);
xnor U8351 (N_8351,N_7022,N_7707);
xor U8352 (N_8352,N_7240,N_7640);
nor U8353 (N_8353,N_7252,N_7280);
xnor U8354 (N_8354,N_7033,N_7457);
nand U8355 (N_8355,N_7574,N_7809);
nor U8356 (N_8356,N_7318,N_7193);
xor U8357 (N_8357,N_7643,N_7600);
or U8358 (N_8358,N_7716,N_7844);
nand U8359 (N_8359,N_7681,N_7975);
and U8360 (N_8360,N_7524,N_7419);
nand U8361 (N_8361,N_7622,N_7593);
xnor U8362 (N_8362,N_7177,N_7444);
xnor U8363 (N_8363,N_7513,N_7129);
or U8364 (N_8364,N_7272,N_7529);
nand U8365 (N_8365,N_7248,N_7127);
and U8366 (N_8366,N_7161,N_7939);
nand U8367 (N_8367,N_7305,N_7610);
nor U8368 (N_8368,N_7800,N_7914);
and U8369 (N_8369,N_7702,N_7687);
xnor U8370 (N_8370,N_7121,N_7568);
nor U8371 (N_8371,N_7896,N_7648);
or U8372 (N_8372,N_7296,N_7005);
nor U8373 (N_8373,N_7607,N_7797);
nand U8374 (N_8374,N_7595,N_7021);
xnor U8375 (N_8375,N_7494,N_7620);
or U8376 (N_8376,N_7818,N_7514);
and U8377 (N_8377,N_7763,N_7638);
xnor U8378 (N_8378,N_7113,N_7505);
nand U8379 (N_8379,N_7603,N_7584);
nand U8380 (N_8380,N_7207,N_7761);
xnor U8381 (N_8381,N_7923,N_7323);
nor U8382 (N_8382,N_7645,N_7266);
nand U8383 (N_8383,N_7460,N_7214);
or U8384 (N_8384,N_7429,N_7115);
xor U8385 (N_8385,N_7138,N_7908);
or U8386 (N_8386,N_7848,N_7277);
and U8387 (N_8387,N_7269,N_7288);
nor U8388 (N_8388,N_7408,N_7891);
and U8389 (N_8389,N_7491,N_7907);
or U8390 (N_8390,N_7157,N_7151);
nand U8391 (N_8391,N_7753,N_7091);
and U8392 (N_8392,N_7474,N_7546);
nand U8393 (N_8393,N_7698,N_7324);
or U8394 (N_8394,N_7450,N_7985);
nor U8395 (N_8395,N_7715,N_7589);
nand U8396 (N_8396,N_7213,N_7028);
xnor U8397 (N_8397,N_7711,N_7092);
xnor U8398 (N_8398,N_7672,N_7512);
nor U8399 (N_8399,N_7700,N_7743);
nor U8400 (N_8400,N_7720,N_7541);
nand U8401 (N_8401,N_7496,N_7930);
xor U8402 (N_8402,N_7619,N_7168);
or U8403 (N_8403,N_7449,N_7924);
nor U8404 (N_8404,N_7355,N_7605);
and U8405 (N_8405,N_7879,N_7899);
nand U8406 (N_8406,N_7794,N_7150);
nor U8407 (N_8407,N_7216,N_7977);
or U8408 (N_8408,N_7321,N_7676);
nand U8409 (N_8409,N_7133,N_7611);
or U8410 (N_8410,N_7649,N_7196);
nand U8411 (N_8411,N_7782,N_7180);
xnor U8412 (N_8412,N_7577,N_7717);
and U8413 (N_8413,N_7302,N_7787);
nand U8414 (N_8414,N_7558,N_7284);
nor U8415 (N_8415,N_7898,N_7386);
and U8416 (N_8416,N_7689,N_7544);
nor U8417 (N_8417,N_7927,N_7247);
or U8418 (N_8418,N_7420,N_7176);
nand U8419 (N_8419,N_7890,N_7361);
and U8420 (N_8420,N_7011,N_7699);
or U8421 (N_8421,N_7009,N_7963);
nand U8422 (N_8422,N_7745,N_7901);
and U8423 (N_8423,N_7949,N_7044);
nand U8424 (N_8424,N_7144,N_7478);
xnor U8425 (N_8425,N_7203,N_7928);
nor U8426 (N_8426,N_7131,N_7051);
nor U8427 (N_8427,N_7053,N_7187);
or U8428 (N_8428,N_7517,N_7889);
nor U8429 (N_8429,N_7004,N_7119);
nand U8430 (N_8430,N_7389,N_7796);
or U8431 (N_8431,N_7448,N_7052);
or U8432 (N_8432,N_7489,N_7533);
or U8433 (N_8433,N_7872,N_7601);
nor U8434 (N_8434,N_7960,N_7236);
nand U8435 (N_8435,N_7401,N_7271);
nand U8436 (N_8436,N_7791,N_7241);
and U8437 (N_8437,N_7760,N_7456);
xnor U8438 (N_8438,N_7235,N_7371);
xor U8439 (N_8439,N_7940,N_7259);
nor U8440 (N_8440,N_7679,N_7966);
nand U8441 (N_8441,N_7978,N_7836);
or U8442 (N_8442,N_7637,N_7991);
nand U8443 (N_8443,N_7023,N_7677);
xor U8444 (N_8444,N_7586,N_7497);
xor U8445 (N_8445,N_7057,N_7171);
or U8446 (N_8446,N_7669,N_7351);
xnor U8447 (N_8447,N_7265,N_7957);
nor U8448 (N_8448,N_7877,N_7767);
and U8449 (N_8449,N_7270,N_7258);
and U8450 (N_8450,N_7312,N_7309);
nand U8451 (N_8451,N_7439,N_7917);
and U8452 (N_8452,N_7522,N_7754);
nor U8453 (N_8453,N_7454,N_7920);
nor U8454 (N_8454,N_7565,N_7431);
or U8455 (N_8455,N_7965,N_7994);
xnor U8456 (N_8456,N_7417,N_7633);
nand U8457 (N_8457,N_7998,N_7383);
nor U8458 (N_8458,N_7938,N_7911);
nand U8459 (N_8459,N_7102,N_7107);
or U8460 (N_8460,N_7212,N_7040);
and U8461 (N_8461,N_7671,N_7047);
or U8462 (N_8462,N_7916,N_7668);
xor U8463 (N_8463,N_7733,N_7472);
or U8464 (N_8464,N_7173,N_7695);
and U8465 (N_8465,N_7281,N_7543);
and U8466 (N_8466,N_7972,N_7530);
nand U8467 (N_8467,N_7971,N_7784);
or U8468 (N_8468,N_7982,N_7231);
nor U8469 (N_8469,N_7283,N_7781);
and U8470 (N_8470,N_7357,N_7735);
and U8471 (N_8471,N_7941,N_7536);
xnor U8472 (N_8472,N_7409,N_7792);
or U8473 (N_8473,N_7748,N_7078);
and U8474 (N_8474,N_7564,N_7334);
nor U8475 (N_8475,N_7117,N_7301);
nand U8476 (N_8476,N_7369,N_7206);
or U8477 (N_8477,N_7631,N_7710);
nand U8478 (N_8478,N_7086,N_7174);
nor U8479 (N_8479,N_7237,N_7292);
nor U8480 (N_8480,N_7980,N_7327);
nand U8481 (N_8481,N_7954,N_7585);
and U8482 (N_8482,N_7256,N_7854);
xor U8483 (N_8483,N_7838,N_7692);
nand U8484 (N_8484,N_7225,N_7590);
nand U8485 (N_8485,N_7201,N_7012);
and U8486 (N_8486,N_7989,N_7080);
xor U8487 (N_8487,N_7549,N_7696);
nor U8488 (N_8488,N_7757,N_7380);
xnor U8489 (N_8489,N_7026,N_7209);
xor U8490 (N_8490,N_7682,N_7476);
nor U8491 (N_8491,N_7039,N_7946);
and U8492 (N_8492,N_7621,N_7024);
nor U8493 (N_8493,N_7347,N_7155);
nor U8494 (N_8494,N_7869,N_7037);
xor U8495 (N_8495,N_7382,N_7007);
nand U8496 (N_8496,N_7801,N_7670);
or U8497 (N_8497,N_7019,N_7990);
nor U8498 (N_8498,N_7962,N_7479);
nor U8499 (N_8499,N_7452,N_7145);
and U8500 (N_8500,N_7168,N_7181);
xnor U8501 (N_8501,N_7821,N_7116);
and U8502 (N_8502,N_7359,N_7370);
or U8503 (N_8503,N_7513,N_7241);
or U8504 (N_8504,N_7945,N_7717);
and U8505 (N_8505,N_7450,N_7730);
nor U8506 (N_8506,N_7353,N_7991);
and U8507 (N_8507,N_7870,N_7311);
xor U8508 (N_8508,N_7071,N_7204);
nor U8509 (N_8509,N_7924,N_7831);
and U8510 (N_8510,N_7944,N_7927);
or U8511 (N_8511,N_7818,N_7785);
or U8512 (N_8512,N_7510,N_7688);
xnor U8513 (N_8513,N_7342,N_7910);
xnor U8514 (N_8514,N_7494,N_7898);
and U8515 (N_8515,N_7472,N_7321);
or U8516 (N_8516,N_7434,N_7064);
nor U8517 (N_8517,N_7306,N_7577);
xnor U8518 (N_8518,N_7774,N_7609);
nand U8519 (N_8519,N_7859,N_7193);
xor U8520 (N_8520,N_7669,N_7504);
and U8521 (N_8521,N_7087,N_7327);
nor U8522 (N_8522,N_7385,N_7030);
or U8523 (N_8523,N_7840,N_7030);
nor U8524 (N_8524,N_7825,N_7405);
or U8525 (N_8525,N_7403,N_7330);
xnor U8526 (N_8526,N_7591,N_7809);
and U8527 (N_8527,N_7434,N_7875);
nand U8528 (N_8528,N_7060,N_7352);
or U8529 (N_8529,N_7321,N_7278);
nand U8530 (N_8530,N_7547,N_7647);
and U8531 (N_8531,N_7024,N_7925);
and U8532 (N_8532,N_7855,N_7559);
xnor U8533 (N_8533,N_7902,N_7866);
xor U8534 (N_8534,N_7300,N_7549);
xor U8535 (N_8535,N_7305,N_7431);
xnor U8536 (N_8536,N_7137,N_7286);
and U8537 (N_8537,N_7538,N_7379);
xnor U8538 (N_8538,N_7147,N_7678);
nand U8539 (N_8539,N_7698,N_7279);
nor U8540 (N_8540,N_7906,N_7898);
or U8541 (N_8541,N_7115,N_7410);
nand U8542 (N_8542,N_7518,N_7136);
nand U8543 (N_8543,N_7533,N_7990);
nand U8544 (N_8544,N_7455,N_7238);
or U8545 (N_8545,N_7795,N_7870);
or U8546 (N_8546,N_7136,N_7719);
nand U8547 (N_8547,N_7075,N_7117);
or U8548 (N_8548,N_7635,N_7283);
or U8549 (N_8549,N_7614,N_7456);
and U8550 (N_8550,N_7897,N_7609);
and U8551 (N_8551,N_7981,N_7470);
xnor U8552 (N_8552,N_7948,N_7923);
xor U8553 (N_8553,N_7316,N_7772);
nor U8554 (N_8554,N_7072,N_7356);
nor U8555 (N_8555,N_7944,N_7369);
nand U8556 (N_8556,N_7437,N_7541);
xor U8557 (N_8557,N_7662,N_7090);
nand U8558 (N_8558,N_7554,N_7743);
nor U8559 (N_8559,N_7353,N_7091);
nand U8560 (N_8560,N_7546,N_7754);
or U8561 (N_8561,N_7759,N_7811);
and U8562 (N_8562,N_7186,N_7517);
and U8563 (N_8563,N_7414,N_7558);
nor U8564 (N_8564,N_7385,N_7084);
and U8565 (N_8565,N_7074,N_7787);
xor U8566 (N_8566,N_7349,N_7552);
nand U8567 (N_8567,N_7856,N_7734);
nand U8568 (N_8568,N_7117,N_7153);
xnor U8569 (N_8569,N_7998,N_7958);
xnor U8570 (N_8570,N_7133,N_7447);
nor U8571 (N_8571,N_7405,N_7266);
nand U8572 (N_8572,N_7867,N_7786);
xor U8573 (N_8573,N_7405,N_7605);
xor U8574 (N_8574,N_7019,N_7342);
and U8575 (N_8575,N_7787,N_7305);
or U8576 (N_8576,N_7211,N_7603);
or U8577 (N_8577,N_7654,N_7022);
xnor U8578 (N_8578,N_7378,N_7807);
xnor U8579 (N_8579,N_7822,N_7173);
xnor U8580 (N_8580,N_7719,N_7231);
xnor U8581 (N_8581,N_7778,N_7346);
xnor U8582 (N_8582,N_7337,N_7857);
and U8583 (N_8583,N_7329,N_7521);
nor U8584 (N_8584,N_7602,N_7975);
or U8585 (N_8585,N_7865,N_7471);
xnor U8586 (N_8586,N_7872,N_7698);
and U8587 (N_8587,N_7726,N_7284);
and U8588 (N_8588,N_7736,N_7846);
nand U8589 (N_8589,N_7612,N_7172);
nor U8590 (N_8590,N_7754,N_7185);
nor U8591 (N_8591,N_7415,N_7738);
and U8592 (N_8592,N_7942,N_7322);
nor U8593 (N_8593,N_7067,N_7664);
xnor U8594 (N_8594,N_7990,N_7607);
nand U8595 (N_8595,N_7131,N_7341);
or U8596 (N_8596,N_7664,N_7060);
nor U8597 (N_8597,N_7813,N_7804);
and U8598 (N_8598,N_7471,N_7872);
or U8599 (N_8599,N_7759,N_7443);
and U8600 (N_8600,N_7140,N_7111);
and U8601 (N_8601,N_7913,N_7562);
nor U8602 (N_8602,N_7818,N_7902);
nand U8603 (N_8603,N_7253,N_7777);
nand U8604 (N_8604,N_7345,N_7799);
nand U8605 (N_8605,N_7586,N_7940);
nor U8606 (N_8606,N_7266,N_7544);
and U8607 (N_8607,N_7717,N_7169);
xnor U8608 (N_8608,N_7450,N_7693);
nand U8609 (N_8609,N_7753,N_7192);
nand U8610 (N_8610,N_7051,N_7940);
xnor U8611 (N_8611,N_7901,N_7104);
and U8612 (N_8612,N_7940,N_7892);
xor U8613 (N_8613,N_7097,N_7433);
nor U8614 (N_8614,N_7151,N_7234);
or U8615 (N_8615,N_7264,N_7772);
xor U8616 (N_8616,N_7546,N_7467);
nand U8617 (N_8617,N_7932,N_7770);
nor U8618 (N_8618,N_7773,N_7967);
or U8619 (N_8619,N_7988,N_7736);
xnor U8620 (N_8620,N_7579,N_7892);
nor U8621 (N_8621,N_7671,N_7408);
nor U8622 (N_8622,N_7366,N_7610);
or U8623 (N_8623,N_7415,N_7140);
nand U8624 (N_8624,N_7014,N_7303);
nand U8625 (N_8625,N_7933,N_7185);
or U8626 (N_8626,N_7244,N_7302);
or U8627 (N_8627,N_7281,N_7267);
and U8628 (N_8628,N_7045,N_7995);
xor U8629 (N_8629,N_7237,N_7268);
or U8630 (N_8630,N_7001,N_7323);
nor U8631 (N_8631,N_7445,N_7688);
nand U8632 (N_8632,N_7776,N_7633);
nand U8633 (N_8633,N_7483,N_7069);
nor U8634 (N_8634,N_7608,N_7281);
or U8635 (N_8635,N_7284,N_7729);
nor U8636 (N_8636,N_7616,N_7574);
and U8637 (N_8637,N_7912,N_7653);
nor U8638 (N_8638,N_7207,N_7162);
xor U8639 (N_8639,N_7440,N_7790);
xor U8640 (N_8640,N_7861,N_7991);
xnor U8641 (N_8641,N_7597,N_7944);
or U8642 (N_8642,N_7514,N_7521);
or U8643 (N_8643,N_7631,N_7038);
nand U8644 (N_8644,N_7618,N_7097);
nand U8645 (N_8645,N_7939,N_7583);
and U8646 (N_8646,N_7078,N_7544);
xnor U8647 (N_8647,N_7130,N_7601);
nand U8648 (N_8648,N_7721,N_7300);
xor U8649 (N_8649,N_7372,N_7894);
nand U8650 (N_8650,N_7706,N_7272);
nand U8651 (N_8651,N_7227,N_7625);
and U8652 (N_8652,N_7957,N_7154);
nor U8653 (N_8653,N_7431,N_7649);
nor U8654 (N_8654,N_7968,N_7765);
nand U8655 (N_8655,N_7780,N_7186);
nand U8656 (N_8656,N_7050,N_7377);
xnor U8657 (N_8657,N_7193,N_7601);
or U8658 (N_8658,N_7004,N_7080);
or U8659 (N_8659,N_7455,N_7808);
nor U8660 (N_8660,N_7599,N_7779);
nor U8661 (N_8661,N_7039,N_7090);
nand U8662 (N_8662,N_7001,N_7649);
nor U8663 (N_8663,N_7123,N_7707);
xnor U8664 (N_8664,N_7469,N_7356);
and U8665 (N_8665,N_7521,N_7687);
nor U8666 (N_8666,N_7909,N_7877);
and U8667 (N_8667,N_7894,N_7026);
xnor U8668 (N_8668,N_7772,N_7677);
or U8669 (N_8669,N_7785,N_7646);
nand U8670 (N_8670,N_7509,N_7401);
and U8671 (N_8671,N_7780,N_7188);
nor U8672 (N_8672,N_7121,N_7813);
nand U8673 (N_8673,N_7883,N_7388);
xor U8674 (N_8674,N_7773,N_7461);
nand U8675 (N_8675,N_7395,N_7170);
nor U8676 (N_8676,N_7779,N_7104);
nor U8677 (N_8677,N_7204,N_7388);
nor U8678 (N_8678,N_7337,N_7238);
or U8679 (N_8679,N_7411,N_7453);
and U8680 (N_8680,N_7546,N_7765);
nor U8681 (N_8681,N_7772,N_7465);
or U8682 (N_8682,N_7930,N_7400);
xor U8683 (N_8683,N_7180,N_7659);
nand U8684 (N_8684,N_7612,N_7425);
nand U8685 (N_8685,N_7732,N_7922);
or U8686 (N_8686,N_7542,N_7517);
or U8687 (N_8687,N_7126,N_7206);
nand U8688 (N_8688,N_7691,N_7599);
or U8689 (N_8689,N_7802,N_7832);
xor U8690 (N_8690,N_7826,N_7579);
and U8691 (N_8691,N_7532,N_7518);
nand U8692 (N_8692,N_7578,N_7369);
xnor U8693 (N_8693,N_7141,N_7613);
and U8694 (N_8694,N_7447,N_7726);
nand U8695 (N_8695,N_7196,N_7405);
or U8696 (N_8696,N_7203,N_7172);
nand U8697 (N_8697,N_7072,N_7504);
and U8698 (N_8698,N_7392,N_7612);
and U8699 (N_8699,N_7928,N_7227);
or U8700 (N_8700,N_7570,N_7281);
nor U8701 (N_8701,N_7033,N_7172);
and U8702 (N_8702,N_7207,N_7364);
or U8703 (N_8703,N_7098,N_7438);
and U8704 (N_8704,N_7974,N_7350);
or U8705 (N_8705,N_7674,N_7999);
nand U8706 (N_8706,N_7395,N_7642);
and U8707 (N_8707,N_7870,N_7627);
or U8708 (N_8708,N_7835,N_7685);
or U8709 (N_8709,N_7409,N_7815);
and U8710 (N_8710,N_7089,N_7478);
xor U8711 (N_8711,N_7615,N_7943);
xnor U8712 (N_8712,N_7470,N_7335);
nand U8713 (N_8713,N_7914,N_7832);
and U8714 (N_8714,N_7883,N_7284);
nor U8715 (N_8715,N_7372,N_7088);
or U8716 (N_8716,N_7556,N_7943);
and U8717 (N_8717,N_7476,N_7854);
nor U8718 (N_8718,N_7125,N_7646);
or U8719 (N_8719,N_7478,N_7692);
nor U8720 (N_8720,N_7876,N_7603);
or U8721 (N_8721,N_7884,N_7116);
and U8722 (N_8722,N_7405,N_7690);
nor U8723 (N_8723,N_7455,N_7710);
xnor U8724 (N_8724,N_7518,N_7334);
nand U8725 (N_8725,N_7397,N_7531);
xnor U8726 (N_8726,N_7192,N_7791);
and U8727 (N_8727,N_7323,N_7274);
xnor U8728 (N_8728,N_7832,N_7179);
nand U8729 (N_8729,N_7724,N_7700);
or U8730 (N_8730,N_7344,N_7957);
nand U8731 (N_8731,N_7378,N_7076);
nand U8732 (N_8732,N_7751,N_7444);
nor U8733 (N_8733,N_7208,N_7149);
and U8734 (N_8734,N_7286,N_7630);
xor U8735 (N_8735,N_7585,N_7832);
nand U8736 (N_8736,N_7775,N_7117);
nand U8737 (N_8737,N_7606,N_7647);
and U8738 (N_8738,N_7127,N_7876);
xor U8739 (N_8739,N_7708,N_7939);
nand U8740 (N_8740,N_7810,N_7750);
or U8741 (N_8741,N_7297,N_7269);
nand U8742 (N_8742,N_7403,N_7300);
nor U8743 (N_8743,N_7568,N_7550);
xnor U8744 (N_8744,N_7145,N_7009);
xor U8745 (N_8745,N_7749,N_7782);
xnor U8746 (N_8746,N_7255,N_7873);
or U8747 (N_8747,N_7809,N_7827);
and U8748 (N_8748,N_7927,N_7366);
nand U8749 (N_8749,N_7012,N_7403);
nand U8750 (N_8750,N_7120,N_7423);
nand U8751 (N_8751,N_7688,N_7672);
nor U8752 (N_8752,N_7801,N_7578);
or U8753 (N_8753,N_7047,N_7683);
or U8754 (N_8754,N_7341,N_7129);
or U8755 (N_8755,N_7216,N_7067);
nand U8756 (N_8756,N_7856,N_7001);
nand U8757 (N_8757,N_7159,N_7882);
nand U8758 (N_8758,N_7241,N_7470);
and U8759 (N_8759,N_7226,N_7683);
nand U8760 (N_8760,N_7989,N_7592);
nand U8761 (N_8761,N_7028,N_7408);
nand U8762 (N_8762,N_7570,N_7008);
and U8763 (N_8763,N_7931,N_7433);
nor U8764 (N_8764,N_7639,N_7485);
and U8765 (N_8765,N_7908,N_7181);
or U8766 (N_8766,N_7911,N_7876);
xnor U8767 (N_8767,N_7305,N_7209);
xor U8768 (N_8768,N_7497,N_7675);
nand U8769 (N_8769,N_7386,N_7475);
nand U8770 (N_8770,N_7670,N_7905);
nand U8771 (N_8771,N_7733,N_7151);
xor U8772 (N_8772,N_7609,N_7255);
nor U8773 (N_8773,N_7985,N_7350);
nor U8774 (N_8774,N_7690,N_7962);
and U8775 (N_8775,N_7955,N_7202);
nor U8776 (N_8776,N_7098,N_7926);
or U8777 (N_8777,N_7655,N_7050);
nand U8778 (N_8778,N_7634,N_7951);
and U8779 (N_8779,N_7701,N_7663);
nand U8780 (N_8780,N_7277,N_7142);
nand U8781 (N_8781,N_7607,N_7938);
and U8782 (N_8782,N_7776,N_7648);
and U8783 (N_8783,N_7235,N_7773);
nand U8784 (N_8784,N_7814,N_7594);
nand U8785 (N_8785,N_7964,N_7546);
xnor U8786 (N_8786,N_7240,N_7982);
and U8787 (N_8787,N_7534,N_7179);
xnor U8788 (N_8788,N_7354,N_7330);
and U8789 (N_8789,N_7683,N_7958);
nand U8790 (N_8790,N_7045,N_7662);
nor U8791 (N_8791,N_7044,N_7327);
xnor U8792 (N_8792,N_7043,N_7076);
nor U8793 (N_8793,N_7205,N_7159);
or U8794 (N_8794,N_7032,N_7054);
nand U8795 (N_8795,N_7548,N_7152);
and U8796 (N_8796,N_7488,N_7154);
or U8797 (N_8797,N_7310,N_7821);
and U8798 (N_8798,N_7458,N_7549);
or U8799 (N_8799,N_7947,N_7023);
nor U8800 (N_8800,N_7704,N_7117);
xnor U8801 (N_8801,N_7484,N_7065);
nand U8802 (N_8802,N_7505,N_7186);
and U8803 (N_8803,N_7555,N_7176);
nand U8804 (N_8804,N_7226,N_7606);
nand U8805 (N_8805,N_7309,N_7618);
nor U8806 (N_8806,N_7456,N_7608);
nand U8807 (N_8807,N_7070,N_7800);
nor U8808 (N_8808,N_7449,N_7963);
nor U8809 (N_8809,N_7390,N_7166);
or U8810 (N_8810,N_7250,N_7864);
nand U8811 (N_8811,N_7634,N_7225);
or U8812 (N_8812,N_7586,N_7417);
and U8813 (N_8813,N_7084,N_7821);
nor U8814 (N_8814,N_7860,N_7252);
nand U8815 (N_8815,N_7847,N_7007);
xor U8816 (N_8816,N_7478,N_7322);
xnor U8817 (N_8817,N_7943,N_7088);
nand U8818 (N_8818,N_7857,N_7741);
xnor U8819 (N_8819,N_7148,N_7521);
xor U8820 (N_8820,N_7819,N_7444);
nand U8821 (N_8821,N_7671,N_7293);
nor U8822 (N_8822,N_7668,N_7101);
or U8823 (N_8823,N_7290,N_7361);
or U8824 (N_8824,N_7384,N_7342);
nand U8825 (N_8825,N_7543,N_7795);
nor U8826 (N_8826,N_7670,N_7534);
nor U8827 (N_8827,N_7234,N_7251);
nand U8828 (N_8828,N_7633,N_7193);
and U8829 (N_8829,N_7408,N_7795);
and U8830 (N_8830,N_7764,N_7688);
nand U8831 (N_8831,N_7941,N_7635);
nand U8832 (N_8832,N_7141,N_7349);
or U8833 (N_8833,N_7526,N_7840);
and U8834 (N_8834,N_7541,N_7708);
or U8835 (N_8835,N_7744,N_7244);
xor U8836 (N_8836,N_7280,N_7366);
nand U8837 (N_8837,N_7879,N_7158);
nor U8838 (N_8838,N_7737,N_7562);
xor U8839 (N_8839,N_7307,N_7208);
xnor U8840 (N_8840,N_7409,N_7191);
xnor U8841 (N_8841,N_7120,N_7072);
nand U8842 (N_8842,N_7987,N_7989);
nand U8843 (N_8843,N_7673,N_7888);
and U8844 (N_8844,N_7309,N_7948);
nand U8845 (N_8845,N_7072,N_7247);
nand U8846 (N_8846,N_7315,N_7224);
nand U8847 (N_8847,N_7263,N_7101);
and U8848 (N_8848,N_7632,N_7000);
or U8849 (N_8849,N_7541,N_7564);
nand U8850 (N_8850,N_7476,N_7101);
nor U8851 (N_8851,N_7995,N_7337);
and U8852 (N_8852,N_7012,N_7107);
nor U8853 (N_8853,N_7792,N_7045);
nand U8854 (N_8854,N_7595,N_7839);
nor U8855 (N_8855,N_7267,N_7469);
nand U8856 (N_8856,N_7294,N_7710);
nand U8857 (N_8857,N_7472,N_7621);
xnor U8858 (N_8858,N_7569,N_7087);
or U8859 (N_8859,N_7133,N_7430);
xnor U8860 (N_8860,N_7415,N_7336);
or U8861 (N_8861,N_7342,N_7674);
nand U8862 (N_8862,N_7283,N_7258);
nand U8863 (N_8863,N_7230,N_7967);
and U8864 (N_8864,N_7805,N_7823);
or U8865 (N_8865,N_7820,N_7278);
nor U8866 (N_8866,N_7356,N_7656);
nand U8867 (N_8867,N_7571,N_7818);
and U8868 (N_8868,N_7631,N_7740);
nand U8869 (N_8869,N_7818,N_7183);
xor U8870 (N_8870,N_7793,N_7235);
or U8871 (N_8871,N_7517,N_7729);
xor U8872 (N_8872,N_7542,N_7668);
nor U8873 (N_8873,N_7652,N_7943);
or U8874 (N_8874,N_7059,N_7165);
nor U8875 (N_8875,N_7443,N_7762);
nand U8876 (N_8876,N_7725,N_7252);
and U8877 (N_8877,N_7417,N_7787);
or U8878 (N_8878,N_7659,N_7278);
xor U8879 (N_8879,N_7737,N_7286);
xor U8880 (N_8880,N_7968,N_7094);
or U8881 (N_8881,N_7485,N_7468);
and U8882 (N_8882,N_7971,N_7699);
or U8883 (N_8883,N_7075,N_7653);
or U8884 (N_8884,N_7536,N_7431);
or U8885 (N_8885,N_7521,N_7500);
nand U8886 (N_8886,N_7557,N_7870);
nor U8887 (N_8887,N_7756,N_7509);
xnor U8888 (N_8888,N_7853,N_7534);
and U8889 (N_8889,N_7018,N_7187);
nor U8890 (N_8890,N_7996,N_7942);
xor U8891 (N_8891,N_7437,N_7266);
nor U8892 (N_8892,N_7638,N_7694);
xor U8893 (N_8893,N_7058,N_7965);
nand U8894 (N_8894,N_7165,N_7013);
or U8895 (N_8895,N_7438,N_7982);
xor U8896 (N_8896,N_7781,N_7383);
nor U8897 (N_8897,N_7872,N_7384);
or U8898 (N_8898,N_7165,N_7311);
and U8899 (N_8899,N_7064,N_7474);
nand U8900 (N_8900,N_7958,N_7448);
nor U8901 (N_8901,N_7443,N_7655);
nor U8902 (N_8902,N_7007,N_7005);
nand U8903 (N_8903,N_7009,N_7030);
and U8904 (N_8904,N_7505,N_7273);
xor U8905 (N_8905,N_7947,N_7818);
nor U8906 (N_8906,N_7112,N_7629);
and U8907 (N_8907,N_7918,N_7566);
and U8908 (N_8908,N_7060,N_7635);
and U8909 (N_8909,N_7935,N_7301);
or U8910 (N_8910,N_7685,N_7405);
nand U8911 (N_8911,N_7557,N_7617);
or U8912 (N_8912,N_7400,N_7061);
nor U8913 (N_8913,N_7128,N_7763);
and U8914 (N_8914,N_7341,N_7438);
nor U8915 (N_8915,N_7965,N_7756);
xnor U8916 (N_8916,N_7582,N_7167);
nand U8917 (N_8917,N_7564,N_7860);
xnor U8918 (N_8918,N_7734,N_7653);
nor U8919 (N_8919,N_7268,N_7682);
or U8920 (N_8920,N_7998,N_7581);
xnor U8921 (N_8921,N_7619,N_7427);
nand U8922 (N_8922,N_7323,N_7437);
xor U8923 (N_8923,N_7602,N_7568);
nand U8924 (N_8924,N_7888,N_7747);
nand U8925 (N_8925,N_7197,N_7095);
and U8926 (N_8926,N_7558,N_7798);
or U8927 (N_8927,N_7929,N_7415);
or U8928 (N_8928,N_7175,N_7994);
xnor U8929 (N_8929,N_7717,N_7589);
or U8930 (N_8930,N_7396,N_7845);
nor U8931 (N_8931,N_7442,N_7312);
nand U8932 (N_8932,N_7639,N_7720);
xnor U8933 (N_8933,N_7673,N_7362);
xor U8934 (N_8934,N_7643,N_7260);
or U8935 (N_8935,N_7167,N_7436);
nand U8936 (N_8936,N_7352,N_7200);
nor U8937 (N_8937,N_7496,N_7975);
and U8938 (N_8938,N_7424,N_7168);
and U8939 (N_8939,N_7252,N_7402);
and U8940 (N_8940,N_7656,N_7316);
nand U8941 (N_8941,N_7099,N_7384);
or U8942 (N_8942,N_7282,N_7433);
nand U8943 (N_8943,N_7504,N_7750);
nor U8944 (N_8944,N_7197,N_7256);
or U8945 (N_8945,N_7151,N_7891);
and U8946 (N_8946,N_7114,N_7222);
xor U8947 (N_8947,N_7954,N_7590);
nor U8948 (N_8948,N_7134,N_7173);
or U8949 (N_8949,N_7953,N_7150);
and U8950 (N_8950,N_7735,N_7912);
and U8951 (N_8951,N_7628,N_7267);
and U8952 (N_8952,N_7987,N_7257);
or U8953 (N_8953,N_7557,N_7251);
nand U8954 (N_8954,N_7087,N_7059);
nor U8955 (N_8955,N_7097,N_7392);
or U8956 (N_8956,N_7158,N_7700);
and U8957 (N_8957,N_7906,N_7544);
nand U8958 (N_8958,N_7096,N_7793);
and U8959 (N_8959,N_7136,N_7912);
nor U8960 (N_8960,N_7240,N_7886);
or U8961 (N_8961,N_7531,N_7563);
nand U8962 (N_8962,N_7132,N_7541);
or U8963 (N_8963,N_7022,N_7540);
nand U8964 (N_8964,N_7514,N_7773);
nor U8965 (N_8965,N_7309,N_7210);
xor U8966 (N_8966,N_7529,N_7134);
or U8967 (N_8967,N_7386,N_7203);
and U8968 (N_8968,N_7535,N_7590);
or U8969 (N_8969,N_7845,N_7945);
or U8970 (N_8970,N_7033,N_7765);
nand U8971 (N_8971,N_7946,N_7434);
nor U8972 (N_8972,N_7067,N_7378);
or U8973 (N_8973,N_7892,N_7121);
and U8974 (N_8974,N_7062,N_7075);
and U8975 (N_8975,N_7185,N_7120);
nand U8976 (N_8976,N_7243,N_7073);
nor U8977 (N_8977,N_7377,N_7510);
nor U8978 (N_8978,N_7452,N_7922);
nand U8979 (N_8979,N_7966,N_7386);
nor U8980 (N_8980,N_7625,N_7520);
or U8981 (N_8981,N_7007,N_7715);
xnor U8982 (N_8982,N_7865,N_7706);
nor U8983 (N_8983,N_7245,N_7021);
nor U8984 (N_8984,N_7278,N_7014);
or U8985 (N_8985,N_7751,N_7284);
and U8986 (N_8986,N_7877,N_7481);
nor U8987 (N_8987,N_7405,N_7901);
and U8988 (N_8988,N_7589,N_7509);
or U8989 (N_8989,N_7933,N_7935);
or U8990 (N_8990,N_7651,N_7729);
and U8991 (N_8991,N_7301,N_7287);
nand U8992 (N_8992,N_7936,N_7513);
xnor U8993 (N_8993,N_7676,N_7971);
nand U8994 (N_8994,N_7578,N_7334);
or U8995 (N_8995,N_7267,N_7424);
and U8996 (N_8996,N_7054,N_7152);
or U8997 (N_8997,N_7716,N_7347);
nand U8998 (N_8998,N_7502,N_7091);
nand U8999 (N_8999,N_7482,N_7867);
xor U9000 (N_9000,N_8663,N_8813);
xor U9001 (N_9001,N_8679,N_8733);
nand U9002 (N_9002,N_8427,N_8062);
or U9003 (N_9003,N_8880,N_8218);
nor U9004 (N_9004,N_8982,N_8351);
and U9005 (N_9005,N_8752,N_8220);
nor U9006 (N_9006,N_8026,N_8369);
or U9007 (N_9007,N_8998,N_8658);
xnor U9008 (N_9008,N_8418,N_8484);
or U9009 (N_9009,N_8232,N_8595);
and U9010 (N_9010,N_8629,N_8670);
xor U9011 (N_9011,N_8296,N_8394);
nor U9012 (N_9012,N_8977,N_8108);
or U9013 (N_9013,N_8975,N_8107);
and U9014 (N_9014,N_8567,N_8959);
or U9015 (N_9015,N_8326,N_8947);
nand U9016 (N_9016,N_8362,N_8198);
or U9017 (N_9017,N_8417,N_8028);
xnor U9018 (N_9018,N_8970,N_8916);
nor U9019 (N_9019,N_8129,N_8908);
or U9020 (N_9020,N_8065,N_8978);
nor U9021 (N_9021,N_8926,N_8050);
and U9022 (N_9022,N_8823,N_8954);
xnor U9023 (N_9023,N_8797,N_8105);
and U9024 (N_9024,N_8973,N_8481);
nor U9025 (N_9025,N_8447,N_8084);
nand U9026 (N_9026,N_8780,N_8127);
xor U9027 (N_9027,N_8390,N_8546);
and U9028 (N_9028,N_8816,N_8715);
nor U9029 (N_9029,N_8821,N_8933);
xor U9030 (N_9030,N_8535,N_8718);
nand U9031 (N_9031,N_8339,N_8864);
xor U9032 (N_9032,N_8126,N_8958);
nand U9033 (N_9033,N_8385,N_8138);
nor U9034 (N_9034,N_8689,N_8241);
nor U9035 (N_9035,N_8896,N_8153);
and U9036 (N_9036,N_8361,N_8005);
and U9037 (N_9037,N_8805,N_8645);
and U9038 (N_9038,N_8726,N_8937);
and U9039 (N_9039,N_8125,N_8891);
or U9040 (N_9040,N_8332,N_8782);
nand U9041 (N_9041,N_8955,N_8435);
and U9042 (N_9042,N_8486,N_8239);
and U9043 (N_9043,N_8961,N_8490);
and U9044 (N_9044,N_8375,N_8191);
and U9045 (N_9045,N_8568,N_8651);
and U9046 (N_9046,N_8060,N_8646);
xnor U9047 (N_9047,N_8628,N_8301);
or U9048 (N_9048,N_8288,N_8969);
or U9049 (N_9049,N_8291,N_8506);
nor U9050 (N_9050,N_8251,N_8092);
nor U9051 (N_9051,N_8921,N_8193);
xor U9052 (N_9052,N_8335,N_8158);
nand U9053 (N_9053,N_8799,N_8470);
xor U9054 (N_9054,N_8465,N_8397);
or U9055 (N_9055,N_8521,N_8340);
or U9056 (N_9056,N_8063,N_8936);
nand U9057 (N_9057,N_8162,N_8508);
or U9058 (N_9058,N_8620,N_8745);
nor U9059 (N_9059,N_8684,N_8210);
nor U9060 (N_9060,N_8184,N_8479);
nand U9061 (N_9061,N_8401,N_8565);
or U9062 (N_9062,N_8122,N_8355);
xnor U9063 (N_9063,N_8284,N_8830);
or U9064 (N_9064,N_8824,N_8110);
and U9065 (N_9065,N_8386,N_8793);
or U9066 (N_9066,N_8650,N_8990);
and U9067 (N_9067,N_8017,N_8784);
or U9068 (N_9068,N_8913,N_8669);
xnor U9069 (N_9069,N_8530,N_8734);
xnor U9070 (N_9070,N_8139,N_8558);
and U9071 (N_9071,N_8308,N_8250);
xnor U9072 (N_9072,N_8133,N_8163);
and U9073 (N_9073,N_8403,N_8722);
or U9074 (N_9074,N_8619,N_8080);
and U9075 (N_9075,N_8667,N_8269);
nor U9076 (N_9076,N_8132,N_8573);
nand U9077 (N_9077,N_8875,N_8614);
nand U9078 (N_9078,N_8388,N_8203);
xnor U9079 (N_9079,N_8898,N_8421);
and U9080 (N_9080,N_8211,N_8069);
or U9081 (N_9081,N_8588,N_8756);
or U9082 (N_9082,N_8295,N_8770);
nor U9083 (N_9083,N_8474,N_8795);
nand U9084 (N_9084,N_8687,N_8324);
xnor U9085 (N_9085,N_8141,N_8984);
and U9086 (N_9086,N_8399,N_8703);
and U9087 (N_9087,N_8807,N_8980);
and U9088 (N_9088,N_8999,N_8837);
nand U9089 (N_9089,N_8556,N_8425);
nand U9090 (N_9090,N_8605,N_8789);
or U9091 (N_9091,N_8720,N_8016);
xor U9092 (N_9092,N_8216,N_8409);
or U9093 (N_9093,N_8723,N_8466);
xnor U9094 (N_9094,N_8102,N_8111);
xor U9095 (N_9095,N_8836,N_8278);
and U9096 (N_9096,N_8510,N_8130);
nand U9097 (N_9097,N_8047,N_8753);
or U9098 (N_9098,N_8682,N_8443);
nand U9099 (N_9099,N_8121,N_8819);
nand U9100 (N_9100,N_8603,N_8685);
and U9101 (N_9101,N_8249,N_8828);
nand U9102 (N_9102,N_8087,N_8265);
and U9103 (N_9103,N_8539,N_8923);
xnor U9104 (N_9104,N_8072,N_8621);
nand U9105 (N_9105,N_8011,N_8302);
xnor U9106 (N_9106,N_8070,N_8634);
xnor U9107 (N_9107,N_8438,N_8440);
or U9108 (N_9108,N_8095,N_8380);
xnor U9109 (N_9109,N_8676,N_8328);
nand U9110 (N_9110,N_8030,N_8106);
and U9111 (N_9111,N_8454,N_8849);
nand U9112 (N_9112,N_8238,N_8868);
xor U9113 (N_9113,N_8648,N_8766);
and U9114 (N_9114,N_8613,N_8342);
nor U9115 (N_9115,N_8548,N_8176);
and U9116 (N_9116,N_8654,N_8117);
nand U9117 (N_9117,N_8177,N_8119);
or U9118 (N_9118,N_8825,N_8943);
or U9119 (N_9119,N_8960,N_8349);
and U9120 (N_9120,N_8416,N_8792);
or U9121 (N_9121,N_8845,N_8590);
nor U9122 (N_9122,N_8895,N_8516);
and U9123 (N_9123,N_8839,N_8275);
nor U9124 (N_9124,N_8915,N_8639);
xnor U9125 (N_9125,N_8396,N_8333);
nor U9126 (N_9126,N_8195,N_8578);
nor U9127 (N_9127,N_8496,N_8584);
xor U9128 (N_9128,N_8346,N_8777);
and U9129 (N_9129,N_8509,N_8909);
nor U9130 (N_9130,N_8967,N_8116);
xnor U9131 (N_9131,N_8609,N_8901);
or U9132 (N_9132,N_8754,N_8531);
nand U9133 (N_9133,N_8931,N_8870);
xor U9134 (N_9134,N_8366,N_8000);
xor U9135 (N_9135,N_8147,N_8817);
nand U9136 (N_9136,N_8897,N_8692);
xnor U9137 (N_9137,N_8906,N_8304);
and U9138 (N_9138,N_8927,N_8942);
and U9139 (N_9139,N_8744,N_8529);
nand U9140 (N_9140,N_8404,N_8693);
and U9141 (N_9141,N_8489,N_8174);
nor U9142 (N_9142,N_8932,N_8918);
nor U9143 (N_9143,N_8449,N_8230);
or U9144 (N_9144,N_8320,N_8061);
nor U9145 (N_9145,N_8538,N_8233);
and U9146 (N_9146,N_8156,N_8665);
nand U9147 (N_9147,N_8844,N_8307);
nor U9148 (N_9148,N_8091,N_8525);
or U9149 (N_9149,N_8809,N_8109);
nand U9150 (N_9150,N_8379,N_8790);
or U9151 (N_9151,N_8869,N_8058);
or U9152 (N_9152,N_8701,N_8096);
xor U9153 (N_9153,N_8704,N_8501);
and U9154 (N_9154,N_8576,N_8928);
nor U9155 (N_9155,N_8995,N_8169);
or U9156 (N_9156,N_8219,N_8422);
and U9157 (N_9157,N_8019,N_8053);
or U9158 (N_9158,N_8575,N_8965);
nand U9159 (N_9159,N_8951,N_8491);
nor U9160 (N_9160,N_8165,N_8175);
xor U9161 (N_9161,N_8264,N_8635);
nor U9162 (N_9162,N_8006,N_8444);
nor U9163 (N_9163,N_8405,N_8245);
nand U9164 (N_9164,N_8524,N_8456);
and U9165 (N_9165,N_8631,N_8852);
xor U9166 (N_9166,N_8820,N_8929);
and U9167 (N_9167,N_8100,N_8647);
nor U9168 (N_9168,N_8043,N_8788);
xnor U9169 (N_9169,N_8856,N_8183);
nand U9170 (N_9170,N_8157,N_8851);
or U9171 (N_9171,N_8545,N_8323);
nand U9172 (N_9172,N_8741,N_8601);
or U9173 (N_9173,N_8561,N_8261);
nor U9174 (N_9174,N_8123,N_8772);
xor U9175 (N_9175,N_8451,N_8585);
and U9176 (N_9176,N_8981,N_8315);
and U9177 (N_9177,N_8549,N_8757);
or U9178 (N_9178,N_8476,N_8986);
or U9179 (N_9179,N_8318,N_8112);
nand U9180 (N_9180,N_8415,N_8972);
nand U9181 (N_9181,N_8583,N_8306);
and U9182 (N_9182,N_8725,N_8528);
and U9183 (N_9183,N_8794,N_8207);
nand U9184 (N_9184,N_8542,N_8433);
nand U9185 (N_9185,N_8483,N_8786);
nor U9186 (N_9186,N_8886,N_8336);
nor U9187 (N_9187,N_8755,N_8137);
nor U9188 (N_9188,N_8957,N_8262);
and U9189 (N_9189,N_8463,N_8426);
xor U9190 (N_9190,N_8638,N_8468);
and U9191 (N_9191,N_8493,N_8858);
and U9192 (N_9192,N_8767,N_8768);
and U9193 (N_9193,N_8518,N_8464);
nor U9194 (N_9194,N_8395,N_8142);
nand U9195 (N_9195,N_8268,N_8254);
xnor U9196 (N_9196,N_8337,N_8334);
and U9197 (N_9197,N_8010,N_8724);
xnor U9198 (N_9198,N_8159,N_8325);
or U9199 (N_9199,N_8796,N_8672);
nor U9200 (N_9200,N_8729,N_8146);
nor U9201 (N_9201,N_8237,N_8271);
xnor U9202 (N_9202,N_8452,N_8743);
nand U9203 (N_9203,N_8553,N_8900);
nor U9204 (N_9204,N_8376,N_8370);
xnor U9205 (N_9205,N_8758,N_8534);
nand U9206 (N_9206,N_8012,N_8423);
or U9207 (N_9207,N_8559,N_8407);
xnor U9208 (N_9208,N_8511,N_8290);
or U9209 (N_9209,N_8359,N_8469);
xnor U9210 (N_9210,N_8574,N_8044);
xnor U9211 (N_9211,N_8419,N_8267);
nor U9212 (N_9212,N_8659,N_8083);
or U9213 (N_9213,N_8094,N_8702);
and U9214 (N_9214,N_8231,N_8987);
or U9215 (N_9215,N_8074,N_8101);
nand U9216 (N_9216,N_8617,N_8877);
xor U9217 (N_9217,N_8537,N_8683);
or U9218 (N_9218,N_8746,N_8356);
xor U9219 (N_9219,N_8103,N_8289);
nand U9220 (N_9220,N_8874,N_8800);
or U9221 (N_9221,N_8167,N_8081);
nand U9222 (N_9222,N_8666,N_8907);
nor U9223 (N_9223,N_8367,N_8164);
and U9224 (N_9224,N_8991,N_8114);
nor U9225 (N_9225,N_8077,N_8208);
or U9226 (N_9226,N_8607,N_8277);
nor U9227 (N_9227,N_8602,N_8042);
xnor U9228 (N_9228,N_8205,N_8360);
or U9229 (N_9229,N_8507,N_8656);
or U9230 (N_9230,N_8482,N_8675);
nand U9231 (N_9231,N_8352,N_8892);
or U9232 (N_9232,N_8013,N_8018);
or U9233 (N_9233,N_8783,N_8652);
nor U9234 (N_9234,N_8850,N_8007);
xor U9235 (N_9235,N_8618,N_8150);
and U9236 (N_9236,N_8387,N_8624);
nand U9237 (N_9237,N_8041,N_8505);
and U9238 (N_9238,N_8696,N_8344);
xnor U9239 (N_9239,N_8597,N_8866);
nand U9240 (N_9240,N_8170,N_8075);
or U9241 (N_9241,N_8544,N_8917);
xnor U9242 (N_9242,N_8616,N_8188);
nor U9243 (N_9243,N_8668,N_8441);
nand U9244 (N_9244,N_8023,N_8252);
xnor U9245 (N_9245,N_8434,N_8637);
and U9246 (N_9246,N_8774,N_8562);
xnor U9247 (N_9247,N_8365,N_8750);
nand U9248 (N_9248,N_8941,N_8678);
nand U9249 (N_9249,N_8118,N_8128);
nor U9250 (N_9250,N_8855,N_8270);
and U9251 (N_9251,N_8467,N_8214);
or U9252 (N_9252,N_8078,N_8178);
nor U9253 (N_9253,N_8206,N_8363);
xnor U9254 (N_9254,N_8912,N_8717);
and U9255 (N_9255,N_8771,N_8259);
nand U9256 (N_9256,N_8009,N_8381);
xnor U9257 (N_9257,N_8377,N_8492);
or U9258 (N_9258,N_8186,N_8226);
nand U9259 (N_9259,N_8950,N_8168);
and U9260 (N_9260,N_8348,N_8229);
xnor U9261 (N_9261,N_8499,N_8217);
or U9262 (N_9262,N_8460,N_8563);
xor U9263 (N_9263,N_8697,N_8925);
nor U9264 (N_9264,N_8842,N_8504);
xor U9265 (N_9265,N_8622,N_8329);
xor U9266 (N_9266,N_8389,N_8861);
and U9267 (N_9267,N_8136,N_8341);
or U9268 (N_9268,N_8224,N_8455);
xnor U9269 (N_9269,N_8256,N_8610);
nand U9270 (N_9270,N_8731,N_8657);
nand U9271 (N_9271,N_8580,N_8904);
xnor U9272 (N_9272,N_8046,N_8402);
nand U9273 (N_9273,N_8632,N_8343);
nor U9274 (N_9274,N_8579,N_8458);
xnor U9275 (N_9275,N_8640,N_8930);
nor U9276 (N_9276,N_8974,N_8773);
nand U9277 (N_9277,N_8812,N_8257);
xor U9278 (N_9278,N_8688,N_8079);
nor U9279 (N_9279,N_8759,N_8453);
or U9280 (N_9280,N_8826,N_8643);
xor U9281 (N_9281,N_8098,N_8939);
nand U9282 (N_9282,N_8694,N_8462);
and U9283 (N_9283,N_8964,N_8283);
nor U9284 (N_9284,N_8540,N_8709);
and U9285 (N_9285,N_8225,N_8089);
or U9286 (N_9286,N_8700,N_8594);
xnor U9287 (N_9287,N_8393,N_8354);
xnor U9288 (N_9288,N_8410,N_8899);
or U9289 (N_9289,N_8699,N_8276);
xnor U9290 (N_9290,N_8330,N_8803);
nand U9291 (N_9291,N_8215,N_8073);
and U9292 (N_9292,N_8680,N_8526);
xor U9293 (N_9293,N_8644,N_8246);
nand U9294 (N_9294,N_8591,N_8242);
nand U9295 (N_9295,N_8949,N_8272);
nor U9296 (N_9296,N_8714,N_8992);
xor U9297 (N_9297,N_8829,N_8835);
xor U9298 (N_9298,N_8885,N_8151);
nand U9299 (N_9299,N_8520,N_8764);
or U9300 (N_9300,N_8626,N_8979);
xnor U9301 (N_9301,N_8873,N_8171);
and U9302 (N_9302,N_8124,N_8134);
or U9303 (N_9303,N_8884,N_8582);
xor U9304 (N_9304,N_8384,N_8003);
or U9305 (N_9305,N_8732,N_8478);
nor U9306 (N_9306,N_8442,N_8924);
or U9307 (N_9307,N_8513,N_8867);
or U9308 (N_9308,N_8876,N_8748);
and U9309 (N_9309,N_8189,N_8309);
nand U9310 (N_9310,N_8859,N_8299);
xnor U9311 (N_9311,N_8555,N_8515);
nor U9312 (N_9312,N_8038,N_8934);
or U9313 (N_9313,N_8814,N_8287);
xnor U9314 (N_9314,N_8681,N_8586);
xor U9315 (N_9315,N_8708,N_8775);
or U9316 (N_9316,N_8331,N_8946);
nand U9317 (N_9317,N_8552,N_8808);
and U9318 (N_9318,N_8727,N_8001);
nand U9319 (N_9319,N_8413,N_8199);
or U9320 (N_9320,N_8040,N_8194);
nand U9321 (N_9321,N_8940,N_8671);
and U9322 (N_9322,N_8893,N_8910);
or U9323 (N_9323,N_8707,N_8067);
xor U9324 (N_9324,N_8636,N_8022);
or U9325 (N_9325,N_8374,N_8461);
nand U9326 (N_9326,N_8751,N_8185);
nand U9327 (N_9327,N_8778,N_8633);
nor U9328 (N_9328,N_8204,N_8604);
and U9329 (N_9329,N_8662,N_8840);
or U9330 (N_9330,N_8804,N_8033);
nand U9331 (N_9331,N_8512,N_8321);
or U9332 (N_9332,N_8414,N_8457);
nor U9333 (N_9333,N_8378,N_8255);
or U9334 (N_9334,N_8625,N_8446);
xor U9335 (N_9335,N_8742,N_8922);
and U9336 (N_9336,N_8201,N_8313);
xnor U9337 (N_9337,N_8408,N_8522);
or U9338 (N_9338,N_8577,N_8311);
and U9339 (N_9339,N_8785,N_8762);
nand U9340 (N_9340,N_8948,N_8068);
and U9341 (N_9341,N_8052,N_8160);
or U9342 (N_9342,N_8316,N_8314);
or U9343 (N_9343,N_8459,N_8533);
nor U9344 (N_9344,N_8223,N_8878);
nor U9345 (N_9345,N_8487,N_8822);
nor U9346 (N_9346,N_8432,N_8879);
and U9347 (N_9347,N_8350,N_8076);
xor U9348 (N_9348,N_8905,N_8547);
and U9349 (N_9349,N_8902,N_8247);
nor U9350 (N_9350,N_8082,N_8935);
or U9351 (N_9351,N_8993,N_8623);
nand U9352 (N_9352,N_8273,N_8541);
nor U9353 (N_9353,N_8810,N_8115);
nand U9354 (N_9354,N_8391,N_8192);
nand U9355 (N_9355,N_8345,N_8274);
nor U9356 (N_9356,N_8209,N_8202);
and U9357 (N_9357,N_8811,N_8887);
nor U9358 (N_9358,N_8860,N_8448);
or U9359 (N_9359,N_8029,N_8606);
and U9360 (N_9360,N_8698,N_8439);
xnor U9361 (N_9361,N_8227,N_8503);
nand U9362 (N_9362,N_8894,N_8514);
and U9363 (N_9363,N_8719,N_8557);
nand U9364 (N_9364,N_8612,N_8711);
xor U9365 (N_9365,N_8347,N_8281);
nor U9366 (N_9366,N_8473,N_8570);
nor U9367 (N_9367,N_8004,N_8445);
xor U9368 (N_9368,N_8608,N_8471);
nand U9369 (N_9369,N_8180,N_8051);
nand U9370 (N_9370,N_8371,N_8236);
nand U9371 (N_9371,N_8920,N_8429);
nand U9372 (N_9372,N_8297,N_8412);
and U9373 (N_9373,N_8190,N_8914);
xor U9374 (N_9374,N_8155,N_8488);
nor U9375 (N_9375,N_8765,N_8056);
xor U9376 (N_9376,N_8266,N_8500);
and U9377 (N_9377,N_8587,N_8956);
xor U9378 (N_9378,N_8599,N_8021);
nand U9379 (N_9379,N_8818,N_8424);
and U9380 (N_9380,N_8364,N_8712);
or U9381 (N_9381,N_8104,N_8131);
or U9382 (N_9382,N_8495,N_8710);
nand U9383 (N_9383,N_8411,N_8066);
nand U9384 (N_9384,N_8550,N_8039);
and U9385 (N_9385,N_8596,N_8172);
or U9386 (N_9386,N_8057,N_8862);
nand U9387 (N_9387,N_8327,N_8228);
or U9388 (N_9388,N_8400,N_8686);
and U9389 (N_9389,N_8200,N_8560);
or U9390 (N_9390,N_8881,N_8593);
nor U9391 (N_9391,N_8853,N_8713);
nor U9392 (N_9392,N_8985,N_8801);
xnor U9393 (N_9393,N_8649,N_8034);
xnor U9394 (N_9394,N_8997,N_8292);
and U9395 (N_9395,N_8962,N_8589);
and U9396 (N_9396,N_8989,N_8234);
nand U9397 (N_9397,N_8747,N_8338);
nand U9398 (N_9398,N_8055,N_8600);
xor U9399 (N_9399,N_8598,N_8197);
or U9400 (N_9400,N_8032,N_8641);
and U9401 (N_9401,N_8838,N_8093);
nand U9402 (N_9402,N_8294,N_8258);
or U9403 (N_9403,N_8882,N_8085);
or U9404 (N_9404,N_8031,N_8730);
nor U9405 (N_9405,N_8863,N_8841);
or U9406 (N_9406,N_8564,N_8368);
nand U9407 (N_9407,N_8890,N_8615);
nand U9408 (N_9408,N_8145,N_8952);
and U9409 (N_9409,N_8406,N_8173);
nand U9410 (N_9410,N_8293,N_8353);
nor U9411 (N_9411,N_8398,N_8791);
nand U9412 (N_9412,N_8088,N_8166);
or U9413 (N_9413,N_8760,N_8502);
nand U9414 (N_9414,N_8148,N_8282);
xor U9415 (N_9415,N_8776,N_8739);
or U9416 (N_9416,N_8498,N_8317);
nor U9417 (N_9417,N_8736,N_8428);
nand U9418 (N_9418,N_8485,N_8472);
nand U9419 (N_9419,N_8944,N_8135);
or U9420 (N_9420,N_8036,N_8015);
nand U9421 (N_9421,N_8871,N_8235);
nand U9422 (N_9422,N_8140,N_8263);
and U9423 (N_9423,N_8431,N_8551);
or U9424 (N_9424,N_8420,N_8322);
nand U9425 (N_9425,N_8020,N_8059);
or U9426 (N_9426,N_8903,N_8749);
or U9427 (N_9427,N_8319,N_8988);
and U9428 (N_9428,N_8781,N_8523);
nor U9429 (N_9429,N_8310,N_8737);
xnor U9430 (N_9430,N_8938,N_8806);
nand U9431 (N_9431,N_8152,N_8611);
nor U9432 (N_9432,N_8677,N_8357);
nor U9433 (N_9433,N_8179,N_8221);
and U9434 (N_9434,N_8832,N_8673);
nand U9435 (N_9435,N_8843,N_8833);
nand U9436 (N_9436,N_8572,N_8695);
xor U9437 (N_9437,N_8543,N_8888);
and U9438 (N_9438,N_8120,N_8161);
xor U9439 (N_9439,N_8035,N_8592);
or U9440 (N_9440,N_8721,N_8802);
or U9441 (N_9441,N_8527,N_8848);
xnor U9442 (N_9442,N_8976,N_8660);
xor U9443 (N_9443,N_8787,N_8008);
or U9444 (N_9444,N_8834,N_8090);
nor U9445 (N_9445,N_8286,N_8690);
nand U9446 (N_9446,N_8532,N_8280);
nor U9447 (N_9447,N_8048,N_8182);
xor U9448 (N_9448,N_8735,N_8519);
or U9449 (N_9449,N_8436,N_8763);
xnor U9450 (N_9450,N_8857,N_8653);
xor U9451 (N_9451,N_8945,N_8373);
xor U9452 (N_9452,N_8437,N_8312);
xor U9453 (N_9453,N_8244,N_8196);
and U9454 (N_9454,N_8831,N_8827);
or U9455 (N_9455,N_8248,N_8705);
nand U9456 (N_9456,N_8883,N_8996);
xnor U9457 (N_9457,N_8054,N_8706);
or U9458 (N_9458,N_8187,N_8664);
nand U9459 (N_9459,N_8674,N_8740);
xor U9460 (N_9460,N_8300,N_8285);
and U9461 (N_9461,N_8994,N_8027);
nand U9462 (N_9462,N_8045,N_8963);
nor U9463 (N_9463,N_8213,N_8581);
xnor U9464 (N_9464,N_8212,N_8480);
nand U9465 (N_9465,N_8779,N_8494);
and U9466 (N_9466,N_8392,N_8630);
or U9467 (N_9467,N_8149,N_8536);
and U9468 (N_9468,N_8260,N_8382);
and U9469 (N_9469,N_8728,N_8847);
nand U9470 (N_9470,N_8086,N_8099);
nor U9471 (N_9471,N_8037,N_8430);
xnor U9472 (N_9472,N_8222,N_8372);
nand U9473 (N_9473,N_8911,N_8554);
nor U9474 (N_9474,N_8024,N_8097);
and U9475 (N_9475,N_8846,N_8181);
and U9476 (N_9476,N_8953,N_8571);
and U9477 (N_9477,N_8477,N_8071);
or U9478 (N_9478,N_8627,N_8450);
and U9479 (N_9479,N_8358,N_8303);
nand U9480 (N_9480,N_8642,N_8240);
nor U9481 (N_9481,N_8143,N_8064);
or U9482 (N_9482,N_8014,N_8968);
nor U9483 (N_9483,N_8691,N_8738);
and U9484 (N_9484,N_8854,N_8298);
nor U9485 (N_9485,N_8569,N_8655);
and U9486 (N_9486,N_8144,N_8798);
nand U9487 (N_9487,N_8049,N_8971);
and U9488 (N_9488,N_8761,N_8253);
nand U9489 (N_9489,N_8966,N_8517);
or U9490 (N_9490,N_8769,N_8002);
nor U9491 (N_9491,N_8716,N_8025);
xnor U9492 (N_9492,N_8983,N_8475);
and U9493 (N_9493,N_8566,N_8919);
or U9494 (N_9494,N_8305,N_8661);
xor U9495 (N_9495,N_8497,N_8243);
nand U9496 (N_9496,N_8154,N_8865);
or U9497 (N_9497,N_8872,N_8383);
xor U9498 (N_9498,N_8815,N_8279);
and U9499 (N_9499,N_8113,N_8889);
or U9500 (N_9500,N_8479,N_8913);
and U9501 (N_9501,N_8535,N_8954);
nand U9502 (N_9502,N_8998,N_8442);
and U9503 (N_9503,N_8521,N_8187);
or U9504 (N_9504,N_8091,N_8193);
or U9505 (N_9505,N_8229,N_8510);
and U9506 (N_9506,N_8121,N_8226);
nand U9507 (N_9507,N_8055,N_8028);
xnor U9508 (N_9508,N_8734,N_8223);
or U9509 (N_9509,N_8274,N_8949);
nand U9510 (N_9510,N_8439,N_8499);
nand U9511 (N_9511,N_8856,N_8851);
or U9512 (N_9512,N_8088,N_8683);
nor U9513 (N_9513,N_8443,N_8487);
and U9514 (N_9514,N_8911,N_8995);
nor U9515 (N_9515,N_8267,N_8648);
xnor U9516 (N_9516,N_8706,N_8813);
and U9517 (N_9517,N_8907,N_8717);
xnor U9518 (N_9518,N_8825,N_8644);
nand U9519 (N_9519,N_8977,N_8368);
or U9520 (N_9520,N_8828,N_8409);
nand U9521 (N_9521,N_8329,N_8082);
xor U9522 (N_9522,N_8999,N_8311);
nand U9523 (N_9523,N_8460,N_8285);
or U9524 (N_9524,N_8728,N_8668);
xnor U9525 (N_9525,N_8548,N_8581);
nand U9526 (N_9526,N_8637,N_8431);
xor U9527 (N_9527,N_8557,N_8904);
xor U9528 (N_9528,N_8892,N_8775);
xor U9529 (N_9529,N_8539,N_8180);
or U9530 (N_9530,N_8375,N_8134);
xnor U9531 (N_9531,N_8036,N_8086);
nand U9532 (N_9532,N_8435,N_8802);
or U9533 (N_9533,N_8034,N_8448);
nand U9534 (N_9534,N_8966,N_8879);
and U9535 (N_9535,N_8104,N_8349);
nand U9536 (N_9536,N_8776,N_8125);
nor U9537 (N_9537,N_8719,N_8411);
xor U9538 (N_9538,N_8212,N_8979);
nor U9539 (N_9539,N_8807,N_8347);
and U9540 (N_9540,N_8779,N_8859);
nand U9541 (N_9541,N_8565,N_8752);
nor U9542 (N_9542,N_8304,N_8021);
nor U9543 (N_9543,N_8365,N_8339);
and U9544 (N_9544,N_8410,N_8026);
and U9545 (N_9545,N_8417,N_8281);
nand U9546 (N_9546,N_8265,N_8709);
or U9547 (N_9547,N_8535,N_8361);
xor U9548 (N_9548,N_8907,N_8726);
nand U9549 (N_9549,N_8342,N_8820);
xor U9550 (N_9550,N_8089,N_8979);
and U9551 (N_9551,N_8889,N_8713);
nand U9552 (N_9552,N_8336,N_8786);
and U9553 (N_9553,N_8082,N_8736);
and U9554 (N_9554,N_8253,N_8108);
and U9555 (N_9555,N_8435,N_8875);
nand U9556 (N_9556,N_8921,N_8892);
nand U9557 (N_9557,N_8131,N_8228);
and U9558 (N_9558,N_8618,N_8029);
xor U9559 (N_9559,N_8825,N_8944);
and U9560 (N_9560,N_8580,N_8999);
and U9561 (N_9561,N_8934,N_8175);
or U9562 (N_9562,N_8596,N_8988);
nand U9563 (N_9563,N_8027,N_8654);
and U9564 (N_9564,N_8559,N_8272);
and U9565 (N_9565,N_8249,N_8024);
nand U9566 (N_9566,N_8471,N_8152);
and U9567 (N_9567,N_8035,N_8293);
or U9568 (N_9568,N_8195,N_8683);
or U9569 (N_9569,N_8418,N_8155);
and U9570 (N_9570,N_8677,N_8068);
nand U9571 (N_9571,N_8490,N_8449);
nor U9572 (N_9572,N_8197,N_8179);
nor U9573 (N_9573,N_8591,N_8927);
or U9574 (N_9574,N_8739,N_8753);
xnor U9575 (N_9575,N_8873,N_8016);
and U9576 (N_9576,N_8050,N_8579);
and U9577 (N_9577,N_8589,N_8331);
nand U9578 (N_9578,N_8548,N_8461);
and U9579 (N_9579,N_8642,N_8381);
xnor U9580 (N_9580,N_8502,N_8132);
xor U9581 (N_9581,N_8665,N_8626);
and U9582 (N_9582,N_8346,N_8727);
and U9583 (N_9583,N_8789,N_8324);
xnor U9584 (N_9584,N_8200,N_8148);
xor U9585 (N_9585,N_8114,N_8151);
xor U9586 (N_9586,N_8863,N_8251);
nand U9587 (N_9587,N_8091,N_8313);
xor U9588 (N_9588,N_8573,N_8672);
or U9589 (N_9589,N_8271,N_8584);
xor U9590 (N_9590,N_8172,N_8075);
xor U9591 (N_9591,N_8425,N_8899);
nand U9592 (N_9592,N_8525,N_8021);
or U9593 (N_9593,N_8080,N_8217);
nand U9594 (N_9594,N_8623,N_8103);
or U9595 (N_9595,N_8089,N_8601);
nand U9596 (N_9596,N_8949,N_8623);
nor U9597 (N_9597,N_8313,N_8536);
or U9598 (N_9598,N_8294,N_8591);
nor U9599 (N_9599,N_8811,N_8878);
or U9600 (N_9600,N_8743,N_8623);
nand U9601 (N_9601,N_8727,N_8323);
nor U9602 (N_9602,N_8119,N_8371);
xor U9603 (N_9603,N_8309,N_8379);
nor U9604 (N_9604,N_8029,N_8650);
or U9605 (N_9605,N_8204,N_8471);
nor U9606 (N_9606,N_8863,N_8038);
and U9607 (N_9607,N_8546,N_8082);
xor U9608 (N_9608,N_8926,N_8526);
nor U9609 (N_9609,N_8924,N_8150);
and U9610 (N_9610,N_8509,N_8440);
and U9611 (N_9611,N_8917,N_8096);
nor U9612 (N_9612,N_8464,N_8345);
nand U9613 (N_9613,N_8467,N_8865);
and U9614 (N_9614,N_8327,N_8998);
or U9615 (N_9615,N_8145,N_8185);
and U9616 (N_9616,N_8914,N_8870);
nand U9617 (N_9617,N_8919,N_8477);
and U9618 (N_9618,N_8986,N_8807);
xnor U9619 (N_9619,N_8865,N_8687);
nor U9620 (N_9620,N_8716,N_8356);
and U9621 (N_9621,N_8833,N_8109);
nor U9622 (N_9622,N_8604,N_8173);
and U9623 (N_9623,N_8359,N_8659);
xor U9624 (N_9624,N_8672,N_8247);
and U9625 (N_9625,N_8797,N_8766);
nor U9626 (N_9626,N_8609,N_8763);
or U9627 (N_9627,N_8944,N_8566);
xor U9628 (N_9628,N_8671,N_8204);
and U9629 (N_9629,N_8983,N_8267);
xor U9630 (N_9630,N_8679,N_8329);
and U9631 (N_9631,N_8075,N_8334);
and U9632 (N_9632,N_8256,N_8870);
nor U9633 (N_9633,N_8763,N_8351);
nand U9634 (N_9634,N_8444,N_8017);
nand U9635 (N_9635,N_8174,N_8918);
nand U9636 (N_9636,N_8256,N_8684);
nor U9637 (N_9637,N_8736,N_8979);
or U9638 (N_9638,N_8685,N_8722);
or U9639 (N_9639,N_8823,N_8984);
or U9640 (N_9640,N_8855,N_8717);
xnor U9641 (N_9641,N_8978,N_8912);
or U9642 (N_9642,N_8914,N_8826);
nor U9643 (N_9643,N_8739,N_8342);
nand U9644 (N_9644,N_8719,N_8815);
or U9645 (N_9645,N_8824,N_8229);
nand U9646 (N_9646,N_8679,N_8779);
nand U9647 (N_9647,N_8886,N_8049);
and U9648 (N_9648,N_8381,N_8815);
nand U9649 (N_9649,N_8106,N_8405);
or U9650 (N_9650,N_8784,N_8411);
nand U9651 (N_9651,N_8737,N_8972);
and U9652 (N_9652,N_8136,N_8575);
nor U9653 (N_9653,N_8540,N_8784);
nand U9654 (N_9654,N_8295,N_8781);
xor U9655 (N_9655,N_8051,N_8654);
nand U9656 (N_9656,N_8276,N_8815);
nand U9657 (N_9657,N_8527,N_8380);
and U9658 (N_9658,N_8815,N_8798);
nor U9659 (N_9659,N_8619,N_8119);
and U9660 (N_9660,N_8171,N_8353);
nor U9661 (N_9661,N_8349,N_8953);
or U9662 (N_9662,N_8309,N_8876);
xnor U9663 (N_9663,N_8333,N_8399);
xor U9664 (N_9664,N_8414,N_8385);
or U9665 (N_9665,N_8911,N_8446);
or U9666 (N_9666,N_8460,N_8501);
or U9667 (N_9667,N_8862,N_8509);
or U9668 (N_9668,N_8881,N_8176);
and U9669 (N_9669,N_8933,N_8046);
or U9670 (N_9670,N_8255,N_8055);
and U9671 (N_9671,N_8485,N_8393);
nor U9672 (N_9672,N_8586,N_8756);
and U9673 (N_9673,N_8445,N_8203);
xnor U9674 (N_9674,N_8701,N_8004);
or U9675 (N_9675,N_8230,N_8078);
or U9676 (N_9676,N_8135,N_8219);
and U9677 (N_9677,N_8492,N_8312);
xnor U9678 (N_9678,N_8299,N_8685);
or U9679 (N_9679,N_8589,N_8443);
and U9680 (N_9680,N_8233,N_8198);
xor U9681 (N_9681,N_8701,N_8661);
or U9682 (N_9682,N_8508,N_8156);
or U9683 (N_9683,N_8403,N_8277);
nor U9684 (N_9684,N_8665,N_8050);
and U9685 (N_9685,N_8111,N_8644);
nand U9686 (N_9686,N_8781,N_8822);
nor U9687 (N_9687,N_8504,N_8793);
nor U9688 (N_9688,N_8164,N_8524);
or U9689 (N_9689,N_8356,N_8829);
xnor U9690 (N_9690,N_8759,N_8579);
xnor U9691 (N_9691,N_8777,N_8027);
nand U9692 (N_9692,N_8710,N_8514);
and U9693 (N_9693,N_8918,N_8664);
xor U9694 (N_9694,N_8060,N_8189);
or U9695 (N_9695,N_8506,N_8451);
xor U9696 (N_9696,N_8140,N_8257);
nor U9697 (N_9697,N_8713,N_8093);
or U9698 (N_9698,N_8736,N_8328);
nor U9699 (N_9699,N_8461,N_8531);
xor U9700 (N_9700,N_8158,N_8775);
or U9701 (N_9701,N_8290,N_8189);
nor U9702 (N_9702,N_8779,N_8541);
and U9703 (N_9703,N_8797,N_8080);
xor U9704 (N_9704,N_8263,N_8385);
xnor U9705 (N_9705,N_8431,N_8384);
nand U9706 (N_9706,N_8122,N_8029);
nand U9707 (N_9707,N_8927,N_8921);
or U9708 (N_9708,N_8828,N_8097);
nor U9709 (N_9709,N_8028,N_8644);
nand U9710 (N_9710,N_8759,N_8636);
nand U9711 (N_9711,N_8608,N_8082);
nand U9712 (N_9712,N_8938,N_8272);
and U9713 (N_9713,N_8102,N_8259);
or U9714 (N_9714,N_8659,N_8019);
nand U9715 (N_9715,N_8167,N_8267);
nand U9716 (N_9716,N_8291,N_8549);
or U9717 (N_9717,N_8609,N_8696);
nand U9718 (N_9718,N_8532,N_8577);
and U9719 (N_9719,N_8732,N_8848);
and U9720 (N_9720,N_8398,N_8278);
xnor U9721 (N_9721,N_8647,N_8371);
or U9722 (N_9722,N_8863,N_8225);
xor U9723 (N_9723,N_8276,N_8754);
and U9724 (N_9724,N_8236,N_8104);
and U9725 (N_9725,N_8022,N_8451);
nand U9726 (N_9726,N_8100,N_8929);
or U9727 (N_9727,N_8104,N_8826);
nor U9728 (N_9728,N_8408,N_8357);
nor U9729 (N_9729,N_8106,N_8014);
and U9730 (N_9730,N_8974,N_8282);
nor U9731 (N_9731,N_8516,N_8208);
nand U9732 (N_9732,N_8215,N_8208);
and U9733 (N_9733,N_8952,N_8078);
nand U9734 (N_9734,N_8823,N_8977);
and U9735 (N_9735,N_8047,N_8883);
and U9736 (N_9736,N_8184,N_8960);
nand U9737 (N_9737,N_8181,N_8297);
xor U9738 (N_9738,N_8320,N_8255);
or U9739 (N_9739,N_8799,N_8786);
and U9740 (N_9740,N_8061,N_8799);
nor U9741 (N_9741,N_8533,N_8783);
nand U9742 (N_9742,N_8594,N_8795);
nor U9743 (N_9743,N_8617,N_8754);
nor U9744 (N_9744,N_8025,N_8020);
xor U9745 (N_9745,N_8403,N_8989);
nor U9746 (N_9746,N_8510,N_8624);
nand U9747 (N_9747,N_8164,N_8163);
nor U9748 (N_9748,N_8378,N_8018);
and U9749 (N_9749,N_8514,N_8605);
xor U9750 (N_9750,N_8042,N_8187);
nor U9751 (N_9751,N_8747,N_8572);
nor U9752 (N_9752,N_8509,N_8033);
and U9753 (N_9753,N_8989,N_8851);
nand U9754 (N_9754,N_8691,N_8212);
nand U9755 (N_9755,N_8984,N_8376);
nor U9756 (N_9756,N_8703,N_8708);
nand U9757 (N_9757,N_8982,N_8421);
or U9758 (N_9758,N_8314,N_8193);
nand U9759 (N_9759,N_8322,N_8073);
nand U9760 (N_9760,N_8594,N_8668);
xor U9761 (N_9761,N_8665,N_8294);
nand U9762 (N_9762,N_8640,N_8621);
nor U9763 (N_9763,N_8457,N_8978);
xor U9764 (N_9764,N_8083,N_8699);
or U9765 (N_9765,N_8187,N_8145);
nor U9766 (N_9766,N_8128,N_8152);
or U9767 (N_9767,N_8087,N_8662);
or U9768 (N_9768,N_8319,N_8677);
and U9769 (N_9769,N_8386,N_8324);
nand U9770 (N_9770,N_8622,N_8470);
nor U9771 (N_9771,N_8520,N_8926);
or U9772 (N_9772,N_8359,N_8760);
nand U9773 (N_9773,N_8908,N_8322);
nand U9774 (N_9774,N_8186,N_8587);
and U9775 (N_9775,N_8940,N_8957);
xor U9776 (N_9776,N_8484,N_8898);
and U9777 (N_9777,N_8579,N_8112);
and U9778 (N_9778,N_8539,N_8019);
xor U9779 (N_9779,N_8452,N_8108);
and U9780 (N_9780,N_8511,N_8191);
or U9781 (N_9781,N_8115,N_8364);
and U9782 (N_9782,N_8919,N_8785);
nor U9783 (N_9783,N_8391,N_8937);
or U9784 (N_9784,N_8707,N_8585);
nor U9785 (N_9785,N_8045,N_8522);
or U9786 (N_9786,N_8640,N_8906);
or U9787 (N_9787,N_8199,N_8666);
xor U9788 (N_9788,N_8740,N_8956);
or U9789 (N_9789,N_8663,N_8922);
nand U9790 (N_9790,N_8816,N_8403);
xor U9791 (N_9791,N_8025,N_8824);
or U9792 (N_9792,N_8580,N_8707);
nand U9793 (N_9793,N_8238,N_8001);
nor U9794 (N_9794,N_8768,N_8753);
xnor U9795 (N_9795,N_8690,N_8955);
or U9796 (N_9796,N_8092,N_8441);
xnor U9797 (N_9797,N_8850,N_8764);
or U9798 (N_9798,N_8087,N_8458);
nand U9799 (N_9799,N_8398,N_8468);
nor U9800 (N_9800,N_8352,N_8098);
nor U9801 (N_9801,N_8936,N_8210);
nor U9802 (N_9802,N_8850,N_8261);
or U9803 (N_9803,N_8142,N_8121);
and U9804 (N_9804,N_8195,N_8316);
nor U9805 (N_9805,N_8009,N_8308);
or U9806 (N_9806,N_8508,N_8345);
xnor U9807 (N_9807,N_8760,N_8327);
and U9808 (N_9808,N_8467,N_8027);
xnor U9809 (N_9809,N_8910,N_8008);
and U9810 (N_9810,N_8314,N_8888);
nor U9811 (N_9811,N_8001,N_8160);
nor U9812 (N_9812,N_8851,N_8602);
nand U9813 (N_9813,N_8773,N_8552);
xnor U9814 (N_9814,N_8835,N_8296);
nor U9815 (N_9815,N_8910,N_8164);
xor U9816 (N_9816,N_8361,N_8312);
and U9817 (N_9817,N_8701,N_8988);
nand U9818 (N_9818,N_8853,N_8514);
and U9819 (N_9819,N_8117,N_8078);
xnor U9820 (N_9820,N_8760,N_8838);
and U9821 (N_9821,N_8105,N_8683);
nor U9822 (N_9822,N_8294,N_8740);
xor U9823 (N_9823,N_8283,N_8357);
or U9824 (N_9824,N_8532,N_8116);
xor U9825 (N_9825,N_8237,N_8504);
nor U9826 (N_9826,N_8194,N_8910);
xnor U9827 (N_9827,N_8963,N_8635);
xnor U9828 (N_9828,N_8667,N_8816);
and U9829 (N_9829,N_8416,N_8946);
nor U9830 (N_9830,N_8206,N_8961);
or U9831 (N_9831,N_8730,N_8461);
nand U9832 (N_9832,N_8603,N_8984);
nand U9833 (N_9833,N_8470,N_8850);
nand U9834 (N_9834,N_8701,N_8841);
xnor U9835 (N_9835,N_8403,N_8643);
nand U9836 (N_9836,N_8252,N_8178);
and U9837 (N_9837,N_8604,N_8898);
and U9838 (N_9838,N_8852,N_8332);
nor U9839 (N_9839,N_8995,N_8917);
xnor U9840 (N_9840,N_8541,N_8418);
or U9841 (N_9841,N_8106,N_8869);
nor U9842 (N_9842,N_8414,N_8938);
nand U9843 (N_9843,N_8862,N_8501);
nand U9844 (N_9844,N_8511,N_8403);
nand U9845 (N_9845,N_8370,N_8257);
and U9846 (N_9846,N_8469,N_8661);
nand U9847 (N_9847,N_8301,N_8831);
nor U9848 (N_9848,N_8448,N_8696);
or U9849 (N_9849,N_8316,N_8916);
and U9850 (N_9850,N_8614,N_8524);
and U9851 (N_9851,N_8419,N_8317);
and U9852 (N_9852,N_8865,N_8068);
nor U9853 (N_9853,N_8974,N_8859);
nand U9854 (N_9854,N_8539,N_8581);
xnor U9855 (N_9855,N_8340,N_8640);
xor U9856 (N_9856,N_8139,N_8046);
nor U9857 (N_9857,N_8480,N_8750);
nand U9858 (N_9858,N_8755,N_8569);
or U9859 (N_9859,N_8166,N_8575);
and U9860 (N_9860,N_8096,N_8441);
nand U9861 (N_9861,N_8468,N_8805);
or U9862 (N_9862,N_8126,N_8335);
xnor U9863 (N_9863,N_8200,N_8178);
nand U9864 (N_9864,N_8380,N_8602);
and U9865 (N_9865,N_8647,N_8199);
xor U9866 (N_9866,N_8174,N_8171);
nor U9867 (N_9867,N_8594,N_8817);
xor U9868 (N_9868,N_8949,N_8662);
and U9869 (N_9869,N_8627,N_8685);
nor U9870 (N_9870,N_8930,N_8358);
xnor U9871 (N_9871,N_8555,N_8185);
or U9872 (N_9872,N_8959,N_8004);
nand U9873 (N_9873,N_8116,N_8606);
xor U9874 (N_9874,N_8920,N_8746);
xor U9875 (N_9875,N_8288,N_8472);
xor U9876 (N_9876,N_8041,N_8800);
xnor U9877 (N_9877,N_8725,N_8434);
nor U9878 (N_9878,N_8948,N_8597);
xnor U9879 (N_9879,N_8952,N_8313);
or U9880 (N_9880,N_8035,N_8762);
and U9881 (N_9881,N_8922,N_8066);
or U9882 (N_9882,N_8528,N_8857);
xnor U9883 (N_9883,N_8261,N_8319);
xor U9884 (N_9884,N_8404,N_8190);
and U9885 (N_9885,N_8265,N_8245);
xnor U9886 (N_9886,N_8213,N_8192);
nor U9887 (N_9887,N_8490,N_8212);
nand U9888 (N_9888,N_8795,N_8010);
nor U9889 (N_9889,N_8576,N_8577);
or U9890 (N_9890,N_8104,N_8364);
nand U9891 (N_9891,N_8791,N_8503);
and U9892 (N_9892,N_8068,N_8333);
nand U9893 (N_9893,N_8911,N_8222);
and U9894 (N_9894,N_8943,N_8337);
or U9895 (N_9895,N_8896,N_8158);
nand U9896 (N_9896,N_8371,N_8830);
nor U9897 (N_9897,N_8580,N_8454);
nand U9898 (N_9898,N_8782,N_8160);
and U9899 (N_9899,N_8000,N_8922);
nand U9900 (N_9900,N_8623,N_8477);
xor U9901 (N_9901,N_8603,N_8914);
nor U9902 (N_9902,N_8958,N_8476);
or U9903 (N_9903,N_8013,N_8464);
and U9904 (N_9904,N_8155,N_8999);
xnor U9905 (N_9905,N_8785,N_8344);
xor U9906 (N_9906,N_8011,N_8484);
or U9907 (N_9907,N_8253,N_8343);
xor U9908 (N_9908,N_8420,N_8023);
xnor U9909 (N_9909,N_8713,N_8362);
or U9910 (N_9910,N_8180,N_8500);
nor U9911 (N_9911,N_8465,N_8442);
and U9912 (N_9912,N_8434,N_8249);
xor U9913 (N_9913,N_8943,N_8169);
nor U9914 (N_9914,N_8461,N_8194);
xnor U9915 (N_9915,N_8431,N_8340);
or U9916 (N_9916,N_8599,N_8876);
or U9917 (N_9917,N_8653,N_8354);
nand U9918 (N_9918,N_8748,N_8950);
nand U9919 (N_9919,N_8616,N_8222);
or U9920 (N_9920,N_8177,N_8006);
and U9921 (N_9921,N_8101,N_8523);
nor U9922 (N_9922,N_8465,N_8912);
or U9923 (N_9923,N_8834,N_8297);
nand U9924 (N_9924,N_8887,N_8819);
or U9925 (N_9925,N_8611,N_8813);
xor U9926 (N_9926,N_8099,N_8980);
xnor U9927 (N_9927,N_8173,N_8093);
and U9928 (N_9928,N_8409,N_8802);
and U9929 (N_9929,N_8850,N_8122);
nand U9930 (N_9930,N_8059,N_8925);
xnor U9931 (N_9931,N_8980,N_8321);
xnor U9932 (N_9932,N_8534,N_8040);
nor U9933 (N_9933,N_8257,N_8288);
or U9934 (N_9934,N_8484,N_8495);
xnor U9935 (N_9935,N_8063,N_8921);
or U9936 (N_9936,N_8972,N_8483);
and U9937 (N_9937,N_8302,N_8900);
and U9938 (N_9938,N_8023,N_8723);
nand U9939 (N_9939,N_8891,N_8721);
nand U9940 (N_9940,N_8734,N_8427);
and U9941 (N_9941,N_8945,N_8651);
or U9942 (N_9942,N_8301,N_8042);
or U9943 (N_9943,N_8193,N_8599);
xor U9944 (N_9944,N_8585,N_8587);
and U9945 (N_9945,N_8426,N_8637);
or U9946 (N_9946,N_8601,N_8430);
or U9947 (N_9947,N_8514,N_8682);
nand U9948 (N_9948,N_8525,N_8646);
or U9949 (N_9949,N_8200,N_8119);
nand U9950 (N_9950,N_8068,N_8946);
xnor U9951 (N_9951,N_8187,N_8408);
nor U9952 (N_9952,N_8167,N_8883);
and U9953 (N_9953,N_8414,N_8546);
nor U9954 (N_9954,N_8699,N_8795);
xnor U9955 (N_9955,N_8300,N_8468);
xnor U9956 (N_9956,N_8590,N_8834);
or U9957 (N_9957,N_8405,N_8394);
nor U9958 (N_9958,N_8630,N_8617);
or U9959 (N_9959,N_8545,N_8497);
nor U9960 (N_9960,N_8519,N_8095);
or U9961 (N_9961,N_8151,N_8836);
and U9962 (N_9962,N_8464,N_8683);
or U9963 (N_9963,N_8409,N_8595);
xnor U9964 (N_9964,N_8164,N_8185);
nand U9965 (N_9965,N_8493,N_8399);
xor U9966 (N_9966,N_8332,N_8205);
nand U9967 (N_9967,N_8555,N_8360);
or U9968 (N_9968,N_8909,N_8207);
or U9969 (N_9969,N_8043,N_8014);
and U9970 (N_9970,N_8182,N_8239);
or U9971 (N_9971,N_8229,N_8656);
nor U9972 (N_9972,N_8708,N_8175);
nor U9973 (N_9973,N_8852,N_8529);
xor U9974 (N_9974,N_8031,N_8181);
or U9975 (N_9975,N_8288,N_8861);
nand U9976 (N_9976,N_8816,N_8997);
and U9977 (N_9977,N_8913,N_8329);
nand U9978 (N_9978,N_8969,N_8703);
or U9979 (N_9979,N_8178,N_8238);
or U9980 (N_9980,N_8791,N_8454);
or U9981 (N_9981,N_8330,N_8547);
nand U9982 (N_9982,N_8930,N_8897);
and U9983 (N_9983,N_8472,N_8149);
nor U9984 (N_9984,N_8032,N_8016);
xor U9985 (N_9985,N_8185,N_8277);
xnor U9986 (N_9986,N_8946,N_8320);
nand U9987 (N_9987,N_8995,N_8524);
or U9988 (N_9988,N_8051,N_8995);
or U9989 (N_9989,N_8893,N_8426);
or U9990 (N_9990,N_8355,N_8673);
xnor U9991 (N_9991,N_8376,N_8853);
nand U9992 (N_9992,N_8127,N_8210);
nor U9993 (N_9993,N_8097,N_8352);
or U9994 (N_9994,N_8744,N_8525);
or U9995 (N_9995,N_8073,N_8423);
xor U9996 (N_9996,N_8545,N_8715);
nand U9997 (N_9997,N_8501,N_8995);
and U9998 (N_9998,N_8736,N_8708);
xor U9999 (N_9999,N_8398,N_8305);
nand U10000 (N_10000,N_9427,N_9366);
nand U10001 (N_10001,N_9925,N_9566);
nand U10002 (N_10002,N_9569,N_9100);
nand U10003 (N_10003,N_9150,N_9837);
or U10004 (N_10004,N_9022,N_9594);
nand U10005 (N_10005,N_9681,N_9843);
nor U10006 (N_10006,N_9216,N_9805);
nand U10007 (N_10007,N_9748,N_9142);
xnor U10008 (N_10008,N_9167,N_9516);
xnor U10009 (N_10009,N_9103,N_9572);
nor U10010 (N_10010,N_9729,N_9510);
or U10011 (N_10011,N_9912,N_9767);
and U10012 (N_10012,N_9463,N_9246);
and U10013 (N_10013,N_9691,N_9061);
xnor U10014 (N_10014,N_9982,N_9906);
or U10015 (N_10015,N_9847,N_9435);
nor U10016 (N_10016,N_9476,N_9720);
nor U10017 (N_10017,N_9485,N_9746);
nor U10018 (N_10018,N_9221,N_9774);
or U10019 (N_10019,N_9094,N_9825);
nor U10020 (N_10020,N_9359,N_9763);
and U10021 (N_10021,N_9351,N_9632);
or U10022 (N_10022,N_9621,N_9669);
or U10023 (N_10023,N_9564,N_9812);
xnor U10024 (N_10024,N_9090,N_9429);
or U10025 (N_10025,N_9307,N_9153);
and U10026 (N_10026,N_9391,N_9078);
nand U10027 (N_10027,N_9299,N_9283);
and U10028 (N_10028,N_9994,N_9101);
and U10029 (N_10029,N_9890,N_9475);
nor U10030 (N_10030,N_9645,N_9617);
nor U10031 (N_10031,N_9135,N_9260);
nor U10032 (N_10032,N_9279,N_9392);
nand U10033 (N_10033,N_9139,N_9570);
or U10034 (N_10034,N_9779,N_9143);
nand U10035 (N_10035,N_9448,N_9926);
nor U10036 (N_10036,N_9769,N_9481);
xor U10037 (N_10037,N_9866,N_9341);
or U10038 (N_10038,N_9338,N_9327);
nor U10039 (N_10039,N_9236,N_9537);
xnor U10040 (N_10040,N_9313,N_9749);
or U10041 (N_10041,N_9724,N_9854);
or U10042 (N_10042,N_9708,N_9131);
or U10043 (N_10043,N_9842,N_9851);
and U10044 (N_10044,N_9863,N_9444);
and U10045 (N_10045,N_9501,N_9950);
nand U10046 (N_10046,N_9477,N_9253);
nand U10047 (N_10047,N_9212,N_9051);
or U10048 (N_10048,N_9525,N_9317);
nand U10049 (N_10049,N_9794,N_9986);
and U10050 (N_10050,N_9507,N_9534);
nor U10051 (N_10051,N_9331,N_9828);
nand U10052 (N_10052,N_9050,N_9290);
xor U10053 (N_10053,N_9705,N_9978);
or U10054 (N_10054,N_9993,N_9919);
xnor U10055 (N_10055,N_9377,N_9040);
and U10056 (N_10056,N_9249,N_9284);
and U10057 (N_10057,N_9562,N_9019);
or U10058 (N_10058,N_9093,N_9213);
nor U10059 (N_10059,N_9014,N_9007);
nor U10060 (N_10060,N_9321,N_9751);
nor U10061 (N_10061,N_9440,N_9160);
nand U10062 (N_10062,N_9031,N_9242);
nand U10063 (N_10063,N_9294,N_9648);
or U10064 (N_10064,N_9309,N_9742);
nor U10065 (N_10065,N_9489,N_9713);
nand U10066 (N_10066,N_9339,N_9776);
nor U10067 (N_10067,N_9578,N_9659);
and U10068 (N_10068,N_9037,N_9816);
and U10069 (N_10069,N_9164,N_9015);
and U10070 (N_10070,N_9302,N_9677);
or U10071 (N_10071,N_9798,N_9496);
nor U10072 (N_10072,N_9208,N_9232);
nor U10073 (N_10073,N_9428,N_9931);
and U10074 (N_10074,N_9091,N_9670);
or U10075 (N_10075,N_9555,N_9647);
xnor U10076 (N_10076,N_9989,N_9155);
or U10077 (N_10077,N_9055,N_9258);
or U10078 (N_10078,N_9158,N_9154);
nand U10079 (N_10079,N_9373,N_9112);
xor U10080 (N_10080,N_9305,N_9161);
nor U10081 (N_10081,N_9030,N_9217);
or U10082 (N_10082,N_9781,N_9757);
nor U10083 (N_10083,N_9330,N_9703);
xor U10084 (N_10084,N_9021,N_9988);
nand U10085 (N_10085,N_9001,N_9360);
or U10086 (N_10086,N_9857,N_9575);
nor U10087 (N_10087,N_9685,N_9412);
nand U10088 (N_10088,N_9881,N_9588);
or U10089 (N_10089,N_9827,N_9075);
nor U10090 (N_10090,N_9025,N_9416);
xor U10091 (N_10091,N_9162,N_9606);
nand U10092 (N_10092,N_9240,N_9581);
nand U10093 (N_10093,N_9174,N_9577);
or U10094 (N_10094,N_9241,N_9601);
nand U10095 (N_10095,N_9747,N_9409);
and U10096 (N_10096,N_9702,N_9374);
nor U10097 (N_10097,N_9710,N_9082);
nor U10098 (N_10098,N_9792,N_9092);
or U10099 (N_10099,N_9974,N_9786);
and U10100 (N_10100,N_9179,N_9607);
xor U10101 (N_10101,N_9222,N_9590);
xor U10102 (N_10102,N_9332,N_9401);
and U10103 (N_10103,N_9627,N_9121);
nor U10104 (N_10104,N_9626,N_9824);
or U10105 (N_10105,N_9303,N_9459);
nor U10106 (N_10106,N_9680,N_9043);
or U10107 (N_10107,N_9324,N_9419);
xor U10108 (N_10108,N_9257,N_9848);
nor U10109 (N_10109,N_9272,N_9946);
or U10110 (N_10110,N_9576,N_9697);
nand U10111 (N_10111,N_9182,N_9999);
nor U10112 (N_10112,N_9894,N_9755);
and U10113 (N_10113,N_9072,N_9549);
or U10114 (N_10114,N_9329,N_9613);
xor U10115 (N_10115,N_9765,N_9415);
nand U10116 (N_10116,N_9296,N_9773);
and U10117 (N_10117,N_9504,N_9337);
xor U10118 (N_10118,N_9418,N_9565);
nor U10119 (N_10119,N_9883,N_9889);
xor U10120 (N_10120,N_9643,N_9264);
and U10121 (N_10121,N_9888,N_9628);
and U10122 (N_10122,N_9084,N_9582);
nor U10123 (N_10123,N_9281,N_9943);
and U10124 (N_10124,N_9148,N_9984);
nor U10125 (N_10125,N_9243,N_9558);
or U10126 (N_10126,N_9116,N_9903);
and U10127 (N_10127,N_9032,N_9300);
nand U10128 (N_10128,N_9519,N_9069);
and U10129 (N_10129,N_9758,N_9494);
or U10130 (N_10130,N_9508,N_9194);
nor U10131 (N_10131,N_9048,N_9417);
or U10132 (N_10132,N_9325,N_9186);
nand U10133 (N_10133,N_9344,N_9102);
nor U10134 (N_10134,N_9612,N_9815);
nor U10135 (N_10135,N_9630,N_9364);
nor U10136 (N_10136,N_9096,N_9687);
nand U10137 (N_10137,N_9822,N_9977);
and U10138 (N_10138,N_9887,N_9698);
xnor U10139 (N_10139,N_9683,N_9721);
nor U10140 (N_10140,N_9214,N_9944);
or U10141 (N_10141,N_9850,N_9656);
xnor U10142 (N_10142,N_9629,N_9191);
nor U10143 (N_10143,N_9455,N_9599);
or U10144 (N_10144,N_9542,N_9423);
and U10145 (N_10145,N_9457,N_9471);
and U10146 (N_10146,N_9134,N_9190);
nor U10147 (N_10147,N_9342,N_9620);
nor U10148 (N_10148,N_9255,N_9878);
and U10149 (N_10149,N_9618,N_9872);
and U10150 (N_10150,N_9288,N_9602);
xor U10151 (N_10151,N_9853,N_9998);
nand U10152 (N_10152,N_9314,N_9130);
or U10153 (N_10153,N_9492,N_9394);
xnor U10154 (N_10154,N_9512,N_9318);
nand U10155 (N_10155,N_9584,N_9526);
nor U10156 (N_10156,N_9376,N_9247);
nand U10157 (N_10157,N_9270,N_9768);
nand U10158 (N_10158,N_9368,N_9388);
or U10159 (N_10159,N_9750,N_9841);
and U10160 (N_10160,N_9736,N_9591);
xor U10161 (N_10161,N_9737,N_9233);
or U10162 (N_10162,N_9954,N_9046);
or U10163 (N_10163,N_9719,N_9961);
xor U10164 (N_10164,N_9083,N_9262);
nand U10165 (N_10165,N_9775,N_9985);
or U10166 (N_10166,N_9634,N_9336);
and U10167 (N_10167,N_9865,N_9111);
nand U10168 (N_10168,N_9668,N_9559);
nand U10169 (N_10169,N_9560,N_9949);
and U10170 (N_10170,N_9505,N_9334);
and U10171 (N_10171,N_9646,N_9070);
nor U10172 (N_10172,N_9308,N_9744);
nor U10173 (N_10173,N_9261,N_9384);
or U10174 (N_10174,N_9382,N_9044);
or U10175 (N_10175,N_9873,N_9722);
nand U10176 (N_10176,N_9219,N_9975);
nand U10177 (N_10177,N_9802,N_9445);
nand U10178 (N_10178,N_9231,N_9229);
nand U10179 (N_10179,N_9530,N_9458);
nand U10180 (N_10180,N_9468,N_9488);
nand U10181 (N_10181,N_9956,N_9657);
xor U10182 (N_10182,N_9395,N_9641);
and U10183 (N_10183,N_9404,N_9655);
and U10184 (N_10184,N_9035,N_9788);
xnor U10185 (N_10185,N_9945,N_9834);
or U10186 (N_10186,N_9686,N_9005);
or U10187 (N_10187,N_9466,N_9852);
or U10188 (N_10188,N_9473,N_9067);
nand U10189 (N_10189,N_9664,N_9169);
or U10190 (N_10190,N_9108,N_9104);
nand U10191 (N_10191,N_9058,N_9206);
and U10192 (N_10192,N_9004,N_9545);
nand U10193 (N_10193,N_9701,N_9992);
or U10194 (N_10194,N_9995,N_9807);
nor U10195 (N_10195,N_9515,N_9034);
or U10196 (N_10196,N_9728,N_9898);
nor U10197 (N_10197,N_9754,N_9402);
nand U10198 (N_10198,N_9552,N_9411);
xnor U10199 (N_10199,N_9784,N_9692);
nor U10200 (N_10200,N_9859,N_9652);
nand U10201 (N_10201,N_9353,N_9573);
and U10202 (N_10202,N_9413,N_9885);
and U10203 (N_10203,N_9624,N_9616);
nor U10204 (N_10204,N_9731,N_9088);
nor U10205 (N_10205,N_9785,N_9474);
nand U10206 (N_10206,N_9123,N_9183);
or U10207 (N_10207,N_9904,N_9009);
nand U10208 (N_10208,N_9266,N_9438);
nor U10209 (N_10209,N_9587,N_9393);
and U10210 (N_10210,N_9937,N_9804);
or U10211 (N_10211,N_9352,N_9536);
xnor U10212 (N_10212,N_9821,N_9235);
nor U10213 (N_10213,N_9844,N_9598);
and U10214 (N_10214,N_9586,N_9527);
nand U10215 (N_10215,N_9958,N_9389);
and U10216 (N_10216,N_9521,N_9018);
xnor U10217 (N_10217,N_9790,N_9876);
xor U10218 (N_10218,N_9163,N_9835);
xor U10219 (N_10219,N_9579,N_9907);
and U10220 (N_10220,N_9660,N_9712);
or U10221 (N_10221,N_9354,N_9465);
xor U10222 (N_10222,N_9363,N_9684);
nand U10223 (N_10223,N_9913,N_9789);
nand U10224 (N_10224,N_9340,N_9414);
xor U10225 (N_10225,N_9089,N_9400);
or U10226 (N_10226,N_9017,N_9073);
xnor U10227 (N_10227,N_9795,N_9625);
or U10228 (N_10228,N_9178,N_9230);
or U10229 (N_10229,N_9787,N_9033);
nor U10230 (N_10230,N_9449,N_9375);
nor U10231 (N_10231,N_9709,N_9097);
and U10232 (N_10232,N_9727,N_9772);
nor U10233 (N_10233,N_9940,N_9951);
nor U10234 (N_10234,N_9304,N_9105);
or U10235 (N_10235,N_9735,N_9311);
and U10236 (N_10236,N_9140,N_9688);
or U10237 (N_10237,N_9743,N_9874);
nand U10238 (N_10238,N_9398,N_9674);
or U10239 (N_10239,N_9614,N_9276);
or U10240 (N_10240,N_9896,N_9464);
nor U10241 (N_10241,N_9533,N_9238);
nand U10242 (N_10242,N_9611,N_9346);
xnor U10243 (N_10243,N_9063,N_9365);
xor U10244 (N_10244,N_9631,N_9503);
xor U10245 (N_10245,N_9271,N_9862);
or U10246 (N_10246,N_9099,N_9436);
nand U10247 (N_10247,N_9871,N_9280);
and U10248 (N_10248,N_9770,N_9690);
and U10249 (N_10249,N_9642,N_9540);
or U10250 (N_10250,N_9239,N_9506);
xnor U10251 (N_10251,N_9472,N_9372);
and U10252 (N_10252,N_9855,N_9973);
nand U10253 (N_10253,N_9152,N_9277);
xnor U10254 (N_10254,N_9589,N_9820);
nor U10255 (N_10255,N_9204,N_9210);
nor U10256 (N_10256,N_9653,N_9518);
or U10257 (N_10257,N_9864,N_9386);
nor U10258 (N_10258,N_9291,N_9195);
or U10259 (N_10259,N_9910,N_9700);
and U10260 (N_10260,N_9500,N_9615);
or U10261 (N_10261,N_9902,N_9585);
and U10262 (N_10262,N_9446,N_9144);
nand U10263 (N_10263,N_9651,N_9740);
xor U10264 (N_10264,N_9965,N_9369);
nand U10265 (N_10265,N_9726,N_9502);
and U10266 (N_10266,N_9410,N_9900);
or U10267 (N_10267,N_9826,N_9006);
or U10268 (N_10268,N_9432,N_9706);
xnor U10269 (N_10269,N_9491,N_9057);
xnor U10270 (N_10270,N_9600,N_9224);
or U10271 (N_10271,N_9544,N_9071);
nor U10272 (N_10272,N_9267,N_9293);
nand U10273 (N_10273,N_9462,N_9326);
xnor U10274 (N_10274,N_9953,N_9892);
nand U10275 (N_10275,N_9133,N_9456);
and U10276 (N_10276,N_9933,N_9292);
or U10277 (N_10277,N_9833,N_9399);
nand U10278 (N_10278,N_9316,N_9054);
nor U10279 (N_10279,N_9132,N_9707);
xnor U10280 (N_10280,N_9278,N_9170);
and U10281 (N_10281,N_9539,N_9875);
or U10282 (N_10282,N_9066,N_9509);
and U10283 (N_10283,N_9367,N_9936);
nor U10284 (N_10284,N_9780,N_9268);
and U10285 (N_10285,N_9320,N_9443);
and U10286 (N_10286,N_9568,N_9064);
and U10287 (N_10287,N_9942,N_9916);
nand U10288 (N_10288,N_9301,N_9490);
or U10289 (N_10289,N_9927,N_9049);
and U10290 (N_10290,N_9312,N_9322);
xnor U10291 (N_10291,N_9189,N_9228);
and U10292 (N_10292,N_9319,N_9350);
and U10293 (N_10293,N_9197,N_9407);
or U10294 (N_10294,N_9605,N_9172);
or U10295 (N_10295,N_9551,N_9146);
nand U10296 (N_10296,N_9287,N_9486);
or U10297 (N_10297,N_9487,N_9858);
nor U10298 (N_10298,N_9085,N_9196);
and U10299 (N_10299,N_9137,N_9420);
nor U10300 (N_10300,N_9110,N_9849);
and U10301 (N_10301,N_9483,N_9593);
and U10302 (N_10302,N_9193,N_9315);
or U10303 (N_10303,N_9884,N_9451);
nor U10304 (N_10304,N_9730,N_9915);
or U10305 (N_10305,N_9114,N_9295);
nor U10306 (N_10306,N_9733,N_9723);
nand U10307 (N_10307,N_9245,N_9125);
or U10308 (N_10308,N_9187,N_9371);
and U10309 (N_10309,N_9557,N_9310);
and U10310 (N_10310,N_9237,N_9306);
xor U10311 (N_10311,N_9996,N_9076);
xor U10312 (N_10312,N_9433,N_9041);
or U10313 (N_10313,N_9126,N_9715);
or U10314 (N_10314,N_9693,N_9948);
or U10315 (N_10315,N_9151,N_9676);
or U10316 (N_10316,N_9205,N_9405);
xnor U10317 (N_10317,N_9358,N_9886);
nand U10318 (N_10318,N_9548,N_9981);
xnor U10319 (N_10319,N_9782,N_9497);
xnor U10320 (N_10320,N_9603,N_9128);
or U10321 (N_10321,N_9543,N_9059);
or U10322 (N_10322,N_9200,N_9285);
or U10323 (N_10323,N_9002,N_9861);
nand U10324 (N_10324,N_9421,N_9831);
nand U10325 (N_10325,N_9036,N_9809);
and U10326 (N_10326,N_9065,N_9914);
and U10327 (N_10327,N_9406,N_9918);
nor U10328 (N_10328,N_9244,N_9962);
nand U10329 (N_10329,N_9397,N_9797);
nand U10330 (N_10330,N_9638,N_9000);
nor U10331 (N_10331,N_9498,N_9106);
and U10332 (N_10332,N_9595,N_9273);
and U10333 (N_10333,N_9553,N_9425);
xnor U10334 (N_10334,N_9493,N_9003);
nand U10335 (N_10335,N_9696,N_9650);
and U10336 (N_10336,N_9047,N_9666);
xnor U10337 (N_10337,N_9667,N_9345);
nand U10338 (N_10338,N_9813,N_9275);
xor U10339 (N_10339,N_9138,N_9868);
and U10340 (N_10340,N_9609,N_9171);
nand U10341 (N_10341,N_9704,N_9513);
xnor U10342 (N_10342,N_9921,N_9959);
and U10343 (N_10343,N_9026,N_9532);
nor U10344 (N_10344,N_9547,N_9752);
and U10345 (N_10345,N_9426,N_9929);
xor U10346 (N_10346,N_9963,N_9348);
or U10347 (N_10347,N_9830,N_9997);
nand U10348 (N_10348,N_9538,N_9251);
nor U10349 (N_10349,N_9370,N_9678);
or U10350 (N_10350,N_9165,N_9385);
and U10351 (N_10351,N_9524,N_9122);
or U10352 (N_10352,N_9020,N_9523);
and U10353 (N_10353,N_9145,N_9571);
xnor U10354 (N_10354,N_9010,N_9349);
xnor U10355 (N_10355,N_9028,N_9467);
and U10356 (N_10356,N_9934,N_9869);
nand U10357 (N_10357,N_9430,N_9269);
or U10358 (N_10358,N_9362,N_9860);
xor U10359 (N_10359,N_9665,N_9636);
nor U10360 (N_10360,N_9136,N_9381);
nor U10361 (N_10361,N_9450,N_9203);
nor U10362 (N_10362,N_9608,N_9932);
nor U10363 (N_10363,N_9920,N_9739);
xor U10364 (N_10364,N_9604,N_9899);
xnor U10365 (N_10365,N_9218,N_9012);
nor U10366 (N_10366,N_9298,N_9732);
nor U10367 (N_10367,N_9147,N_9226);
or U10368 (N_10368,N_9819,N_9909);
nand U10369 (N_10369,N_9771,N_9441);
nand U10370 (N_10370,N_9528,N_9248);
or U10371 (N_10371,N_9469,N_9972);
nor U10372 (N_10372,N_9380,N_9597);
xnor U10373 (N_10373,N_9199,N_9453);
xor U10374 (N_10374,N_9484,N_9176);
nor U10375 (N_10375,N_9554,N_9791);
xnor U10376 (N_10376,N_9013,N_9546);
nand U10377 (N_10377,N_9928,N_9356);
xor U10378 (N_10378,N_9008,N_9141);
nor U10379 (N_10379,N_9220,N_9762);
nor U10380 (N_10380,N_9157,N_9766);
xor U10381 (N_10381,N_9390,N_9180);
and U10382 (N_10382,N_9938,N_9793);
and U10383 (N_10383,N_9991,N_9511);
nand U10384 (N_10384,N_9107,N_9149);
xnor U10385 (N_10385,N_9838,N_9117);
nor U10386 (N_10386,N_9960,N_9970);
or U10387 (N_10387,N_9202,N_9734);
xor U10388 (N_10388,N_9738,N_9623);
or U10389 (N_10389,N_9810,N_9663);
xor U10390 (N_10390,N_9911,N_9355);
or U10391 (N_10391,N_9673,N_9596);
and U10392 (N_10392,N_9038,N_9198);
and U10393 (N_10393,N_9403,N_9761);
xor U10394 (N_10394,N_9957,N_9556);
nor U10395 (N_10395,N_9181,N_9764);
and U10396 (N_10396,N_9396,N_9286);
nand U10397 (N_10397,N_9478,N_9966);
or U10398 (N_10398,N_9297,N_9045);
xor U10399 (N_10399,N_9649,N_9333);
nand U10400 (N_10400,N_9361,N_9118);
nand U10401 (N_10401,N_9166,N_9357);
and U10402 (N_10402,N_9424,N_9967);
xnor U10403 (N_10403,N_9561,N_9832);
or U10404 (N_10404,N_9905,N_9563);
and U10405 (N_10405,N_9756,N_9759);
or U10406 (N_10406,N_9387,N_9679);
nand U10407 (N_10407,N_9188,N_9482);
or U10408 (N_10408,N_9592,N_9935);
nand U10409 (N_10409,N_9201,N_9461);
nor U10410 (N_10410,N_9753,N_9074);
xor U10411 (N_10411,N_9029,N_9964);
nor U10412 (N_10412,N_9550,N_9947);
nand U10413 (N_10413,N_9745,N_9808);
nand U10414 (N_10414,N_9109,N_9893);
or U10415 (N_10415,N_9159,N_9800);
or U10416 (N_10416,N_9250,N_9454);
xnor U10417 (N_10417,N_9062,N_9610);
nand U10418 (N_10418,N_9803,N_9976);
and U10419 (N_10419,N_9725,N_9077);
xnor U10420 (N_10420,N_9289,N_9823);
nor U10421 (N_10421,N_9801,N_9635);
nand U10422 (N_10422,N_9347,N_9522);
and U10423 (N_10423,N_9840,N_9495);
and U10424 (N_10424,N_9119,N_9567);
nand U10425 (N_10425,N_9856,N_9979);
xnor U10426 (N_10426,N_9806,N_9127);
nand U10427 (N_10427,N_9129,N_9917);
or U10428 (N_10428,N_9952,N_9175);
nand U10429 (N_10429,N_9177,N_9777);
or U10430 (N_10430,N_9675,N_9990);
and U10431 (N_10431,N_9256,N_9225);
or U10432 (N_10432,N_9654,N_9115);
nand U10433 (N_10433,N_9434,N_9839);
or U10434 (N_10434,N_9053,N_9796);
nand U10435 (N_10435,N_9930,N_9227);
nand U10436 (N_10436,N_9081,N_9880);
nand U10437 (N_10437,N_9343,N_9694);
and U10438 (N_10438,N_9924,N_9265);
and U10439 (N_10439,N_9922,N_9867);
xor U10440 (N_10440,N_9955,N_9470);
and U10441 (N_10441,N_9829,N_9968);
or U10442 (N_10442,N_9215,N_9846);
and U10443 (N_10443,N_9439,N_9662);
nand U10444 (N_10444,N_9060,N_9583);
xor U10445 (N_10445,N_9633,N_9207);
xnor U10446 (N_10446,N_9901,N_9223);
xor U10447 (N_10447,N_9682,N_9499);
or U10448 (N_10448,N_9908,N_9328);
nor U10449 (N_10449,N_9541,N_9039);
or U10450 (N_10450,N_9079,N_9323);
or U10451 (N_10451,N_9480,N_9335);
or U10452 (N_10452,N_9923,N_9783);
nor U10453 (N_10453,N_9383,N_9168);
and U10454 (N_10454,N_9052,N_9941);
and U10455 (N_10455,N_9520,N_9185);
xnor U10456 (N_10456,N_9818,N_9259);
and U10457 (N_10457,N_9408,N_9514);
nor U10458 (N_10458,N_9778,N_9879);
nor U10459 (N_10459,N_9184,N_9460);
nor U10460 (N_10460,N_9814,N_9939);
nand U10461 (N_10461,N_9234,N_9192);
and U10462 (N_10462,N_9895,N_9086);
xnor U10463 (N_10463,N_9817,N_9987);
and U10464 (N_10464,N_9983,N_9011);
xnor U10465 (N_10465,N_9442,N_9447);
xnor U10466 (N_10466,N_9845,N_9209);
xor U10467 (N_10467,N_9897,N_9971);
nor U10468 (N_10468,N_9098,N_9811);
nor U10469 (N_10469,N_9027,N_9714);
xor U10470 (N_10470,N_9437,N_9087);
or U10471 (N_10471,N_9580,N_9378);
xor U10472 (N_10472,N_9891,N_9431);
nor U10473 (N_10473,N_9672,N_9760);
xor U10474 (N_10474,N_9080,N_9124);
and U10475 (N_10475,N_9263,N_9619);
or U10476 (N_10476,N_9422,N_9718);
nor U10477 (N_10477,N_9274,N_9252);
and U10478 (N_10478,N_9452,N_9113);
nand U10479 (N_10479,N_9056,N_9024);
or U10480 (N_10480,N_9870,N_9799);
nor U10481 (N_10481,N_9671,N_9622);
nor U10482 (N_10482,N_9877,N_9023);
and U10483 (N_10483,N_9016,N_9741);
xnor U10484 (N_10484,N_9120,N_9574);
or U10485 (N_10485,N_9379,N_9529);
xnor U10486 (N_10486,N_9637,N_9095);
xor U10487 (N_10487,N_9156,N_9068);
and U10488 (N_10488,N_9661,N_9535);
xor U10489 (N_10489,N_9699,N_9479);
xnor U10490 (N_10490,N_9695,N_9717);
nand U10491 (N_10491,N_9689,N_9254);
xnor U10492 (N_10492,N_9658,N_9644);
and U10493 (N_10493,N_9711,N_9531);
xor U10494 (N_10494,N_9042,N_9517);
nand U10495 (N_10495,N_9211,N_9716);
xnor U10496 (N_10496,N_9980,N_9173);
and U10497 (N_10497,N_9282,N_9969);
nor U10498 (N_10498,N_9640,N_9882);
nand U10499 (N_10499,N_9639,N_9836);
or U10500 (N_10500,N_9437,N_9210);
nor U10501 (N_10501,N_9967,N_9279);
nand U10502 (N_10502,N_9629,N_9292);
xnor U10503 (N_10503,N_9618,N_9595);
xnor U10504 (N_10504,N_9725,N_9645);
nor U10505 (N_10505,N_9296,N_9116);
nand U10506 (N_10506,N_9469,N_9204);
nor U10507 (N_10507,N_9722,N_9842);
and U10508 (N_10508,N_9887,N_9054);
xor U10509 (N_10509,N_9178,N_9518);
nor U10510 (N_10510,N_9833,N_9676);
nand U10511 (N_10511,N_9369,N_9776);
nand U10512 (N_10512,N_9469,N_9810);
xnor U10513 (N_10513,N_9042,N_9010);
nor U10514 (N_10514,N_9733,N_9068);
and U10515 (N_10515,N_9485,N_9387);
nor U10516 (N_10516,N_9164,N_9592);
nand U10517 (N_10517,N_9362,N_9759);
or U10518 (N_10518,N_9802,N_9450);
and U10519 (N_10519,N_9059,N_9544);
or U10520 (N_10520,N_9401,N_9972);
or U10521 (N_10521,N_9091,N_9462);
xor U10522 (N_10522,N_9529,N_9023);
and U10523 (N_10523,N_9481,N_9551);
nand U10524 (N_10524,N_9277,N_9930);
nor U10525 (N_10525,N_9770,N_9059);
nand U10526 (N_10526,N_9962,N_9699);
nand U10527 (N_10527,N_9885,N_9515);
xor U10528 (N_10528,N_9255,N_9780);
nor U10529 (N_10529,N_9370,N_9354);
or U10530 (N_10530,N_9440,N_9798);
xor U10531 (N_10531,N_9528,N_9280);
xnor U10532 (N_10532,N_9851,N_9492);
nand U10533 (N_10533,N_9315,N_9391);
xor U10534 (N_10534,N_9662,N_9945);
or U10535 (N_10535,N_9945,N_9890);
nor U10536 (N_10536,N_9928,N_9123);
nor U10537 (N_10537,N_9985,N_9370);
or U10538 (N_10538,N_9558,N_9904);
and U10539 (N_10539,N_9074,N_9692);
or U10540 (N_10540,N_9231,N_9450);
nand U10541 (N_10541,N_9844,N_9971);
or U10542 (N_10542,N_9028,N_9547);
or U10543 (N_10543,N_9249,N_9199);
nand U10544 (N_10544,N_9208,N_9319);
or U10545 (N_10545,N_9033,N_9613);
nor U10546 (N_10546,N_9571,N_9765);
nand U10547 (N_10547,N_9940,N_9838);
and U10548 (N_10548,N_9606,N_9286);
nand U10549 (N_10549,N_9388,N_9831);
nand U10550 (N_10550,N_9198,N_9167);
or U10551 (N_10551,N_9673,N_9896);
or U10552 (N_10552,N_9742,N_9050);
nor U10553 (N_10553,N_9286,N_9938);
nand U10554 (N_10554,N_9136,N_9108);
nand U10555 (N_10555,N_9589,N_9084);
or U10556 (N_10556,N_9025,N_9425);
and U10557 (N_10557,N_9718,N_9902);
and U10558 (N_10558,N_9633,N_9745);
and U10559 (N_10559,N_9534,N_9696);
and U10560 (N_10560,N_9711,N_9774);
nand U10561 (N_10561,N_9622,N_9606);
and U10562 (N_10562,N_9023,N_9590);
and U10563 (N_10563,N_9697,N_9878);
nor U10564 (N_10564,N_9588,N_9735);
xnor U10565 (N_10565,N_9719,N_9138);
or U10566 (N_10566,N_9266,N_9137);
xnor U10567 (N_10567,N_9509,N_9919);
xnor U10568 (N_10568,N_9560,N_9857);
or U10569 (N_10569,N_9575,N_9618);
xnor U10570 (N_10570,N_9997,N_9699);
nor U10571 (N_10571,N_9092,N_9522);
or U10572 (N_10572,N_9750,N_9189);
nor U10573 (N_10573,N_9433,N_9176);
and U10574 (N_10574,N_9109,N_9307);
nor U10575 (N_10575,N_9450,N_9862);
nor U10576 (N_10576,N_9364,N_9320);
and U10577 (N_10577,N_9001,N_9665);
or U10578 (N_10578,N_9876,N_9052);
nor U10579 (N_10579,N_9571,N_9382);
nor U10580 (N_10580,N_9501,N_9422);
nand U10581 (N_10581,N_9743,N_9580);
and U10582 (N_10582,N_9162,N_9190);
or U10583 (N_10583,N_9060,N_9830);
nand U10584 (N_10584,N_9649,N_9287);
nor U10585 (N_10585,N_9836,N_9642);
nor U10586 (N_10586,N_9220,N_9606);
nand U10587 (N_10587,N_9451,N_9530);
nor U10588 (N_10588,N_9061,N_9976);
and U10589 (N_10589,N_9848,N_9850);
xnor U10590 (N_10590,N_9525,N_9529);
and U10591 (N_10591,N_9356,N_9344);
nand U10592 (N_10592,N_9958,N_9914);
nor U10593 (N_10593,N_9997,N_9894);
xnor U10594 (N_10594,N_9145,N_9897);
and U10595 (N_10595,N_9233,N_9640);
nor U10596 (N_10596,N_9871,N_9019);
or U10597 (N_10597,N_9553,N_9680);
nand U10598 (N_10598,N_9040,N_9577);
and U10599 (N_10599,N_9612,N_9270);
nand U10600 (N_10600,N_9166,N_9503);
nand U10601 (N_10601,N_9185,N_9069);
or U10602 (N_10602,N_9824,N_9571);
nor U10603 (N_10603,N_9396,N_9715);
nor U10604 (N_10604,N_9534,N_9361);
nor U10605 (N_10605,N_9403,N_9601);
or U10606 (N_10606,N_9265,N_9552);
or U10607 (N_10607,N_9000,N_9276);
xnor U10608 (N_10608,N_9483,N_9121);
or U10609 (N_10609,N_9423,N_9076);
nand U10610 (N_10610,N_9685,N_9479);
and U10611 (N_10611,N_9267,N_9693);
xnor U10612 (N_10612,N_9502,N_9022);
xnor U10613 (N_10613,N_9558,N_9444);
nand U10614 (N_10614,N_9990,N_9199);
or U10615 (N_10615,N_9981,N_9807);
nor U10616 (N_10616,N_9494,N_9651);
nand U10617 (N_10617,N_9572,N_9193);
or U10618 (N_10618,N_9822,N_9386);
nand U10619 (N_10619,N_9651,N_9571);
nor U10620 (N_10620,N_9462,N_9081);
or U10621 (N_10621,N_9442,N_9771);
nand U10622 (N_10622,N_9093,N_9763);
nand U10623 (N_10623,N_9169,N_9609);
nor U10624 (N_10624,N_9530,N_9876);
or U10625 (N_10625,N_9471,N_9659);
nand U10626 (N_10626,N_9986,N_9180);
nand U10627 (N_10627,N_9247,N_9132);
nor U10628 (N_10628,N_9483,N_9145);
xor U10629 (N_10629,N_9591,N_9244);
nand U10630 (N_10630,N_9370,N_9362);
or U10631 (N_10631,N_9641,N_9746);
nand U10632 (N_10632,N_9509,N_9966);
xor U10633 (N_10633,N_9589,N_9373);
nand U10634 (N_10634,N_9161,N_9629);
xnor U10635 (N_10635,N_9383,N_9011);
and U10636 (N_10636,N_9699,N_9797);
nor U10637 (N_10637,N_9382,N_9436);
or U10638 (N_10638,N_9135,N_9669);
nor U10639 (N_10639,N_9033,N_9109);
nor U10640 (N_10640,N_9296,N_9512);
nand U10641 (N_10641,N_9974,N_9044);
nor U10642 (N_10642,N_9606,N_9577);
and U10643 (N_10643,N_9325,N_9738);
nor U10644 (N_10644,N_9684,N_9552);
or U10645 (N_10645,N_9051,N_9748);
nor U10646 (N_10646,N_9893,N_9726);
xor U10647 (N_10647,N_9945,N_9776);
or U10648 (N_10648,N_9520,N_9721);
and U10649 (N_10649,N_9500,N_9094);
and U10650 (N_10650,N_9825,N_9850);
and U10651 (N_10651,N_9482,N_9948);
nor U10652 (N_10652,N_9210,N_9935);
and U10653 (N_10653,N_9602,N_9033);
nand U10654 (N_10654,N_9437,N_9009);
and U10655 (N_10655,N_9295,N_9970);
nor U10656 (N_10656,N_9651,N_9761);
and U10657 (N_10657,N_9362,N_9413);
and U10658 (N_10658,N_9575,N_9123);
or U10659 (N_10659,N_9936,N_9793);
or U10660 (N_10660,N_9307,N_9569);
nand U10661 (N_10661,N_9016,N_9065);
and U10662 (N_10662,N_9861,N_9771);
nand U10663 (N_10663,N_9269,N_9765);
nand U10664 (N_10664,N_9411,N_9094);
nand U10665 (N_10665,N_9779,N_9613);
nor U10666 (N_10666,N_9064,N_9315);
and U10667 (N_10667,N_9990,N_9341);
or U10668 (N_10668,N_9926,N_9127);
and U10669 (N_10669,N_9617,N_9715);
nor U10670 (N_10670,N_9376,N_9040);
and U10671 (N_10671,N_9572,N_9102);
nand U10672 (N_10672,N_9852,N_9850);
or U10673 (N_10673,N_9871,N_9228);
nand U10674 (N_10674,N_9185,N_9836);
xnor U10675 (N_10675,N_9847,N_9778);
nand U10676 (N_10676,N_9767,N_9529);
or U10677 (N_10677,N_9393,N_9175);
nor U10678 (N_10678,N_9076,N_9438);
xor U10679 (N_10679,N_9067,N_9147);
and U10680 (N_10680,N_9962,N_9929);
or U10681 (N_10681,N_9309,N_9424);
or U10682 (N_10682,N_9882,N_9893);
or U10683 (N_10683,N_9300,N_9061);
nand U10684 (N_10684,N_9037,N_9122);
xnor U10685 (N_10685,N_9150,N_9454);
nand U10686 (N_10686,N_9783,N_9027);
xnor U10687 (N_10687,N_9147,N_9754);
xor U10688 (N_10688,N_9623,N_9395);
and U10689 (N_10689,N_9524,N_9904);
nor U10690 (N_10690,N_9842,N_9122);
xnor U10691 (N_10691,N_9566,N_9755);
xnor U10692 (N_10692,N_9580,N_9162);
and U10693 (N_10693,N_9385,N_9645);
nor U10694 (N_10694,N_9608,N_9499);
nor U10695 (N_10695,N_9569,N_9755);
or U10696 (N_10696,N_9897,N_9260);
xor U10697 (N_10697,N_9831,N_9336);
nand U10698 (N_10698,N_9275,N_9086);
xnor U10699 (N_10699,N_9763,N_9162);
nand U10700 (N_10700,N_9225,N_9030);
nand U10701 (N_10701,N_9237,N_9106);
or U10702 (N_10702,N_9751,N_9689);
or U10703 (N_10703,N_9463,N_9689);
and U10704 (N_10704,N_9193,N_9723);
nand U10705 (N_10705,N_9627,N_9867);
nand U10706 (N_10706,N_9743,N_9488);
or U10707 (N_10707,N_9767,N_9035);
and U10708 (N_10708,N_9527,N_9896);
xnor U10709 (N_10709,N_9476,N_9403);
nand U10710 (N_10710,N_9794,N_9493);
and U10711 (N_10711,N_9361,N_9742);
and U10712 (N_10712,N_9122,N_9092);
nand U10713 (N_10713,N_9889,N_9100);
nand U10714 (N_10714,N_9841,N_9550);
nand U10715 (N_10715,N_9758,N_9673);
or U10716 (N_10716,N_9164,N_9983);
nor U10717 (N_10717,N_9989,N_9247);
or U10718 (N_10718,N_9321,N_9845);
and U10719 (N_10719,N_9758,N_9512);
and U10720 (N_10720,N_9158,N_9902);
and U10721 (N_10721,N_9218,N_9818);
nor U10722 (N_10722,N_9951,N_9052);
nor U10723 (N_10723,N_9602,N_9278);
xor U10724 (N_10724,N_9583,N_9120);
xor U10725 (N_10725,N_9061,N_9672);
and U10726 (N_10726,N_9434,N_9162);
nor U10727 (N_10727,N_9606,N_9278);
and U10728 (N_10728,N_9729,N_9945);
nor U10729 (N_10729,N_9102,N_9394);
xor U10730 (N_10730,N_9580,N_9680);
and U10731 (N_10731,N_9656,N_9300);
or U10732 (N_10732,N_9920,N_9293);
nor U10733 (N_10733,N_9219,N_9823);
or U10734 (N_10734,N_9627,N_9282);
or U10735 (N_10735,N_9051,N_9840);
and U10736 (N_10736,N_9265,N_9221);
and U10737 (N_10737,N_9838,N_9136);
and U10738 (N_10738,N_9608,N_9097);
and U10739 (N_10739,N_9063,N_9759);
xnor U10740 (N_10740,N_9802,N_9373);
nor U10741 (N_10741,N_9151,N_9256);
or U10742 (N_10742,N_9954,N_9933);
nor U10743 (N_10743,N_9158,N_9715);
nor U10744 (N_10744,N_9334,N_9283);
or U10745 (N_10745,N_9787,N_9108);
xnor U10746 (N_10746,N_9989,N_9721);
nand U10747 (N_10747,N_9794,N_9720);
nor U10748 (N_10748,N_9547,N_9669);
nor U10749 (N_10749,N_9246,N_9672);
and U10750 (N_10750,N_9057,N_9710);
or U10751 (N_10751,N_9000,N_9148);
xnor U10752 (N_10752,N_9602,N_9185);
nand U10753 (N_10753,N_9989,N_9428);
xnor U10754 (N_10754,N_9487,N_9218);
or U10755 (N_10755,N_9176,N_9668);
or U10756 (N_10756,N_9335,N_9614);
or U10757 (N_10757,N_9200,N_9532);
and U10758 (N_10758,N_9939,N_9702);
nor U10759 (N_10759,N_9072,N_9202);
or U10760 (N_10760,N_9594,N_9669);
and U10761 (N_10761,N_9401,N_9001);
or U10762 (N_10762,N_9773,N_9159);
nor U10763 (N_10763,N_9875,N_9699);
xnor U10764 (N_10764,N_9231,N_9264);
or U10765 (N_10765,N_9326,N_9762);
xor U10766 (N_10766,N_9153,N_9356);
xnor U10767 (N_10767,N_9783,N_9462);
or U10768 (N_10768,N_9973,N_9995);
nor U10769 (N_10769,N_9287,N_9731);
nor U10770 (N_10770,N_9682,N_9082);
xor U10771 (N_10771,N_9233,N_9501);
xor U10772 (N_10772,N_9613,N_9373);
nor U10773 (N_10773,N_9890,N_9706);
or U10774 (N_10774,N_9217,N_9712);
nor U10775 (N_10775,N_9992,N_9493);
nand U10776 (N_10776,N_9645,N_9544);
xnor U10777 (N_10777,N_9798,N_9006);
xor U10778 (N_10778,N_9379,N_9804);
xor U10779 (N_10779,N_9587,N_9858);
and U10780 (N_10780,N_9812,N_9437);
and U10781 (N_10781,N_9222,N_9657);
xnor U10782 (N_10782,N_9392,N_9469);
and U10783 (N_10783,N_9666,N_9021);
and U10784 (N_10784,N_9863,N_9476);
nor U10785 (N_10785,N_9865,N_9200);
xnor U10786 (N_10786,N_9255,N_9398);
or U10787 (N_10787,N_9738,N_9186);
nand U10788 (N_10788,N_9527,N_9715);
or U10789 (N_10789,N_9131,N_9813);
xnor U10790 (N_10790,N_9045,N_9318);
and U10791 (N_10791,N_9510,N_9606);
and U10792 (N_10792,N_9432,N_9669);
and U10793 (N_10793,N_9345,N_9984);
nand U10794 (N_10794,N_9200,N_9171);
and U10795 (N_10795,N_9127,N_9373);
and U10796 (N_10796,N_9223,N_9367);
nor U10797 (N_10797,N_9011,N_9340);
nor U10798 (N_10798,N_9093,N_9793);
xnor U10799 (N_10799,N_9407,N_9315);
nor U10800 (N_10800,N_9886,N_9527);
xor U10801 (N_10801,N_9462,N_9798);
nand U10802 (N_10802,N_9316,N_9732);
and U10803 (N_10803,N_9487,N_9285);
xor U10804 (N_10804,N_9137,N_9406);
nor U10805 (N_10805,N_9629,N_9231);
xnor U10806 (N_10806,N_9341,N_9343);
and U10807 (N_10807,N_9003,N_9484);
nand U10808 (N_10808,N_9233,N_9154);
or U10809 (N_10809,N_9646,N_9029);
and U10810 (N_10810,N_9146,N_9368);
or U10811 (N_10811,N_9522,N_9457);
nand U10812 (N_10812,N_9196,N_9179);
or U10813 (N_10813,N_9308,N_9615);
nor U10814 (N_10814,N_9829,N_9028);
nand U10815 (N_10815,N_9084,N_9379);
or U10816 (N_10816,N_9243,N_9793);
nand U10817 (N_10817,N_9342,N_9057);
nand U10818 (N_10818,N_9089,N_9755);
or U10819 (N_10819,N_9176,N_9571);
nor U10820 (N_10820,N_9825,N_9341);
xnor U10821 (N_10821,N_9382,N_9047);
and U10822 (N_10822,N_9621,N_9301);
xnor U10823 (N_10823,N_9180,N_9223);
or U10824 (N_10824,N_9610,N_9035);
nand U10825 (N_10825,N_9156,N_9365);
or U10826 (N_10826,N_9184,N_9562);
or U10827 (N_10827,N_9571,N_9950);
and U10828 (N_10828,N_9821,N_9298);
and U10829 (N_10829,N_9204,N_9847);
nand U10830 (N_10830,N_9613,N_9381);
nor U10831 (N_10831,N_9006,N_9805);
or U10832 (N_10832,N_9878,N_9964);
or U10833 (N_10833,N_9527,N_9466);
nor U10834 (N_10834,N_9712,N_9384);
xor U10835 (N_10835,N_9316,N_9281);
nor U10836 (N_10836,N_9786,N_9904);
nor U10837 (N_10837,N_9775,N_9875);
nor U10838 (N_10838,N_9107,N_9402);
nor U10839 (N_10839,N_9254,N_9418);
xor U10840 (N_10840,N_9571,N_9237);
xnor U10841 (N_10841,N_9939,N_9326);
nor U10842 (N_10842,N_9942,N_9085);
or U10843 (N_10843,N_9255,N_9753);
nand U10844 (N_10844,N_9739,N_9499);
nor U10845 (N_10845,N_9551,N_9477);
or U10846 (N_10846,N_9017,N_9957);
or U10847 (N_10847,N_9953,N_9621);
and U10848 (N_10848,N_9517,N_9522);
or U10849 (N_10849,N_9495,N_9992);
and U10850 (N_10850,N_9747,N_9423);
nor U10851 (N_10851,N_9722,N_9648);
or U10852 (N_10852,N_9712,N_9644);
nor U10853 (N_10853,N_9113,N_9909);
xor U10854 (N_10854,N_9050,N_9588);
and U10855 (N_10855,N_9259,N_9230);
and U10856 (N_10856,N_9551,N_9486);
and U10857 (N_10857,N_9974,N_9032);
nor U10858 (N_10858,N_9365,N_9957);
xor U10859 (N_10859,N_9493,N_9152);
and U10860 (N_10860,N_9440,N_9397);
xor U10861 (N_10861,N_9101,N_9106);
xnor U10862 (N_10862,N_9862,N_9419);
and U10863 (N_10863,N_9550,N_9045);
or U10864 (N_10864,N_9036,N_9625);
or U10865 (N_10865,N_9019,N_9532);
xor U10866 (N_10866,N_9880,N_9572);
nand U10867 (N_10867,N_9893,N_9385);
nand U10868 (N_10868,N_9456,N_9931);
nor U10869 (N_10869,N_9191,N_9007);
nor U10870 (N_10870,N_9386,N_9470);
nand U10871 (N_10871,N_9303,N_9214);
nor U10872 (N_10872,N_9682,N_9869);
nor U10873 (N_10873,N_9686,N_9404);
or U10874 (N_10874,N_9140,N_9200);
xnor U10875 (N_10875,N_9470,N_9492);
nand U10876 (N_10876,N_9516,N_9239);
nand U10877 (N_10877,N_9497,N_9469);
or U10878 (N_10878,N_9496,N_9291);
or U10879 (N_10879,N_9270,N_9417);
and U10880 (N_10880,N_9976,N_9899);
and U10881 (N_10881,N_9539,N_9775);
nand U10882 (N_10882,N_9146,N_9773);
or U10883 (N_10883,N_9831,N_9053);
nor U10884 (N_10884,N_9634,N_9753);
xnor U10885 (N_10885,N_9690,N_9140);
and U10886 (N_10886,N_9752,N_9850);
xor U10887 (N_10887,N_9658,N_9939);
and U10888 (N_10888,N_9246,N_9837);
and U10889 (N_10889,N_9541,N_9955);
nor U10890 (N_10890,N_9410,N_9098);
and U10891 (N_10891,N_9021,N_9437);
or U10892 (N_10892,N_9202,N_9778);
xor U10893 (N_10893,N_9912,N_9530);
or U10894 (N_10894,N_9314,N_9422);
xor U10895 (N_10895,N_9256,N_9898);
or U10896 (N_10896,N_9001,N_9307);
or U10897 (N_10897,N_9122,N_9809);
or U10898 (N_10898,N_9424,N_9061);
nand U10899 (N_10899,N_9292,N_9323);
nand U10900 (N_10900,N_9684,N_9540);
nor U10901 (N_10901,N_9236,N_9960);
xnor U10902 (N_10902,N_9272,N_9226);
xnor U10903 (N_10903,N_9416,N_9003);
or U10904 (N_10904,N_9780,N_9676);
nor U10905 (N_10905,N_9988,N_9170);
nand U10906 (N_10906,N_9329,N_9114);
or U10907 (N_10907,N_9650,N_9881);
or U10908 (N_10908,N_9739,N_9200);
and U10909 (N_10909,N_9398,N_9794);
nand U10910 (N_10910,N_9000,N_9162);
xor U10911 (N_10911,N_9683,N_9563);
nand U10912 (N_10912,N_9448,N_9573);
nand U10913 (N_10913,N_9893,N_9051);
xnor U10914 (N_10914,N_9798,N_9377);
and U10915 (N_10915,N_9395,N_9233);
nand U10916 (N_10916,N_9600,N_9452);
nor U10917 (N_10917,N_9048,N_9407);
nand U10918 (N_10918,N_9955,N_9232);
or U10919 (N_10919,N_9590,N_9615);
or U10920 (N_10920,N_9337,N_9649);
nand U10921 (N_10921,N_9833,N_9906);
or U10922 (N_10922,N_9740,N_9535);
nand U10923 (N_10923,N_9470,N_9361);
nor U10924 (N_10924,N_9087,N_9158);
or U10925 (N_10925,N_9644,N_9313);
or U10926 (N_10926,N_9016,N_9095);
nand U10927 (N_10927,N_9925,N_9480);
nand U10928 (N_10928,N_9674,N_9206);
or U10929 (N_10929,N_9454,N_9289);
nor U10930 (N_10930,N_9504,N_9059);
and U10931 (N_10931,N_9738,N_9762);
xor U10932 (N_10932,N_9311,N_9436);
nand U10933 (N_10933,N_9894,N_9686);
or U10934 (N_10934,N_9133,N_9183);
xor U10935 (N_10935,N_9482,N_9200);
or U10936 (N_10936,N_9989,N_9929);
nor U10937 (N_10937,N_9192,N_9591);
and U10938 (N_10938,N_9905,N_9199);
or U10939 (N_10939,N_9525,N_9007);
or U10940 (N_10940,N_9763,N_9229);
nand U10941 (N_10941,N_9692,N_9699);
or U10942 (N_10942,N_9946,N_9333);
nand U10943 (N_10943,N_9895,N_9108);
xnor U10944 (N_10944,N_9549,N_9840);
xnor U10945 (N_10945,N_9473,N_9988);
or U10946 (N_10946,N_9459,N_9818);
nand U10947 (N_10947,N_9181,N_9216);
and U10948 (N_10948,N_9039,N_9490);
nor U10949 (N_10949,N_9110,N_9651);
and U10950 (N_10950,N_9348,N_9617);
and U10951 (N_10951,N_9753,N_9955);
xnor U10952 (N_10952,N_9514,N_9087);
or U10953 (N_10953,N_9330,N_9345);
nand U10954 (N_10954,N_9889,N_9519);
nand U10955 (N_10955,N_9812,N_9296);
xnor U10956 (N_10956,N_9417,N_9915);
and U10957 (N_10957,N_9256,N_9439);
nor U10958 (N_10958,N_9751,N_9040);
and U10959 (N_10959,N_9426,N_9205);
nand U10960 (N_10960,N_9064,N_9434);
nor U10961 (N_10961,N_9676,N_9107);
nor U10962 (N_10962,N_9070,N_9456);
or U10963 (N_10963,N_9000,N_9742);
nor U10964 (N_10964,N_9567,N_9326);
nand U10965 (N_10965,N_9873,N_9227);
and U10966 (N_10966,N_9082,N_9462);
nor U10967 (N_10967,N_9451,N_9447);
nor U10968 (N_10968,N_9066,N_9765);
xor U10969 (N_10969,N_9122,N_9470);
and U10970 (N_10970,N_9131,N_9938);
nor U10971 (N_10971,N_9249,N_9623);
and U10972 (N_10972,N_9747,N_9178);
or U10973 (N_10973,N_9921,N_9120);
xor U10974 (N_10974,N_9994,N_9599);
nand U10975 (N_10975,N_9934,N_9994);
nor U10976 (N_10976,N_9254,N_9049);
and U10977 (N_10977,N_9302,N_9830);
nand U10978 (N_10978,N_9093,N_9670);
nor U10979 (N_10979,N_9848,N_9836);
nand U10980 (N_10980,N_9272,N_9832);
nand U10981 (N_10981,N_9222,N_9172);
or U10982 (N_10982,N_9640,N_9305);
nor U10983 (N_10983,N_9516,N_9780);
or U10984 (N_10984,N_9043,N_9820);
nor U10985 (N_10985,N_9724,N_9508);
nand U10986 (N_10986,N_9014,N_9632);
and U10987 (N_10987,N_9946,N_9380);
xnor U10988 (N_10988,N_9507,N_9080);
or U10989 (N_10989,N_9750,N_9197);
nor U10990 (N_10990,N_9140,N_9047);
or U10991 (N_10991,N_9026,N_9665);
nor U10992 (N_10992,N_9006,N_9952);
or U10993 (N_10993,N_9456,N_9488);
xor U10994 (N_10994,N_9433,N_9338);
and U10995 (N_10995,N_9547,N_9819);
nand U10996 (N_10996,N_9132,N_9945);
xor U10997 (N_10997,N_9738,N_9336);
and U10998 (N_10998,N_9946,N_9687);
nor U10999 (N_10999,N_9648,N_9001);
xnor U11000 (N_11000,N_10611,N_10471);
and U11001 (N_11001,N_10053,N_10932);
nand U11002 (N_11002,N_10113,N_10051);
nand U11003 (N_11003,N_10501,N_10757);
nor U11004 (N_11004,N_10411,N_10015);
nor U11005 (N_11005,N_10499,N_10055);
and U11006 (N_11006,N_10769,N_10068);
or U11007 (N_11007,N_10763,N_10802);
xnor U11008 (N_11008,N_10473,N_10584);
xor U11009 (N_11009,N_10493,N_10884);
xnor U11010 (N_11010,N_10096,N_10014);
or U11011 (N_11011,N_10753,N_10520);
and U11012 (N_11012,N_10309,N_10651);
xnor U11013 (N_11013,N_10925,N_10380);
nor U11014 (N_11014,N_10736,N_10696);
xnor U11015 (N_11015,N_10590,N_10893);
or U11016 (N_11016,N_10995,N_10886);
and U11017 (N_11017,N_10953,N_10999);
nand U11018 (N_11018,N_10549,N_10990);
nor U11019 (N_11019,N_10514,N_10193);
or U11020 (N_11020,N_10556,N_10301);
nand U11021 (N_11021,N_10997,N_10125);
nand U11022 (N_11022,N_10949,N_10324);
xnor U11023 (N_11023,N_10466,N_10412);
or U11024 (N_11024,N_10658,N_10405);
or U11025 (N_11025,N_10421,N_10791);
nand U11026 (N_11026,N_10417,N_10735);
xnor U11027 (N_11027,N_10866,N_10547);
and U11028 (N_11028,N_10021,N_10407);
or U11029 (N_11029,N_10657,N_10740);
and U11030 (N_11030,N_10079,N_10099);
or U11031 (N_11031,N_10858,N_10531);
nor U11032 (N_11032,N_10550,N_10626);
or U11033 (N_11033,N_10379,N_10354);
and U11034 (N_11034,N_10455,N_10574);
nor U11035 (N_11035,N_10027,N_10840);
and U11036 (N_11036,N_10882,N_10320);
nand U11037 (N_11037,N_10679,N_10878);
and U11038 (N_11038,N_10646,N_10891);
xnor U11039 (N_11039,N_10287,N_10154);
nor U11040 (N_11040,N_10152,N_10994);
or U11041 (N_11041,N_10821,N_10451);
nand U11042 (N_11042,N_10219,N_10857);
nand U11043 (N_11043,N_10395,N_10209);
nand U11044 (N_11044,N_10559,N_10159);
or U11045 (N_11045,N_10943,N_10067);
xor U11046 (N_11046,N_10048,N_10138);
xor U11047 (N_11047,N_10686,N_10269);
xnor U11048 (N_11048,N_10930,N_10025);
or U11049 (N_11049,N_10393,N_10042);
nand U11050 (N_11050,N_10355,N_10707);
xnor U11051 (N_11051,N_10117,N_10723);
xnor U11052 (N_11052,N_10522,N_10837);
nor U11053 (N_11053,N_10288,N_10290);
or U11054 (N_11054,N_10634,N_10302);
or U11055 (N_11055,N_10873,N_10533);
nor U11056 (N_11056,N_10947,N_10182);
nand U11057 (N_11057,N_10924,N_10698);
or U11058 (N_11058,N_10765,N_10464);
or U11059 (N_11059,N_10635,N_10912);
nand U11060 (N_11060,N_10390,N_10817);
xor U11061 (N_11061,N_10557,N_10359);
nand U11062 (N_11062,N_10631,N_10221);
or U11063 (N_11063,N_10551,N_10712);
and U11064 (N_11064,N_10612,N_10622);
xor U11065 (N_11065,N_10709,N_10268);
xnor U11066 (N_11066,N_10730,N_10311);
and U11067 (N_11067,N_10582,N_10196);
and U11068 (N_11068,N_10328,N_10486);
nor U11069 (N_11069,N_10992,N_10650);
and U11070 (N_11070,N_10800,N_10123);
xor U11071 (N_11071,N_10711,N_10607);
nor U11072 (N_11072,N_10564,N_10777);
nor U11073 (N_11073,N_10695,N_10868);
nor U11074 (N_11074,N_10491,N_10251);
nand U11075 (N_11075,N_10006,N_10112);
xnor U11076 (N_11076,N_10676,N_10316);
xor U11077 (N_11077,N_10020,N_10392);
xor U11078 (N_11078,N_10373,N_10109);
or U11079 (N_11079,N_10512,N_10326);
nor U11080 (N_11080,N_10605,N_10974);
and U11081 (N_11081,N_10576,N_10385);
or U11082 (N_11082,N_10639,N_10342);
and U11083 (N_11083,N_10865,N_10616);
nor U11084 (N_11084,N_10538,N_10589);
or U11085 (N_11085,N_10917,N_10304);
or U11086 (N_11086,N_10293,N_10744);
nand U11087 (N_11087,N_10186,N_10828);
or U11088 (N_11088,N_10643,N_10835);
xor U11089 (N_11089,N_10376,N_10315);
nor U11090 (N_11090,N_10236,N_10961);
xnor U11091 (N_11091,N_10456,N_10084);
xor U11092 (N_11092,N_10749,N_10495);
or U11093 (N_11093,N_10194,N_10128);
or U11094 (N_11094,N_10286,N_10629);
and U11095 (N_11095,N_10400,N_10191);
nand U11096 (N_11096,N_10850,N_10246);
nand U11097 (N_11097,N_10671,N_10727);
xor U11098 (N_11098,N_10742,N_10497);
nor U11099 (N_11099,N_10216,N_10815);
xnor U11100 (N_11100,N_10841,N_10165);
or U11101 (N_11101,N_10434,N_10477);
and U11102 (N_11102,N_10632,N_10710);
nand U11103 (N_11103,N_10500,N_10608);
nand U11104 (N_11104,N_10463,N_10820);
or U11105 (N_11105,N_10056,N_10579);
and U11106 (N_11106,N_10374,N_10889);
xor U11107 (N_11107,N_10829,N_10085);
xor U11108 (N_11108,N_10010,N_10604);
nor U11109 (N_11109,N_10162,N_10510);
nand U11110 (N_11110,N_10901,N_10274);
or U11111 (N_11111,N_10339,N_10694);
nand U11112 (N_11112,N_10103,N_10419);
and U11113 (N_11113,N_10602,N_10494);
nor U11114 (N_11114,N_10532,N_10936);
xor U11115 (N_11115,N_10016,N_10911);
or U11116 (N_11116,N_10567,N_10244);
xor U11117 (N_11117,N_10278,N_10996);
and U11118 (N_11118,N_10131,N_10641);
or U11119 (N_11119,N_10823,N_10066);
nand U11120 (N_11120,N_10271,N_10610);
and U11121 (N_11121,N_10728,N_10908);
nand U11122 (N_11122,N_10317,N_10964);
nand U11123 (N_11123,N_10472,N_10137);
nand U11124 (N_11124,N_10349,N_10738);
and U11125 (N_11125,N_10931,N_10171);
and U11126 (N_11126,N_10615,N_10807);
nor U11127 (N_11127,N_10313,N_10950);
xor U11128 (N_11128,N_10562,N_10516);
xnor U11129 (N_11129,N_10599,N_10227);
xnor U11130 (N_11130,N_10166,N_10009);
nand U11131 (N_11131,N_10852,N_10235);
xnor U11132 (N_11132,N_10060,N_10369);
or U11133 (N_11133,N_10970,N_10797);
nor U11134 (N_11134,N_10387,N_10179);
nand U11135 (N_11135,N_10654,N_10173);
and U11136 (N_11136,N_10024,N_10687);
xnor U11137 (N_11137,N_10625,N_10031);
xor U11138 (N_11138,N_10050,N_10151);
or U11139 (N_11139,N_10264,N_10764);
nor U11140 (N_11140,N_10693,N_10644);
and U11141 (N_11141,N_10503,N_10366);
nor U11142 (N_11142,N_10289,N_10967);
xnor U11143 (N_11143,N_10778,N_10000);
xor U11144 (N_11144,N_10413,N_10759);
xnor U11145 (N_11145,N_10443,N_10101);
or U11146 (N_11146,N_10169,N_10250);
nor U11147 (N_11147,N_10747,N_10254);
nor U11148 (N_11148,N_10662,N_10902);
and U11149 (N_11149,N_10591,N_10141);
or U11150 (N_11150,N_10799,N_10842);
or U11151 (N_11151,N_10669,N_10459);
nor U11152 (N_11152,N_10665,N_10299);
or U11153 (N_11153,N_10063,N_10170);
xor U11154 (N_11154,N_10448,N_10825);
xor U11155 (N_11155,N_10575,N_10720);
nor U11156 (N_11156,N_10088,N_10052);
and U11157 (N_11157,N_10795,N_10836);
nor U11158 (N_11158,N_10578,N_10869);
nand U11159 (N_11159,N_10982,N_10790);
nor U11160 (N_11160,N_10808,N_10207);
xnor U11161 (N_11161,N_10384,N_10144);
and U11162 (N_11162,N_10715,N_10900);
nor U11163 (N_11163,N_10418,N_10701);
nand U11164 (N_11164,N_10102,N_10150);
or U11165 (N_11165,N_10894,N_10260);
nor U11166 (N_11166,N_10108,N_10259);
or U11167 (N_11167,N_10047,N_10430);
nand U11168 (N_11168,N_10424,N_10176);
nor U11169 (N_11169,N_10167,N_10404);
xor U11170 (N_11170,N_10638,N_10957);
nand U11171 (N_11171,N_10005,N_10240);
nand U11172 (N_11172,N_10896,N_10073);
and U11173 (N_11173,N_10318,N_10548);
and U11174 (N_11174,N_10683,N_10540);
xor U11175 (N_11175,N_10076,N_10517);
nand U11176 (N_11176,N_10043,N_10838);
or U11177 (N_11177,N_10663,N_10297);
nand U11178 (N_11178,N_10595,N_10719);
nor U11179 (N_11179,N_10938,N_10788);
nand U11180 (N_11180,N_10239,N_10205);
and U11181 (N_11181,N_10708,N_10617);
and U11182 (N_11182,N_10426,N_10397);
xor U11183 (N_11183,N_10918,N_10238);
nand U11184 (N_11184,N_10436,N_10175);
nand U11185 (N_11185,N_10987,N_10812);
xnor U11186 (N_11186,N_10204,N_10489);
nand U11187 (N_11187,N_10098,N_10751);
nor U11188 (N_11188,N_10453,N_10139);
and U11189 (N_11189,N_10248,N_10787);
nand U11190 (N_11190,N_10078,N_10656);
nor U11191 (N_11191,N_10202,N_10475);
or U11192 (N_11192,N_10414,N_10245);
nor U11193 (N_11193,N_10529,N_10081);
nor U11194 (N_11194,N_10481,N_10870);
nand U11195 (N_11195,N_10855,N_10779);
or U11196 (N_11196,N_10781,N_10192);
or U11197 (N_11197,N_10523,N_10619);
and U11198 (N_11198,N_10678,N_10070);
nand U11199 (N_11199,N_10653,N_10766);
xor U11200 (N_11200,N_10539,N_10655);
nand U11201 (N_11201,N_10114,N_10846);
nand U11202 (N_11202,N_10899,N_10361);
and U11203 (N_11203,N_10187,N_10926);
or U11204 (N_11204,N_10381,N_10682);
xnor U11205 (N_11205,N_10089,N_10794);
and U11206 (N_11206,N_10774,N_10809);
xnor U11207 (N_11207,N_10630,N_10403);
nand U11208 (N_11208,N_10155,N_10163);
and U11209 (N_11209,N_10482,N_10094);
or U11210 (N_11210,N_10214,N_10046);
and U11211 (N_11211,N_10929,N_10983);
or U11212 (N_11212,N_10168,N_10129);
or U11213 (N_11213,N_10573,N_10319);
nand U11214 (N_11214,N_10793,N_10100);
nand U11215 (N_11215,N_10038,N_10391);
nor U11216 (N_11216,N_10986,N_10824);
xor U11217 (N_11217,N_10325,N_10519);
or U11218 (N_11218,N_10511,N_10199);
or U11219 (N_11219,N_10340,N_10241);
nor U11220 (N_11220,N_10770,N_10441);
nor U11221 (N_11221,N_10365,N_10859);
and U11222 (N_11222,N_10596,N_10093);
or U11223 (N_11223,N_10944,N_10367);
nor U11224 (N_11224,N_10569,N_10518);
and U11225 (N_11225,N_10963,N_10064);
nor U11226 (N_11226,N_10746,N_10554);
xor U11227 (N_11227,N_10724,N_10962);
nand U11228 (N_11228,N_10338,N_10853);
xnor U11229 (N_11229,N_10272,N_10939);
or U11230 (N_11230,N_10704,N_10849);
xnor U11231 (N_11231,N_10661,N_10228);
or U11232 (N_11232,N_10691,N_10305);
nand U11233 (N_11233,N_10335,N_10416);
xor U11234 (N_11234,N_10447,N_10558);
nand U11235 (N_11235,N_10713,N_10498);
nor U11236 (N_11236,N_10904,N_10348);
and U11237 (N_11237,N_10215,N_10314);
and U11238 (N_11238,N_10011,N_10600);
xnor U11239 (N_11239,N_10035,N_10968);
xnor U11240 (N_11240,N_10153,N_10624);
or U11241 (N_11241,N_10524,N_10773);
nand U11242 (N_11242,N_10822,N_10989);
xor U11243 (N_11243,N_10664,N_10796);
and U11244 (N_11244,N_10606,N_10892);
nor U11245 (N_11245,N_10845,N_10537);
nand U11246 (N_11246,N_10504,N_10479);
xor U11247 (N_11247,N_10118,N_10308);
and U11248 (N_11248,N_10382,N_10368);
or U11249 (N_11249,N_10754,N_10910);
nand U11250 (N_11250,N_10592,N_10372);
and U11251 (N_11251,N_10022,N_10871);
xor U11252 (N_11252,N_10371,N_10383);
nor U11253 (N_11253,N_10860,N_10729);
xnor U11254 (N_11254,N_10126,N_10803);
or U11255 (N_11255,N_10277,N_10267);
xnor U11256 (N_11256,N_10408,N_10976);
nor U11257 (N_11257,N_10688,N_10012);
or U11258 (N_11258,N_10030,N_10689);
or U11259 (N_11259,N_10916,N_10143);
and U11260 (N_11260,N_10190,N_10454);
or U11261 (N_11261,N_10065,N_10083);
or U11262 (N_11262,N_10633,N_10530);
and U11263 (N_11263,N_10680,N_10298);
and U11264 (N_11264,N_10146,N_10356);
nand U11265 (N_11265,N_10212,N_10705);
and U11266 (N_11266,N_10174,N_10566);
and U11267 (N_11267,N_10226,N_10568);
xor U11268 (N_11268,N_10922,N_10786);
and U11269 (N_11269,N_10703,N_10394);
or U11270 (N_11270,N_10645,N_10178);
nor U11271 (N_11271,N_10127,N_10438);
xor U11272 (N_11272,N_10462,N_10572);
nor U11273 (N_11273,N_10284,N_10375);
xnor U11274 (N_11274,N_10946,N_10077);
and U11275 (N_11275,N_10898,N_10580);
or U11276 (N_11276,N_10225,N_10352);
and U11277 (N_11277,N_10377,N_10188);
or U11278 (N_11278,N_10667,N_10249);
and U11279 (N_11279,N_10935,N_10649);
or U11280 (N_11280,N_10230,N_10810);
and U11281 (N_11281,N_10675,N_10862);
or U11282 (N_11282,N_10603,N_10734);
xor U11283 (N_11283,N_10013,N_10091);
nand U11284 (N_11284,N_10984,N_10333);
xnor U11285 (N_11285,N_10452,N_10527);
nor U11286 (N_11286,N_10552,N_10200);
nor U11287 (N_11287,N_10061,N_10581);
and U11288 (N_11288,N_10541,N_10714);
xnor U11289 (N_11289,N_10266,N_10149);
nand U11290 (N_11290,N_10023,N_10856);
nor U11291 (N_11291,N_10307,N_10074);
and U11292 (N_11292,N_10208,N_10457);
nor U11293 (N_11293,N_10280,N_10033);
nand U11294 (N_11294,N_10270,N_10353);
xor U11295 (N_11295,N_10909,N_10439);
xnor U11296 (N_11296,N_10410,N_10593);
xnor U11297 (N_11297,N_10161,N_10940);
or U11298 (N_11298,N_10201,N_10621);
nand U11299 (N_11299,N_10095,N_10130);
or U11300 (N_11300,N_10433,N_10934);
xnor U11301 (N_11301,N_10597,N_10652);
and U11302 (N_11302,N_10756,N_10121);
and U11303 (N_11303,N_10402,N_10156);
xnor U11304 (N_11304,N_10180,N_10396);
and U11305 (N_11305,N_10814,N_10036);
and U11306 (N_11306,N_10296,N_10233);
or U11307 (N_11307,N_10933,N_10496);
and U11308 (N_11308,N_10195,N_10758);
nor U11309 (N_11309,N_10872,N_10229);
xor U11310 (N_11310,N_10642,N_10613);
or U11311 (N_11311,N_10087,N_10732);
nor U11312 (N_11312,N_10801,N_10563);
and U11313 (N_11313,N_10183,N_10223);
nor U11314 (N_11314,N_10623,N_10906);
and U11315 (N_11315,N_10848,N_10028);
xor U11316 (N_11316,N_10627,N_10132);
xnor U11317 (N_11317,N_10881,N_10805);
nor U11318 (N_11318,N_10903,N_10185);
or U11319 (N_11319,N_10737,N_10745);
nor U11320 (N_11320,N_10105,N_10423);
nand U11321 (N_11321,N_10609,N_10468);
xnor U11322 (N_11322,N_10389,N_10864);
or U11323 (N_11323,N_10071,N_10851);
xor U11324 (N_11324,N_10344,N_10148);
xnor U11325 (N_11325,N_10692,N_10197);
nand U11326 (N_11326,N_10256,N_10276);
and U11327 (N_11327,N_10378,N_10306);
nand U11328 (N_11328,N_10262,N_10415);
nor U11329 (N_11329,N_10543,N_10003);
xnor U11330 (N_11330,N_10772,N_10386);
nand U11331 (N_11331,N_10040,N_10677);
and U11332 (N_11332,N_10347,N_10637);
and U11333 (N_11333,N_10092,N_10674);
and U11334 (N_11334,N_10560,N_10485);
nand U11335 (N_11335,N_10506,N_10134);
nor U11336 (N_11336,N_10553,N_10037);
nor U11337 (N_11337,N_10952,N_10577);
xor U11338 (N_11338,N_10257,N_10819);
nor U11339 (N_11339,N_10097,N_10670);
xor U11340 (N_11340,N_10292,N_10975);
nor U11341 (N_11341,N_10508,N_10685);
nor U11342 (N_11342,N_10958,N_10941);
nand U11343 (N_11343,N_10830,N_10542);
nor U11344 (N_11344,N_10771,N_10492);
and U11345 (N_11345,N_10798,N_10211);
or U11346 (N_11346,N_10672,N_10666);
and U11347 (N_11347,N_10444,N_10358);
and U11348 (N_11348,N_10755,N_10111);
xnor U11349 (N_11349,N_10782,N_10460);
and U11350 (N_11350,N_10336,N_10806);
nand U11351 (N_11351,N_10534,N_10699);
nand U11352 (N_11352,N_10965,N_10446);
nor U11353 (N_11353,N_10945,N_10488);
nand U11354 (N_11354,N_10034,N_10467);
xnor U11355 (N_11355,N_10640,N_10673);
or U11356 (N_11356,N_10913,N_10258);
nor U11357 (N_11357,N_10887,N_10861);
or U11358 (N_11358,N_10733,N_10750);
nor U11359 (N_11359,N_10157,N_10854);
and U11360 (N_11360,N_10080,N_10721);
xor U11361 (N_11361,N_10090,N_10717);
and U11362 (N_11362,N_10140,N_10279);
nor U11363 (N_11363,N_10263,N_10978);
nand U11364 (N_11364,N_10470,N_10981);
nor U11365 (N_11365,N_10334,N_10401);
xor U11366 (N_11366,N_10461,N_10331);
xnor U11367 (N_11367,N_10697,N_10420);
nand U11368 (N_11368,N_10741,N_10484);
or U11369 (N_11369,N_10690,N_10505);
xnor U11370 (N_11370,N_10045,N_10019);
nor U11371 (N_11371,N_10181,N_10007);
and U11372 (N_11372,N_10370,N_10594);
and U11373 (N_11373,N_10177,N_10437);
xnor U11374 (N_11374,N_10440,N_10136);
and U11375 (N_11375,N_10923,N_10921);
nor U11376 (N_11376,N_10210,N_10160);
xnor U11377 (N_11377,N_10614,N_10458);
nor U11378 (N_11378,N_10907,N_10888);
xor U11379 (N_11379,N_10469,N_10588);
and U11380 (N_11380,N_10867,N_10004);
xor U11381 (N_11381,N_10726,N_10875);
or U11382 (N_11382,N_10785,N_10069);
nor U11383 (N_11383,N_10057,N_10017);
and U11384 (N_11384,N_10222,N_10059);
nor U11385 (N_11385,N_10350,N_10261);
nor U11386 (N_11386,N_10337,N_10224);
nand U11387 (N_11387,N_10847,N_10716);
or U11388 (N_11388,N_10509,N_10811);
nand U11389 (N_11389,N_10535,N_10768);
nand U11390 (N_11390,N_10507,N_10561);
nor U11391 (N_11391,N_10026,N_10874);
nor U11392 (N_11392,N_10748,N_10363);
nor U11393 (N_11393,N_10586,N_10776);
and U11394 (N_11394,N_10832,N_10158);
nor U11395 (N_11395,N_10760,N_10813);
nor U11396 (N_11396,N_10265,N_10502);
xnor U11397 (N_11397,N_10321,N_10839);
nand U11398 (N_11398,N_10145,N_10804);
and U11399 (N_11399,N_10762,N_10971);
or U11400 (N_11400,N_10341,N_10648);
nor U11401 (N_11401,N_10008,N_10956);
xor U11402 (N_11402,N_10189,N_10636);
or U11403 (N_11403,N_10476,N_10243);
or U11404 (N_11404,N_10110,N_10218);
or U11405 (N_11405,N_10291,N_10583);
or U11406 (N_11406,N_10203,N_10834);
and U11407 (N_11407,N_10425,N_10480);
xnor U11408 (N_11408,N_10570,N_10818);
and U11409 (N_11409,N_10104,N_10273);
xor U11410 (N_11410,N_10915,N_10877);
nand U11411 (N_11411,N_10029,N_10998);
and U11412 (N_11412,N_10432,N_10281);
nor U11413 (N_11413,N_10979,N_10660);
nand U11414 (N_11414,N_10345,N_10928);
nand U11415 (N_11415,N_10731,N_10431);
nand U11416 (N_11416,N_10429,N_10133);
xnor U11417 (N_11417,N_10106,N_10330);
and U11418 (N_11418,N_10303,N_10890);
or U11419 (N_11419,N_10525,N_10598);
xnor U11420 (N_11420,N_10844,N_10513);
and U11421 (N_11421,N_10951,N_10357);
or U11422 (N_11422,N_10044,N_10743);
and U11423 (N_11423,N_10075,N_10546);
xnor U11424 (N_11424,N_10885,N_10919);
nand U11425 (N_11425,N_10360,N_10147);
xor U11426 (N_11426,N_10115,N_10285);
and U11427 (N_11427,N_10942,N_10536);
or U11428 (N_11428,N_10565,N_10959);
nand U11429 (N_11429,N_10969,N_10980);
xnor U11430 (N_11430,N_10119,N_10172);
nor U11431 (N_11431,N_10920,N_10427);
and U11432 (N_11432,N_10442,N_10490);
or U11433 (N_11433,N_10295,N_10107);
nor U11434 (N_11434,N_10585,N_10388);
or U11435 (N_11435,N_10237,N_10310);
and U11436 (N_11436,N_10780,N_10973);
and U11437 (N_11437,N_10478,N_10450);
or U11438 (N_11438,N_10445,N_10364);
xor U11439 (N_11439,N_10993,N_10955);
or U11440 (N_11440,N_10752,N_10816);
and U11441 (N_11441,N_10487,N_10300);
nand U11442 (N_11442,N_10876,N_10164);
and U11443 (N_11443,N_10972,N_10954);
nand U11444 (N_11444,N_10406,N_10883);
or U11445 (N_11445,N_10322,N_10895);
and U11446 (N_11446,N_10792,N_10041);
or U11447 (N_11447,N_10398,N_10062);
and U11448 (N_11448,N_10966,N_10252);
and U11449 (N_11449,N_10312,N_10054);
or U11450 (N_11450,N_10618,N_10647);
nand U11451 (N_11451,N_10213,N_10880);
and U11452 (N_11452,N_10700,N_10905);
nor U11453 (N_11453,N_10668,N_10879);
and U11454 (N_11454,N_10275,N_10247);
xnor U11455 (N_11455,N_10659,N_10601);
nand U11456 (N_11456,N_10474,N_10937);
or U11457 (N_11457,N_10283,N_10831);
nand U11458 (N_11458,N_10329,N_10521);
and U11459 (N_11459,N_10988,N_10120);
nand U11460 (N_11460,N_10409,N_10827);
nand U11461 (N_11461,N_10960,N_10833);
or U11462 (N_11462,N_10544,N_10362);
nand U11463 (N_11463,N_10327,N_10927);
and U11464 (N_11464,N_10702,N_10826);
or U11465 (N_11465,N_10232,N_10739);
nor U11466 (N_11466,N_10449,N_10399);
and U11467 (N_11467,N_10039,N_10526);
xnor U11468 (N_11468,N_10789,N_10863);
and U11469 (N_11469,N_10684,N_10914);
nor U11470 (N_11470,N_10242,N_10897);
nor U11471 (N_11471,N_10767,N_10124);
nor U11472 (N_11472,N_10775,N_10072);
nand U11473 (N_11473,N_10032,N_10122);
or U11474 (N_11474,N_10428,N_10948);
nand U11475 (N_11475,N_10231,N_10483);
nor U11476 (N_11476,N_10234,N_10198);
and U11477 (N_11477,N_10783,N_10515);
nor U11478 (N_11478,N_10255,N_10985);
nand U11479 (N_11479,N_10761,N_10784);
xnor U11480 (N_11480,N_10082,N_10346);
nor U11481 (N_11481,N_10545,N_10116);
xor U11482 (N_11482,N_10217,N_10018);
and U11483 (N_11483,N_10465,N_10323);
or U11484 (N_11484,N_10351,N_10843);
xnor U11485 (N_11485,N_10706,N_10002);
and U11486 (N_11486,N_10722,N_10571);
nor U11487 (N_11487,N_10332,N_10620);
xor U11488 (N_11488,N_10142,N_10628);
xnor U11489 (N_11489,N_10587,N_10422);
or U11490 (N_11490,N_10220,N_10718);
and U11491 (N_11491,N_10282,N_10528);
xnor U11492 (N_11492,N_10184,N_10294);
nand U11493 (N_11493,N_10343,N_10725);
or U11494 (N_11494,N_10435,N_10991);
or U11495 (N_11495,N_10135,N_10086);
xnor U11496 (N_11496,N_10058,N_10681);
nor U11497 (N_11497,N_10049,N_10001);
xor U11498 (N_11498,N_10253,N_10206);
nor U11499 (N_11499,N_10977,N_10555);
nor U11500 (N_11500,N_10000,N_10171);
nand U11501 (N_11501,N_10941,N_10872);
xor U11502 (N_11502,N_10080,N_10655);
nand U11503 (N_11503,N_10181,N_10996);
nor U11504 (N_11504,N_10970,N_10994);
nand U11505 (N_11505,N_10909,N_10932);
and U11506 (N_11506,N_10133,N_10889);
xor U11507 (N_11507,N_10962,N_10250);
or U11508 (N_11508,N_10637,N_10804);
or U11509 (N_11509,N_10517,N_10051);
nand U11510 (N_11510,N_10742,N_10289);
or U11511 (N_11511,N_10785,N_10042);
xnor U11512 (N_11512,N_10033,N_10293);
and U11513 (N_11513,N_10354,N_10161);
or U11514 (N_11514,N_10662,N_10198);
nor U11515 (N_11515,N_10548,N_10701);
and U11516 (N_11516,N_10033,N_10950);
xnor U11517 (N_11517,N_10819,N_10157);
xor U11518 (N_11518,N_10996,N_10219);
xnor U11519 (N_11519,N_10957,N_10235);
nand U11520 (N_11520,N_10707,N_10144);
or U11521 (N_11521,N_10202,N_10403);
xnor U11522 (N_11522,N_10036,N_10309);
nand U11523 (N_11523,N_10459,N_10829);
xor U11524 (N_11524,N_10106,N_10746);
or U11525 (N_11525,N_10314,N_10395);
and U11526 (N_11526,N_10887,N_10594);
nor U11527 (N_11527,N_10847,N_10253);
and U11528 (N_11528,N_10337,N_10672);
xor U11529 (N_11529,N_10851,N_10405);
xor U11530 (N_11530,N_10932,N_10166);
nand U11531 (N_11531,N_10301,N_10376);
nor U11532 (N_11532,N_10500,N_10907);
nor U11533 (N_11533,N_10177,N_10529);
or U11534 (N_11534,N_10301,N_10443);
nor U11535 (N_11535,N_10861,N_10169);
nand U11536 (N_11536,N_10920,N_10346);
nand U11537 (N_11537,N_10413,N_10007);
or U11538 (N_11538,N_10265,N_10643);
or U11539 (N_11539,N_10434,N_10847);
nor U11540 (N_11540,N_10240,N_10799);
and U11541 (N_11541,N_10214,N_10422);
nand U11542 (N_11542,N_10341,N_10644);
or U11543 (N_11543,N_10776,N_10577);
nand U11544 (N_11544,N_10207,N_10560);
nand U11545 (N_11545,N_10745,N_10743);
and U11546 (N_11546,N_10954,N_10624);
nor U11547 (N_11547,N_10685,N_10443);
and U11548 (N_11548,N_10731,N_10276);
xor U11549 (N_11549,N_10775,N_10800);
nor U11550 (N_11550,N_10642,N_10878);
nor U11551 (N_11551,N_10740,N_10423);
or U11552 (N_11552,N_10318,N_10944);
and U11553 (N_11553,N_10323,N_10849);
and U11554 (N_11554,N_10467,N_10383);
or U11555 (N_11555,N_10263,N_10644);
nand U11556 (N_11556,N_10842,N_10806);
xnor U11557 (N_11557,N_10545,N_10033);
and U11558 (N_11558,N_10732,N_10505);
or U11559 (N_11559,N_10643,N_10842);
xnor U11560 (N_11560,N_10932,N_10950);
or U11561 (N_11561,N_10147,N_10947);
xnor U11562 (N_11562,N_10060,N_10860);
or U11563 (N_11563,N_10134,N_10621);
xnor U11564 (N_11564,N_10401,N_10942);
or U11565 (N_11565,N_10381,N_10620);
or U11566 (N_11566,N_10043,N_10257);
and U11567 (N_11567,N_10779,N_10620);
and U11568 (N_11568,N_10122,N_10990);
nor U11569 (N_11569,N_10736,N_10904);
nor U11570 (N_11570,N_10046,N_10373);
nand U11571 (N_11571,N_10798,N_10621);
xor U11572 (N_11572,N_10920,N_10937);
nand U11573 (N_11573,N_10065,N_10160);
nor U11574 (N_11574,N_10692,N_10444);
nor U11575 (N_11575,N_10155,N_10445);
nand U11576 (N_11576,N_10234,N_10942);
xnor U11577 (N_11577,N_10912,N_10932);
and U11578 (N_11578,N_10347,N_10942);
or U11579 (N_11579,N_10979,N_10682);
nor U11580 (N_11580,N_10190,N_10642);
or U11581 (N_11581,N_10528,N_10171);
nand U11582 (N_11582,N_10365,N_10297);
nor U11583 (N_11583,N_10331,N_10137);
or U11584 (N_11584,N_10602,N_10884);
or U11585 (N_11585,N_10681,N_10237);
xor U11586 (N_11586,N_10057,N_10704);
and U11587 (N_11587,N_10413,N_10041);
and U11588 (N_11588,N_10517,N_10164);
and U11589 (N_11589,N_10328,N_10647);
nor U11590 (N_11590,N_10723,N_10666);
xor U11591 (N_11591,N_10778,N_10608);
or U11592 (N_11592,N_10764,N_10155);
nand U11593 (N_11593,N_10498,N_10653);
nand U11594 (N_11594,N_10778,N_10472);
and U11595 (N_11595,N_10878,N_10693);
or U11596 (N_11596,N_10434,N_10227);
and U11597 (N_11597,N_10795,N_10092);
xnor U11598 (N_11598,N_10330,N_10098);
xnor U11599 (N_11599,N_10890,N_10467);
nor U11600 (N_11600,N_10079,N_10754);
nor U11601 (N_11601,N_10316,N_10243);
and U11602 (N_11602,N_10248,N_10792);
and U11603 (N_11603,N_10328,N_10067);
nand U11604 (N_11604,N_10829,N_10844);
nand U11605 (N_11605,N_10466,N_10388);
and U11606 (N_11606,N_10819,N_10374);
nor U11607 (N_11607,N_10929,N_10080);
or U11608 (N_11608,N_10329,N_10721);
nor U11609 (N_11609,N_10546,N_10137);
nor U11610 (N_11610,N_10767,N_10774);
or U11611 (N_11611,N_10365,N_10853);
nor U11612 (N_11612,N_10710,N_10384);
or U11613 (N_11613,N_10776,N_10015);
xor U11614 (N_11614,N_10248,N_10784);
nor U11615 (N_11615,N_10614,N_10831);
xnor U11616 (N_11616,N_10218,N_10654);
xnor U11617 (N_11617,N_10611,N_10320);
nand U11618 (N_11618,N_10456,N_10962);
and U11619 (N_11619,N_10325,N_10747);
xor U11620 (N_11620,N_10064,N_10996);
and U11621 (N_11621,N_10626,N_10437);
xor U11622 (N_11622,N_10256,N_10512);
nand U11623 (N_11623,N_10299,N_10040);
nor U11624 (N_11624,N_10865,N_10597);
or U11625 (N_11625,N_10891,N_10281);
and U11626 (N_11626,N_10989,N_10505);
nor U11627 (N_11627,N_10781,N_10519);
nor U11628 (N_11628,N_10080,N_10074);
and U11629 (N_11629,N_10599,N_10010);
nor U11630 (N_11630,N_10141,N_10040);
and U11631 (N_11631,N_10581,N_10746);
and U11632 (N_11632,N_10865,N_10098);
or U11633 (N_11633,N_10103,N_10005);
xnor U11634 (N_11634,N_10341,N_10737);
or U11635 (N_11635,N_10744,N_10542);
nand U11636 (N_11636,N_10729,N_10543);
nor U11637 (N_11637,N_10419,N_10020);
nand U11638 (N_11638,N_10455,N_10164);
nor U11639 (N_11639,N_10490,N_10175);
nand U11640 (N_11640,N_10562,N_10933);
nand U11641 (N_11641,N_10671,N_10376);
or U11642 (N_11642,N_10665,N_10281);
xnor U11643 (N_11643,N_10166,N_10362);
nor U11644 (N_11644,N_10744,N_10099);
and U11645 (N_11645,N_10843,N_10404);
and U11646 (N_11646,N_10821,N_10286);
and U11647 (N_11647,N_10197,N_10726);
xor U11648 (N_11648,N_10932,N_10705);
nand U11649 (N_11649,N_10104,N_10185);
xor U11650 (N_11650,N_10824,N_10948);
xnor U11651 (N_11651,N_10849,N_10031);
nand U11652 (N_11652,N_10266,N_10153);
or U11653 (N_11653,N_10012,N_10800);
nand U11654 (N_11654,N_10372,N_10943);
xor U11655 (N_11655,N_10658,N_10356);
or U11656 (N_11656,N_10682,N_10639);
nand U11657 (N_11657,N_10027,N_10763);
nand U11658 (N_11658,N_10783,N_10496);
or U11659 (N_11659,N_10088,N_10413);
or U11660 (N_11660,N_10332,N_10982);
and U11661 (N_11661,N_10937,N_10153);
nor U11662 (N_11662,N_10163,N_10652);
xor U11663 (N_11663,N_10710,N_10748);
nor U11664 (N_11664,N_10094,N_10292);
and U11665 (N_11665,N_10301,N_10888);
nand U11666 (N_11666,N_10684,N_10635);
nor U11667 (N_11667,N_10016,N_10827);
or U11668 (N_11668,N_10028,N_10231);
or U11669 (N_11669,N_10900,N_10001);
xor U11670 (N_11670,N_10218,N_10422);
nor U11671 (N_11671,N_10230,N_10031);
xor U11672 (N_11672,N_10447,N_10035);
xor U11673 (N_11673,N_10425,N_10671);
or U11674 (N_11674,N_10802,N_10888);
xnor U11675 (N_11675,N_10211,N_10099);
or U11676 (N_11676,N_10105,N_10782);
xnor U11677 (N_11677,N_10602,N_10648);
and U11678 (N_11678,N_10117,N_10300);
xnor U11679 (N_11679,N_10648,N_10368);
and U11680 (N_11680,N_10096,N_10757);
nand U11681 (N_11681,N_10503,N_10400);
and U11682 (N_11682,N_10453,N_10186);
nand U11683 (N_11683,N_10301,N_10760);
or U11684 (N_11684,N_10510,N_10559);
nand U11685 (N_11685,N_10139,N_10758);
nand U11686 (N_11686,N_10575,N_10498);
nor U11687 (N_11687,N_10389,N_10301);
or U11688 (N_11688,N_10394,N_10069);
xnor U11689 (N_11689,N_10733,N_10572);
or U11690 (N_11690,N_10020,N_10412);
nor U11691 (N_11691,N_10803,N_10455);
xnor U11692 (N_11692,N_10367,N_10248);
nor U11693 (N_11693,N_10117,N_10971);
xnor U11694 (N_11694,N_10369,N_10734);
nor U11695 (N_11695,N_10687,N_10515);
nor U11696 (N_11696,N_10277,N_10199);
and U11697 (N_11697,N_10330,N_10420);
nor U11698 (N_11698,N_10924,N_10984);
xor U11699 (N_11699,N_10822,N_10871);
nor U11700 (N_11700,N_10041,N_10886);
nand U11701 (N_11701,N_10027,N_10308);
or U11702 (N_11702,N_10600,N_10621);
nor U11703 (N_11703,N_10534,N_10068);
and U11704 (N_11704,N_10389,N_10793);
nor U11705 (N_11705,N_10260,N_10906);
nor U11706 (N_11706,N_10086,N_10397);
xnor U11707 (N_11707,N_10700,N_10879);
xnor U11708 (N_11708,N_10840,N_10948);
or U11709 (N_11709,N_10255,N_10979);
xor U11710 (N_11710,N_10078,N_10967);
or U11711 (N_11711,N_10224,N_10383);
xnor U11712 (N_11712,N_10313,N_10563);
or U11713 (N_11713,N_10854,N_10046);
and U11714 (N_11714,N_10640,N_10998);
nand U11715 (N_11715,N_10531,N_10526);
or U11716 (N_11716,N_10816,N_10822);
nand U11717 (N_11717,N_10368,N_10874);
nand U11718 (N_11718,N_10620,N_10906);
xor U11719 (N_11719,N_10290,N_10980);
nand U11720 (N_11720,N_10032,N_10330);
and U11721 (N_11721,N_10943,N_10359);
nor U11722 (N_11722,N_10071,N_10565);
and U11723 (N_11723,N_10110,N_10822);
nor U11724 (N_11724,N_10074,N_10222);
or U11725 (N_11725,N_10460,N_10990);
or U11726 (N_11726,N_10674,N_10754);
or U11727 (N_11727,N_10180,N_10082);
or U11728 (N_11728,N_10182,N_10253);
or U11729 (N_11729,N_10733,N_10013);
or U11730 (N_11730,N_10924,N_10632);
xor U11731 (N_11731,N_10851,N_10051);
or U11732 (N_11732,N_10101,N_10239);
and U11733 (N_11733,N_10851,N_10754);
nor U11734 (N_11734,N_10301,N_10540);
and U11735 (N_11735,N_10036,N_10371);
nor U11736 (N_11736,N_10929,N_10622);
nand U11737 (N_11737,N_10408,N_10673);
xnor U11738 (N_11738,N_10757,N_10589);
or U11739 (N_11739,N_10493,N_10539);
or U11740 (N_11740,N_10436,N_10757);
and U11741 (N_11741,N_10462,N_10607);
nor U11742 (N_11742,N_10843,N_10010);
or U11743 (N_11743,N_10989,N_10439);
nand U11744 (N_11744,N_10810,N_10873);
nor U11745 (N_11745,N_10343,N_10607);
or U11746 (N_11746,N_10944,N_10568);
or U11747 (N_11747,N_10766,N_10268);
or U11748 (N_11748,N_10837,N_10491);
nand U11749 (N_11749,N_10158,N_10319);
xnor U11750 (N_11750,N_10293,N_10770);
nand U11751 (N_11751,N_10838,N_10164);
nor U11752 (N_11752,N_10716,N_10706);
nand U11753 (N_11753,N_10941,N_10188);
or U11754 (N_11754,N_10701,N_10187);
xor U11755 (N_11755,N_10767,N_10454);
xor U11756 (N_11756,N_10052,N_10534);
nand U11757 (N_11757,N_10572,N_10018);
nand U11758 (N_11758,N_10775,N_10034);
nand U11759 (N_11759,N_10932,N_10068);
nand U11760 (N_11760,N_10979,N_10483);
nand U11761 (N_11761,N_10754,N_10747);
nor U11762 (N_11762,N_10620,N_10152);
nor U11763 (N_11763,N_10457,N_10046);
nand U11764 (N_11764,N_10908,N_10616);
nor U11765 (N_11765,N_10815,N_10989);
nand U11766 (N_11766,N_10443,N_10084);
or U11767 (N_11767,N_10838,N_10792);
nand U11768 (N_11768,N_10594,N_10234);
nand U11769 (N_11769,N_10768,N_10302);
and U11770 (N_11770,N_10361,N_10860);
nand U11771 (N_11771,N_10295,N_10627);
nand U11772 (N_11772,N_10656,N_10320);
and U11773 (N_11773,N_10728,N_10442);
or U11774 (N_11774,N_10613,N_10801);
nor U11775 (N_11775,N_10296,N_10214);
nor U11776 (N_11776,N_10857,N_10650);
xnor U11777 (N_11777,N_10882,N_10807);
xnor U11778 (N_11778,N_10182,N_10922);
nor U11779 (N_11779,N_10427,N_10968);
xor U11780 (N_11780,N_10191,N_10089);
nand U11781 (N_11781,N_10568,N_10803);
or U11782 (N_11782,N_10014,N_10094);
nor U11783 (N_11783,N_10143,N_10202);
and U11784 (N_11784,N_10822,N_10955);
nor U11785 (N_11785,N_10454,N_10369);
or U11786 (N_11786,N_10545,N_10010);
nor U11787 (N_11787,N_10521,N_10496);
and U11788 (N_11788,N_10093,N_10328);
and U11789 (N_11789,N_10660,N_10802);
nand U11790 (N_11790,N_10164,N_10965);
or U11791 (N_11791,N_10954,N_10343);
and U11792 (N_11792,N_10749,N_10979);
nand U11793 (N_11793,N_10210,N_10841);
and U11794 (N_11794,N_10711,N_10606);
and U11795 (N_11795,N_10017,N_10984);
nand U11796 (N_11796,N_10847,N_10235);
and U11797 (N_11797,N_10919,N_10250);
or U11798 (N_11798,N_10567,N_10593);
nor U11799 (N_11799,N_10237,N_10048);
nand U11800 (N_11800,N_10052,N_10047);
nand U11801 (N_11801,N_10315,N_10682);
nor U11802 (N_11802,N_10303,N_10595);
nor U11803 (N_11803,N_10133,N_10241);
xnor U11804 (N_11804,N_10847,N_10910);
nor U11805 (N_11805,N_10161,N_10201);
xor U11806 (N_11806,N_10480,N_10511);
xnor U11807 (N_11807,N_10330,N_10052);
and U11808 (N_11808,N_10745,N_10598);
and U11809 (N_11809,N_10494,N_10123);
nand U11810 (N_11810,N_10607,N_10817);
nand U11811 (N_11811,N_10506,N_10612);
nor U11812 (N_11812,N_10026,N_10660);
or U11813 (N_11813,N_10791,N_10095);
nor U11814 (N_11814,N_10995,N_10616);
or U11815 (N_11815,N_10967,N_10465);
and U11816 (N_11816,N_10541,N_10788);
nor U11817 (N_11817,N_10924,N_10977);
or U11818 (N_11818,N_10638,N_10694);
nand U11819 (N_11819,N_10500,N_10731);
or U11820 (N_11820,N_10996,N_10345);
or U11821 (N_11821,N_10998,N_10379);
xnor U11822 (N_11822,N_10254,N_10075);
or U11823 (N_11823,N_10414,N_10420);
nand U11824 (N_11824,N_10157,N_10463);
or U11825 (N_11825,N_10906,N_10341);
and U11826 (N_11826,N_10401,N_10824);
nor U11827 (N_11827,N_10597,N_10472);
nand U11828 (N_11828,N_10179,N_10691);
xor U11829 (N_11829,N_10520,N_10336);
or U11830 (N_11830,N_10439,N_10347);
or U11831 (N_11831,N_10817,N_10515);
nand U11832 (N_11832,N_10260,N_10577);
xor U11833 (N_11833,N_10248,N_10461);
or U11834 (N_11834,N_10491,N_10237);
nor U11835 (N_11835,N_10741,N_10546);
xor U11836 (N_11836,N_10520,N_10455);
or U11837 (N_11837,N_10364,N_10682);
and U11838 (N_11838,N_10041,N_10177);
nand U11839 (N_11839,N_10358,N_10072);
nor U11840 (N_11840,N_10193,N_10541);
and U11841 (N_11841,N_10146,N_10814);
nand U11842 (N_11842,N_10252,N_10580);
xor U11843 (N_11843,N_10926,N_10353);
nor U11844 (N_11844,N_10384,N_10309);
or U11845 (N_11845,N_10114,N_10723);
nand U11846 (N_11846,N_10080,N_10554);
xnor U11847 (N_11847,N_10972,N_10987);
or U11848 (N_11848,N_10914,N_10786);
xnor U11849 (N_11849,N_10660,N_10735);
or U11850 (N_11850,N_10514,N_10871);
nand U11851 (N_11851,N_10709,N_10282);
and U11852 (N_11852,N_10127,N_10463);
or U11853 (N_11853,N_10147,N_10648);
nor U11854 (N_11854,N_10459,N_10070);
and U11855 (N_11855,N_10732,N_10562);
xor U11856 (N_11856,N_10795,N_10477);
xor U11857 (N_11857,N_10574,N_10995);
xor U11858 (N_11858,N_10370,N_10076);
xnor U11859 (N_11859,N_10094,N_10709);
nand U11860 (N_11860,N_10237,N_10046);
and U11861 (N_11861,N_10789,N_10801);
nand U11862 (N_11862,N_10524,N_10047);
or U11863 (N_11863,N_10750,N_10374);
or U11864 (N_11864,N_10189,N_10286);
or U11865 (N_11865,N_10135,N_10440);
and U11866 (N_11866,N_10423,N_10600);
and U11867 (N_11867,N_10656,N_10694);
or U11868 (N_11868,N_10938,N_10994);
nor U11869 (N_11869,N_10527,N_10341);
xor U11870 (N_11870,N_10118,N_10480);
nor U11871 (N_11871,N_10108,N_10326);
xnor U11872 (N_11872,N_10146,N_10552);
xnor U11873 (N_11873,N_10860,N_10886);
or U11874 (N_11874,N_10816,N_10936);
nand U11875 (N_11875,N_10858,N_10093);
or U11876 (N_11876,N_10783,N_10047);
and U11877 (N_11877,N_10523,N_10650);
nor U11878 (N_11878,N_10595,N_10030);
xnor U11879 (N_11879,N_10489,N_10589);
or U11880 (N_11880,N_10324,N_10025);
nand U11881 (N_11881,N_10524,N_10940);
nand U11882 (N_11882,N_10775,N_10156);
xnor U11883 (N_11883,N_10493,N_10192);
xnor U11884 (N_11884,N_10714,N_10157);
nand U11885 (N_11885,N_10538,N_10239);
nand U11886 (N_11886,N_10926,N_10744);
or U11887 (N_11887,N_10808,N_10120);
nor U11888 (N_11888,N_10055,N_10698);
nand U11889 (N_11889,N_10534,N_10545);
nor U11890 (N_11890,N_10445,N_10258);
or U11891 (N_11891,N_10770,N_10323);
and U11892 (N_11892,N_10182,N_10249);
and U11893 (N_11893,N_10862,N_10272);
nor U11894 (N_11894,N_10127,N_10412);
xor U11895 (N_11895,N_10315,N_10599);
xor U11896 (N_11896,N_10130,N_10748);
nand U11897 (N_11897,N_10934,N_10364);
nand U11898 (N_11898,N_10109,N_10279);
nor U11899 (N_11899,N_10029,N_10316);
and U11900 (N_11900,N_10155,N_10387);
or U11901 (N_11901,N_10544,N_10440);
or U11902 (N_11902,N_10314,N_10083);
nor U11903 (N_11903,N_10021,N_10192);
nand U11904 (N_11904,N_10984,N_10062);
xnor U11905 (N_11905,N_10545,N_10144);
nand U11906 (N_11906,N_10195,N_10077);
nand U11907 (N_11907,N_10875,N_10145);
and U11908 (N_11908,N_10040,N_10322);
nand U11909 (N_11909,N_10516,N_10323);
and U11910 (N_11910,N_10782,N_10547);
nor U11911 (N_11911,N_10207,N_10781);
nand U11912 (N_11912,N_10381,N_10439);
and U11913 (N_11913,N_10063,N_10082);
and U11914 (N_11914,N_10265,N_10865);
xor U11915 (N_11915,N_10882,N_10883);
or U11916 (N_11916,N_10621,N_10683);
and U11917 (N_11917,N_10786,N_10829);
xor U11918 (N_11918,N_10661,N_10713);
nand U11919 (N_11919,N_10792,N_10545);
nand U11920 (N_11920,N_10522,N_10512);
xor U11921 (N_11921,N_10756,N_10187);
or U11922 (N_11922,N_10229,N_10121);
and U11923 (N_11923,N_10963,N_10300);
nand U11924 (N_11924,N_10877,N_10264);
and U11925 (N_11925,N_10771,N_10395);
and U11926 (N_11926,N_10720,N_10846);
and U11927 (N_11927,N_10479,N_10186);
or U11928 (N_11928,N_10723,N_10378);
nand U11929 (N_11929,N_10610,N_10183);
nor U11930 (N_11930,N_10077,N_10231);
xnor U11931 (N_11931,N_10175,N_10400);
xor U11932 (N_11932,N_10529,N_10524);
and U11933 (N_11933,N_10420,N_10009);
nand U11934 (N_11934,N_10363,N_10770);
and U11935 (N_11935,N_10306,N_10581);
nand U11936 (N_11936,N_10790,N_10656);
xor U11937 (N_11937,N_10810,N_10491);
or U11938 (N_11938,N_10056,N_10763);
nand U11939 (N_11939,N_10066,N_10520);
xnor U11940 (N_11940,N_10552,N_10444);
or U11941 (N_11941,N_10532,N_10129);
nand U11942 (N_11942,N_10871,N_10914);
nor U11943 (N_11943,N_10070,N_10457);
nor U11944 (N_11944,N_10882,N_10571);
or U11945 (N_11945,N_10897,N_10703);
and U11946 (N_11946,N_10264,N_10878);
or U11947 (N_11947,N_10223,N_10369);
nor U11948 (N_11948,N_10203,N_10292);
xnor U11949 (N_11949,N_10852,N_10658);
or U11950 (N_11950,N_10866,N_10404);
nand U11951 (N_11951,N_10328,N_10701);
xnor U11952 (N_11952,N_10536,N_10263);
nor U11953 (N_11953,N_10204,N_10774);
and U11954 (N_11954,N_10188,N_10982);
or U11955 (N_11955,N_10999,N_10771);
nor U11956 (N_11956,N_10286,N_10248);
xnor U11957 (N_11957,N_10746,N_10836);
xnor U11958 (N_11958,N_10105,N_10864);
nor U11959 (N_11959,N_10167,N_10348);
nand U11960 (N_11960,N_10039,N_10020);
nor U11961 (N_11961,N_10754,N_10959);
nand U11962 (N_11962,N_10911,N_10917);
or U11963 (N_11963,N_10216,N_10692);
xor U11964 (N_11964,N_10049,N_10361);
or U11965 (N_11965,N_10156,N_10001);
and U11966 (N_11966,N_10644,N_10505);
and U11967 (N_11967,N_10112,N_10599);
nand U11968 (N_11968,N_10607,N_10131);
or U11969 (N_11969,N_10925,N_10564);
xnor U11970 (N_11970,N_10496,N_10892);
nor U11971 (N_11971,N_10435,N_10731);
nor U11972 (N_11972,N_10438,N_10469);
nand U11973 (N_11973,N_10632,N_10276);
or U11974 (N_11974,N_10430,N_10156);
xor U11975 (N_11975,N_10602,N_10262);
nor U11976 (N_11976,N_10798,N_10311);
nand U11977 (N_11977,N_10871,N_10651);
nand U11978 (N_11978,N_10360,N_10001);
nand U11979 (N_11979,N_10664,N_10184);
nand U11980 (N_11980,N_10121,N_10778);
nand U11981 (N_11981,N_10142,N_10848);
nor U11982 (N_11982,N_10821,N_10237);
xor U11983 (N_11983,N_10037,N_10065);
nand U11984 (N_11984,N_10534,N_10523);
and U11985 (N_11985,N_10475,N_10866);
nor U11986 (N_11986,N_10554,N_10188);
xor U11987 (N_11987,N_10206,N_10127);
and U11988 (N_11988,N_10901,N_10044);
nand U11989 (N_11989,N_10909,N_10187);
and U11990 (N_11990,N_10684,N_10158);
nor U11991 (N_11991,N_10341,N_10587);
or U11992 (N_11992,N_10849,N_10567);
nor U11993 (N_11993,N_10618,N_10034);
xor U11994 (N_11994,N_10973,N_10490);
xnor U11995 (N_11995,N_10722,N_10851);
xnor U11996 (N_11996,N_10707,N_10923);
nor U11997 (N_11997,N_10859,N_10746);
nor U11998 (N_11998,N_10107,N_10346);
or U11999 (N_11999,N_10314,N_10364);
and U12000 (N_12000,N_11944,N_11035);
or U12001 (N_12001,N_11263,N_11248);
and U12002 (N_12002,N_11283,N_11197);
and U12003 (N_12003,N_11294,N_11576);
and U12004 (N_12004,N_11304,N_11847);
xor U12005 (N_12005,N_11861,N_11746);
or U12006 (N_12006,N_11175,N_11392);
nand U12007 (N_12007,N_11716,N_11968);
and U12008 (N_12008,N_11395,N_11137);
xor U12009 (N_12009,N_11505,N_11676);
nor U12010 (N_12010,N_11829,N_11951);
nor U12011 (N_12011,N_11367,N_11754);
nor U12012 (N_12012,N_11914,N_11209);
nand U12013 (N_12013,N_11350,N_11489);
xor U12014 (N_12014,N_11625,N_11622);
or U12015 (N_12015,N_11040,N_11110);
or U12016 (N_12016,N_11067,N_11539);
or U12017 (N_12017,N_11899,N_11860);
nor U12018 (N_12018,N_11938,N_11745);
nand U12019 (N_12019,N_11901,N_11726);
nor U12020 (N_12020,N_11271,N_11379);
or U12021 (N_12021,N_11663,N_11877);
nor U12022 (N_12022,N_11984,N_11297);
and U12023 (N_12023,N_11493,N_11713);
or U12024 (N_12024,N_11051,N_11991);
and U12025 (N_12025,N_11955,N_11074);
and U12026 (N_12026,N_11657,N_11133);
and U12027 (N_12027,N_11315,N_11347);
nor U12028 (N_12028,N_11520,N_11690);
nand U12029 (N_12029,N_11403,N_11206);
nand U12030 (N_12030,N_11875,N_11849);
nor U12031 (N_12031,N_11118,N_11391);
xnor U12032 (N_12032,N_11130,N_11019);
nand U12033 (N_12033,N_11141,N_11753);
xnor U12034 (N_12034,N_11302,N_11522);
and U12035 (N_12035,N_11354,N_11099);
nand U12036 (N_12036,N_11364,N_11455);
nand U12037 (N_12037,N_11805,N_11958);
xor U12038 (N_12038,N_11487,N_11219);
and U12039 (N_12039,N_11729,N_11086);
nor U12040 (N_12040,N_11033,N_11058);
or U12041 (N_12041,N_11836,N_11000);
nor U12042 (N_12042,N_11770,N_11266);
nand U12043 (N_12043,N_11160,N_11566);
nor U12044 (N_12044,N_11767,N_11925);
or U12045 (N_12045,N_11837,N_11010);
xor U12046 (N_12046,N_11939,N_11497);
xnor U12047 (N_12047,N_11377,N_11540);
nand U12048 (N_12048,N_11360,N_11411);
or U12049 (N_12049,N_11859,N_11976);
xnor U12050 (N_12050,N_11414,N_11208);
xnor U12051 (N_12051,N_11390,N_11254);
and U12052 (N_12052,N_11992,N_11060);
nand U12053 (N_12053,N_11748,N_11891);
and U12054 (N_12054,N_11115,N_11180);
or U12055 (N_12055,N_11541,N_11948);
nand U12056 (N_12056,N_11797,N_11814);
and U12057 (N_12057,N_11839,N_11016);
xnor U12058 (N_12058,N_11677,N_11006);
nand U12059 (N_12059,N_11473,N_11365);
and U12060 (N_12060,N_11022,N_11399);
or U12061 (N_12061,N_11819,N_11343);
nor U12062 (N_12062,N_11102,N_11339);
xnor U12063 (N_12063,N_11607,N_11237);
nand U12064 (N_12064,N_11659,N_11904);
and U12065 (N_12065,N_11766,N_11883);
or U12066 (N_12066,N_11635,N_11385);
and U12067 (N_12067,N_11896,N_11789);
or U12068 (N_12068,N_11561,N_11953);
and U12069 (N_12069,N_11557,N_11637);
or U12070 (N_12070,N_11503,N_11563);
nand U12071 (N_12071,N_11780,N_11038);
nor U12072 (N_12072,N_11112,N_11843);
or U12073 (N_12073,N_11162,N_11508);
nor U12074 (N_12074,N_11710,N_11671);
or U12075 (N_12075,N_11863,N_11879);
nand U12076 (N_12076,N_11422,N_11017);
or U12077 (N_12077,N_11446,N_11476);
or U12078 (N_12078,N_11370,N_11567);
and U12079 (N_12079,N_11207,N_11873);
and U12080 (N_12080,N_11096,N_11678);
nand U12081 (N_12081,N_11947,N_11182);
nand U12082 (N_12082,N_11256,N_11428);
or U12083 (N_12083,N_11787,N_11047);
xor U12084 (N_12084,N_11876,N_11545);
nor U12085 (N_12085,N_11649,N_11725);
nand U12086 (N_12086,N_11501,N_11617);
nand U12087 (N_12087,N_11185,N_11507);
nand U12088 (N_12088,N_11830,N_11187);
and U12089 (N_12089,N_11982,N_11090);
or U12090 (N_12090,N_11164,N_11903);
and U12091 (N_12091,N_11462,N_11550);
or U12092 (N_12092,N_11089,N_11580);
nand U12093 (N_12093,N_11867,N_11815);
nand U12094 (N_12094,N_11813,N_11855);
or U12095 (N_12095,N_11255,N_11838);
nand U12096 (N_12096,N_11981,N_11629);
xnor U12097 (N_12097,N_11675,N_11620);
xor U12098 (N_12098,N_11920,N_11149);
nand U12099 (N_12099,N_11394,N_11465);
nor U12100 (N_12100,N_11500,N_11223);
nand U12101 (N_12101,N_11973,N_11078);
and U12102 (N_12102,N_11094,N_11568);
and U12103 (N_12103,N_11652,N_11159);
xnor U12104 (N_12104,N_11851,N_11760);
nor U12105 (N_12105,N_11513,N_11193);
and U12106 (N_12106,N_11932,N_11850);
and U12107 (N_12107,N_11802,N_11028);
xor U12108 (N_12108,N_11273,N_11612);
nor U12109 (N_12109,N_11764,N_11436);
and U12110 (N_12110,N_11695,N_11282);
and U12111 (N_12111,N_11107,N_11077);
and U12112 (N_12112,N_11258,N_11795);
nand U12113 (N_12113,N_11081,N_11643);
xor U12114 (N_12114,N_11630,N_11387);
and U12115 (N_12115,N_11234,N_11080);
nor U12116 (N_12116,N_11585,N_11529);
xnor U12117 (N_12117,N_11449,N_11526);
or U12118 (N_12118,N_11167,N_11718);
nor U12119 (N_12119,N_11872,N_11480);
or U12120 (N_12120,N_11897,N_11531);
nand U12121 (N_12121,N_11834,N_11554);
nor U12122 (N_12122,N_11970,N_11655);
and U12123 (N_12123,N_11744,N_11311);
and U12124 (N_12124,N_11574,N_11322);
nand U12125 (N_12125,N_11692,N_11742);
and U12126 (N_12126,N_11220,N_11919);
nand U12127 (N_12127,N_11225,N_11316);
and U12128 (N_12128,N_11427,N_11001);
nand U12129 (N_12129,N_11573,N_11148);
or U12130 (N_12130,N_11884,N_11964);
xor U12131 (N_12131,N_11435,N_11290);
or U12132 (N_12132,N_11723,N_11980);
nand U12133 (N_12133,N_11827,N_11998);
or U12134 (N_12134,N_11845,N_11609);
xnor U12135 (N_12135,N_11986,N_11471);
or U12136 (N_12136,N_11453,N_11577);
xor U12137 (N_12137,N_11289,N_11353);
and U12138 (N_12138,N_11268,N_11023);
and U12139 (N_12139,N_11600,N_11553);
nand U12140 (N_12140,N_11842,N_11717);
nand U12141 (N_12141,N_11111,N_11810);
and U12142 (N_12142,N_11781,N_11665);
and U12143 (N_12143,N_11405,N_11504);
nor U12144 (N_12144,N_11011,N_11619);
xor U12145 (N_12145,N_11204,N_11494);
nand U12146 (N_12146,N_11288,N_11582);
nor U12147 (N_12147,N_11700,N_11962);
and U12148 (N_12148,N_11596,N_11232);
or U12149 (N_12149,N_11472,N_11482);
and U12150 (N_12150,N_11946,N_11581);
nor U12151 (N_12151,N_11579,N_11739);
xnor U12152 (N_12152,N_11794,N_11603);
nand U12153 (N_12153,N_11997,N_11224);
nor U12154 (N_12154,N_11702,N_11608);
nand U12155 (N_12155,N_11900,N_11790);
and U12156 (N_12156,N_11535,N_11865);
nor U12157 (N_12157,N_11378,N_11857);
xor U12158 (N_12158,N_11025,N_11915);
xor U12159 (N_12159,N_11034,N_11201);
nand U12160 (N_12160,N_11153,N_11388);
and U12161 (N_12161,N_11943,N_11119);
or U12162 (N_12162,N_11050,N_11833);
nor U12163 (N_12163,N_11999,N_11154);
nand U12164 (N_12164,N_11728,N_11045);
or U12165 (N_12165,N_11763,N_11687);
nor U12166 (N_12166,N_11601,N_11004);
and U12167 (N_12167,N_11812,N_11173);
or U12168 (N_12168,N_11961,N_11898);
and U12169 (N_12169,N_11368,N_11544);
nand U12170 (N_12170,N_11751,N_11253);
xnor U12171 (N_12171,N_11602,N_11046);
or U12172 (N_12172,N_11599,N_11731);
xnor U12173 (N_12173,N_11073,N_11909);
or U12174 (N_12174,N_11189,N_11406);
xnor U12175 (N_12175,N_11934,N_11869);
or U12176 (N_12176,N_11092,N_11648);
nand U12177 (N_12177,N_11595,N_11068);
nand U12178 (N_12178,N_11211,N_11194);
nand U12179 (N_12179,N_11908,N_11285);
xnor U12180 (N_12180,N_11260,N_11015);
xnor U12181 (N_12181,N_11989,N_11606);
nand U12182 (N_12182,N_11362,N_11926);
or U12183 (N_12183,N_11486,N_11262);
and U12184 (N_12184,N_11397,N_11460);
xnor U12185 (N_12185,N_11969,N_11594);
xor U12186 (N_12186,N_11181,N_11216);
nor U12187 (N_12187,N_11880,N_11831);
or U12188 (N_12188,N_11008,N_11135);
xor U12189 (N_12189,N_11251,N_11064);
or U12190 (N_12190,N_11707,N_11604);
xor U12191 (N_12191,N_11136,N_11854);
or U12192 (N_12192,N_11933,N_11518);
xnor U12193 (N_12193,N_11711,N_11881);
and U12194 (N_12194,N_11269,N_11506);
and U12195 (N_12195,N_11656,N_11424);
nor U12196 (N_12196,N_11348,N_11684);
nor U12197 (N_12197,N_11215,N_11227);
nand U12198 (N_12198,N_11994,N_11103);
and U12199 (N_12199,N_11457,N_11213);
nand U12200 (N_12200,N_11483,N_11546);
xnor U12201 (N_12201,N_11280,N_11720);
and U12202 (N_12202,N_11688,N_11168);
xnor U12203 (N_12203,N_11470,N_11287);
nor U12204 (N_12204,N_11129,N_11029);
nand U12205 (N_12205,N_11321,N_11514);
nand U12206 (N_12206,N_11757,N_11139);
nand U12207 (N_12207,N_11257,N_11383);
and U12208 (N_12208,N_11037,N_11170);
or U12209 (N_12209,N_11306,N_11323);
nand U12210 (N_12210,N_11091,N_11236);
or U12211 (N_12211,N_11404,N_11856);
and U12212 (N_12212,N_11724,N_11523);
nor U12213 (N_12213,N_11222,N_11432);
or U12214 (N_12214,N_11335,N_11515);
nor U12215 (N_12215,N_11464,N_11373);
xor U12216 (N_12216,N_11990,N_11924);
xnor U12217 (N_12217,N_11642,N_11584);
nor U12218 (N_12218,N_11907,N_11361);
nand U12219 (N_12219,N_11020,N_11041);
or U12220 (N_12220,N_11844,N_11210);
and U12221 (N_12221,N_11715,N_11542);
and U12222 (N_12222,N_11888,N_11138);
and U12223 (N_12223,N_11670,N_11988);
nand U12224 (N_12224,N_11987,N_11491);
nand U12225 (N_12225,N_11150,N_11634);
xor U12226 (N_12226,N_11698,N_11192);
nor U12227 (N_12227,N_11727,N_11440);
or U12228 (N_12228,N_11330,N_11931);
xnor U12229 (N_12229,N_11169,N_11799);
nor U12230 (N_12230,N_11828,N_11171);
or U12231 (N_12231,N_11562,N_11587);
or U12232 (N_12232,N_11380,N_11841);
nand U12233 (N_12233,N_11543,N_11735);
or U12234 (N_12234,N_11680,N_11292);
nor U12235 (N_12235,N_11755,N_11765);
nand U12236 (N_12236,N_11226,N_11940);
and U12237 (N_12237,N_11509,N_11127);
nor U12238 (N_12238,N_11699,N_11202);
or U12239 (N_12239,N_11570,N_11804);
nand U12240 (N_12240,N_11806,N_11488);
nand U12241 (N_12241,N_11826,N_11685);
or U12242 (N_12242,N_11305,N_11752);
nor U12243 (N_12243,N_11633,N_11442);
nor U12244 (N_12244,N_11691,N_11434);
and U12245 (N_12245,N_11293,N_11800);
xnor U12246 (N_12246,N_11113,N_11417);
xnor U12247 (N_12247,N_11184,N_11076);
nor U12248 (N_12248,N_11126,N_11104);
nand U12249 (N_12249,N_11108,N_11341);
and U12250 (N_12250,N_11221,N_11062);
xor U12251 (N_12251,N_11469,N_11605);
xor U12252 (N_12252,N_11758,N_11005);
nor U12253 (N_12253,N_11532,N_11333);
or U12254 (N_12254,N_11425,N_11142);
xor U12255 (N_12255,N_11179,N_11199);
xnor U12256 (N_12256,N_11668,N_11195);
or U12257 (N_12257,N_11935,N_11575);
and U12258 (N_12258,N_11451,N_11479);
nor U12259 (N_12259,N_11071,N_11929);
xnor U12260 (N_12260,N_11578,N_11589);
nand U12261 (N_12261,N_11384,N_11444);
or U12262 (N_12262,N_11618,N_11332);
xnor U12263 (N_12263,N_11552,N_11415);
xnor U12264 (N_12264,N_11636,N_11477);
xor U12265 (N_12265,N_11351,N_11949);
nor U12266 (N_12266,N_11349,N_11967);
nand U12267 (N_12267,N_11534,N_11172);
and U12268 (N_12268,N_11116,N_11918);
nand U12269 (N_12269,N_11053,N_11043);
xnor U12270 (N_12270,N_11291,N_11188);
nor U12271 (N_12271,N_11906,N_11018);
and U12272 (N_12272,N_11244,N_11416);
nor U12273 (N_12273,N_11125,N_11703);
or U12274 (N_12274,N_11864,N_11673);
nand U12275 (N_12275,N_11079,N_11913);
xor U12276 (N_12276,N_11134,N_11774);
or U12277 (N_12277,N_11014,N_11300);
xnor U12278 (N_12278,N_11959,N_11161);
xor U12279 (N_12279,N_11689,N_11274);
or U12280 (N_12280,N_11960,N_11709);
and U12281 (N_12281,N_11978,N_11610);
xor U12282 (N_12282,N_11042,N_11070);
xnor U12283 (N_12283,N_11654,N_11627);
and U12284 (N_12284,N_11923,N_11921);
and U12285 (N_12285,N_11312,N_11510);
nor U12286 (N_12286,N_11624,N_11147);
nor U12287 (N_12287,N_11628,N_11975);
xor U12288 (N_12288,N_11217,N_11463);
and U12289 (N_12289,N_11614,N_11893);
xor U12290 (N_12290,N_11517,N_11088);
nor U12291 (N_12291,N_11556,N_11722);
and U12292 (N_12292,N_11928,N_11538);
xor U12293 (N_12293,N_11808,N_11816);
nor U12294 (N_12294,N_11106,N_11205);
or U12295 (N_12295,N_11075,N_11146);
or U12296 (N_12296,N_11336,N_11985);
or U12297 (N_12297,N_11551,N_11597);
and U12298 (N_12298,N_11196,N_11536);
or U12299 (N_12299,N_11063,N_11467);
nand U12300 (N_12300,N_11298,N_11155);
nor U12301 (N_12301,N_11165,N_11905);
xor U12302 (N_12302,N_11952,N_11441);
and U12303 (N_12303,N_11026,N_11747);
or U12304 (N_12304,N_11007,N_11623);
nand U12305 (N_12305,N_11890,N_11308);
nor U12306 (N_12306,N_11342,N_11866);
nand U12307 (N_12307,N_11085,N_11771);
nand U12308 (N_12308,N_11400,N_11886);
nor U12309 (N_12309,N_11740,N_11295);
nor U12310 (N_12310,N_11681,N_11445);
or U12311 (N_12311,N_11301,N_11558);
nor U12312 (N_12312,N_11817,N_11957);
or U12313 (N_12313,N_11922,N_11738);
or U12314 (N_12314,N_11683,N_11803);
xnor U12315 (N_12315,N_11334,N_11299);
or U12316 (N_12316,N_11669,N_11374);
and U12317 (N_12317,N_11419,N_11835);
xor U12318 (N_12318,N_11097,N_11478);
or U12319 (N_12319,N_11328,N_11936);
and U12320 (N_12320,N_11183,N_11525);
and U12321 (N_12321,N_11458,N_11429);
nand U12322 (N_12322,N_11927,N_11966);
and U12323 (N_12323,N_11344,N_11521);
or U12324 (N_12324,N_11357,N_11426);
or U12325 (N_12325,N_11950,N_11484);
nand U12326 (N_12326,N_11013,N_11631);
nor U12327 (N_12327,N_11036,N_11917);
or U12328 (N_12328,N_11447,N_11977);
nor U12329 (N_12329,N_11069,N_11247);
and U12330 (N_12330,N_11363,N_11275);
and U12331 (N_12331,N_11591,N_11818);
or U12332 (N_12332,N_11235,N_11547);
or U12333 (N_12333,N_11701,N_11459);
xor U12334 (N_12334,N_11359,N_11231);
xnor U12335 (N_12335,N_11250,N_11396);
xor U12336 (N_12336,N_11303,N_11012);
and U12337 (N_12337,N_11796,N_11401);
nor U12338 (N_12338,N_11044,N_11559);
xnor U12339 (N_12339,N_11882,N_11002);
or U12340 (N_12340,N_11320,N_11793);
xor U12341 (N_12341,N_11945,N_11072);
nor U12342 (N_12342,N_11296,N_11265);
xor U12343 (N_12343,N_11971,N_11448);
nand U12344 (N_12344,N_11307,N_11052);
or U12345 (N_12345,N_11996,N_11032);
nor U12346 (N_12346,N_11832,N_11474);
or U12347 (N_12347,N_11569,N_11124);
and U12348 (N_12348,N_11972,N_11768);
nand U12349 (N_12349,N_11356,N_11246);
nand U12350 (N_12350,N_11286,N_11667);
nand U12351 (N_12351,N_11337,N_11495);
nor U12352 (N_12352,N_11120,N_11853);
nor U12353 (N_12353,N_11679,N_11598);
nor U12354 (N_12354,N_11788,N_11564);
and U12355 (N_12355,N_11761,N_11456);
and U12356 (N_12356,N_11249,N_11166);
xnor U12357 (N_12357,N_11369,N_11887);
or U12358 (N_12358,N_11346,N_11156);
nand U12359 (N_12359,N_11593,N_11721);
and U12360 (N_12360,N_11704,N_11241);
nor U12361 (N_12361,N_11439,N_11512);
and U12362 (N_12362,N_11862,N_11331);
and U12363 (N_12363,N_11065,N_11705);
and U12364 (N_12364,N_11885,N_11059);
nor U12365 (N_12365,N_11277,N_11548);
nor U12366 (N_12366,N_11481,N_11143);
and U12367 (N_12367,N_11565,N_11621);
or U12368 (N_12368,N_11466,N_11109);
nand U12369 (N_12369,N_11145,N_11734);
nand U12370 (N_12370,N_11736,N_11712);
nand U12371 (N_12371,N_11528,N_11242);
nand U12372 (N_12372,N_11054,N_11430);
xor U12373 (N_12373,N_11965,N_11782);
nand U12374 (N_12374,N_11749,N_11228);
and U12375 (N_12375,N_11682,N_11661);
nor U12376 (N_12376,N_11105,N_11338);
nor U12377 (N_12377,N_11502,N_11381);
nor U12378 (N_12378,N_11057,N_11658);
or U12379 (N_12379,N_11660,N_11646);
or U12380 (N_12380,N_11775,N_11386);
xnor U12381 (N_12381,N_11912,N_11792);
or U12382 (N_12382,N_11941,N_11772);
nor U12383 (N_12383,N_11176,N_11314);
and U12384 (N_12384,N_11706,N_11776);
and U12385 (N_12385,N_11499,N_11438);
nand U12386 (N_12386,N_11101,N_11811);
xor U12387 (N_12387,N_11352,N_11954);
and U12388 (N_12388,N_11995,N_11431);
and U12389 (N_12389,N_11530,N_11309);
nand U12390 (N_12390,N_11555,N_11413);
nand U12391 (N_12391,N_11402,N_11233);
or U12392 (N_12392,N_11737,N_11993);
xnor U12393 (N_12393,N_11031,N_11777);
and U12394 (N_12394,N_11327,N_11714);
xnor U12395 (N_12395,N_11611,N_11243);
xnor U12396 (N_12396,N_11372,N_11583);
and U12397 (N_12397,N_11393,N_11756);
and U12398 (N_12398,N_11412,N_11519);
nor U12399 (N_12399,N_11791,N_11039);
and U12400 (N_12400,N_11056,N_11144);
and U12401 (N_12401,N_11340,N_11590);
nand U12402 (N_12402,N_11003,N_11894);
nand U12403 (N_12403,N_11279,N_11778);
nand U12404 (N_12404,N_11686,N_11398);
nor U12405 (N_12405,N_11807,N_11930);
nor U12406 (N_12406,N_11892,N_11027);
xor U12407 (N_12407,N_11345,N_11693);
xnor U12408 (N_12408,N_11902,N_11586);
nor U12409 (N_12409,N_11653,N_11132);
or U12410 (N_12410,N_11496,N_11871);
nand U12411 (N_12411,N_11030,N_11592);
nor U12412 (N_12412,N_11730,N_11571);
nor U12413 (N_12413,N_11190,N_11200);
nand U12414 (N_12414,N_11759,N_11140);
nand U12415 (N_12415,N_11672,N_11318);
xor U12416 (N_12416,N_11666,N_11638);
nand U12417 (N_12417,N_11874,N_11868);
nor U12418 (N_12418,N_11284,N_11762);
nor U12419 (N_12419,N_11152,N_11889);
or U12420 (N_12420,N_11157,N_11021);
nor U12421 (N_12421,N_11177,N_11895);
xnor U12422 (N_12422,N_11267,N_11093);
nor U12423 (N_12423,N_11613,N_11743);
and U12424 (N_12424,N_11240,N_11641);
xnor U12425 (N_12425,N_11082,N_11490);
xor U12426 (N_12426,N_11117,N_11650);
nor U12427 (N_12427,N_11632,N_11358);
or U12428 (N_12428,N_11066,N_11492);
nor U12429 (N_12429,N_11375,N_11645);
or U12430 (N_12430,N_11218,N_11259);
nor U12431 (N_12431,N_11572,N_11910);
or U12432 (N_12432,N_11640,N_11820);
nor U12433 (N_12433,N_11916,N_11389);
nand U12434 (N_12434,N_11773,N_11616);
and U12435 (N_12435,N_11178,N_11329);
nand U12436 (N_12436,N_11979,N_11264);
and U12437 (N_12437,N_11870,N_11983);
nor U12438 (N_12438,N_11048,N_11418);
nand U12439 (N_12439,N_11785,N_11647);
and U12440 (N_12440,N_11639,N_11355);
or U12441 (N_12441,N_11098,N_11485);
or U12442 (N_12442,N_11696,N_11750);
xnor U12443 (N_12443,N_11261,N_11852);
xnor U12444 (N_12444,N_11741,N_11840);
or U12445 (N_12445,N_11848,N_11252);
xor U12446 (N_12446,N_11809,N_11158);
and U12447 (N_12447,N_11270,N_11450);
and U12448 (N_12448,N_11516,N_11163);
nor U12449 (N_12449,N_11313,N_11433);
nor U12450 (N_12450,N_11822,N_11786);
xor U12451 (N_12451,N_11376,N_11524);
nor U12452 (N_12452,N_11382,N_11511);
xor U12453 (N_12453,N_11203,N_11674);
and U12454 (N_12454,N_11823,N_11694);
or U12455 (N_12455,N_11733,N_11533);
and U12456 (N_12456,N_11324,N_11212);
xor U12457 (N_12457,N_11095,N_11662);
and U12458 (N_12458,N_11560,N_11100);
nand U12459 (N_12459,N_11131,N_11783);
nand U12460 (N_12460,N_11664,N_11407);
xnor U12461 (N_12461,N_11719,N_11408);
nand U12462 (N_12462,N_11651,N_11825);
nand U12463 (N_12463,N_11644,N_11174);
xnor U12464 (N_12464,N_11061,N_11937);
nand U12465 (N_12465,N_11878,N_11697);
nand U12466 (N_12466,N_11371,N_11214);
and U12467 (N_12467,N_11461,N_11549);
and U12468 (N_12468,N_11588,N_11310);
nand U12469 (N_12469,N_11421,N_11281);
nor U12470 (N_12470,N_11527,N_11769);
nor U12471 (N_12471,N_11272,N_11911);
and U12472 (N_12472,N_11974,N_11239);
and U12473 (N_12473,N_11452,N_11024);
nor U12474 (N_12474,N_11420,N_11410);
xor U12475 (N_12475,N_11186,N_11409);
nand U12476 (N_12476,N_11087,N_11325);
and U12477 (N_12477,N_11326,N_11366);
nor U12478 (N_12478,N_11475,N_11084);
xor U12479 (N_12479,N_11151,N_11437);
and U12480 (N_12480,N_11276,N_11230);
nor U12481 (N_12481,N_11858,N_11128);
nor U12482 (N_12482,N_11498,N_11114);
nand U12483 (N_12483,N_11191,N_11732);
and U12484 (N_12484,N_11238,N_11821);
xnor U12485 (N_12485,N_11801,N_11278);
or U12486 (N_12486,N_11454,N_11824);
and U12487 (N_12487,N_11245,N_11319);
or U12488 (N_12488,N_11083,N_11443);
xor U12489 (N_12489,N_11779,N_11009);
or U12490 (N_12490,N_11537,N_11942);
nand U12491 (N_12491,N_11229,N_11198);
xor U12492 (N_12492,N_11122,N_11049);
or U12493 (N_12493,N_11798,N_11708);
nand U12494 (N_12494,N_11123,N_11956);
xor U12495 (N_12495,N_11784,N_11963);
xnor U12496 (N_12496,N_11615,N_11468);
or U12497 (N_12497,N_11055,N_11121);
xor U12498 (N_12498,N_11846,N_11626);
nor U12499 (N_12499,N_11317,N_11423);
and U12500 (N_12500,N_11074,N_11845);
xor U12501 (N_12501,N_11900,N_11087);
and U12502 (N_12502,N_11758,N_11345);
and U12503 (N_12503,N_11004,N_11661);
nand U12504 (N_12504,N_11147,N_11707);
xor U12505 (N_12505,N_11052,N_11230);
and U12506 (N_12506,N_11536,N_11281);
or U12507 (N_12507,N_11734,N_11118);
nor U12508 (N_12508,N_11145,N_11756);
and U12509 (N_12509,N_11099,N_11570);
xor U12510 (N_12510,N_11515,N_11348);
nand U12511 (N_12511,N_11810,N_11942);
xor U12512 (N_12512,N_11494,N_11437);
nor U12513 (N_12513,N_11449,N_11540);
or U12514 (N_12514,N_11485,N_11173);
nand U12515 (N_12515,N_11395,N_11844);
and U12516 (N_12516,N_11899,N_11255);
nor U12517 (N_12517,N_11006,N_11036);
nor U12518 (N_12518,N_11038,N_11839);
and U12519 (N_12519,N_11403,N_11096);
xor U12520 (N_12520,N_11953,N_11405);
and U12521 (N_12521,N_11358,N_11214);
xnor U12522 (N_12522,N_11933,N_11881);
nand U12523 (N_12523,N_11769,N_11220);
nand U12524 (N_12524,N_11492,N_11701);
nand U12525 (N_12525,N_11512,N_11719);
and U12526 (N_12526,N_11012,N_11741);
or U12527 (N_12527,N_11784,N_11080);
xor U12528 (N_12528,N_11246,N_11409);
xor U12529 (N_12529,N_11856,N_11484);
nand U12530 (N_12530,N_11868,N_11536);
xnor U12531 (N_12531,N_11121,N_11828);
xnor U12532 (N_12532,N_11133,N_11252);
nor U12533 (N_12533,N_11187,N_11744);
nor U12534 (N_12534,N_11731,N_11393);
and U12535 (N_12535,N_11284,N_11826);
and U12536 (N_12536,N_11247,N_11443);
xnor U12537 (N_12537,N_11518,N_11345);
nor U12538 (N_12538,N_11638,N_11599);
nand U12539 (N_12539,N_11673,N_11457);
nor U12540 (N_12540,N_11664,N_11323);
nand U12541 (N_12541,N_11213,N_11080);
xor U12542 (N_12542,N_11312,N_11231);
nor U12543 (N_12543,N_11818,N_11798);
xnor U12544 (N_12544,N_11911,N_11323);
nor U12545 (N_12545,N_11029,N_11294);
nor U12546 (N_12546,N_11598,N_11581);
or U12547 (N_12547,N_11897,N_11804);
xnor U12548 (N_12548,N_11958,N_11890);
nor U12549 (N_12549,N_11464,N_11336);
and U12550 (N_12550,N_11543,N_11893);
nand U12551 (N_12551,N_11975,N_11762);
nor U12552 (N_12552,N_11249,N_11296);
xnor U12553 (N_12553,N_11212,N_11628);
nor U12554 (N_12554,N_11979,N_11818);
nor U12555 (N_12555,N_11308,N_11867);
and U12556 (N_12556,N_11785,N_11349);
nor U12557 (N_12557,N_11701,N_11872);
and U12558 (N_12558,N_11298,N_11712);
nand U12559 (N_12559,N_11308,N_11079);
xnor U12560 (N_12560,N_11689,N_11341);
and U12561 (N_12561,N_11060,N_11258);
nor U12562 (N_12562,N_11188,N_11682);
xnor U12563 (N_12563,N_11729,N_11456);
or U12564 (N_12564,N_11607,N_11483);
nor U12565 (N_12565,N_11707,N_11108);
nand U12566 (N_12566,N_11260,N_11611);
or U12567 (N_12567,N_11739,N_11738);
and U12568 (N_12568,N_11043,N_11644);
and U12569 (N_12569,N_11642,N_11440);
nor U12570 (N_12570,N_11520,N_11098);
nand U12571 (N_12571,N_11301,N_11160);
or U12572 (N_12572,N_11227,N_11402);
nand U12573 (N_12573,N_11260,N_11042);
and U12574 (N_12574,N_11873,N_11490);
or U12575 (N_12575,N_11055,N_11927);
nor U12576 (N_12576,N_11897,N_11848);
xnor U12577 (N_12577,N_11788,N_11603);
nand U12578 (N_12578,N_11091,N_11265);
nor U12579 (N_12579,N_11578,N_11049);
and U12580 (N_12580,N_11240,N_11454);
or U12581 (N_12581,N_11207,N_11792);
or U12582 (N_12582,N_11496,N_11575);
nand U12583 (N_12583,N_11160,N_11836);
and U12584 (N_12584,N_11799,N_11123);
xor U12585 (N_12585,N_11653,N_11582);
nor U12586 (N_12586,N_11337,N_11232);
or U12587 (N_12587,N_11114,N_11902);
nand U12588 (N_12588,N_11048,N_11870);
or U12589 (N_12589,N_11665,N_11966);
xor U12590 (N_12590,N_11464,N_11791);
or U12591 (N_12591,N_11275,N_11524);
nand U12592 (N_12592,N_11219,N_11863);
nand U12593 (N_12593,N_11964,N_11248);
or U12594 (N_12594,N_11421,N_11775);
xor U12595 (N_12595,N_11782,N_11689);
nor U12596 (N_12596,N_11999,N_11422);
nand U12597 (N_12597,N_11669,N_11309);
or U12598 (N_12598,N_11676,N_11830);
xor U12599 (N_12599,N_11659,N_11860);
or U12600 (N_12600,N_11069,N_11494);
and U12601 (N_12601,N_11689,N_11876);
and U12602 (N_12602,N_11071,N_11660);
or U12603 (N_12603,N_11333,N_11541);
and U12604 (N_12604,N_11927,N_11427);
nor U12605 (N_12605,N_11338,N_11660);
or U12606 (N_12606,N_11863,N_11081);
and U12607 (N_12607,N_11166,N_11974);
nor U12608 (N_12608,N_11522,N_11689);
or U12609 (N_12609,N_11445,N_11187);
xnor U12610 (N_12610,N_11406,N_11084);
and U12611 (N_12611,N_11194,N_11752);
nand U12612 (N_12612,N_11228,N_11237);
and U12613 (N_12613,N_11716,N_11826);
nand U12614 (N_12614,N_11001,N_11465);
and U12615 (N_12615,N_11190,N_11583);
and U12616 (N_12616,N_11462,N_11872);
or U12617 (N_12617,N_11929,N_11784);
xnor U12618 (N_12618,N_11106,N_11451);
nor U12619 (N_12619,N_11962,N_11272);
nand U12620 (N_12620,N_11541,N_11042);
xor U12621 (N_12621,N_11247,N_11767);
xor U12622 (N_12622,N_11011,N_11256);
nor U12623 (N_12623,N_11887,N_11221);
or U12624 (N_12624,N_11061,N_11372);
or U12625 (N_12625,N_11819,N_11478);
xnor U12626 (N_12626,N_11251,N_11874);
nand U12627 (N_12627,N_11552,N_11116);
and U12628 (N_12628,N_11772,N_11117);
nand U12629 (N_12629,N_11373,N_11303);
and U12630 (N_12630,N_11845,N_11020);
nor U12631 (N_12631,N_11762,N_11712);
xnor U12632 (N_12632,N_11569,N_11412);
nand U12633 (N_12633,N_11507,N_11913);
nand U12634 (N_12634,N_11311,N_11236);
nand U12635 (N_12635,N_11162,N_11181);
nand U12636 (N_12636,N_11716,N_11051);
nand U12637 (N_12637,N_11719,N_11104);
and U12638 (N_12638,N_11398,N_11553);
nor U12639 (N_12639,N_11419,N_11626);
xnor U12640 (N_12640,N_11027,N_11225);
nand U12641 (N_12641,N_11073,N_11984);
nor U12642 (N_12642,N_11815,N_11223);
or U12643 (N_12643,N_11681,N_11473);
xor U12644 (N_12644,N_11249,N_11792);
and U12645 (N_12645,N_11865,N_11216);
xnor U12646 (N_12646,N_11688,N_11210);
xor U12647 (N_12647,N_11550,N_11188);
nand U12648 (N_12648,N_11861,N_11811);
nand U12649 (N_12649,N_11051,N_11309);
and U12650 (N_12650,N_11371,N_11358);
or U12651 (N_12651,N_11538,N_11903);
nand U12652 (N_12652,N_11504,N_11980);
xnor U12653 (N_12653,N_11518,N_11220);
or U12654 (N_12654,N_11625,N_11796);
or U12655 (N_12655,N_11479,N_11883);
and U12656 (N_12656,N_11090,N_11682);
nand U12657 (N_12657,N_11442,N_11366);
or U12658 (N_12658,N_11747,N_11057);
and U12659 (N_12659,N_11411,N_11565);
xnor U12660 (N_12660,N_11839,N_11278);
or U12661 (N_12661,N_11317,N_11692);
nor U12662 (N_12662,N_11648,N_11732);
nand U12663 (N_12663,N_11634,N_11184);
xor U12664 (N_12664,N_11144,N_11825);
nand U12665 (N_12665,N_11500,N_11031);
xor U12666 (N_12666,N_11417,N_11094);
xor U12667 (N_12667,N_11261,N_11424);
xnor U12668 (N_12668,N_11430,N_11232);
and U12669 (N_12669,N_11823,N_11437);
nor U12670 (N_12670,N_11666,N_11475);
nand U12671 (N_12671,N_11963,N_11058);
nand U12672 (N_12672,N_11934,N_11315);
nor U12673 (N_12673,N_11362,N_11352);
nor U12674 (N_12674,N_11051,N_11657);
or U12675 (N_12675,N_11768,N_11145);
nor U12676 (N_12676,N_11409,N_11977);
nor U12677 (N_12677,N_11788,N_11857);
nand U12678 (N_12678,N_11095,N_11770);
nand U12679 (N_12679,N_11588,N_11755);
and U12680 (N_12680,N_11071,N_11566);
nand U12681 (N_12681,N_11169,N_11704);
nand U12682 (N_12682,N_11934,N_11471);
or U12683 (N_12683,N_11134,N_11272);
or U12684 (N_12684,N_11046,N_11240);
nor U12685 (N_12685,N_11368,N_11461);
or U12686 (N_12686,N_11129,N_11257);
and U12687 (N_12687,N_11899,N_11321);
nand U12688 (N_12688,N_11790,N_11594);
and U12689 (N_12689,N_11635,N_11199);
xnor U12690 (N_12690,N_11843,N_11163);
or U12691 (N_12691,N_11110,N_11372);
xor U12692 (N_12692,N_11142,N_11906);
xor U12693 (N_12693,N_11451,N_11068);
xnor U12694 (N_12694,N_11637,N_11576);
nand U12695 (N_12695,N_11254,N_11455);
nor U12696 (N_12696,N_11015,N_11830);
or U12697 (N_12697,N_11389,N_11950);
or U12698 (N_12698,N_11708,N_11317);
nand U12699 (N_12699,N_11804,N_11085);
nor U12700 (N_12700,N_11970,N_11053);
nor U12701 (N_12701,N_11573,N_11565);
and U12702 (N_12702,N_11091,N_11562);
nor U12703 (N_12703,N_11300,N_11478);
or U12704 (N_12704,N_11786,N_11165);
nand U12705 (N_12705,N_11394,N_11169);
nor U12706 (N_12706,N_11506,N_11844);
nand U12707 (N_12707,N_11445,N_11742);
nor U12708 (N_12708,N_11583,N_11011);
nor U12709 (N_12709,N_11965,N_11837);
xor U12710 (N_12710,N_11771,N_11199);
nor U12711 (N_12711,N_11691,N_11547);
and U12712 (N_12712,N_11769,N_11635);
and U12713 (N_12713,N_11626,N_11387);
and U12714 (N_12714,N_11008,N_11139);
or U12715 (N_12715,N_11847,N_11953);
xnor U12716 (N_12716,N_11465,N_11271);
or U12717 (N_12717,N_11441,N_11323);
xnor U12718 (N_12718,N_11187,N_11728);
xnor U12719 (N_12719,N_11846,N_11804);
xor U12720 (N_12720,N_11862,N_11208);
or U12721 (N_12721,N_11526,N_11438);
nand U12722 (N_12722,N_11434,N_11939);
and U12723 (N_12723,N_11360,N_11662);
nor U12724 (N_12724,N_11734,N_11530);
xor U12725 (N_12725,N_11676,N_11852);
or U12726 (N_12726,N_11596,N_11019);
nor U12727 (N_12727,N_11892,N_11428);
xor U12728 (N_12728,N_11232,N_11579);
or U12729 (N_12729,N_11902,N_11367);
xnor U12730 (N_12730,N_11929,N_11006);
xor U12731 (N_12731,N_11644,N_11969);
nand U12732 (N_12732,N_11680,N_11531);
xor U12733 (N_12733,N_11137,N_11333);
nand U12734 (N_12734,N_11532,N_11527);
nor U12735 (N_12735,N_11427,N_11125);
xor U12736 (N_12736,N_11788,N_11398);
and U12737 (N_12737,N_11995,N_11664);
and U12738 (N_12738,N_11522,N_11155);
nor U12739 (N_12739,N_11684,N_11262);
nand U12740 (N_12740,N_11181,N_11173);
nor U12741 (N_12741,N_11217,N_11909);
or U12742 (N_12742,N_11512,N_11913);
or U12743 (N_12743,N_11252,N_11815);
and U12744 (N_12744,N_11462,N_11729);
and U12745 (N_12745,N_11947,N_11446);
xnor U12746 (N_12746,N_11929,N_11816);
xnor U12747 (N_12747,N_11756,N_11839);
xor U12748 (N_12748,N_11211,N_11600);
xor U12749 (N_12749,N_11873,N_11589);
nand U12750 (N_12750,N_11353,N_11206);
or U12751 (N_12751,N_11587,N_11038);
or U12752 (N_12752,N_11257,N_11615);
xor U12753 (N_12753,N_11348,N_11147);
nor U12754 (N_12754,N_11740,N_11721);
and U12755 (N_12755,N_11447,N_11732);
or U12756 (N_12756,N_11072,N_11543);
or U12757 (N_12757,N_11788,N_11463);
nand U12758 (N_12758,N_11904,N_11556);
and U12759 (N_12759,N_11868,N_11838);
or U12760 (N_12760,N_11307,N_11709);
nand U12761 (N_12761,N_11268,N_11941);
nor U12762 (N_12762,N_11600,N_11676);
nand U12763 (N_12763,N_11672,N_11838);
and U12764 (N_12764,N_11843,N_11140);
xnor U12765 (N_12765,N_11821,N_11568);
nand U12766 (N_12766,N_11564,N_11486);
xnor U12767 (N_12767,N_11225,N_11421);
xor U12768 (N_12768,N_11436,N_11510);
and U12769 (N_12769,N_11815,N_11982);
xor U12770 (N_12770,N_11831,N_11680);
nor U12771 (N_12771,N_11639,N_11769);
or U12772 (N_12772,N_11824,N_11438);
nand U12773 (N_12773,N_11083,N_11254);
nand U12774 (N_12774,N_11650,N_11366);
nand U12775 (N_12775,N_11975,N_11531);
xor U12776 (N_12776,N_11521,N_11774);
and U12777 (N_12777,N_11288,N_11810);
xor U12778 (N_12778,N_11642,N_11236);
nand U12779 (N_12779,N_11530,N_11288);
and U12780 (N_12780,N_11859,N_11046);
xnor U12781 (N_12781,N_11353,N_11458);
or U12782 (N_12782,N_11176,N_11270);
nor U12783 (N_12783,N_11910,N_11028);
or U12784 (N_12784,N_11872,N_11485);
xor U12785 (N_12785,N_11197,N_11628);
or U12786 (N_12786,N_11530,N_11332);
nand U12787 (N_12787,N_11612,N_11064);
xor U12788 (N_12788,N_11367,N_11059);
and U12789 (N_12789,N_11295,N_11411);
nand U12790 (N_12790,N_11000,N_11850);
or U12791 (N_12791,N_11663,N_11995);
or U12792 (N_12792,N_11819,N_11654);
xnor U12793 (N_12793,N_11497,N_11738);
or U12794 (N_12794,N_11045,N_11916);
or U12795 (N_12795,N_11428,N_11168);
nor U12796 (N_12796,N_11138,N_11353);
nand U12797 (N_12797,N_11740,N_11521);
nor U12798 (N_12798,N_11304,N_11341);
or U12799 (N_12799,N_11834,N_11694);
xor U12800 (N_12800,N_11960,N_11140);
nor U12801 (N_12801,N_11550,N_11547);
nor U12802 (N_12802,N_11309,N_11106);
or U12803 (N_12803,N_11594,N_11764);
nand U12804 (N_12804,N_11946,N_11729);
nor U12805 (N_12805,N_11668,N_11953);
or U12806 (N_12806,N_11848,N_11999);
xor U12807 (N_12807,N_11019,N_11752);
or U12808 (N_12808,N_11635,N_11396);
nand U12809 (N_12809,N_11114,N_11732);
or U12810 (N_12810,N_11765,N_11936);
and U12811 (N_12811,N_11793,N_11695);
xor U12812 (N_12812,N_11464,N_11866);
nand U12813 (N_12813,N_11423,N_11119);
nand U12814 (N_12814,N_11895,N_11183);
xnor U12815 (N_12815,N_11918,N_11742);
xor U12816 (N_12816,N_11399,N_11194);
xor U12817 (N_12817,N_11037,N_11606);
or U12818 (N_12818,N_11619,N_11117);
or U12819 (N_12819,N_11693,N_11747);
nand U12820 (N_12820,N_11482,N_11735);
nor U12821 (N_12821,N_11061,N_11075);
or U12822 (N_12822,N_11597,N_11348);
or U12823 (N_12823,N_11047,N_11051);
nor U12824 (N_12824,N_11845,N_11550);
nand U12825 (N_12825,N_11764,N_11103);
and U12826 (N_12826,N_11032,N_11380);
or U12827 (N_12827,N_11500,N_11816);
xor U12828 (N_12828,N_11342,N_11818);
nor U12829 (N_12829,N_11259,N_11204);
or U12830 (N_12830,N_11919,N_11579);
nor U12831 (N_12831,N_11668,N_11955);
and U12832 (N_12832,N_11329,N_11622);
nand U12833 (N_12833,N_11599,N_11176);
and U12834 (N_12834,N_11836,N_11918);
or U12835 (N_12835,N_11379,N_11716);
nand U12836 (N_12836,N_11933,N_11671);
and U12837 (N_12837,N_11226,N_11868);
nor U12838 (N_12838,N_11141,N_11448);
or U12839 (N_12839,N_11977,N_11149);
xnor U12840 (N_12840,N_11975,N_11598);
nand U12841 (N_12841,N_11463,N_11296);
nor U12842 (N_12842,N_11083,N_11424);
xor U12843 (N_12843,N_11025,N_11418);
and U12844 (N_12844,N_11051,N_11993);
nor U12845 (N_12845,N_11766,N_11212);
nor U12846 (N_12846,N_11487,N_11398);
xnor U12847 (N_12847,N_11830,N_11590);
xor U12848 (N_12848,N_11276,N_11962);
and U12849 (N_12849,N_11427,N_11347);
or U12850 (N_12850,N_11485,N_11288);
nor U12851 (N_12851,N_11150,N_11020);
nor U12852 (N_12852,N_11905,N_11877);
nand U12853 (N_12853,N_11717,N_11414);
or U12854 (N_12854,N_11022,N_11464);
nor U12855 (N_12855,N_11138,N_11329);
and U12856 (N_12856,N_11700,N_11075);
and U12857 (N_12857,N_11992,N_11737);
nand U12858 (N_12858,N_11166,N_11404);
or U12859 (N_12859,N_11245,N_11966);
and U12860 (N_12860,N_11230,N_11035);
and U12861 (N_12861,N_11317,N_11131);
or U12862 (N_12862,N_11659,N_11338);
nor U12863 (N_12863,N_11033,N_11120);
xor U12864 (N_12864,N_11015,N_11392);
xnor U12865 (N_12865,N_11265,N_11065);
or U12866 (N_12866,N_11163,N_11672);
nor U12867 (N_12867,N_11048,N_11769);
and U12868 (N_12868,N_11599,N_11975);
nand U12869 (N_12869,N_11524,N_11887);
nand U12870 (N_12870,N_11828,N_11165);
and U12871 (N_12871,N_11718,N_11438);
and U12872 (N_12872,N_11586,N_11164);
nor U12873 (N_12873,N_11028,N_11131);
nor U12874 (N_12874,N_11734,N_11787);
nand U12875 (N_12875,N_11950,N_11705);
nand U12876 (N_12876,N_11985,N_11227);
nand U12877 (N_12877,N_11942,N_11399);
nor U12878 (N_12878,N_11045,N_11415);
nor U12879 (N_12879,N_11261,N_11029);
nor U12880 (N_12880,N_11538,N_11020);
and U12881 (N_12881,N_11281,N_11467);
nand U12882 (N_12882,N_11890,N_11006);
xnor U12883 (N_12883,N_11701,N_11533);
nand U12884 (N_12884,N_11231,N_11877);
nand U12885 (N_12885,N_11380,N_11721);
nor U12886 (N_12886,N_11828,N_11208);
and U12887 (N_12887,N_11092,N_11259);
xor U12888 (N_12888,N_11757,N_11853);
and U12889 (N_12889,N_11623,N_11712);
or U12890 (N_12890,N_11453,N_11197);
or U12891 (N_12891,N_11311,N_11411);
or U12892 (N_12892,N_11678,N_11339);
and U12893 (N_12893,N_11703,N_11980);
and U12894 (N_12894,N_11271,N_11201);
xor U12895 (N_12895,N_11747,N_11824);
or U12896 (N_12896,N_11964,N_11201);
nor U12897 (N_12897,N_11927,N_11388);
or U12898 (N_12898,N_11451,N_11594);
xor U12899 (N_12899,N_11834,N_11173);
xor U12900 (N_12900,N_11160,N_11977);
and U12901 (N_12901,N_11973,N_11291);
or U12902 (N_12902,N_11287,N_11703);
xnor U12903 (N_12903,N_11757,N_11616);
and U12904 (N_12904,N_11080,N_11127);
nor U12905 (N_12905,N_11114,N_11700);
nand U12906 (N_12906,N_11590,N_11526);
nor U12907 (N_12907,N_11545,N_11881);
and U12908 (N_12908,N_11439,N_11982);
xnor U12909 (N_12909,N_11062,N_11624);
nor U12910 (N_12910,N_11096,N_11275);
nand U12911 (N_12911,N_11424,N_11186);
nor U12912 (N_12912,N_11998,N_11913);
nor U12913 (N_12913,N_11263,N_11403);
or U12914 (N_12914,N_11493,N_11544);
and U12915 (N_12915,N_11416,N_11666);
nand U12916 (N_12916,N_11126,N_11517);
nor U12917 (N_12917,N_11193,N_11163);
xor U12918 (N_12918,N_11337,N_11738);
nor U12919 (N_12919,N_11501,N_11482);
nand U12920 (N_12920,N_11358,N_11573);
or U12921 (N_12921,N_11738,N_11149);
nand U12922 (N_12922,N_11969,N_11883);
nand U12923 (N_12923,N_11498,N_11828);
or U12924 (N_12924,N_11633,N_11815);
nand U12925 (N_12925,N_11768,N_11868);
nand U12926 (N_12926,N_11593,N_11371);
or U12927 (N_12927,N_11249,N_11653);
nor U12928 (N_12928,N_11923,N_11133);
or U12929 (N_12929,N_11758,N_11693);
or U12930 (N_12930,N_11516,N_11556);
xor U12931 (N_12931,N_11382,N_11551);
xnor U12932 (N_12932,N_11220,N_11581);
nor U12933 (N_12933,N_11938,N_11873);
and U12934 (N_12934,N_11506,N_11432);
or U12935 (N_12935,N_11621,N_11376);
xor U12936 (N_12936,N_11747,N_11038);
nand U12937 (N_12937,N_11950,N_11585);
and U12938 (N_12938,N_11093,N_11081);
and U12939 (N_12939,N_11750,N_11423);
or U12940 (N_12940,N_11463,N_11471);
xor U12941 (N_12941,N_11921,N_11932);
nor U12942 (N_12942,N_11314,N_11980);
xor U12943 (N_12943,N_11279,N_11108);
nand U12944 (N_12944,N_11034,N_11167);
nand U12945 (N_12945,N_11109,N_11864);
nor U12946 (N_12946,N_11505,N_11818);
xnor U12947 (N_12947,N_11069,N_11142);
nand U12948 (N_12948,N_11183,N_11541);
and U12949 (N_12949,N_11604,N_11452);
nor U12950 (N_12950,N_11832,N_11356);
or U12951 (N_12951,N_11453,N_11992);
or U12952 (N_12952,N_11031,N_11551);
xnor U12953 (N_12953,N_11899,N_11031);
xnor U12954 (N_12954,N_11087,N_11726);
nand U12955 (N_12955,N_11205,N_11105);
xnor U12956 (N_12956,N_11611,N_11845);
xor U12957 (N_12957,N_11469,N_11513);
xor U12958 (N_12958,N_11551,N_11185);
nand U12959 (N_12959,N_11412,N_11530);
xor U12960 (N_12960,N_11742,N_11841);
and U12961 (N_12961,N_11084,N_11498);
nand U12962 (N_12962,N_11571,N_11909);
and U12963 (N_12963,N_11881,N_11524);
nor U12964 (N_12964,N_11106,N_11178);
xnor U12965 (N_12965,N_11165,N_11109);
nor U12966 (N_12966,N_11577,N_11946);
nor U12967 (N_12967,N_11535,N_11714);
nand U12968 (N_12968,N_11580,N_11187);
xor U12969 (N_12969,N_11928,N_11855);
nand U12970 (N_12970,N_11894,N_11056);
nand U12971 (N_12971,N_11293,N_11409);
and U12972 (N_12972,N_11134,N_11453);
xnor U12973 (N_12973,N_11199,N_11615);
xor U12974 (N_12974,N_11280,N_11016);
and U12975 (N_12975,N_11911,N_11343);
nand U12976 (N_12976,N_11017,N_11083);
nor U12977 (N_12977,N_11830,N_11886);
nand U12978 (N_12978,N_11039,N_11530);
xnor U12979 (N_12979,N_11351,N_11962);
nand U12980 (N_12980,N_11258,N_11398);
and U12981 (N_12981,N_11926,N_11867);
nor U12982 (N_12982,N_11013,N_11747);
xor U12983 (N_12983,N_11041,N_11118);
or U12984 (N_12984,N_11890,N_11899);
xnor U12985 (N_12985,N_11872,N_11281);
xor U12986 (N_12986,N_11674,N_11707);
or U12987 (N_12987,N_11254,N_11846);
nand U12988 (N_12988,N_11978,N_11746);
or U12989 (N_12989,N_11658,N_11773);
or U12990 (N_12990,N_11479,N_11822);
or U12991 (N_12991,N_11141,N_11622);
nor U12992 (N_12992,N_11373,N_11365);
nand U12993 (N_12993,N_11144,N_11074);
or U12994 (N_12994,N_11639,N_11759);
nand U12995 (N_12995,N_11730,N_11835);
or U12996 (N_12996,N_11370,N_11209);
xnor U12997 (N_12997,N_11985,N_11718);
and U12998 (N_12998,N_11334,N_11428);
nor U12999 (N_12999,N_11015,N_11587);
nor U13000 (N_13000,N_12593,N_12587);
xnor U13001 (N_13001,N_12340,N_12537);
xnor U13002 (N_13002,N_12014,N_12444);
nand U13003 (N_13003,N_12591,N_12749);
or U13004 (N_13004,N_12582,N_12220);
nor U13005 (N_13005,N_12736,N_12830);
or U13006 (N_13006,N_12823,N_12527);
nor U13007 (N_13007,N_12311,N_12520);
or U13008 (N_13008,N_12882,N_12304);
xor U13009 (N_13009,N_12975,N_12091);
nor U13010 (N_13010,N_12495,N_12522);
nand U13011 (N_13011,N_12499,N_12891);
and U13012 (N_13012,N_12068,N_12667);
or U13013 (N_13013,N_12894,N_12023);
and U13014 (N_13014,N_12654,N_12528);
and U13015 (N_13015,N_12008,N_12459);
or U13016 (N_13016,N_12341,N_12945);
nand U13017 (N_13017,N_12208,N_12908);
and U13018 (N_13018,N_12717,N_12511);
and U13019 (N_13019,N_12431,N_12984);
nor U13020 (N_13020,N_12079,N_12930);
nor U13021 (N_13021,N_12623,N_12964);
nand U13022 (N_13022,N_12162,N_12506);
xor U13023 (N_13023,N_12962,N_12998);
and U13024 (N_13024,N_12138,N_12308);
nor U13025 (N_13025,N_12575,N_12886);
xor U13026 (N_13026,N_12562,N_12172);
and U13027 (N_13027,N_12036,N_12057);
nand U13028 (N_13028,N_12405,N_12484);
nor U13029 (N_13029,N_12878,N_12094);
nor U13030 (N_13030,N_12106,N_12325);
xor U13031 (N_13031,N_12584,N_12293);
and U13032 (N_13032,N_12224,N_12988);
and U13033 (N_13033,N_12326,N_12342);
nor U13034 (N_13034,N_12135,N_12842);
xor U13035 (N_13035,N_12912,N_12190);
nor U13036 (N_13036,N_12048,N_12229);
nor U13037 (N_13037,N_12982,N_12480);
or U13038 (N_13038,N_12486,N_12840);
or U13039 (N_13039,N_12577,N_12195);
or U13040 (N_13040,N_12096,N_12493);
xor U13041 (N_13041,N_12409,N_12365);
and U13042 (N_13042,N_12946,N_12099);
or U13043 (N_13043,N_12532,N_12555);
xnor U13044 (N_13044,N_12884,N_12940);
nand U13045 (N_13045,N_12943,N_12056);
or U13046 (N_13046,N_12624,N_12191);
and U13047 (N_13047,N_12569,N_12395);
or U13048 (N_13048,N_12179,N_12777);
or U13049 (N_13049,N_12595,N_12148);
nand U13050 (N_13050,N_12944,N_12927);
nand U13051 (N_13051,N_12935,N_12959);
nor U13052 (N_13052,N_12501,N_12931);
and U13053 (N_13053,N_12235,N_12170);
xor U13054 (N_13054,N_12016,N_12820);
nand U13055 (N_13055,N_12917,N_12489);
or U13056 (N_13056,N_12372,N_12774);
nor U13057 (N_13057,N_12967,N_12803);
or U13058 (N_13058,N_12411,N_12349);
and U13059 (N_13059,N_12323,N_12044);
xor U13060 (N_13060,N_12380,N_12523);
or U13061 (N_13061,N_12165,N_12760);
nand U13062 (N_13062,N_12080,N_12812);
nor U13063 (N_13063,N_12674,N_12512);
nor U13064 (N_13064,N_12619,N_12403);
or U13065 (N_13065,N_12111,N_12333);
xnor U13066 (N_13066,N_12620,N_12184);
xnor U13067 (N_13067,N_12526,N_12579);
xnor U13068 (N_13068,N_12542,N_12059);
nand U13069 (N_13069,N_12804,N_12926);
xnor U13070 (N_13070,N_12354,N_12299);
and U13071 (N_13071,N_12686,N_12280);
and U13072 (N_13072,N_12189,N_12706);
nand U13073 (N_13073,N_12055,N_12492);
nand U13074 (N_13074,N_12206,N_12618);
and U13075 (N_13075,N_12129,N_12535);
nand U13076 (N_13076,N_12734,N_12490);
and U13077 (N_13077,N_12767,N_12589);
xnor U13078 (N_13078,N_12090,N_12565);
and U13079 (N_13079,N_12219,N_12652);
and U13080 (N_13080,N_12656,N_12413);
nor U13081 (N_13081,N_12617,N_12320);
and U13082 (N_13082,N_12100,N_12695);
xor U13083 (N_13083,N_12780,N_12548);
nand U13084 (N_13084,N_12784,N_12061);
or U13085 (N_13085,N_12929,N_12525);
xnor U13086 (N_13086,N_12387,N_12054);
and U13087 (N_13087,N_12478,N_12420);
and U13088 (N_13088,N_12028,N_12045);
nand U13089 (N_13089,N_12288,N_12136);
nor U13090 (N_13090,N_12980,N_12400);
nand U13091 (N_13091,N_12228,N_12762);
and U13092 (N_13092,N_12861,N_12192);
and U13093 (N_13093,N_12601,N_12146);
nor U13094 (N_13094,N_12669,N_12266);
xnor U13095 (N_13095,N_12473,N_12176);
nand U13096 (N_13096,N_12401,N_12211);
nor U13097 (N_13097,N_12246,N_12270);
and U13098 (N_13098,N_12105,N_12441);
xor U13099 (N_13099,N_12704,N_12049);
or U13100 (N_13100,N_12564,N_12806);
nand U13101 (N_13101,N_12263,N_12729);
and U13102 (N_13102,N_12067,N_12360);
and U13103 (N_13103,N_12075,N_12672);
nor U13104 (N_13104,N_12000,N_12267);
and U13105 (N_13105,N_12494,N_12050);
and U13106 (N_13106,N_12924,N_12845);
or U13107 (N_13107,N_12212,N_12633);
or U13108 (N_13108,N_12974,N_12328);
nand U13109 (N_13109,N_12378,N_12871);
and U13110 (N_13110,N_12539,N_12121);
xnor U13111 (N_13111,N_12201,N_12417);
or U13112 (N_13112,N_12802,N_12433);
nand U13113 (N_13113,N_12261,N_12665);
or U13114 (N_13114,N_12113,N_12755);
xor U13115 (N_13115,N_12453,N_12025);
nor U13116 (N_13116,N_12163,N_12086);
nor U13117 (N_13117,N_12622,N_12107);
and U13118 (N_13118,N_12249,N_12868);
xor U13119 (N_13119,N_12483,N_12279);
nand U13120 (N_13120,N_12640,N_12870);
nand U13121 (N_13121,N_12007,N_12084);
and U13122 (N_13122,N_12688,N_12356);
nor U13123 (N_13123,N_12561,N_12697);
and U13124 (N_13124,N_12995,N_12603);
nand U13125 (N_13125,N_12230,N_12218);
or U13126 (N_13126,N_12382,N_12673);
xor U13127 (N_13127,N_12251,N_12447);
and U13128 (N_13128,N_12268,N_12787);
nor U13129 (N_13129,N_12725,N_12765);
nand U13130 (N_13130,N_12596,N_12104);
or U13131 (N_13131,N_12416,N_12352);
nand U13132 (N_13132,N_12541,N_12297);
xnor U13133 (N_13133,N_12322,N_12324);
and U13134 (N_13134,N_12809,N_12747);
and U13135 (N_13135,N_12215,N_12074);
and U13136 (N_13136,N_12456,N_12970);
or U13137 (N_13137,N_12602,N_12037);
or U13138 (N_13138,N_12318,N_12452);
xor U13139 (N_13139,N_12609,N_12728);
xnor U13140 (N_13140,N_12630,N_12936);
xnor U13141 (N_13141,N_12553,N_12437);
and U13142 (N_13142,N_12794,N_12002);
nand U13143 (N_13143,N_12782,N_12247);
nand U13144 (N_13144,N_12689,N_12125);
and U13145 (N_13145,N_12012,N_12766);
or U13146 (N_13146,N_12773,N_12758);
or U13147 (N_13147,N_12126,N_12530);
xnor U13148 (N_13148,N_12419,N_12465);
nor U13149 (N_13149,N_12240,N_12078);
nand U13150 (N_13150,N_12408,N_12987);
and U13151 (N_13151,N_12292,N_12149);
or U13152 (N_13152,N_12137,N_12114);
xnor U13153 (N_13153,N_12790,N_12432);
nand U13154 (N_13154,N_12415,N_12488);
nor U13155 (N_13155,N_12544,N_12879);
nor U13156 (N_13156,N_12637,N_12559);
nor U13157 (N_13157,N_12171,N_12402);
xnor U13158 (N_13158,N_12142,N_12497);
or U13159 (N_13159,N_12029,N_12344);
xor U13160 (N_13160,N_12981,N_12978);
nor U13161 (N_13161,N_12938,N_12883);
or U13162 (N_13162,N_12715,N_12200);
xor U13163 (N_13163,N_12072,N_12685);
xor U13164 (N_13164,N_12810,N_12046);
nor U13165 (N_13165,N_12899,N_12414);
and U13166 (N_13166,N_12710,N_12347);
or U13167 (N_13167,N_12626,N_12629);
and U13168 (N_13168,N_12157,N_12143);
or U13169 (N_13169,N_12881,N_12284);
nand U13170 (N_13170,N_12188,N_12664);
nand U13171 (N_13171,N_12952,N_12556);
nand U13172 (N_13172,N_12887,N_12009);
or U13173 (N_13173,N_12960,N_12731);
nand U13174 (N_13174,N_12031,N_12684);
nor U13175 (N_13175,N_12900,N_12203);
or U13176 (N_13176,N_12145,N_12262);
nor U13177 (N_13177,N_12771,N_12902);
xnor U13178 (N_13178,N_12832,N_12273);
xnor U13179 (N_13179,N_12193,N_12017);
nor U13180 (N_13180,N_12177,N_12600);
nand U13181 (N_13181,N_12425,N_12849);
nor U13182 (N_13182,N_12379,N_12885);
nor U13183 (N_13183,N_12321,N_12651);
or U13184 (N_13184,N_12957,N_12127);
nor U13185 (N_13185,N_12257,N_12566);
nand U13186 (N_13186,N_12448,N_12101);
xnor U13187 (N_13187,N_12001,N_12892);
and U13188 (N_13188,N_12457,N_12546);
xor U13189 (N_13189,N_12350,N_12828);
nand U13190 (N_13190,N_12300,N_12083);
xnor U13191 (N_13191,N_12999,N_12791);
xor U13192 (N_13192,N_12876,N_12648);
xnor U13193 (N_13193,N_12214,N_12663);
and U13194 (N_13194,N_12965,N_12516);
and U13195 (N_13195,N_12646,N_12032);
and U13196 (N_13196,N_12788,N_12997);
xor U13197 (N_13197,N_12576,N_12335);
nor U13198 (N_13198,N_12909,N_12314);
xnor U13199 (N_13199,N_12786,N_12196);
xor U13200 (N_13200,N_12968,N_12337);
and U13201 (N_13201,N_12131,N_12116);
xnor U13202 (N_13202,N_12181,N_12289);
or U13203 (N_13203,N_12973,N_12034);
nor U13204 (N_13204,N_12503,N_12446);
xor U13205 (N_13205,N_12154,N_12421);
xnor U13206 (N_13206,N_12854,N_12355);
nand U13207 (N_13207,N_12724,N_12963);
and U13208 (N_13208,N_12122,N_12843);
and U13209 (N_13209,N_12156,N_12644);
or U13210 (N_13210,N_12653,N_12740);
nand U13211 (N_13211,N_12258,N_12581);
xnor U13212 (N_13212,N_12655,N_12918);
nand U13213 (N_13213,N_12875,N_12703);
nor U13214 (N_13214,N_12366,N_12514);
xnor U13215 (N_13215,N_12475,N_12385);
and U13216 (N_13216,N_12159,N_12313);
or U13217 (N_13217,N_12920,N_12916);
or U13218 (N_13218,N_12937,N_12814);
and U13219 (N_13219,N_12496,N_12811);
nor U13220 (N_13220,N_12066,N_12334);
nand U13221 (N_13221,N_12781,N_12255);
or U13222 (N_13222,N_12397,N_12151);
or U13223 (N_13223,N_12594,N_12799);
and U13224 (N_13224,N_12574,N_12407);
nand U13225 (N_13225,N_12969,N_12161);
nor U13226 (N_13226,N_12947,N_12241);
nand U13227 (N_13227,N_12058,N_12932);
nand U13228 (N_13228,N_12634,N_12702);
or U13229 (N_13229,N_12460,N_12088);
and U13230 (N_13230,N_12616,N_12837);
xor U13231 (N_13231,N_12907,N_12911);
nor U13232 (N_13232,N_12815,N_12979);
nor U13233 (N_13233,N_12705,N_12426);
nand U13234 (N_13234,N_12117,N_12676);
or U13235 (N_13235,N_12223,N_12976);
xor U13236 (N_13236,N_12357,N_12307);
or U13237 (N_13237,N_12950,N_12586);
or U13238 (N_13238,N_12166,N_12836);
and U13239 (N_13239,N_12035,N_12245);
or U13240 (N_13240,N_12021,N_12906);
xor U13241 (N_13241,N_12775,N_12921);
or U13242 (N_13242,N_12558,N_12521);
xnor U13243 (N_13243,N_12855,N_12238);
or U13244 (N_13244,N_12042,N_12041);
nand U13245 (N_13245,N_12233,N_12750);
nor U13246 (N_13246,N_12123,N_12632);
nand U13247 (N_13247,N_12610,N_12390);
or U13248 (N_13248,N_12312,N_12461);
nand U13249 (N_13249,N_12714,N_12467);
nand U13250 (N_13250,N_12560,N_12852);
nor U13251 (N_13251,N_12063,N_12485);
nor U13252 (N_13252,N_12252,N_12278);
xnor U13253 (N_13253,N_12643,N_12642);
nand U13254 (N_13254,N_12197,N_12018);
xor U13255 (N_13255,N_12185,N_12482);
or U13256 (N_13256,N_12679,N_12573);
or U13257 (N_13257,N_12040,N_12259);
or U13258 (N_13258,N_12449,N_12737);
nand U13259 (N_13259,N_12631,N_12670);
and U13260 (N_13260,N_12800,N_12770);
xor U13261 (N_13261,N_12339,N_12680);
nor U13262 (N_13262,N_12256,N_12666);
nand U13263 (N_13263,N_12645,N_12627);
nor U13264 (N_13264,N_12949,N_12282);
nor U13265 (N_13265,N_12612,N_12598);
and U13266 (N_13266,N_12795,N_12391);
and U13267 (N_13267,N_12826,N_12897);
and U13268 (N_13268,N_12047,N_12423);
or U13269 (N_13269,N_12721,N_12692);
xor U13270 (N_13270,N_12316,N_12701);
nand U13271 (N_13271,N_12716,N_12509);
or U13272 (N_13272,N_12112,N_12353);
and U13273 (N_13273,N_12250,N_12660);
nand U13274 (N_13274,N_12412,N_12368);
and U13275 (N_13275,N_12277,N_12343);
xnor U13276 (N_13276,N_12903,N_12169);
or U13277 (N_13277,N_12462,N_12662);
nor U13278 (N_13278,N_12108,N_12829);
or U13279 (N_13279,N_12427,N_12797);
nand U13280 (N_13280,N_12739,N_12636);
xor U13281 (N_13281,N_12607,N_12064);
and U13282 (N_13282,N_12399,N_12585);
nand U13283 (N_13283,N_12719,N_12529);
and U13284 (N_13284,N_12635,N_12118);
nor U13285 (N_13285,N_12792,N_12371);
nand U13286 (N_13286,N_12264,N_12003);
or U13287 (N_13287,N_12272,N_12168);
nand U13288 (N_13288,N_12153,N_12827);
and U13289 (N_13289,N_12180,N_12778);
or U13290 (N_13290,N_12650,N_12134);
nand U13291 (N_13291,N_12182,N_12869);
xnor U13292 (N_13292,N_12087,N_12071);
nand U13293 (N_13293,N_12373,N_12451);
nand U13294 (N_13294,N_12377,N_12860);
or U13295 (N_13295,N_12691,N_12428);
or U13296 (N_13296,N_12597,N_12076);
and U13297 (N_13297,N_12638,N_12540);
nor U13298 (N_13298,N_12986,N_12948);
nand U13299 (N_13299,N_12178,N_12835);
nor U13300 (N_13300,N_12236,N_12498);
and U13301 (N_13301,N_12690,N_12914);
or U13302 (N_13302,N_12841,N_12092);
nor U13303 (N_13303,N_12455,N_12367);
and U13304 (N_13304,N_12536,N_12346);
or U13305 (N_13305,N_12510,N_12269);
nand U13306 (N_13306,N_12232,N_12880);
or U13307 (N_13307,N_12393,N_12848);
nand U13308 (N_13308,N_12422,N_12039);
or U13309 (N_13309,N_12730,N_12531);
nand U13310 (N_13310,N_12202,N_12386);
nor U13311 (N_13311,N_12306,N_12374);
or U13312 (N_13312,N_12102,N_12013);
and U13313 (N_13313,N_12103,N_12291);
or U13314 (N_13314,N_12410,N_12647);
or U13315 (N_13315,N_12294,N_12759);
xnor U13316 (N_13316,N_12060,N_12798);
xor U13317 (N_13317,N_12351,N_12972);
and U13318 (N_13318,N_12015,N_12989);
xor U13319 (N_13319,N_12712,N_12991);
and U13320 (N_13320,N_12913,N_12557);
nor U13321 (N_13321,N_12332,N_12939);
and U13322 (N_13322,N_12951,N_12085);
xnor U13323 (N_13323,N_12376,N_12783);
nor U13324 (N_13324,N_12851,N_12824);
or U13325 (N_13325,N_12744,N_12274);
nor U13326 (N_13326,N_12604,N_12813);
nor U13327 (N_13327,N_12183,N_12834);
nand U13328 (N_13328,N_12793,N_12150);
xor U13329 (N_13329,N_12051,N_12155);
and U13330 (N_13330,N_12808,N_12639);
xnor U13331 (N_13331,N_12990,N_12859);
nor U13332 (N_13332,N_12174,N_12005);
nand U13333 (N_13333,N_12375,N_12445);
nand U13334 (N_13334,N_12713,N_12024);
nand U13335 (N_13335,N_12052,N_12020);
and U13336 (N_13336,N_12271,N_12026);
xor U13337 (N_13337,N_12850,N_12934);
or U13338 (N_13338,N_12296,N_12693);
and U13339 (N_13339,N_12905,N_12006);
and U13340 (N_13340,N_12550,N_12727);
nand U13341 (N_13341,N_12732,N_12533);
and U13342 (N_13342,N_12507,N_12895);
xnor U13343 (N_13343,N_12668,N_12234);
xor U13344 (N_13344,N_12801,N_12825);
and U13345 (N_13345,N_12216,N_12140);
nand U13346 (N_13346,N_12500,N_12866);
nand U13347 (N_13347,N_12471,N_12303);
and U13348 (N_13348,N_12361,N_12160);
nor U13349 (N_13349,N_12450,N_12817);
nand U13350 (N_13350,N_12502,N_12839);
and U13351 (N_13351,N_12327,N_12204);
xnor U13352 (N_13352,N_12130,N_12383);
nand U13353 (N_13353,N_12095,N_12923);
and U13354 (N_13354,N_12305,N_12022);
nand U13355 (N_13355,N_12298,N_12776);
or U13356 (N_13356,N_12889,N_12276);
and U13357 (N_13357,N_12865,N_12756);
xor U13358 (N_13358,N_12504,N_12173);
or U13359 (N_13359,N_12745,N_12062);
and U13360 (N_13360,N_12853,N_12772);
or U13361 (N_13361,N_12534,N_12658);
or U13362 (N_13362,N_12519,N_12443);
nor U13363 (N_13363,N_12207,N_12115);
xnor U13364 (N_13364,N_12043,N_12389);
nand U13365 (N_13365,N_12198,N_12033);
nand U13366 (N_13366,N_12070,N_12682);
xnor U13367 (N_13367,N_12910,N_12833);
nand U13368 (N_13368,N_12831,N_12983);
and U13369 (N_13369,N_12124,N_12468);
xor U13370 (N_13370,N_12733,N_12789);
xnor U13371 (N_13371,N_12928,N_12439);
and U13372 (N_13372,N_12992,N_12711);
or U13373 (N_13373,N_12606,N_12081);
or U13374 (N_13374,N_12898,N_12515);
nand U13375 (N_13375,N_12707,N_12217);
and U13376 (N_13376,N_12890,N_12821);
nand U13377 (N_13377,N_12567,N_12764);
nand U13378 (N_13378,N_12369,N_12547);
nor U13379 (N_13379,N_12144,N_12877);
and U13380 (N_13380,N_12649,N_12552);
or U13381 (N_13381,N_12491,N_12286);
or U13382 (N_13382,N_12364,N_12753);
or U13383 (N_13383,N_12743,N_12454);
nor U13384 (N_13384,N_12641,N_12011);
xor U13385 (N_13385,N_12466,N_12132);
xor U13386 (N_13386,N_12867,N_12093);
or U13387 (N_13387,N_12977,N_12210);
nor U13388 (N_13388,N_12678,N_12242);
nand U13389 (N_13389,N_12370,N_12838);
nor U13390 (N_13390,N_12430,N_12681);
xnor U13391 (N_13391,N_12147,N_12757);
and U13392 (N_13392,N_12605,N_12694);
nor U13393 (N_13393,N_12287,N_12481);
xnor U13394 (N_13394,N_12396,N_12543);
and U13395 (N_13395,N_12738,N_12901);
nand U13396 (N_13396,N_12985,N_12438);
nor U13397 (N_13397,N_12508,N_12139);
or U13398 (N_13398,N_12763,N_12819);
nor U13399 (N_13399,N_12700,N_12120);
and U13400 (N_13400,N_12338,N_12283);
nand U13401 (N_13401,N_12164,N_12822);
or U13402 (N_13402,N_12384,N_12621);
nand U13403 (N_13403,N_12073,N_12709);
or U13404 (N_13404,N_12551,N_12231);
xnor U13405 (N_13405,N_12440,N_12254);
nor U13406 (N_13406,N_12696,N_12392);
or U13407 (N_13407,N_12030,N_12479);
nor U13408 (N_13408,N_12578,N_12590);
or U13409 (N_13409,N_12027,N_12019);
or U13410 (N_13410,N_12718,N_12253);
xnor U13411 (N_13411,N_12608,N_12818);
xnor U13412 (N_13412,N_12097,N_12677);
or U13413 (N_13413,N_12583,N_12227);
xnor U13414 (N_13414,N_12708,N_12675);
xnor U13415 (N_13415,N_12434,N_12614);
or U13416 (N_13416,N_12243,N_12625);
nor U13417 (N_13417,N_12752,N_12476);
nand U13418 (N_13418,N_12128,N_12563);
or U13419 (N_13419,N_12888,N_12082);
nand U13420 (N_13420,N_12069,N_12904);
or U13421 (N_13421,N_12194,N_12119);
nand U13422 (N_13422,N_12175,N_12199);
xor U13423 (N_13423,N_12687,N_12919);
and U13424 (N_13424,N_12768,N_12698);
nand U13425 (N_13425,N_12167,N_12599);
or U13426 (N_13426,N_12331,N_12110);
or U13427 (N_13427,N_12133,N_12435);
xnor U13428 (N_13428,N_12477,N_12065);
nand U13429 (N_13429,N_12954,N_12470);
or U13430 (N_13430,N_12748,N_12319);
nand U13431 (N_13431,N_12345,N_12513);
nor U13432 (N_13432,N_12295,N_12796);
or U13433 (N_13433,N_12518,N_12761);
nand U13434 (N_13434,N_12571,N_12722);
nand U13435 (N_13435,N_12244,N_12874);
xnor U13436 (N_13436,N_12141,N_12816);
xnor U13437 (N_13437,N_12077,N_12863);
xnor U13438 (N_13438,N_12330,N_12442);
nor U13439 (N_13439,N_12398,N_12158);
nand U13440 (N_13440,N_12329,N_12864);
xor U13441 (N_13441,N_12186,N_12010);
and U13442 (N_13442,N_12925,N_12358);
nand U13443 (N_13443,N_12857,N_12588);
and U13444 (N_13444,N_12098,N_12915);
nand U13445 (N_13445,N_12464,N_12538);
nand U13446 (N_13446,N_12961,N_12205);
and U13447 (N_13447,N_12873,N_12237);
nand U13448 (N_13448,N_12956,N_12779);
nand U13449 (N_13449,N_12592,N_12615);
xnor U13450 (N_13450,N_12661,N_12953);
nand U13451 (N_13451,N_12580,N_12893);
nor U13452 (N_13452,N_12436,N_12671);
nor U13453 (N_13453,N_12315,N_12469);
nand U13454 (N_13454,N_12611,N_12746);
xor U13455 (N_13455,N_12302,N_12213);
or U13456 (N_13456,N_12517,N_12933);
xor U13457 (N_13457,N_12458,N_12741);
nor U13458 (N_13458,N_12699,N_12856);
nand U13459 (N_13459,N_12388,N_12844);
xor U13460 (N_13460,N_12742,N_12089);
nand U13461 (N_13461,N_12285,N_12424);
nor U13462 (N_13462,N_12720,N_12221);
nor U13463 (N_13463,N_12505,N_12404);
nand U13464 (N_13464,N_12971,N_12362);
nor U13465 (N_13465,N_12265,N_12922);
nor U13466 (N_13466,N_12209,N_12570);
nor U13467 (N_13467,N_12785,N_12735);
and U13468 (N_13468,N_12657,N_12348);
or U13469 (N_13469,N_12038,N_12996);
nor U13470 (N_13470,N_12053,N_12472);
nand U13471 (N_13471,N_12394,N_12336);
nor U13472 (N_13472,N_12281,N_12805);
and U13473 (N_13473,N_12659,N_12222);
nand U13474 (N_13474,N_12109,N_12463);
nand U13475 (N_13475,N_12549,N_12226);
nand U13476 (N_13476,N_12187,N_12004);
xor U13477 (N_13477,N_12754,N_12807);
and U13478 (N_13478,N_12554,N_12872);
xnor U13479 (N_13479,N_12955,N_12993);
xor U13480 (N_13480,N_12152,N_12474);
nor U13481 (N_13481,N_12275,N_12309);
nor U13482 (N_13482,N_12723,N_12260);
or U13483 (N_13483,N_12572,N_12363);
nand U13484 (N_13484,N_12858,N_12683);
nor U13485 (N_13485,N_12239,N_12941);
xor U13486 (N_13486,N_12301,N_12769);
and U13487 (N_13487,N_12310,N_12487);
nor U13488 (N_13488,N_12359,N_12418);
nor U13489 (N_13489,N_12994,N_12524);
and U13490 (N_13490,N_12896,N_12613);
or U13491 (N_13491,N_12317,N_12429);
nand U13492 (N_13492,N_12942,N_12628);
nand U13493 (N_13493,N_12290,N_12406);
nor U13494 (N_13494,N_12726,N_12847);
and U13495 (N_13495,N_12545,N_12966);
nand U13496 (N_13496,N_12751,N_12225);
nand U13497 (N_13497,N_12958,N_12568);
xnor U13498 (N_13498,N_12381,N_12862);
or U13499 (N_13499,N_12846,N_12248);
xnor U13500 (N_13500,N_12437,N_12245);
nor U13501 (N_13501,N_12114,N_12633);
nand U13502 (N_13502,N_12656,N_12519);
nand U13503 (N_13503,N_12328,N_12088);
xnor U13504 (N_13504,N_12109,N_12046);
nor U13505 (N_13505,N_12389,N_12599);
nand U13506 (N_13506,N_12923,N_12345);
xor U13507 (N_13507,N_12436,N_12499);
nand U13508 (N_13508,N_12139,N_12296);
xnor U13509 (N_13509,N_12845,N_12770);
nor U13510 (N_13510,N_12857,N_12957);
nand U13511 (N_13511,N_12020,N_12992);
or U13512 (N_13512,N_12148,N_12937);
or U13513 (N_13513,N_12492,N_12834);
and U13514 (N_13514,N_12728,N_12355);
nand U13515 (N_13515,N_12441,N_12910);
xor U13516 (N_13516,N_12326,N_12426);
or U13517 (N_13517,N_12290,N_12309);
xnor U13518 (N_13518,N_12509,N_12815);
or U13519 (N_13519,N_12951,N_12967);
nand U13520 (N_13520,N_12875,N_12770);
xnor U13521 (N_13521,N_12496,N_12745);
or U13522 (N_13522,N_12031,N_12461);
nor U13523 (N_13523,N_12044,N_12157);
xnor U13524 (N_13524,N_12199,N_12111);
or U13525 (N_13525,N_12145,N_12326);
nand U13526 (N_13526,N_12822,N_12416);
and U13527 (N_13527,N_12431,N_12933);
xnor U13528 (N_13528,N_12334,N_12710);
xnor U13529 (N_13529,N_12926,N_12158);
nand U13530 (N_13530,N_12205,N_12822);
and U13531 (N_13531,N_12101,N_12105);
nand U13532 (N_13532,N_12732,N_12738);
nor U13533 (N_13533,N_12021,N_12306);
xor U13534 (N_13534,N_12415,N_12963);
and U13535 (N_13535,N_12942,N_12175);
xor U13536 (N_13536,N_12616,N_12330);
nor U13537 (N_13537,N_12352,N_12327);
nor U13538 (N_13538,N_12622,N_12856);
and U13539 (N_13539,N_12843,N_12368);
xor U13540 (N_13540,N_12081,N_12544);
and U13541 (N_13541,N_12686,N_12896);
and U13542 (N_13542,N_12823,N_12523);
nor U13543 (N_13543,N_12762,N_12875);
xor U13544 (N_13544,N_12149,N_12818);
nand U13545 (N_13545,N_12336,N_12014);
xnor U13546 (N_13546,N_12742,N_12849);
xor U13547 (N_13547,N_12947,N_12651);
or U13548 (N_13548,N_12247,N_12085);
nand U13549 (N_13549,N_12747,N_12426);
or U13550 (N_13550,N_12922,N_12399);
xnor U13551 (N_13551,N_12110,N_12957);
and U13552 (N_13552,N_12664,N_12155);
xnor U13553 (N_13553,N_12141,N_12835);
or U13554 (N_13554,N_12093,N_12525);
xor U13555 (N_13555,N_12211,N_12361);
nand U13556 (N_13556,N_12957,N_12872);
or U13557 (N_13557,N_12712,N_12033);
and U13558 (N_13558,N_12388,N_12990);
nor U13559 (N_13559,N_12886,N_12791);
nand U13560 (N_13560,N_12461,N_12455);
and U13561 (N_13561,N_12592,N_12491);
and U13562 (N_13562,N_12636,N_12357);
xnor U13563 (N_13563,N_12900,N_12583);
or U13564 (N_13564,N_12250,N_12229);
and U13565 (N_13565,N_12988,N_12771);
nand U13566 (N_13566,N_12000,N_12090);
nand U13567 (N_13567,N_12470,N_12547);
or U13568 (N_13568,N_12643,N_12312);
or U13569 (N_13569,N_12947,N_12890);
xnor U13570 (N_13570,N_12599,N_12764);
nand U13571 (N_13571,N_12427,N_12438);
or U13572 (N_13572,N_12069,N_12228);
and U13573 (N_13573,N_12415,N_12533);
nand U13574 (N_13574,N_12789,N_12615);
or U13575 (N_13575,N_12574,N_12831);
or U13576 (N_13576,N_12165,N_12775);
or U13577 (N_13577,N_12150,N_12248);
nand U13578 (N_13578,N_12163,N_12065);
nor U13579 (N_13579,N_12937,N_12000);
and U13580 (N_13580,N_12439,N_12413);
nand U13581 (N_13581,N_12932,N_12616);
and U13582 (N_13582,N_12877,N_12517);
and U13583 (N_13583,N_12348,N_12235);
and U13584 (N_13584,N_12712,N_12212);
xnor U13585 (N_13585,N_12971,N_12475);
and U13586 (N_13586,N_12427,N_12981);
nor U13587 (N_13587,N_12715,N_12568);
and U13588 (N_13588,N_12021,N_12628);
or U13589 (N_13589,N_12336,N_12943);
nand U13590 (N_13590,N_12544,N_12385);
and U13591 (N_13591,N_12313,N_12257);
nand U13592 (N_13592,N_12488,N_12301);
and U13593 (N_13593,N_12293,N_12728);
or U13594 (N_13594,N_12992,N_12759);
nor U13595 (N_13595,N_12635,N_12647);
or U13596 (N_13596,N_12702,N_12095);
nand U13597 (N_13597,N_12516,N_12808);
or U13598 (N_13598,N_12864,N_12787);
and U13599 (N_13599,N_12657,N_12859);
and U13600 (N_13600,N_12212,N_12640);
or U13601 (N_13601,N_12177,N_12527);
nand U13602 (N_13602,N_12312,N_12754);
nor U13603 (N_13603,N_12255,N_12319);
nor U13604 (N_13604,N_12912,N_12431);
and U13605 (N_13605,N_12312,N_12651);
xnor U13606 (N_13606,N_12911,N_12938);
nand U13607 (N_13607,N_12266,N_12430);
xnor U13608 (N_13608,N_12997,N_12727);
or U13609 (N_13609,N_12847,N_12371);
xnor U13610 (N_13610,N_12776,N_12399);
nor U13611 (N_13611,N_12649,N_12806);
and U13612 (N_13612,N_12793,N_12435);
xor U13613 (N_13613,N_12958,N_12699);
nor U13614 (N_13614,N_12170,N_12518);
or U13615 (N_13615,N_12784,N_12977);
nand U13616 (N_13616,N_12791,N_12695);
and U13617 (N_13617,N_12356,N_12593);
or U13618 (N_13618,N_12991,N_12797);
and U13619 (N_13619,N_12112,N_12021);
and U13620 (N_13620,N_12191,N_12508);
xnor U13621 (N_13621,N_12168,N_12353);
and U13622 (N_13622,N_12883,N_12421);
or U13623 (N_13623,N_12768,N_12914);
and U13624 (N_13624,N_12689,N_12183);
nor U13625 (N_13625,N_12547,N_12219);
nor U13626 (N_13626,N_12477,N_12200);
xnor U13627 (N_13627,N_12682,N_12520);
nand U13628 (N_13628,N_12539,N_12486);
or U13629 (N_13629,N_12360,N_12001);
or U13630 (N_13630,N_12198,N_12505);
or U13631 (N_13631,N_12956,N_12415);
xor U13632 (N_13632,N_12418,N_12406);
xnor U13633 (N_13633,N_12924,N_12824);
xor U13634 (N_13634,N_12163,N_12997);
or U13635 (N_13635,N_12660,N_12750);
and U13636 (N_13636,N_12117,N_12562);
and U13637 (N_13637,N_12180,N_12687);
nand U13638 (N_13638,N_12302,N_12938);
and U13639 (N_13639,N_12923,N_12211);
nand U13640 (N_13640,N_12454,N_12605);
nor U13641 (N_13641,N_12380,N_12929);
or U13642 (N_13642,N_12614,N_12241);
or U13643 (N_13643,N_12606,N_12608);
or U13644 (N_13644,N_12671,N_12154);
or U13645 (N_13645,N_12554,N_12348);
and U13646 (N_13646,N_12030,N_12607);
or U13647 (N_13647,N_12146,N_12875);
nor U13648 (N_13648,N_12721,N_12020);
xnor U13649 (N_13649,N_12811,N_12825);
nand U13650 (N_13650,N_12783,N_12265);
xor U13651 (N_13651,N_12205,N_12458);
nor U13652 (N_13652,N_12704,N_12311);
and U13653 (N_13653,N_12492,N_12835);
nand U13654 (N_13654,N_12357,N_12160);
xor U13655 (N_13655,N_12345,N_12867);
nand U13656 (N_13656,N_12541,N_12923);
xnor U13657 (N_13657,N_12293,N_12497);
xnor U13658 (N_13658,N_12601,N_12426);
nand U13659 (N_13659,N_12005,N_12866);
or U13660 (N_13660,N_12280,N_12185);
nand U13661 (N_13661,N_12897,N_12508);
xor U13662 (N_13662,N_12556,N_12962);
and U13663 (N_13663,N_12951,N_12546);
or U13664 (N_13664,N_12922,N_12798);
and U13665 (N_13665,N_12368,N_12479);
nand U13666 (N_13666,N_12505,N_12572);
xnor U13667 (N_13667,N_12720,N_12649);
or U13668 (N_13668,N_12745,N_12608);
and U13669 (N_13669,N_12494,N_12314);
xor U13670 (N_13670,N_12884,N_12426);
nor U13671 (N_13671,N_12513,N_12480);
nor U13672 (N_13672,N_12118,N_12100);
nor U13673 (N_13673,N_12197,N_12191);
nor U13674 (N_13674,N_12626,N_12681);
nand U13675 (N_13675,N_12922,N_12611);
nand U13676 (N_13676,N_12933,N_12507);
nor U13677 (N_13677,N_12689,N_12487);
or U13678 (N_13678,N_12397,N_12536);
nand U13679 (N_13679,N_12515,N_12476);
nand U13680 (N_13680,N_12639,N_12457);
or U13681 (N_13681,N_12066,N_12397);
nor U13682 (N_13682,N_12887,N_12380);
and U13683 (N_13683,N_12886,N_12019);
or U13684 (N_13684,N_12119,N_12023);
or U13685 (N_13685,N_12912,N_12767);
nand U13686 (N_13686,N_12764,N_12993);
xor U13687 (N_13687,N_12634,N_12493);
nand U13688 (N_13688,N_12431,N_12118);
or U13689 (N_13689,N_12401,N_12531);
nor U13690 (N_13690,N_12217,N_12539);
nor U13691 (N_13691,N_12220,N_12883);
or U13692 (N_13692,N_12922,N_12449);
and U13693 (N_13693,N_12704,N_12426);
nor U13694 (N_13694,N_12897,N_12645);
nand U13695 (N_13695,N_12519,N_12288);
and U13696 (N_13696,N_12703,N_12245);
xnor U13697 (N_13697,N_12028,N_12844);
nor U13698 (N_13698,N_12912,N_12525);
or U13699 (N_13699,N_12888,N_12101);
or U13700 (N_13700,N_12501,N_12198);
or U13701 (N_13701,N_12990,N_12017);
or U13702 (N_13702,N_12862,N_12166);
or U13703 (N_13703,N_12639,N_12456);
xor U13704 (N_13704,N_12772,N_12846);
nand U13705 (N_13705,N_12176,N_12742);
and U13706 (N_13706,N_12424,N_12316);
or U13707 (N_13707,N_12209,N_12783);
nand U13708 (N_13708,N_12464,N_12282);
xnor U13709 (N_13709,N_12817,N_12760);
and U13710 (N_13710,N_12959,N_12848);
nand U13711 (N_13711,N_12856,N_12799);
or U13712 (N_13712,N_12988,N_12232);
xnor U13713 (N_13713,N_12097,N_12740);
and U13714 (N_13714,N_12006,N_12981);
nor U13715 (N_13715,N_12733,N_12359);
and U13716 (N_13716,N_12822,N_12706);
xnor U13717 (N_13717,N_12677,N_12610);
xor U13718 (N_13718,N_12269,N_12126);
nor U13719 (N_13719,N_12467,N_12772);
or U13720 (N_13720,N_12436,N_12869);
nor U13721 (N_13721,N_12561,N_12260);
nor U13722 (N_13722,N_12201,N_12476);
nand U13723 (N_13723,N_12997,N_12968);
and U13724 (N_13724,N_12881,N_12907);
and U13725 (N_13725,N_12314,N_12881);
xnor U13726 (N_13726,N_12382,N_12889);
and U13727 (N_13727,N_12293,N_12147);
xor U13728 (N_13728,N_12342,N_12058);
or U13729 (N_13729,N_12771,N_12607);
and U13730 (N_13730,N_12072,N_12090);
nor U13731 (N_13731,N_12643,N_12273);
nor U13732 (N_13732,N_12567,N_12989);
nor U13733 (N_13733,N_12940,N_12475);
and U13734 (N_13734,N_12515,N_12383);
or U13735 (N_13735,N_12731,N_12188);
nor U13736 (N_13736,N_12317,N_12299);
nor U13737 (N_13737,N_12854,N_12052);
xor U13738 (N_13738,N_12688,N_12477);
or U13739 (N_13739,N_12419,N_12744);
nor U13740 (N_13740,N_12293,N_12357);
nand U13741 (N_13741,N_12239,N_12925);
or U13742 (N_13742,N_12186,N_12857);
and U13743 (N_13743,N_12907,N_12695);
xor U13744 (N_13744,N_12968,N_12378);
xor U13745 (N_13745,N_12598,N_12646);
nand U13746 (N_13746,N_12797,N_12595);
or U13747 (N_13747,N_12938,N_12080);
or U13748 (N_13748,N_12585,N_12495);
nand U13749 (N_13749,N_12246,N_12068);
or U13750 (N_13750,N_12272,N_12562);
xor U13751 (N_13751,N_12586,N_12462);
or U13752 (N_13752,N_12387,N_12281);
nor U13753 (N_13753,N_12644,N_12741);
and U13754 (N_13754,N_12367,N_12226);
and U13755 (N_13755,N_12338,N_12825);
xor U13756 (N_13756,N_12632,N_12594);
nand U13757 (N_13757,N_12938,N_12701);
xnor U13758 (N_13758,N_12855,N_12766);
nor U13759 (N_13759,N_12973,N_12403);
or U13760 (N_13760,N_12091,N_12414);
or U13761 (N_13761,N_12797,N_12872);
xnor U13762 (N_13762,N_12769,N_12128);
xor U13763 (N_13763,N_12240,N_12397);
and U13764 (N_13764,N_12731,N_12686);
nand U13765 (N_13765,N_12302,N_12379);
xor U13766 (N_13766,N_12891,N_12504);
nand U13767 (N_13767,N_12092,N_12426);
xor U13768 (N_13768,N_12594,N_12961);
or U13769 (N_13769,N_12679,N_12596);
nand U13770 (N_13770,N_12637,N_12828);
nand U13771 (N_13771,N_12874,N_12336);
xor U13772 (N_13772,N_12518,N_12031);
or U13773 (N_13773,N_12236,N_12750);
or U13774 (N_13774,N_12573,N_12447);
or U13775 (N_13775,N_12804,N_12399);
nor U13776 (N_13776,N_12455,N_12597);
xnor U13777 (N_13777,N_12504,N_12612);
nand U13778 (N_13778,N_12728,N_12619);
nand U13779 (N_13779,N_12596,N_12964);
nand U13780 (N_13780,N_12284,N_12253);
nand U13781 (N_13781,N_12628,N_12018);
and U13782 (N_13782,N_12656,N_12165);
nor U13783 (N_13783,N_12884,N_12798);
nand U13784 (N_13784,N_12436,N_12891);
nor U13785 (N_13785,N_12752,N_12616);
nand U13786 (N_13786,N_12569,N_12521);
or U13787 (N_13787,N_12576,N_12344);
and U13788 (N_13788,N_12706,N_12048);
and U13789 (N_13789,N_12099,N_12416);
or U13790 (N_13790,N_12614,N_12570);
xor U13791 (N_13791,N_12188,N_12528);
nor U13792 (N_13792,N_12346,N_12495);
or U13793 (N_13793,N_12602,N_12909);
nand U13794 (N_13794,N_12117,N_12535);
nand U13795 (N_13795,N_12058,N_12999);
or U13796 (N_13796,N_12431,N_12227);
or U13797 (N_13797,N_12159,N_12697);
xor U13798 (N_13798,N_12554,N_12989);
or U13799 (N_13799,N_12481,N_12118);
nand U13800 (N_13800,N_12130,N_12497);
xor U13801 (N_13801,N_12348,N_12588);
nor U13802 (N_13802,N_12499,N_12770);
nand U13803 (N_13803,N_12816,N_12673);
nor U13804 (N_13804,N_12035,N_12622);
and U13805 (N_13805,N_12063,N_12266);
nor U13806 (N_13806,N_12213,N_12217);
nor U13807 (N_13807,N_12919,N_12429);
xnor U13808 (N_13808,N_12111,N_12531);
xor U13809 (N_13809,N_12759,N_12997);
or U13810 (N_13810,N_12280,N_12077);
or U13811 (N_13811,N_12204,N_12334);
and U13812 (N_13812,N_12289,N_12648);
xnor U13813 (N_13813,N_12142,N_12695);
and U13814 (N_13814,N_12961,N_12308);
xnor U13815 (N_13815,N_12514,N_12404);
and U13816 (N_13816,N_12513,N_12397);
or U13817 (N_13817,N_12986,N_12908);
nand U13818 (N_13818,N_12217,N_12887);
or U13819 (N_13819,N_12311,N_12309);
nor U13820 (N_13820,N_12923,N_12505);
xnor U13821 (N_13821,N_12818,N_12708);
nand U13822 (N_13822,N_12503,N_12079);
xnor U13823 (N_13823,N_12745,N_12399);
xnor U13824 (N_13824,N_12443,N_12525);
xor U13825 (N_13825,N_12512,N_12154);
xnor U13826 (N_13826,N_12581,N_12887);
nand U13827 (N_13827,N_12491,N_12818);
xor U13828 (N_13828,N_12568,N_12066);
or U13829 (N_13829,N_12536,N_12983);
or U13830 (N_13830,N_12710,N_12098);
xor U13831 (N_13831,N_12208,N_12448);
and U13832 (N_13832,N_12569,N_12720);
or U13833 (N_13833,N_12293,N_12259);
nand U13834 (N_13834,N_12237,N_12298);
nand U13835 (N_13835,N_12731,N_12790);
or U13836 (N_13836,N_12301,N_12095);
and U13837 (N_13837,N_12452,N_12769);
or U13838 (N_13838,N_12652,N_12004);
xor U13839 (N_13839,N_12771,N_12166);
or U13840 (N_13840,N_12263,N_12044);
nor U13841 (N_13841,N_12660,N_12162);
or U13842 (N_13842,N_12409,N_12306);
nor U13843 (N_13843,N_12696,N_12306);
xor U13844 (N_13844,N_12417,N_12931);
nor U13845 (N_13845,N_12806,N_12959);
nand U13846 (N_13846,N_12085,N_12506);
nand U13847 (N_13847,N_12367,N_12646);
and U13848 (N_13848,N_12874,N_12026);
or U13849 (N_13849,N_12747,N_12471);
xor U13850 (N_13850,N_12456,N_12459);
nand U13851 (N_13851,N_12903,N_12257);
nor U13852 (N_13852,N_12334,N_12873);
nor U13853 (N_13853,N_12407,N_12488);
or U13854 (N_13854,N_12814,N_12754);
or U13855 (N_13855,N_12486,N_12204);
nand U13856 (N_13856,N_12472,N_12841);
nor U13857 (N_13857,N_12933,N_12293);
and U13858 (N_13858,N_12265,N_12043);
and U13859 (N_13859,N_12814,N_12620);
or U13860 (N_13860,N_12555,N_12172);
and U13861 (N_13861,N_12590,N_12153);
and U13862 (N_13862,N_12163,N_12614);
nand U13863 (N_13863,N_12561,N_12273);
nor U13864 (N_13864,N_12552,N_12724);
and U13865 (N_13865,N_12674,N_12166);
nand U13866 (N_13866,N_12240,N_12675);
xor U13867 (N_13867,N_12421,N_12981);
nor U13868 (N_13868,N_12550,N_12356);
xor U13869 (N_13869,N_12127,N_12069);
xnor U13870 (N_13870,N_12069,N_12213);
nand U13871 (N_13871,N_12691,N_12284);
nor U13872 (N_13872,N_12426,N_12032);
nor U13873 (N_13873,N_12425,N_12463);
or U13874 (N_13874,N_12189,N_12598);
nand U13875 (N_13875,N_12288,N_12212);
xnor U13876 (N_13876,N_12466,N_12488);
nand U13877 (N_13877,N_12166,N_12877);
or U13878 (N_13878,N_12772,N_12272);
or U13879 (N_13879,N_12746,N_12124);
nand U13880 (N_13880,N_12932,N_12477);
and U13881 (N_13881,N_12077,N_12261);
or U13882 (N_13882,N_12714,N_12411);
nor U13883 (N_13883,N_12748,N_12006);
and U13884 (N_13884,N_12234,N_12534);
or U13885 (N_13885,N_12346,N_12829);
nor U13886 (N_13886,N_12292,N_12010);
or U13887 (N_13887,N_12786,N_12784);
xnor U13888 (N_13888,N_12122,N_12461);
nand U13889 (N_13889,N_12597,N_12133);
and U13890 (N_13890,N_12845,N_12081);
nor U13891 (N_13891,N_12251,N_12226);
nor U13892 (N_13892,N_12155,N_12093);
nand U13893 (N_13893,N_12778,N_12873);
nor U13894 (N_13894,N_12095,N_12650);
and U13895 (N_13895,N_12704,N_12938);
or U13896 (N_13896,N_12135,N_12210);
nand U13897 (N_13897,N_12431,N_12377);
nand U13898 (N_13898,N_12675,N_12575);
and U13899 (N_13899,N_12821,N_12044);
nor U13900 (N_13900,N_12457,N_12796);
and U13901 (N_13901,N_12969,N_12237);
and U13902 (N_13902,N_12015,N_12650);
or U13903 (N_13903,N_12527,N_12466);
nor U13904 (N_13904,N_12753,N_12054);
and U13905 (N_13905,N_12677,N_12589);
xor U13906 (N_13906,N_12556,N_12582);
or U13907 (N_13907,N_12478,N_12692);
nand U13908 (N_13908,N_12429,N_12013);
nor U13909 (N_13909,N_12530,N_12789);
xor U13910 (N_13910,N_12722,N_12367);
nand U13911 (N_13911,N_12461,N_12476);
nor U13912 (N_13912,N_12840,N_12916);
or U13913 (N_13913,N_12739,N_12326);
nand U13914 (N_13914,N_12664,N_12726);
xnor U13915 (N_13915,N_12990,N_12319);
or U13916 (N_13916,N_12822,N_12451);
nand U13917 (N_13917,N_12745,N_12465);
and U13918 (N_13918,N_12571,N_12674);
nand U13919 (N_13919,N_12398,N_12596);
xor U13920 (N_13920,N_12840,N_12102);
nand U13921 (N_13921,N_12994,N_12825);
xor U13922 (N_13922,N_12294,N_12281);
nor U13923 (N_13923,N_12272,N_12520);
and U13924 (N_13924,N_12290,N_12852);
nand U13925 (N_13925,N_12101,N_12307);
nor U13926 (N_13926,N_12065,N_12053);
nor U13927 (N_13927,N_12937,N_12362);
or U13928 (N_13928,N_12598,N_12940);
nor U13929 (N_13929,N_12097,N_12971);
nor U13930 (N_13930,N_12021,N_12916);
xnor U13931 (N_13931,N_12541,N_12743);
xor U13932 (N_13932,N_12514,N_12032);
or U13933 (N_13933,N_12689,N_12001);
and U13934 (N_13934,N_12942,N_12854);
nor U13935 (N_13935,N_12622,N_12524);
nand U13936 (N_13936,N_12813,N_12694);
or U13937 (N_13937,N_12904,N_12243);
xnor U13938 (N_13938,N_12103,N_12650);
or U13939 (N_13939,N_12180,N_12749);
nand U13940 (N_13940,N_12538,N_12025);
nand U13941 (N_13941,N_12172,N_12142);
and U13942 (N_13942,N_12930,N_12552);
and U13943 (N_13943,N_12407,N_12026);
or U13944 (N_13944,N_12172,N_12743);
xnor U13945 (N_13945,N_12058,N_12395);
nand U13946 (N_13946,N_12981,N_12241);
nor U13947 (N_13947,N_12025,N_12923);
xor U13948 (N_13948,N_12169,N_12545);
nor U13949 (N_13949,N_12837,N_12032);
nor U13950 (N_13950,N_12521,N_12970);
nand U13951 (N_13951,N_12602,N_12133);
nor U13952 (N_13952,N_12325,N_12485);
nor U13953 (N_13953,N_12917,N_12746);
or U13954 (N_13954,N_12840,N_12248);
or U13955 (N_13955,N_12904,N_12692);
or U13956 (N_13956,N_12343,N_12050);
nor U13957 (N_13957,N_12630,N_12017);
and U13958 (N_13958,N_12752,N_12480);
and U13959 (N_13959,N_12351,N_12910);
or U13960 (N_13960,N_12390,N_12193);
or U13961 (N_13961,N_12542,N_12328);
or U13962 (N_13962,N_12581,N_12698);
nor U13963 (N_13963,N_12664,N_12786);
or U13964 (N_13964,N_12144,N_12342);
and U13965 (N_13965,N_12281,N_12110);
xor U13966 (N_13966,N_12992,N_12897);
or U13967 (N_13967,N_12223,N_12282);
or U13968 (N_13968,N_12568,N_12714);
xor U13969 (N_13969,N_12484,N_12838);
or U13970 (N_13970,N_12190,N_12532);
nor U13971 (N_13971,N_12202,N_12760);
nand U13972 (N_13972,N_12624,N_12140);
or U13973 (N_13973,N_12325,N_12956);
and U13974 (N_13974,N_12695,N_12576);
nor U13975 (N_13975,N_12321,N_12743);
nor U13976 (N_13976,N_12014,N_12825);
xnor U13977 (N_13977,N_12634,N_12226);
nand U13978 (N_13978,N_12350,N_12362);
and U13979 (N_13979,N_12900,N_12562);
or U13980 (N_13980,N_12651,N_12845);
xor U13981 (N_13981,N_12709,N_12954);
and U13982 (N_13982,N_12283,N_12047);
nand U13983 (N_13983,N_12063,N_12459);
nand U13984 (N_13984,N_12536,N_12872);
nor U13985 (N_13985,N_12034,N_12201);
nand U13986 (N_13986,N_12516,N_12043);
and U13987 (N_13987,N_12669,N_12586);
or U13988 (N_13988,N_12598,N_12770);
or U13989 (N_13989,N_12284,N_12129);
nor U13990 (N_13990,N_12885,N_12283);
and U13991 (N_13991,N_12249,N_12903);
nor U13992 (N_13992,N_12566,N_12374);
nor U13993 (N_13993,N_12945,N_12969);
and U13994 (N_13994,N_12881,N_12464);
nor U13995 (N_13995,N_12292,N_12897);
nor U13996 (N_13996,N_12687,N_12109);
nor U13997 (N_13997,N_12899,N_12146);
and U13998 (N_13998,N_12209,N_12139);
nor U13999 (N_13999,N_12653,N_12030);
and U14000 (N_14000,N_13064,N_13602);
xnor U14001 (N_14001,N_13437,N_13541);
xor U14002 (N_14002,N_13399,N_13781);
nor U14003 (N_14003,N_13154,N_13691);
nand U14004 (N_14004,N_13992,N_13877);
xnor U14005 (N_14005,N_13755,N_13645);
xnor U14006 (N_14006,N_13463,N_13943);
and U14007 (N_14007,N_13585,N_13606);
nor U14008 (N_14008,N_13939,N_13707);
nor U14009 (N_14009,N_13044,N_13546);
and U14010 (N_14010,N_13816,N_13516);
and U14011 (N_14011,N_13205,N_13689);
and U14012 (N_14012,N_13977,N_13754);
or U14013 (N_14013,N_13176,N_13016);
or U14014 (N_14014,N_13747,N_13396);
or U14015 (N_14015,N_13037,N_13393);
nor U14016 (N_14016,N_13252,N_13532);
or U14017 (N_14017,N_13423,N_13690);
nand U14018 (N_14018,N_13530,N_13562);
and U14019 (N_14019,N_13628,N_13626);
xor U14020 (N_14020,N_13269,N_13674);
nand U14021 (N_14021,N_13948,N_13245);
nand U14022 (N_14022,N_13542,N_13419);
xnor U14023 (N_14023,N_13919,N_13930);
nor U14024 (N_14024,N_13327,N_13696);
or U14025 (N_14025,N_13354,N_13957);
nor U14026 (N_14026,N_13923,N_13384);
and U14027 (N_14027,N_13027,N_13882);
xnor U14028 (N_14028,N_13501,N_13879);
nand U14029 (N_14029,N_13139,N_13905);
xor U14030 (N_14030,N_13869,N_13475);
nor U14031 (N_14031,N_13584,N_13296);
nand U14032 (N_14032,N_13819,N_13920);
and U14033 (N_14033,N_13109,N_13328);
or U14034 (N_14034,N_13211,N_13650);
nand U14035 (N_14035,N_13589,N_13307);
or U14036 (N_14036,N_13389,N_13439);
nor U14037 (N_14037,N_13941,N_13732);
nor U14038 (N_14038,N_13421,N_13518);
or U14039 (N_14039,N_13828,N_13420);
xnor U14040 (N_14040,N_13125,N_13914);
and U14041 (N_14041,N_13052,N_13092);
nand U14042 (N_14042,N_13592,N_13167);
or U14043 (N_14043,N_13374,N_13385);
nor U14044 (N_14044,N_13694,N_13442);
and U14045 (N_14045,N_13314,N_13901);
or U14046 (N_14046,N_13752,N_13241);
or U14047 (N_14047,N_13034,N_13731);
xor U14048 (N_14048,N_13257,N_13803);
nor U14049 (N_14049,N_13579,N_13196);
and U14050 (N_14050,N_13168,N_13062);
and U14051 (N_14051,N_13112,N_13020);
xnor U14052 (N_14052,N_13505,N_13724);
nor U14053 (N_14053,N_13456,N_13593);
and U14054 (N_14054,N_13447,N_13985);
or U14055 (N_14055,N_13911,N_13331);
and U14056 (N_14056,N_13410,N_13527);
and U14057 (N_14057,N_13906,N_13619);
xor U14058 (N_14058,N_13093,N_13630);
xor U14059 (N_14059,N_13843,N_13443);
or U14060 (N_14060,N_13534,N_13433);
and U14061 (N_14061,N_13487,N_13591);
xor U14062 (N_14062,N_13657,N_13868);
nor U14063 (N_14063,N_13067,N_13637);
or U14064 (N_14064,N_13239,N_13286);
nand U14065 (N_14065,N_13232,N_13348);
or U14066 (N_14066,N_13959,N_13672);
nand U14067 (N_14067,N_13976,N_13150);
nand U14068 (N_14068,N_13537,N_13636);
or U14069 (N_14069,N_13345,N_13012);
nand U14070 (N_14070,N_13357,N_13807);
and U14071 (N_14071,N_13453,N_13272);
and U14072 (N_14072,N_13055,N_13426);
or U14073 (N_14073,N_13014,N_13318);
xor U14074 (N_14074,N_13370,N_13369);
or U14075 (N_14075,N_13207,N_13829);
and U14076 (N_14076,N_13367,N_13342);
nand U14077 (N_14077,N_13573,N_13336);
xor U14078 (N_14078,N_13146,N_13737);
nor U14079 (N_14079,N_13451,N_13152);
nor U14080 (N_14080,N_13326,N_13551);
and U14081 (N_14081,N_13667,N_13559);
and U14082 (N_14082,N_13665,N_13851);
nand U14083 (N_14083,N_13801,N_13123);
and U14084 (N_14084,N_13263,N_13891);
xor U14085 (N_14085,N_13346,N_13655);
nand U14086 (N_14086,N_13835,N_13547);
and U14087 (N_14087,N_13065,N_13250);
nand U14088 (N_14088,N_13554,N_13225);
and U14089 (N_14089,N_13129,N_13646);
xnor U14090 (N_14090,N_13108,N_13821);
nand U14091 (N_14091,N_13942,N_13254);
or U14092 (N_14092,N_13928,N_13022);
and U14093 (N_14093,N_13508,N_13251);
or U14094 (N_14094,N_13805,N_13446);
nand U14095 (N_14095,N_13838,N_13716);
xnor U14096 (N_14096,N_13074,N_13302);
nand U14097 (N_14097,N_13767,N_13049);
nor U14098 (N_14098,N_13436,N_13826);
nand U14099 (N_14099,N_13746,N_13347);
nor U14100 (N_14100,N_13811,N_13409);
and U14101 (N_14101,N_13961,N_13684);
xnor U14102 (N_14102,N_13395,N_13733);
xor U14103 (N_14103,N_13777,N_13535);
nor U14104 (N_14104,N_13790,N_13968);
nor U14105 (N_14105,N_13709,N_13122);
xnor U14106 (N_14106,N_13687,N_13742);
and U14107 (N_14107,N_13308,N_13333);
nor U14108 (N_14108,N_13043,N_13170);
xnor U14109 (N_14109,N_13749,N_13499);
nor U14110 (N_14110,N_13855,N_13414);
nand U14111 (N_14111,N_13768,N_13236);
nor U14112 (N_14112,N_13915,N_13373);
nand U14113 (N_14113,N_13633,N_13330);
nor U14114 (N_14114,N_13470,N_13886);
or U14115 (N_14115,N_13735,N_13116);
nor U14116 (N_14116,N_13040,N_13932);
or U14117 (N_14117,N_13320,N_13360);
nor U14118 (N_14118,N_13009,N_13458);
nor U14119 (N_14119,N_13235,N_13944);
nand U14120 (N_14120,N_13144,N_13185);
nor U14121 (N_14121,N_13676,N_13722);
xnor U14122 (N_14122,N_13836,N_13918);
nor U14123 (N_14123,N_13169,N_13000);
nand U14124 (N_14124,N_13311,N_13564);
xnor U14125 (N_14125,N_13188,N_13153);
or U14126 (N_14126,N_13391,N_13402);
and U14127 (N_14127,N_13025,N_13625);
and U14128 (N_14128,N_13164,N_13779);
xor U14129 (N_14129,N_13529,N_13947);
and U14130 (N_14130,N_13179,N_13230);
nand U14131 (N_14131,N_13117,N_13723);
xnor U14132 (N_14132,N_13449,N_13576);
nand U14133 (N_14133,N_13216,N_13292);
xor U14134 (N_14134,N_13841,N_13708);
xnor U14135 (N_14135,N_13830,N_13862);
xnor U14136 (N_14136,N_13006,N_13791);
or U14137 (N_14137,N_13114,N_13917);
nor U14138 (N_14138,N_13995,N_13435);
and U14139 (N_14139,N_13111,N_13846);
nand U14140 (N_14140,N_13989,N_13969);
nor U14141 (N_14141,N_13951,N_13197);
xor U14142 (N_14142,N_13804,N_13351);
nand U14143 (N_14143,N_13519,N_13823);
nor U14144 (N_14144,N_13679,N_13643);
and U14145 (N_14145,N_13668,N_13387);
xor U14146 (N_14146,N_13334,N_13894);
or U14147 (N_14147,N_13454,N_13990);
nor U14148 (N_14148,N_13916,N_13343);
nor U14149 (N_14149,N_13743,N_13660);
nand U14150 (N_14150,N_13595,N_13898);
or U14151 (N_14151,N_13653,N_13946);
and U14152 (N_14152,N_13087,N_13960);
nand U14153 (N_14153,N_13448,N_13215);
or U14154 (N_14154,N_13753,N_13670);
or U14155 (N_14155,N_13011,N_13121);
or U14156 (N_14156,N_13935,N_13432);
and U14157 (N_14157,N_13528,N_13945);
nor U14158 (N_14158,N_13962,N_13227);
and U14159 (N_14159,N_13166,N_13353);
nor U14160 (N_14160,N_13762,N_13477);
nor U14161 (N_14161,N_13714,N_13605);
or U14162 (N_14162,N_13986,N_13118);
xnor U14163 (N_14163,N_13113,N_13305);
and U14164 (N_14164,N_13566,N_13912);
or U14165 (N_14165,N_13298,N_13688);
and U14166 (N_14166,N_13558,N_13023);
or U14167 (N_14167,N_13485,N_13588);
or U14168 (N_14168,N_13904,N_13213);
nor U14169 (N_14169,N_13967,N_13194);
nor U14170 (N_14170,N_13865,N_13775);
nor U14171 (N_14171,N_13618,N_13332);
nor U14172 (N_14172,N_13431,N_13565);
and U14173 (N_14173,N_13563,N_13103);
nor U14174 (N_14174,N_13497,N_13469);
nor U14175 (N_14175,N_13950,N_13147);
xor U14176 (N_14176,N_13323,N_13725);
or U14177 (N_14177,N_13897,N_13763);
nor U14178 (N_14178,N_13210,N_13165);
nor U14179 (N_14179,N_13623,N_13979);
and U14180 (N_14180,N_13099,N_13089);
nor U14181 (N_14181,N_13524,N_13892);
xor U14182 (N_14182,N_13603,N_13030);
and U14183 (N_14183,N_13736,N_13693);
xnor U14184 (N_14184,N_13137,N_13727);
and U14185 (N_14185,N_13284,N_13772);
and U14186 (N_14186,N_13671,N_13617);
xnor U14187 (N_14187,N_13440,N_13751);
nor U14188 (N_14188,N_13304,N_13711);
and U14189 (N_14189,N_13638,N_13640);
xnor U14190 (N_14190,N_13664,N_13577);
and U14191 (N_14191,N_13492,N_13549);
or U14192 (N_14192,N_13158,N_13494);
and U14193 (N_14193,N_13789,N_13632);
nand U14194 (N_14194,N_13063,N_13466);
nand U14195 (N_14195,N_13024,N_13856);
and U14196 (N_14196,N_13248,N_13299);
nor U14197 (N_14197,N_13130,N_13783);
xor U14198 (N_14198,N_13622,N_13875);
nor U14199 (N_14199,N_13276,N_13583);
nand U14200 (N_14200,N_13788,N_13091);
or U14201 (N_14201,N_13261,N_13859);
xor U14202 (N_14202,N_13329,N_13386);
or U14203 (N_14203,N_13656,N_13090);
nand U14204 (N_14204,N_13096,N_13321);
or U14205 (N_14205,N_13569,N_13922);
xnor U14206 (N_14206,N_13008,N_13193);
or U14207 (N_14207,N_13186,N_13933);
nand U14208 (N_14208,N_13580,N_13766);
nor U14209 (N_14209,N_13195,N_13212);
xnor U14210 (N_14210,N_13774,N_13548);
nand U14211 (N_14211,N_13682,N_13019);
xnor U14212 (N_14212,N_13428,N_13502);
xnor U14213 (N_14213,N_13110,N_13240);
nor U14214 (N_14214,N_13281,N_13315);
nand U14215 (N_14215,N_13837,N_13010);
nand U14216 (N_14216,N_13124,N_13231);
nand U14217 (N_14217,N_13247,N_13713);
xor U14218 (N_14218,N_13870,N_13078);
or U14219 (N_14219,N_13127,N_13417);
and U14220 (N_14220,N_13057,N_13764);
nand U14221 (N_14221,N_13316,N_13552);
nand U14222 (N_14222,N_13517,N_13770);
xor U14223 (N_14223,N_13203,N_13474);
xnor U14224 (N_14224,N_13457,N_13940);
or U14225 (N_14225,N_13018,N_13536);
and U14226 (N_14226,N_13913,N_13441);
xnor U14227 (N_14227,N_13059,N_13931);
nor U14228 (N_14228,N_13756,N_13377);
and U14229 (N_14229,N_13082,N_13309);
xnor U14230 (N_14230,N_13482,N_13980);
nand U14231 (N_14231,N_13480,N_13275);
nand U14232 (N_14232,N_13553,N_13219);
nand U14233 (N_14233,N_13253,N_13578);
and U14234 (N_14234,N_13404,N_13523);
xnor U14235 (N_14235,N_13809,N_13908);
and U14236 (N_14236,N_13380,N_13242);
nor U14237 (N_14237,N_13860,N_13975);
and U14238 (N_14238,N_13413,N_13228);
nor U14239 (N_14239,N_13984,N_13184);
nor U14240 (N_14240,N_13647,N_13484);
and U14241 (N_14241,N_13631,N_13700);
nand U14242 (N_14242,N_13629,N_13155);
or U14243 (N_14243,N_13526,N_13949);
or U14244 (N_14244,N_13422,N_13854);
or U14245 (N_14245,N_13221,N_13080);
and U14246 (N_14246,N_13408,N_13368);
nand U14247 (N_14247,N_13738,N_13258);
or U14248 (N_14248,N_13782,N_13274);
or U14249 (N_14249,N_13310,N_13681);
nand U14250 (N_14250,N_13467,N_13596);
xnor U14251 (N_14251,N_13148,N_13827);
or U14252 (N_14252,N_13704,N_13649);
nor U14253 (N_14253,N_13105,N_13157);
and U14254 (N_14254,N_13133,N_13478);
or U14255 (N_14255,N_13863,N_13615);
xor U14256 (N_14256,N_13450,N_13001);
and U14257 (N_14257,N_13703,N_13255);
xnor U14258 (N_14258,N_13972,N_13509);
nor U14259 (N_14259,N_13680,N_13060);
nor U14260 (N_14260,N_13178,N_13512);
nor U14261 (N_14261,N_13268,N_13459);
nand U14262 (N_14262,N_13493,N_13295);
nand U14263 (N_14263,N_13156,N_13319);
and U14264 (N_14264,N_13107,N_13683);
and U14265 (N_14265,N_13607,N_13717);
xor U14266 (N_14266,N_13120,N_13445);
nor U14267 (N_14267,N_13895,N_13608);
nor U14268 (N_14268,N_13223,N_13085);
or U14269 (N_14269,N_13266,N_13802);
nor U14270 (N_14270,N_13748,N_13934);
nor U14271 (N_14271,N_13719,N_13925);
xor U14272 (N_14272,N_13135,N_13356);
nand U14273 (N_14273,N_13287,N_13624);
or U14274 (N_14274,N_13866,N_13238);
nor U14275 (N_14275,N_13705,N_13698);
xnor U14276 (N_14276,N_13887,N_13013);
nor U14277 (N_14277,N_13372,N_13411);
and U14278 (N_14278,N_13106,N_13045);
or U14279 (N_14279,N_13094,N_13893);
xor U14280 (N_14280,N_13036,N_13204);
nand U14281 (N_14281,N_13283,N_13639);
or U14282 (N_14282,N_13574,N_13233);
xnor U14283 (N_14283,N_13744,N_13398);
xnor U14284 (N_14284,N_13531,N_13504);
or U14285 (N_14285,N_13427,N_13002);
nor U14286 (N_14286,N_13822,N_13198);
xnor U14287 (N_14287,N_13889,N_13510);
nand U14288 (N_14288,N_13750,N_13361);
or U14289 (N_14289,N_13814,N_13614);
and U14290 (N_14290,N_13359,N_13648);
nor U14291 (N_14291,N_13817,N_13175);
xnor U14292 (N_14292,N_13026,N_13952);
or U14293 (N_14293,N_13780,N_13539);
nor U14294 (N_14294,N_13885,N_13881);
and U14295 (N_14295,N_13192,N_13871);
or U14296 (N_14296,N_13191,N_13695);
and U14297 (N_14297,N_13128,N_13878);
or U14298 (N_14298,N_13760,N_13824);
xnor U14299 (N_14299,N_13813,N_13134);
and U14300 (N_14300,N_13180,N_13567);
and U14301 (N_14301,N_13349,N_13726);
nor U14302 (N_14302,N_13903,N_13046);
nand U14303 (N_14303,N_13503,N_13799);
or U14304 (N_14304,N_13187,N_13340);
or U14305 (N_14305,N_13362,N_13634);
nor U14306 (N_14306,N_13997,N_13425);
xnor U14307 (N_14307,N_13874,N_13787);
or U14308 (N_14308,N_13429,N_13061);
nand U14309 (N_14309,N_13481,N_13661);
or U14310 (N_14310,N_13488,N_13850);
and U14311 (N_14311,N_13872,N_13270);
or U14312 (N_14312,N_13285,N_13430);
and U14313 (N_14313,N_13966,N_13438);
xor U14314 (N_14314,N_13452,N_13610);
or U14315 (N_14315,N_13658,N_13963);
nor U14316 (N_14316,N_13273,N_13303);
xor U14317 (N_14317,N_13005,N_13621);
nand U14318 (N_14318,N_13352,N_13675);
or U14319 (N_14319,N_13325,N_13808);
nand U14320 (N_14320,N_13379,N_13070);
nand U14321 (N_14321,N_13476,N_13172);
and U14322 (N_14322,N_13490,N_13224);
and U14323 (N_14323,N_13810,N_13594);
nand U14324 (N_14324,N_13383,N_13142);
nand U14325 (N_14325,N_13282,N_13699);
nand U14326 (N_14326,N_13978,N_13145);
xnor U14327 (N_14327,N_13246,N_13294);
nand U14328 (N_14328,N_13183,N_13797);
nor U14329 (N_14329,N_13104,N_13338);
and U14330 (N_14330,N_13132,N_13712);
nand U14331 (N_14331,N_13820,N_13279);
xnor U14332 (N_14332,N_13720,N_13991);
nor U14333 (N_14333,N_13056,N_13394);
nand U14334 (N_14334,N_13785,N_13601);
and U14335 (N_14335,N_13867,N_13496);
nand U14336 (N_14336,N_13514,N_13642);
or U14337 (N_14337,N_13718,N_13407);
and U14338 (N_14338,N_13289,N_13842);
and U14339 (N_14339,N_13757,N_13815);
nand U14340 (N_14340,N_13831,N_13138);
xnor U14341 (N_14341,N_13079,N_13858);
xor U14342 (N_14342,N_13769,N_13460);
or U14343 (N_14343,N_13806,N_13249);
nand U14344 (N_14344,N_13201,N_13500);
nand U14345 (N_14345,N_13265,N_13880);
nand U14346 (N_14346,N_13344,N_13378);
or U14347 (N_14347,N_13115,N_13035);
xor U14348 (N_14348,N_13256,N_13126);
or U14349 (N_14349,N_13371,N_13987);
and U14350 (N_14350,N_13088,N_13406);
nor U14351 (N_14351,N_13277,N_13927);
or U14352 (N_14352,N_13861,N_13786);
xnor U14353 (N_14353,N_13392,N_13416);
or U14354 (N_14354,N_13208,N_13054);
and U14355 (N_14355,N_13084,N_13173);
nor U14356 (N_14356,N_13513,N_13613);
nor U14357 (N_14357,N_13243,N_13555);
nor U14358 (N_14358,N_13654,N_13021);
nand U14359 (N_14359,N_13560,N_13050);
nand U14360 (N_14360,N_13652,N_13635);
nor U14361 (N_14361,N_13489,N_13483);
and U14362 (N_14362,N_13032,N_13572);
or U14363 (N_14363,N_13244,N_13031);
nand U14364 (N_14364,N_13515,N_13520);
or U14365 (N_14365,N_13974,N_13970);
nand U14366 (N_14366,N_13793,N_13400);
or U14367 (N_14367,N_13401,N_13715);
nor U14368 (N_14368,N_13234,N_13069);
nand U14369 (N_14369,N_13812,N_13921);
and U14370 (N_14370,N_13883,N_13119);
and U14371 (N_14371,N_13073,N_13382);
xor U14372 (N_14372,N_13051,N_13616);
xnor U14373 (N_14373,N_13728,N_13486);
or U14374 (N_14374,N_13544,N_13954);
nand U14375 (N_14375,N_13086,N_13988);
nor U14376 (N_14376,N_13907,N_13190);
nand U14377 (N_14377,N_13053,N_13834);
xnor U14378 (N_14378,N_13557,N_13376);
or U14379 (N_14379,N_13609,N_13202);
nor U14380 (N_14380,N_13507,N_13038);
nand U14381 (N_14381,N_13561,N_13405);
nand U14382 (N_14382,N_13206,N_13271);
and U14383 (N_14383,N_13926,N_13424);
or U14384 (N_14384,N_13160,N_13097);
nand U14385 (N_14385,N_13259,N_13182);
xor U14386 (N_14386,N_13522,N_13083);
and U14387 (N_14387,N_13100,N_13996);
xnor U14388 (N_14388,N_13909,N_13971);
or U14389 (N_14389,N_13355,N_13076);
nor U14390 (N_14390,N_13390,N_13288);
nor U14391 (N_14391,N_13844,N_13773);
xnor U14392 (N_14392,N_13312,N_13095);
nor U14393 (N_14393,N_13998,N_13776);
nor U14394 (N_14394,N_13848,N_13464);
or U14395 (N_14395,N_13759,N_13042);
nor U14396 (N_14396,N_13301,N_13039);
and U14397 (N_14397,N_13599,N_13291);
and U14398 (N_14398,N_13899,N_13910);
nor U14399 (N_14399,N_13644,N_13041);
and U14400 (N_14400,N_13545,N_13597);
nand U14401 (N_14401,N_13058,N_13543);
nand U14402 (N_14402,N_13778,N_13677);
nand U14403 (N_14403,N_13651,N_13798);
nand U14404 (N_14404,N_13163,N_13101);
xor U14405 (N_14405,N_13800,N_13506);
and U14406 (N_14406,N_13612,N_13784);
and U14407 (N_14407,N_13701,N_13324);
or U14408 (N_14408,N_13556,N_13571);
and U14409 (N_14409,N_13833,N_13364);
or U14410 (N_14410,N_13604,N_13162);
xor U14411 (N_14411,N_13847,N_13840);
or U14412 (N_14412,N_13365,N_13418);
nand U14413 (N_14413,N_13993,N_13350);
or U14414 (N_14414,N_13159,N_13958);
nand U14415 (N_14415,N_13662,N_13412);
nor U14416 (N_14416,N_13171,N_13741);
nand U14417 (N_14417,N_13048,N_13358);
xor U14418 (N_14418,N_13761,N_13953);
nor U14419 (N_14419,N_13825,N_13028);
and U14420 (N_14420,N_13697,N_13888);
nor U14421 (N_14421,N_13669,N_13538);
nand U14422 (N_14422,N_13666,N_13397);
nand U14423 (N_14423,N_13465,N_13590);
or U14424 (N_14424,N_13745,N_13140);
nand U14425 (N_14425,N_13280,N_13794);
nand U14426 (N_14426,N_13226,N_13568);
or U14427 (N_14427,N_13363,N_13857);
nand U14428 (N_14428,N_13017,N_13004);
nor U14429 (N_14429,N_13322,N_13900);
or U14430 (N_14430,N_13143,N_13290);
xor U14431 (N_14431,N_13381,N_13199);
or U14432 (N_14432,N_13511,N_13102);
nand U14433 (N_14433,N_13771,N_13994);
nand U14434 (N_14434,N_13181,N_13721);
nand U14435 (N_14435,N_13278,N_13229);
nand U14436 (N_14436,N_13796,N_13479);
and U14437 (N_14437,N_13938,N_13792);
xor U14438 (N_14438,N_13077,N_13983);
and U14439 (N_14439,N_13313,N_13071);
nor U14440 (N_14440,N_13853,N_13066);
nand U14441 (N_14441,N_13317,N_13673);
nor U14442 (N_14442,N_13678,N_13765);
or U14443 (N_14443,N_13864,N_13471);
nand U14444 (N_14444,N_13525,N_13686);
nor U14445 (N_14445,N_13982,N_13260);
and U14446 (N_14446,N_13575,N_13141);
xnor U14447 (N_14447,N_13267,N_13174);
or U14448 (N_14448,N_13600,N_13706);
and U14449 (N_14449,N_13586,N_13964);
or U14450 (N_14450,N_13849,N_13293);
xnor U14451 (N_14451,N_13209,N_13692);
or U14452 (N_14452,N_13029,N_13047);
and U14453 (N_14453,N_13461,N_13220);
and U14454 (N_14454,N_13729,N_13003);
nand U14455 (N_14455,N_13300,N_13068);
and U14456 (N_14456,N_13902,N_13710);
nor U14457 (N_14457,N_13177,N_13341);
nand U14458 (N_14458,N_13415,N_13237);
nand U14459 (N_14459,N_13582,N_13873);
or U14460 (N_14460,N_13955,N_13473);
nand U14461 (N_14461,N_13075,N_13161);
and U14462 (N_14462,N_13081,N_13550);
nand U14463 (N_14463,N_13533,N_13015);
xnor U14464 (N_14464,N_13999,N_13521);
nor U14465 (N_14465,N_13462,N_13734);
or U14466 (N_14466,N_13956,N_13262);
nand U14467 (N_14467,N_13098,N_13007);
nand U14468 (N_14468,N_13965,N_13217);
and U14469 (N_14469,N_13896,N_13659);
nor U14470 (N_14470,N_13200,N_13620);
nand U14471 (N_14471,N_13876,N_13758);
nor U14472 (N_14472,N_13149,N_13685);
and U14473 (N_14473,N_13598,N_13730);
or U14474 (N_14474,N_13339,N_13335);
or U14475 (N_14475,N_13839,N_13366);
nand U14476 (N_14476,N_13375,N_13214);
and U14477 (N_14477,N_13627,N_13740);
xnor U14478 (N_14478,N_13929,N_13388);
and U14479 (N_14479,N_13337,N_13570);
and U14480 (N_14480,N_13498,N_13491);
xnor U14481 (N_14481,N_13434,N_13587);
nor U14482 (N_14482,N_13136,N_13937);
nor U14483 (N_14483,N_13884,N_13297);
or U14484 (N_14484,N_13189,N_13218);
nor U14485 (N_14485,N_13832,N_13033);
nor U14486 (N_14486,N_13455,N_13981);
xor U14487 (N_14487,N_13818,N_13581);
and U14488 (N_14488,N_13472,N_13936);
and U14489 (N_14489,N_13468,N_13795);
xnor U14490 (N_14490,N_13495,N_13973);
nor U14491 (N_14491,N_13540,N_13924);
and U14492 (N_14492,N_13131,N_13641);
nand U14493 (N_14493,N_13151,N_13444);
and U14494 (N_14494,N_13702,N_13890);
or U14495 (N_14495,N_13072,N_13222);
nor U14496 (N_14496,N_13403,N_13611);
xor U14497 (N_14497,N_13306,N_13264);
nand U14498 (N_14498,N_13852,N_13663);
xnor U14499 (N_14499,N_13845,N_13739);
and U14500 (N_14500,N_13557,N_13114);
nand U14501 (N_14501,N_13514,N_13391);
nand U14502 (N_14502,N_13267,N_13366);
nor U14503 (N_14503,N_13480,N_13775);
xor U14504 (N_14504,N_13386,N_13879);
xor U14505 (N_14505,N_13677,N_13382);
nand U14506 (N_14506,N_13758,N_13861);
and U14507 (N_14507,N_13345,N_13108);
and U14508 (N_14508,N_13032,N_13199);
nor U14509 (N_14509,N_13950,N_13852);
or U14510 (N_14510,N_13181,N_13205);
nand U14511 (N_14511,N_13899,N_13573);
xor U14512 (N_14512,N_13689,N_13072);
nor U14513 (N_14513,N_13211,N_13068);
and U14514 (N_14514,N_13608,N_13490);
and U14515 (N_14515,N_13128,N_13139);
nor U14516 (N_14516,N_13624,N_13385);
xor U14517 (N_14517,N_13330,N_13366);
nor U14518 (N_14518,N_13130,N_13711);
nor U14519 (N_14519,N_13254,N_13505);
and U14520 (N_14520,N_13906,N_13229);
xnor U14521 (N_14521,N_13456,N_13452);
nand U14522 (N_14522,N_13650,N_13099);
nand U14523 (N_14523,N_13950,N_13580);
or U14524 (N_14524,N_13575,N_13317);
and U14525 (N_14525,N_13171,N_13365);
or U14526 (N_14526,N_13553,N_13221);
or U14527 (N_14527,N_13768,N_13327);
xor U14528 (N_14528,N_13981,N_13445);
nand U14529 (N_14529,N_13905,N_13120);
xnor U14530 (N_14530,N_13552,N_13409);
nand U14531 (N_14531,N_13823,N_13005);
or U14532 (N_14532,N_13596,N_13293);
xnor U14533 (N_14533,N_13122,N_13667);
nor U14534 (N_14534,N_13561,N_13474);
nand U14535 (N_14535,N_13346,N_13886);
nand U14536 (N_14536,N_13030,N_13700);
or U14537 (N_14537,N_13148,N_13973);
or U14538 (N_14538,N_13020,N_13503);
or U14539 (N_14539,N_13118,N_13121);
and U14540 (N_14540,N_13526,N_13761);
and U14541 (N_14541,N_13102,N_13108);
xnor U14542 (N_14542,N_13703,N_13600);
and U14543 (N_14543,N_13344,N_13162);
and U14544 (N_14544,N_13816,N_13395);
nand U14545 (N_14545,N_13673,N_13192);
nand U14546 (N_14546,N_13098,N_13389);
xnor U14547 (N_14547,N_13170,N_13380);
nor U14548 (N_14548,N_13265,N_13529);
nand U14549 (N_14549,N_13267,N_13804);
or U14550 (N_14550,N_13645,N_13628);
nor U14551 (N_14551,N_13261,N_13321);
nand U14552 (N_14552,N_13319,N_13445);
and U14553 (N_14553,N_13886,N_13526);
nand U14554 (N_14554,N_13079,N_13433);
xor U14555 (N_14555,N_13311,N_13165);
nand U14556 (N_14556,N_13558,N_13124);
nor U14557 (N_14557,N_13142,N_13376);
nand U14558 (N_14558,N_13419,N_13398);
or U14559 (N_14559,N_13656,N_13318);
nand U14560 (N_14560,N_13837,N_13444);
nor U14561 (N_14561,N_13030,N_13308);
and U14562 (N_14562,N_13893,N_13646);
or U14563 (N_14563,N_13038,N_13996);
nor U14564 (N_14564,N_13523,N_13692);
or U14565 (N_14565,N_13140,N_13901);
xnor U14566 (N_14566,N_13173,N_13279);
and U14567 (N_14567,N_13155,N_13432);
xor U14568 (N_14568,N_13356,N_13994);
xnor U14569 (N_14569,N_13768,N_13316);
and U14570 (N_14570,N_13506,N_13624);
nor U14571 (N_14571,N_13117,N_13693);
xnor U14572 (N_14572,N_13511,N_13563);
nor U14573 (N_14573,N_13463,N_13162);
and U14574 (N_14574,N_13321,N_13043);
nand U14575 (N_14575,N_13840,N_13694);
nand U14576 (N_14576,N_13111,N_13726);
nor U14577 (N_14577,N_13239,N_13949);
nand U14578 (N_14578,N_13478,N_13816);
nand U14579 (N_14579,N_13403,N_13740);
nor U14580 (N_14580,N_13411,N_13126);
or U14581 (N_14581,N_13596,N_13428);
and U14582 (N_14582,N_13484,N_13959);
and U14583 (N_14583,N_13896,N_13863);
xor U14584 (N_14584,N_13290,N_13282);
or U14585 (N_14585,N_13776,N_13719);
nor U14586 (N_14586,N_13389,N_13194);
xnor U14587 (N_14587,N_13234,N_13754);
and U14588 (N_14588,N_13962,N_13203);
nor U14589 (N_14589,N_13022,N_13184);
nand U14590 (N_14590,N_13721,N_13219);
nor U14591 (N_14591,N_13571,N_13743);
xnor U14592 (N_14592,N_13451,N_13911);
or U14593 (N_14593,N_13006,N_13661);
nor U14594 (N_14594,N_13460,N_13353);
xor U14595 (N_14595,N_13238,N_13270);
nand U14596 (N_14596,N_13725,N_13917);
and U14597 (N_14597,N_13514,N_13487);
nand U14598 (N_14598,N_13582,N_13012);
nand U14599 (N_14599,N_13001,N_13572);
or U14600 (N_14600,N_13037,N_13615);
and U14601 (N_14601,N_13551,N_13838);
xor U14602 (N_14602,N_13386,N_13627);
xor U14603 (N_14603,N_13077,N_13095);
nor U14604 (N_14604,N_13251,N_13178);
xnor U14605 (N_14605,N_13466,N_13998);
and U14606 (N_14606,N_13513,N_13892);
and U14607 (N_14607,N_13367,N_13112);
xor U14608 (N_14608,N_13332,N_13573);
nor U14609 (N_14609,N_13896,N_13479);
xor U14610 (N_14610,N_13707,N_13568);
xnor U14611 (N_14611,N_13842,N_13860);
and U14612 (N_14612,N_13555,N_13920);
and U14613 (N_14613,N_13580,N_13582);
nand U14614 (N_14614,N_13157,N_13372);
nor U14615 (N_14615,N_13937,N_13985);
nor U14616 (N_14616,N_13479,N_13308);
or U14617 (N_14617,N_13196,N_13833);
nor U14618 (N_14618,N_13697,N_13427);
or U14619 (N_14619,N_13229,N_13827);
and U14620 (N_14620,N_13974,N_13187);
and U14621 (N_14621,N_13132,N_13909);
and U14622 (N_14622,N_13372,N_13455);
or U14623 (N_14623,N_13528,N_13279);
nand U14624 (N_14624,N_13707,N_13678);
nand U14625 (N_14625,N_13490,N_13556);
nor U14626 (N_14626,N_13080,N_13268);
nor U14627 (N_14627,N_13051,N_13945);
nand U14628 (N_14628,N_13801,N_13419);
nor U14629 (N_14629,N_13377,N_13358);
nand U14630 (N_14630,N_13409,N_13479);
xnor U14631 (N_14631,N_13098,N_13534);
or U14632 (N_14632,N_13663,N_13831);
or U14633 (N_14633,N_13326,N_13284);
nor U14634 (N_14634,N_13948,N_13740);
xor U14635 (N_14635,N_13167,N_13747);
and U14636 (N_14636,N_13787,N_13696);
nand U14637 (N_14637,N_13039,N_13665);
nand U14638 (N_14638,N_13273,N_13781);
nor U14639 (N_14639,N_13470,N_13851);
and U14640 (N_14640,N_13510,N_13520);
and U14641 (N_14641,N_13587,N_13405);
nor U14642 (N_14642,N_13484,N_13796);
and U14643 (N_14643,N_13103,N_13122);
or U14644 (N_14644,N_13694,N_13846);
nand U14645 (N_14645,N_13050,N_13836);
xor U14646 (N_14646,N_13815,N_13421);
nor U14647 (N_14647,N_13213,N_13536);
or U14648 (N_14648,N_13506,N_13829);
and U14649 (N_14649,N_13324,N_13207);
and U14650 (N_14650,N_13954,N_13984);
or U14651 (N_14651,N_13626,N_13334);
nor U14652 (N_14652,N_13074,N_13397);
nor U14653 (N_14653,N_13587,N_13617);
and U14654 (N_14654,N_13954,N_13757);
and U14655 (N_14655,N_13546,N_13129);
nor U14656 (N_14656,N_13455,N_13773);
xnor U14657 (N_14657,N_13862,N_13581);
xor U14658 (N_14658,N_13149,N_13265);
and U14659 (N_14659,N_13192,N_13089);
xor U14660 (N_14660,N_13973,N_13858);
nor U14661 (N_14661,N_13901,N_13840);
nor U14662 (N_14662,N_13370,N_13254);
or U14663 (N_14663,N_13291,N_13441);
and U14664 (N_14664,N_13818,N_13247);
nor U14665 (N_14665,N_13888,N_13746);
nor U14666 (N_14666,N_13068,N_13902);
and U14667 (N_14667,N_13159,N_13978);
nor U14668 (N_14668,N_13439,N_13569);
nand U14669 (N_14669,N_13785,N_13284);
or U14670 (N_14670,N_13409,N_13901);
nor U14671 (N_14671,N_13579,N_13839);
xnor U14672 (N_14672,N_13834,N_13766);
and U14673 (N_14673,N_13989,N_13230);
or U14674 (N_14674,N_13434,N_13722);
nor U14675 (N_14675,N_13594,N_13949);
and U14676 (N_14676,N_13714,N_13637);
nand U14677 (N_14677,N_13647,N_13621);
nor U14678 (N_14678,N_13159,N_13720);
xnor U14679 (N_14679,N_13416,N_13538);
nand U14680 (N_14680,N_13867,N_13934);
nor U14681 (N_14681,N_13090,N_13193);
or U14682 (N_14682,N_13398,N_13225);
or U14683 (N_14683,N_13173,N_13823);
xor U14684 (N_14684,N_13236,N_13109);
xnor U14685 (N_14685,N_13009,N_13090);
xor U14686 (N_14686,N_13998,N_13247);
nand U14687 (N_14687,N_13114,N_13422);
nand U14688 (N_14688,N_13400,N_13986);
nor U14689 (N_14689,N_13606,N_13383);
nand U14690 (N_14690,N_13881,N_13136);
and U14691 (N_14691,N_13102,N_13204);
nand U14692 (N_14692,N_13953,N_13321);
nand U14693 (N_14693,N_13764,N_13434);
xnor U14694 (N_14694,N_13317,N_13656);
xnor U14695 (N_14695,N_13519,N_13999);
and U14696 (N_14696,N_13222,N_13131);
or U14697 (N_14697,N_13768,N_13738);
xnor U14698 (N_14698,N_13608,N_13228);
and U14699 (N_14699,N_13420,N_13799);
nand U14700 (N_14700,N_13448,N_13222);
and U14701 (N_14701,N_13759,N_13482);
nand U14702 (N_14702,N_13275,N_13759);
nor U14703 (N_14703,N_13135,N_13096);
nand U14704 (N_14704,N_13326,N_13173);
xnor U14705 (N_14705,N_13579,N_13683);
nor U14706 (N_14706,N_13373,N_13047);
and U14707 (N_14707,N_13710,N_13240);
nor U14708 (N_14708,N_13235,N_13408);
and U14709 (N_14709,N_13981,N_13072);
xor U14710 (N_14710,N_13481,N_13939);
nand U14711 (N_14711,N_13764,N_13738);
nand U14712 (N_14712,N_13825,N_13623);
or U14713 (N_14713,N_13988,N_13610);
or U14714 (N_14714,N_13054,N_13295);
nand U14715 (N_14715,N_13513,N_13597);
xnor U14716 (N_14716,N_13392,N_13880);
and U14717 (N_14717,N_13073,N_13296);
or U14718 (N_14718,N_13779,N_13901);
or U14719 (N_14719,N_13522,N_13592);
nor U14720 (N_14720,N_13921,N_13481);
or U14721 (N_14721,N_13233,N_13973);
nand U14722 (N_14722,N_13054,N_13215);
xnor U14723 (N_14723,N_13131,N_13235);
xor U14724 (N_14724,N_13075,N_13462);
and U14725 (N_14725,N_13001,N_13997);
nor U14726 (N_14726,N_13416,N_13156);
xnor U14727 (N_14727,N_13160,N_13787);
nor U14728 (N_14728,N_13782,N_13221);
xnor U14729 (N_14729,N_13646,N_13109);
nand U14730 (N_14730,N_13920,N_13784);
and U14731 (N_14731,N_13692,N_13931);
nand U14732 (N_14732,N_13492,N_13079);
and U14733 (N_14733,N_13233,N_13428);
nand U14734 (N_14734,N_13733,N_13443);
and U14735 (N_14735,N_13930,N_13956);
and U14736 (N_14736,N_13501,N_13802);
xor U14737 (N_14737,N_13740,N_13034);
nor U14738 (N_14738,N_13562,N_13564);
xor U14739 (N_14739,N_13156,N_13594);
or U14740 (N_14740,N_13605,N_13031);
xor U14741 (N_14741,N_13110,N_13630);
nand U14742 (N_14742,N_13446,N_13474);
nor U14743 (N_14743,N_13695,N_13119);
xnor U14744 (N_14744,N_13764,N_13873);
or U14745 (N_14745,N_13082,N_13163);
nand U14746 (N_14746,N_13411,N_13770);
or U14747 (N_14747,N_13269,N_13968);
or U14748 (N_14748,N_13305,N_13572);
or U14749 (N_14749,N_13703,N_13070);
xor U14750 (N_14750,N_13005,N_13153);
nor U14751 (N_14751,N_13362,N_13262);
xor U14752 (N_14752,N_13658,N_13437);
or U14753 (N_14753,N_13464,N_13866);
nor U14754 (N_14754,N_13722,N_13963);
xor U14755 (N_14755,N_13879,N_13404);
or U14756 (N_14756,N_13598,N_13477);
or U14757 (N_14757,N_13043,N_13791);
or U14758 (N_14758,N_13988,N_13391);
and U14759 (N_14759,N_13473,N_13331);
or U14760 (N_14760,N_13394,N_13724);
nand U14761 (N_14761,N_13942,N_13102);
nand U14762 (N_14762,N_13260,N_13514);
nand U14763 (N_14763,N_13859,N_13357);
or U14764 (N_14764,N_13117,N_13539);
nand U14765 (N_14765,N_13634,N_13581);
and U14766 (N_14766,N_13534,N_13297);
xnor U14767 (N_14767,N_13606,N_13496);
and U14768 (N_14768,N_13542,N_13442);
nand U14769 (N_14769,N_13113,N_13329);
xnor U14770 (N_14770,N_13071,N_13459);
xnor U14771 (N_14771,N_13560,N_13869);
or U14772 (N_14772,N_13917,N_13228);
xnor U14773 (N_14773,N_13092,N_13338);
xor U14774 (N_14774,N_13270,N_13051);
or U14775 (N_14775,N_13368,N_13914);
nor U14776 (N_14776,N_13827,N_13543);
or U14777 (N_14777,N_13421,N_13576);
or U14778 (N_14778,N_13368,N_13653);
and U14779 (N_14779,N_13850,N_13322);
and U14780 (N_14780,N_13326,N_13447);
nand U14781 (N_14781,N_13194,N_13685);
nor U14782 (N_14782,N_13213,N_13856);
nor U14783 (N_14783,N_13693,N_13006);
nor U14784 (N_14784,N_13618,N_13600);
or U14785 (N_14785,N_13681,N_13553);
nor U14786 (N_14786,N_13786,N_13935);
nand U14787 (N_14787,N_13364,N_13309);
xnor U14788 (N_14788,N_13788,N_13344);
xor U14789 (N_14789,N_13125,N_13743);
and U14790 (N_14790,N_13996,N_13218);
and U14791 (N_14791,N_13905,N_13984);
or U14792 (N_14792,N_13135,N_13113);
nor U14793 (N_14793,N_13427,N_13030);
nor U14794 (N_14794,N_13902,N_13292);
nor U14795 (N_14795,N_13349,N_13763);
and U14796 (N_14796,N_13108,N_13451);
nand U14797 (N_14797,N_13535,N_13501);
or U14798 (N_14798,N_13661,N_13806);
or U14799 (N_14799,N_13527,N_13033);
xor U14800 (N_14800,N_13288,N_13550);
and U14801 (N_14801,N_13529,N_13797);
and U14802 (N_14802,N_13212,N_13157);
and U14803 (N_14803,N_13217,N_13615);
nand U14804 (N_14804,N_13256,N_13179);
nand U14805 (N_14805,N_13651,N_13687);
nand U14806 (N_14806,N_13439,N_13172);
or U14807 (N_14807,N_13022,N_13784);
nor U14808 (N_14808,N_13268,N_13670);
and U14809 (N_14809,N_13356,N_13299);
nand U14810 (N_14810,N_13835,N_13748);
nor U14811 (N_14811,N_13894,N_13922);
nor U14812 (N_14812,N_13232,N_13586);
xnor U14813 (N_14813,N_13087,N_13658);
or U14814 (N_14814,N_13771,N_13702);
nand U14815 (N_14815,N_13819,N_13842);
xor U14816 (N_14816,N_13865,N_13770);
or U14817 (N_14817,N_13770,N_13664);
xnor U14818 (N_14818,N_13076,N_13583);
and U14819 (N_14819,N_13962,N_13488);
nand U14820 (N_14820,N_13880,N_13729);
xnor U14821 (N_14821,N_13807,N_13814);
xor U14822 (N_14822,N_13792,N_13555);
nand U14823 (N_14823,N_13855,N_13349);
or U14824 (N_14824,N_13072,N_13324);
nand U14825 (N_14825,N_13625,N_13252);
nand U14826 (N_14826,N_13714,N_13234);
nor U14827 (N_14827,N_13920,N_13506);
and U14828 (N_14828,N_13004,N_13966);
nand U14829 (N_14829,N_13931,N_13907);
nor U14830 (N_14830,N_13580,N_13533);
xnor U14831 (N_14831,N_13995,N_13456);
or U14832 (N_14832,N_13086,N_13081);
and U14833 (N_14833,N_13986,N_13407);
xnor U14834 (N_14834,N_13406,N_13607);
xor U14835 (N_14835,N_13848,N_13907);
and U14836 (N_14836,N_13452,N_13470);
xor U14837 (N_14837,N_13812,N_13132);
nand U14838 (N_14838,N_13891,N_13936);
nand U14839 (N_14839,N_13519,N_13981);
nor U14840 (N_14840,N_13863,N_13229);
or U14841 (N_14841,N_13931,N_13727);
or U14842 (N_14842,N_13191,N_13579);
xor U14843 (N_14843,N_13547,N_13969);
and U14844 (N_14844,N_13979,N_13278);
nor U14845 (N_14845,N_13728,N_13606);
and U14846 (N_14846,N_13999,N_13911);
nor U14847 (N_14847,N_13009,N_13058);
xnor U14848 (N_14848,N_13845,N_13807);
and U14849 (N_14849,N_13653,N_13388);
nand U14850 (N_14850,N_13486,N_13232);
nor U14851 (N_14851,N_13575,N_13327);
nand U14852 (N_14852,N_13132,N_13110);
nor U14853 (N_14853,N_13923,N_13690);
xnor U14854 (N_14854,N_13433,N_13248);
xor U14855 (N_14855,N_13960,N_13946);
xor U14856 (N_14856,N_13843,N_13570);
nand U14857 (N_14857,N_13701,N_13240);
nor U14858 (N_14858,N_13279,N_13859);
xor U14859 (N_14859,N_13030,N_13673);
nand U14860 (N_14860,N_13404,N_13867);
or U14861 (N_14861,N_13777,N_13358);
and U14862 (N_14862,N_13578,N_13636);
or U14863 (N_14863,N_13889,N_13106);
xnor U14864 (N_14864,N_13354,N_13337);
and U14865 (N_14865,N_13529,N_13349);
nand U14866 (N_14866,N_13030,N_13269);
nand U14867 (N_14867,N_13606,N_13202);
xnor U14868 (N_14868,N_13146,N_13157);
or U14869 (N_14869,N_13092,N_13680);
nand U14870 (N_14870,N_13795,N_13042);
nand U14871 (N_14871,N_13367,N_13552);
nand U14872 (N_14872,N_13141,N_13473);
xor U14873 (N_14873,N_13546,N_13265);
nand U14874 (N_14874,N_13435,N_13087);
xor U14875 (N_14875,N_13551,N_13635);
xor U14876 (N_14876,N_13764,N_13931);
nand U14877 (N_14877,N_13763,N_13663);
and U14878 (N_14878,N_13375,N_13099);
and U14879 (N_14879,N_13525,N_13852);
nand U14880 (N_14880,N_13668,N_13356);
nor U14881 (N_14881,N_13455,N_13550);
or U14882 (N_14882,N_13249,N_13484);
or U14883 (N_14883,N_13247,N_13316);
and U14884 (N_14884,N_13781,N_13701);
nand U14885 (N_14885,N_13930,N_13727);
or U14886 (N_14886,N_13404,N_13896);
or U14887 (N_14887,N_13063,N_13210);
xnor U14888 (N_14888,N_13372,N_13430);
and U14889 (N_14889,N_13193,N_13368);
or U14890 (N_14890,N_13077,N_13037);
or U14891 (N_14891,N_13044,N_13296);
nand U14892 (N_14892,N_13300,N_13568);
xnor U14893 (N_14893,N_13324,N_13288);
xnor U14894 (N_14894,N_13334,N_13014);
nand U14895 (N_14895,N_13428,N_13810);
nand U14896 (N_14896,N_13436,N_13760);
nor U14897 (N_14897,N_13949,N_13514);
and U14898 (N_14898,N_13691,N_13826);
and U14899 (N_14899,N_13143,N_13576);
or U14900 (N_14900,N_13023,N_13968);
and U14901 (N_14901,N_13493,N_13957);
and U14902 (N_14902,N_13265,N_13879);
or U14903 (N_14903,N_13855,N_13371);
nor U14904 (N_14904,N_13212,N_13680);
and U14905 (N_14905,N_13942,N_13885);
xor U14906 (N_14906,N_13581,N_13128);
and U14907 (N_14907,N_13730,N_13357);
nor U14908 (N_14908,N_13174,N_13328);
nand U14909 (N_14909,N_13698,N_13898);
nand U14910 (N_14910,N_13189,N_13033);
xor U14911 (N_14911,N_13502,N_13029);
xnor U14912 (N_14912,N_13886,N_13905);
nor U14913 (N_14913,N_13139,N_13599);
or U14914 (N_14914,N_13325,N_13699);
or U14915 (N_14915,N_13684,N_13712);
nand U14916 (N_14916,N_13462,N_13094);
and U14917 (N_14917,N_13285,N_13086);
nor U14918 (N_14918,N_13256,N_13324);
and U14919 (N_14919,N_13393,N_13184);
or U14920 (N_14920,N_13093,N_13183);
and U14921 (N_14921,N_13768,N_13592);
xor U14922 (N_14922,N_13477,N_13889);
nor U14923 (N_14923,N_13267,N_13943);
or U14924 (N_14924,N_13363,N_13137);
nor U14925 (N_14925,N_13443,N_13216);
or U14926 (N_14926,N_13542,N_13529);
nand U14927 (N_14927,N_13920,N_13328);
xor U14928 (N_14928,N_13961,N_13093);
nand U14929 (N_14929,N_13371,N_13512);
xor U14930 (N_14930,N_13640,N_13687);
nand U14931 (N_14931,N_13949,N_13777);
and U14932 (N_14932,N_13628,N_13413);
nand U14933 (N_14933,N_13849,N_13758);
nor U14934 (N_14934,N_13813,N_13340);
nor U14935 (N_14935,N_13653,N_13425);
nand U14936 (N_14936,N_13077,N_13275);
or U14937 (N_14937,N_13199,N_13836);
and U14938 (N_14938,N_13296,N_13138);
xor U14939 (N_14939,N_13121,N_13050);
nand U14940 (N_14940,N_13013,N_13324);
and U14941 (N_14941,N_13570,N_13699);
and U14942 (N_14942,N_13209,N_13502);
nand U14943 (N_14943,N_13112,N_13907);
nand U14944 (N_14944,N_13780,N_13984);
nor U14945 (N_14945,N_13585,N_13519);
nand U14946 (N_14946,N_13354,N_13153);
xor U14947 (N_14947,N_13836,N_13999);
nand U14948 (N_14948,N_13224,N_13034);
and U14949 (N_14949,N_13931,N_13493);
nor U14950 (N_14950,N_13730,N_13543);
and U14951 (N_14951,N_13079,N_13452);
and U14952 (N_14952,N_13945,N_13448);
nor U14953 (N_14953,N_13552,N_13273);
xor U14954 (N_14954,N_13847,N_13677);
nand U14955 (N_14955,N_13627,N_13466);
and U14956 (N_14956,N_13054,N_13200);
and U14957 (N_14957,N_13660,N_13175);
nor U14958 (N_14958,N_13424,N_13230);
or U14959 (N_14959,N_13390,N_13763);
nor U14960 (N_14960,N_13380,N_13935);
nor U14961 (N_14961,N_13164,N_13451);
and U14962 (N_14962,N_13557,N_13609);
nor U14963 (N_14963,N_13313,N_13057);
nor U14964 (N_14964,N_13248,N_13336);
nand U14965 (N_14965,N_13992,N_13855);
xnor U14966 (N_14966,N_13676,N_13232);
or U14967 (N_14967,N_13267,N_13054);
or U14968 (N_14968,N_13380,N_13255);
and U14969 (N_14969,N_13909,N_13238);
nand U14970 (N_14970,N_13417,N_13207);
nor U14971 (N_14971,N_13675,N_13998);
or U14972 (N_14972,N_13662,N_13593);
and U14973 (N_14973,N_13564,N_13846);
or U14974 (N_14974,N_13732,N_13751);
nand U14975 (N_14975,N_13374,N_13413);
or U14976 (N_14976,N_13231,N_13529);
xnor U14977 (N_14977,N_13998,N_13116);
nor U14978 (N_14978,N_13840,N_13866);
xnor U14979 (N_14979,N_13657,N_13039);
xor U14980 (N_14980,N_13368,N_13287);
nand U14981 (N_14981,N_13621,N_13509);
nor U14982 (N_14982,N_13339,N_13859);
or U14983 (N_14983,N_13453,N_13480);
or U14984 (N_14984,N_13159,N_13807);
nand U14985 (N_14985,N_13464,N_13163);
and U14986 (N_14986,N_13067,N_13012);
nor U14987 (N_14987,N_13343,N_13105);
xnor U14988 (N_14988,N_13586,N_13659);
or U14989 (N_14989,N_13231,N_13850);
xnor U14990 (N_14990,N_13983,N_13546);
nand U14991 (N_14991,N_13163,N_13545);
nor U14992 (N_14992,N_13757,N_13468);
xnor U14993 (N_14993,N_13292,N_13409);
xor U14994 (N_14994,N_13347,N_13026);
nor U14995 (N_14995,N_13224,N_13410);
xor U14996 (N_14996,N_13583,N_13597);
nor U14997 (N_14997,N_13108,N_13892);
xor U14998 (N_14998,N_13241,N_13695);
and U14999 (N_14999,N_13128,N_13422);
nor U15000 (N_15000,N_14584,N_14282);
nand U15001 (N_15001,N_14905,N_14109);
nand U15002 (N_15002,N_14654,N_14438);
and U15003 (N_15003,N_14789,N_14658);
nor U15004 (N_15004,N_14195,N_14866);
or U15005 (N_15005,N_14279,N_14451);
nand U15006 (N_15006,N_14168,N_14842);
and U15007 (N_15007,N_14000,N_14064);
and U15008 (N_15008,N_14904,N_14704);
nand U15009 (N_15009,N_14854,N_14865);
and U15010 (N_15010,N_14699,N_14399);
nand U15011 (N_15011,N_14370,N_14656);
nand U15012 (N_15012,N_14734,N_14456);
nand U15013 (N_15013,N_14809,N_14986);
xor U15014 (N_15014,N_14479,N_14029);
and U15015 (N_15015,N_14291,N_14690);
xor U15016 (N_15016,N_14600,N_14055);
and U15017 (N_15017,N_14929,N_14803);
and U15018 (N_15018,N_14048,N_14397);
xor U15019 (N_15019,N_14092,N_14976);
and U15020 (N_15020,N_14042,N_14559);
nand U15021 (N_15021,N_14806,N_14616);
or U15022 (N_15022,N_14820,N_14705);
nor U15023 (N_15023,N_14623,N_14535);
or U15024 (N_15024,N_14878,N_14469);
nand U15025 (N_15025,N_14999,N_14298);
xnor U15026 (N_15026,N_14326,N_14108);
nand U15027 (N_15027,N_14828,N_14489);
xnor U15028 (N_15028,N_14744,N_14271);
nand U15029 (N_15029,N_14299,N_14977);
or U15030 (N_15030,N_14363,N_14194);
or U15031 (N_15031,N_14421,N_14202);
or U15032 (N_15032,N_14918,N_14991);
and U15033 (N_15033,N_14831,N_14761);
nor U15034 (N_15034,N_14107,N_14666);
and U15035 (N_15035,N_14180,N_14963);
nor U15036 (N_15036,N_14182,N_14898);
or U15037 (N_15037,N_14056,N_14464);
nand U15038 (N_15038,N_14151,N_14773);
nor U15039 (N_15039,N_14375,N_14333);
and U15040 (N_15040,N_14780,N_14241);
nand U15041 (N_15041,N_14113,N_14617);
and U15042 (N_15042,N_14433,N_14070);
xor U15043 (N_15043,N_14852,N_14590);
or U15044 (N_15044,N_14261,N_14077);
or U15045 (N_15045,N_14344,N_14133);
and U15046 (N_15046,N_14791,N_14971);
and U15047 (N_15047,N_14651,N_14418);
nand U15048 (N_15048,N_14013,N_14412);
or U15049 (N_15049,N_14150,N_14829);
or U15050 (N_15050,N_14115,N_14609);
xnor U15051 (N_15051,N_14622,N_14085);
or U15052 (N_15052,N_14642,N_14360);
nand U15053 (N_15053,N_14844,N_14361);
nand U15054 (N_15054,N_14557,N_14275);
nor U15055 (N_15055,N_14355,N_14367);
nand U15056 (N_15056,N_14309,N_14737);
xor U15057 (N_15057,N_14119,N_14340);
or U15058 (N_15058,N_14942,N_14447);
xor U15059 (N_15059,N_14619,N_14722);
or U15060 (N_15060,N_14288,N_14516);
nor U15061 (N_15061,N_14439,N_14634);
nand U15062 (N_15062,N_14745,N_14927);
and U15063 (N_15063,N_14206,N_14838);
nor U15064 (N_15064,N_14330,N_14718);
and U15065 (N_15065,N_14346,N_14243);
and U15066 (N_15066,N_14037,N_14318);
nor U15067 (N_15067,N_14294,N_14964);
nor U15068 (N_15068,N_14967,N_14117);
nand U15069 (N_15069,N_14235,N_14205);
nor U15070 (N_15070,N_14242,N_14802);
or U15071 (N_15071,N_14143,N_14824);
xnor U15072 (N_15072,N_14930,N_14511);
and U15073 (N_15073,N_14125,N_14250);
nor U15074 (N_15074,N_14139,N_14425);
xor U15075 (N_15075,N_14747,N_14371);
and U15076 (N_15076,N_14601,N_14922);
nor U15077 (N_15077,N_14572,N_14214);
nor U15078 (N_15078,N_14138,N_14075);
xor U15079 (N_15079,N_14548,N_14532);
and U15080 (N_15080,N_14515,N_14233);
nand U15081 (N_15081,N_14045,N_14210);
and U15082 (N_15082,N_14493,N_14017);
and U15083 (N_15083,N_14675,N_14380);
nor U15084 (N_15084,N_14952,N_14307);
nor U15085 (N_15085,N_14627,N_14174);
or U15086 (N_15086,N_14767,N_14568);
nand U15087 (N_15087,N_14413,N_14506);
and U15088 (N_15088,N_14453,N_14083);
xnor U15089 (N_15089,N_14207,N_14980);
nor U15090 (N_15090,N_14801,N_14006);
xnor U15091 (N_15091,N_14173,N_14677);
nor U15092 (N_15092,N_14522,N_14847);
or U15093 (N_15093,N_14219,N_14259);
xnor U15094 (N_15094,N_14782,N_14751);
or U15095 (N_15095,N_14834,N_14420);
and U15096 (N_15096,N_14653,N_14742);
nor U15097 (N_15097,N_14434,N_14303);
xor U15098 (N_15098,N_14902,N_14545);
or U15099 (N_15099,N_14059,N_14962);
or U15100 (N_15100,N_14758,N_14714);
nand U15101 (N_15101,N_14474,N_14321);
or U15102 (N_15102,N_14983,N_14179);
and U15103 (N_15103,N_14289,N_14381);
or U15104 (N_15104,N_14644,N_14222);
and U15105 (N_15105,N_14940,N_14050);
and U15106 (N_15106,N_14430,N_14931);
or U15107 (N_15107,N_14657,N_14337);
or U15108 (N_15108,N_14953,N_14002);
nor U15109 (N_15109,N_14351,N_14992);
nand U15110 (N_15110,N_14188,N_14081);
and U15111 (N_15111,N_14156,N_14629);
nand U15112 (N_15112,N_14273,N_14229);
or U15113 (N_15113,N_14883,N_14533);
nand U15114 (N_15114,N_14163,N_14888);
and U15115 (N_15115,N_14018,N_14246);
nand U15116 (N_15116,N_14350,N_14890);
or U15117 (N_15117,N_14571,N_14165);
nor U15118 (N_15118,N_14404,N_14814);
and U15119 (N_15119,N_14885,N_14638);
nand U15120 (N_15120,N_14621,N_14662);
and U15121 (N_15121,N_14448,N_14015);
nand U15122 (N_15122,N_14477,N_14353);
xnor U15123 (N_15123,N_14014,N_14567);
xor U15124 (N_15124,N_14216,N_14785);
nor U15125 (N_15125,N_14924,N_14341);
or U15126 (N_15126,N_14668,N_14221);
nand U15127 (N_15127,N_14892,N_14848);
and U15128 (N_15128,N_14843,N_14851);
nor U15129 (N_15129,N_14035,N_14939);
nor U15130 (N_15130,N_14480,N_14716);
and U15131 (N_15131,N_14209,N_14463);
xor U15132 (N_15132,N_14120,N_14011);
nor U15133 (N_15133,N_14440,N_14470);
nor U15134 (N_15134,N_14449,N_14605);
and U15135 (N_15135,N_14135,N_14252);
and U15136 (N_15136,N_14041,N_14523);
and U15137 (N_15137,N_14850,N_14706);
and U15138 (N_15138,N_14428,N_14912);
xor U15139 (N_15139,N_14228,N_14023);
and U15140 (N_15140,N_14503,N_14102);
nand U15141 (N_15141,N_14673,N_14756);
and U15142 (N_15142,N_14260,N_14944);
or U15143 (N_15143,N_14938,N_14682);
nor U15144 (N_15144,N_14712,N_14123);
nand U15145 (N_15145,N_14383,N_14359);
nand U15146 (N_15146,N_14274,N_14155);
and U15147 (N_15147,N_14869,N_14840);
xor U15148 (N_15148,N_14272,N_14721);
or U15149 (N_15149,N_14646,N_14226);
nand U15150 (N_15150,N_14454,N_14431);
nor U15151 (N_15151,N_14204,N_14192);
and U15152 (N_15152,N_14717,N_14588);
or U15153 (N_15153,N_14184,N_14429);
xnor U15154 (N_15154,N_14507,N_14066);
or U15155 (N_15155,N_14100,N_14741);
and U15156 (N_15156,N_14845,N_14103);
nor U15157 (N_15157,N_14001,N_14458);
xor U15158 (N_15158,N_14599,N_14937);
xnor U15159 (N_15159,N_14777,N_14074);
and U15160 (N_15160,N_14961,N_14762);
nand U15161 (N_15161,N_14604,N_14364);
and U15162 (N_15162,N_14876,N_14794);
or U15163 (N_15163,N_14234,N_14864);
nor U15164 (N_15164,N_14024,N_14973);
nand U15165 (N_15165,N_14089,N_14916);
and U15166 (N_15166,N_14552,N_14293);
and U15167 (N_15167,N_14862,N_14262);
xor U15168 (N_15168,N_14612,N_14643);
nand U15169 (N_15169,N_14324,N_14020);
nor U15170 (N_15170,N_14191,N_14415);
or U15171 (N_15171,N_14147,N_14435);
and U15172 (N_15172,N_14499,N_14417);
nand U15173 (N_15173,N_14392,N_14157);
xnor U15174 (N_15174,N_14543,N_14894);
xor U15175 (N_15175,N_14594,N_14466);
xor U15176 (N_15176,N_14678,N_14054);
nor U15177 (N_15177,N_14396,N_14684);
or U15178 (N_15178,N_14031,N_14365);
xnor U15179 (N_15179,N_14224,N_14086);
nor U15180 (N_15180,N_14713,N_14492);
and U15181 (N_15181,N_14422,N_14240);
nor U15182 (N_15182,N_14748,N_14573);
xor U15183 (N_15183,N_14674,N_14387);
xor U15184 (N_15184,N_14671,N_14827);
xnor U15185 (N_15185,N_14841,N_14798);
xor U15186 (N_15186,N_14302,N_14542);
nor U15187 (N_15187,N_14078,N_14790);
and U15188 (N_15188,N_14026,N_14591);
or U15189 (N_15189,N_14659,N_14546);
or U15190 (N_15190,N_14561,N_14719);
nor U15191 (N_15191,N_14197,N_14036);
xnor U15192 (N_15192,N_14193,N_14911);
and U15193 (N_15193,N_14424,N_14951);
xnor U15194 (N_15194,N_14407,N_14322);
xor U15195 (N_15195,N_14183,N_14948);
nand U15196 (N_15196,N_14076,N_14781);
nor U15197 (N_15197,N_14304,N_14501);
and U15198 (N_15198,N_14832,N_14129);
and U15199 (N_15199,N_14636,N_14907);
or U15200 (N_15200,N_14839,N_14116);
nand U15201 (N_15201,N_14121,N_14130);
nand U15202 (N_15202,N_14947,N_14702);
xor U15203 (N_15203,N_14372,N_14171);
xor U15204 (N_15204,N_14258,N_14158);
nor U15205 (N_15205,N_14645,N_14826);
and U15206 (N_15206,N_14534,N_14080);
nand U15207 (N_15207,N_14032,N_14319);
or U15208 (N_15208,N_14140,N_14393);
nor U15209 (N_15209,N_14185,N_14459);
or U15210 (N_15210,N_14539,N_14283);
and U15211 (N_15211,N_14595,N_14386);
or U15212 (N_15212,N_14873,N_14253);
and U15213 (N_15213,N_14549,N_14169);
xor U15214 (N_15214,N_14491,N_14889);
and U15215 (N_15215,N_14989,N_14073);
and U15216 (N_15216,N_14725,N_14146);
xor U15217 (N_15217,N_14886,N_14486);
nor U15218 (N_15218,N_14028,N_14517);
nand U15219 (N_15219,N_14943,N_14765);
xnor U15220 (N_15220,N_14112,N_14606);
nor U15221 (N_15221,N_14587,N_14932);
xor U15222 (N_15222,N_14484,N_14596);
nor U15223 (N_15223,N_14731,N_14611);
or U15224 (N_15224,N_14166,N_14749);
nor U15225 (N_15225,N_14019,N_14715);
nand U15226 (N_15226,N_14007,N_14558);
and U15227 (N_15227,N_14555,N_14471);
nand U15228 (N_15228,N_14368,N_14170);
nor U15229 (N_15229,N_14703,N_14728);
nor U15230 (N_15230,N_14053,N_14483);
xor U15231 (N_15231,N_14536,N_14597);
and U15232 (N_15232,N_14452,N_14118);
nor U15233 (N_15233,N_14954,N_14342);
nand U15234 (N_15234,N_14087,N_14084);
or U15235 (N_15235,N_14547,N_14095);
and U15236 (N_15236,N_14974,N_14488);
nand U15237 (N_15237,N_14910,N_14349);
nor U15238 (N_15238,N_14046,N_14735);
and U15239 (N_15239,N_14215,N_14290);
or U15240 (N_15240,N_14966,N_14540);
xnor U15241 (N_15241,N_14317,N_14090);
xnor U15242 (N_15242,N_14105,N_14004);
nor U15243 (N_15243,N_14723,N_14186);
nand U15244 (N_15244,N_14720,N_14960);
and U15245 (N_15245,N_14338,N_14040);
and U15246 (N_15246,N_14859,N_14237);
and U15247 (N_15247,N_14647,N_14855);
nor U15248 (N_15248,N_14799,N_14267);
nand U15249 (N_15249,N_14835,N_14443);
xor U15250 (N_15250,N_14891,N_14683);
or U15251 (N_15251,N_14672,N_14804);
nor U15252 (N_15252,N_14411,N_14232);
xnor U15253 (N_15253,N_14097,N_14959);
nor U15254 (N_15254,N_14154,N_14467);
nand U15255 (N_15255,N_14524,N_14010);
nand U15256 (N_15256,N_14212,N_14352);
and U15257 (N_15257,N_14265,N_14061);
or U15258 (N_15258,N_14500,N_14926);
nor U15259 (N_15259,N_14776,N_14822);
nor U15260 (N_15260,N_14856,N_14336);
nand U15261 (N_15261,N_14389,N_14475);
and U15262 (N_15262,N_14689,N_14867);
and U15263 (N_15263,N_14378,N_14920);
and U15264 (N_15264,N_14661,N_14465);
nand U15265 (N_15265,N_14498,N_14200);
or U15266 (N_15266,N_14710,N_14917);
nand U15267 (N_15267,N_14268,N_14903);
nand U15268 (N_15268,N_14377,N_14313);
nor U15269 (N_15269,N_14223,N_14199);
or U15270 (N_15270,N_14863,N_14257);
or U15271 (N_15271,N_14247,N_14494);
xor U15272 (N_15272,N_14805,N_14630);
and U15273 (N_15273,N_14476,N_14461);
nand U15274 (N_15274,N_14110,N_14314);
and U15275 (N_15275,N_14795,N_14187);
and U15276 (N_15276,N_14400,N_14663);
or U15277 (N_15277,N_14472,N_14356);
xnor U15278 (N_15278,N_14022,N_14641);
nor U15279 (N_15279,N_14774,N_14667);
nand U15280 (N_15280,N_14877,N_14172);
nand U15281 (N_15281,N_14057,N_14857);
and U15282 (N_15282,N_14906,N_14047);
and U15283 (N_15283,N_14764,N_14589);
or U15284 (N_15284,N_14733,N_14519);
nor U15285 (N_15285,N_14949,N_14408);
or U15286 (N_15286,N_14152,N_14382);
nand U15287 (N_15287,N_14039,N_14044);
nand U15288 (N_15288,N_14414,N_14784);
nor U15289 (N_15289,N_14320,N_14132);
xnor U15290 (N_15290,N_14496,N_14769);
and U15291 (N_15291,N_14525,N_14460);
xor U15292 (N_15292,N_14513,N_14264);
or U15293 (N_15293,N_14993,N_14608);
xnor U15294 (N_15294,N_14763,N_14306);
xor U15295 (N_15295,N_14148,N_14021);
nand U15296 (N_15296,N_14965,N_14141);
nand U15297 (N_15297,N_14373,N_14779);
nor U15298 (N_15298,N_14520,N_14175);
and U15299 (N_15299,N_14950,N_14553);
xnor U15300 (N_15300,N_14398,N_14094);
nand U15301 (N_15301,N_14227,N_14391);
nand U15302 (N_15302,N_14946,N_14681);
and U15303 (N_15303,N_14676,N_14550);
or U15304 (N_15304,N_14565,N_14305);
and U15305 (N_15305,N_14560,N_14694);
nor U15306 (N_15306,N_14446,N_14490);
xor U15307 (N_15307,N_14664,N_14755);
and U15308 (N_15308,N_14575,N_14285);
and U15309 (N_15309,N_14708,N_14248);
xnor U15310 (N_15310,N_14379,N_14481);
or U15311 (N_15311,N_14921,N_14928);
nand U15312 (N_15312,N_14376,N_14374);
nand U15313 (N_15313,N_14698,N_14692);
nor U15314 (N_15314,N_14582,N_14104);
nand U15315 (N_15315,N_14908,N_14727);
nor U15316 (N_15316,N_14062,N_14730);
nand U15317 (N_15317,N_14065,N_14402);
xnor U15318 (N_15318,N_14091,N_14615);
xor U15319 (N_15319,N_14786,N_14310);
xnor U15320 (N_15320,N_14278,N_14697);
nor U15321 (N_15321,N_14846,N_14203);
or U15322 (N_15322,N_14334,N_14537);
and U15323 (N_15323,N_14693,N_14280);
and U15324 (N_15324,N_14236,N_14137);
and U15325 (N_15325,N_14300,N_14518);
xnor U15326 (N_15326,N_14406,N_14551);
nand U15327 (N_15327,N_14362,N_14628);
or U15328 (N_15328,N_14729,N_14936);
nor U15329 (N_15329,N_14872,N_14711);
xnor U15330 (N_15330,N_14860,N_14580);
or U15331 (N_15331,N_14098,N_14998);
and U15332 (N_15332,N_14388,N_14159);
xnor U15333 (N_15333,N_14450,N_14201);
and U15334 (N_15334,N_14957,N_14189);
and U15335 (N_15335,N_14879,N_14923);
or U15336 (N_15336,N_14444,N_14256);
or U15337 (N_15337,N_14301,N_14161);
or U15338 (N_15338,N_14625,N_14984);
or U15339 (N_15339,N_14836,N_14660);
and U15340 (N_15340,N_14049,N_14255);
nand U15341 (N_15341,N_14919,N_14823);
nor U15342 (N_15342,N_14316,N_14632);
xnor U15343 (N_15343,N_14160,N_14251);
nor U15344 (N_15344,N_14030,N_14401);
nand U15345 (N_15345,N_14178,N_14566);
or U15346 (N_15346,N_14423,N_14585);
nand U15347 (N_15347,N_14153,N_14487);
nor U15348 (N_15348,N_14686,N_14167);
and U15349 (N_15349,N_14384,N_14956);
nor U15350 (N_15350,N_14882,N_14410);
and U15351 (N_15351,N_14685,N_14136);
and U15352 (N_15352,N_14972,N_14441);
nand U15353 (N_15353,N_14270,N_14812);
nor U15354 (N_15354,N_14564,N_14357);
xor U15355 (N_15355,N_14696,N_14164);
nor U15356 (N_15356,N_14510,N_14997);
nor U15357 (N_15357,N_14995,N_14088);
nor U15358 (N_15358,N_14740,N_14009);
nand U15359 (N_15359,N_14881,N_14987);
or U15360 (N_15360,N_14071,N_14849);
or U15361 (N_15361,N_14933,N_14707);
nand U15362 (N_15362,N_14544,N_14695);
and U15363 (N_15363,N_14114,N_14008);
xor U15364 (N_15364,N_14655,N_14665);
and U15365 (N_15365,N_14620,N_14060);
and U15366 (N_15366,N_14868,N_14315);
xnor U15367 (N_15367,N_14016,N_14286);
nor U15368 (N_15368,N_14126,N_14874);
nor U15369 (N_15369,N_14211,N_14145);
nand U15370 (N_15370,N_14586,N_14482);
xor U15371 (N_15371,N_14810,N_14277);
and U15372 (N_15372,N_14754,N_14648);
nor U15373 (N_15373,N_14502,N_14578);
nand U15374 (N_15374,N_14871,N_14770);
nand U15375 (N_15375,N_14052,N_14230);
nor U15376 (N_15376,N_14649,N_14759);
or U15377 (N_15377,N_14614,N_14436);
xor U15378 (N_15378,N_14680,N_14875);
nor U15379 (N_15379,N_14082,N_14577);
xor U15380 (N_15380,N_14732,N_14395);
and U15381 (N_15381,N_14245,N_14249);
xor U15382 (N_15382,N_14527,N_14468);
and U15383 (N_15383,N_14811,N_14366);
nand U15384 (N_15384,N_14347,N_14101);
nor U15385 (N_15385,N_14909,N_14941);
xor U15386 (N_15386,N_14297,N_14994);
and U15387 (N_15387,N_14816,N_14331);
nand U15388 (N_15388,N_14478,N_14354);
or U15389 (N_15389,N_14739,N_14602);
nor U15390 (N_15390,N_14043,N_14473);
nand U15391 (N_15391,N_14244,N_14530);
or U15392 (N_15392,N_14462,N_14508);
nand U15393 (N_15393,N_14531,N_14409);
nand U15394 (N_15394,N_14106,N_14012);
nor U15395 (N_15395,N_14914,N_14217);
or U15396 (N_15396,N_14269,N_14896);
nor U15397 (N_15397,N_14603,N_14162);
nand U15398 (N_15398,N_14514,N_14815);
or U15399 (N_15399,N_14072,N_14807);
or U15400 (N_15400,N_14724,N_14529);
xnor U15401 (N_15401,N_14752,N_14311);
nor U15402 (N_15402,N_14526,N_14208);
nand U15403 (N_15403,N_14198,N_14281);
xnor U15404 (N_15404,N_14335,N_14284);
and U15405 (N_15405,N_14419,N_14554);
nand U15406 (N_15406,N_14025,N_14981);
nand U15407 (N_15407,N_14633,N_14295);
and U15408 (N_15408,N_14339,N_14652);
and U15409 (N_15409,N_14593,N_14969);
xor U15410 (N_15410,N_14427,N_14127);
or U15411 (N_15411,N_14821,N_14058);
xor U15412 (N_15412,N_14687,N_14432);
and U15413 (N_15413,N_14771,N_14394);
and U15414 (N_15414,N_14128,N_14562);
or U15415 (N_15415,N_14901,N_14345);
nor U15416 (N_15416,N_14775,N_14935);
xnor U15417 (N_15417,N_14970,N_14592);
nor U15418 (N_15418,N_14880,N_14497);
nand U15419 (N_15419,N_14034,N_14817);
nand U15420 (N_15420,N_14778,N_14583);
or U15421 (N_15421,N_14607,N_14067);
and U15422 (N_15422,N_14003,N_14738);
and U15423 (N_15423,N_14788,N_14505);
or U15424 (N_15424,N_14181,N_14985);
or U15425 (N_15425,N_14099,N_14726);
nand U15426 (N_15426,N_14131,N_14390);
nand U15427 (N_15427,N_14743,N_14005);
and U15428 (N_15428,N_14858,N_14144);
and U15429 (N_15429,N_14818,N_14640);
xor U15430 (N_15430,N_14079,N_14783);
or U15431 (N_15431,N_14753,N_14975);
nor U15432 (N_15432,N_14238,N_14988);
nor U15433 (N_15433,N_14650,N_14833);
nor U15434 (N_15434,N_14669,N_14093);
xor U15435 (N_15435,N_14563,N_14955);
nor U15436 (N_15436,N_14292,N_14038);
or U15437 (N_15437,N_14837,N_14887);
nor U15438 (N_15438,N_14688,N_14541);
xnor U15439 (N_15439,N_14149,N_14793);
or U15440 (N_15440,N_14254,N_14915);
nor U15441 (N_15441,N_14736,N_14618);
xor U15442 (N_15442,N_14700,N_14457);
nand U15443 (N_15443,N_14239,N_14870);
nand U15444 (N_15444,N_14925,N_14637);
nand U15445 (N_15445,N_14631,N_14512);
or U15446 (N_15446,N_14797,N_14343);
nor U15447 (N_15447,N_14405,N_14895);
nor U15448 (N_15448,N_14124,N_14796);
and U15449 (N_15449,N_14403,N_14979);
and U15450 (N_15450,N_14308,N_14670);
or U15451 (N_15451,N_14639,N_14220);
nor U15452 (N_15452,N_14416,N_14445);
and U15453 (N_15453,N_14613,N_14581);
nor U15454 (N_15454,N_14576,N_14358);
nor U15455 (N_15455,N_14332,N_14033);
and U15456 (N_15456,N_14027,N_14800);
or U15457 (N_15457,N_14190,N_14177);
and U15458 (N_15458,N_14096,N_14111);
nand U15459 (N_15459,N_14825,N_14853);
nand U15460 (N_15460,N_14830,N_14968);
or U15461 (N_15461,N_14122,N_14610);
nand U15462 (N_15462,N_14142,N_14495);
nor U15463 (N_15463,N_14899,N_14574);
nand U15464 (N_15464,N_14772,N_14934);
and U15465 (N_15465,N_14068,N_14982);
or U15466 (N_15466,N_14263,N_14455);
and U15467 (N_15467,N_14808,N_14900);
nor U15468 (N_15468,N_14323,N_14813);
or U15469 (N_15469,N_14196,N_14787);
xnor U15470 (N_15470,N_14884,N_14329);
nand U15471 (N_15471,N_14792,N_14176);
xnor U15472 (N_15472,N_14287,N_14624);
or U15473 (N_15473,N_14276,N_14485);
nand U15474 (N_15474,N_14861,N_14750);
nand U15475 (N_15475,N_14231,N_14579);
nand U15476 (N_15476,N_14635,N_14509);
xor U15477 (N_15477,N_14213,N_14691);
nand U15478 (N_15478,N_14528,N_14063);
nand U15479 (N_15479,N_14709,N_14369);
xor U15480 (N_15480,N_14760,N_14312);
nand U15481 (N_15481,N_14069,N_14569);
xnor U15482 (N_15482,N_14679,N_14521);
and U15483 (N_15483,N_14225,N_14958);
xnor U15484 (N_15484,N_14757,N_14327);
xor U15485 (N_15485,N_14437,N_14266);
nand U15486 (N_15486,N_14819,N_14945);
nor U15487 (N_15487,N_14766,N_14296);
nor U15488 (N_15488,N_14598,N_14701);
xnor U15489 (N_15489,N_14746,N_14051);
and U15490 (N_15490,N_14978,N_14538);
nand U15491 (N_15491,N_14996,N_14626);
nor U15492 (N_15492,N_14426,N_14768);
xor U15493 (N_15493,N_14897,N_14218);
or U15494 (N_15494,N_14570,N_14325);
xnor U15495 (N_15495,N_14385,N_14348);
xnor U15496 (N_15496,N_14893,N_14913);
nor U15497 (N_15497,N_14556,N_14442);
xor U15498 (N_15498,N_14134,N_14990);
or U15499 (N_15499,N_14504,N_14328);
xnor U15500 (N_15500,N_14021,N_14830);
and U15501 (N_15501,N_14566,N_14739);
xnor U15502 (N_15502,N_14422,N_14158);
nand U15503 (N_15503,N_14293,N_14334);
and U15504 (N_15504,N_14800,N_14007);
and U15505 (N_15505,N_14687,N_14984);
or U15506 (N_15506,N_14965,N_14488);
nand U15507 (N_15507,N_14652,N_14218);
or U15508 (N_15508,N_14896,N_14425);
and U15509 (N_15509,N_14901,N_14663);
nor U15510 (N_15510,N_14694,N_14016);
nor U15511 (N_15511,N_14676,N_14924);
nor U15512 (N_15512,N_14555,N_14465);
or U15513 (N_15513,N_14068,N_14104);
nor U15514 (N_15514,N_14698,N_14722);
or U15515 (N_15515,N_14896,N_14799);
nor U15516 (N_15516,N_14506,N_14621);
and U15517 (N_15517,N_14401,N_14551);
xor U15518 (N_15518,N_14973,N_14040);
nand U15519 (N_15519,N_14435,N_14959);
nand U15520 (N_15520,N_14594,N_14689);
and U15521 (N_15521,N_14344,N_14838);
xnor U15522 (N_15522,N_14806,N_14950);
nand U15523 (N_15523,N_14271,N_14959);
or U15524 (N_15524,N_14129,N_14934);
nor U15525 (N_15525,N_14074,N_14683);
nor U15526 (N_15526,N_14250,N_14816);
nand U15527 (N_15527,N_14156,N_14765);
and U15528 (N_15528,N_14573,N_14028);
nor U15529 (N_15529,N_14672,N_14337);
nor U15530 (N_15530,N_14755,N_14487);
nand U15531 (N_15531,N_14055,N_14098);
and U15532 (N_15532,N_14532,N_14382);
nand U15533 (N_15533,N_14880,N_14117);
nand U15534 (N_15534,N_14218,N_14059);
nor U15535 (N_15535,N_14102,N_14933);
nand U15536 (N_15536,N_14572,N_14055);
xor U15537 (N_15537,N_14802,N_14168);
xor U15538 (N_15538,N_14430,N_14210);
and U15539 (N_15539,N_14223,N_14757);
or U15540 (N_15540,N_14399,N_14501);
and U15541 (N_15541,N_14962,N_14929);
xor U15542 (N_15542,N_14457,N_14456);
and U15543 (N_15543,N_14949,N_14770);
nor U15544 (N_15544,N_14863,N_14310);
nand U15545 (N_15545,N_14591,N_14899);
or U15546 (N_15546,N_14953,N_14788);
or U15547 (N_15547,N_14661,N_14933);
nand U15548 (N_15548,N_14504,N_14327);
nand U15549 (N_15549,N_14979,N_14308);
or U15550 (N_15550,N_14014,N_14751);
or U15551 (N_15551,N_14961,N_14395);
nand U15552 (N_15552,N_14110,N_14194);
or U15553 (N_15553,N_14571,N_14941);
nand U15554 (N_15554,N_14947,N_14627);
or U15555 (N_15555,N_14134,N_14533);
and U15556 (N_15556,N_14080,N_14975);
nand U15557 (N_15557,N_14809,N_14011);
nand U15558 (N_15558,N_14080,N_14083);
nor U15559 (N_15559,N_14945,N_14884);
nand U15560 (N_15560,N_14972,N_14223);
and U15561 (N_15561,N_14808,N_14985);
nor U15562 (N_15562,N_14182,N_14536);
nor U15563 (N_15563,N_14792,N_14054);
nand U15564 (N_15564,N_14294,N_14257);
xor U15565 (N_15565,N_14512,N_14287);
and U15566 (N_15566,N_14280,N_14915);
xor U15567 (N_15567,N_14870,N_14441);
and U15568 (N_15568,N_14267,N_14603);
nor U15569 (N_15569,N_14504,N_14523);
nand U15570 (N_15570,N_14401,N_14377);
nand U15571 (N_15571,N_14361,N_14675);
nor U15572 (N_15572,N_14063,N_14737);
xor U15573 (N_15573,N_14945,N_14152);
or U15574 (N_15574,N_14045,N_14292);
nand U15575 (N_15575,N_14540,N_14480);
nand U15576 (N_15576,N_14396,N_14253);
or U15577 (N_15577,N_14841,N_14968);
and U15578 (N_15578,N_14801,N_14497);
and U15579 (N_15579,N_14929,N_14928);
nand U15580 (N_15580,N_14413,N_14679);
xor U15581 (N_15581,N_14428,N_14603);
xnor U15582 (N_15582,N_14980,N_14215);
nor U15583 (N_15583,N_14278,N_14131);
or U15584 (N_15584,N_14222,N_14315);
xor U15585 (N_15585,N_14587,N_14235);
xnor U15586 (N_15586,N_14451,N_14134);
xor U15587 (N_15587,N_14045,N_14250);
nand U15588 (N_15588,N_14210,N_14392);
xor U15589 (N_15589,N_14636,N_14429);
nand U15590 (N_15590,N_14501,N_14751);
nor U15591 (N_15591,N_14723,N_14755);
nor U15592 (N_15592,N_14363,N_14118);
xor U15593 (N_15593,N_14864,N_14669);
nor U15594 (N_15594,N_14378,N_14441);
and U15595 (N_15595,N_14735,N_14618);
and U15596 (N_15596,N_14583,N_14883);
nand U15597 (N_15597,N_14339,N_14340);
and U15598 (N_15598,N_14265,N_14734);
xnor U15599 (N_15599,N_14733,N_14147);
nand U15600 (N_15600,N_14330,N_14623);
nor U15601 (N_15601,N_14234,N_14357);
and U15602 (N_15602,N_14405,N_14193);
xor U15603 (N_15603,N_14636,N_14488);
nand U15604 (N_15604,N_14972,N_14718);
and U15605 (N_15605,N_14625,N_14549);
nand U15606 (N_15606,N_14388,N_14967);
or U15607 (N_15607,N_14198,N_14494);
and U15608 (N_15608,N_14013,N_14218);
nor U15609 (N_15609,N_14377,N_14616);
nand U15610 (N_15610,N_14645,N_14872);
nor U15611 (N_15611,N_14034,N_14266);
or U15612 (N_15612,N_14495,N_14954);
nor U15613 (N_15613,N_14961,N_14929);
or U15614 (N_15614,N_14916,N_14362);
nand U15615 (N_15615,N_14777,N_14246);
and U15616 (N_15616,N_14415,N_14383);
nand U15617 (N_15617,N_14729,N_14461);
nand U15618 (N_15618,N_14763,N_14661);
and U15619 (N_15619,N_14720,N_14985);
nor U15620 (N_15620,N_14377,N_14276);
and U15621 (N_15621,N_14509,N_14446);
or U15622 (N_15622,N_14414,N_14270);
xnor U15623 (N_15623,N_14048,N_14343);
and U15624 (N_15624,N_14566,N_14190);
or U15625 (N_15625,N_14700,N_14175);
nand U15626 (N_15626,N_14051,N_14550);
xor U15627 (N_15627,N_14417,N_14680);
xor U15628 (N_15628,N_14247,N_14868);
nor U15629 (N_15629,N_14622,N_14436);
nand U15630 (N_15630,N_14598,N_14921);
or U15631 (N_15631,N_14630,N_14431);
xnor U15632 (N_15632,N_14100,N_14555);
nor U15633 (N_15633,N_14273,N_14123);
and U15634 (N_15634,N_14147,N_14443);
or U15635 (N_15635,N_14426,N_14732);
xnor U15636 (N_15636,N_14468,N_14232);
xor U15637 (N_15637,N_14701,N_14590);
nor U15638 (N_15638,N_14836,N_14094);
and U15639 (N_15639,N_14715,N_14590);
and U15640 (N_15640,N_14026,N_14571);
and U15641 (N_15641,N_14916,N_14793);
or U15642 (N_15642,N_14457,N_14191);
nand U15643 (N_15643,N_14268,N_14810);
xnor U15644 (N_15644,N_14365,N_14620);
nor U15645 (N_15645,N_14730,N_14900);
or U15646 (N_15646,N_14692,N_14781);
xor U15647 (N_15647,N_14065,N_14589);
nand U15648 (N_15648,N_14840,N_14211);
xor U15649 (N_15649,N_14034,N_14714);
and U15650 (N_15650,N_14001,N_14599);
nor U15651 (N_15651,N_14413,N_14917);
xnor U15652 (N_15652,N_14694,N_14057);
and U15653 (N_15653,N_14555,N_14501);
nand U15654 (N_15654,N_14792,N_14633);
or U15655 (N_15655,N_14175,N_14424);
xnor U15656 (N_15656,N_14950,N_14196);
nand U15657 (N_15657,N_14287,N_14797);
and U15658 (N_15658,N_14223,N_14322);
nand U15659 (N_15659,N_14026,N_14761);
and U15660 (N_15660,N_14510,N_14253);
nand U15661 (N_15661,N_14771,N_14897);
xnor U15662 (N_15662,N_14586,N_14320);
xnor U15663 (N_15663,N_14684,N_14175);
or U15664 (N_15664,N_14874,N_14217);
xor U15665 (N_15665,N_14807,N_14329);
nand U15666 (N_15666,N_14085,N_14202);
nor U15667 (N_15667,N_14737,N_14184);
nor U15668 (N_15668,N_14004,N_14487);
nand U15669 (N_15669,N_14493,N_14186);
or U15670 (N_15670,N_14564,N_14974);
nor U15671 (N_15671,N_14621,N_14239);
xor U15672 (N_15672,N_14872,N_14938);
nand U15673 (N_15673,N_14038,N_14677);
xor U15674 (N_15674,N_14571,N_14432);
xor U15675 (N_15675,N_14522,N_14523);
nor U15676 (N_15676,N_14097,N_14984);
xnor U15677 (N_15677,N_14950,N_14696);
and U15678 (N_15678,N_14926,N_14184);
and U15679 (N_15679,N_14353,N_14228);
or U15680 (N_15680,N_14368,N_14906);
nand U15681 (N_15681,N_14023,N_14192);
nand U15682 (N_15682,N_14291,N_14215);
nor U15683 (N_15683,N_14426,N_14333);
or U15684 (N_15684,N_14366,N_14337);
and U15685 (N_15685,N_14665,N_14537);
nand U15686 (N_15686,N_14391,N_14972);
or U15687 (N_15687,N_14388,N_14548);
xor U15688 (N_15688,N_14865,N_14896);
nand U15689 (N_15689,N_14553,N_14937);
nor U15690 (N_15690,N_14478,N_14445);
xnor U15691 (N_15691,N_14981,N_14053);
or U15692 (N_15692,N_14558,N_14437);
nand U15693 (N_15693,N_14337,N_14748);
and U15694 (N_15694,N_14023,N_14442);
and U15695 (N_15695,N_14173,N_14940);
xor U15696 (N_15696,N_14796,N_14083);
nor U15697 (N_15697,N_14714,N_14430);
nor U15698 (N_15698,N_14424,N_14802);
xnor U15699 (N_15699,N_14625,N_14779);
or U15700 (N_15700,N_14415,N_14774);
and U15701 (N_15701,N_14495,N_14207);
or U15702 (N_15702,N_14082,N_14387);
xor U15703 (N_15703,N_14711,N_14041);
nor U15704 (N_15704,N_14763,N_14368);
xnor U15705 (N_15705,N_14640,N_14110);
or U15706 (N_15706,N_14205,N_14403);
xor U15707 (N_15707,N_14218,N_14809);
xnor U15708 (N_15708,N_14979,N_14932);
or U15709 (N_15709,N_14895,N_14930);
nor U15710 (N_15710,N_14645,N_14932);
nand U15711 (N_15711,N_14964,N_14009);
or U15712 (N_15712,N_14586,N_14994);
nand U15713 (N_15713,N_14318,N_14908);
nor U15714 (N_15714,N_14911,N_14406);
nand U15715 (N_15715,N_14318,N_14804);
nand U15716 (N_15716,N_14856,N_14213);
or U15717 (N_15717,N_14401,N_14709);
and U15718 (N_15718,N_14309,N_14201);
nand U15719 (N_15719,N_14639,N_14486);
nor U15720 (N_15720,N_14161,N_14046);
or U15721 (N_15721,N_14615,N_14807);
nand U15722 (N_15722,N_14243,N_14322);
nor U15723 (N_15723,N_14440,N_14041);
or U15724 (N_15724,N_14954,N_14382);
nand U15725 (N_15725,N_14821,N_14746);
xnor U15726 (N_15726,N_14162,N_14753);
nand U15727 (N_15727,N_14998,N_14604);
or U15728 (N_15728,N_14537,N_14119);
xnor U15729 (N_15729,N_14243,N_14464);
xnor U15730 (N_15730,N_14499,N_14182);
nand U15731 (N_15731,N_14831,N_14634);
or U15732 (N_15732,N_14524,N_14471);
and U15733 (N_15733,N_14285,N_14015);
xor U15734 (N_15734,N_14765,N_14831);
xor U15735 (N_15735,N_14441,N_14198);
nand U15736 (N_15736,N_14681,N_14881);
nor U15737 (N_15737,N_14344,N_14961);
and U15738 (N_15738,N_14443,N_14658);
nand U15739 (N_15739,N_14295,N_14526);
nor U15740 (N_15740,N_14225,N_14273);
and U15741 (N_15741,N_14414,N_14294);
or U15742 (N_15742,N_14855,N_14974);
and U15743 (N_15743,N_14123,N_14375);
nand U15744 (N_15744,N_14937,N_14873);
nand U15745 (N_15745,N_14478,N_14394);
or U15746 (N_15746,N_14947,N_14282);
nand U15747 (N_15747,N_14882,N_14673);
or U15748 (N_15748,N_14751,N_14404);
nor U15749 (N_15749,N_14239,N_14625);
and U15750 (N_15750,N_14632,N_14422);
nor U15751 (N_15751,N_14489,N_14084);
xor U15752 (N_15752,N_14220,N_14489);
nand U15753 (N_15753,N_14433,N_14482);
or U15754 (N_15754,N_14232,N_14947);
nor U15755 (N_15755,N_14521,N_14208);
and U15756 (N_15756,N_14426,N_14212);
and U15757 (N_15757,N_14804,N_14606);
nand U15758 (N_15758,N_14090,N_14007);
xnor U15759 (N_15759,N_14751,N_14151);
xor U15760 (N_15760,N_14240,N_14991);
and U15761 (N_15761,N_14182,N_14503);
nand U15762 (N_15762,N_14511,N_14198);
nor U15763 (N_15763,N_14008,N_14395);
nor U15764 (N_15764,N_14558,N_14890);
or U15765 (N_15765,N_14265,N_14425);
and U15766 (N_15766,N_14656,N_14985);
or U15767 (N_15767,N_14438,N_14334);
nor U15768 (N_15768,N_14845,N_14562);
and U15769 (N_15769,N_14546,N_14931);
xnor U15770 (N_15770,N_14965,N_14922);
or U15771 (N_15771,N_14801,N_14897);
or U15772 (N_15772,N_14732,N_14163);
and U15773 (N_15773,N_14606,N_14610);
nor U15774 (N_15774,N_14043,N_14584);
or U15775 (N_15775,N_14468,N_14042);
nor U15776 (N_15776,N_14928,N_14889);
nor U15777 (N_15777,N_14396,N_14607);
nor U15778 (N_15778,N_14285,N_14753);
and U15779 (N_15779,N_14795,N_14463);
or U15780 (N_15780,N_14243,N_14579);
nand U15781 (N_15781,N_14889,N_14552);
or U15782 (N_15782,N_14846,N_14542);
and U15783 (N_15783,N_14859,N_14274);
or U15784 (N_15784,N_14014,N_14821);
nand U15785 (N_15785,N_14706,N_14322);
xor U15786 (N_15786,N_14021,N_14167);
or U15787 (N_15787,N_14385,N_14306);
and U15788 (N_15788,N_14931,N_14155);
or U15789 (N_15789,N_14305,N_14556);
xnor U15790 (N_15790,N_14689,N_14450);
nor U15791 (N_15791,N_14900,N_14593);
nand U15792 (N_15792,N_14691,N_14036);
xnor U15793 (N_15793,N_14117,N_14873);
xnor U15794 (N_15794,N_14864,N_14402);
nand U15795 (N_15795,N_14926,N_14955);
and U15796 (N_15796,N_14530,N_14900);
and U15797 (N_15797,N_14382,N_14626);
or U15798 (N_15798,N_14569,N_14573);
and U15799 (N_15799,N_14440,N_14222);
or U15800 (N_15800,N_14590,N_14609);
xnor U15801 (N_15801,N_14577,N_14406);
nand U15802 (N_15802,N_14847,N_14349);
nand U15803 (N_15803,N_14217,N_14220);
xor U15804 (N_15804,N_14971,N_14990);
xor U15805 (N_15805,N_14486,N_14632);
and U15806 (N_15806,N_14838,N_14562);
nor U15807 (N_15807,N_14492,N_14559);
nor U15808 (N_15808,N_14847,N_14875);
nand U15809 (N_15809,N_14104,N_14288);
and U15810 (N_15810,N_14523,N_14815);
nor U15811 (N_15811,N_14590,N_14971);
xnor U15812 (N_15812,N_14332,N_14026);
xor U15813 (N_15813,N_14901,N_14653);
nor U15814 (N_15814,N_14681,N_14866);
and U15815 (N_15815,N_14812,N_14951);
nor U15816 (N_15816,N_14511,N_14651);
xnor U15817 (N_15817,N_14025,N_14133);
nand U15818 (N_15818,N_14659,N_14133);
and U15819 (N_15819,N_14979,N_14975);
and U15820 (N_15820,N_14558,N_14926);
nor U15821 (N_15821,N_14982,N_14381);
nand U15822 (N_15822,N_14964,N_14651);
and U15823 (N_15823,N_14948,N_14638);
nor U15824 (N_15824,N_14149,N_14548);
nor U15825 (N_15825,N_14365,N_14709);
nand U15826 (N_15826,N_14688,N_14449);
nand U15827 (N_15827,N_14227,N_14533);
nor U15828 (N_15828,N_14012,N_14282);
xor U15829 (N_15829,N_14364,N_14081);
and U15830 (N_15830,N_14295,N_14998);
xor U15831 (N_15831,N_14053,N_14022);
or U15832 (N_15832,N_14364,N_14021);
and U15833 (N_15833,N_14353,N_14041);
or U15834 (N_15834,N_14578,N_14997);
and U15835 (N_15835,N_14887,N_14595);
nor U15836 (N_15836,N_14348,N_14763);
nand U15837 (N_15837,N_14243,N_14849);
xor U15838 (N_15838,N_14922,N_14227);
and U15839 (N_15839,N_14769,N_14789);
xnor U15840 (N_15840,N_14176,N_14317);
xor U15841 (N_15841,N_14908,N_14169);
nor U15842 (N_15842,N_14238,N_14169);
and U15843 (N_15843,N_14648,N_14834);
and U15844 (N_15844,N_14486,N_14504);
and U15845 (N_15845,N_14789,N_14576);
xor U15846 (N_15846,N_14759,N_14114);
xnor U15847 (N_15847,N_14482,N_14747);
xnor U15848 (N_15848,N_14862,N_14907);
and U15849 (N_15849,N_14225,N_14715);
nor U15850 (N_15850,N_14655,N_14440);
xor U15851 (N_15851,N_14252,N_14467);
xnor U15852 (N_15852,N_14761,N_14234);
or U15853 (N_15853,N_14741,N_14658);
or U15854 (N_15854,N_14759,N_14357);
nor U15855 (N_15855,N_14136,N_14016);
xor U15856 (N_15856,N_14205,N_14627);
xnor U15857 (N_15857,N_14034,N_14193);
nand U15858 (N_15858,N_14644,N_14786);
xor U15859 (N_15859,N_14393,N_14929);
nand U15860 (N_15860,N_14080,N_14458);
and U15861 (N_15861,N_14182,N_14289);
nor U15862 (N_15862,N_14117,N_14134);
xnor U15863 (N_15863,N_14708,N_14421);
and U15864 (N_15864,N_14164,N_14883);
nand U15865 (N_15865,N_14947,N_14354);
xnor U15866 (N_15866,N_14450,N_14247);
nor U15867 (N_15867,N_14360,N_14500);
and U15868 (N_15868,N_14985,N_14883);
xnor U15869 (N_15869,N_14096,N_14870);
and U15870 (N_15870,N_14277,N_14504);
nand U15871 (N_15871,N_14971,N_14118);
nand U15872 (N_15872,N_14182,N_14029);
or U15873 (N_15873,N_14439,N_14762);
and U15874 (N_15874,N_14605,N_14536);
or U15875 (N_15875,N_14901,N_14627);
nand U15876 (N_15876,N_14126,N_14510);
or U15877 (N_15877,N_14032,N_14854);
or U15878 (N_15878,N_14320,N_14845);
xor U15879 (N_15879,N_14402,N_14626);
nor U15880 (N_15880,N_14910,N_14253);
nor U15881 (N_15881,N_14814,N_14634);
nand U15882 (N_15882,N_14672,N_14106);
nor U15883 (N_15883,N_14360,N_14567);
nand U15884 (N_15884,N_14926,N_14366);
nand U15885 (N_15885,N_14318,N_14462);
nand U15886 (N_15886,N_14612,N_14435);
and U15887 (N_15887,N_14513,N_14215);
and U15888 (N_15888,N_14278,N_14407);
nand U15889 (N_15889,N_14297,N_14068);
nand U15890 (N_15890,N_14005,N_14976);
nand U15891 (N_15891,N_14068,N_14261);
nor U15892 (N_15892,N_14404,N_14578);
xor U15893 (N_15893,N_14439,N_14224);
and U15894 (N_15894,N_14328,N_14565);
nand U15895 (N_15895,N_14550,N_14514);
xor U15896 (N_15896,N_14329,N_14875);
nor U15897 (N_15897,N_14693,N_14309);
or U15898 (N_15898,N_14007,N_14180);
or U15899 (N_15899,N_14136,N_14328);
or U15900 (N_15900,N_14368,N_14456);
xor U15901 (N_15901,N_14369,N_14503);
or U15902 (N_15902,N_14358,N_14815);
xnor U15903 (N_15903,N_14704,N_14228);
or U15904 (N_15904,N_14569,N_14192);
nor U15905 (N_15905,N_14717,N_14434);
xor U15906 (N_15906,N_14749,N_14108);
xnor U15907 (N_15907,N_14142,N_14015);
nand U15908 (N_15908,N_14304,N_14983);
or U15909 (N_15909,N_14100,N_14195);
xor U15910 (N_15910,N_14597,N_14395);
nand U15911 (N_15911,N_14382,N_14018);
xor U15912 (N_15912,N_14966,N_14013);
nand U15913 (N_15913,N_14551,N_14911);
nand U15914 (N_15914,N_14740,N_14079);
and U15915 (N_15915,N_14718,N_14083);
nor U15916 (N_15916,N_14994,N_14550);
nand U15917 (N_15917,N_14261,N_14501);
xnor U15918 (N_15918,N_14869,N_14139);
and U15919 (N_15919,N_14470,N_14466);
nor U15920 (N_15920,N_14302,N_14564);
or U15921 (N_15921,N_14400,N_14941);
and U15922 (N_15922,N_14039,N_14959);
nor U15923 (N_15923,N_14344,N_14402);
nor U15924 (N_15924,N_14207,N_14930);
or U15925 (N_15925,N_14173,N_14553);
nor U15926 (N_15926,N_14992,N_14138);
or U15927 (N_15927,N_14851,N_14838);
xor U15928 (N_15928,N_14107,N_14891);
xor U15929 (N_15929,N_14215,N_14321);
xnor U15930 (N_15930,N_14051,N_14145);
xnor U15931 (N_15931,N_14380,N_14054);
and U15932 (N_15932,N_14660,N_14983);
and U15933 (N_15933,N_14597,N_14356);
and U15934 (N_15934,N_14735,N_14761);
xor U15935 (N_15935,N_14430,N_14036);
nor U15936 (N_15936,N_14065,N_14983);
xor U15937 (N_15937,N_14929,N_14895);
or U15938 (N_15938,N_14900,N_14242);
or U15939 (N_15939,N_14528,N_14435);
nand U15940 (N_15940,N_14601,N_14121);
or U15941 (N_15941,N_14610,N_14913);
nor U15942 (N_15942,N_14779,N_14739);
or U15943 (N_15943,N_14180,N_14252);
or U15944 (N_15944,N_14718,N_14239);
and U15945 (N_15945,N_14393,N_14020);
nand U15946 (N_15946,N_14056,N_14905);
xor U15947 (N_15947,N_14116,N_14460);
and U15948 (N_15948,N_14764,N_14367);
and U15949 (N_15949,N_14504,N_14391);
nand U15950 (N_15950,N_14273,N_14949);
xnor U15951 (N_15951,N_14371,N_14173);
nand U15952 (N_15952,N_14724,N_14055);
or U15953 (N_15953,N_14534,N_14079);
nand U15954 (N_15954,N_14316,N_14954);
and U15955 (N_15955,N_14451,N_14231);
and U15956 (N_15956,N_14254,N_14008);
and U15957 (N_15957,N_14544,N_14105);
xnor U15958 (N_15958,N_14390,N_14407);
xnor U15959 (N_15959,N_14130,N_14043);
and U15960 (N_15960,N_14465,N_14984);
or U15961 (N_15961,N_14190,N_14162);
nor U15962 (N_15962,N_14280,N_14716);
and U15963 (N_15963,N_14621,N_14898);
xor U15964 (N_15964,N_14638,N_14865);
and U15965 (N_15965,N_14362,N_14337);
and U15966 (N_15966,N_14466,N_14967);
nor U15967 (N_15967,N_14073,N_14692);
xnor U15968 (N_15968,N_14604,N_14104);
nand U15969 (N_15969,N_14942,N_14750);
or U15970 (N_15970,N_14251,N_14714);
nand U15971 (N_15971,N_14053,N_14760);
and U15972 (N_15972,N_14271,N_14896);
or U15973 (N_15973,N_14132,N_14250);
or U15974 (N_15974,N_14991,N_14117);
nand U15975 (N_15975,N_14563,N_14445);
nand U15976 (N_15976,N_14179,N_14976);
or U15977 (N_15977,N_14412,N_14081);
nor U15978 (N_15978,N_14633,N_14490);
xor U15979 (N_15979,N_14928,N_14789);
nor U15980 (N_15980,N_14868,N_14196);
nor U15981 (N_15981,N_14500,N_14123);
nor U15982 (N_15982,N_14158,N_14451);
nand U15983 (N_15983,N_14939,N_14066);
xnor U15984 (N_15984,N_14163,N_14321);
nor U15985 (N_15985,N_14878,N_14258);
or U15986 (N_15986,N_14106,N_14285);
nand U15987 (N_15987,N_14776,N_14394);
nand U15988 (N_15988,N_14546,N_14667);
or U15989 (N_15989,N_14674,N_14395);
and U15990 (N_15990,N_14149,N_14293);
or U15991 (N_15991,N_14956,N_14253);
or U15992 (N_15992,N_14670,N_14703);
nand U15993 (N_15993,N_14780,N_14362);
nand U15994 (N_15994,N_14514,N_14039);
nand U15995 (N_15995,N_14728,N_14212);
xnor U15996 (N_15996,N_14388,N_14809);
or U15997 (N_15997,N_14436,N_14444);
nor U15998 (N_15998,N_14424,N_14126);
xnor U15999 (N_15999,N_14631,N_14203);
nand U16000 (N_16000,N_15101,N_15738);
xnor U16001 (N_16001,N_15424,N_15077);
nand U16002 (N_16002,N_15399,N_15090);
nor U16003 (N_16003,N_15108,N_15201);
xnor U16004 (N_16004,N_15755,N_15074);
nand U16005 (N_16005,N_15457,N_15986);
or U16006 (N_16006,N_15121,N_15223);
xor U16007 (N_16007,N_15066,N_15430);
nor U16008 (N_16008,N_15858,N_15254);
nor U16009 (N_16009,N_15282,N_15174);
and U16010 (N_16010,N_15132,N_15651);
and U16011 (N_16011,N_15652,N_15219);
or U16012 (N_16012,N_15106,N_15646);
xor U16013 (N_16013,N_15823,N_15727);
xnor U16014 (N_16014,N_15281,N_15486);
nor U16015 (N_16015,N_15972,N_15530);
xor U16016 (N_16016,N_15177,N_15175);
xor U16017 (N_16017,N_15683,N_15600);
and U16018 (N_16018,N_15521,N_15190);
nor U16019 (N_16019,N_15470,N_15673);
and U16020 (N_16020,N_15148,N_15788);
and U16021 (N_16021,N_15447,N_15191);
nand U16022 (N_16022,N_15978,N_15378);
nand U16023 (N_16023,N_15348,N_15333);
or U16024 (N_16024,N_15273,N_15178);
and U16025 (N_16025,N_15630,N_15908);
nand U16026 (N_16026,N_15815,N_15428);
or U16027 (N_16027,N_15199,N_15360);
nor U16028 (N_16028,N_15163,N_15770);
and U16029 (N_16029,N_15809,N_15312);
or U16030 (N_16030,N_15393,N_15391);
and U16031 (N_16031,N_15371,N_15446);
xor U16032 (N_16032,N_15344,N_15276);
nor U16033 (N_16033,N_15542,N_15316);
xor U16034 (N_16034,N_15395,N_15822);
xor U16035 (N_16035,N_15413,N_15568);
nand U16036 (N_16036,N_15492,N_15362);
nand U16037 (N_16037,N_15329,N_15930);
or U16038 (N_16038,N_15143,N_15971);
or U16039 (N_16039,N_15136,N_15948);
nor U16040 (N_16040,N_15152,N_15602);
xnor U16041 (N_16041,N_15490,N_15476);
nor U16042 (N_16042,N_15789,N_15123);
xor U16043 (N_16043,N_15583,N_15050);
or U16044 (N_16044,N_15648,N_15624);
xnor U16045 (N_16045,N_15157,N_15252);
nand U16046 (N_16046,N_15386,N_15150);
nand U16047 (N_16047,N_15968,N_15024);
xnor U16048 (N_16048,N_15692,N_15512);
nor U16049 (N_16049,N_15133,N_15883);
or U16050 (N_16050,N_15632,N_15766);
and U16051 (N_16051,N_15647,N_15695);
nor U16052 (N_16052,N_15072,N_15185);
or U16053 (N_16053,N_15843,N_15380);
nand U16054 (N_16054,N_15603,N_15880);
or U16055 (N_16055,N_15627,N_15240);
nor U16056 (N_16056,N_15062,N_15158);
or U16057 (N_16057,N_15573,N_15100);
or U16058 (N_16058,N_15529,N_15722);
xnor U16059 (N_16059,N_15308,N_15743);
and U16060 (N_16060,N_15554,N_15332);
or U16061 (N_16061,N_15239,N_15419);
and U16062 (N_16062,N_15297,N_15144);
xnor U16063 (N_16063,N_15608,N_15562);
nand U16064 (N_16064,N_15207,N_15225);
nor U16065 (N_16065,N_15059,N_15742);
nand U16066 (N_16066,N_15941,N_15083);
xor U16067 (N_16067,N_15925,N_15350);
nand U16068 (N_16068,N_15286,N_15913);
nor U16069 (N_16069,N_15844,N_15811);
nand U16070 (N_16070,N_15641,N_15991);
xor U16071 (N_16071,N_15871,N_15764);
or U16072 (N_16072,N_15345,N_15688);
nor U16073 (N_16073,N_15214,N_15576);
xor U16074 (N_16074,N_15650,N_15656);
or U16075 (N_16075,N_15759,N_15537);
nor U16076 (N_16076,N_15967,N_15266);
and U16077 (N_16077,N_15054,N_15610);
and U16078 (N_16078,N_15716,N_15454);
and U16079 (N_16079,N_15127,N_15633);
or U16080 (N_16080,N_15729,N_15825);
nand U16081 (N_16081,N_15712,N_15515);
or U16082 (N_16082,N_15795,N_15997);
nor U16083 (N_16083,N_15028,N_15230);
xnor U16084 (N_16084,N_15096,N_15078);
nand U16085 (N_16085,N_15593,N_15741);
and U16086 (N_16086,N_15998,N_15920);
xnor U16087 (N_16087,N_15414,N_15000);
nand U16088 (N_16088,N_15499,N_15249);
nor U16089 (N_16089,N_15406,N_15812);
or U16090 (N_16090,N_15315,N_15945);
nand U16091 (N_16091,N_15791,N_15325);
nor U16092 (N_16092,N_15305,N_15487);
and U16093 (N_16093,N_15820,N_15776);
nand U16094 (N_16094,N_15319,N_15995);
nand U16095 (N_16095,N_15217,N_15346);
and U16096 (N_16096,N_15241,N_15409);
nor U16097 (N_16097,N_15005,N_15942);
xnor U16098 (N_16098,N_15122,N_15555);
nand U16099 (N_16099,N_15668,N_15167);
xnor U16100 (N_16100,N_15556,N_15804);
or U16101 (N_16101,N_15619,N_15238);
or U16102 (N_16102,N_15452,N_15450);
or U16103 (N_16103,N_15489,N_15359);
xor U16104 (N_16104,N_15002,N_15003);
or U16105 (N_16105,N_15464,N_15643);
nand U16106 (N_16106,N_15361,N_15257);
nand U16107 (N_16107,N_15307,N_15436);
or U16108 (N_16108,N_15453,N_15543);
xnor U16109 (N_16109,N_15782,N_15874);
xnor U16110 (N_16110,N_15418,N_15417);
xor U16111 (N_16111,N_15203,N_15887);
xor U16112 (N_16112,N_15828,N_15025);
nor U16113 (N_16113,N_15434,N_15001);
or U16114 (N_16114,N_15717,N_15895);
and U16115 (N_16115,N_15445,N_15700);
nor U16116 (N_16116,N_15611,N_15046);
and U16117 (N_16117,N_15351,N_15889);
or U16118 (N_16118,N_15721,N_15277);
nor U16119 (N_16119,N_15037,N_15243);
nand U16120 (N_16120,N_15231,N_15961);
nand U16121 (N_16121,N_15279,N_15213);
nor U16122 (N_16122,N_15129,N_15671);
and U16123 (N_16123,N_15161,N_15228);
nor U16124 (N_16124,N_15410,N_15058);
nor U16125 (N_16125,N_15372,N_15118);
and U16126 (N_16126,N_15732,N_15735);
or U16127 (N_16127,N_15964,N_15979);
and U16128 (N_16128,N_15119,N_15658);
xor U16129 (N_16129,N_15864,N_15128);
or U16130 (N_16130,N_15038,N_15196);
nor U16131 (N_16131,N_15120,N_15839);
or U16132 (N_16132,N_15027,N_15993);
and U16133 (N_16133,N_15097,N_15443);
xnor U16134 (N_16134,N_15425,N_15909);
xor U16135 (N_16135,N_15299,N_15509);
nor U16136 (N_16136,N_15481,N_15339);
and U16137 (N_16137,N_15797,N_15900);
and U16138 (N_16138,N_15637,N_15757);
nand U16139 (N_16139,N_15621,N_15879);
nand U16140 (N_16140,N_15438,N_15403);
xnor U16141 (N_16141,N_15540,N_15309);
and U16142 (N_16142,N_15326,N_15165);
or U16143 (N_16143,N_15469,N_15639);
nor U16144 (N_16144,N_15687,N_15954);
nor U16145 (N_16145,N_15884,N_15153);
nand U16146 (N_16146,N_15194,N_15682);
nand U16147 (N_16147,N_15007,N_15892);
xnor U16148 (N_16148,N_15661,N_15578);
nor U16149 (N_16149,N_15726,N_15155);
nand U16150 (N_16150,N_15951,N_15181);
and U16151 (N_16151,N_15963,N_15367);
or U16152 (N_16152,N_15752,N_15253);
or U16153 (N_16153,N_15672,N_15754);
nor U16154 (N_16154,N_15176,N_15160);
nor U16155 (N_16155,N_15218,N_15278);
xor U16156 (N_16156,N_15775,N_15922);
or U16157 (N_16157,N_15517,N_15131);
and U16158 (N_16158,N_15209,N_15761);
or U16159 (N_16159,N_15534,N_15533);
xnor U16160 (N_16160,N_15818,N_15349);
or U16161 (N_16161,N_15455,N_15705);
or U16162 (N_16162,N_15549,N_15079);
nor U16163 (N_16163,N_15103,N_15494);
nor U16164 (N_16164,N_15869,N_15426);
xor U16165 (N_16165,N_15435,N_15935);
nand U16166 (N_16166,N_15875,N_15644);
xnor U16167 (N_16167,N_15965,N_15065);
nand U16168 (N_16168,N_15793,N_15599);
or U16169 (N_16169,N_15873,N_15669);
and U16170 (N_16170,N_15164,N_15114);
and U16171 (N_16171,N_15328,N_15220);
xor U16172 (N_16172,N_15711,N_15865);
and U16173 (N_16173,N_15753,N_15064);
xnor U16174 (N_16174,N_15575,N_15248);
nand U16175 (N_16175,N_15032,N_15989);
nand U16176 (N_16176,N_15431,N_15283);
or U16177 (N_16177,N_15660,N_15667);
nand U16178 (N_16178,N_15388,N_15786);
nor U16179 (N_16179,N_15642,N_15597);
and U16180 (N_16180,N_15045,N_15352);
and U16181 (N_16181,N_15068,N_15763);
or U16182 (N_16182,N_15698,N_15511);
nand U16183 (N_16183,N_15044,N_15336);
xnor U16184 (N_16184,N_15681,N_15347);
xnor U16185 (N_16185,N_15561,N_15794);
xor U16186 (N_16186,N_15290,N_15676);
and U16187 (N_16187,N_15557,N_15212);
nor U16188 (N_16188,N_15029,N_15265);
xor U16189 (N_16189,N_15594,N_15317);
or U16190 (N_16190,N_15284,N_15094);
nand U16191 (N_16191,N_15514,N_15723);
or U16192 (N_16192,N_15442,N_15507);
and U16193 (N_16193,N_15084,N_15462);
nand U16194 (N_16194,N_15404,N_15545);
or U16195 (N_16195,N_15595,N_15060);
or U16196 (N_16196,N_15402,N_15192);
and U16197 (N_16197,N_15306,N_15746);
or U16198 (N_16198,N_15973,N_15082);
nand U16199 (N_16199,N_15725,N_15500);
and U16200 (N_16200,N_15970,N_15737);
nand U16201 (N_16201,N_15992,N_15829);
nor U16202 (N_16202,N_15977,N_15141);
and U16203 (N_16203,N_15769,N_15852);
xnor U16204 (N_16204,N_15547,N_15894);
xor U16205 (N_16205,N_15510,N_15899);
nor U16206 (N_16206,N_15915,N_15061);
nor U16207 (N_16207,N_15876,N_15645);
nor U16208 (N_16208,N_15242,N_15466);
nand U16209 (N_16209,N_15536,N_15800);
and U16210 (N_16210,N_15354,N_15444);
nor U16211 (N_16211,N_15370,N_15188);
xnor U16212 (N_16212,N_15051,N_15006);
xor U16213 (N_16213,N_15893,N_15193);
nor U16214 (N_16214,N_15382,N_15373);
and U16215 (N_16215,N_15923,N_15826);
or U16216 (N_16216,N_15338,N_15056);
xor U16217 (N_16217,N_15861,N_15092);
xor U16218 (N_16218,N_15496,N_15206);
nand U16219 (N_16219,N_15936,N_15982);
and U16220 (N_16220,N_15246,N_15098);
nor U16221 (N_16221,N_15969,N_15263);
and U16222 (N_16222,N_15151,N_15974);
nand U16223 (N_16223,N_15842,N_15030);
xor U16224 (N_16224,N_15919,N_15606);
nand U16225 (N_16225,N_15017,N_15535);
nor U16226 (N_16226,N_15985,N_15670);
and U16227 (N_16227,N_15034,N_15484);
nor U16228 (N_16228,N_15748,N_15385);
and U16229 (N_16229,N_15762,N_15322);
nor U16230 (N_16230,N_15256,N_15983);
nand U16231 (N_16231,N_15270,N_15172);
nand U16232 (N_16232,N_15262,N_15693);
or U16233 (N_16233,N_15204,N_15719);
or U16234 (N_16234,N_15314,N_15666);
and U16235 (N_16235,N_15421,N_15888);
nand U16236 (N_16236,N_15657,N_15622);
xor U16237 (N_16237,N_15665,N_15335);
nand U16238 (N_16238,N_15837,N_15043);
xnor U16239 (N_16239,N_15427,N_15856);
xnor U16240 (N_16240,N_15095,N_15806);
nand U16241 (N_16241,N_15955,N_15853);
and U16242 (N_16242,N_15664,N_15471);
xnor U16243 (N_16243,N_15113,N_15274);
nor U16244 (N_16244,N_15012,N_15659);
xnor U16245 (N_16245,N_15949,N_15311);
or U16246 (N_16246,N_15004,N_15126);
xnor U16247 (N_16247,N_15291,N_15912);
xor U16248 (N_16248,N_15886,N_15574);
or U16249 (N_16249,N_15300,N_15878);
and U16250 (N_16250,N_15778,N_15411);
nor U16251 (N_16251,N_15750,N_15039);
nor U16252 (N_16252,N_15473,N_15703);
nor U16253 (N_16253,N_15298,N_15287);
nand U16254 (N_16254,N_15740,N_15903);
or U16255 (N_16255,N_15774,N_15321);
xor U16256 (N_16256,N_15042,N_15397);
and U16257 (N_16257,N_15546,N_15898);
xor U16258 (N_16258,N_15891,N_15468);
nor U16259 (N_16259,N_15847,N_15707);
nor U16260 (N_16260,N_15293,N_15405);
xnor U16261 (N_16261,N_15495,N_15805);
nand U16262 (N_16262,N_15882,N_15690);
and U16263 (N_16263,N_15572,N_15803);
or U16264 (N_16264,N_15186,N_15343);
xor U16265 (N_16265,N_15130,N_15474);
or U16266 (N_16266,N_15099,N_15744);
nand U16267 (N_16267,N_15526,N_15171);
nor U16268 (N_16268,N_15053,N_15689);
xor U16269 (N_16269,N_15790,N_15866);
or U16270 (N_16270,N_15236,N_15303);
or U16271 (N_16271,N_15234,N_15701);
nor U16272 (N_16272,N_15137,N_15959);
and U16273 (N_16273,N_15168,N_15943);
nor U16274 (N_16274,N_15439,N_15341);
and U16275 (N_16275,N_15760,N_15902);
or U16276 (N_16276,N_15244,N_15467);
nor U16277 (N_16277,N_15086,N_15394);
nor U16278 (N_16278,N_15662,N_15553);
xnor U16279 (N_16279,N_15010,N_15679);
nor U16280 (N_16280,N_15233,N_15585);
or U16281 (N_16281,N_15988,N_15751);
xnor U16282 (N_16282,N_15859,N_15586);
and U16283 (N_16283,N_15697,N_15292);
and U16284 (N_16284,N_15807,N_15071);
xor U16285 (N_16285,N_15960,N_15264);
nand U16286 (N_16286,N_15756,N_15590);
nor U16287 (N_16287,N_15867,N_15182);
and U16288 (N_16288,N_15928,N_15035);
or U16289 (N_16289,N_15226,N_15532);
and U16290 (N_16290,N_15901,N_15015);
nor U16291 (N_16291,N_15834,N_15838);
nor U16292 (N_16292,N_15835,N_15910);
xnor U16293 (N_16293,N_15854,N_15376);
nand U16294 (N_16294,N_15550,N_15523);
xnor U16295 (N_16295,N_15541,N_15166);
or U16296 (N_16296,N_15851,N_15475);
xor U16297 (N_16297,N_15832,N_15635);
nor U16298 (N_16298,N_15483,N_15294);
and U16299 (N_16299,N_15868,N_15390);
nor U16300 (N_16300,N_15433,N_15357);
and U16301 (N_16301,N_15567,N_15031);
nor U16302 (N_16302,N_15154,N_15944);
and U16303 (N_16303,N_15195,N_15544);
and U16304 (N_16304,N_15479,N_15021);
or U16305 (N_16305,N_15087,N_15816);
nor U16306 (N_16306,N_15009,N_15911);
or U16307 (N_16307,N_15200,N_15401);
and U16308 (N_16308,N_15677,N_15310);
and U16309 (N_16309,N_15458,N_15708);
nor U16310 (N_16310,N_15503,N_15674);
or U16311 (N_16311,N_15288,N_15558);
and U16312 (N_16312,N_15680,N_15840);
xnor U16313 (N_16313,N_15745,N_15598);
and U16314 (N_16314,N_15771,N_15147);
xor U16315 (N_16315,N_15956,N_15724);
or U16316 (N_16316,N_15491,N_15999);
xnor U16317 (N_16317,N_15379,N_15250);
nand U16318 (N_16318,N_15846,N_15613);
and U16319 (N_16319,N_15581,N_15862);
xor U16320 (N_16320,N_15105,N_15441);
and U16321 (N_16321,N_15437,N_15636);
and U16322 (N_16322,N_15366,N_15259);
and U16323 (N_16323,N_15596,N_15145);
nand U16324 (N_16324,N_15396,N_15653);
and U16325 (N_16325,N_15781,N_15987);
or U16326 (N_16326,N_15601,N_15626);
nand U16327 (N_16327,N_15422,N_15519);
and U16328 (N_16328,N_15318,N_15261);
or U16329 (N_16329,N_15728,N_15159);
or U16330 (N_16330,N_15146,N_15041);
and U16331 (N_16331,N_15472,N_15398);
and U16332 (N_16332,N_15821,N_15216);
nor U16333 (N_16333,N_15081,N_15953);
xor U16334 (N_16334,N_15202,N_15358);
and U16335 (N_16335,N_15817,N_15747);
or U16336 (N_16336,N_15400,N_15224);
nor U16337 (N_16337,N_15827,N_15940);
nor U16338 (N_16338,N_15587,N_15089);
nor U16339 (N_16339,N_15720,N_15055);
and U16340 (N_16340,N_15088,N_15138);
nor U16341 (N_16341,N_15552,N_15980);
xor U16342 (N_16342,N_15631,N_15020);
nor U16343 (N_16343,N_15407,N_15124);
and U16344 (N_16344,N_15104,N_15932);
nor U16345 (N_16345,N_15018,N_15432);
xnor U16346 (N_16346,N_15531,N_15918);
nand U16347 (N_16347,N_15654,N_15275);
xor U16348 (N_16348,N_15251,N_15420);
nand U16349 (N_16349,N_15260,N_15460);
nor U16350 (N_16350,N_15779,N_15237);
and U16351 (N_16351,N_15872,N_15787);
and U16352 (N_16352,N_15502,N_15501);
nand U16353 (N_16353,N_15247,N_15258);
nor U16354 (N_16354,N_15620,N_15845);
xor U16355 (N_16355,N_15210,N_15629);
and U16356 (N_16356,N_15208,N_15736);
and U16357 (N_16357,N_15589,N_15461);
xnor U16358 (N_16358,N_15485,N_15327);
nand U16359 (N_16359,N_15022,N_15855);
or U16360 (N_16360,N_15966,N_15924);
and U16361 (N_16361,N_15836,N_15819);
xnor U16362 (N_16362,N_15798,N_15429);
and U16363 (N_16363,N_15885,N_15189);
nor U16364 (N_16364,N_15772,N_15684);
and U16365 (N_16365,N_15075,N_15733);
or U16366 (N_16366,N_15374,N_15093);
xnor U16367 (N_16367,N_15423,N_15504);
nor U16368 (N_16368,N_15235,N_15881);
nor U16369 (N_16369,N_15296,N_15267);
or U16370 (N_16370,N_15506,N_15984);
nor U16371 (N_16371,N_15571,N_15580);
or U16372 (N_16372,N_15917,N_15057);
and U16373 (N_16373,N_15134,N_15369);
and U16374 (N_16374,N_15187,N_15841);
or U16375 (N_16375,N_15933,N_15067);
and U16376 (N_16376,N_15952,N_15814);
and U16377 (N_16377,N_15634,N_15169);
nor U16378 (N_16378,N_15033,N_15564);
and U16379 (N_16379,N_15280,N_15527);
and U16380 (N_16380,N_15715,N_15111);
nor U16381 (N_16381,N_15582,N_15649);
and U16382 (N_16382,N_15850,N_15295);
nand U16383 (N_16383,N_15459,N_15478);
xor U16384 (N_16384,N_15813,N_15440);
and U16385 (N_16385,N_15768,N_15675);
nand U16386 (N_16386,N_15073,N_15498);
or U16387 (N_16387,N_15016,N_15508);
or U16388 (N_16388,N_15205,N_15023);
or U16389 (N_16389,N_15849,N_15686);
nor U16390 (N_16390,N_15916,N_15831);
or U16391 (N_16391,N_15363,N_15896);
nand U16392 (N_16392,N_15416,N_15616);
or U16393 (N_16393,N_15019,N_15516);
xor U16394 (N_16394,N_15767,N_15914);
and U16395 (N_16395,N_15116,N_15785);
nand U16396 (N_16396,N_15342,N_15139);
nand U16397 (N_16397,N_15824,N_15758);
xor U16398 (N_16398,N_15625,N_15389);
or U16399 (N_16399,N_15232,N_15691);
and U16400 (N_16400,N_15539,N_15493);
or U16401 (N_16401,N_15008,N_15921);
or U16402 (N_16402,N_15513,N_15857);
nand U16403 (N_16403,N_15245,N_15927);
nand U16404 (N_16404,N_15730,N_15694);
xnor U16405 (N_16405,N_15799,N_15377);
nor U16406 (N_16406,N_15482,N_15356);
and U16407 (N_16407,N_15699,N_15860);
and U16408 (N_16408,N_15777,N_15184);
nand U16409 (N_16409,N_15962,N_15947);
nor U16410 (N_16410,N_15183,N_15591);
xor U16411 (N_16411,N_15375,N_15117);
nor U16412 (N_16412,N_15323,N_15085);
and U16413 (N_16413,N_15149,N_15520);
and U16414 (N_16414,N_15331,N_15285);
nand U16415 (N_16415,N_15609,N_15802);
nor U16416 (N_16416,N_15488,N_15518);
xnor U16417 (N_16417,N_15638,N_15463);
nor U16418 (N_16418,N_15938,N_15710);
xnor U16419 (N_16419,N_15497,N_15412);
xor U16420 (N_16420,N_15026,N_15939);
and U16421 (N_16421,N_15528,N_15222);
nand U16422 (N_16422,N_15135,N_15538);
nor U16423 (N_16423,N_15477,N_15091);
and U16424 (N_16424,N_15272,N_15566);
nor U16425 (N_16425,N_15731,N_15465);
or U16426 (N_16426,N_15355,N_15069);
or U16427 (N_16427,N_15353,N_15907);
nand U16428 (N_16428,N_15702,N_15289);
xnor U16429 (N_16429,N_15052,N_15047);
xor U16430 (N_16430,N_15340,N_15456);
and U16431 (N_16431,N_15584,N_15180);
xnor U16432 (N_16432,N_15269,N_15313);
xnor U16433 (N_16433,N_15107,N_15381);
and U16434 (N_16434,N_15227,N_15783);
and U16435 (N_16435,N_15996,N_15931);
or U16436 (N_16436,N_15480,N_15976);
or U16437 (N_16437,N_15063,N_15368);
nand U16438 (N_16438,N_15897,N_15615);
xor U16439 (N_16439,N_15696,N_15179);
nor U16440 (N_16440,N_15801,N_15577);
nor U16441 (N_16441,N_15014,N_15870);
xor U16442 (N_16442,N_15229,N_15565);
and U16443 (N_16443,N_15848,N_15387);
xor U16444 (N_16444,N_15579,N_15364);
and U16445 (N_16445,N_15011,N_15448);
nor U16446 (N_16446,N_15877,N_15392);
or U16447 (N_16447,N_15102,N_15173);
or U16448 (N_16448,N_15830,N_15330);
nand U16449 (N_16449,N_15994,N_15334);
nor U16450 (N_16450,N_15551,N_15505);
and U16451 (N_16451,N_15904,N_15569);
and U16452 (N_16452,N_15588,N_15934);
nand U16453 (N_16453,N_15142,N_15605);
and U16454 (N_16454,N_15780,N_15663);
nand U16455 (N_16455,N_15162,N_15324);
and U16456 (N_16456,N_15950,N_15833);
or U16457 (N_16457,N_15975,N_15906);
xnor U16458 (N_16458,N_15685,N_15607);
xnor U16459 (N_16459,N_15614,N_15125);
xor U16460 (N_16460,N_15784,N_15524);
and U16461 (N_16461,N_15990,N_15320);
and U16462 (N_16462,N_15773,N_15604);
nand U16463 (N_16463,N_15678,N_15156);
or U16464 (N_16464,N_15765,N_15628);
and U16465 (N_16465,N_15080,N_15640);
nor U16466 (N_16466,N_15709,N_15749);
nor U16467 (N_16467,N_15548,N_15617);
nor U16468 (N_16468,N_15383,N_15215);
and U16469 (N_16469,N_15076,N_15040);
xor U16470 (N_16470,N_15559,N_15714);
nand U16471 (N_16471,N_15890,N_15796);
nor U16472 (N_16472,N_15197,N_15937);
or U16473 (N_16473,N_15449,N_15563);
and U16474 (N_16474,N_15365,N_15618);
xnor U16475 (N_16475,N_15704,N_15926);
nor U16476 (N_16476,N_15109,N_15255);
and U16477 (N_16477,N_15958,N_15036);
nand U16478 (N_16478,N_15792,N_15302);
nor U16479 (N_16479,N_15221,N_15592);
xor U16480 (N_16480,N_15301,N_15946);
nand U16481 (N_16481,N_15451,N_15408);
xnor U16482 (N_16482,N_15810,N_15713);
and U16483 (N_16483,N_15905,N_15337);
xor U16484 (N_16484,N_15304,N_15110);
nor U16485 (N_16485,N_15612,N_15718);
nor U16486 (N_16486,N_15115,N_15981);
nand U16487 (N_16487,N_15049,N_15522);
or U16488 (N_16488,N_15706,N_15268);
xnor U16489 (N_16489,N_15525,N_15929);
and U16490 (N_16490,N_15739,N_15560);
or U16491 (N_16491,N_15957,N_15140);
nand U16492 (N_16492,N_15863,N_15048);
or U16493 (N_16493,N_15198,N_15415);
nor U16494 (N_16494,N_15734,N_15623);
and U16495 (N_16495,N_15808,N_15570);
nand U16496 (N_16496,N_15013,N_15070);
or U16497 (N_16497,N_15112,N_15655);
nand U16498 (N_16498,N_15170,N_15271);
nor U16499 (N_16499,N_15211,N_15384);
xnor U16500 (N_16500,N_15659,N_15899);
or U16501 (N_16501,N_15149,N_15663);
nor U16502 (N_16502,N_15448,N_15536);
xnor U16503 (N_16503,N_15050,N_15252);
or U16504 (N_16504,N_15419,N_15404);
nand U16505 (N_16505,N_15905,N_15947);
nor U16506 (N_16506,N_15831,N_15513);
and U16507 (N_16507,N_15654,N_15261);
xnor U16508 (N_16508,N_15353,N_15561);
or U16509 (N_16509,N_15542,N_15272);
nor U16510 (N_16510,N_15825,N_15617);
or U16511 (N_16511,N_15243,N_15562);
nor U16512 (N_16512,N_15057,N_15355);
or U16513 (N_16513,N_15928,N_15834);
and U16514 (N_16514,N_15592,N_15048);
nor U16515 (N_16515,N_15459,N_15513);
nor U16516 (N_16516,N_15371,N_15499);
nor U16517 (N_16517,N_15766,N_15165);
xnor U16518 (N_16518,N_15336,N_15443);
xor U16519 (N_16519,N_15796,N_15366);
nor U16520 (N_16520,N_15087,N_15567);
or U16521 (N_16521,N_15289,N_15004);
nand U16522 (N_16522,N_15559,N_15388);
nand U16523 (N_16523,N_15719,N_15828);
nand U16524 (N_16524,N_15206,N_15100);
or U16525 (N_16525,N_15061,N_15676);
nand U16526 (N_16526,N_15791,N_15939);
or U16527 (N_16527,N_15946,N_15483);
xor U16528 (N_16528,N_15210,N_15800);
or U16529 (N_16529,N_15479,N_15289);
nor U16530 (N_16530,N_15410,N_15494);
nor U16531 (N_16531,N_15559,N_15062);
or U16532 (N_16532,N_15850,N_15021);
xor U16533 (N_16533,N_15889,N_15556);
xor U16534 (N_16534,N_15039,N_15656);
or U16535 (N_16535,N_15647,N_15093);
or U16536 (N_16536,N_15049,N_15003);
nor U16537 (N_16537,N_15669,N_15293);
and U16538 (N_16538,N_15994,N_15167);
nand U16539 (N_16539,N_15582,N_15235);
and U16540 (N_16540,N_15559,N_15100);
and U16541 (N_16541,N_15599,N_15845);
nor U16542 (N_16542,N_15751,N_15764);
or U16543 (N_16543,N_15928,N_15813);
or U16544 (N_16544,N_15964,N_15087);
nor U16545 (N_16545,N_15178,N_15725);
and U16546 (N_16546,N_15454,N_15386);
and U16547 (N_16547,N_15133,N_15754);
nand U16548 (N_16548,N_15920,N_15305);
nor U16549 (N_16549,N_15499,N_15943);
xnor U16550 (N_16550,N_15754,N_15267);
nor U16551 (N_16551,N_15596,N_15125);
xnor U16552 (N_16552,N_15632,N_15931);
nand U16553 (N_16553,N_15794,N_15592);
nor U16554 (N_16554,N_15983,N_15366);
and U16555 (N_16555,N_15046,N_15413);
nor U16556 (N_16556,N_15644,N_15855);
nand U16557 (N_16557,N_15710,N_15583);
and U16558 (N_16558,N_15743,N_15069);
or U16559 (N_16559,N_15694,N_15605);
or U16560 (N_16560,N_15404,N_15415);
or U16561 (N_16561,N_15291,N_15050);
xnor U16562 (N_16562,N_15087,N_15947);
nor U16563 (N_16563,N_15071,N_15548);
xor U16564 (N_16564,N_15799,N_15797);
nand U16565 (N_16565,N_15139,N_15352);
nand U16566 (N_16566,N_15569,N_15387);
nor U16567 (N_16567,N_15382,N_15398);
and U16568 (N_16568,N_15123,N_15938);
nor U16569 (N_16569,N_15652,N_15459);
and U16570 (N_16570,N_15715,N_15074);
nor U16571 (N_16571,N_15108,N_15417);
nor U16572 (N_16572,N_15205,N_15316);
or U16573 (N_16573,N_15265,N_15105);
or U16574 (N_16574,N_15028,N_15484);
and U16575 (N_16575,N_15205,N_15893);
nor U16576 (N_16576,N_15997,N_15954);
and U16577 (N_16577,N_15551,N_15353);
nand U16578 (N_16578,N_15875,N_15928);
nor U16579 (N_16579,N_15110,N_15820);
or U16580 (N_16580,N_15999,N_15297);
or U16581 (N_16581,N_15491,N_15125);
or U16582 (N_16582,N_15338,N_15614);
nor U16583 (N_16583,N_15177,N_15861);
or U16584 (N_16584,N_15280,N_15811);
nor U16585 (N_16585,N_15455,N_15415);
xor U16586 (N_16586,N_15199,N_15333);
or U16587 (N_16587,N_15714,N_15543);
and U16588 (N_16588,N_15006,N_15858);
nor U16589 (N_16589,N_15306,N_15916);
nand U16590 (N_16590,N_15313,N_15813);
and U16591 (N_16591,N_15562,N_15790);
or U16592 (N_16592,N_15168,N_15836);
nand U16593 (N_16593,N_15805,N_15611);
and U16594 (N_16594,N_15930,N_15111);
nor U16595 (N_16595,N_15277,N_15494);
xnor U16596 (N_16596,N_15235,N_15428);
or U16597 (N_16597,N_15710,N_15181);
nand U16598 (N_16598,N_15414,N_15695);
or U16599 (N_16599,N_15282,N_15518);
or U16600 (N_16600,N_15811,N_15489);
or U16601 (N_16601,N_15539,N_15356);
nand U16602 (N_16602,N_15792,N_15197);
and U16603 (N_16603,N_15670,N_15303);
or U16604 (N_16604,N_15876,N_15976);
nor U16605 (N_16605,N_15978,N_15056);
nor U16606 (N_16606,N_15026,N_15876);
nand U16607 (N_16607,N_15354,N_15966);
nand U16608 (N_16608,N_15981,N_15066);
xnor U16609 (N_16609,N_15446,N_15933);
xor U16610 (N_16610,N_15284,N_15228);
nand U16611 (N_16611,N_15238,N_15358);
nand U16612 (N_16612,N_15259,N_15837);
and U16613 (N_16613,N_15949,N_15367);
nand U16614 (N_16614,N_15101,N_15370);
nand U16615 (N_16615,N_15224,N_15958);
xor U16616 (N_16616,N_15727,N_15670);
nor U16617 (N_16617,N_15793,N_15822);
or U16618 (N_16618,N_15832,N_15456);
xor U16619 (N_16619,N_15978,N_15385);
and U16620 (N_16620,N_15294,N_15176);
nand U16621 (N_16621,N_15434,N_15795);
xor U16622 (N_16622,N_15026,N_15998);
and U16623 (N_16623,N_15540,N_15981);
nor U16624 (N_16624,N_15745,N_15012);
nor U16625 (N_16625,N_15222,N_15233);
and U16626 (N_16626,N_15875,N_15236);
nand U16627 (N_16627,N_15486,N_15603);
nor U16628 (N_16628,N_15183,N_15793);
xor U16629 (N_16629,N_15312,N_15640);
xnor U16630 (N_16630,N_15091,N_15673);
and U16631 (N_16631,N_15246,N_15605);
or U16632 (N_16632,N_15432,N_15019);
xnor U16633 (N_16633,N_15345,N_15022);
nand U16634 (N_16634,N_15605,N_15764);
nor U16635 (N_16635,N_15215,N_15231);
nor U16636 (N_16636,N_15706,N_15139);
nor U16637 (N_16637,N_15125,N_15225);
xor U16638 (N_16638,N_15997,N_15098);
or U16639 (N_16639,N_15544,N_15206);
and U16640 (N_16640,N_15753,N_15412);
xnor U16641 (N_16641,N_15647,N_15019);
or U16642 (N_16642,N_15332,N_15235);
nor U16643 (N_16643,N_15400,N_15331);
nor U16644 (N_16644,N_15522,N_15127);
xnor U16645 (N_16645,N_15684,N_15908);
nor U16646 (N_16646,N_15858,N_15395);
nand U16647 (N_16647,N_15992,N_15019);
nor U16648 (N_16648,N_15541,N_15277);
nor U16649 (N_16649,N_15954,N_15331);
nand U16650 (N_16650,N_15255,N_15976);
nor U16651 (N_16651,N_15915,N_15537);
nand U16652 (N_16652,N_15511,N_15002);
xor U16653 (N_16653,N_15422,N_15794);
xor U16654 (N_16654,N_15049,N_15760);
nor U16655 (N_16655,N_15430,N_15318);
or U16656 (N_16656,N_15767,N_15676);
xor U16657 (N_16657,N_15100,N_15458);
and U16658 (N_16658,N_15812,N_15826);
nor U16659 (N_16659,N_15385,N_15668);
and U16660 (N_16660,N_15845,N_15340);
xnor U16661 (N_16661,N_15659,N_15067);
xnor U16662 (N_16662,N_15603,N_15248);
nand U16663 (N_16663,N_15003,N_15184);
or U16664 (N_16664,N_15614,N_15013);
or U16665 (N_16665,N_15189,N_15003);
or U16666 (N_16666,N_15190,N_15292);
nor U16667 (N_16667,N_15351,N_15206);
or U16668 (N_16668,N_15155,N_15485);
nand U16669 (N_16669,N_15865,N_15791);
nand U16670 (N_16670,N_15853,N_15206);
xnor U16671 (N_16671,N_15648,N_15814);
nand U16672 (N_16672,N_15561,N_15094);
and U16673 (N_16673,N_15563,N_15207);
or U16674 (N_16674,N_15087,N_15756);
nor U16675 (N_16675,N_15540,N_15147);
xor U16676 (N_16676,N_15632,N_15655);
nor U16677 (N_16677,N_15254,N_15689);
xor U16678 (N_16678,N_15143,N_15776);
xnor U16679 (N_16679,N_15480,N_15656);
and U16680 (N_16680,N_15721,N_15147);
and U16681 (N_16681,N_15928,N_15204);
and U16682 (N_16682,N_15960,N_15707);
nor U16683 (N_16683,N_15310,N_15524);
nand U16684 (N_16684,N_15589,N_15977);
or U16685 (N_16685,N_15261,N_15937);
nor U16686 (N_16686,N_15125,N_15746);
nand U16687 (N_16687,N_15297,N_15710);
nor U16688 (N_16688,N_15036,N_15050);
xnor U16689 (N_16689,N_15480,N_15693);
nor U16690 (N_16690,N_15467,N_15162);
xnor U16691 (N_16691,N_15948,N_15177);
xor U16692 (N_16692,N_15366,N_15763);
nor U16693 (N_16693,N_15302,N_15935);
nor U16694 (N_16694,N_15643,N_15128);
or U16695 (N_16695,N_15588,N_15307);
xor U16696 (N_16696,N_15464,N_15009);
or U16697 (N_16697,N_15278,N_15354);
nor U16698 (N_16698,N_15538,N_15736);
nor U16699 (N_16699,N_15952,N_15372);
and U16700 (N_16700,N_15754,N_15009);
xnor U16701 (N_16701,N_15326,N_15567);
and U16702 (N_16702,N_15770,N_15134);
and U16703 (N_16703,N_15088,N_15734);
nand U16704 (N_16704,N_15026,N_15893);
xor U16705 (N_16705,N_15699,N_15194);
nor U16706 (N_16706,N_15713,N_15857);
nor U16707 (N_16707,N_15015,N_15118);
nor U16708 (N_16708,N_15095,N_15001);
nor U16709 (N_16709,N_15708,N_15826);
or U16710 (N_16710,N_15509,N_15107);
xnor U16711 (N_16711,N_15927,N_15195);
and U16712 (N_16712,N_15852,N_15468);
nor U16713 (N_16713,N_15417,N_15576);
and U16714 (N_16714,N_15463,N_15775);
and U16715 (N_16715,N_15134,N_15462);
and U16716 (N_16716,N_15396,N_15388);
or U16717 (N_16717,N_15290,N_15309);
nand U16718 (N_16718,N_15042,N_15332);
and U16719 (N_16719,N_15935,N_15257);
nor U16720 (N_16720,N_15856,N_15893);
xnor U16721 (N_16721,N_15051,N_15962);
or U16722 (N_16722,N_15340,N_15923);
xor U16723 (N_16723,N_15052,N_15325);
nor U16724 (N_16724,N_15503,N_15599);
or U16725 (N_16725,N_15524,N_15016);
nand U16726 (N_16726,N_15907,N_15857);
xor U16727 (N_16727,N_15029,N_15505);
nand U16728 (N_16728,N_15668,N_15946);
and U16729 (N_16729,N_15800,N_15346);
or U16730 (N_16730,N_15354,N_15943);
xnor U16731 (N_16731,N_15605,N_15784);
nor U16732 (N_16732,N_15517,N_15766);
nand U16733 (N_16733,N_15057,N_15412);
nor U16734 (N_16734,N_15362,N_15048);
nand U16735 (N_16735,N_15263,N_15273);
or U16736 (N_16736,N_15284,N_15708);
and U16737 (N_16737,N_15731,N_15253);
xor U16738 (N_16738,N_15580,N_15440);
xor U16739 (N_16739,N_15686,N_15129);
and U16740 (N_16740,N_15070,N_15751);
xnor U16741 (N_16741,N_15629,N_15692);
nand U16742 (N_16742,N_15797,N_15750);
xor U16743 (N_16743,N_15953,N_15390);
nand U16744 (N_16744,N_15776,N_15046);
or U16745 (N_16745,N_15982,N_15762);
and U16746 (N_16746,N_15376,N_15281);
or U16747 (N_16747,N_15908,N_15914);
or U16748 (N_16748,N_15158,N_15503);
nand U16749 (N_16749,N_15390,N_15303);
nand U16750 (N_16750,N_15567,N_15833);
or U16751 (N_16751,N_15933,N_15232);
and U16752 (N_16752,N_15628,N_15084);
xnor U16753 (N_16753,N_15177,N_15400);
or U16754 (N_16754,N_15215,N_15757);
nand U16755 (N_16755,N_15908,N_15598);
nand U16756 (N_16756,N_15421,N_15322);
xor U16757 (N_16757,N_15054,N_15565);
nand U16758 (N_16758,N_15665,N_15969);
nor U16759 (N_16759,N_15317,N_15707);
and U16760 (N_16760,N_15889,N_15387);
nand U16761 (N_16761,N_15647,N_15769);
xnor U16762 (N_16762,N_15738,N_15149);
nor U16763 (N_16763,N_15506,N_15380);
and U16764 (N_16764,N_15291,N_15145);
and U16765 (N_16765,N_15555,N_15041);
nand U16766 (N_16766,N_15942,N_15048);
or U16767 (N_16767,N_15590,N_15632);
or U16768 (N_16768,N_15446,N_15188);
or U16769 (N_16769,N_15727,N_15244);
xor U16770 (N_16770,N_15033,N_15000);
xor U16771 (N_16771,N_15203,N_15172);
xnor U16772 (N_16772,N_15659,N_15542);
xnor U16773 (N_16773,N_15668,N_15250);
or U16774 (N_16774,N_15122,N_15651);
nand U16775 (N_16775,N_15895,N_15088);
xor U16776 (N_16776,N_15221,N_15869);
nand U16777 (N_16777,N_15204,N_15821);
and U16778 (N_16778,N_15911,N_15410);
nor U16779 (N_16779,N_15342,N_15605);
nand U16780 (N_16780,N_15854,N_15754);
and U16781 (N_16781,N_15239,N_15061);
xnor U16782 (N_16782,N_15230,N_15150);
xnor U16783 (N_16783,N_15711,N_15549);
nand U16784 (N_16784,N_15906,N_15551);
and U16785 (N_16785,N_15636,N_15162);
xnor U16786 (N_16786,N_15113,N_15123);
nand U16787 (N_16787,N_15416,N_15798);
or U16788 (N_16788,N_15792,N_15211);
and U16789 (N_16789,N_15070,N_15393);
or U16790 (N_16790,N_15863,N_15633);
nand U16791 (N_16791,N_15935,N_15644);
and U16792 (N_16792,N_15977,N_15775);
xor U16793 (N_16793,N_15421,N_15721);
xnor U16794 (N_16794,N_15501,N_15443);
nor U16795 (N_16795,N_15144,N_15696);
nor U16796 (N_16796,N_15672,N_15401);
nor U16797 (N_16797,N_15721,N_15397);
and U16798 (N_16798,N_15067,N_15442);
nor U16799 (N_16799,N_15097,N_15716);
or U16800 (N_16800,N_15238,N_15225);
nand U16801 (N_16801,N_15416,N_15642);
and U16802 (N_16802,N_15510,N_15452);
nor U16803 (N_16803,N_15142,N_15404);
xnor U16804 (N_16804,N_15052,N_15802);
nor U16805 (N_16805,N_15491,N_15133);
nor U16806 (N_16806,N_15062,N_15429);
or U16807 (N_16807,N_15878,N_15605);
or U16808 (N_16808,N_15896,N_15132);
nor U16809 (N_16809,N_15752,N_15638);
nor U16810 (N_16810,N_15139,N_15564);
nand U16811 (N_16811,N_15328,N_15082);
nor U16812 (N_16812,N_15290,N_15406);
nand U16813 (N_16813,N_15573,N_15109);
nor U16814 (N_16814,N_15822,N_15580);
nor U16815 (N_16815,N_15828,N_15366);
nor U16816 (N_16816,N_15856,N_15036);
xor U16817 (N_16817,N_15326,N_15860);
nor U16818 (N_16818,N_15945,N_15115);
and U16819 (N_16819,N_15498,N_15049);
or U16820 (N_16820,N_15138,N_15166);
or U16821 (N_16821,N_15427,N_15129);
xnor U16822 (N_16822,N_15375,N_15920);
and U16823 (N_16823,N_15625,N_15354);
nor U16824 (N_16824,N_15748,N_15181);
nor U16825 (N_16825,N_15034,N_15576);
or U16826 (N_16826,N_15317,N_15736);
nor U16827 (N_16827,N_15192,N_15142);
nand U16828 (N_16828,N_15031,N_15182);
and U16829 (N_16829,N_15679,N_15113);
nand U16830 (N_16830,N_15818,N_15051);
xor U16831 (N_16831,N_15427,N_15926);
or U16832 (N_16832,N_15276,N_15503);
xnor U16833 (N_16833,N_15365,N_15925);
or U16834 (N_16834,N_15099,N_15803);
nand U16835 (N_16835,N_15137,N_15760);
nand U16836 (N_16836,N_15467,N_15053);
nand U16837 (N_16837,N_15749,N_15144);
and U16838 (N_16838,N_15602,N_15463);
nor U16839 (N_16839,N_15111,N_15420);
and U16840 (N_16840,N_15211,N_15932);
or U16841 (N_16841,N_15749,N_15774);
nand U16842 (N_16842,N_15753,N_15120);
xnor U16843 (N_16843,N_15033,N_15264);
or U16844 (N_16844,N_15953,N_15643);
nand U16845 (N_16845,N_15237,N_15636);
nor U16846 (N_16846,N_15443,N_15602);
and U16847 (N_16847,N_15804,N_15118);
or U16848 (N_16848,N_15289,N_15929);
or U16849 (N_16849,N_15803,N_15002);
nor U16850 (N_16850,N_15279,N_15072);
nand U16851 (N_16851,N_15203,N_15408);
or U16852 (N_16852,N_15197,N_15665);
nand U16853 (N_16853,N_15401,N_15546);
nor U16854 (N_16854,N_15391,N_15968);
nor U16855 (N_16855,N_15668,N_15176);
or U16856 (N_16856,N_15429,N_15960);
nor U16857 (N_16857,N_15198,N_15099);
nand U16858 (N_16858,N_15146,N_15423);
and U16859 (N_16859,N_15384,N_15619);
or U16860 (N_16860,N_15470,N_15791);
nand U16861 (N_16861,N_15984,N_15857);
or U16862 (N_16862,N_15693,N_15605);
nand U16863 (N_16863,N_15661,N_15336);
nor U16864 (N_16864,N_15008,N_15448);
nand U16865 (N_16865,N_15946,N_15043);
or U16866 (N_16866,N_15818,N_15206);
or U16867 (N_16867,N_15102,N_15065);
nand U16868 (N_16868,N_15048,N_15956);
nand U16869 (N_16869,N_15772,N_15065);
or U16870 (N_16870,N_15447,N_15569);
nand U16871 (N_16871,N_15521,N_15666);
nand U16872 (N_16872,N_15974,N_15016);
and U16873 (N_16873,N_15766,N_15561);
xnor U16874 (N_16874,N_15180,N_15098);
nand U16875 (N_16875,N_15877,N_15558);
and U16876 (N_16876,N_15107,N_15319);
or U16877 (N_16877,N_15341,N_15579);
and U16878 (N_16878,N_15621,N_15622);
or U16879 (N_16879,N_15965,N_15780);
xor U16880 (N_16880,N_15817,N_15266);
nor U16881 (N_16881,N_15558,N_15682);
nor U16882 (N_16882,N_15530,N_15813);
nor U16883 (N_16883,N_15522,N_15412);
or U16884 (N_16884,N_15749,N_15736);
nor U16885 (N_16885,N_15338,N_15092);
or U16886 (N_16886,N_15074,N_15815);
nor U16887 (N_16887,N_15443,N_15784);
and U16888 (N_16888,N_15839,N_15116);
and U16889 (N_16889,N_15579,N_15089);
or U16890 (N_16890,N_15366,N_15424);
or U16891 (N_16891,N_15495,N_15959);
xnor U16892 (N_16892,N_15687,N_15619);
nand U16893 (N_16893,N_15709,N_15751);
or U16894 (N_16894,N_15295,N_15556);
and U16895 (N_16895,N_15659,N_15284);
xnor U16896 (N_16896,N_15035,N_15156);
and U16897 (N_16897,N_15704,N_15565);
and U16898 (N_16898,N_15674,N_15047);
nand U16899 (N_16899,N_15215,N_15856);
nand U16900 (N_16900,N_15092,N_15130);
nand U16901 (N_16901,N_15359,N_15468);
nor U16902 (N_16902,N_15831,N_15644);
or U16903 (N_16903,N_15647,N_15657);
xnor U16904 (N_16904,N_15037,N_15596);
nor U16905 (N_16905,N_15772,N_15142);
nand U16906 (N_16906,N_15096,N_15622);
and U16907 (N_16907,N_15067,N_15322);
xor U16908 (N_16908,N_15111,N_15293);
or U16909 (N_16909,N_15548,N_15474);
nand U16910 (N_16910,N_15270,N_15796);
nor U16911 (N_16911,N_15853,N_15596);
nor U16912 (N_16912,N_15930,N_15140);
nor U16913 (N_16913,N_15949,N_15467);
nor U16914 (N_16914,N_15682,N_15942);
or U16915 (N_16915,N_15875,N_15327);
and U16916 (N_16916,N_15229,N_15961);
nand U16917 (N_16917,N_15070,N_15381);
nand U16918 (N_16918,N_15795,N_15717);
or U16919 (N_16919,N_15605,N_15054);
xor U16920 (N_16920,N_15288,N_15980);
xnor U16921 (N_16921,N_15950,N_15037);
nand U16922 (N_16922,N_15665,N_15173);
nor U16923 (N_16923,N_15496,N_15501);
nor U16924 (N_16924,N_15089,N_15879);
nand U16925 (N_16925,N_15048,N_15769);
and U16926 (N_16926,N_15924,N_15817);
nor U16927 (N_16927,N_15115,N_15119);
nor U16928 (N_16928,N_15518,N_15053);
nor U16929 (N_16929,N_15223,N_15096);
xor U16930 (N_16930,N_15153,N_15948);
nand U16931 (N_16931,N_15546,N_15738);
and U16932 (N_16932,N_15354,N_15500);
and U16933 (N_16933,N_15316,N_15381);
or U16934 (N_16934,N_15558,N_15478);
or U16935 (N_16935,N_15989,N_15475);
nor U16936 (N_16936,N_15027,N_15337);
nand U16937 (N_16937,N_15797,N_15765);
or U16938 (N_16938,N_15423,N_15045);
nor U16939 (N_16939,N_15385,N_15858);
nand U16940 (N_16940,N_15850,N_15858);
nor U16941 (N_16941,N_15504,N_15074);
xnor U16942 (N_16942,N_15391,N_15378);
xnor U16943 (N_16943,N_15421,N_15907);
nor U16944 (N_16944,N_15279,N_15759);
and U16945 (N_16945,N_15760,N_15388);
and U16946 (N_16946,N_15083,N_15117);
nor U16947 (N_16947,N_15767,N_15210);
nor U16948 (N_16948,N_15280,N_15161);
nor U16949 (N_16949,N_15380,N_15122);
or U16950 (N_16950,N_15853,N_15520);
xor U16951 (N_16951,N_15809,N_15762);
nand U16952 (N_16952,N_15814,N_15088);
xnor U16953 (N_16953,N_15795,N_15205);
nand U16954 (N_16954,N_15932,N_15998);
nor U16955 (N_16955,N_15520,N_15610);
and U16956 (N_16956,N_15201,N_15249);
and U16957 (N_16957,N_15914,N_15616);
nor U16958 (N_16958,N_15140,N_15542);
nor U16959 (N_16959,N_15496,N_15621);
xnor U16960 (N_16960,N_15039,N_15296);
xor U16961 (N_16961,N_15609,N_15021);
or U16962 (N_16962,N_15094,N_15371);
or U16963 (N_16963,N_15741,N_15853);
nor U16964 (N_16964,N_15864,N_15163);
xor U16965 (N_16965,N_15567,N_15987);
or U16966 (N_16966,N_15168,N_15094);
nor U16967 (N_16967,N_15360,N_15563);
or U16968 (N_16968,N_15884,N_15597);
nand U16969 (N_16969,N_15484,N_15987);
nor U16970 (N_16970,N_15683,N_15974);
nand U16971 (N_16971,N_15648,N_15947);
xnor U16972 (N_16972,N_15111,N_15717);
nor U16973 (N_16973,N_15191,N_15490);
xor U16974 (N_16974,N_15807,N_15757);
and U16975 (N_16975,N_15997,N_15708);
nand U16976 (N_16976,N_15423,N_15135);
nor U16977 (N_16977,N_15163,N_15871);
or U16978 (N_16978,N_15214,N_15885);
nand U16979 (N_16979,N_15173,N_15217);
nand U16980 (N_16980,N_15653,N_15331);
or U16981 (N_16981,N_15708,N_15743);
xnor U16982 (N_16982,N_15047,N_15446);
or U16983 (N_16983,N_15582,N_15027);
nor U16984 (N_16984,N_15673,N_15738);
nor U16985 (N_16985,N_15438,N_15056);
nand U16986 (N_16986,N_15806,N_15626);
nor U16987 (N_16987,N_15429,N_15894);
and U16988 (N_16988,N_15584,N_15868);
nand U16989 (N_16989,N_15945,N_15633);
xor U16990 (N_16990,N_15831,N_15095);
xnor U16991 (N_16991,N_15098,N_15544);
xor U16992 (N_16992,N_15131,N_15088);
nand U16993 (N_16993,N_15127,N_15991);
nor U16994 (N_16994,N_15816,N_15808);
xor U16995 (N_16995,N_15564,N_15817);
and U16996 (N_16996,N_15541,N_15941);
and U16997 (N_16997,N_15997,N_15791);
and U16998 (N_16998,N_15764,N_15238);
xnor U16999 (N_16999,N_15345,N_15565);
and U17000 (N_17000,N_16919,N_16446);
nand U17001 (N_17001,N_16754,N_16966);
nor U17002 (N_17002,N_16553,N_16421);
or U17003 (N_17003,N_16520,N_16471);
xor U17004 (N_17004,N_16793,N_16029);
or U17005 (N_17005,N_16870,N_16608);
nor U17006 (N_17006,N_16698,N_16363);
or U17007 (N_17007,N_16210,N_16152);
or U17008 (N_17008,N_16240,N_16759);
or U17009 (N_17009,N_16319,N_16587);
xor U17010 (N_17010,N_16264,N_16565);
xor U17011 (N_17011,N_16099,N_16519);
or U17012 (N_17012,N_16756,N_16622);
nor U17013 (N_17013,N_16073,N_16493);
or U17014 (N_17014,N_16418,N_16991);
or U17015 (N_17015,N_16138,N_16393);
xnor U17016 (N_17016,N_16570,N_16525);
nor U17017 (N_17017,N_16299,N_16241);
nor U17018 (N_17018,N_16344,N_16464);
and U17019 (N_17019,N_16329,N_16889);
nand U17020 (N_17020,N_16150,N_16262);
nand U17021 (N_17021,N_16239,N_16287);
nand U17022 (N_17022,N_16310,N_16107);
xor U17023 (N_17023,N_16528,N_16989);
and U17024 (N_17024,N_16395,N_16088);
and U17025 (N_17025,N_16452,N_16591);
xnor U17026 (N_17026,N_16062,N_16868);
xor U17027 (N_17027,N_16423,N_16821);
and U17028 (N_17028,N_16653,N_16281);
or U17029 (N_17029,N_16635,N_16920);
or U17030 (N_17030,N_16361,N_16054);
xnor U17031 (N_17031,N_16067,N_16223);
and U17032 (N_17032,N_16752,N_16709);
and U17033 (N_17033,N_16804,N_16613);
nor U17034 (N_17034,N_16391,N_16888);
nor U17035 (N_17035,N_16585,N_16031);
xor U17036 (N_17036,N_16738,N_16964);
xnor U17037 (N_17037,N_16288,N_16069);
nor U17038 (N_17038,N_16090,N_16135);
or U17039 (N_17039,N_16339,N_16245);
nand U17040 (N_17040,N_16687,N_16316);
xor U17041 (N_17041,N_16522,N_16753);
and U17042 (N_17042,N_16774,N_16488);
nor U17043 (N_17043,N_16662,N_16259);
nor U17044 (N_17044,N_16872,N_16751);
xnor U17045 (N_17045,N_16289,N_16524);
or U17046 (N_17046,N_16517,N_16529);
nor U17047 (N_17047,N_16096,N_16768);
nor U17048 (N_17048,N_16030,N_16449);
and U17049 (N_17049,N_16475,N_16847);
nor U17050 (N_17050,N_16283,N_16611);
and U17051 (N_17051,N_16624,N_16006);
xnor U17052 (N_17052,N_16408,N_16185);
and U17053 (N_17053,N_16175,N_16448);
xor U17054 (N_17054,N_16468,N_16645);
nor U17055 (N_17055,N_16479,N_16829);
and U17056 (N_17056,N_16817,N_16758);
nor U17057 (N_17057,N_16658,N_16132);
nor U17058 (N_17058,N_16322,N_16762);
and U17059 (N_17059,N_16595,N_16318);
nor U17060 (N_17060,N_16231,N_16269);
or U17061 (N_17061,N_16302,N_16313);
nand U17062 (N_17062,N_16673,N_16696);
nand U17063 (N_17063,N_16236,N_16828);
nand U17064 (N_17064,N_16874,N_16140);
nand U17065 (N_17065,N_16854,N_16807);
and U17066 (N_17066,N_16757,N_16438);
nand U17067 (N_17067,N_16413,N_16497);
nor U17068 (N_17068,N_16101,N_16199);
xor U17069 (N_17069,N_16548,N_16005);
nand U17070 (N_17070,N_16426,N_16655);
or U17071 (N_17071,N_16536,N_16945);
nand U17072 (N_17072,N_16083,N_16389);
nand U17073 (N_17073,N_16461,N_16184);
nand U17074 (N_17074,N_16098,N_16417);
xnor U17075 (N_17075,N_16230,N_16061);
and U17076 (N_17076,N_16415,N_16977);
and U17077 (N_17077,N_16727,N_16547);
and U17078 (N_17078,N_16345,N_16050);
or U17079 (N_17079,N_16782,N_16711);
and U17080 (N_17080,N_16370,N_16952);
xor U17081 (N_17081,N_16484,N_16351);
nor U17082 (N_17082,N_16725,N_16724);
xor U17083 (N_17083,N_16158,N_16542);
nand U17084 (N_17084,N_16082,N_16374);
nand U17085 (N_17085,N_16350,N_16496);
or U17086 (N_17086,N_16961,N_16197);
xor U17087 (N_17087,N_16047,N_16016);
or U17088 (N_17088,N_16720,N_16642);
nor U17089 (N_17089,N_16348,N_16632);
nor U17090 (N_17090,N_16789,N_16224);
nand U17091 (N_17091,N_16671,N_16597);
nand U17092 (N_17092,N_16242,N_16078);
nor U17093 (N_17093,N_16124,N_16060);
and U17094 (N_17094,N_16271,N_16787);
xnor U17095 (N_17095,N_16692,N_16155);
xnor U17096 (N_17096,N_16649,N_16890);
and U17097 (N_17097,N_16809,N_16434);
or U17098 (N_17098,N_16499,N_16786);
or U17099 (N_17099,N_16588,N_16358);
and U17100 (N_17100,N_16730,N_16041);
nand U17101 (N_17101,N_16561,N_16250);
and U17102 (N_17102,N_16676,N_16081);
nand U17103 (N_17103,N_16353,N_16679);
xnor U17104 (N_17104,N_16557,N_16644);
nand U17105 (N_17105,N_16229,N_16760);
or U17106 (N_17106,N_16396,N_16965);
or U17107 (N_17107,N_16215,N_16397);
and U17108 (N_17108,N_16707,N_16309);
xor U17109 (N_17109,N_16144,N_16274);
nand U17110 (N_17110,N_16718,N_16902);
or U17111 (N_17111,N_16867,N_16182);
xor U17112 (N_17112,N_16303,N_16306);
nor U17113 (N_17113,N_16295,N_16770);
nand U17114 (N_17114,N_16656,N_16168);
or U17115 (N_17115,N_16490,N_16097);
or U17116 (N_17116,N_16717,N_16279);
nor U17117 (N_17117,N_16944,N_16857);
xnor U17118 (N_17118,N_16292,N_16716);
nor U17119 (N_17119,N_16648,N_16129);
xor U17120 (N_17120,N_16419,N_16428);
and U17121 (N_17121,N_16327,N_16494);
and U17122 (N_17122,N_16476,N_16880);
or U17123 (N_17123,N_16071,N_16256);
nand U17124 (N_17124,N_16684,N_16704);
or U17125 (N_17125,N_16905,N_16399);
nand U17126 (N_17126,N_16409,N_16743);
nand U17127 (N_17127,N_16599,N_16922);
nor U17128 (N_17128,N_16291,N_16928);
xnor U17129 (N_17129,N_16609,N_16560);
or U17130 (N_17130,N_16102,N_16992);
and U17131 (N_17131,N_16228,N_16394);
nand U17132 (N_17132,N_16092,N_16219);
nor U17133 (N_17133,N_16507,N_16474);
nand U17134 (N_17134,N_16906,N_16504);
or U17135 (N_17135,N_16003,N_16436);
nand U17136 (N_17136,N_16012,N_16921);
or U17137 (N_17137,N_16123,N_16206);
nor U17138 (N_17138,N_16544,N_16951);
nor U17139 (N_17139,N_16583,N_16487);
nor U17140 (N_17140,N_16830,N_16312);
nor U17141 (N_17141,N_16975,N_16871);
xor U17142 (N_17142,N_16806,N_16369);
or U17143 (N_17143,N_16148,N_16639);
nand U17144 (N_17144,N_16328,N_16246);
xnor U17145 (N_17145,N_16967,N_16424);
or U17146 (N_17146,N_16217,N_16796);
and U17147 (N_17147,N_16546,N_16483);
or U17148 (N_17148,N_16015,N_16323);
nand U17149 (N_17149,N_16297,N_16443);
and U17150 (N_17150,N_16926,N_16066);
nor U17151 (N_17151,N_16338,N_16925);
nand U17152 (N_17152,N_16664,N_16349);
and U17153 (N_17153,N_16188,N_16201);
and U17154 (N_17154,N_16477,N_16521);
nor U17155 (N_17155,N_16315,N_16916);
xnor U17156 (N_17156,N_16437,N_16462);
xnor U17157 (N_17157,N_16892,N_16482);
xor U17158 (N_17158,N_16994,N_16359);
xor U17159 (N_17159,N_16453,N_16190);
nand U17160 (N_17160,N_16347,N_16111);
nor U17161 (N_17161,N_16933,N_16332);
xor U17162 (N_17162,N_16205,N_16420);
nor U17163 (N_17163,N_16669,N_16068);
xor U17164 (N_17164,N_16954,N_16136);
nand U17165 (N_17165,N_16552,N_16341);
nand U17166 (N_17166,N_16272,N_16680);
nor U17167 (N_17167,N_16538,N_16032);
xnor U17168 (N_17168,N_16678,N_16234);
xor U17169 (N_17169,N_16105,N_16910);
xor U17170 (N_17170,N_16220,N_16076);
or U17171 (N_17171,N_16859,N_16070);
and U17172 (N_17172,N_16600,N_16625);
or U17173 (N_17173,N_16741,N_16263);
nor U17174 (N_17174,N_16130,N_16275);
nor U17175 (N_17175,N_16444,N_16960);
and U17176 (N_17176,N_16675,N_16566);
and U17177 (N_17177,N_16017,N_16674);
nor U17178 (N_17178,N_16790,N_16976);
or U17179 (N_17179,N_16710,N_16573);
or U17180 (N_17180,N_16203,N_16589);
nand U17181 (N_17181,N_16955,N_16593);
xnor U17182 (N_17182,N_16917,N_16534);
and U17183 (N_17183,N_16844,N_16503);
xnor U17184 (N_17184,N_16677,N_16610);
nand U17185 (N_17185,N_16657,N_16875);
nand U17186 (N_17186,N_16192,N_16747);
nor U17187 (N_17187,N_16151,N_16265);
xor U17188 (N_17188,N_16301,N_16093);
nor U17189 (N_17189,N_16783,N_16849);
and U17190 (N_17190,N_16109,N_16887);
nor U17191 (N_17191,N_16576,N_16586);
nor U17192 (N_17192,N_16941,N_16178);
or U17193 (N_17193,N_16400,N_16043);
xnor U17194 (N_17194,N_16280,N_16267);
xnor U17195 (N_17195,N_16851,N_16154);
and U17196 (N_17196,N_16072,N_16654);
nand U17197 (N_17197,N_16159,N_16311);
nand U17198 (N_17198,N_16581,N_16442);
nor U17199 (N_17199,N_16968,N_16131);
or U17200 (N_17200,N_16958,N_16174);
nand U17201 (N_17201,N_16321,N_16149);
and U17202 (N_17202,N_16579,N_16033);
and U17203 (N_17203,N_16406,N_16024);
nand U17204 (N_17204,N_16104,N_16000);
nand U17205 (N_17205,N_16571,N_16886);
and U17206 (N_17206,N_16640,N_16455);
nor U17207 (N_17207,N_16688,N_16606);
and U17208 (N_17208,N_16682,N_16286);
and U17209 (N_17209,N_16626,N_16852);
nand U17210 (N_17210,N_16835,N_16085);
or U17211 (N_17211,N_16700,N_16660);
and U17212 (N_17212,N_16163,N_16532);
or U17213 (N_17213,N_16162,N_16866);
or U17214 (N_17214,N_16337,N_16858);
and U17215 (N_17215,N_16294,N_16403);
or U17216 (N_17216,N_16410,N_16196);
xnor U17217 (N_17217,N_16284,N_16414);
and U17218 (N_17218,N_16861,N_16079);
nand U17219 (N_17219,N_16077,N_16094);
xnor U17220 (N_17220,N_16742,N_16946);
xor U17221 (N_17221,N_16038,N_16918);
or U17222 (N_17222,N_16346,N_16034);
and U17223 (N_17223,N_16198,N_16822);
xnor U17224 (N_17224,N_16364,N_16422);
or U17225 (N_17225,N_16512,N_16802);
xnor U17226 (N_17226,N_16384,N_16333);
nand U17227 (N_17227,N_16266,N_16372);
and U17228 (N_17228,N_16630,N_16900);
xnor U17229 (N_17229,N_16736,N_16371);
nor U17230 (N_17230,N_16035,N_16164);
nand U17231 (N_17231,N_16848,N_16993);
xnor U17232 (N_17232,N_16996,N_16990);
nor U17233 (N_17233,N_16686,N_16411);
nor U17234 (N_17234,N_16506,N_16550);
xor U17235 (N_17235,N_16053,N_16979);
nand U17236 (N_17236,N_16074,N_16904);
and U17237 (N_17237,N_16431,N_16556);
or U17238 (N_17238,N_16026,N_16878);
nor U17239 (N_17239,N_16732,N_16100);
and U17240 (N_17240,N_16873,N_16939);
or U17241 (N_17241,N_16084,N_16114);
or U17242 (N_17242,N_16143,N_16458);
or U17243 (N_17243,N_16763,N_16260);
xor U17244 (N_17244,N_16794,N_16145);
nand U17245 (N_17245,N_16883,N_16354);
nor U17246 (N_17246,N_16691,N_16180);
and U17247 (N_17247,N_16832,N_16620);
or U17248 (N_17248,N_16278,N_16235);
nand U17249 (N_17249,N_16983,N_16931);
xnor U17250 (N_17250,N_16864,N_16059);
xor U17251 (N_17251,N_16469,N_16563);
or U17252 (N_17252,N_16950,N_16028);
nand U17253 (N_17253,N_16969,N_16695);
nor U17254 (N_17254,N_16670,N_16018);
and U17255 (N_17255,N_16480,N_16478);
xor U17256 (N_17256,N_16533,N_16456);
nand U17257 (N_17257,N_16784,N_16492);
and U17258 (N_17258,N_16451,N_16010);
or U17259 (N_17259,N_16202,N_16011);
xnor U17260 (N_17260,N_16971,N_16980);
nor U17261 (N_17261,N_16491,N_16986);
xnor U17262 (N_17262,N_16590,N_16631);
xnor U17263 (N_17263,N_16209,N_16767);
nor U17264 (N_17264,N_16304,N_16666);
nand U17265 (N_17265,N_16814,N_16334);
and U17266 (N_17266,N_16603,N_16366);
nand U17267 (N_17267,N_16080,N_16501);
nor U17268 (N_17268,N_16340,N_16853);
and U17269 (N_17269,N_16799,N_16997);
and U17270 (N_17270,N_16237,N_16013);
or U17271 (N_17271,N_16596,N_16020);
xnor U17272 (N_17272,N_16156,N_16834);
nand U17273 (N_17273,N_16728,N_16863);
nand U17274 (N_17274,N_16661,N_16002);
nand U17275 (N_17275,N_16489,N_16619);
nor U17276 (N_17276,N_16392,N_16785);
nor U17277 (N_17277,N_16296,N_16379);
nor U17278 (N_17278,N_16485,N_16745);
or U17279 (N_17279,N_16126,N_16502);
or U17280 (N_17280,N_16058,N_16122);
xor U17281 (N_17281,N_16731,N_16580);
xor U17282 (N_17282,N_16116,N_16412);
or U17283 (N_17283,N_16541,N_16911);
or U17284 (N_17284,N_16694,N_16470);
nand U17285 (N_17285,N_16404,N_16244);
nor U17286 (N_17286,N_16025,N_16282);
nand U17287 (N_17287,N_16831,N_16427);
nor U17288 (N_17288,N_16447,N_16120);
and U17289 (N_17289,N_16232,N_16841);
and U17290 (N_17290,N_16153,N_16401);
and U17291 (N_17291,N_16936,N_16803);
nand U17292 (N_17292,N_16293,N_16598);
xor U17293 (N_17293,N_16134,N_16454);
nand U17294 (N_17294,N_16326,N_16450);
xor U17295 (N_17295,N_16169,N_16562);
nor U17296 (N_17296,N_16923,N_16137);
or U17297 (N_17297,N_16646,N_16027);
xnor U17298 (N_17298,N_16530,N_16022);
nand U17299 (N_17299,N_16974,N_16559);
or U17300 (N_17300,N_16368,N_16750);
and U17301 (N_17301,N_16051,N_16064);
nand U17302 (N_17302,N_16091,N_16445);
nor U17303 (N_17303,N_16914,N_16697);
nand U17304 (N_17304,N_16771,N_16825);
or U17305 (N_17305,N_16765,N_16367);
xor U17306 (N_17306,N_16407,N_16811);
nand U17307 (N_17307,N_16773,N_16518);
nor U17308 (N_17308,N_16865,N_16171);
xnor U17309 (N_17309,N_16042,N_16247);
xnor U17310 (N_17310,N_16769,N_16672);
nor U17311 (N_17311,N_16932,N_16176);
nand U17312 (N_17312,N_16509,N_16930);
nand U17313 (N_17313,N_16737,N_16584);
nand U17314 (N_17314,N_16810,N_16170);
nand U17315 (N_17315,N_16879,N_16141);
xor U17316 (N_17316,N_16699,N_16276);
or U17317 (N_17317,N_16935,N_16009);
xnor U17318 (N_17318,N_16740,N_16924);
or U17319 (N_17319,N_16435,N_16390);
and U17320 (N_17320,N_16008,N_16972);
xnor U17321 (N_17321,N_16860,N_16195);
xor U17322 (N_17322,N_16252,N_16856);
nand U17323 (N_17323,N_16194,N_16947);
xnor U17324 (N_17324,N_16837,N_16592);
xor U17325 (N_17325,N_16405,N_16824);
nand U17326 (N_17326,N_16998,N_16113);
xnor U17327 (N_17327,N_16615,N_16987);
or U17328 (N_17328,N_16881,N_16508);
nand U17329 (N_17329,N_16956,N_16617);
nand U17330 (N_17330,N_16948,N_16708);
nor U17331 (N_17331,N_16602,N_16795);
nand U17332 (N_17332,N_16995,N_16441);
nor U17333 (N_17333,N_16183,N_16087);
or U17334 (N_17334,N_16416,N_16940);
xor U17335 (N_17335,N_16776,N_16999);
nand U17336 (N_17336,N_16775,N_16398);
xnor U17337 (N_17337,N_16285,N_16385);
and U17338 (N_17338,N_16962,N_16612);
nor U17339 (N_17339,N_16929,N_16057);
or U17340 (N_17340,N_16685,N_16733);
nor U17341 (N_17341,N_16121,N_16526);
xor U17342 (N_17342,N_16869,N_16147);
or U17343 (N_17343,N_16040,N_16665);
or U17344 (N_17344,N_16701,N_16815);
and U17345 (N_17345,N_16212,N_16772);
nor U17346 (N_17346,N_16894,N_16360);
and U17347 (N_17347,N_16937,N_16627);
xnor U17348 (N_17348,N_16749,N_16179);
nand U17349 (N_17349,N_16706,N_16459);
and U17350 (N_17350,N_16637,N_16204);
xnor U17351 (N_17351,N_16375,N_16982);
nor U17352 (N_17352,N_16623,N_16387);
nor U17353 (N_17353,N_16988,N_16118);
or U17354 (N_17354,N_16643,N_16248);
nand U17355 (N_17355,N_16689,N_16049);
and U17356 (N_17356,N_16290,N_16934);
xnor U17357 (N_17357,N_16693,N_16128);
xor U17358 (N_17358,N_16957,N_16777);
and U17359 (N_17359,N_16908,N_16125);
xnor U17360 (N_17360,N_16298,N_16086);
xnor U17361 (N_17361,N_16177,N_16915);
nand U17362 (N_17362,N_16255,N_16495);
nor U17363 (N_17363,N_16568,N_16913);
nor U17364 (N_17364,N_16582,N_16705);
and U17365 (N_17365,N_16575,N_16505);
nor U17366 (N_17366,N_16226,N_16621);
or U17367 (N_17367,N_16840,N_16882);
or U17368 (N_17368,N_16211,N_16681);
nor U17369 (N_17369,N_16305,N_16667);
nand U17370 (N_17370,N_16901,N_16792);
and U17371 (N_17371,N_16095,N_16780);
nor U17372 (N_17372,N_16187,N_16253);
or U17373 (N_17373,N_16554,N_16055);
or U17374 (N_17374,N_16540,N_16778);
xor U17375 (N_17375,N_16139,N_16324);
and U17376 (N_17376,N_16007,N_16897);
nand U17377 (N_17377,N_16895,N_16636);
or U17378 (N_17378,N_16300,N_16891);
or U17379 (N_17379,N_16373,N_16826);
and U17380 (N_17380,N_16335,N_16764);
nor U17381 (N_17381,N_16896,N_16791);
nor U17382 (N_17382,N_16044,N_16052);
xor U17383 (N_17383,N_16021,N_16641);
nor U17384 (N_17384,N_16167,N_16089);
or U17385 (N_17385,N_16207,N_16261);
and U17386 (N_17386,N_16605,N_16473);
nand U17387 (N_17387,N_16112,N_16330);
nand U17388 (N_17388,N_16616,N_16481);
or U17389 (N_17389,N_16110,N_16193);
and U17390 (N_17390,N_16486,N_16208);
nand U17391 (N_17391,N_16981,N_16703);
or U17392 (N_17392,N_16739,N_16165);
nor U17393 (N_17393,N_16903,N_16383);
or U17394 (N_17394,N_16663,N_16818);
xnor U17395 (N_17395,N_16307,N_16045);
xor U17396 (N_17396,N_16761,N_16713);
or U17397 (N_17397,N_16376,N_16885);
nor U17398 (N_17398,N_16225,N_16943);
and U17399 (N_17399,N_16065,N_16801);
and U17400 (N_17400,N_16516,N_16734);
xor U17401 (N_17401,N_16146,N_16877);
nand U17402 (N_17402,N_16117,N_16800);
xnor U17403 (N_17403,N_16722,N_16317);
and U17404 (N_17404,N_16628,N_16647);
nand U17405 (N_17405,N_16798,N_16222);
or U17406 (N_17406,N_16651,N_16467);
nand U17407 (N_17407,N_16823,N_16555);
or U17408 (N_17408,N_16604,N_16650);
nand U17409 (N_17409,N_16172,N_16004);
nand U17410 (N_17410,N_16106,N_16909);
nor U17411 (N_17411,N_16214,N_16254);
nor U17412 (N_17412,N_16320,N_16539);
or U17413 (N_17413,N_16668,N_16463);
xor U17414 (N_17414,N_16001,N_16978);
xnor U17415 (N_17415,N_16515,N_16161);
xnor U17416 (N_17416,N_16166,N_16607);
xnor U17417 (N_17417,N_16963,N_16249);
nor U17418 (N_17418,N_16046,N_16633);
nor U17419 (N_17419,N_16659,N_16820);
nor U17420 (N_17420,N_16465,N_16514);
xnor U17421 (N_17421,N_16381,N_16543);
or U17422 (N_17422,N_16277,N_16838);
nor U17423 (N_17423,N_16862,N_16402);
and U17424 (N_17424,N_16523,N_16014);
and U17425 (N_17425,N_16601,N_16430);
nand U17426 (N_17426,N_16382,N_16238);
xor U17427 (N_17427,N_16377,N_16558);
nor U17428 (N_17428,N_16748,N_16766);
nand U17429 (N_17429,N_16425,N_16893);
and U17430 (N_17430,N_16103,N_16970);
and U17431 (N_17431,N_16380,N_16690);
or U17432 (N_17432,N_16652,N_16735);
nor U17433 (N_17433,N_16712,N_16898);
xnor U17434 (N_17434,N_16805,N_16702);
xor U17435 (N_17435,N_16535,N_16343);
xnor U17436 (N_17436,N_16439,N_16812);
and U17437 (N_17437,N_16308,N_16115);
nor U17438 (N_17438,N_16233,N_16549);
and U17439 (N_17439,N_16912,N_16746);
xor U17440 (N_17440,N_16594,N_16843);
nor U17441 (N_17441,N_16833,N_16191);
xor U17442 (N_17442,N_16075,N_16634);
nor U17443 (N_17443,N_16846,N_16781);
xor U17444 (N_17444,N_16186,N_16719);
nor U17445 (N_17445,N_16839,N_16744);
or U17446 (N_17446,N_16984,N_16362);
xnor U17447 (N_17447,N_16567,N_16797);
and U17448 (N_17448,N_16365,N_16133);
nor U17449 (N_17449,N_16243,N_16355);
nor U17450 (N_17450,N_16356,N_16827);
xnor U17451 (N_17451,N_16715,N_16850);
nand U17452 (N_17452,N_16432,N_16440);
and U17453 (N_17453,N_16884,N_16907);
and U17454 (N_17454,N_16388,N_16855);
nor U17455 (N_17455,N_16336,N_16227);
xor U17456 (N_17456,N_16726,N_16779);
xnor U17457 (N_17457,N_16938,N_16258);
or U17458 (N_17458,N_16638,N_16498);
or U17459 (N_17459,N_16500,N_16836);
nor U17460 (N_17460,N_16899,N_16574);
and U17461 (N_17461,N_16314,N_16942);
nand U17462 (N_17462,N_16036,N_16842);
and U17463 (N_17463,N_16331,N_16466);
nor U17464 (N_17464,N_16268,N_16816);
nand U17465 (N_17465,N_16531,N_16819);
xnor U17466 (N_17466,N_16572,N_16953);
nand U17467 (N_17467,N_16845,N_16683);
nand U17468 (N_17468,N_16714,N_16251);
nand U17469 (N_17469,N_16048,N_16723);
or U17470 (N_17470,N_16577,N_16160);
xnor U17471 (N_17471,N_16457,N_16578);
nand U17472 (N_17472,N_16357,N_16927);
xnor U17473 (N_17473,N_16876,N_16221);
nand U17474 (N_17474,N_16564,N_16510);
and U17475 (N_17475,N_16108,N_16433);
nand U17476 (N_17476,N_16189,N_16429);
or U17477 (N_17477,N_16039,N_16270);
and U17478 (N_17478,N_16157,N_16142);
or U17479 (N_17479,N_16019,N_16537);
nor U17480 (N_17480,N_16618,N_16545);
nor U17481 (N_17481,N_16119,N_16257);
xor U17482 (N_17482,N_16813,N_16614);
nand U17483 (N_17483,N_16200,N_16513);
xnor U17484 (N_17484,N_16527,N_16342);
nor U17485 (N_17485,N_16569,N_16181);
or U17486 (N_17486,N_16378,N_16511);
nand U17487 (N_17487,N_16218,N_16949);
nor U17488 (N_17488,N_16460,N_16127);
xnor U17489 (N_17489,N_16216,N_16985);
nor U17490 (N_17490,N_16721,N_16023);
xor U17491 (N_17491,N_16959,N_16173);
or U17492 (N_17492,N_16386,N_16213);
xor U17493 (N_17493,N_16352,N_16788);
xnor U17494 (N_17494,N_16808,N_16273);
nand U17495 (N_17495,N_16037,N_16325);
and U17496 (N_17496,N_16472,N_16551);
nor U17497 (N_17497,N_16973,N_16063);
and U17498 (N_17498,N_16755,N_16729);
xnor U17499 (N_17499,N_16629,N_16056);
or U17500 (N_17500,N_16058,N_16227);
xnor U17501 (N_17501,N_16931,N_16305);
nor U17502 (N_17502,N_16668,N_16756);
xnor U17503 (N_17503,N_16299,N_16468);
nand U17504 (N_17504,N_16065,N_16410);
xnor U17505 (N_17505,N_16562,N_16131);
or U17506 (N_17506,N_16035,N_16106);
nor U17507 (N_17507,N_16933,N_16007);
nor U17508 (N_17508,N_16817,N_16291);
xnor U17509 (N_17509,N_16903,N_16464);
xnor U17510 (N_17510,N_16747,N_16645);
xor U17511 (N_17511,N_16382,N_16283);
nand U17512 (N_17512,N_16005,N_16789);
xnor U17513 (N_17513,N_16133,N_16950);
xor U17514 (N_17514,N_16873,N_16320);
nand U17515 (N_17515,N_16513,N_16460);
nand U17516 (N_17516,N_16116,N_16466);
nand U17517 (N_17517,N_16032,N_16304);
and U17518 (N_17518,N_16155,N_16910);
and U17519 (N_17519,N_16002,N_16485);
and U17520 (N_17520,N_16329,N_16251);
nor U17521 (N_17521,N_16588,N_16272);
nor U17522 (N_17522,N_16910,N_16924);
nor U17523 (N_17523,N_16832,N_16519);
xor U17524 (N_17524,N_16593,N_16039);
nor U17525 (N_17525,N_16994,N_16403);
nand U17526 (N_17526,N_16717,N_16212);
xor U17527 (N_17527,N_16368,N_16946);
nand U17528 (N_17528,N_16424,N_16480);
nor U17529 (N_17529,N_16952,N_16456);
or U17530 (N_17530,N_16823,N_16901);
nand U17531 (N_17531,N_16115,N_16471);
nand U17532 (N_17532,N_16299,N_16290);
or U17533 (N_17533,N_16635,N_16542);
or U17534 (N_17534,N_16740,N_16638);
or U17535 (N_17535,N_16085,N_16166);
or U17536 (N_17536,N_16059,N_16126);
nand U17537 (N_17537,N_16224,N_16700);
or U17538 (N_17538,N_16335,N_16710);
nand U17539 (N_17539,N_16381,N_16237);
nor U17540 (N_17540,N_16538,N_16664);
and U17541 (N_17541,N_16594,N_16799);
xnor U17542 (N_17542,N_16230,N_16290);
nor U17543 (N_17543,N_16445,N_16065);
nand U17544 (N_17544,N_16513,N_16554);
nor U17545 (N_17545,N_16271,N_16825);
nor U17546 (N_17546,N_16901,N_16581);
and U17547 (N_17547,N_16468,N_16664);
or U17548 (N_17548,N_16091,N_16283);
xor U17549 (N_17549,N_16104,N_16748);
or U17550 (N_17550,N_16885,N_16278);
nor U17551 (N_17551,N_16333,N_16860);
or U17552 (N_17552,N_16816,N_16825);
or U17553 (N_17553,N_16485,N_16567);
or U17554 (N_17554,N_16331,N_16947);
nor U17555 (N_17555,N_16970,N_16332);
nand U17556 (N_17556,N_16578,N_16916);
or U17557 (N_17557,N_16123,N_16724);
and U17558 (N_17558,N_16630,N_16974);
or U17559 (N_17559,N_16130,N_16709);
xor U17560 (N_17560,N_16990,N_16341);
and U17561 (N_17561,N_16596,N_16532);
xnor U17562 (N_17562,N_16066,N_16981);
nor U17563 (N_17563,N_16236,N_16282);
and U17564 (N_17564,N_16328,N_16413);
nor U17565 (N_17565,N_16854,N_16481);
and U17566 (N_17566,N_16813,N_16798);
nand U17567 (N_17567,N_16916,N_16752);
xor U17568 (N_17568,N_16466,N_16540);
or U17569 (N_17569,N_16056,N_16743);
nand U17570 (N_17570,N_16862,N_16167);
and U17571 (N_17571,N_16675,N_16633);
xnor U17572 (N_17572,N_16500,N_16784);
xor U17573 (N_17573,N_16607,N_16648);
nor U17574 (N_17574,N_16911,N_16482);
nor U17575 (N_17575,N_16390,N_16088);
xnor U17576 (N_17576,N_16040,N_16101);
or U17577 (N_17577,N_16005,N_16317);
or U17578 (N_17578,N_16210,N_16887);
nand U17579 (N_17579,N_16459,N_16480);
or U17580 (N_17580,N_16954,N_16512);
xor U17581 (N_17581,N_16031,N_16637);
nand U17582 (N_17582,N_16073,N_16132);
nor U17583 (N_17583,N_16663,N_16626);
nand U17584 (N_17584,N_16959,N_16310);
or U17585 (N_17585,N_16852,N_16744);
or U17586 (N_17586,N_16435,N_16107);
nand U17587 (N_17587,N_16616,N_16722);
nand U17588 (N_17588,N_16063,N_16078);
or U17589 (N_17589,N_16313,N_16941);
nor U17590 (N_17590,N_16465,N_16683);
and U17591 (N_17591,N_16458,N_16962);
xnor U17592 (N_17592,N_16818,N_16787);
nand U17593 (N_17593,N_16575,N_16620);
xor U17594 (N_17594,N_16458,N_16885);
and U17595 (N_17595,N_16690,N_16694);
nor U17596 (N_17596,N_16066,N_16591);
or U17597 (N_17597,N_16912,N_16774);
xor U17598 (N_17598,N_16517,N_16816);
nand U17599 (N_17599,N_16482,N_16541);
and U17600 (N_17600,N_16021,N_16602);
nand U17601 (N_17601,N_16278,N_16816);
nand U17602 (N_17602,N_16902,N_16575);
xnor U17603 (N_17603,N_16405,N_16547);
or U17604 (N_17604,N_16594,N_16730);
nor U17605 (N_17605,N_16130,N_16744);
nor U17606 (N_17606,N_16285,N_16672);
or U17607 (N_17607,N_16938,N_16011);
and U17608 (N_17608,N_16577,N_16626);
nand U17609 (N_17609,N_16042,N_16914);
or U17610 (N_17610,N_16586,N_16779);
nor U17611 (N_17611,N_16979,N_16006);
and U17612 (N_17612,N_16006,N_16517);
xnor U17613 (N_17613,N_16530,N_16186);
xnor U17614 (N_17614,N_16913,N_16759);
or U17615 (N_17615,N_16890,N_16876);
or U17616 (N_17616,N_16015,N_16754);
nor U17617 (N_17617,N_16602,N_16008);
nand U17618 (N_17618,N_16013,N_16897);
and U17619 (N_17619,N_16710,N_16803);
nor U17620 (N_17620,N_16897,N_16277);
and U17621 (N_17621,N_16941,N_16782);
nand U17622 (N_17622,N_16138,N_16463);
nor U17623 (N_17623,N_16523,N_16538);
xor U17624 (N_17624,N_16976,N_16147);
nand U17625 (N_17625,N_16100,N_16534);
xor U17626 (N_17626,N_16386,N_16438);
and U17627 (N_17627,N_16167,N_16056);
xor U17628 (N_17628,N_16167,N_16358);
and U17629 (N_17629,N_16892,N_16391);
or U17630 (N_17630,N_16735,N_16570);
nor U17631 (N_17631,N_16511,N_16088);
nor U17632 (N_17632,N_16500,N_16495);
or U17633 (N_17633,N_16306,N_16362);
xor U17634 (N_17634,N_16557,N_16566);
nand U17635 (N_17635,N_16231,N_16800);
or U17636 (N_17636,N_16131,N_16298);
xor U17637 (N_17637,N_16997,N_16974);
nor U17638 (N_17638,N_16824,N_16297);
xnor U17639 (N_17639,N_16598,N_16309);
and U17640 (N_17640,N_16389,N_16294);
xor U17641 (N_17641,N_16374,N_16277);
or U17642 (N_17642,N_16202,N_16688);
nor U17643 (N_17643,N_16357,N_16058);
nand U17644 (N_17644,N_16532,N_16062);
or U17645 (N_17645,N_16118,N_16197);
and U17646 (N_17646,N_16074,N_16532);
or U17647 (N_17647,N_16684,N_16164);
nand U17648 (N_17648,N_16404,N_16086);
xnor U17649 (N_17649,N_16411,N_16729);
and U17650 (N_17650,N_16918,N_16129);
or U17651 (N_17651,N_16239,N_16800);
or U17652 (N_17652,N_16703,N_16726);
nor U17653 (N_17653,N_16911,N_16593);
nand U17654 (N_17654,N_16147,N_16248);
nor U17655 (N_17655,N_16536,N_16786);
nor U17656 (N_17656,N_16860,N_16721);
nor U17657 (N_17657,N_16457,N_16530);
xnor U17658 (N_17658,N_16987,N_16827);
xor U17659 (N_17659,N_16180,N_16712);
nor U17660 (N_17660,N_16074,N_16925);
nor U17661 (N_17661,N_16429,N_16581);
nand U17662 (N_17662,N_16107,N_16208);
nor U17663 (N_17663,N_16976,N_16531);
and U17664 (N_17664,N_16367,N_16378);
and U17665 (N_17665,N_16538,N_16922);
nor U17666 (N_17666,N_16555,N_16092);
and U17667 (N_17667,N_16918,N_16254);
and U17668 (N_17668,N_16397,N_16291);
nand U17669 (N_17669,N_16797,N_16870);
nor U17670 (N_17670,N_16605,N_16902);
nand U17671 (N_17671,N_16439,N_16300);
xnor U17672 (N_17672,N_16271,N_16261);
nor U17673 (N_17673,N_16901,N_16930);
and U17674 (N_17674,N_16579,N_16008);
nor U17675 (N_17675,N_16078,N_16447);
and U17676 (N_17676,N_16502,N_16030);
or U17677 (N_17677,N_16735,N_16390);
nor U17678 (N_17678,N_16894,N_16734);
xnor U17679 (N_17679,N_16704,N_16114);
nor U17680 (N_17680,N_16000,N_16277);
nand U17681 (N_17681,N_16996,N_16993);
or U17682 (N_17682,N_16572,N_16756);
or U17683 (N_17683,N_16169,N_16257);
xor U17684 (N_17684,N_16358,N_16650);
nor U17685 (N_17685,N_16156,N_16654);
or U17686 (N_17686,N_16395,N_16157);
or U17687 (N_17687,N_16959,N_16744);
and U17688 (N_17688,N_16244,N_16255);
nor U17689 (N_17689,N_16364,N_16611);
nand U17690 (N_17690,N_16236,N_16259);
or U17691 (N_17691,N_16403,N_16002);
nand U17692 (N_17692,N_16065,N_16554);
nand U17693 (N_17693,N_16978,N_16282);
nor U17694 (N_17694,N_16883,N_16047);
nor U17695 (N_17695,N_16054,N_16550);
nand U17696 (N_17696,N_16505,N_16466);
nor U17697 (N_17697,N_16917,N_16250);
nor U17698 (N_17698,N_16134,N_16812);
nor U17699 (N_17699,N_16814,N_16608);
and U17700 (N_17700,N_16348,N_16430);
xor U17701 (N_17701,N_16540,N_16385);
and U17702 (N_17702,N_16713,N_16406);
or U17703 (N_17703,N_16630,N_16968);
nand U17704 (N_17704,N_16554,N_16113);
xor U17705 (N_17705,N_16455,N_16521);
nand U17706 (N_17706,N_16734,N_16996);
nand U17707 (N_17707,N_16399,N_16554);
nor U17708 (N_17708,N_16043,N_16862);
or U17709 (N_17709,N_16867,N_16973);
and U17710 (N_17710,N_16035,N_16579);
or U17711 (N_17711,N_16302,N_16555);
xnor U17712 (N_17712,N_16441,N_16411);
or U17713 (N_17713,N_16075,N_16033);
and U17714 (N_17714,N_16891,N_16658);
and U17715 (N_17715,N_16831,N_16925);
xnor U17716 (N_17716,N_16631,N_16340);
nor U17717 (N_17717,N_16498,N_16166);
nor U17718 (N_17718,N_16950,N_16714);
xnor U17719 (N_17719,N_16482,N_16969);
and U17720 (N_17720,N_16787,N_16257);
and U17721 (N_17721,N_16956,N_16284);
and U17722 (N_17722,N_16080,N_16574);
nand U17723 (N_17723,N_16092,N_16074);
xnor U17724 (N_17724,N_16048,N_16605);
xor U17725 (N_17725,N_16691,N_16328);
and U17726 (N_17726,N_16743,N_16077);
nand U17727 (N_17727,N_16558,N_16953);
or U17728 (N_17728,N_16245,N_16998);
nor U17729 (N_17729,N_16007,N_16307);
nor U17730 (N_17730,N_16470,N_16490);
nor U17731 (N_17731,N_16809,N_16425);
xnor U17732 (N_17732,N_16010,N_16732);
nor U17733 (N_17733,N_16161,N_16466);
xnor U17734 (N_17734,N_16699,N_16321);
and U17735 (N_17735,N_16494,N_16468);
and U17736 (N_17736,N_16250,N_16583);
or U17737 (N_17737,N_16654,N_16599);
or U17738 (N_17738,N_16864,N_16598);
or U17739 (N_17739,N_16933,N_16527);
or U17740 (N_17740,N_16538,N_16761);
and U17741 (N_17741,N_16470,N_16356);
or U17742 (N_17742,N_16918,N_16678);
nand U17743 (N_17743,N_16387,N_16187);
or U17744 (N_17744,N_16201,N_16151);
and U17745 (N_17745,N_16874,N_16197);
and U17746 (N_17746,N_16565,N_16617);
xnor U17747 (N_17747,N_16885,N_16954);
xor U17748 (N_17748,N_16705,N_16868);
or U17749 (N_17749,N_16517,N_16693);
nor U17750 (N_17750,N_16891,N_16494);
xnor U17751 (N_17751,N_16244,N_16230);
xor U17752 (N_17752,N_16346,N_16512);
and U17753 (N_17753,N_16159,N_16336);
nand U17754 (N_17754,N_16143,N_16380);
or U17755 (N_17755,N_16440,N_16551);
and U17756 (N_17756,N_16456,N_16162);
nand U17757 (N_17757,N_16139,N_16591);
or U17758 (N_17758,N_16196,N_16086);
or U17759 (N_17759,N_16282,N_16513);
and U17760 (N_17760,N_16551,N_16309);
or U17761 (N_17761,N_16899,N_16960);
or U17762 (N_17762,N_16155,N_16024);
or U17763 (N_17763,N_16246,N_16741);
nor U17764 (N_17764,N_16917,N_16334);
or U17765 (N_17765,N_16732,N_16522);
nand U17766 (N_17766,N_16573,N_16353);
or U17767 (N_17767,N_16548,N_16364);
or U17768 (N_17768,N_16298,N_16555);
nor U17769 (N_17769,N_16904,N_16191);
nor U17770 (N_17770,N_16471,N_16145);
and U17771 (N_17771,N_16377,N_16272);
and U17772 (N_17772,N_16385,N_16109);
nor U17773 (N_17773,N_16351,N_16040);
nor U17774 (N_17774,N_16625,N_16146);
nand U17775 (N_17775,N_16426,N_16740);
nor U17776 (N_17776,N_16287,N_16256);
nand U17777 (N_17777,N_16659,N_16507);
nor U17778 (N_17778,N_16048,N_16600);
or U17779 (N_17779,N_16383,N_16488);
xnor U17780 (N_17780,N_16964,N_16238);
and U17781 (N_17781,N_16896,N_16642);
nor U17782 (N_17782,N_16156,N_16933);
nor U17783 (N_17783,N_16141,N_16313);
or U17784 (N_17784,N_16874,N_16809);
and U17785 (N_17785,N_16950,N_16946);
xor U17786 (N_17786,N_16647,N_16089);
or U17787 (N_17787,N_16526,N_16826);
or U17788 (N_17788,N_16210,N_16035);
and U17789 (N_17789,N_16553,N_16252);
nor U17790 (N_17790,N_16040,N_16707);
or U17791 (N_17791,N_16452,N_16762);
nand U17792 (N_17792,N_16444,N_16024);
nor U17793 (N_17793,N_16483,N_16579);
xor U17794 (N_17794,N_16479,N_16252);
xnor U17795 (N_17795,N_16121,N_16125);
xor U17796 (N_17796,N_16640,N_16903);
xor U17797 (N_17797,N_16701,N_16821);
xnor U17798 (N_17798,N_16229,N_16014);
nor U17799 (N_17799,N_16027,N_16210);
or U17800 (N_17800,N_16994,N_16591);
nand U17801 (N_17801,N_16878,N_16414);
nor U17802 (N_17802,N_16038,N_16291);
xnor U17803 (N_17803,N_16473,N_16694);
nor U17804 (N_17804,N_16919,N_16926);
xnor U17805 (N_17805,N_16802,N_16155);
or U17806 (N_17806,N_16066,N_16623);
or U17807 (N_17807,N_16339,N_16179);
nor U17808 (N_17808,N_16716,N_16032);
nand U17809 (N_17809,N_16027,N_16003);
and U17810 (N_17810,N_16146,N_16518);
and U17811 (N_17811,N_16407,N_16570);
nor U17812 (N_17812,N_16612,N_16732);
and U17813 (N_17813,N_16890,N_16746);
or U17814 (N_17814,N_16058,N_16383);
nand U17815 (N_17815,N_16040,N_16895);
xnor U17816 (N_17816,N_16153,N_16518);
nor U17817 (N_17817,N_16055,N_16584);
and U17818 (N_17818,N_16957,N_16915);
or U17819 (N_17819,N_16810,N_16923);
nand U17820 (N_17820,N_16603,N_16555);
and U17821 (N_17821,N_16202,N_16715);
or U17822 (N_17822,N_16939,N_16917);
nor U17823 (N_17823,N_16986,N_16503);
nand U17824 (N_17824,N_16403,N_16877);
xnor U17825 (N_17825,N_16368,N_16628);
xnor U17826 (N_17826,N_16249,N_16576);
nor U17827 (N_17827,N_16843,N_16466);
xnor U17828 (N_17828,N_16548,N_16708);
and U17829 (N_17829,N_16203,N_16535);
and U17830 (N_17830,N_16983,N_16602);
nand U17831 (N_17831,N_16472,N_16522);
or U17832 (N_17832,N_16542,N_16660);
nand U17833 (N_17833,N_16386,N_16655);
or U17834 (N_17834,N_16088,N_16059);
xor U17835 (N_17835,N_16237,N_16030);
or U17836 (N_17836,N_16548,N_16192);
and U17837 (N_17837,N_16544,N_16706);
or U17838 (N_17838,N_16110,N_16919);
or U17839 (N_17839,N_16850,N_16948);
nand U17840 (N_17840,N_16721,N_16225);
or U17841 (N_17841,N_16395,N_16657);
nand U17842 (N_17842,N_16690,N_16807);
or U17843 (N_17843,N_16958,N_16062);
nor U17844 (N_17844,N_16975,N_16065);
xor U17845 (N_17845,N_16868,N_16890);
xnor U17846 (N_17846,N_16805,N_16041);
xnor U17847 (N_17847,N_16752,N_16445);
xnor U17848 (N_17848,N_16118,N_16969);
and U17849 (N_17849,N_16754,N_16407);
or U17850 (N_17850,N_16708,N_16019);
and U17851 (N_17851,N_16025,N_16468);
or U17852 (N_17852,N_16090,N_16590);
nor U17853 (N_17853,N_16668,N_16573);
and U17854 (N_17854,N_16233,N_16186);
xnor U17855 (N_17855,N_16958,N_16291);
nor U17856 (N_17856,N_16053,N_16891);
nor U17857 (N_17857,N_16811,N_16309);
and U17858 (N_17858,N_16039,N_16451);
nor U17859 (N_17859,N_16318,N_16101);
nor U17860 (N_17860,N_16318,N_16666);
nor U17861 (N_17861,N_16767,N_16879);
or U17862 (N_17862,N_16369,N_16221);
and U17863 (N_17863,N_16699,N_16950);
and U17864 (N_17864,N_16995,N_16331);
xnor U17865 (N_17865,N_16936,N_16810);
and U17866 (N_17866,N_16355,N_16023);
nor U17867 (N_17867,N_16379,N_16001);
or U17868 (N_17868,N_16740,N_16820);
xnor U17869 (N_17869,N_16003,N_16586);
nand U17870 (N_17870,N_16961,N_16271);
xnor U17871 (N_17871,N_16766,N_16757);
xnor U17872 (N_17872,N_16499,N_16916);
nand U17873 (N_17873,N_16116,N_16898);
nor U17874 (N_17874,N_16278,N_16920);
xnor U17875 (N_17875,N_16155,N_16385);
xor U17876 (N_17876,N_16989,N_16437);
and U17877 (N_17877,N_16192,N_16817);
nand U17878 (N_17878,N_16412,N_16940);
or U17879 (N_17879,N_16687,N_16032);
and U17880 (N_17880,N_16348,N_16267);
nand U17881 (N_17881,N_16943,N_16124);
nor U17882 (N_17882,N_16067,N_16875);
or U17883 (N_17883,N_16226,N_16775);
nand U17884 (N_17884,N_16715,N_16487);
nand U17885 (N_17885,N_16651,N_16502);
nand U17886 (N_17886,N_16151,N_16824);
and U17887 (N_17887,N_16580,N_16838);
or U17888 (N_17888,N_16265,N_16966);
and U17889 (N_17889,N_16390,N_16826);
or U17890 (N_17890,N_16845,N_16529);
or U17891 (N_17891,N_16854,N_16501);
xnor U17892 (N_17892,N_16471,N_16402);
nand U17893 (N_17893,N_16213,N_16011);
nand U17894 (N_17894,N_16889,N_16600);
or U17895 (N_17895,N_16799,N_16077);
or U17896 (N_17896,N_16695,N_16311);
or U17897 (N_17897,N_16847,N_16187);
or U17898 (N_17898,N_16389,N_16359);
nor U17899 (N_17899,N_16540,N_16310);
xnor U17900 (N_17900,N_16671,N_16899);
nor U17901 (N_17901,N_16412,N_16320);
nor U17902 (N_17902,N_16798,N_16151);
xor U17903 (N_17903,N_16027,N_16149);
xnor U17904 (N_17904,N_16178,N_16695);
nor U17905 (N_17905,N_16757,N_16553);
nand U17906 (N_17906,N_16108,N_16546);
nor U17907 (N_17907,N_16038,N_16938);
and U17908 (N_17908,N_16810,N_16507);
xor U17909 (N_17909,N_16211,N_16183);
nor U17910 (N_17910,N_16359,N_16421);
or U17911 (N_17911,N_16464,N_16954);
and U17912 (N_17912,N_16489,N_16570);
xnor U17913 (N_17913,N_16175,N_16705);
xnor U17914 (N_17914,N_16335,N_16581);
and U17915 (N_17915,N_16102,N_16127);
nor U17916 (N_17916,N_16444,N_16837);
nor U17917 (N_17917,N_16365,N_16718);
nor U17918 (N_17918,N_16851,N_16818);
xor U17919 (N_17919,N_16150,N_16970);
nor U17920 (N_17920,N_16160,N_16400);
nand U17921 (N_17921,N_16616,N_16555);
nor U17922 (N_17922,N_16997,N_16156);
nand U17923 (N_17923,N_16494,N_16385);
xor U17924 (N_17924,N_16839,N_16651);
nand U17925 (N_17925,N_16930,N_16259);
or U17926 (N_17926,N_16266,N_16881);
nor U17927 (N_17927,N_16131,N_16600);
and U17928 (N_17928,N_16735,N_16747);
nand U17929 (N_17929,N_16768,N_16283);
xor U17930 (N_17930,N_16057,N_16107);
nand U17931 (N_17931,N_16508,N_16011);
nor U17932 (N_17932,N_16077,N_16584);
nor U17933 (N_17933,N_16796,N_16990);
and U17934 (N_17934,N_16895,N_16564);
nor U17935 (N_17935,N_16509,N_16598);
nand U17936 (N_17936,N_16845,N_16983);
nand U17937 (N_17937,N_16173,N_16060);
or U17938 (N_17938,N_16859,N_16710);
xnor U17939 (N_17939,N_16840,N_16172);
and U17940 (N_17940,N_16250,N_16475);
nor U17941 (N_17941,N_16604,N_16736);
nand U17942 (N_17942,N_16759,N_16008);
nand U17943 (N_17943,N_16671,N_16493);
nand U17944 (N_17944,N_16022,N_16722);
nor U17945 (N_17945,N_16128,N_16480);
nand U17946 (N_17946,N_16417,N_16970);
nor U17947 (N_17947,N_16127,N_16753);
nand U17948 (N_17948,N_16521,N_16358);
xor U17949 (N_17949,N_16448,N_16866);
nor U17950 (N_17950,N_16182,N_16311);
nand U17951 (N_17951,N_16333,N_16793);
xor U17952 (N_17952,N_16157,N_16425);
nand U17953 (N_17953,N_16581,N_16940);
nand U17954 (N_17954,N_16489,N_16969);
nand U17955 (N_17955,N_16086,N_16808);
xnor U17956 (N_17956,N_16141,N_16772);
nor U17957 (N_17957,N_16954,N_16341);
nor U17958 (N_17958,N_16015,N_16225);
nor U17959 (N_17959,N_16865,N_16566);
nand U17960 (N_17960,N_16829,N_16728);
nor U17961 (N_17961,N_16918,N_16082);
xor U17962 (N_17962,N_16909,N_16202);
or U17963 (N_17963,N_16833,N_16623);
xnor U17964 (N_17964,N_16168,N_16050);
nand U17965 (N_17965,N_16624,N_16564);
nand U17966 (N_17966,N_16314,N_16430);
nand U17967 (N_17967,N_16339,N_16412);
nand U17968 (N_17968,N_16569,N_16089);
or U17969 (N_17969,N_16132,N_16763);
and U17970 (N_17970,N_16910,N_16057);
or U17971 (N_17971,N_16418,N_16356);
or U17972 (N_17972,N_16003,N_16711);
and U17973 (N_17973,N_16400,N_16488);
and U17974 (N_17974,N_16211,N_16699);
nand U17975 (N_17975,N_16417,N_16029);
nand U17976 (N_17976,N_16782,N_16900);
and U17977 (N_17977,N_16141,N_16888);
xnor U17978 (N_17978,N_16919,N_16048);
nand U17979 (N_17979,N_16255,N_16807);
or U17980 (N_17980,N_16418,N_16696);
nand U17981 (N_17981,N_16759,N_16806);
xnor U17982 (N_17982,N_16952,N_16750);
xnor U17983 (N_17983,N_16833,N_16632);
nand U17984 (N_17984,N_16782,N_16827);
nand U17985 (N_17985,N_16824,N_16000);
xnor U17986 (N_17986,N_16767,N_16888);
nor U17987 (N_17987,N_16694,N_16515);
or U17988 (N_17988,N_16423,N_16398);
or U17989 (N_17989,N_16564,N_16820);
and U17990 (N_17990,N_16366,N_16882);
nand U17991 (N_17991,N_16346,N_16059);
nand U17992 (N_17992,N_16116,N_16336);
and U17993 (N_17993,N_16665,N_16985);
nand U17994 (N_17994,N_16869,N_16874);
or U17995 (N_17995,N_16729,N_16920);
nor U17996 (N_17996,N_16714,N_16759);
nand U17997 (N_17997,N_16312,N_16116);
or U17998 (N_17998,N_16481,N_16363);
and U17999 (N_17999,N_16321,N_16722);
nor U18000 (N_18000,N_17180,N_17081);
xnor U18001 (N_18001,N_17888,N_17433);
nor U18002 (N_18002,N_17969,N_17718);
or U18003 (N_18003,N_17508,N_17754);
and U18004 (N_18004,N_17052,N_17287);
xor U18005 (N_18005,N_17842,N_17610);
nand U18006 (N_18006,N_17203,N_17424);
or U18007 (N_18007,N_17390,N_17809);
or U18008 (N_18008,N_17353,N_17825);
and U18009 (N_18009,N_17705,N_17944);
or U18010 (N_18010,N_17557,N_17444);
nor U18011 (N_18011,N_17979,N_17876);
xor U18012 (N_18012,N_17284,N_17331);
nand U18013 (N_18013,N_17847,N_17161);
nor U18014 (N_18014,N_17495,N_17430);
or U18015 (N_18015,N_17870,N_17271);
or U18016 (N_18016,N_17612,N_17669);
nand U18017 (N_18017,N_17733,N_17563);
xnor U18018 (N_18018,N_17596,N_17348);
nand U18019 (N_18019,N_17558,N_17550);
or U18020 (N_18020,N_17282,N_17060);
nor U18021 (N_18021,N_17240,N_17651);
and U18022 (N_18022,N_17208,N_17780);
nor U18023 (N_18023,N_17379,N_17073);
or U18024 (N_18024,N_17176,N_17694);
nand U18025 (N_18025,N_17013,N_17128);
or U18026 (N_18026,N_17385,N_17947);
and U18027 (N_18027,N_17113,N_17542);
xor U18028 (N_18028,N_17742,N_17318);
nor U18029 (N_18029,N_17878,N_17711);
xor U18030 (N_18030,N_17023,N_17342);
nor U18031 (N_18031,N_17791,N_17359);
nand U18032 (N_18032,N_17998,N_17577);
and U18033 (N_18033,N_17639,N_17633);
nand U18034 (N_18034,N_17374,N_17098);
nor U18035 (N_18035,N_17327,N_17887);
nor U18036 (N_18036,N_17166,N_17048);
xor U18037 (N_18037,N_17786,N_17659);
and U18038 (N_18038,N_17003,N_17991);
or U18039 (N_18039,N_17478,N_17360);
or U18040 (N_18040,N_17107,N_17506);
nor U18041 (N_18041,N_17942,N_17518);
nor U18042 (N_18042,N_17986,N_17362);
nor U18043 (N_18043,N_17093,N_17338);
or U18044 (N_18044,N_17623,N_17578);
xnor U18045 (N_18045,N_17441,N_17635);
nand U18046 (N_18046,N_17871,N_17761);
xnor U18047 (N_18047,N_17447,N_17598);
xor U18048 (N_18048,N_17975,N_17957);
nand U18049 (N_18049,N_17469,N_17946);
or U18050 (N_18050,N_17905,N_17728);
and U18051 (N_18051,N_17296,N_17425);
or U18052 (N_18052,N_17426,N_17212);
or U18053 (N_18053,N_17658,N_17350);
and U18054 (N_18054,N_17756,N_17798);
and U18055 (N_18055,N_17361,N_17152);
xor U18056 (N_18056,N_17094,N_17706);
nand U18057 (N_18057,N_17608,N_17216);
nor U18058 (N_18058,N_17923,N_17267);
and U18059 (N_18059,N_17459,N_17178);
nand U18060 (N_18060,N_17914,N_17984);
xor U18061 (N_18061,N_17642,N_17647);
xor U18062 (N_18062,N_17953,N_17421);
nand U18063 (N_18063,N_17885,N_17020);
nor U18064 (N_18064,N_17845,N_17268);
nand U18065 (N_18065,N_17813,N_17238);
nor U18066 (N_18066,N_17988,N_17033);
nand U18067 (N_18067,N_17653,N_17482);
and U18068 (N_18068,N_17521,N_17964);
xnor U18069 (N_18069,N_17114,N_17265);
or U18070 (N_18070,N_17803,N_17209);
nor U18071 (N_18071,N_17131,N_17129);
or U18072 (N_18072,N_17865,N_17170);
nand U18073 (N_18073,N_17740,N_17371);
xor U18074 (N_18074,N_17739,N_17965);
or U18075 (N_18075,N_17922,N_17758);
xor U18076 (N_18076,N_17648,N_17179);
xnor U18077 (N_18077,N_17355,N_17788);
nor U18078 (N_18078,N_17677,N_17399);
nand U18079 (N_18079,N_17115,N_17898);
nand U18080 (N_18080,N_17784,N_17637);
nor U18081 (N_18081,N_17283,N_17043);
and U18082 (N_18082,N_17005,N_17262);
nand U18083 (N_18083,N_17218,N_17732);
xnor U18084 (N_18084,N_17859,N_17483);
nand U18085 (N_18085,N_17785,N_17276);
nor U18086 (N_18086,N_17402,N_17802);
nor U18087 (N_18087,N_17047,N_17833);
or U18088 (N_18088,N_17621,N_17800);
xnor U18089 (N_18089,N_17717,N_17294);
nor U18090 (N_18090,N_17886,N_17310);
or U18091 (N_18091,N_17032,N_17877);
nor U18092 (N_18092,N_17553,N_17416);
or U18093 (N_18093,N_17997,N_17008);
nand U18094 (N_18094,N_17231,N_17151);
nor U18095 (N_18095,N_17630,N_17691);
nand U18096 (N_18096,N_17470,N_17099);
xnor U18097 (N_18097,N_17417,N_17408);
nor U18098 (N_18098,N_17415,N_17852);
nor U18099 (N_18099,N_17229,N_17773);
nand U18100 (N_18100,N_17239,N_17146);
nor U18101 (N_18101,N_17450,N_17202);
xnor U18102 (N_18102,N_17423,N_17243);
xor U18103 (N_18103,N_17219,N_17215);
nand U18104 (N_18104,N_17201,N_17256);
nand U18105 (N_18105,N_17745,N_17794);
or U18106 (N_18106,N_17150,N_17461);
nand U18107 (N_18107,N_17588,N_17681);
xor U18108 (N_18108,N_17321,N_17737);
and U18109 (N_18109,N_17398,N_17792);
xor U18110 (N_18110,N_17400,N_17344);
and U18111 (N_18111,N_17382,N_17827);
nor U18112 (N_18112,N_17925,N_17729);
nor U18113 (N_18113,N_17144,N_17473);
nand U18114 (N_18114,N_17041,N_17959);
and U18115 (N_18115,N_17292,N_17096);
and U18116 (N_18116,N_17304,N_17451);
or U18117 (N_18117,N_17019,N_17090);
nor U18118 (N_18118,N_17396,N_17365);
or U18119 (N_18119,N_17184,N_17832);
nand U18120 (N_18120,N_17725,N_17332);
nor U18121 (N_18121,N_17091,N_17194);
nor U18122 (N_18122,N_17100,N_17299);
xor U18123 (N_18123,N_17274,N_17667);
and U18124 (N_18124,N_17641,N_17738);
nand U18125 (N_18125,N_17743,N_17475);
nand U18126 (N_18126,N_17222,N_17199);
nand U18127 (N_18127,N_17968,N_17934);
nand U18128 (N_18128,N_17657,N_17987);
nor U18129 (N_18129,N_17936,N_17586);
xnor U18130 (N_18130,N_17118,N_17607);
xor U18131 (N_18131,N_17797,N_17941);
nor U18132 (N_18132,N_17901,N_17103);
nor U18133 (N_18133,N_17490,N_17566);
nand U18134 (N_18134,N_17962,N_17600);
nand U18135 (N_18135,N_17252,N_17367);
and U18136 (N_18136,N_17322,N_17235);
and U18137 (N_18137,N_17030,N_17401);
and U18138 (N_18138,N_17722,N_17333);
xor U18139 (N_18139,N_17339,N_17029);
or U18140 (N_18140,N_17909,N_17080);
and U18141 (N_18141,N_17237,N_17526);
or U18142 (N_18142,N_17714,N_17241);
or U18143 (N_18143,N_17655,N_17049);
xnor U18144 (N_18144,N_17255,N_17077);
or U18145 (N_18145,N_17719,N_17516);
xnor U18146 (N_18146,N_17109,N_17171);
or U18147 (N_18147,N_17851,N_17807);
xor U18148 (N_18148,N_17846,N_17445);
or U18149 (N_18149,N_17801,N_17661);
and U18150 (N_18150,N_17242,N_17016);
and U18151 (N_18151,N_17038,N_17844);
xnor U18152 (N_18152,N_17181,N_17306);
nor U18153 (N_18153,N_17311,N_17042);
or U18154 (N_18154,N_17198,N_17308);
xor U18155 (N_18155,N_17232,N_17976);
xnor U18156 (N_18156,N_17145,N_17892);
and U18157 (N_18157,N_17177,N_17187);
nor U18158 (N_18158,N_17875,N_17864);
nand U18159 (N_18159,N_17319,N_17487);
or U18160 (N_18160,N_17514,N_17026);
xor U18161 (N_18161,N_17907,N_17337);
xor U18162 (N_18162,N_17768,N_17406);
nor U18163 (N_18163,N_17760,N_17996);
nor U18164 (N_18164,N_17403,N_17329);
nor U18165 (N_18165,N_17254,N_17443);
xnor U18166 (N_18166,N_17731,N_17662);
and U18167 (N_18167,N_17629,N_17244);
xnor U18168 (N_18168,N_17498,N_17142);
or U18169 (N_18169,N_17650,N_17505);
and U18170 (N_18170,N_17480,N_17716);
xor U18171 (N_18171,N_17536,N_17465);
xor U18172 (N_18172,N_17228,N_17172);
xor U18173 (N_18173,N_17519,N_17771);
and U18174 (N_18174,N_17044,N_17468);
nand U18175 (N_18175,N_17313,N_17420);
xnor U18176 (N_18176,N_17804,N_17446);
and U18177 (N_18177,N_17057,N_17250);
and U18178 (N_18178,N_17897,N_17952);
nor U18179 (N_18179,N_17314,N_17105);
and U18180 (N_18180,N_17200,N_17948);
and U18181 (N_18181,N_17169,N_17162);
nor U18182 (N_18182,N_17701,N_17766);
and U18183 (N_18183,N_17741,N_17912);
nor U18184 (N_18184,N_17812,N_17393);
nor U18185 (N_18185,N_17675,N_17700);
nand U18186 (N_18186,N_17497,N_17626);
and U18187 (N_18187,N_17850,N_17966);
xor U18188 (N_18188,N_17568,N_17974);
nand U18189 (N_18189,N_17665,N_17460);
and U18190 (N_18190,N_17839,N_17205);
nand U18191 (N_18191,N_17175,N_17059);
xor U18192 (N_18192,N_17015,N_17230);
nand U18193 (N_18193,N_17702,N_17084);
nand U18194 (N_18194,N_17206,N_17695);
xnor U18195 (N_18195,N_17672,N_17358);
nor U18196 (N_18196,N_17001,N_17493);
nand U18197 (N_18197,N_17474,N_17715);
nor U18198 (N_18198,N_17918,N_17410);
or U18199 (N_18199,N_17924,N_17624);
nand U18200 (N_18200,N_17606,N_17106);
or U18201 (N_18201,N_17853,N_17652);
and U18202 (N_18202,N_17576,N_17945);
xor U18203 (N_18203,N_17346,N_17189);
nand U18204 (N_18204,N_17890,N_17491);
xnor U18205 (N_18205,N_17328,N_17046);
or U18206 (N_18206,N_17050,N_17572);
nand U18207 (N_18207,N_17755,N_17915);
nand U18208 (N_18208,N_17213,N_17245);
xnor U18209 (N_18209,N_17605,N_17438);
nand U18210 (N_18210,N_17211,N_17375);
and U18211 (N_18211,N_17273,N_17783);
or U18212 (N_18212,N_17156,N_17591);
and U18213 (N_18213,N_17867,N_17806);
nor U18214 (N_18214,N_17025,N_17971);
and U18215 (N_18215,N_17838,N_17502);
or U18216 (N_18216,N_17000,N_17823);
nand U18217 (N_18217,N_17625,N_17779);
xnor U18218 (N_18218,N_17489,N_17031);
xnor U18219 (N_18219,N_17501,N_17906);
nand U18220 (N_18220,N_17594,N_17949);
or U18221 (N_18221,N_17039,N_17009);
and U18222 (N_18222,N_17072,N_17618);
nand U18223 (N_18223,N_17749,N_17727);
nor U18224 (N_18224,N_17532,N_17334);
or U18225 (N_18225,N_17893,N_17427);
nand U18226 (N_18226,N_17500,N_17253);
or U18227 (N_18227,N_17186,N_17158);
or U18228 (N_18228,N_17076,N_17750);
nor U18229 (N_18229,N_17615,N_17108);
nor U18230 (N_18230,N_17117,N_17614);
or U18231 (N_18231,N_17210,N_17682);
nand U18232 (N_18232,N_17824,N_17432);
xor U18233 (N_18233,N_17574,N_17492);
nor U18234 (N_18234,N_17581,N_17448);
nor U18235 (N_18235,N_17165,N_17139);
nor U18236 (N_18236,N_17699,N_17275);
nand U18237 (N_18237,N_17082,N_17869);
nor U18238 (N_18238,N_17884,N_17819);
nor U18239 (N_18239,N_17775,N_17751);
and U18240 (N_18240,N_17278,N_17926);
nand U18241 (N_18241,N_17730,N_17195);
nand U18242 (N_18242,N_17554,N_17654);
xnor U18243 (N_18243,N_17599,N_17370);
nand U18244 (N_18244,N_17649,N_17196);
nand U18245 (N_18245,N_17354,N_17685);
nand U18246 (N_18246,N_17762,N_17668);
or U18247 (N_18247,N_17343,N_17481);
xnor U18248 (N_18248,N_17836,N_17961);
nand U18249 (N_18249,N_17056,N_17110);
and U18250 (N_18250,N_17386,N_17297);
and U18251 (N_18251,N_17676,N_17330);
or U18252 (N_18252,N_17437,N_17787);
or U18253 (N_18253,N_17562,N_17479);
nor U18254 (N_18254,N_17028,N_17351);
nand U18255 (N_18255,N_17548,N_17613);
and U18256 (N_18256,N_17167,N_17021);
xor U18257 (N_18257,N_17970,N_17656);
or U18258 (N_18258,N_17088,N_17690);
and U18259 (N_18259,N_17678,N_17340);
nand U18260 (N_18260,N_17266,N_17644);
xor U18261 (N_18261,N_17397,N_17193);
xor U18262 (N_18262,N_17246,N_17494);
nand U18263 (N_18263,N_17006,N_17617);
nand U18264 (N_18264,N_17551,N_17584);
xor U18265 (N_18265,N_17204,N_17312);
nand U18266 (N_18266,N_17281,N_17272);
and U18267 (N_18267,N_17593,N_17759);
nor U18268 (N_18268,N_17055,N_17191);
nor U18269 (N_18269,N_17795,N_17325);
or U18270 (N_18270,N_17589,N_17973);
or U18271 (N_18271,N_17620,N_17697);
and U18272 (N_18272,N_17980,N_17774);
and U18273 (N_18273,N_17636,N_17781);
or U18274 (N_18274,N_17776,N_17680);
or U18275 (N_18275,N_17127,N_17356);
and U18276 (N_18276,N_17570,N_17111);
and U18277 (N_18277,N_17429,N_17036);
nor U18278 (N_18278,N_17157,N_17018);
and U18279 (N_18279,N_17561,N_17102);
nor U18280 (N_18280,N_17830,N_17069);
nand U18281 (N_18281,N_17671,N_17686);
and U18282 (N_18282,N_17580,N_17054);
and U18283 (N_18283,N_17486,N_17476);
xnor U18284 (N_18284,N_17814,N_17249);
and U18285 (N_18285,N_17264,N_17790);
nor U18286 (N_18286,N_17645,N_17627);
xor U18287 (N_18287,N_17866,N_17748);
and U18288 (N_18288,N_17937,N_17067);
nor U18289 (N_18289,N_17684,N_17539);
and U18290 (N_18290,N_17512,N_17455);
xnor U18291 (N_18291,N_17251,N_17065);
and U18292 (N_18292,N_17225,N_17873);
and U18293 (N_18293,N_17323,N_17511);
or U18294 (N_18294,N_17646,N_17543);
xnor U18295 (N_18295,N_17035,N_17247);
and U18296 (N_18296,N_17289,N_17525);
or U18297 (N_18297,N_17902,N_17805);
nor U18298 (N_18298,N_17510,N_17917);
nand U18299 (N_18299,N_17452,N_17528);
nor U18300 (N_18300,N_17467,N_17777);
or U18301 (N_18301,N_17995,N_17457);
xnor U18302 (N_18302,N_17515,N_17520);
or U18303 (N_18303,N_17002,N_17037);
nand U18304 (N_18304,N_17395,N_17141);
xor U18305 (N_18305,N_17236,N_17933);
or U18306 (N_18306,N_17928,N_17585);
nor U18307 (N_18307,N_17704,N_17155);
nand U18308 (N_18308,N_17992,N_17810);
or U18309 (N_18309,N_17471,N_17364);
or U18310 (N_18310,N_17604,N_17341);
and U18311 (N_18311,N_17384,N_17595);
nand U18312 (N_18312,N_17619,N_17083);
nand U18313 (N_18313,N_17960,N_17290);
xor U18314 (N_18314,N_17197,N_17855);
xnor U18315 (N_18315,N_17376,N_17135);
and U18316 (N_18316,N_17703,N_17575);
nor U18317 (N_18317,N_17439,N_17414);
and U18318 (N_18318,N_17582,N_17927);
nor U18319 (N_18319,N_17349,N_17164);
xnor U18320 (N_18320,N_17010,N_17214);
or U18321 (N_18321,N_17453,N_17860);
xor U18322 (N_18322,N_17380,N_17808);
nand U18323 (N_18323,N_17990,N_17541);
xnor U18324 (N_18324,N_17903,N_17316);
and U18325 (N_18325,N_17609,N_17880);
or U18326 (N_18326,N_17772,N_17303);
nand U18327 (N_18327,N_17079,N_17413);
or U18328 (N_18328,N_17434,N_17537);
or U18329 (N_18329,N_17387,N_17422);
xnor U18330 (N_18330,N_17440,N_17357);
and U18331 (N_18331,N_17565,N_17829);
or U18332 (N_18332,N_17078,N_17889);
and U18333 (N_18333,N_17874,N_17064);
xor U18334 (N_18334,N_17721,N_17981);
nor U18335 (N_18335,N_17217,N_17280);
xnor U18336 (N_18336,N_17336,N_17027);
xnor U18337 (N_18337,N_17908,N_17854);
nand U18338 (N_18338,N_17631,N_17564);
or U18339 (N_18339,N_17590,N_17985);
nor U18340 (N_18340,N_17752,N_17963);
or U18341 (N_18341,N_17305,N_17567);
nand U18342 (N_18342,N_17435,N_17696);
and U18343 (N_18343,N_17904,N_17683);
or U18344 (N_18344,N_17378,N_17999);
and U18345 (N_18345,N_17726,N_17286);
nor U18346 (N_18346,N_17882,N_17883);
xnor U18347 (N_18347,N_17221,N_17309);
nor U18348 (N_18348,N_17993,N_17017);
nor U18349 (N_18349,N_17956,N_17517);
or U18350 (N_18350,N_17503,N_17938);
or U18351 (N_18351,N_17368,N_17140);
or U18352 (N_18352,N_17404,N_17921);
nand U18353 (N_18353,N_17012,N_17087);
or U18354 (N_18354,N_17789,N_17134);
and U18355 (N_18355,N_17449,N_17664);
nand U18356 (N_18356,N_17817,N_17513);
and U18357 (N_18357,N_17307,N_17587);
xor U18358 (N_18358,N_17125,N_17720);
or U18359 (N_18359,N_17377,N_17916);
and U18360 (N_18360,N_17763,N_17552);
nand U18361 (N_18361,N_17724,N_17837);
nand U18362 (N_18362,N_17063,N_17687);
or U18363 (N_18363,N_17463,N_17062);
or U18364 (N_18364,N_17534,N_17747);
and U18365 (N_18365,N_17821,N_17939);
and U18366 (N_18366,N_17549,N_17616);
and U18367 (N_18367,N_17147,N_17507);
nand U18368 (N_18368,N_17220,N_17138);
nor U18369 (N_18369,N_17058,N_17392);
and U18370 (N_18370,N_17116,N_17394);
and U18371 (N_18371,N_17345,N_17547);
nor U18372 (N_18372,N_17472,N_17769);
or U18373 (N_18373,N_17840,N_17061);
nor U18374 (N_18374,N_17014,N_17488);
and U18375 (N_18375,N_17227,N_17920);
nand U18376 (N_18376,N_17736,N_17185);
xor U18377 (N_18377,N_17931,N_17383);
or U18378 (N_18378,N_17796,N_17955);
and U18379 (N_18379,N_17101,N_17688);
nand U18380 (N_18380,N_17982,N_17632);
and U18381 (N_18381,N_17381,N_17746);
and U18382 (N_18382,N_17291,N_17143);
and U18383 (N_18383,N_17753,N_17089);
or U18384 (N_18384,N_17431,N_17815);
xnor U18385 (N_18385,N_17458,N_17260);
xnor U18386 (N_18386,N_17707,N_17863);
nand U18387 (N_18387,N_17841,N_17086);
xnor U18388 (N_18388,N_17462,N_17799);
or U18389 (N_18389,N_17045,N_17120);
xnor U18390 (N_18390,N_17248,N_17123);
nor U18391 (N_18391,N_17277,N_17279);
and U18392 (N_18392,N_17622,N_17689);
and U18393 (N_18393,N_17112,N_17085);
or U18394 (N_18394,N_17744,N_17051);
nand U18395 (N_18395,N_17713,N_17259);
nand U18396 (N_18396,N_17660,N_17270);
nand U18397 (N_18397,N_17545,N_17666);
and U18398 (N_18398,N_17556,N_17640);
and U18399 (N_18399,N_17634,N_17958);
nand U18400 (N_18400,N_17477,N_17133);
xnor U18401 (N_18401,N_17159,N_17428);
nor U18402 (N_18402,N_17315,N_17950);
nand U18403 (N_18403,N_17929,N_17710);
and U18404 (N_18404,N_17831,N_17258);
xor U18405 (N_18405,N_17592,N_17670);
nor U18406 (N_18406,N_17302,N_17095);
and U18407 (N_18407,N_17075,N_17411);
nor U18408 (N_18408,N_17967,N_17011);
nand U18409 (N_18409,N_17464,N_17989);
xnor U18410 (N_18410,N_17484,N_17940);
xor U18411 (N_18411,N_17285,N_17442);
and U18412 (N_18412,N_17224,N_17538);
nor U18413 (N_18413,N_17391,N_17288);
xnor U18414 (N_18414,N_17192,N_17068);
xnor U18415 (N_18415,N_17295,N_17007);
nand U18416 (N_18416,N_17173,N_17363);
and U18417 (N_18417,N_17735,N_17919);
nand U18418 (N_18418,N_17977,N_17301);
or U18419 (N_18419,N_17040,N_17602);
nand U18420 (N_18420,N_17712,N_17182);
nand U18421 (N_18421,N_17074,N_17540);
or U18422 (N_18422,N_17261,N_17136);
and U18423 (N_18423,N_17811,N_17709);
xnor U18424 (N_18424,N_17263,N_17862);
or U18425 (N_18425,N_17663,N_17820);
or U18426 (N_18426,N_17053,N_17674);
nand U18427 (N_18427,N_17698,N_17868);
nor U18428 (N_18428,N_17895,N_17530);
nor U18429 (N_18429,N_17555,N_17782);
or U18430 (N_18430,N_17896,N_17972);
nor U18431 (N_18431,N_17174,N_17132);
nand U18432 (N_18432,N_17022,N_17419);
nor U18433 (N_18433,N_17188,N_17603);
and U18434 (N_18434,N_17190,N_17372);
xnor U18435 (N_18435,N_17223,N_17913);
and U18436 (N_18436,N_17579,N_17436);
xnor U18437 (N_18437,N_17881,N_17573);
or U18438 (N_18438,N_17693,N_17092);
or U18439 (N_18439,N_17148,N_17034);
nor U18440 (N_18440,N_17816,N_17168);
xor U18441 (N_18441,N_17104,N_17335);
nand U18442 (N_18442,N_17366,N_17418);
or U18443 (N_18443,N_17122,N_17638);
nor U18444 (N_18444,N_17834,N_17757);
nor U18445 (N_18445,N_17137,N_17951);
nor U18446 (N_18446,N_17571,N_17849);
or U18447 (N_18447,N_17793,N_17544);
nor U18448 (N_18448,N_17894,N_17533);
or U18449 (N_18449,N_17559,N_17160);
xnor U18450 (N_18450,N_17835,N_17679);
or U18451 (N_18451,N_17770,N_17767);
or U18452 (N_18452,N_17911,N_17269);
xnor U18453 (N_18453,N_17527,N_17024);
and U18454 (N_18454,N_17407,N_17496);
xor U18455 (N_18455,N_17778,N_17879);
or U18456 (N_18456,N_17765,N_17535);
nand U18457 (N_18457,N_17293,N_17764);
or U18458 (N_18458,N_17546,N_17900);
or U18459 (N_18459,N_17723,N_17529);
nand U18460 (N_18460,N_17149,N_17734);
or U18461 (N_18461,N_17843,N_17523);
xnor U18462 (N_18462,N_17233,N_17560);
or U18463 (N_18463,N_17943,N_17861);
xnor U18464 (N_18464,N_17352,N_17643);
or U18465 (N_18465,N_17466,N_17389);
or U18466 (N_18466,N_17097,N_17070);
and U18467 (N_18467,N_17298,N_17597);
nor U18468 (N_18468,N_17066,N_17456);
nand U18469 (N_18469,N_17257,N_17994);
or U18470 (N_18470,N_17119,N_17601);
nand U18471 (N_18471,N_17673,N_17153);
and U18472 (N_18472,N_17856,N_17300);
xnor U18473 (N_18473,N_17183,N_17524);
or U18474 (N_18474,N_17320,N_17409);
or U18475 (N_18475,N_17930,N_17509);
or U18476 (N_18476,N_17899,N_17130);
or U18477 (N_18477,N_17504,N_17326);
and U18478 (N_18478,N_17828,N_17954);
and U18479 (N_18479,N_17124,N_17207);
xnor U18480 (N_18480,N_17347,N_17848);
nand U18481 (N_18481,N_17412,N_17454);
nand U18482 (N_18482,N_17499,N_17121);
and U18483 (N_18483,N_17935,N_17891);
or U18484 (N_18484,N_17818,N_17910);
xnor U18485 (N_18485,N_17163,N_17126);
xnor U18486 (N_18486,N_17611,N_17583);
nand U18487 (N_18487,N_17983,N_17826);
xor U18488 (N_18488,N_17485,N_17324);
nand U18489 (N_18489,N_17858,N_17692);
and U18490 (N_18490,N_17154,N_17522);
nand U18491 (N_18491,N_17369,N_17388);
and U18492 (N_18492,N_17317,N_17234);
or U18493 (N_18493,N_17405,N_17628);
xnor U18494 (N_18494,N_17531,N_17708);
xnor U18495 (N_18495,N_17872,N_17857);
or U18496 (N_18496,N_17071,N_17373);
or U18497 (N_18497,N_17004,N_17569);
nor U18498 (N_18498,N_17226,N_17822);
nor U18499 (N_18499,N_17932,N_17978);
nor U18500 (N_18500,N_17400,N_17375);
or U18501 (N_18501,N_17310,N_17524);
and U18502 (N_18502,N_17466,N_17450);
or U18503 (N_18503,N_17385,N_17969);
nand U18504 (N_18504,N_17200,N_17864);
nor U18505 (N_18505,N_17109,N_17395);
nor U18506 (N_18506,N_17966,N_17730);
xor U18507 (N_18507,N_17587,N_17196);
nand U18508 (N_18508,N_17545,N_17870);
xor U18509 (N_18509,N_17523,N_17684);
and U18510 (N_18510,N_17459,N_17219);
nor U18511 (N_18511,N_17837,N_17926);
xnor U18512 (N_18512,N_17877,N_17634);
nor U18513 (N_18513,N_17678,N_17877);
xor U18514 (N_18514,N_17870,N_17063);
and U18515 (N_18515,N_17375,N_17965);
nand U18516 (N_18516,N_17188,N_17190);
xor U18517 (N_18517,N_17571,N_17613);
nand U18518 (N_18518,N_17962,N_17755);
xnor U18519 (N_18519,N_17028,N_17772);
or U18520 (N_18520,N_17620,N_17240);
nand U18521 (N_18521,N_17926,N_17540);
or U18522 (N_18522,N_17487,N_17935);
nor U18523 (N_18523,N_17112,N_17070);
nand U18524 (N_18524,N_17756,N_17079);
xor U18525 (N_18525,N_17731,N_17589);
nor U18526 (N_18526,N_17060,N_17012);
nand U18527 (N_18527,N_17666,N_17389);
xnor U18528 (N_18528,N_17018,N_17232);
xnor U18529 (N_18529,N_17360,N_17578);
and U18530 (N_18530,N_17306,N_17537);
xor U18531 (N_18531,N_17822,N_17357);
nor U18532 (N_18532,N_17033,N_17872);
nor U18533 (N_18533,N_17654,N_17817);
xor U18534 (N_18534,N_17101,N_17278);
and U18535 (N_18535,N_17837,N_17905);
nor U18536 (N_18536,N_17007,N_17916);
xor U18537 (N_18537,N_17881,N_17851);
or U18538 (N_18538,N_17120,N_17003);
xor U18539 (N_18539,N_17219,N_17024);
and U18540 (N_18540,N_17675,N_17996);
nand U18541 (N_18541,N_17257,N_17062);
or U18542 (N_18542,N_17557,N_17742);
nor U18543 (N_18543,N_17375,N_17418);
xor U18544 (N_18544,N_17587,N_17876);
and U18545 (N_18545,N_17367,N_17883);
nor U18546 (N_18546,N_17848,N_17874);
nor U18547 (N_18547,N_17621,N_17991);
nand U18548 (N_18548,N_17836,N_17329);
and U18549 (N_18549,N_17391,N_17663);
nor U18550 (N_18550,N_17215,N_17345);
nand U18551 (N_18551,N_17526,N_17888);
nand U18552 (N_18552,N_17569,N_17508);
nand U18553 (N_18553,N_17495,N_17792);
and U18554 (N_18554,N_17794,N_17077);
nor U18555 (N_18555,N_17871,N_17956);
or U18556 (N_18556,N_17836,N_17082);
and U18557 (N_18557,N_17546,N_17276);
or U18558 (N_18558,N_17848,N_17062);
and U18559 (N_18559,N_17998,N_17697);
xnor U18560 (N_18560,N_17243,N_17624);
nand U18561 (N_18561,N_17175,N_17691);
xor U18562 (N_18562,N_17019,N_17898);
nand U18563 (N_18563,N_17113,N_17751);
xor U18564 (N_18564,N_17820,N_17393);
and U18565 (N_18565,N_17545,N_17358);
xnor U18566 (N_18566,N_17373,N_17694);
nor U18567 (N_18567,N_17167,N_17982);
xnor U18568 (N_18568,N_17442,N_17054);
xnor U18569 (N_18569,N_17220,N_17944);
and U18570 (N_18570,N_17476,N_17190);
nand U18571 (N_18571,N_17876,N_17338);
nor U18572 (N_18572,N_17381,N_17297);
xnor U18573 (N_18573,N_17106,N_17138);
nand U18574 (N_18574,N_17618,N_17801);
and U18575 (N_18575,N_17069,N_17646);
nand U18576 (N_18576,N_17471,N_17564);
nand U18577 (N_18577,N_17120,N_17762);
and U18578 (N_18578,N_17278,N_17448);
nand U18579 (N_18579,N_17183,N_17396);
or U18580 (N_18580,N_17319,N_17754);
or U18581 (N_18581,N_17842,N_17552);
nor U18582 (N_18582,N_17390,N_17505);
and U18583 (N_18583,N_17113,N_17490);
nor U18584 (N_18584,N_17706,N_17522);
and U18585 (N_18585,N_17892,N_17444);
nand U18586 (N_18586,N_17477,N_17597);
nor U18587 (N_18587,N_17074,N_17474);
nand U18588 (N_18588,N_17304,N_17449);
xor U18589 (N_18589,N_17506,N_17271);
and U18590 (N_18590,N_17579,N_17006);
and U18591 (N_18591,N_17393,N_17646);
nand U18592 (N_18592,N_17015,N_17516);
xnor U18593 (N_18593,N_17710,N_17108);
nand U18594 (N_18594,N_17126,N_17292);
or U18595 (N_18595,N_17585,N_17023);
or U18596 (N_18596,N_17195,N_17413);
or U18597 (N_18597,N_17317,N_17242);
nor U18598 (N_18598,N_17854,N_17205);
nand U18599 (N_18599,N_17639,N_17637);
and U18600 (N_18600,N_17547,N_17608);
and U18601 (N_18601,N_17145,N_17108);
or U18602 (N_18602,N_17770,N_17757);
nand U18603 (N_18603,N_17463,N_17240);
and U18604 (N_18604,N_17149,N_17172);
nor U18605 (N_18605,N_17625,N_17458);
nand U18606 (N_18606,N_17964,N_17427);
nor U18607 (N_18607,N_17243,N_17787);
xnor U18608 (N_18608,N_17547,N_17990);
nand U18609 (N_18609,N_17544,N_17221);
nor U18610 (N_18610,N_17624,N_17580);
nor U18611 (N_18611,N_17916,N_17514);
or U18612 (N_18612,N_17040,N_17355);
or U18613 (N_18613,N_17833,N_17823);
nor U18614 (N_18614,N_17054,N_17584);
or U18615 (N_18615,N_17226,N_17257);
xnor U18616 (N_18616,N_17418,N_17019);
nand U18617 (N_18617,N_17724,N_17293);
xnor U18618 (N_18618,N_17714,N_17867);
or U18619 (N_18619,N_17381,N_17182);
xor U18620 (N_18620,N_17094,N_17426);
or U18621 (N_18621,N_17898,N_17406);
or U18622 (N_18622,N_17739,N_17646);
or U18623 (N_18623,N_17800,N_17109);
or U18624 (N_18624,N_17924,N_17168);
xor U18625 (N_18625,N_17915,N_17649);
and U18626 (N_18626,N_17374,N_17985);
or U18627 (N_18627,N_17837,N_17051);
nand U18628 (N_18628,N_17153,N_17996);
xnor U18629 (N_18629,N_17216,N_17960);
nor U18630 (N_18630,N_17314,N_17637);
xor U18631 (N_18631,N_17745,N_17843);
nand U18632 (N_18632,N_17433,N_17477);
xor U18633 (N_18633,N_17958,N_17876);
nor U18634 (N_18634,N_17516,N_17113);
or U18635 (N_18635,N_17046,N_17867);
and U18636 (N_18636,N_17056,N_17769);
nand U18637 (N_18637,N_17221,N_17017);
and U18638 (N_18638,N_17037,N_17088);
nor U18639 (N_18639,N_17816,N_17748);
nand U18640 (N_18640,N_17177,N_17141);
nor U18641 (N_18641,N_17991,N_17700);
xor U18642 (N_18642,N_17556,N_17516);
and U18643 (N_18643,N_17751,N_17914);
xor U18644 (N_18644,N_17129,N_17311);
or U18645 (N_18645,N_17421,N_17455);
nor U18646 (N_18646,N_17199,N_17183);
xnor U18647 (N_18647,N_17681,N_17018);
or U18648 (N_18648,N_17742,N_17871);
nor U18649 (N_18649,N_17958,N_17916);
and U18650 (N_18650,N_17716,N_17173);
nor U18651 (N_18651,N_17081,N_17663);
nand U18652 (N_18652,N_17725,N_17643);
or U18653 (N_18653,N_17862,N_17222);
or U18654 (N_18654,N_17694,N_17196);
nand U18655 (N_18655,N_17920,N_17422);
nand U18656 (N_18656,N_17828,N_17054);
nand U18657 (N_18657,N_17438,N_17361);
and U18658 (N_18658,N_17155,N_17537);
or U18659 (N_18659,N_17253,N_17953);
or U18660 (N_18660,N_17479,N_17901);
or U18661 (N_18661,N_17282,N_17425);
nor U18662 (N_18662,N_17596,N_17266);
and U18663 (N_18663,N_17754,N_17573);
and U18664 (N_18664,N_17323,N_17389);
or U18665 (N_18665,N_17722,N_17750);
xnor U18666 (N_18666,N_17221,N_17775);
nor U18667 (N_18667,N_17025,N_17081);
nand U18668 (N_18668,N_17057,N_17924);
and U18669 (N_18669,N_17126,N_17918);
xnor U18670 (N_18670,N_17258,N_17473);
xnor U18671 (N_18671,N_17262,N_17378);
xnor U18672 (N_18672,N_17306,N_17271);
and U18673 (N_18673,N_17902,N_17688);
xnor U18674 (N_18674,N_17598,N_17928);
and U18675 (N_18675,N_17902,N_17364);
and U18676 (N_18676,N_17875,N_17185);
nand U18677 (N_18677,N_17115,N_17355);
and U18678 (N_18678,N_17015,N_17893);
nor U18679 (N_18679,N_17353,N_17146);
nand U18680 (N_18680,N_17857,N_17231);
xnor U18681 (N_18681,N_17782,N_17303);
nand U18682 (N_18682,N_17610,N_17140);
and U18683 (N_18683,N_17698,N_17007);
xnor U18684 (N_18684,N_17084,N_17536);
nor U18685 (N_18685,N_17117,N_17014);
and U18686 (N_18686,N_17998,N_17102);
or U18687 (N_18687,N_17691,N_17491);
nand U18688 (N_18688,N_17690,N_17904);
nand U18689 (N_18689,N_17919,N_17725);
nor U18690 (N_18690,N_17166,N_17332);
nand U18691 (N_18691,N_17594,N_17465);
and U18692 (N_18692,N_17507,N_17491);
xnor U18693 (N_18693,N_17820,N_17898);
xor U18694 (N_18694,N_17868,N_17737);
nand U18695 (N_18695,N_17857,N_17750);
nor U18696 (N_18696,N_17379,N_17273);
and U18697 (N_18697,N_17519,N_17608);
nand U18698 (N_18698,N_17260,N_17064);
nor U18699 (N_18699,N_17598,N_17795);
nor U18700 (N_18700,N_17230,N_17185);
nor U18701 (N_18701,N_17472,N_17962);
and U18702 (N_18702,N_17352,N_17596);
and U18703 (N_18703,N_17863,N_17270);
and U18704 (N_18704,N_17599,N_17692);
and U18705 (N_18705,N_17395,N_17514);
and U18706 (N_18706,N_17189,N_17689);
or U18707 (N_18707,N_17127,N_17841);
or U18708 (N_18708,N_17624,N_17503);
xor U18709 (N_18709,N_17715,N_17673);
and U18710 (N_18710,N_17813,N_17174);
or U18711 (N_18711,N_17192,N_17693);
nor U18712 (N_18712,N_17414,N_17939);
nand U18713 (N_18713,N_17256,N_17783);
nand U18714 (N_18714,N_17747,N_17258);
and U18715 (N_18715,N_17566,N_17094);
and U18716 (N_18716,N_17317,N_17750);
nor U18717 (N_18717,N_17818,N_17155);
nand U18718 (N_18718,N_17659,N_17086);
or U18719 (N_18719,N_17275,N_17100);
xnor U18720 (N_18720,N_17131,N_17767);
nand U18721 (N_18721,N_17111,N_17622);
nor U18722 (N_18722,N_17969,N_17177);
nor U18723 (N_18723,N_17443,N_17250);
or U18724 (N_18724,N_17911,N_17712);
nand U18725 (N_18725,N_17482,N_17259);
xnor U18726 (N_18726,N_17420,N_17926);
nand U18727 (N_18727,N_17412,N_17307);
and U18728 (N_18728,N_17063,N_17121);
and U18729 (N_18729,N_17323,N_17236);
or U18730 (N_18730,N_17790,N_17605);
xor U18731 (N_18731,N_17054,N_17177);
and U18732 (N_18732,N_17577,N_17067);
xnor U18733 (N_18733,N_17697,N_17984);
xor U18734 (N_18734,N_17666,N_17265);
xor U18735 (N_18735,N_17621,N_17464);
nor U18736 (N_18736,N_17566,N_17904);
nand U18737 (N_18737,N_17704,N_17279);
nor U18738 (N_18738,N_17122,N_17457);
nor U18739 (N_18739,N_17547,N_17129);
nor U18740 (N_18740,N_17545,N_17080);
xnor U18741 (N_18741,N_17384,N_17866);
nand U18742 (N_18742,N_17743,N_17264);
and U18743 (N_18743,N_17509,N_17963);
and U18744 (N_18744,N_17495,N_17433);
and U18745 (N_18745,N_17102,N_17877);
and U18746 (N_18746,N_17419,N_17153);
or U18747 (N_18747,N_17413,N_17827);
and U18748 (N_18748,N_17063,N_17337);
nand U18749 (N_18749,N_17120,N_17124);
nor U18750 (N_18750,N_17458,N_17001);
or U18751 (N_18751,N_17179,N_17735);
and U18752 (N_18752,N_17690,N_17641);
nand U18753 (N_18753,N_17518,N_17072);
nand U18754 (N_18754,N_17016,N_17333);
or U18755 (N_18755,N_17209,N_17947);
and U18756 (N_18756,N_17073,N_17134);
and U18757 (N_18757,N_17392,N_17770);
and U18758 (N_18758,N_17757,N_17900);
and U18759 (N_18759,N_17526,N_17546);
and U18760 (N_18760,N_17850,N_17267);
xnor U18761 (N_18761,N_17577,N_17159);
nand U18762 (N_18762,N_17072,N_17255);
or U18763 (N_18763,N_17615,N_17754);
xnor U18764 (N_18764,N_17432,N_17471);
nand U18765 (N_18765,N_17203,N_17513);
xor U18766 (N_18766,N_17468,N_17251);
xnor U18767 (N_18767,N_17346,N_17155);
or U18768 (N_18768,N_17170,N_17267);
nor U18769 (N_18769,N_17235,N_17568);
and U18770 (N_18770,N_17584,N_17242);
nor U18771 (N_18771,N_17061,N_17895);
xor U18772 (N_18772,N_17962,N_17941);
xnor U18773 (N_18773,N_17802,N_17332);
nand U18774 (N_18774,N_17148,N_17946);
nor U18775 (N_18775,N_17344,N_17549);
or U18776 (N_18776,N_17490,N_17846);
nand U18777 (N_18777,N_17133,N_17100);
and U18778 (N_18778,N_17203,N_17477);
xor U18779 (N_18779,N_17951,N_17409);
xor U18780 (N_18780,N_17108,N_17562);
and U18781 (N_18781,N_17152,N_17176);
xor U18782 (N_18782,N_17343,N_17419);
nor U18783 (N_18783,N_17455,N_17189);
xor U18784 (N_18784,N_17270,N_17348);
nand U18785 (N_18785,N_17828,N_17323);
and U18786 (N_18786,N_17630,N_17966);
and U18787 (N_18787,N_17690,N_17146);
and U18788 (N_18788,N_17449,N_17457);
and U18789 (N_18789,N_17913,N_17731);
and U18790 (N_18790,N_17447,N_17253);
nand U18791 (N_18791,N_17663,N_17682);
nor U18792 (N_18792,N_17109,N_17410);
nor U18793 (N_18793,N_17372,N_17117);
nor U18794 (N_18794,N_17162,N_17706);
and U18795 (N_18795,N_17351,N_17878);
nor U18796 (N_18796,N_17240,N_17518);
nor U18797 (N_18797,N_17289,N_17100);
xor U18798 (N_18798,N_17497,N_17069);
xnor U18799 (N_18799,N_17408,N_17959);
xor U18800 (N_18800,N_17931,N_17652);
nand U18801 (N_18801,N_17184,N_17613);
nor U18802 (N_18802,N_17034,N_17167);
nand U18803 (N_18803,N_17713,N_17487);
nand U18804 (N_18804,N_17801,N_17003);
xor U18805 (N_18805,N_17386,N_17128);
nand U18806 (N_18806,N_17205,N_17034);
or U18807 (N_18807,N_17327,N_17406);
nor U18808 (N_18808,N_17478,N_17922);
nor U18809 (N_18809,N_17802,N_17142);
nand U18810 (N_18810,N_17944,N_17851);
nand U18811 (N_18811,N_17121,N_17118);
and U18812 (N_18812,N_17668,N_17666);
and U18813 (N_18813,N_17955,N_17102);
xor U18814 (N_18814,N_17251,N_17380);
nor U18815 (N_18815,N_17690,N_17457);
nand U18816 (N_18816,N_17850,N_17569);
nand U18817 (N_18817,N_17369,N_17556);
xor U18818 (N_18818,N_17712,N_17718);
xor U18819 (N_18819,N_17756,N_17816);
xnor U18820 (N_18820,N_17963,N_17906);
or U18821 (N_18821,N_17393,N_17289);
nor U18822 (N_18822,N_17180,N_17934);
or U18823 (N_18823,N_17395,N_17748);
nor U18824 (N_18824,N_17272,N_17908);
or U18825 (N_18825,N_17224,N_17413);
nand U18826 (N_18826,N_17894,N_17865);
nor U18827 (N_18827,N_17611,N_17588);
xnor U18828 (N_18828,N_17757,N_17529);
and U18829 (N_18829,N_17703,N_17266);
nand U18830 (N_18830,N_17869,N_17785);
or U18831 (N_18831,N_17628,N_17361);
xor U18832 (N_18832,N_17644,N_17862);
xor U18833 (N_18833,N_17433,N_17777);
or U18834 (N_18834,N_17267,N_17200);
nand U18835 (N_18835,N_17477,N_17484);
and U18836 (N_18836,N_17327,N_17417);
nand U18837 (N_18837,N_17075,N_17143);
nor U18838 (N_18838,N_17354,N_17880);
nand U18839 (N_18839,N_17072,N_17741);
nand U18840 (N_18840,N_17595,N_17260);
nor U18841 (N_18841,N_17401,N_17475);
xnor U18842 (N_18842,N_17441,N_17450);
or U18843 (N_18843,N_17538,N_17707);
or U18844 (N_18844,N_17476,N_17661);
and U18845 (N_18845,N_17124,N_17858);
nor U18846 (N_18846,N_17784,N_17300);
or U18847 (N_18847,N_17154,N_17733);
nand U18848 (N_18848,N_17984,N_17462);
xnor U18849 (N_18849,N_17462,N_17675);
and U18850 (N_18850,N_17617,N_17085);
xnor U18851 (N_18851,N_17321,N_17109);
or U18852 (N_18852,N_17588,N_17548);
nor U18853 (N_18853,N_17095,N_17960);
or U18854 (N_18854,N_17781,N_17963);
nand U18855 (N_18855,N_17934,N_17373);
or U18856 (N_18856,N_17889,N_17626);
or U18857 (N_18857,N_17927,N_17529);
or U18858 (N_18858,N_17596,N_17192);
nand U18859 (N_18859,N_17746,N_17903);
nor U18860 (N_18860,N_17725,N_17855);
and U18861 (N_18861,N_17615,N_17757);
nand U18862 (N_18862,N_17110,N_17802);
nor U18863 (N_18863,N_17914,N_17552);
nand U18864 (N_18864,N_17377,N_17892);
and U18865 (N_18865,N_17225,N_17097);
nand U18866 (N_18866,N_17155,N_17755);
and U18867 (N_18867,N_17705,N_17380);
or U18868 (N_18868,N_17262,N_17239);
and U18869 (N_18869,N_17449,N_17838);
xor U18870 (N_18870,N_17242,N_17895);
or U18871 (N_18871,N_17635,N_17620);
nand U18872 (N_18872,N_17206,N_17635);
xor U18873 (N_18873,N_17067,N_17080);
and U18874 (N_18874,N_17599,N_17169);
and U18875 (N_18875,N_17832,N_17743);
xor U18876 (N_18876,N_17383,N_17891);
xnor U18877 (N_18877,N_17371,N_17238);
nand U18878 (N_18878,N_17551,N_17896);
nor U18879 (N_18879,N_17455,N_17811);
or U18880 (N_18880,N_17133,N_17325);
or U18881 (N_18881,N_17278,N_17502);
or U18882 (N_18882,N_17598,N_17697);
nand U18883 (N_18883,N_17076,N_17456);
nand U18884 (N_18884,N_17456,N_17627);
nor U18885 (N_18885,N_17509,N_17387);
nor U18886 (N_18886,N_17195,N_17864);
nor U18887 (N_18887,N_17365,N_17561);
nor U18888 (N_18888,N_17683,N_17980);
nor U18889 (N_18889,N_17487,N_17893);
and U18890 (N_18890,N_17837,N_17409);
nand U18891 (N_18891,N_17027,N_17420);
xor U18892 (N_18892,N_17687,N_17144);
or U18893 (N_18893,N_17673,N_17931);
and U18894 (N_18894,N_17446,N_17892);
nor U18895 (N_18895,N_17118,N_17997);
or U18896 (N_18896,N_17577,N_17493);
or U18897 (N_18897,N_17646,N_17969);
or U18898 (N_18898,N_17717,N_17569);
xor U18899 (N_18899,N_17314,N_17302);
nor U18900 (N_18900,N_17449,N_17997);
nand U18901 (N_18901,N_17397,N_17183);
nand U18902 (N_18902,N_17092,N_17411);
and U18903 (N_18903,N_17324,N_17187);
xnor U18904 (N_18904,N_17048,N_17787);
and U18905 (N_18905,N_17115,N_17708);
xnor U18906 (N_18906,N_17458,N_17043);
xor U18907 (N_18907,N_17306,N_17623);
nor U18908 (N_18908,N_17842,N_17142);
or U18909 (N_18909,N_17248,N_17080);
and U18910 (N_18910,N_17733,N_17888);
nand U18911 (N_18911,N_17591,N_17860);
nor U18912 (N_18912,N_17605,N_17837);
nand U18913 (N_18913,N_17294,N_17935);
xor U18914 (N_18914,N_17947,N_17376);
nand U18915 (N_18915,N_17712,N_17238);
nor U18916 (N_18916,N_17448,N_17792);
xnor U18917 (N_18917,N_17948,N_17130);
and U18918 (N_18918,N_17465,N_17331);
and U18919 (N_18919,N_17066,N_17690);
nor U18920 (N_18920,N_17469,N_17324);
nor U18921 (N_18921,N_17343,N_17408);
nor U18922 (N_18922,N_17094,N_17082);
nand U18923 (N_18923,N_17847,N_17224);
nor U18924 (N_18924,N_17996,N_17707);
or U18925 (N_18925,N_17430,N_17278);
or U18926 (N_18926,N_17683,N_17906);
or U18927 (N_18927,N_17970,N_17623);
xor U18928 (N_18928,N_17016,N_17623);
nor U18929 (N_18929,N_17203,N_17164);
nand U18930 (N_18930,N_17667,N_17152);
nand U18931 (N_18931,N_17619,N_17840);
xnor U18932 (N_18932,N_17392,N_17038);
xnor U18933 (N_18933,N_17897,N_17815);
nand U18934 (N_18934,N_17607,N_17194);
and U18935 (N_18935,N_17936,N_17737);
nand U18936 (N_18936,N_17959,N_17699);
nor U18937 (N_18937,N_17647,N_17294);
or U18938 (N_18938,N_17932,N_17209);
and U18939 (N_18939,N_17731,N_17127);
and U18940 (N_18940,N_17913,N_17565);
or U18941 (N_18941,N_17946,N_17229);
nand U18942 (N_18942,N_17466,N_17080);
or U18943 (N_18943,N_17630,N_17352);
nor U18944 (N_18944,N_17799,N_17775);
xor U18945 (N_18945,N_17467,N_17151);
xnor U18946 (N_18946,N_17015,N_17781);
nand U18947 (N_18947,N_17554,N_17227);
nor U18948 (N_18948,N_17130,N_17671);
or U18949 (N_18949,N_17863,N_17159);
or U18950 (N_18950,N_17159,N_17600);
nand U18951 (N_18951,N_17966,N_17085);
or U18952 (N_18952,N_17421,N_17798);
nand U18953 (N_18953,N_17694,N_17767);
xor U18954 (N_18954,N_17317,N_17830);
nor U18955 (N_18955,N_17465,N_17177);
and U18956 (N_18956,N_17579,N_17443);
nand U18957 (N_18957,N_17852,N_17263);
nor U18958 (N_18958,N_17739,N_17962);
nor U18959 (N_18959,N_17133,N_17082);
or U18960 (N_18960,N_17421,N_17794);
or U18961 (N_18961,N_17733,N_17305);
and U18962 (N_18962,N_17185,N_17500);
and U18963 (N_18963,N_17868,N_17157);
xor U18964 (N_18964,N_17880,N_17592);
nor U18965 (N_18965,N_17062,N_17130);
and U18966 (N_18966,N_17660,N_17875);
nor U18967 (N_18967,N_17441,N_17964);
nand U18968 (N_18968,N_17426,N_17836);
and U18969 (N_18969,N_17999,N_17132);
and U18970 (N_18970,N_17533,N_17595);
or U18971 (N_18971,N_17105,N_17538);
or U18972 (N_18972,N_17334,N_17080);
and U18973 (N_18973,N_17945,N_17667);
nor U18974 (N_18974,N_17260,N_17818);
or U18975 (N_18975,N_17697,N_17857);
and U18976 (N_18976,N_17023,N_17644);
nor U18977 (N_18977,N_17517,N_17512);
nand U18978 (N_18978,N_17190,N_17250);
nor U18979 (N_18979,N_17441,N_17924);
nor U18980 (N_18980,N_17812,N_17304);
nor U18981 (N_18981,N_17021,N_17352);
and U18982 (N_18982,N_17345,N_17766);
nand U18983 (N_18983,N_17710,N_17801);
xnor U18984 (N_18984,N_17114,N_17399);
and U18985 (N_18985,N_17131,N_17787);
nand U18986 (N_18986,N_17757,N_17485);
and U18987 (N_18987,N_17235,N_17655);
nand U18988 (N_18988,N_17301,N_17347);
or U18989 (N_18989,N_17116,N_17678);
nand U18990 (N_18990,N_17162,N_17198);
or U18991 (N_18991,N_17320,N_17554);
and U18992 (N_18992,N_17540,N_17556);
xnor U18993 (N_18993,N_17947,N_17852);
nand U18994 (N_18994,N_17864,N_17787);
and U18995 (N_18995,N_17472,N_17979);
nor U18996 (N_18996,N_17691,N_17258);
and U18997 (N_18997,N_17019,N_17053);
nand U18998 (N_18998,N_17769,N_17099);
xor U18999 (N_18999,N_17583,N_17627);
nand U19000 (N_19000,N_18410,N_18160);
or U19001 (N_19001,N_18645,N_18346);
nand U19002 (N_19002,N_18916,N_18469);
nand U19003 (N_19003,N_18845,N_18405);
nand U19004 (N_19004,N_18579,N_18178);
nand U19005 (N_19005,N_18045,N_18978);
or U19006 (N_19006,N_18325,N_18058);
and U19007 (N_19007,N_18561,N_18092);
nand U19008 (N_19008,N_18713,N_18698);
xnor U19009 (N_19009,N_18049,N_18208);
nor U19010 (N_19010,N_18486,N_18803);
nand U19011 (N_19011,N_18913,N_18467);
nor U19012 (N_19012,N_18810,N_18417);
or U19013 (N_19013,N_18548,N_18905);
or U19014 (N_19014,N_18990,N_18890);
nand U19015 (N_19015,N_18127,N_18695);
and U19016 (N_19016,N_18195,N_18466);
nand U19017 (N_19017,N_18721,N_18289);
nor U19018 (N_19018,N_18910,N_18353);
nand U19019 (N_19019,N_18416,N_18511);
or U19020 (N_19020,N_18196,N_18229);
and U19021 (N_19021,N_18936,N_18595);
and U19022 (N_19022,N_18268,N_18024);
and U19023 (N_19023,N_18534,N_18737);
nand U19024 (N_19024,N_18016,N_18758);
xnor U19025 (N_19025,N_18538,N_18349);
nand U19026 (N_19026,N_18621,N_18592);
xnor U19027 (N_19027,N_18658,N_18980);
xor U19028 (N_19028,N_18309,N_18821);
nand U19029 (N_19029,N_18902,N_18025);
xor U19030 (N_19030,N_18341,N_18888);
or U19031 (N_19031,N_18661,N_18403);
nor U19032 (N_19032,N_18773,N_18081);
and U19033 (N_19033,N_18272,N_18568);
or U19034 (N_19034,N_18523,N_18026);
or U19035 (N_19035,N_18998,N_18763);
and U19036 (N_19036,N_18542,N_18067);
nand U19037 (N_19037,N_18626,N_18391);
and U19038 (N_19038,N_18857,N_18720);
nand U19039 (N_19039,N_18787,N_18244);
or U19040 (N_19040,N_18488,N_18679);
or U19041 (N_19041,N_18318,N_18370);
or U19042 (N_19042,N_18076,N_18334);
nand U19043 (N_19043,N_18572,N_18893);
nand U19044 (N_19044,N_18085,N_18168);
nand U19045 (N_19045,N_18751,N_18671);
or U19046 (N_19046,N_18456,N_18735);
nand U19047 (N_19047,N_18977,N_18828);
or U19048 (N_19048,N_18940,N_18146);
nand U19049 (N_19049,N_18794,N_18419);
xnor U19050 (N_19050,N_18443,N_18131);
nor U19051 (N_19051,N_18322,N_18220);
nand U19052 (N_19052,N_18188,N_18840);
or U19053 (N_19053,N_18526,N_18447);
and U19054 (N_19054,N_18429,N_18694);
xnor U19055 (N_19055,N_18313,N_18264);
or U19056 (N_19056,N_18675,N_18424);
and U19057 (N_19057,N_18769,N_18212);
or U19058 (N_19058,N_18701,N_18121);
xor U19059 (N_19059,N_18051,N_18225);
or U19060 (N_19060,N_18554,N_18906);
nor U19061 (N_19061,N_18964,N_18152);
nand U19062 (N_19062,N_18907,N_18169);
nand U19063 (N_19063,N_18375,N_18932);
xor U19064 (N_19064,N_18861,N_18185);
or U19065 (N_19065,N_18749,N_18125);
nand U19066 (N_19066,N_18611,N_18569);
nor U19067 (N_19067,N_18173,N_18966);
and U19068 (N_19068,N_18428,N_18480);
nand U19069 (N_19069,N_18000,N_18851);
nand U19070 (N_19070,N_18544,N_18266);
xnor U19071 (N_19071,N_18054,N_18603);
nand U19072 (N_19072,N_18514,N_18065);
nand U19073 (N_19073,N_18759,N_18528);
xnor U19074 (N_19074,N_18609,N_18471);
and U19075 (N_19075,N_18598,N_18764);
or U19076 (N_19076,N_18739,N_18925);
nand U19077 (N_19077,N_18032,N_18604);
and U19078 (N_19078,N_18638,N_18068);
and U19079 (N_19079,N_18882,N_18060);
xnor U19080 (N_19080,N_18253,N_18867);
xnor U19081 (N_19081,N_18394,N_18435);
xnor U19082 (N_19082,N_18733,N_18439);
or U19083 (N_19083,N_18754,N_18690);
and U19084 (N_19084,N_18014,N_18423);
and U19085 (N_19085,N_18223,N_18580);
nand U19086 (N_19086,N_18130,N_18513);
nand U19087 (N_19087,N_18159,N_18140);
or U19088 (N_19088,N_18390,N_18649);
xnor U19089 (N_19089,N_18317,N_18702);
nand U19090 (N_19090,N_18101,N_18899);
xor U19091 (N_19091,N_18897,N_18617);
nand U19092 (N_19092,N_18942,N_18019);
xor U19093 (N_19093,N_18669,N_18260);
nand U19094 (N_19094,N_18033,N_18017);
and U19095 (N_19095,N_18935,N_18814);
nor U19096 (N_19096,N_18245,N_18472);
nor U19097 (N_19097,N_18089,N_18426);
or U19098 (N_19098,N_18967,N_18619);
xor U19099 (N_19099,N_18321,N_18635);
or U19100 (N_19100,N_18983,N_18445);
or U19101 (N_19101,N_18862,N_18597);
nor U19102 (N_19102,N_18686,N_18736);
nor U19103 (N_19103,N_18356,N_18079);
nor U19104 (N_19104,N_18292,N_18252);
nor U19105 (N_19105,N_18262,N_18396);
xor U19106 (N_19106,N_18459,N_18107);
nor U19107 (N_19107,N_18271,N_18704);
nor U19108 (N_19108,N_18259,N_18373);
nor U19109 (N_19109,N_18361,N_18997);
xnor U19110 (N_19110,N_18103,N_18796);
nand U19111 (N_19111,N_18230,N_18194);
nor U19112 (N_19112,N_18279,N_18996);
xnor U19113 (N_19113,N_18023,N_18301);
nand U19114 (N_19114,N_18781,N_18440);
nand U19115 (N_19115,N_18329,N_18873);
xnor U19116 (N_19116,N_18525,N_18653);
or U19117 (N_19117,N_18385,N_18408);
nand U19118 (N_19118,N_18532,N_18643);
nand U19119 (N_19119,N_18712,N_18696);
nor U19120 (N_19120,N_18955,N_18654);
nand U19121 (N_19121,N_18143,N_18540);
and U19122 (N_19122,N_18562,N_18216);
xor U19123 (N_19123,N_18491,N_18944);
nand U19124 (N_19124,N_18400,N_18108);
xor U19125 (N_19125,N_18874,N_18833);
nor U19126 (N_19126,N_18859,N_18830);
and U19127 (N_19127,N_18080,N_18098);
nor U19128 (N_19128,N_18126,N_18247);
and U19129 (N_19129,N_18084,N_18614);
nand U19130 (N_19130,N_18295,N_18601);
and U19131 (N_19131,N_18053,N_18241);
xnor U19132 (N_19132,N_18791,N_18824);
nand U19133 (N_19133,N_18703,N_18633);
and U19134 (N_19134,N_18100,N_18520);
xor U19135 (N_19135,N_18900,N_18681);
xor U19136 (N_19136,N_18761,N_18015);
and U19137 (N_19137,N_18345,N_18339);
xor U19138 (N_19138,N_18254,N_18729);
or U19139 (N_19139,N_18879,N_18506);
and U19140 (N_19140,N_18946,N_18772);
nand U19141 (N_19141,N_18485,N_18564);
and U19142 (N_19142,N_18657,N_18812);
and U19143 (N_19143,N_18574,N_18179);
or U19144 (N_19144,N_18782,N_18578);
and U19145 (N_19145,N_18697,N_18515);
and U19146 (N_19146,N_18559,N_18217);
nand U19147 (N_19147,N_18573,N_18246);
and U19148 (N_19148,N_18880,N_18930);
nor U19149 (N_19149,N_18755,N_18096);
and U19150 (N_19150,N_18853,N_18470);
nor U19151 (N_19151,N_18211,N_18717);
or U19152 (N_19152,N_18363,N_18489);
nor U19153 (N_19153,N_18043,N_18004);
nor U19154 (N_19154,N_18433,N_18995);
nor U19155 (N_19155,N_18668,N_18006);
or U19156 (N_19156,N_18177,N_18516);
nand U19157 (N_19157,N_18806,N_18502);
nand U19158 (N_19158,N_18786,N_18748);
nand U19159 (N_19159,N_18818,N_18872);
xor U19160 (N_19160,N_18756,N_18109);
nand U19161 (N_19161,N_18113,N_18093);
and U19162 (N_19162,N_18347,N_18765);
and U19163 (N_19163,N_18280,N_18778);
nor U19164 (N_19164,N_18293,N_18151);
nand U19165 (N_19165,N_18915,N_18959);
xnor U19166 (N_19166,N_18308,N_18413);
or U19167 (N_19167,N_18310,N_18945);
or U19168 (N_19168,N_18644,N_18009);
xor U19169 (N_19169,N_18921,N_18203);
xor U19170 (N_19170,N_18599,N_18714);
nand U19171 (N_19171,N_18487,N_18226);
or U19172 (N_19172,N_18961,N_18802);
xnor U19173 (N_19173,N_18029,N_18444);
and U19174 (N_19174,N_18987,N_18132);
xor U19175 (N_19175,N_18425,N_18138);
or U19176 (N_19176,N_18332,N_18157);
xor U19177 (N_19177,N_18665,N_18844);
nor U19178 (N_19178,N_18637,N_18040);
nor U19179 (N_19179,N_18003,N_18360);
nand U19180 (N_19180,N_18210,N_18519);
xor U19181 (N_19181,N_18917,N_18243);
and U19182 (N_19182,N_18744,N_18642);
and U19183 (N_19183,N_18077,N_18402);
and U19184 (N_19184,N_18176,N_18386);
and U19185 (N_19185,N_18650,N_18134);
and U19186 (N_19186,N_18481,N_18204);
or U19187 (N_19187,N_18228,N_18021);
or U19188 (N_19188,N_18904,N_18933);
nor U19189 (N_19189,N_18767,N_18112);
nand U19190 (N_19190,N_18458,N_18284);
or U19191 (N_19191,N_18829,N_18815);
and U19192 (N_19192,N_18792,N_18330);
or U19193 (N_19193,N_18813,N_18876);
xnor U19194 (N_19194,N_18706,N_18894);
nor U19195 (N_19195,N_18656,N_18672);
or U19196 (N_19196,N_18199,N_18999);
and U19197 (N_19197,N_18071,N_18184);
or U19198 (N_19198,N_18478,N_18455);
or U19199 (N_19199,N_18868,N_18030);
nand U19200 (N_19200,N_18197,N_18651);
xor U19201 (N_19201,N_18474,N_18594);
and U19202 (N_19202,N_18809,N_18187);
or U19203 (N_19203,N_18832,N_18354);
nor U19204 (N_19204,N_18583,N_18401);
nand U19205 (N_19205,N_18605,N_18531);
nand U19206 (N_19206,N_18189,N_18901);
or U19207 (N_19207,N_18898,N_18783);
and U19208 (N_19208,N_18920,N_18951);
nor U19209 (N_19209,N_18608,N_18409);
xor U19210 (N_19210,N_18547,N_18378);
nor U19211 (N_19211,N_18732,N_18008);
xnor U19212 (N_19212,N_18965,N_18392);
nand U19213 (N_19213,N_18239,N_18726);
xnor U19214 (N_19214,N_18475,N_18227);
or U19215 (N_19215,N_18529,N_18911);
xor U19216 (N_19216,N_18251,N_18105);
xor U19217 (N_19217,N_18206,N_18541);
nand U19218 (N_19218,N_18962,N_18753);
nand U19219 (N_19219,N_18683,N_18795);
or U19220 (N_19220,N_18171,N_18827);
xnor U19221 (N_19221,N_18034,N_18294);
or U19222 (N_19222,N_18070,N_18078);
or U19223 (N_19223,N_18120,N_18449);
nor U19224 (N_19224,N_18490,N_18062);
xnor U19225 (N_19225,N_18274,N_18563);
xnor U19226 (N_19226,N_18046,N_18358);
nor U19227 (N_19227,N_18148,N_18492);
nand U19228 (N_19228,N_18104,N_18261);
or U19229 (N_19229,N_18981,N_18826);
and U19230 (N_19230,N_18359,N_18707);
nand U19231 (N_19231,N_18133,N_18161);
nor U19232 (N_19232,N_18369,N_18170);
nor U19233 (N_19233,N_18750,N_18760);
nand U19234 (N_19234,N_18938,N_18350);
nor U19235 (N_19235,N_18086,N_18801);
or U19236 (N_19236,N_18892,N_18452);
or U19237 (N_19237,N_18632,N_18949);
nand U19238 (N_19238,N_18610,N_18789);
or U19239 (N_19239,N_18710,N_18504);
xor U19240 (N_19240,N_18200,N_18718);
nor U19241 (N_19241,N_18822,N_18856);
xnor U19242 (N_19242,N_18943,N_18087);
or U19243 (N_19243,N_18565,N_18010);
xnor U19244 (N_19244,N_18135,N_18865);
nor U19245 (N_19245,N_18839,N_18670);
nand U19246 (N_19246,N_18473,N_18871);
nor U19247 (N_19247,N_18468,N_18885);
nor U19248 (N_19248,N_18929,N_18555);
xnor U19249 (N_19249,N_18923,N_18287);
or U19250 (N_19250,N_18442,N_18012);
nand U19251 (N_19251,N_18676,N_18388);
xor U19252 (N_19252,N_18201,N_18242);
and U19253 (N_19253,N_18265,N_18664);
xor U19254 (N_19254,N_18588,N_18602);
xor U19255 (N_19255,N_18041,N_18166);
xor U19256 (N_19256,N_18205,N_18835);
xnor U19257 (N_19257,N_18799,N_18581);
or U19258 (N_19258,N_18174,N_18122);
xnor U19259 (N_19259,N_18479,N_18202);
nor U19260 (N_19260,N_18482,N_18465);
xnor U19261 (N_19261,N_18854,N_18512);
xnor U19262 (N_19262,N_18437,N_18947);
xor U19263 (N_19263,N_18631,N_18889);
nand U19264 (N_19264,N_18117,N_18307);
and U19265 (N_19265,N_18044,N_18677);
or U19266 (N_19266,N_18838,N_18807);
xor U19267 (N_19267,N_18155,N_18556);
nand U19268 (N_19268,N_18823,N_18368);
nor U19269 (N_19269,N_18855,N_18537);
xnor U19270 (N_19270,N_18625,N_18319);
nor U19271 (N_19271,N_18118,N_18629);
nand U19272 (N_19272,N_18774,N_18052);
or U19273 (N_19273,N_18066,N_18436);
nor U19274 (N_19274,N_18421,N_18190);
nand U19275 (N_19275,N_18527,N_18285);
and U19276 (N_19276,N_18928,N_18878);
and U19277 (N_19277,N_18454,N_18175);
or U19278 (N_19278,N_18156,N_18150);
and U19279 (N_19279,N_18327,N_18647);
and U19280 (N_19280,N_18976,N_18785);
nor U19281 (N_19281,N_18509,N_18495);
nand U19282 (N_19282,N_18387,N_18914);
or U19283 (N_19283,N_18847,N_18496);
or U19284 (N_19284,N_18498,N_18673);
and U19285 (N_19285,N_18276,N_18711);
xnor U19286 (N_19286,N_18384,N_18142);
nand U19287 (N_19287,N_18110,N_18038);
xor U19288 (N_19288,N_18877,N_18587);
xnor U19289 (N_19289,N_18805,N_18059);
or U19290 (N_19290,N_18094,N_18042);
or U19291 (N_19291,N_18727,N_18483);
nand U19292 (N_19292,N_18970,N_18145);
xnor U19293 (N_19293,N_18887,N_18715);
or U19294 (N_19294,N_18627,N_18406);
xnor U19295 (N_19295,N_18198,N_18517);
nand U19296 (N_19296,N_18881,N_18508);
nand U19297 (N_19297,N_18811,N_18969);
nand U19298 (N_19298,N_18180,N_18507);
and U19299 (N_19299,N_18639,N_18666);
nand U19300 (N_19300,N_18430,N_18357);
nor U19301 (N_19301,N_18992,N_18376);
and U19302 (N_19302,N_18352,N_18411);
xor U19303 (N_19303,N_18766,N_18278);
nor U19304 (N_19304,N_18441,N_18518);
nor U19305 (N_19305,N_18256,N_18323);
nand U19306 (N_19306,N_18734,N_18816);
or U19307 (N_19307,N_18777,N_18738);
xnor U19308 (N_19308,N_18926,N_18073);
xor U19309 (N_19309,N_18493,N_18461);
and U19310 (N_19310,N_18484,N_18628);
nand U19311 (N_19311,N_18343,N_18432);
and U19312 (N_19312,N_18891,N_18296);
xor U19313 (N_19313,N_18404,N_18954);
nor U19314 (N_19314,N_18687,N_18606);
nand U19315 (N_19315,N_18001,N_18640);
and U19316 (N_19316,N_18770,N_18743);
or U19317 (N_19317,N_18273,N_18808);
xor U19318 (N_19318,N_18340,N_18215);
xor U19319 (N_19319,N_18300,N_18374);
nor U19320 (N_19320,N_18072,N_18600);
or U19321 (N_19321,N_18234,N_18963);
or U19322 (N_19322,N_18596,N_18288);
or U19323 (N_19323,N_18699,N_18971);
nand U19324 (N_19324,N_18716,N_18883);
or U19325 (N_19325,N_18613,N_18267);
nand U19326 (N_19326,N_18636,N_18158);
xor U19327 (N_19327,N_18237,N_18018);
and U19328 (N_19328,N_18298,N_18521);
nor U19329 (N_19329,N_18875,N_18324);
nor U19330 (N_19330,N_18972,N_18576);
nand U19331 (N_19331,N_18290,N_18884);
nand U19332 (N_19332,N_18123,N_18377);
nand U19333 (N_19333,N_18869,N_18037);
or U19334 (N_19334,N_18730,N_18723);
nand U19335 (N_19335,N_18922,N_18752);
nand U19336 (N_19336,N_18364,N_18927);
xor U19337 (N_19337,N_18846,N_18589);
or U19338 (N_19338,N_18450,N_18678);
or U19339 (N_19339,N_18591,N_18383);
nor U19340 (N_19340,N_18684,N_18477);
nor U19341 (N_19341,N_18747,N_18530);
nand U19342 (N_19342,N_18870,N_18700);
and U19343 (N_19343,N_18850,N_18372);
nor U19344 (N_19344,N_18790,N_18434);
and U19345 (N_19345,N_18367,N_18616);
and U19346 (N_19346,N_18316,N_18149);
xor U19347 (N_19347,N_18539,N_18007);
nor U19348 (N_19348,N_18866,N_18074);
nor U19349 (N_19349,N_18986,N_18503);
nor U19350 (N_19350,N_18797,N_18097);
and U19351 (N_19351,N_18355,N_18119);
nand U19352 (N_19352,N_18837,N_18545);
nand U19353 (N_19353,N_18849,N_18463);
nand U19354 (N_19354,N_18630,N_18144);
xor U19355 (N_19355,N_18305,N_18039);
xor U19356 (N_19356,N_18618,N_18167);
nand U19357 (N_19357,N_18233,N_18982);
xor U19358 (N_19358,N_18705,N_18036);
and U19359 (N_19359,N_18820,N_18106);
or U19360 (N_19360,N_18584,N_18586);
or U19361 (N_19361,N_18075,N_18953);
nand U19362 (N_19362,N_18800,N_18993);
or U19363 (N_19363,N_18895,N_18934);
or U19364 (N_19364,N_18139,N_18438);
nand U19365 (N_19365,N_18533,N_18543);
nand U19366 (N_19366,N_18379,N_18306);
and U19367 (N_19367,N_18570,N_18817);
nand U19368 (N_19368,N_18919,N_18622);
or U19369 (N_19369,N_18115,N_18741);
nor U19370 (N_19370,N_18864,N_18398);
nand U19371 (N_19371,N_18960,N_18566);
or U19372 (N_19372,N_18218,N_18291);
nor U19373 (N_19373,N_18536,N_18326);
nor U19374 (N_19374,N_18776,N_18956);
xor U19375 (N_19375,N_18431,N_18172);
nand U19376 (N_19376,N_18742,N_18129);
xor U19377 (N_19377,N_18136,N_18240);
or U19378 (N_19378,N_18099,N_18297);
nor U19379 (N_19379,N_18304,N_18090);
nand U19380 (N_19380,N_18775,N_18908);
or U19381 (N_19381,N_18337,N_18446);
xnor U19382 (N_19382,N_18163,N_18623);
and U19383 (N_19383,N_18249,N_18250);
or U19384 (N_19384,N_18020,N_18842);
and U19385 (N_19385,N_18939,N_18724);
nor U19386 (N_19386,N_18464,N_18063);
xor U19387 (N_19387,N_18380,N_18731);
nand U19388 (N_19388,N_18191,N_18371);
xor U19389 (N_19389,N_18111,N_18560);
nor U19390 (N_19390,N_18192,N_18988);
nor U19391 (N_19391,N_18181,N_18558);
nor U19392 (N_19392,N_18153,N_18662);
nor U19393 (N_19393,N_18607,N_18612);
and U19394 (N_19394,N_18255,N_18336);
nor U19395 (N_19395,N_18397,N_18941);
and U19396 (N_19396,N_18083,N_18680);
or U19397 (N_19397,N_18725,N_18270);
nor U19398 (N_19398,N_18128,N_18667);
nor U19399 (N_19399,N_18315,N_18841);
xor U19400 (N_19400,N_18091,N_18193);
and U19401 (N_19401,N_18768,N_18286);
and U19402 (N_19402,N_18395,N_18834);
xor U19403 (N_19403,N_18427,N_18582);
and U19404 (N_19404,N_18975,N_18335);
nor U19405 (N_19405,N_18344,N_18183);
xor U19406 (N_19406,N_18451,N_18028);
or U19407 (N_19407,N_18549,N_18590);
xnor U19408 (N_19408,N_18858,N_18709);
xnor U19409 (N_19409,N_18005,N_18248);
nor U19410 (N_19410,N_18389,N_18641);
xor U19411 (N_19411,N_18674,N_18263);
nor U19412 (N_19412,N_18958,N_18164);
nand U19413 (N_19413,N_18719,N_18124);
or U19414 (N_19414,N_18652,N_18064);
nand U19415 (N_19415,N_18886,N_18303);
and U19416 (N_19416,N_18460,N_18659);
nand U19417 (N_19417,N_18214,N_18994);
xnor U19418 (N_19418,N_18788,N_18277);
or U19419 (N_19419,N_18968,N_18338);
xnor U19420 (N_19420,N_18088,N_18162);
nand U19421 (N_19421,N_18655,N_18989);
and U19422 (N_19422,N_18728,N_18258);
or U19423 (N_19423,N_18047,N_18011);
xor U19424 (N_19424,N_18407,N_18762);
nand U19425 (N_19425,N_18282,N_18804);
nor U19426 (N_19426,N_18550,N_18535);
nor U19427 (N_19427,N_18979,N_18991);
nand U19428 (N_19428,N_18235,N_18257);
nand U19429 (N_19429,N_18577,N_18692);
nand U19430 (N_19430,N_18102,N_18924);
nor U19431 (N_19431,N_18918,N_18974);
nand U19432 (N_19432,N_18333,N_18141);
or U19433 (N_19433,N_18524,N_18056);
nor U19434 (N_19434,N_18620,N_18985);
nor U19435 (N_19435,N_18950,N_18222);
xnor U19436 (N_19436,N_18362,N_18746);
nand U19437 (N_19437,N_18116,N_18784);
xnor U19438 (N_19438,N_18366,N_18476);
nor U19439 (N_19439,N_18311,N_18182);
nand U19440 (N_19440,N_18722,N_18557);
nand U19441 (N_19441,N_18793,N_18412);
nand U19442 (N_19442,N_18740,N_18165);
and U19443 (N_19443,N_18399,N_18660);
nand U19444 (N_19444,N_18422,N_18453);
xnor U19445 (N_19445,N_18779,N_18798);
nor U19446 (N_19446,N_18415,N_18312);
or U19447 (N_19447,N_18448,N_18973);
nand U19448 (N_19448,N_18957,N_18236);
nor U19449 (N_19449,N_18013,N_18393);
xnor U19450 (N_19450,N_18500,N_18382);
or U19451 (N_19451,N_18499,N_18457);
xor U19452 (N_19452,N_18462,N_18501);
or U19453 (N_19453,N_18843,N_18552);
nand U19454 (N_19454,N_18095,N_18615);
nand U19455 (N_19455,N_18551,N_18224);
and U19456 (N_19456,N_18231,N_18624);
nand U19457 (N_19457,N_18320,N_18342);
nand U19458 (N_19458,N_18693,N_18219);
nand U19459 (N_19459,N_18819,N_18546);
nand U19460 (N_19460,N_18348,N_18685);
nand U19461 (N_19461,N_18420,N_18771);
or U19462 (N_19462,N_18909,N_18061);
xor U19463 (N_19463,N_18585,N_18137);
or U19464 (N_19464,N_18836,N_18863);
xor U19465 (N_19465,N_18553,N_18931);
nor U19466 (N_19466,N_18831,N_18522);
nor U19467 (N_19467,N_18069,N_18825);
xor U19468 (N_19468,N_18952,N_18281);
or U19469 (N_19469,N_18213,N_18283);
nor U19470 (N_19470,N_18682,N_18186);
and U19471 (N_19471,N_18351,N_18035);
nand U19472 (N_19472,N_18302,N_18154);
nand U19473 (N_19473,N_18757,N_18494);
or U19474 (N_19474,N_18663,N_18238);
or U19475 (N_19475,N_18057,N_18299);
xor U19476 (N_19476,N_18147,N_18207);
nor U19477 (N_19477,N_18328,N_18984);
or U19478 (N_19478,N_18567,N_18209);
or U19479 (N_19479,N_18593,N_18275);
xnor U19480 (N_19480,N_18221,N_18418);
and U19481 (N_19481,N_18848,N_18708);
nand U19482 (N_19482,N_18575,N_18691);
nor U19483 (N_19483,N_18780,N_18688);
and U19484 (N_19484,N_18912,N_18896);
xor U19485 (N_19485,N_18022,N_18414);
xnor U19486 (N_19486,N_18634,N_18745);
nand U19487 (N_19487,N_18055,N_18027);
and U19488 (N_19488,N_18331,N_18510);
nand U19489 (N_19489,N_18571,N_18852);
or U19490 (N_19490,N_18937,N_18903);
or U19491 (N_19491,N_18948,N_18269);
or U19492 (N_19492,N_18860,N_18381);
and U19493 (N_19493,N_18689,N_18497);
and U19494 (N_19494,N_18114,N_18048);
xor U19495 (N_19495,N_18050,N_18314);
xnor U19496 (N_19496,N_18365,N_18646);
nand U19497 (N_19497,N_18505,N_18031);
or U19498 (N_19498,N_18002,N_18648);
xnor U19499 (N_19499,N_18232,N_18082);
xor U19500 (N_19500,N_18615,N_18640);
nor U19501 (N_19501,N_18952,N_18399);
or U19502 (N_19502,N_18301,N_18731);
nand U19503 (N_19503,N_18653,N_18409);
and U19504 (N_19504,N_18419,N_18640);
xnor U19505 (N_19505,N_18621,N_18912);
xor U19506 (N_19506,N_18875,N_18567);
nor U19507 (N_19507,N_18890,N_18498);
or U19508 (N_19508,N_18952,N_18887);
nor U19509 (N_19509,N_18599,N_18947);
nor U19510 (N_19510,N_18237,N_18719);
nor U19511 (N_19511,N_18685,N_18480);
nand U19512 (N_19512,N_18281,N_18850);
or U19513 (N_19513,N_18201,N_18497);
and U19514 (N_19514,N_18862,N_18751);
xnor U19515 (N_19515,N_18564,N_18588);
nand U19516 (N_19516,N_18389,N_18315);
or U19517 (N_19517,N_18898,N_18090);
xor U19518 (N_19518,N_18650,N_18943);
or U19519 (N_19519,N_18016,N_18734);
xnor U19520 (N_19520,N_18925,N_18995);
and U19521 (N_19521,N_18112,N_18297);
nand U19522 (N_19522,N_18493,N_18148);
and U19523 (N_19523,N_18205,N_18220);
xnor U19524 (N_19524,N_18077,N_18460);
xor U19525 (N_19525,N_18618,N_18071);
nand U19526 (N_19526,N_18024,N_18589);
and U19527 (N_19527,N_18626,N_18379);
nor U19528 (N_19528,N_18554,N_18621);
xnor U19529 (N_19529,N_18020,N_18185);
nand U19530 (N_19530,N_18096,N_18666);
nand U19531 (N_19531,N_18937,N_18915);
or U19532 (N_19532,N_18252,N_18332);
nand U19533 (N_19533,N_18208,N_18864);
nand U19534 (N_19534,N_18453,N_18061);
or U19535 (N_19535,N_18674,N_18310);
nor U19536 (N_19536,N_18331,N_18847);
and U19537 (N_19537,N_18074,N_18726);
nand U19538 (N_19538,N_18594,N_18231);
nand U19539 (N_19539,N_18239,N_18220);
nor U19540 (N_19540,N_18973,N_18702);
or U19541 (N_19541,N_18261,N_18834);
or U19542 (N_19542,N_18309,N_18186);
nor U19543 (N_19543,N_18613,N_18909);
and U19544 (N_19544,N_18261,N_18662);
nor U19545 (N_19545,N_18748,N_18086);
or U19546 (N_19546,N_18584,N_18128);
nand U19547 (N_19547,N_18868,N_18634);
nand U19548 (N_19548,N_18837,N_18979);
xnor U19549 (N_19549,N_18522,N_18142);
nor U19550 (N_19550,N_18837,N_18086);
and U19551 (N_19551,N_18295,N_18574);
or U19552 (N_19552,N_18986,N_18088);
nand U19553 (N_19553,N_18637,N_18638);
nor U19554 (N_19554,N_18165,N_18560);
nor U19555 (N_19555,N_18955,N_18502);
xnor U19556 (N_19556,N_18301,N_18263);
nor U19557 (N_19557,N_18921,N_18408);
and U19558 (N_19558,N_18222,N_18736);
and U19559 (N_19559,N_18477,N_18837);
nand U19560 (N_19560,N_18318,N_18797);
xnor U19561 (N_19561,N_18084,N_18639);
xor U19562 (N_19562,N_18382,N_18602);
and U19563 (N_19563,N_18566,N_18028);
nand U19564 (N_19564,N_18096,N_18091);
nor U19565 (N_19565,N_18291,N_18648);
or U19566 (N_19566,N_18460,N_18591);
xnor U19567 (N_19567,N_18721,N_18888);
nand U19568 (N_19568,N_18114,N_18482);
nor U19569 (N_19569,N_18245,N_18994);
and U19570 (N_19570,N_18405,N_18623);
nand U19571 (N_19571,N_18196,N_18664);
or U19572 (N_19572,N_18819,N_18281);
and U19573 (N_19573,N_18939,N_18065);
nor U19574 (N_19574,N_18824,N_18048);
and U19575 (N_19575,N_18186,N_18165);
xnor U19576 (N_19576,N_18910,N_18145);
xor U19577 (N_19577,N_18172,N_18103);
or U19578 (N_19578,N_18584,N_18555);
or U19579 (N_19579,N_18325,N_18005);
nor U19580 (N_19580,N_18604,N_18445);
xnor U19581 (N_19581,N_18719,N_18806);
nand U19582 (N_19582,N_18955,N_18593);
or U19583 (N_19583,N_18333,N_18847);
and U19584 (N_19584,N_18466,N_18999);
nor U19585 (N_19585,N_18587,N_18478);
nor U19586 (N_19586,N_18417,N_18012);
and U19587 (N_19587,N_18564,N_18771);
and U19588 (N_19588,N_18331,N_18919);
nand U19589 (N_19589,N_18559,N_18581);
and U19590 (N_19590,N_18037,N_18727);
nand U19591 (N_19591,N_18279,N_18861);
nor U19592 (N_19592,N_18628,N_18360);
and U19593 (N_19593,N_18719,N_18422);
or U19594 (N_19594,N_18206,N_18198);
nor U19595 (N_19595,N_18303,N_18148);
xnor U19596 (N_19596,N_18984,N_18921);
and U19597 (N_19597,N_18601,N_18987);
or U19598 (N_19598,N_18518,N_18891);
or U19599 (N_19599,N_18699,N_18713);
or U19600 (N_19600,N_18543,N_18953);
xor U19601 (N_19601,N_18429,N_18521);
or U19602 (N_19602,N_18925,N_18773);
and U19603 (N_19603,N_18744,N_18631);
nand U19604 (N_19604,N_18012,N_18824);
or U19605 (N_19605,N_18704,N_18490);
and U19606 (N_19606,N_18462,N_18095);
nand U19607 (N_19607,N_18338,N_18289);
nand U19608 (N_19608,N_18341,N_18355);
nand U19609 (N_19609,N_18559,N_18930);
nor U19610 (N_19610,N_18774,N_18546);
or U19611 (N_19611,N_18209,N_18159);
xnor U19612 (N_19612,N_18510,N_18758);
nor U19613 (N_19613,N_18371,N_18238);
nand U19614 (N_19614,N_18693,N_18614);
and U19615 (N_19615,N_18977,N_18898);
and U19616 (N_19616,N_18901,N_18678);
nor U19617 (N_19617,N_18238,N_18456);
xor U19618 (N_19618,N_18126,N_18175);
nor U19619 (N_19619,N_18676,N_18453);
and U19620 (N_19620,N_18398,N_18929);
xnor U19621 (N_19621,N_18755,N_18587);
nand U19622 (N_19622,N_18674,N_18006);
and U19623 (N_19623,N_18781,N_18305);
nor U19624 (N_19624,N_18641,N_18172);
nor U19625 (N_19625,N_18671,N_18745);
nand U19626 (N_19626,N_18154,N_18386);
and U19627 (N_19627,N_18382,N_18634);
nor U19628 (N_19628,N_18168,N_18891);
and U19629 (N_19629,N_18105,N_18997);
or U19630 (N_19630,N_18732,N_18742);
and U19631 (N_19631,N_18951,N_18469);
nand U19632 (N_19632,N_18257,N_18983);
or U19633 (N_19633,N_18653,N_18550);
and U19634 (N_19634,N_18451,N_18447);
nor U19635 (N_19635,N_18161,N_18321);
xnor U19636 (N_19636,N_18246,N_18097);
nand U19637 (N_19637,N_18212,N_18771);
and U19638 (N_19638,N_18839,N_18160);
or U19639 (N_19639,N_18483,N_18153);
nand U19640 (N_19640,N_18325,N_18598);
nor U19641 (N_19641,N_18359,N_18784);
and U19642 (N_19642,N_18616,N_18031);
nand U19643 (N_19643,N_18487,N_18249);
nor U19644 (N_19644,N_18257,N_18113);
or U19645 (N_19645,N_18166,N_18979);
nor U19646 (N_19646,N_18081,N_18434);
or U19647 (N_19647,N_18010,N_18950);
or U19648 (N_19648,N_18861,N_18921);
and U19649 (N_19649,N_18328,N_18357);
xor U19650 (N_19650,N_18917,N_18017);
nand U19651 (N_19651,N_18401,N_18846);
or U19652 (N_19652,N_18413,N_18500);
nor U19653 (N_19653,N_18531,N_18242);
or U19654 (N_19654,N_18993,N_18185);
nor U19655 (N_19655,N_18950,N_18722);
nand U19656 (N_19656,N_18467,N_18802);
nand U19657 (N_19657,N_18218,N_18119);
nand U19658 (N_19658,N_18964,N_18809);
nand U19659 (N_19659,N_18078,N_18896);
and U19660 (N_19660,N_18137,N_18370);
or U19661 (N_19661,N_18261,N_18273);
nand U19662 (N_19662,N_18349,N_18351);
or U19663 (N_19663,N_18025,N_18012);
xnor U19664 (N_19664,N_18832,N_18891);
and U19665 (N_19665,N_18248,N_18499);
nand U19666 (N_19666,N_18711,N_18196);
xor U19667 (N_19667,N_18030,N_18478);
and U19668 (N_19668,N_18824,N_18826);
nor U19669 (N_19669,N_18782,N_18773);
or U19670 (N_19670,N_18848,N_18503);
nor U19671 (N_19671,N_18932,N_18056);
xor U19672 (N_19672,N_18749,N_18265);
and U19673 (N_19673,N_18736,N_18894);
nand U19674 (N_19674,N_18346,N_18392);
nand U19675 (N_19675,N_18554,N_18095);
and U19676 (N_19676,N_18198,N_18561);
nand U19677 (N_19677,N_18383,N_18759);
xnor U19678 (N_19678,N_18078,N_18671);
nor U19679 (N_19679,N_18465,N_18724);
and U19680 (N_19680,N_18628,N_18778);
nor U19681 (N_19681,N_18958,N_18070);
or U19682 (N_19682,N_18190,N_18260);
xor U19683 (N_19683,N_18905,N_18103);
or U19684 (N_19684,N_18791,N_18650);
nand U19685 (N_19685,N_18026,N_18636);
nor U19686 (N_19686,N_18542,N_18226);
xor U19687 (N_19687,N_18637,N_18236);
and U19688 (N_19688,N_18323,N_18252);
or U19689 (N_19689,N_18148,N_18762);
and U19690 (N_19690,N_18272,N_18021);
xor U19691 (N_19691,N_18184,N_18159);
nor U19692 (N_19692,N_18149,N_18839);
and U19693 (N_19693,N_18644,N_18042);
and U19694 (N_19694,N_18127,N_18943);
and U19695 (N_19695,N_18630,N_18619);
xor U19696 (N_19696,N_18860,N_18309);
or U19697 (N_19697,N_18801,N_18995);
nand U19698 (N_19698,N_18179,N_18692);
nand U19699 (N_19699,N_18006,N_18411);
xnor U19700 (N_19700,N_18884,N_18094);
and U19701 (N_19701,N_18785,N_18104);
xor U19702 (N_19702,N_18972,N_18834);
xor U19703 (N_19703,N_18263,N_18576);
nor U19704 (N_19704,N_18318,N_18001);
nor U19705 (N_19705,N_18943,N_18640);
and U19706 (N_19706,N_18103,N_18819);
and U19707 (N_19707,N_18897,N_18416);
nand U19708 (N_19708,N_18327,N_18211);
xnor U19709 (N_19709,N_18639,N_18795);
xor U19710 (N_19710,N_18847,N_18926);
xor U19711 (N_19711,N_18832,N_18682);
xor U19712 (N_19712,N_18312,N_18116);
and U19713 (N_19713,N_18503,N_18464);
xnor U19714 (N_19714,N_18113,N_18722);
nor U19715 (N_19715,N_18033,N_18726);
or U19716 (N_19716,N_18152,N_18795);
nand U19717 (N_19717,N_18497,N_18229);
and U19718 (N_19718,N_18394,N_18500);
nor U19719 (N_19719,N_18129,N_18064);
or U19720 (N_19720,N_18015,N_18587);
or U19721 (N_19721,N_18970,N_18543);
nor U19722 (N_19722,N_18501,N_18438);
xor U19723 (N_19723,N_18561,N_18840);
nor U19724 (N_19724,N_18849,N_18599);
nand U19725 (N_19725,N_18694,N_18877);
xor U19726 (N_19726,N_18627,N_18922);
nand U19727 (N_19727,N_18870,N_18215);
and U19728 (N_19728,N_18034,N_18676);
nor U19729 (N_19729,N_18072,N_18412);
and U19730 (N_19730,N_18905,N_18443);
or U19731 (N_19731,N_18567,N_18634);
nand U19732 (N_19732,N_18226,N_18435);
and U19733 (N_19733,N_18658,N_18179);
and U19734 (N_19734,N_18843,N_18518);
nor U19735 (N_19735,N_18579,N_18844);
nor U19736 (N_19736,N_18670,N_18733);
nor U19737 (N_19737,N_18340,N_18348);
nor U19738 (N_19738,N_18214,N_18339);
xnor U19739 (N_19739,N_18794,N_18366);
nand U19740 (N_19740,N_18603,N_18164);
nand U19741 (N_19741,N_18104,N_18908);
or U19742 (N_19742,N_18064,N_18230);
and U19743 (N_19743,N_18761,N_18763);
and U19744 (N_19744,N_18682,N_18201);
nor U19745 (N_19745,N_18946,N_18646);
xor U19746 (N_19746,N_18505,N_18995);
and U19747 (N_19747,N_18495,N_18266);
or U19748 (N_19748,N_18378,N_18644);
and U19749 (N_19749,N_18898,N_18350);
nand U19750 (N_19750,N_18124,N_18034);
nor U19751 (N_19751,N_18338,N_18254);
xor U19752 (N_19752,N_18919,N_18499);
nor U19753 (N_19753,N_18876,N_18486);
or U19754 (N_19754,N_18766,N_18236);
and U19755 (N_19755,N_18624,N_18002);
nand U19756 (N_19756,N_18521,N_18630);
xor U19757 (N_19757,N_18876,N_18614);
nor U19758 (N_19758,N_18226,N_18843);
xnor U19759 (N_19759,N_18882,N_18816);
nand U19760 (N_19760,N_18261,N_18259);
nand U19761 (N_19761,N_18346,N_18251);
nor U19762 (N_19762,N_18200,N_18352);
nor U19763 (N_19763,N_18967,N_18429);
xor U19764 (N_19764,N_18750,N_18579);
nand U19765 (N_19765,N_18399,N_18424);
or U19766 (N_19766,N_18977,N_18190);
or U19767 (N_19767,N_18405,N_18362);
or U19768 (N_19768,N_18173,N_18552);
nand U19769 (N_19769,N_18915,N_18359);
or U19770 (N_19770,N_18748,N_18179);
xnor U19771 (N_19771,N_18563,N_18768);
nand U19772 (N_19772,N_18743,N_18217);
nor U19773 (N_19773,N_18771,N_18072);
nand U19774 (N_19774,N_18088,N_18286);
nand U19775 (N_19775,N_18565,N_18154);
nor U19776 (N_19776,N_18781,N_18908);
nand U19777 (N_19777,N_18263,N_18014);
or U19778 (N_19778,N_18970,N_18826);
nand U19779 (N_19779,N_18839,N_18515);
and U19780 (N_19780,N_18062,N_18980);
xor U19781 (N_19781,N_18473,N_18551);
nor U19782 (N_19782,N_18398,N_18418);
and U19783 (N_19783,N_18882,N_18796);
xor U19784 (N_19784,N_18434,N_18919);
or U19785 (N_19785,N_18425,N_18207);
or U19786 (N_19786,N_18621,N_18197);
xor U19787 (N_19787,N_18754,N_18675);
nand U19788 (N_19788,N_18933,N_18670);
or U19789 (N_19789,N_18075,N_18354);
nand U19790 (N_19790,N_18752,N_18627);
nor U19791 (N_19791,N_18971,N_18205);
xor U19792 (N_19792,N_18236,N_18133);
or U19793 (N_19793,N_18294,N_18982);
nor U19794 (N_19794,N_18989,N_18614);
nor U19795 (N_19795,N_18165,N_18574);
xor U19796 (N_19796,N_18628,N_18624);
nor U19797 (N_19797,N_18258,N_18445);
xor U19798 (N_19798,N_18051,N_18442);
or U19799 (N_19799,N_18989,N_18421);
and U19800 (N_19800,N_18384,N_18748);
or U19801 (N_19801,N_18966,N_18704);
or U19802 (N_19802,N_18331,N_18302);
nand U19803 (N_19803,N_18599,N_18056);
and U19804 (N_19804,N_18717,N_18746);
and U19805 (N_19805,N_18525,N_18941);
and U19806 (N_19806,N_18395,N_18513);
or U19807 (N_19807,N_18913,N_18452);
xnor U19808 (N_19808,N_18210,N_18875);
or U19809 (N_19809,N_18206,N_18497);
nor U19810 (N_19810,N_18257,N_18616);
nand U19811 (N_19811,N_18276,N_18247);
and U19812 (N_19812,N_18214,N_18496);
or U19813 (N_19813,N_18499,N_18312);
and U19814 (N_19814,N_18467,N_18905);
nand U19815 (N_19815,N_18518,N_18866);
and U19816 (N_19816,N_18477,N_18307);
nor U19817 (N_19817,N_18484,N_18015);
xor U19818 (N_19818,N_18755,N_18514);
nand U19819 (N_19819,N_18858,N_18851);
xnor U19820 (N_19820,N_18148,N_18083);
and U19821 (N_19821,N_18193,N_18200);
and U19822 (N_19822,N_18129,N_18601);
and U19823 (N_19823,N_18553,N_18007);
xor U19824 (N_19824,N_18268,N_18600);
or U19825 (N_19825,N_18088,N_18838);
xor U19826 (N_19826,N_18580,N_18405);
nand U19827 (N_19827,N_18680,N_18648);
xor U19828 (N_19828,N_18197,N_18414);
nor U19829 (N_19829,N_18886,N_18792);
and U19830 (N_19830,N_18191,N_18047);
xnor U19831 (N_19831,N_18391,N_18569);
nand U19832 (N_19832,N_18076,N_18952);
xnor U19833 (N_19833,N_18571,N_18033);
xnor U19834 (N_19834,N_18895,N_18894);
or U19835 (N_19835,N_18687,N_18453);
nor U19836 (N_19836,N_18542,N_18408);
nor U19837 (N_19837,N_18052,N_18437);
and U19838 (N_19838,N_18630,N_18180);
or U19839 (N_19839,N_18896,N_18976);
nand U19840 (N_19840,N_18733,N_18849);
and U19841 (N_19841,N_18693,N_18109);
nand U19842 (N_19842,N_18913,N_18618);
and U19843 (N_19843,N_18233,N_18606);
nor U19844 (N_19844,N_18975,N_18046);
or U19845 (N_19845,N_18362,N_18830);
xnor U19846 (N_19846,N_18597,N_18654);
nor U19847 (N_19847,N_18964,N_18773);
xnor U19848 (N_19848,N_18249,N_18595);
nor U19849 (N_19849,N_18009,N_18424);
or U19850 (N_19850,N_18912,N_18430);
nand U19851 (N_19851,N_18137,N_18580);
and U19852 (N_19852,N_18734,N_18120);
xnor U19853 (N_19853,N_18386,N_18707);
xor U19854 (N_19854,N_18111,N_18535);
xor U19855 (N_19855,N_18168,N_18548);
nand U19856 (N_19856,N_18493,N_18196);
xor U19857 (N_19857,N_18842,N_18745);
and U19858 (N_19858,N_18420,N_18763);
nor U19859 (N_19859,N_18735,N_18092);
nor U19860 (N_19860,N_18264,N_18085);
and U19861 (N_19861,N_18427,N_18443);
xor U19862 (N_19862,N_18252,N_18369);
or U19863 (N_19863,N_18011,N_18031);
nand U19864 (N_19864,N_18803,N_18575);
xnor U19865 (N_19865,N_18311,N_18849);
xnor U19866 (N_19866,N_18216,N_18302);
nand U19867 (N_19867,N_18134,N_18094);
and U19868 (N_19868,N_18651,N_18473);
nor U19869 (N_19869,N_18649,N_18682);
xor U19870 (N_19870,N_18649,N_18096);
nor U19871 (N_19871,N_18683,N_18012);
and U19872 (N_19872,N_18222,N_18730);
nor U19873 (N_19873,N_18880,N_18534);
xnor U19874 (N_19874,N_18865,N_18954);
and U19875 (N_19875,N_18310,N_18797);
and U19876 (N_19876,N_18767,N_18110);
or U19877 (N_19877,N_18927,N_18846);
nor U19878 (N_19878,N_18460,N_18158);
or U19879 (N_19879,N_18451,N_18159);
and U19880 (N_19880,N_18668,N_18957);
xnor U19881 (N_19881,N_18617,N_18586);
nor U19882 (N_19882,N_18505,N_18996);
nand U19883 (N_19883,N_18154,N_18028);
nand U19884 (N_19884,N_18678,N_18459);
nor U19885 (N_19885,N_18688,N_18386);
or U19886 (N_19886,N_18926,N_18027);
nand U19887 (N_19887,N_18318,N_18664);
xor U19888 (N_19888,N_18242,N_18694);
and U19889 (N_19889,N_18719,N_18991);
and U19890 (N_19890,N_18120,N_18752);
or U19891 (N_19891,N_18241,N_18920);
and U19892 (N_19892,N_18470,N_18453);
xor U19893 (N_19893,N_18956,N_18717);
or U19894 (N_19894,N_18869,N_18653);
or U19895 (N_19895,N_18131,N_18734);
nand U19896 (N_19896,N_18657,N_18112);
xnor U19897 (N_19897,N_18114,N_18739);
nand U19898 (N_19898,N_18001,N_18829);
or U19899 (N_19899,N_18328,N_18151);
nor U19900 (N_19900,N_18001,N_18326);
and U19901 (N_19901,N_18850,N_18923);
and U19902 (N_19902,N_18497,N_18049);
and U19903 (N_19903,N_18367,N_18012);
nand U19904 (N_19904,N_18413,N_18296);
and U19905 (N_19905,N_18772,N_18822);
nand U19906 (N_19906,N_18585,N_18545);
or U19907 (N_19907,N_18883,N_18776);
or U19908 (N_19908,N_18379,N_18946);
xor U19909 (N_19909,N_18052,N_18941);
xor U19910 (N_19910,N_18305,N_18532);
and U19911 (N_19911,N_18037,N_18153);
or U19912 (N_19912,N_18765,N_18642);
xor U19913 (N_19913,N_18099,N_18261);
and U19914 (N_19914,N_18517,N_18970);
and U19915 (N_19915,N_18235,N_18682);
nor U19916 (N_19916,N_18845,N_18033);
nor U19917 (N_19917,N_18863,N_18970);
or U19918 (N_19918,N_18370,N_18349);
xor U19919 (N_19919,N_18371,N_18385);
nor U19920 (N_19920,N_18055,N_18890);
and U19921 (N_19921,N_18857,N_18867);
or U19922 (N_19922,N_18882,N_18843);
nand U19923 (N_19923,N_18197,N_18151);
nor U19924 (N_19924,N_18153,N_18261);
or U19925 (N_19925,N_18336,N_18625);
nand U19926 (N_19926,N_18052,N_18786);
nor U19927 (N_19927,N_18981,N_18987);
and U19928 (N_19928,N_18860,N_18256);
or U19929 (N_19929,N_18142,N_18872);
xor U19930 (N_19930,N_18407,N_18989);
nand U19931 (N_19931,N_18580,N_18176);
xnor U19932 (N_19932,N_18493,N_18864);
nor U19933 (N_19933,N_18751,N_18082);
nor U19934 (N_19934,N_18365,N_18097);
nor U19935 (N_19935,N_18050,N_18352);
or U19936 (N_19936,N_18560,N_18720);
or U19937 (N_19937,N_18380,N_18093);
xor U19938 (N_19938,N_18177,N_18666);
nor U19939 (N_19939,N_18437,N_18534);
nand U19940 (N_19940,N_18699,N_18965);
and U19941 (N_19941,N_18489,N_18744);
nor U19942 (N_19942,N_18617,N_18771);
nor U19943 (N_19943,N_18549,N_18536);
nor U19944 (N_19944,N_18231,N_18406);
and U19945 (N_19945,N_18577,N_18000);
or U19946 (N_19946,N_18955,N_18258);
xnor U19947 (N_19947,N_18038,N_18620);
or U19948 (N_19948,N_18753,N_18161);
nor U19949 (N_19949,N_18056,N_18491);
nor U19950 (N_19950,N_18953,N_18094);
xor U19951 (N_19951,N_18468,N_18692);
nand U19952 (N_19952,N_18238,N_18147);
xnor U19953 (N_19953,N_18442,N_18541);
or U19954 (N_19954,N_18975,N_18438);
or U19955 (N_19955,N_18438,N_18958);
nand U19956 (N_19956,N_18276,N_18332);
nand U19957 (N_19957,N_18469,N_18115);
and U19958 (N_19958,N_18645,N_18545);
nor U19959 (N_19959,N_18905,N_18282);
nor U19960 (N_19960,N_18493,N_18301);
or U19961 (N_19961,N_18774,N_18445);
nor U19962 (N_19962,N_18262,N_18600);
and U19963 (N_19963,N_18107,N_18643);
nor U19964 (N_19964,N_18820,N_18729);
xor U19965 (N_19965,N_18282,N_18693);
and U19966 (N_19966,N_18495,N_18008);
and U19967 (N_19967,N_18592,N_18522);
nand U19968 (N_19968,N_18796,N_18974);
and U19969 (N_19969,N_18000,N_18937);
xor U19970 (N_19970,N_18681,N_18114);
and U19971 (N_19971,N_18043,N_18677);
xnor U19972 (N_19972,N_18436,N_18237);
xnor U19973 (N_19973,N_18001,N_18653);
nand U19974 (N_19974,N_18617,N_18403);
nand U19975 (N_19975,N_18022,N_18126);
xnor U19976 (N_19976,N_18282,N_18876);
and U19977 (N_19977,N_18874,N_18228);
or U19978 (N_19978,N_18209,N_18892);
or U19979 (N_19979,N_18513,N_18865);
and U19980 (N_19980,N_18047,N_18154);
or U19981 (N_19981,N_18780,N_18644);
or U19982 (N_19982,N_18170,N_18010);
or U19983 (N_19983,N_18335,N_18505);
nor U19984 (N_19984,N_18399,N_18701);
and U19985 (N_19985,N_18396,N_18420);
nor U19986 (N_19986,N_18133,N_18000);
nand U19987 (N_19987,N_18185,N_18680);
xor U19988 (N_19988,N_18744,N_18187);
nor U19989 (N_19989,N_18853,N_18481);
nor U19990 (N_19990,N_18474,N_18440);
nor U19991 (N_19991,N_18769,N_18436);
or U19992 (N_19992,N_18749,N_18640);
nor U19993 (N_19993,N_18152,N_18495);
or U19994 (N_19994,N_18269,N_18526);
nand U19995 (N_19995,N_18724,N_18452);
and U19996 (N_19996,N_18492,N_18212);
or U19997 (N_19997,N_18719,N_18240);
nor U19998 (N_19998,N_18878,N_18638);
xnor U19999 (N_19999,N_18443,N_18433);
nor U20000 (N_20000,N_19902,N_19919);
nor U20001 (N_20001,N_19948,N_19509);
and U20002 (N_20002,N_19885,N_19558);
nand U20003 (N_20003,N_19114,N_19251);
nand U20004 (N_20004,N_19533,N_19088);
xnor U20005 (N_20005,N_19563,N_19975);
or U20006 (N_20006,N_19889,N_19953);
xnor U20007 (N_20007,N_19551,N_19484);
and U20008 (N_20008,N_19673,N_19606);
or U20009 (N_20009,N_19577,N_19810);
or U20010 (N_20010,N_19772,N_19464);
and U20011 (N_20011,N_19207,N_19575);
xnor U20012 (N_20012,N_19498,N_19694);
and U20013 (N_20013,N_19915,N_19028);
xor U20014 (N_20014,N_19246,N_19029);
xor U20015 (N_20015,N_19908,N_19934);
or U20016 (N_20016,N_19540,N_19706);
nor U20017 (N_20017,N_19235,N_19117);
xnor U20018 (N_20018,N_19593,N_19229);
and U20019 (N_20019,N_19596,N_19044);
or U20020 (N_20020,N_19475,N_19064);
xnor U20021 (N_20021,N_19234,N_19972);
nor U20022 (N_20022,N_19600,N_19869);
or U20023 (N_20023,N_19411,N_19590);
nand U20024 (N_20024,N_19249,N_19984);
nor U20025 (N_20025,N_19944,N_19609);
or U20026 (N_20026,N_19047,N_19657);
nor U20027 (N_20027,N_19298,N_19252);
nand U20028 (N_20028,N_19347,N_19004);
xor U20029 (N_20029,N_19806,N_19959);
nand U20030 (N_20030,N_19069,N_19259);
xnor U20031 (N_20031,N_19928,N_19424);
and U20032 (N_20032,N_19713,N_19541);
xor U20033 (N_20033,N_19999,N_19724);
or U20034 (N_20034,N_19491,N_19794);
xor U20035 (N_20035,N_19880,N_19704);
and U20036 (N_20036,N_19272,N_19050);
nand U20037 (N_20037,N_19082,N_19168);
nor U20038 (N_20038,N_19552,N_19749);
or U20039 (N_20039,N_19032,N_19173);
nand U20040 (N_20040,N_19709,N_19874);
xnor U20041 (N_20041,N_19436,N_19774);
nor U20042 (N_20042,N_19012,N_19583);
or U20043 (N_20043,N_19895,N_19400);
xnor U20044 (N_20044,N_19691,N_19814);
nand U20045 (N_20045,N_19578,N_19568);
nand U20046 (N_20046,N_19977,N_19019);
or U20047 (N_20047,N_19043,N_19375);
nand U20048 (N_20048,N_19800,N_19838);
nand U20049 (N_20049,N_19927,N_19700);
nor U20050 (N_20050,N_19520,N_19398);
xnor U20051 (N_20051,N_19936,N_19039);
nand U20052 (N_20052,N_19397,N_19684);
and U20053 (N_20053,N_19904,N_19042);
and U20054 (N_20054,N_19000,N_19026);
and U20055 (N_20055,N_19282,N_19487);
xnor U20056 (N_20056,N_19320,N_19963);
or U20057 (N_20057,N_19642,N_19284);
or U20058 (N_20058,N_19655,N_19736);
nand U20059 (N_20059,N_19864,N_19137);
xnor U20060 (N_20060,N_19478,N_19631);
xor U20061 (N_20061,N_19792,N_19066);
or U20062 (N_20062,N_19485,N_19231);
and U20063 (N_20063,N_19450,N_19460);
xnor U20064 (N_20064,N_19532,N_19636);
xor U20065 (N_20065,N_19931,N_19516);
nand U20066 (N_20066,N_19356,N_19993);
xor U20067 (N_20067,N_19134,N_19413);
nand U20068 (N_20068,N_19265,N_19214);
nor U20069 (N_20069,N_19494,N_19690);
or U20070 (N_20070,N_19385,N_19926);
nand U20071 (N_20071,N_19705,N_19518);
nor U20072 (N_20072,N_19909,N_19967);
nor U20073 (N_20073,N_19285,N_19729);
and U20074 (N_20074,N_19365,N_19421);
nand U20075 (N_20075,N_19635,N_19095);
xor U20076 (N_20076,N_19799,N_19399);
nand U20077 (N_20077,N_19348,N_19403);
nor U20078 (N_20078,N_19830,N_19712);
or U20079 (N_20079,N_19796,N_19887);
nand U20080 (N_20080,N_19773,N_19942);
nor U20081 (N_20081,N_19198,N_19315);
or U20082 (N_20082,N_19527,N_19384);
or U20083 (N_20083,N_19428,N_19415);
and U20084 (N_20084,N_19689,N_19326);
nand U20085 (N_20085,N_19409,N_19493);
and U20086 (N_20086,N_19731,N_19051);
or U20087 (N_20087,N_19112,N_19130);
nor U20088 (N_20088,N_19359,N_19813);
nor U20089 (N_20089,N_19750,N_19857);
xor U20090 (N_20090,N_19239,N_19727);
xnor U20091 (N_20091,N_19555,N_19101);
or U20092 (N_20092,N_19534,N_19978);
and U20093 (N_20093,N_19495,N_19401);
nor U20094 (N_20094,N_19269,N_19430);
xor U20095 (N_20095,N_19218,N_19544);
nand U20096 (N_20096,N_19276,N_19548);
nor U20097 (N_20097,N_19623,N_19528);
xnor U20098 (N_20098,N_19804,N_19361);
or U20099 (N_20099,N_19063,N_19052);
or U20100 (N_20100,N_19718,N_19273);
nor U20101 (N_20101,N_19539,N_19075);
xor U20102 (N_20102,N_19158,N_19716);
and U20103 (N_20103,N_19938,N_19213);
nand U20104 (N_20104,N_19441,N_19859);
nor U20105 (N_20105,N_19784,N_19679);
and U20106 (N_20106,N_19790,N_19038);
nand U20107 (N_20107,N_19786,N_19416);
and U20108 (N_20108,N_19092,N_19871);
or U20109 (N_20109,N_19512,N_19440);
and U20110 (N_20110,N_19672,N_19654);
nor U20111 (N_20111,N_19087,N_19395);
and U20112 (N_20112,N_19678,N_19858);
nor U20113 (N_20113,N_19763,N_19225);
nand U20114 (N_20114,N_19581,N_19369);
and U20115 (N_20115,N_19305,N_19837);
xor U20116 (N_20116,N_19935,N_19988);
xnor U20117 (N_20117,N_19976,N_19888);
xor U20118 (N_20118,N_19681,N_19007);
or U20119 (N_20119,N_19328,N_19514);
or U20120 (N_20120,N_19970,N_19383);
or U20121 (N_20121,N_19492,N_19200);
nor U20122 (N_20122,N_19671,N_19835);
or U20123 (N_20123,N_19892,N_19956);
nor U20124 (N_20124,N_19536,N_19439);
or U20125 (N_20125,N_19056,N_19426);
or U20126 (N_20126,N_19027,N_19040);
nand U20127 (N_20127,N_19381,N_19876);
xor U20128 (N_20128,N_19852,N_19649);
or U20129 (N_20129,N_19417,N_19291);
or U20130 (N_20130,N_19925,N_19994);
nand U20131 (N_20131,N_19571,N_19856);
or U20132 (N_20132,N_19429,N_19319);
or U20133 (N_20133,N_19390,N_19998);
nand U20134 (N_20134,N_19625,N_19448);
xnor U20135 (N_20135,N_19878,N_19715);
or U20136 (N_20136,N_19989,N_19768);
or U20137 (N_20137,N_19634,N_19839);
or U20138 (N_20138,N_19071,N_19031);
nor U20139 (N_20139,N_19022,N_19181);
nand U20140 (N_20140,N_19849,N_19288);
nor U20141 (N_20141,N_19233,N_19363);
and U20142 (N_20142,N_19331,N_19477);
nand U20143 (N_20143,N_19041,N_19661);
and U20144 (N_20144,N_19990,N_19789);
nor U20145 (N_20145,N_19697,N_19638);
nor U20146 (N_20146,N_19923,N_19821);
nand U20147 (N_20147,N_19180,N_19054);
nor U20148 (N_20148,N_19483,N_19238);
nand U20149 (N_20149,N_19920,N_19129);
and U20150 (N_20150,N_19525,N_19605);
xor U20151 (N_20151,N_19243,N_19145);
nor U20152 (N_20152,N_19542,N_19916);
nor U20153 (N_20153,N_19313,N_19556);
xor U20154 (N_20154,N_19685,N_19738);
nand U20155 (N_20155,N_19201,N_19010);
xor U20156 (N_20156,N_19550,N_19451);
and U20157 (N_20157,N_19209,N_19622);
nand U20158 (N_20158,N_19072,N_19300);
xor U20159 (N_20159,N_19604,N_19135);
nand U20160 (N_20160,N_19437,N_19929);
nand U20161 (N_20161,N_19143,N_19619);
and U20162 (N_20162,N_19912,N_19937);
xnor U20163 (N_20163,N_19947,N_19688);
or U20164 (N_20164,N_19127,N_19023);
or U20165 (N_20165,N_19264,N_19324);
or U20166 (N_20166,N_19643,N_19488);
nor U20167 (N_20167,N_19759,N_19035);
xor U20168 (N_20168,N_19003,N_19997);
or U20169 (N_20169,N_19133,N_19442);
or U20170 (N_20170,N_19569,N_19292);
nand U20171 (N_20171,N_19797,N_19312);
nor U20172 (N_20172,N_19250,N_19378);
and U20173 (N_20173,N_19254,N_19021);
nand U20174 (N_20174,N_19189,N_19817);
nor U20175 (N_20175,N_19553,N_19388);
nor U20176 (N_20176,N_19179,N_19163);
and U20177 (N_20177,N_19677,N_19194);
nand U20178 (N_20178,N_19325,N_19002);
or U20179 (N_20179,N_19462,N_19711);
or U20180 (N_20180,N_19930,N_19220);
nand U20181 (N_20181,N_19662,N_19840);
nand U20182 (N_20182,N_19795,N_19503);
nor U20183 (N_20183,N_19960,N_19873);
or U20184 (N_20184,N_19076,N_19391);
nand U20185 (N_20185,N_19579,N_19248);
xor U20186 (N_20186,N_19376,N_19367);
and U20187 (N_20187,N_19107,N_19819);
xnor U20188 (N_20188,N_19296,N_19455);
and U20189 (N_20189,N_19394,N_19206);
or U20190 (N_20190,N_19756,N_19256);
and U20191 (N_20191,N_19323,N_19008);
and U20192 (N_20192,N_19161,N_19081);
nand U20193 (N_20193,N_19853,N_19422);
or U20194 (N_20194,N_19446,N_19992);
nand U20195 (N_20195,N_19346,N_19393);
nor U20196 (N_20196,N_19106,N_19482);
and U20197 (N_20197,N_19588,N_19263);
nor U20198 (N_20198,N_19221,N_19996);
and U20199 (N_20199,N_19392,N_19500);
and U20200 (N_20200,N_19585,N_19240);
nand U20201 (N_20201,N_19103,N_19974);
xor U20202 (N_20202,N_19809,N_19981);
xor U20203 (N_20203,N_19102,N_19211);
xor U20204 (N_20204,N_19743,N_19203);
xor U20205 (N_20205,N_19150,N_19979);
nor U20206 (N_20206,N_19722,N_19607);
nand U20207 (N_20207,N_19836,N_19077);
nand U20208 (N_20208,N_19434,N_19167);
or U20209 (N_20209,N_19445,N_19486);
nand U20210 (N_20210,N_19834,N_19405);
xor U20211 (N_20211,N_19612,N_19262);
nand U20212 (N_20212,N_19222,N_19005);
nand U20213 (N_20213,N_19624,N_19037);
or U20214 (N_20214,N_19641,N_19782);
nor U20215 (N_20215,N_19844,N_19224);
xnor U20216 (N_20216,N_19253,N_19302);
xor U20217 (N_20217,N_19099,N_19734);
nand U20218 (N_20218,N_19884,N_19699);
or U20219 (N_20219,N_19244,N_19310);
and U20220 (N_20220,N_19097,N_19511);
xor U20221 (N_20221,N_19766,N_19753);
and U20222 (N_20222,N_19109,N_19961);
or U20223 (N_20223,N_19893,N_19538);
or U20224 (N_20224,N_19205,N_19952);
and U20225 (N_20225,N_19785,N_19757);
and U20226 (N_20226,N_19073,N_19223);
or U20227 (N_20227,N_19543,N_19245);
xnor U20228 (N_20228,N_19847,N_19185);
xor U20229 (N_20229,N_19862,N_19215);
nand U20230 (N_20230,N_19781,N_19123);
or U20231 (N_20231,N_19725,N_19720);
xnor U20232 (N_20232,N_19277,N_19197);
nand U20233 (N_20233,N_19057,N_19140);
nand U20234 (N_20234,N_19640,N_19921);
and U20235 (N_20235,N_19687,N_19212);
and U20236 (N_20236,N_19427,N_19666);
and U20237 (N_20237,N_19444,N_19208);
nand U20238 (N_20238,N_19771,N_19062);
nand U20239 (N_20239,N_19693,N_19061);
nor U20240 (N_20240,N_19172,N_19337);
nand U20241 (N_20241,N_19680,N_19025);
and U20242 (N_20242,N_19922,N_19329);
nand U20243 (N_20243,N_19589,N_19560);
nor U20244 (N_20244,N_19184,N_19602);
nor U20245 (N_20245,N_19190,N_19945);
nand U20246 (N_20246,N_19177,N_19803);
nor U20247 (N_20247,N_19456,N_19954);
xor U20248 (N_20248,N_19898,N_19615);
nand U20249 (N_20249,N_19971,N_19675);
and U20250 (N_20250,N_19472,N_19469);
xnor U20251 (N_20251,N_19116,N_19940);
and U20252 (N_20252,N_19522,N_19595);
xor U20253 (N_20253,N_19695,N_19053);
xnor U20254 (N_20254,N_19741,N_19812);
nor U20255 (N_20255,N_19169,N_19121);
xor U20256 (N_20256,N_19196,N_19747);
nor U20257 (N_20257,N_19537,N_19316);
or U20258 (N_20258,N_19610,N_19386);
nand U20259 (N_20259,N_19780,N_19255);
xnor U20260 (N_20260,N_19015,N_19648);
xor U20261 (N_20261,N_19351,N_19119);
and U20262 (N_20262,N_19170,N_19174);
xor U20263 (N_20263,N_19530,N_19358);
and U20264 (N_20264,N_19350,N_19601);
xnor U20265 (N_20265,N_19890,N_19149);
xor U20266 (N_20266,N_19085,N_19122);
or U20267 (N_20267,N_19549,N_19059);
xor U20268 (N_20268,N_19461,N_19124);
and U20269 (N_20269,N_19823,N_19968);
nand U20270 (N_20270,N_19899,N_19281);
nand U20271 (N_20271,N_19219,N_19710);
nor U20272 (N_20272,N_19188,N_19176);
nor U20273 (N_20273,N_19089,N_19973);
nand U20274 (N_20274,N_19828,N_19090);
nand U20275 (N_20275,N_19354,N_19497);
nand U20276 (N_20276,N_19848,N_19656);
or U20277 (N_20277,N_19321,N_19438);
nor U20278 (N_20278,N_19913,N_19567);
nor U20279 (N_20279,N_19807,N_19311);
or U20280 (N_20280,N_19764,N_19815);
or U20281 (N_20281,N_19271,N_19125);
and U20282 (N_20282,N_19418,N_19557);
or U20283 (N_20283,N_19192,N_19258);
and U20284 (N_20284,N_19805,N_19524);
nand U20285 (N_20285,N_19676,N_19816);
xor U20286 (N_20286,N_19113,N_19084);
or U20287 (N_20287,N_19660,N_19138);
and U20288 (N_20288,N_19286,N_19098);
xor U20289 (N_20289,N_19307,N_19481);
nor U20290 (N_20290,N_19074,N_19746);
and U20291 (N_20291,N_19969,N_19613);
and U20292 (N_20292,N_19686,N_19868);
or U20293 (N_20293,N_19330,N_19778);
xnor U20294 (N_20294,N_19572,N_19132);
or U20295 (N_20295,N_19187,N_19030);
xnor U20296 (N_20296,N_19658,N_19183);
and U20297 (N_20297,N_19983,N_19299);
xnor U20298 (N_20298,N_19476,N_19006);
nand U20299 (N_20299,N_19001,N_19637);
and U20300 (N_20300,N_19410,N_19779);
xnor U20301 (N_20301,N_19278,N_19824);
nand U20302 (N_20302,N_19279,N_19408);
or U20303 (N_20303,N_19344,N_19745);
or U20304 (N_20304,N_19216,N_19850);
nand U20305 (N_20305,N_19142,N_19698);
xnor U20306 (N_20306,N_19570,N_19626);
xnor U20307 (N_20307,N_19452,N_19742);
xor U20308 (N_20308,N_19034,N_19651);
nor U20309 (N_20309,N_19268,N_19371);
xnor U20310 (N_20310,N_19515,N_19217);
or U20311 (N_20311,N_19175,N_19941);
or U20312 (N_20312,N_19151,N_19573);
nand U20313 (N_20313,N_19517,N_19078);
nor U20314 (N_20314,N_19080,N_19751);
xnor U20315 (N_20315,N_19147,N_19650);
nand U20316 (N_20316,N_19295,N_19160);
and U20317 (N_20317,N_19368,N_19389);
nor U20318 (N_20318,N_19357,N_19707);
or U20319 (N_20319,N_19431,N_19237);
or U20320 (N_20320,N_19236,N_19526);
xor U20321 (N_20321,N_19752,N_19165);
or U20322 (N_20322,N_19854,N_19886);
nor U20323 (N_20323,N_19918,N_19270);
nand U20324 (N_20324,N_19621,N_19104);
and U20325 (N_20325,N_19760,N_19280);
and U20326 (N_20326,N_19939,N_19740);
nor U20327 (N_20327,N_19274,N_19701);
and U20328 (N_20328,N_19195,N_19349);
nor U20329 (N_20329,N_19507,N_19414);
and U20330 (N_20330,N_19545,N_19566);
or U20331 (N_20331,N_19728,N_19499);
nor U20332 (N_20332,N_19755,N_19591);
nor U20333 (N_20333,N_19412,N_19338);
xor U20334 (N_20334,N_19714,N_19985);
and U20335 (N_20335,N_19597,N_19370);
or U20336 (N_20336,N_19667,N_19110);
nor U20337 (N_20337,N_19907,N_19881);
xnor U20338 (N_20338,N_19721,N_19297);
nor U20339 (N_20339,N_19341,N_19633);
or U20340 (N_20340,N_19776,N_19046);
or U20341 (N_20341,N_19407,N_19793);
xor U20342 (N_20342,N_19843,N_19293);
nor U20343 (N_20343,N_19060,N_19128);
and U20344 (N_20344,N_19618,N_19501);
nor U20345 (N_20345,N_19458,N_19290);
or U20346 (N_20346,N_19906,N_19199);
and U20347 (N_20347,N_19327,N_19423);
nand U20348 (N_20348,N_19171,N_19565);
and U20349 (N_20349,N_19334,N_19962);
or U20350 (N_20350,N_19943,N_19480);
nor U20351 (N_20351,N_19362,N_19382);
and U20352 (N_20352,N_19105,N_19574);
xor U20353 (N_20353,N_19958,N_19627);
xor U20354 (N_20354,N_19049,N_19846);
and U20355 (N_20355,N_19732,N_19283);
and U20356 (N_20356,N_19340,N_19991);
xor U20357 (N_20357,N_19901,N_19467);
xor U20358 (N_20358,N_19966,N_19360);
xor U20359 (N_20359,N_19965,N_19617);
xor U20360 (N_20360,N_19825,N_19865);
nor U20361 (N_20361,N_19374,N_19014);
nand U20362 (N_20362,N_19910,N_19559);
nor U20363 (N_20363,N_19950,N_19466);
xnor U20364 (N_20364,N_19519,N_19096);
or U20365 (N_20365,N_19986,N_19562);
nand U20366 (N_20366,N_19833,N_19287);
nand U20367 (N_20367,N_19178,N_19425);
and U20368 (N_20368,N_19093,N_19111);
or U20369 (N_20369,N_19683,N_19758);
or U20370 (N_20370,N_19739,N_19159);
nor U20371 (N_20371,N_19582,N_19141);
and U20372 (N_20372,N_19336,N_19332);
nor U20373 (N_20373,N_19335,N_19146);
or U20374 (N_20374,N_19860,N_19402);
or U20375 (N_20375,N_19017,N_19406);
xnor U20376 (N_20376,N_19659,N_19896);
nand U20377 (N_20377,N_19016,N_19584);
xnor U20378 (N_20378,N_19308,N_19447);
or U20379 (N_20379,N_19762,N_19156);
and U20380 (N_20380,N_19911,N_19013);
and U20381 (N_20381,N_19343,N_19465);
or U20382 (N_20382,N_19879,N_19730);
nand U20383 (N_20383,N_19304,N_19802);
and U20384 (N_20384,N_19645,N_19045);
and U20385 (N_20385,N_19702,N_19261);
xnor U20386 (N_20386,N_19506,N_19523);
and U20387 (N_20387,N_19420,N_19663);
xor U20388 (N_20388,N_19614,N_19067);
xnor U20389 (N_20389,N_19933,N_19761);
xor U20390 (N_20390,N_19957,N_19257);
and U20391 (N_20391,N_19513,N_19342);
nor U20392 (N_20392,N_19470,N_19692);
nor U20393 (N_20393,N_19301,N_19275);
nand U20394 (N_20394,N_19419,N_19668);
nand U20395 (N_20395,N_19831,N_19387);
nor U20396 (N_20396,N_19033,N_19289);
xor U20397 (N_20397,N_19191,N_19317);
xnor U20398 (N_20398,N_19586,N_19818);
xnor U20399 (N_20399,N_19576,N_19696);
xnor U20400 (N_20400,N_19787,N_19309);
and U20401 (N_20401,N_19894,N_19510);
nand U20402 (N_20402,N_19496,N_19083);
xor U20403 (N_20403,N_19877,N_19435);
nand U20404 (N_20404,N_19791,N_19079);
or U20405 (N_20405,N_19166,N_19202);
nor U20406 (N_20406,N_19164,N_19230);
and U20407 (N_20407,N_19318,N_19474);
or U20408 (N_20408,N_19726,N_19647);
xor U20409 (N_20409,N_19744,N_19210);
xor U20410 (N_20410,N_19842,N_19748);
xor U20411 (N_20411,N_19628,N_19162);
and U20412 (N_20412,N_19100,N_19580);
or U20413 (N_20413,N_19951,N_19903);
or U20414 (N_20414,N_19872,N_19153);
nand U20415 (N_20415,N_19775,N_19306);
nand U20416 (N_20416,N_19155,N_19674);
nor U20417 (N_20417,N_19242,N_19788);
nand U20418 (N_20418,N_19036,N_19154);
nand U20419 (N_20419,N_19769,N_19851);
nor U20420 (N_20420,N_19598,N_19120);
nand U20421 (N_20421,N_19379,N_19737);
nor U20422 (N_20422,N_19531,N_19345);
nand U20423 (N_20423,N_19068,N_19443);
nand U20424 (N_20424,N_19396,N_19870);
nand U20425 (N_20425,N_19353,N_19490);
or U20426 (N_20426,N_19995,N_19294);
nor U20427 (N_20427,N_19653,N_19152);
nand U20428 (N_20428,N_19629,N_19682);
and U20429 (N_20429,N_19867,N_19204);
nor U20430 (N_20430,N_19664,N_19070);
or U20431 (N_20431,N_19646,N_19917);
xor U20432 (N_20432,N_19144,N_19065);
nor U20433 (N_20433,N_19822,N_19665);
or U20434 (N_20434,N_19827,N_19863);
or U20435 (N_20435,N_19267,N_19987);
and U20436 (N_20436,N_19599,N_19955);
nand U20437 (N_20437,N_19266,N_19980);
nor U20438 (N_20438,N_19489,N_19770);
nor U20439 (N_20439,N_19020,N_19433);
nor U20440 (N_20440,N_19946,N_19454);
and U20441 (N_20441,N_19767,N_19964);
nor U20442 (N_20442,N_19058,N_19808);
or U20443 (N_20443,N_19639,N_19048);
nor U20444 (N_20444,N_19882,N_19502);
or U20445 (N_20445,N_19457,N_19468);
xnor U20446 (N_20446,N_19949,N_19554);
nor U20447 (N_20447,N_19463,N_19086);
and U20448 (N_20448,N_19193,N_19723);
nor U20449 (N_20449,N_19018,N_19644);
nand U20450 (N_20450,N_19924,N_19735);
or U20451 (N_20451,N_19670,N_19829);
xor U20452 (N_20452,N_19024,N_19459);
or U20453 (N_20453,N_19449,N_19333);
nand U20454 (N_20454,N_19131,N_19303);
xor U20455 (N_20455,N_19364,N_19733);
xnor U20456 (N_20456,N_19473,N_19508);
nand U20457 (N_20457,N_19226,N_19479);
or U20458 (N_20458,N_19564,N_19900);
nor U20459 (N_20459,N_19982,N_19355);
or U20460 (N_20460,N_19841,N_19754);
and U20461 (N_20461,N_19546,N_19826);
or U20462 (N_20462,N_19432,N_19811);
nand U20463 (N_20463,N_19875,N_19866);
xnor U20464 (N_20464,N_19832,N_19703);
nand U20465 (N_20465,N_19009,N_19228);
and U20466 (N_20466,N_19157,N_19380);
and U20467 (N_20467,N_19801,N_19783);
nand U20468 (N_20468,N_19453,N_19247);
and U20469 (N_20469,N_19765,N_19905);
xor U20470 (N_20470,N_19504,N_19352);
or U20471 (N_20471,N_19529,N_19535);
or U20472 (N_20472,N_19373,N_19719);
nand U20473 (N_20473,N_19611,N_19108);
nand U20474 (N_20474,N_19861,N_19055);
and U20475 (N_20475,N_19182,N_19136);
nor U20476 (N_20476,N_19669,N_19708);
xor U20477 (N_20477,N_19186,N_19616);
nand U20478 (N_20478,N_19115,N_19471);
or U20479 (N_20479,N_19404,N_19314);
or U20480 (N_20480,N_19630,N_19322);
and U20481 (N_20481,N_19547,N_19652);
or U20482 (N_20482,N_19632,N_19118);
xnor U20483 (N_20483,N_19592,N_19620);
nor U20484 (N_20484,N_19521,N_19227);
nand U20485 (N_20485,N_19148,N_19603);
and U20486 (N_20486,N_19505,N_19897);
nand U20487 (N_20487,N_19717,N_19366);
nor U20488 (N_20488,N_19377,N_19241);
xor U20489 (N_20489,N_19091,N_19587);
and U20490 (N_20490,N_19126,N_19798);
and U20491 (N_20491,N_19339,N_19608);
or U20492 (N_20492,N_19561,N_19845);
nor U20493 (N_20493,N_19139,N_19883);
xor U20494 (N_20494,N_19932,N_19232);
or U20495 (N_20495,N_19372,N_19914);
nor U20496 (N_20496,N_19820,N_19094);
xnor U20497 (N_20497,N_19594,N_19855);
or U20498 (N_20498,N_19891,N_19260);
xnor U20499 (N_20499,N_19777,N_19011);
and U20500 (N_20500,N_19663,N_19271);
and U20501 (N_20501,N_19813,N_19939);
nand U20502 (N_20502,N_19972,N_19527);
nor U20503 (N_20503,N_19143,N_19612);
nand U20504 (N_20504,N_19497,N_19752);
xnor U20505 (N_20505,N_19245,N_19063);
or U20506 (N_20506,N_19478,N_19332);
or U20507 (N_20507,N_19783,N_19718);
and U20508 (N_20508,N_19453,N_19082);
nand U20509 (N_20509,N_19478,N_19255);
or U20510 (N_20510,N_19483,N_19497);
nor U20511 (N_20511,N_19952,N_19957);
nor U20512 (N_20512,N_19354,N_19200);
nor U20513 (N_20513,N_19111,N_19470);
nand U20514 (N_20514,N_19742,N_19578);
xor U20515 (N_20515,N_19955,N_19077);
and U20516 (N_20516,N_19548,N_19797);
nand U20517 (N_20517,N_19610,N_19500);
and U20518 (N_20518,N_19024,N_19455);
or U20519 (N_20519,N_19469,N_19924);
nor U20520 (N_20520,N_19365,N_19284);
nand U20521 (N_20521,N_19446,N_19157);
xor U20522 (N_20522,N_19825,N_19010);
and U20523 (N_20523,N_19249,N_19999);
nor U20524 (N_20524,N_19062,N_19146);
nand U20525 (N_20525,N_19558,N_19701);
or U20526 (N_20526,N_19927,N_19838);
xnor U20527 (N_20527,N_19048,N_19719);
or U20528 (N_20528,N_19483,N_19461);
or U20529 (N_20529,N_19167,N_19046);
or U20530 (N_20530,N_19477,N_19564);
nand U20531 (N_20531,N_19592,N_19868);
and U20532 (N_20532,N_19855,N_19153);
nand U20533 (N_20533,N_19763,N_19915);
nand U20534 (N_20534,N_19447,N_19178);
and U20535 (N_20535,N_19582,N_19970);
or U20536 (N_20536,N_19057,N_19485);
xnor U20537 (N_20537,N_19737,N_19644);
nand U20538 (N_20538,N_19931,N_19596);
or U20539 (N_20539,N_19182,N_19364);
or U20540 (N_20540,N_19267,N_19337);
nand U20541 (N_20541,N_19727,N_19110);
or U20542 (N_20542,N_19515,N_19791);
and U20543 (N_20543,N_19309,N_19221);
and U20544 (N_20544,N_19170,N_19266);
or U20545 (N_20545,N_19764,N_19715);
and U20546 (N_20546,N_19273,N_19359);
xnor U20547 (N_20547,N_19832,N_19108);
nor U20548 (N_20548,N_19305,N_19166);
or U20549 (N_20549,N_19250,N_19247);
nand U20550 (N_20550,N_19633,N_19598);
or U20551 (N_20551,N_19420,N_19297);
and U20552 (N_20552,N_19150,N_19832);
and U20553 (N_20553,N_19218,N_19750);
xor U20554 (N_20554,N_19700,N_19163);
nor U20555 (N_20555,N_19072,N_19670);
or U20556 (N_20556,N_19207,N_19981);
and U20557 (N_20557,N_19622,N_19427);
nor U20558 (N_20558,N_19244,N_19995);
xnor U20559 (N_20559,N_19997,N_19201);
nand U20560 (N_20560,N_19819,N_19215);
xor U20561 (N_20561,N_19504,N_19766);
nor U20562 (N_20562,N_19986,N_19672);
or U20563 (N_20563,N_19976,N_19521);
xor U20564 (N_20564,N_19427,N_19974);
nor U20565 (N_20565,N_19399,N_19689);
and U20566 (N_20566,N_19619,N_19547);
or U20567 (N_20567,N_19958,N_19699);
or U20568 (N_20568,N_19039,N_19899);
nand U20569 (N_20569,N_19353,N_19406);
and U20570 (N_20570,N_19293,N_19370);
xnor U20571 (N_20571,N_19495,N_19193);
xor U20572 (N_20572,N_19560,N_19617);
nor U20573 (N_20573,N_19388,N_19590);
nor U20574 (N_20574,N_19821,N_19559);
nor U20575 (N_20575,N_19760,N_19290);
nand U20576 (N_20576,N_19924,N_19789);
nand U20577 (N_20577,N_19537,N_19207);
nand U20578 (N_20578,N_19086,N_19816);
or U20579 (N_20579,N_19376,N_19054);
and U20580 (N_20580,N_19911,N_19527);
and U20581 (N_20581,N_19427,N_19265);
or U20582 (N_20582,N_19036,N_19904);
nor U20583 (N_20583,N_19744,N_19592);
or U20584 (N_20584,N_19005,N_19353);
nand U20585 (N_20585,N_19858,N_19232);
or U20586 (N_20586,N_19243,N_19234);
and U20587 (N_20587,N_19845,N_19182);
nor U20588 (N_20588,N_19576,N_19607);
and U20589 (N_20589,N_19595,N_19401);
nand U20590 (N_20590,N_19979,N_19953);
nand U20591 (N_20591,N_19557,N_19779);
and U20592 (N_20592,N_19356,N_19849);
xor U20593 (N_20593,N_19029,N_19358);
and U20594 (N_20594,N_19433,N_19939);
nand U20595 (N_20595,N_19332,N_19050);
nand U20596 (N_20596,N_19300,N_19690);
or U20597 (N_20597,N_19503,N_19701);
and U20598 (N_20598,N_19323,N_19626);
xor U20599 (N_20599,N_19975,N_19655);
or U20600 (N_20600,N_19767,N_19922);
xor U20601 (N_20601,N_19743,N_19543);
nand U20602 (N_20602,N_19645,N_19760);
xor U20603 (N_20603,N_19844,N_19208);
nor U20604 (N_20604,N_19101,N_19604);
and U20605 (N_20605,N_19056,N_19555);
xor U20606 (N_20606,N_19037,N_19350);
nor U20607 (N_20607,N_19361,N_19322);
nor U20608 (N_20608,N_19695,N_19321);
or U20609 (N_20609,N_19124,N_19528);
nand U20610 (N_20610,N_19665,N_19352);
or U20611 (N_20611,N_19377,N_19042);
and U20612 (N_20612,N_19337,N_19598);
nor U20613 (N_20613,N_19152,N_19899);
or U20614 (N_20614,N_19771,N_19354);
nor U20615 (N_20615,N_19164,N_19807);
xor U20616 (N_20616,N_19344,N_19920);
xnor U20617 (N_20617,N_19308,N_19835);
or U20618 (N_20618,N_19574,N_19112);
nand U20619 (N_20619,N_19929,N_19974);
xnor U20620 (N_20620,N_19074,N_19169);
and U20621 (N_20621,N_19424,N_19387);
or U20622 (N_20622,N_19366,N_19092);
or U20623 (N_20623,N_19582,N_19061);
xor U20624 (N_20624,N_19788,N_19409);
or U20625 (N_20625,N_19964,N_19400);
nand U20626 (N_20626,N_19778,N_19602);
and U20627 (N_20627,N_19598,N_19874);
nand U20628 (N_20628,N_19665,N_19449);
and U20629 (N_20629,N_19075,N_19293);
nor U20630 (N_20630,N_19442,N_19335);
xor U20631 (N_20631,N_19891,N_19964);
and U20632 (N_20632,N_19497,N_19798);
and U20633 (N_20633,N_19237,N_19822);
or U20634 (N_20634,N_19116,N_19054);
and U20635 (N_20635,N_19112,N_19957);
or U20636 (N_20636,N_19029,N_19389);
and U20637 (N_20637,N_19562,N_19699);
or U20638 (N_20638,N_19046,N_19710);
nand U20639 (N_20639,N_19208,N_19210);
or U20640 (N_20640,N_19927,N_19934);
nor U20641 (N_20641,N_19961,N_19200);
or U20642 (N_20642,N_19044,N_19156);
nand U20643 (N_20643,N_19039,N_19811);
nand U20644 (N_20644,N_19448,N_19319);
nor U20645 (N_20645,N_19528,N_19194);
nand U20646 (N_20646,N_19132,N_19419);
nand U20647 (N_20647,N_19845,N_19675);
xnor U20648 (N_20648,N_19244,N_19069);
and U20649 (N_20649,N_19338,N_19837);
or U20650 (N_20650,N_19862,N_19503);
nand U20651 (N_20651,N_19696,N_19945);
or U20652 (N_20652,N_19989,N_19642);
or U20653 (N_20653,N_19936,N_19494);
nand U20654 (N_20654,N_19163,N_19934);
nor U20655 (N_20655,N_19328,N_19446);
xor U20656 (N_20656,N_19229,N_19785);
nand U20657 (N_20657,N_19214,N_19992);
nand U20658 (N_20658,N_19650,N_19516);
or U20659 (N_20659,N_19234,N_19421);
xnor U20660 (N_20660,N_19285,N_19160);
nand U20661 (N_20661,N_19887,N_19398);
and U20662 (N_20662,N_19739,N_19705);
xor U20663 (N_20663,N_19708,N_19739);
xnor U20664 (N_20664,N_19905,N_19291);
nor U20665 (N_20665,N_19776,N_19622);
xor U20666 (N_20666,N_19978,N_19259);
and U20667 (N_20667,N_19971,N_19804);
nand U20668 (N_20668,N_19924,N_19292);
or U20669 (N_20669,N_19836,N_19493);
and U20670 (N_20670,N_19211,N_19642);
nor U20671 (N_20671,N_19546,N_19973);
and U20672 (N_20672,N_19332,N_19326);
and U20673 (N_20673,N_19279,N_19036);
and U20674 (N_20674,N_19670,N_19799);
and U20675 (N_20675,N_19064,N_19177);
nor U20676 (N_20676,N_19042,N_19341);
nand U20677 (N_20677,N_19474,N_19011);
or U20678 (N_20678,N_19111,N_19635);
xnor U20679 (N_20679,N_19923,N_19640);
nor U20680 (N_20680,N_19984,N_19472);
nor U20681 (N_20681,N_19274,N_19277);
and U20682 (N_20682,N_19057,N_19294);
xnor U20683 (N_20683,N_19022,N_19219);
xnor U20684 (N_20684,N_19856,N_19695);
or U20685 (N_20685,N_19509,N_19850);
and U20686 (N_20686,N_19667,N_19485);
nor U20687 (N_20687,N_19746,N_19642);
or U20688 (N_20688,N_19639,N_19858);
or U20689 (N_20689,N_19736,N_19249);
or U20690 (N_20690,N_19307,N_19653);
nand U20691 (N_20691,N_19833,N_19968);
nand U20692 (N_20692,N_19653,N_19922);
nand U20693 (N_20693,N_19254,N_19940);
nand U20694 (N_20694,N_19507,N_19708);
and U20695 (N_20695,N_19833,N_19863);
nand U20696 (N_20696,N_19100,N_19428);
or U20697 (N_20697,N_19407,N_19638);
nand U20698 (N_20698,N_19723,N_19468);
nand U20699 (N_20699,N_19127,N_19700);
xor U20700 (N_20700,N_19168,N_19327);
xnor U20701 (N_20701,N_19062,N_19044);
nor U20702 (N_20702,N_19722,N_19293);
or U20703 (N_20703,N_19870,N_19569);
and U20704 (N_20704,N_19804,N_19653);
and U20705 (N_20705,N_19769,N_19775);
or U20706 (N_20706,N_19019,N_19618);
xnor U20707 (N_20707,N_19938,N_19059);
or U20708 (N_20708,N_19565,N_19205);
nor U20709 (N_20709,N_19868,N_19217);
nor U20710 (N_20710,N_19140,N_19776);
nand U20711 (N_20711,N_19826,N_19155);
or U20712 (N_20712,N_19389,N_19645);
or U20713 (N_20713,N_19879,N_19281);
nor U20714 (N_20714,N_19000,N_19896);
xnor U20715 (N_20715,N_19071,N_19455);
xor U20716 (N_20716,N_19020,N_19671);
nand U20717 (N_20717,N_19200,N_19254);
and U20718 (N_20718,N_19417,N_19534);
nand U20719 (N_20719,N_19440,N_19812);
xor U20720 (N_20720,N_19774,N_19352);
nand U20721 (N_20721,N_19398,N_19281);
and U20722 (N_20722,N_19151,N_19595);
nand U20723 (N_20723,N_19544,N_19098);
nor U20724 (N_20724,N_19215,N_19421);
or U20725 (N_20725,N_19236,N_19706);
or U20726 (N_20726,N_19923,N_19636);
nor U20727 (N_20727,N_19449,N_19332);
nand U20728 (N_20728,N_19689,N_19783);
nor U20729 (N_20729,N_19679,N_19625);
xnor U20730 (N_20730,N_19045,N_19845);
nand U20731 (N_20731,N_19042,N_19393);
nand U20732 (N_20732,N_19078,N_19280);
nor U20733 (N_20733,N_19620,N_19634);
nand U20734 (N_20734,N_19476,N_19496);
or U20735 (N_20735,N_19251,N_19683);
nand U20736 (N_20736,N_19311,N_19257);
or U20737 (N_20737,N_19629,N_19026);
and U20738 (N_20738,N_19435,N_19621);
nand U20739 (N_20739,N_19360,N_19535);
nand U20740 (N_20740,N_19445,N_19384);
xor U20741 (N_20741,N_19939,N_19129);
and U20742 (N_20742,N_19253,N_19937);
or U20743 (N_20743,N_19526,N_19106);
and U20744 (N_20744,N_19658,N_19198);
nor U20745 (N_20745,N_19582,N_19553);
nand U20746 (N_20746,N_19804,N_19282);
nand U20747 (N_20747,N_19131,N_19980);
xor U20748 (N_20748,N_19247,N_19551);
nor U20749 (N_20749,N_19579,N_19627);
nor U20750 (N_20750,N_19537,N_19139);
and U20751 (N_20751,N_19483,N_19903);
nor U20752 (N_20752,N_19879,N_19590);
xnor U20753 (N_20753,N_19437,N_19165);
or U20754 (N_20754,N_19623,N_19606);
or U20755 (N_20755,N_19271,N_19703);
nor U20756 (N_20756,N_19262,N_19030);
or U20757 (N_20757,N_19698,N_19565);
or U20758 (N_20758,N_19471,N_19671);
and U20759 (N_20759,N_19936,N_19422);
xor U20760 (N_20760,N_19403,N_19743);
xnor U20761 (N_20761,N_19684,N_19621);
nand U20762 (N_20762,N_19758,N_19334);
nand U20763 (N_20763,N_19118,N_19305);
nor U20764 (N_20764,N_19480,N_19860);
and U20765 (N_20765,N_19835,N_19254);
nor U20766 (N_20766,N_19266,N_19735);
and U20767 (N_20767,N_19842,N_19693);
and U20768 (N_20768,N_19820,N_19447);
or U20769 (N_20769,N_19816,N_19052);
or U20770 (N_20770,N_19136,N_19749);
or U20771 (N_20771,N_19148,N_19528);
and U20772 (N_20772,N_19380,N_19459);
or U20773 (N_20773,N_19036,N_19685);
xnor U20774 (N_20774,N_19837,N_19919);
nand U20775 (N_20775,N_19147,N_19231);
or U20776 (N_20776,N_19363,N_19254);
nor U20777 (N_20777,N_19879,N_19689);
or U20778 (N_20778,N_19270,N_19729);
nand U20779 (N_20779,N_19125,N_19472);
nand U20780 (N_20780,N_19133,N_19298);
and U20781 (N_20781,N_19491,N_19533);
or U20782 (N_20782,N_19940,N_19054);
xnor U20783 (N_20783,N_19720,N_19640);
xor U20784 (N_20784,N_19636,N_19075);
or U20785 (N_20785,N_19747,N_19154);
nand U20786 (N_20786,N_19677,N_19039);
nand U20787 (N_20787,N_19276,N_19319);
and U20788 (N_20788,N_19899,N_19096);
xnor U20789 (N_20789,N_19724,N_19367);
nor U20790 (N_20790,N_19831,N_19058);
nand U20791 (N_20791,N_19028,N_19688);
or U20792 (N_20792,N_19850,N_19262);
nor U20793 (N_20793,N_19504,N_19039);
nand U20794 (N_20794,N_19868,N_19645);
nand U20795 (N_20795,N_19296,N_19551);
xnor U20796 (N_20796,N_19464,N_19785);
or U20797 (N_20797,N_19712,N_19026);
and U20798 (N_20798,N_19556,N_19101);
or U20799 (N_20799,N_19889,N_19522);
or U20800 (N_20800,N_19200,N_19926);
or U20801 (N_20801,N_19044,N_19245);
or U20802 (N_20802,N_19497,N_19321);
or U20803 (N_20803,N_19612,N_19847);
nor U20804 (N_20804,N_19107,N_19604);
and U20805 (N_20805,N_19347,N_19392);
nand U20806 (N_20806,N_19219,N_19777);
and U20807 (N_20807,N_19607,N_19410);
or U20808 (N_20808,N_19571,N_19699);
xnor U20809 (N_20809,N_19569,N_19196);
nor U20810 (N_20810,N_19043,N_19252);
or U20811 (N_20811,N_19325,N_19941);
nand U20812 (N_20812,N_19137,N_19190);
and U20813 (N_20813,N_19045,N_19925);
nor U20814 (N_20814,N_19397,N_19301);
and U20815 (N_20815,N_19091,N_19626);
nand U20816 (N_20816,N_19202,N_19076);
nand U20817 (N_20817,N_19097,N_19124);
nor U20818 (N_20818,N_19412,N_19280);
or U20819 (N_20819,N_19718,N_19954);
nor U20820 (N_20820,N_19574,N_19294);
nor U20821 (N_20821,N_19058,N_19684);
or U20822 (N_20822,N_19991,N_19568);
and U20823 (N_20823,N_19817,N_19103);
or U20824 (N_20824,N_19832,N_19921);
xnor U20825 (N_20825,N_19113,N_19671);
and U20826 (N_20826,N_19623,N_19544);
xnor U20827 (N_20827,N_19317,N_19734);
nor U20828 (N_20828,N_19984,N_19089);
nor U20829 (N_20829,N_19189,N_19529);
nand U20830 (N_20830,N_19776,N_19637);
nor U20831 (N_20831,N_19977,N_19751);
and U20832 (N_20832,N_19927,N_19170);
or U20833 (N_20833,N_19137,N_19992);
nand U20834 (N_20834,N_19089,N_19150);
nor U20835 (N_20835,N_19975,N_19990);
nor U20836 (N_20836,N_19164,N_19540);
and U20837 (N_20837,N_19173,N_19738);
nor U20838 (N_20838,N_19693,N_19001);
xor U20839 (N_20839,N_19419,N_19313);
nand U20840 (N_20840,N_19676,N_19197);
or U20841 (N_20841,N_19358,N_19751);
xnor U20842 (N_20842,N_19842,N_19286);
xnor U20843 (N_20843,N_19720,N_19321);
nand U20844 (N_20844,N_19530,N_19591);
or U20845 (N_20845,N_19210,N_19811);
xor U20846 (N_20846,N_19269,N_19786);
xnor U20847 (N_20847,N_19555,N_19834);
and U20848 (N_20848,N_19485,N_19968);
nor U20849 (N_20849,N_19216,N_19383);
nand U20850 (N_20850,N_19252,N_19358);
xnor U20851 (N_20851,N_19868,N_19041);
nor U20852 (N_20852,N_19946,N_19049);
and U20853 (N_20853,N_19984,N_19242);
xor U20854 (N_20854,N_19995,N_19070);
nor U20855 (N_20855,N_19780,N_19515);
or U20856 (N_20856,N_19731,N_19028);
xor U20857 (N_20857,N_19881,N_19979);
or U20858 (N_20858,N_19218,N_19242);
nor U20859 (N_20859,N_19020,N_19244);
nor U20860 (N_20860,N_19554,N_19139);
xnor U20861 (N_20861,N_19882,N_19006);
xnor U20862 (N_20862,N_19108,N_19939);
and U20863 (N_20863,N_19202,N_19043);
or U20864 (N_20864,N_19187,N_19344);
nand U20865 (N_20865,N_19326,N_19296);
and U20866 (N_20866,N_19023,N_19478);
xor U20867 (N_20867,N_19137,N_19881);
and U20868 (N_20868,N_19032,N_19551);
nor U20869 (N_20869,N_19338,N_19354);
xnor U20870 (N_20870,N_19769,N_19398);
xor U20871 (N_20871,N_19741,N_19759);
xnor U20872 (N_20872,N_19465,N_19315);
nand U20873 (N_20873,N_19396,N_19527);
nand U20874 (N_20874,N_19775,N_19620);
xor U20875 (N_20875,N_19236,N_19452);
and U20876 (N_20876,N_19690,N_19393);
nand U20877 (N_20877,N_19672,N_19295);
nand U20878 (N_20878,N_19963,N_19816);
or U20879 (N_20879,N_19943,N_19434);
or U20880 (N_20880,N_19313,N_19056);
nand U20881 (N_20881,N_19356,N_19643);
nor U20882 (N_20882,N_19207,N_19189);
nand U20883 (N_20883,N_19547,N_19822);
or U20884 (N_20884,N_19425,N_19017);
nand U20885 (N_20885,N_19809,N_19336);
and U20886 (N_20886,N_19158,N_19628);
nand U20887 (N_20887,N_19122,N_19356);
nand U20888 (N_20888,N_19217,N_19062);
and U20889 (N_20889,N_19692,N_19754);
and U20890 (N_20890,N_19190,N_19628);
xor U20891 (N_20891,N_19353,N_19412);
xnor U20892 (N_20892,N_19706,N_19747);
and U20893 (N_20893,N_19132,N_19251);
or U20894 (N_20894,N_19866,N_19499);
xor U20895 (N_20895,N_19087,N_19250);
nand U20896 (N_20896,N_19219,N_19198);
xor U20897 (N_20897,N_19536,N_19326);
nor U20898 (N_20898,N_19585,N_19830);
xor U20899 (N_20899,N_19820,N_19837);
nor U20900 (N_20900,N_19957,N_19735);
and U20901 (N_20901,N_19456,N_19148);
xnor U20902 (N_20902,N_19514,N_19143);
or U20903 (N_20903,N_19590,N_19156);
xnor U20904 (N_20904,N_19346,N_19720);
or U20905 (N_20905,N_19225,N_19811);
nor U20906 (N_20906,N_19660,N_19888);
xor U20907 (N_20907,N_19308,N_19380);
and U20908 (N_20908,N_19592,N_19613);
and U20909 (N_20909,N_19251,N_19239);
or U20910 (N_20910,N_19508,N_19299);
xnor U20911 (N_20911,N_19786,N_19056);
nand U20912 (N_20912,N_19223,N_19548);
nand U20913 (N_20913,N_19400,N_19659);
nor U20914 (N_20914,N_19373,N_19411);
xor U20915 (N_20915,N_19113,N_19476);
and U20916 (N_20916,N_19518,N_19710);
nor U20917 (N_20917,N_19309,N_19770);
or U20918 (N_20918,N_19333,N_19356);
or U20919 (N_20919,N_19993,N_19994);
or U20920 (N_20920,N_19999,N_19663);
nand U20921 (N_20921,N_19018,N_19967);
nand U20922 (N_20922,N_19829,N_19590);
or U20923 (N_20923,N_19003,N_19234);
nand U20924 (N_20924,N_19329,N_19802);
or U20925 (N_20925,N_19160,N_19904);
and U20926 (N_20926,N_19814,N_19338);
and U20927 (N_20927,N_19999,N_19177);
or U20928 (N_20928,N_19475,N_19730);
nor U20929 (N_20929,N_19620,N_19088);
or U20930 (N_20930,N_19738,N_19813);
or U20931 (N_20931,N_19293,N_19766);
nor U20932 (N_20932,N_19751,N_19826);
nor U20933 (N_20933,N_19604,N_19383);
xnor U20934 (N_20934,N_19704,N_19424);
nand U20935 (N_20935,N_19473,N_19157);
nand U20936 (N_20936,N_19147,N_19696);
xor U20937 (N_20937,N_19949,N_19541);
xnor U20938 (N_20938,N_19720,N_19455);
nor U20939 (N_20939,N_19993,N_19814);
nand U20940 (N_20940,N_19588,N_19111);
nand U20941 (N_20941,N_19253,N_19842);
or U20942 (N_20942,N_19174,N_19294);
and U20943 (N_20943,N_19109,N_19673);
and U20944 (N_20944,N_19120,N_19515);
and U20945 (N_20945,N_19090,N_19790);
or U20946 (N_20946,N_19042,N_19670);
nand U20947 (N_20947,N_19368,N_19621);
xnor U20948 (N_20948,N_19537,N_19364);
nor U20949 (N_20949,N_19593,N_19278);
and U20950 (N_20950,N_19785,N_19453);
and U20951 (N_20951,N_19678,N_19205);
or U20952 (N_20952,N_19945,N_19245);
or U20953 (N_20953,N_19335,N_19365);
nand U20954 (N_20954,N_19037,N_19814);
or U20955 (N_20955,N_19838,N_19128);
xnor U20956 (N_20956,N_19104,N_19455);
nor U20957 (N_20957,N_19448,N_19583);
nand U20958 (N_20958,N_19409,N_19308);
and U20959 (N_20959,N_19528,N_19746);
xnor U20960 (N_20960,N_19352,N_19192);
nand U20961 (N_20961,N_19412,N_19102);
nand U20962 (N_20962,N_19695,N_19009);
nand U20963 (N_20963,N_19960,N_19161);
xnor U20964 (N_20964,N_19280,N_19003);
and U20965 (N_20965,N_19452,N_19271);
and U20966 (N_20966,N_19179,N_19481);
or U20967 (N_20967,N_19414,N_19972);
and U20968 (N_20968,N_19395,N_19834);
xor U20969 (N_20969,N_19692,N_19909);
xor U20970 (N_20970,N_19156,N_19689);
xor U20971 (N_20971,N_19809,N_19654);
or U20972 (N_20972,N_19312,N_19027);
nand U20973 (N_20973,N_19841,N_19623);
and U20974 (N_20974,N_19006,N_19967);
nor U20975 (N_20975,N_19622,N_19717);
nand U20976 (N_20976,N_19945,N_19599);
or U20977 (N_20977,N_19900,N_19579);
xor U20978 (N_20978,N_19707,N_19891);
and U20979 (N_20979,N_19932,N_19165);
nand U20980 (N_20980,N_19178,N_19012);
nor U20981 (N_20981,N_19445,N_19820);
xnor U20982 (N_20982,N_19670,N_19498);
nand U20983 (N_20983,N_19101,N_19432);
and U20984 (N_20984,N_19183,N_19126);
or U20985 (N_20985,N_19800,N_19667);
or U20986 (N_20986,N_19240,N_19013);
and U20987 (N_20987,N_19127,N_19044);
and U20988 (N_20988,N_19651,N_19132);
nor U20989 (N_20989,N_19990,N_19148);
or U20990 (N_20990,N_19684,N_19735);
nand U20991 (N_20991,N_19757,N_19931);
and U20992 (N_20992,N_19518,N_19840);
or U20993 (N_20993,N_19444,N_19650);
nor U20994 (N_20994,N_19217,N_19903);
xnor U20995 (N_20995,N_19239,N_19010);
nand U20996 (N_20996,N_19767,N_19498);
and U20997 (N_20997,N_19070,N_19495);
and U20998 (N_20998,N_19747,N_19680);
xnor U20999 (N_20999,N_19501,N_19109);
and U21000 (N_21000,N_20338,N_20104);
xnor U21001 (N_21001,N_20337,N_20709);
nor U21002 (N_21002,N_20750,N_20230);
xnor U21003 (N_21003,N_20902,N_20050);
nor U21004 (N_21004,N_20445,N_20650);
or U21005 (N_21005,N_20314,N_20683);
nor U21006 (N_21006,N_20165,N_20033);
and U21007 (N_21007,N_20823,N_20257);
xor U21008 (N_21008,N_20686,N_20935);
nor U21009 (N_21009,N_20582,N_20382);
xor U21010 (N_21010,N_20105,N_20118);
and U21011 (N_21011,N_20941,N_20255);
and U21012 (N_21012,N_20364,N_20990);
and U21013 (N_21013,N_20981,N_20208);
and U21014 (N_21014,N_20646,N_20614);
and U21015 (N_21015,N_20507,N_20845);
nor U21016 (N_21016,N_20980,N_20161);
or U21017 (N_21017,N_20631,N_20626);
xor U21018 (N_21018,N_20694,N_20867);
xor U21019 (N_21019,N_20818,N_20802);
xnor U21020 (N_21020,N_20567,N_20404);
xor U21021 (N_21021,N_20399,N_20770);
and U21022 (N_21022,N_20788,N_20217);
nand U21023 (N_21023,N_20137,N_20253);
nand U21024 (N_21024,N_20463,N_20679);
or U21025 (N_21025,N_20380,N_20886);
nor U21026 (N_21026,N_20263,N_20659);
nand U21027 (N_21027,N_20405,N_20114);
xor U21028 (N_21028,N_20784,N_20157);
xnor U21029 (N_21029,N_20058,N_20147);
and U21030 (N_21030,N_20417,N_20484);
nor U21031 (N_21031,N_20919,N_20304);
xor U21032 (N_21032,N_20123,N_20330);
nand U21033 (N_21033,N_20976,N_20632);
nand U21034 (N_21034,N_20475,N_20102);
or U21035 (N_21035,N_20030,N_20251);
nand U21036 (N_21036,N_20227,N_20052);
nor U21037 (N_21037,N_20651,N_20583);
nand U21038 (N_21038,N_20712,N_20434);
xnor U21039 (N_21039,N_20135,N_20989);
or U21040 (N_21040,N_20863,N_20617);
nor U21041 (N_21041,N_20909,N_20765);
xnor U21042 (N_21042,N_20891,N_20408);
nand U21043 (N_21043,N_20497,N_20495);
xor U21044 (N_21044,N_20645,N_20848);
nor U21045 (N_21045,N_20810,N_20930);
nor U21046 (N_21046,N_20865,N_20874);
or U21047 (N_21047,N_20478,N_20900);
or U21048 (N_21048,N_20799,N_20496);
xnor U21049 (N_21049,N_20216,N_20218);
xor U21050 (N_21050,N_20388,N_20534);
nand U21051 (N_21051,N_20957,N_20668);
xor U21052 (N_21052,N_20093,N_20516);
nand U21053 (N_21053,N_20665,N_20244);
nor U21054 (N_21054,N_20034,N_20661);
xnor U21055 (N_21055,N_20016,N_20013);
nor U21056 (N_21056,N_20004,N_20270);
xor U21057 (N_21057,N_20213,N_20853);
and U21058 (N_21058,N_20524,N_20077);
nor U21059 (N_21059,N_20731,N_20885);
nor U21060 (N_21060,N_20852,N_20793);
nand U21061 (N_21061,N_20097,N_20603);
xor U21062 (N_21062,N_20080,N_20803);
nand U21063 (N_21063,N_20616,N_20317);
or U21064 (N_21064,N_20038,N_20882);
nor U21065 (N_21065,N_20132,N_20881);
or U21066 (N_21066,N_20795,N_20889);
and U21067 (N_21067,N_20069,N_20819);
xor U21068 (N_21068,N_20535,N_20772);
xor U21069 (N_21069,N_20681,N_20978);
nand U21070 (N_21070,N_20843,N_20483);
nand U21071 (N_21071,N_20527,N_20136);
and U21072 (N_21072,N_20986,N_20083);
or U21073 (N_21073,N_20861,N_20271);
or U21074 (N_21074,N_20315,N_20350);
nor U21075 (N_21075,N_20296,N_20760);
and U21076 (N_21076,N_20283,N_20966);
nand U21077 (N_21077,N_20787,N_20722);
or U21078 (N_21078,N_20796,N_20998);
nor U21079 (N_21079,N_20204,N_20313);
nand U21080 (N_21080,N_20736,N_20751);
nor U21081 (N_21081,N_20950,N_20830);
xor U21082 (N_21082,N_20252,N_20409);
nor U21083 (N_21083,N_20566,N_20910);
nand U21084 (N_21084,N_20719,N_20654);
and U21085 (N_21085,N_20913,N_20814);
or U21086 (N_21086,N_20533,N_20997);
and U21087 (N_21087,N_20438,N_20677);
or U21088 (N_21088,N_20492,N_20860);
xor U21089 (N_21089,N_20241,N_20139);
nand U21090 (N_21090,N_20588,N_20844);
or U21091 (N_21091,N_20229,N_20499);
or U21092 (N_21092,N_20285,N_20232);
or U21093 (N_21093,N_20066,N_20074);
nor U21094 (N_21094,N_20329,N_20240);
xor U21095 (N_21095,N_20007,N_20854);
and U21096 (N_21096,N_20243,N_20246);
or U21097 (N_21097,N_20570,N_20426);
nand U21098 (N_21098,N_20505,N_20441);
nand U21099 (N_21099,N_20849,N_20663);
nor U21100 (N_21100,N_20187,N_20647);
or U21101 (N_21101,N_20028,N_20081);
and U21102 (N_21102,N_20198,N_20706);
xor U21103 (N_21103,N_20993,N_20808);
xnor U21104 (N_21104,N_20390,N_20185);
and U21105 (N_21105,N_20444,N_20248);
and U21106 (N_21106,N_20179,N_20847);
nor U21107 (N_21107,N_20413,N_20125);
or U21108 (N_21108,N_20435,N_20449);
or U21109 (N_21109,N_20267,N_20912);
or U21110 (N_21110,N_20121,N_20360);
nand U21111 (N_21111,N_20301,N_20402);
and U21112 (N_21112,N_20658,N_20559);
nor U21113 (N_21113,N_20630,N_20391);
and U21114 (N_21114,N_20932,N_20268);
and U21115 (N_21115,N_20821,N_20831);
and U21116 (N_21116,N_20826,N_20906);
xnor U21117 (N_21117,N_20653,N_20600);
nor U21118 (N_21118,N_20357,N_20711);
nor U21119 (N_21119,N_20680,N_20581);
xor U21120 (N_21120,N_20837,N_20893);
nand U21121 (N_21121,N_20734,N_20374);
nor U21122 (N_21122,N_20988,N_20407);
nor U21123 (N_21123,N_20397,N_20965);
xnor U21124 (N_21124,N_20173,N_20064);
nor U21125 (N_21125,N_20446,N_20688);
nand U21126 (N_21126,N_20384,N_20937);
nor U21127 (N_21127,N_20394,N_20529);
nand U21128 (N_21128,N_20071,N_20816);
xor U21129 (N_21129,N_20353,N_20465);
or U21130 (N_21130,N_20303,N_20592);
nor U21131 (N_21131,N_20428,N_20473);
xor U21132 (N_21132,N_20880,N_20197);
and U21133 (N_21133,N_20541,N_20113);
xor U21134 (N_21134,N_20396,N_20738);
or U21135 (N_21135,N_20487,N_20927);
nor U21136 (N_21136,N_20747,N_20554);
xor U21137 (N_21137,N_20633,N_20172);
nor U21138 (N_21138,N_20648,N_20265);
xnor U21139 (N_21139,N_20723,N_20348);
nand U21140 (N_21140,N_20783,N_20887);
nor U21141 (N_21141,N_20961,N_20207);
or U21142 (N_21142,N_20331,N_20641);
and U21143 (N_21143,N_20078,N_20278);
or U21144 (N_21144,N_20211,N_20203);
nor U21145 (N_21145,N_20868,N_20585);
nand U21146 (N_21146,N_20234,N_20326);
or U21147 (N_21147,N_20356,N_20228);
xor U21148 (N_21148,N_20440,N_20128);
or U21149 (N_21149,N_20596,N_20299);
xor U21150 (N_21150,N_20576,N_20355);
nand U21151 (N_21151,N_20578,N_20838);
nor U21152 (N_21152,N_20580,N_20901);
or U21153 (N_21153,N_20225,N_20460);
and U21154 (N_21154,N_20842,N_20851);
nand U21155 (N_21155,N_20752,N_20850);
or U21156 (N_21156,N_20079,N_20115);
and U21157 (N_21157,N_20552,N_20972);
and U21158 (N_21158,N_20914,N_20491);
and U21159 (N_21159,N_20628,N_20528);
nand U21160 (N_21160,N_20643,N_20133);
or U21161 (N_21161,N_20419,N_20450);
nor U21162 (N_21162,N_20884,N_20824);
or U21163 (N_21163,N_20298,N_20352);
nand U21164 (N_21164,N_20154,N_20952);
xnor U21165 (N_21165,N_20320,N_20468);
nand U21166 (N_21166,N_20876,N_20652);
xor U21167 (N_21167,N_20032,N_20939);
or U21168 (N_21168,N_20191,N_20024);
and U21169 (N_21169,N_20822,N_20755);
and U21170 (N_21170,N_20781,N_20017);
xor U21171 (N_21171,N_20467,N_20649);
nor U21172 (N_21172,N_20942,N_20691);
and U21173 (N_21173,N_20743,N_20547);
xor U21174 (N_21174,N_20864,N_20040);
nor U21175 (N_21175,N_20656,N_20277);
and U21176 (N_21176,N_20716,N_20510);
nand U21177 (N_21177,N_20143,N_20809);
nand U21178 (N_21178,N_20642,N_20447);
nand U21179 (N_21179,N_20586,N_20488);
or U21180 (N_21180,N_20070,N_20205);
xor U21181 (N_21181,N_20292,N_20183);
nor U21182 (N_21182,N_20708,N_20958);
nor U21183 (N_21183,N_20526,N_20142);
xor U21184 (N_21184,N_20372,N_20572);
xor U21185 (N_21185,N_20127,N_20065);
nand U21186 (N_21186,N_20044,N_20046);
or U21187 (N_21187,N_20740,N_20639);
nand U21188 (N_21188,N_20026,N_20791);
and U21189 (N_21189,N_20037,N_20938);
and U21190 (N_21190,N_20280,N_20905);
and U21191 (N_21191,N_20060,N_20875);
or U21192 (N_21192,N_20427,N_20797);
nand U21193 (N_21193,N_20341,N_20202);
nor U21194 (N_21194,N_20525,N_20908);
nor U21195 (N_21195,N_20532,N_20857);
nand U21196 (N_21196,N_20666,N_20917);
nor U21197 (N_21197,N_20381,N_20929);
nand U21198 (N_21198,N_20289,N_20514);
or U21199 (N_21199,N_20715,N_20335);
nand U21200 (N_21200,N_20171,N_20247);
nor U21201 (N_21201,N_20332,N_20856);
nand U21202 (N_21202,N_20945,N_20474);
nor U21203 (N_21203,N_20964,N_20710);
nand U21204 (N_21204,N_20726,N_20778);
nor U21205 (N_21205,N_20705,N_20373);
nor U21206 (N_21206,N_20481,N_20131);
and U21207 (N_21207,N_20221,N_20109);
and U21208 (N_21208,N_20174,N_20602);
nor U21209 (N_21209,N_20879,N_20226);
nor U21210 (N_21210,N_20601,N_20422);
xor U21211 (N_21211,N_20178,N_20180);
xnor U21212 (N_21212,N_20924,N_20604);
nand U21213 (N_21213,N_20798,N_20523);
or U21214 (N_21214,N_20455,N_20089);
nor U21215 (N_21215,N_20704,N_20310);
and U21216 (N_21216,N_20739,N_20223);
nand U21217 (N_21217,N_20212,N_20764);
and U21218 (N_21218,N_20622,N_20748);
xor U21219 (N_21219,N_20318,N_20775);
nor U21220 (N_21220,N_20983,N_20569);
nor U21221 (N_21221,N_20564,N_20005);
nor U21222 (N_21222,N_20101,N_20056);
or U21223 (N_21223,N_20258,N_20521);
nor U21224 (N_21224,N_20866,N_20279);
nand U21225 (N_21225,N_20249,N_20611);
xor U21226 (N_21226,N_20144,N_20480);
xnor U21227 (N_21227,N_20431,N_20951);
nand U21228 (N_21228,N_20994,N_20169);
xnor U21229 (N_21229,N_20266,N_20490);
or U21230 (N_21230,N_20832,N_20073);
xor U21231 (N_21231,N_20464,N_20922);
or U21232 (N_21232,N_20090,N_20638);
and U21233 (N_21233,N_20546,N_20817);
and U21234 (N_21234,N_20012,N_20502);
or U21235 (N_21235,N_20055,N_20053);
and U21236 (N_21236,N_20272,N_20124);
and U21237 (N_21237,N_20096,N_20769);
xnor U21238 (N_21238,N_20327,N_20392);
or U21239 (N_21239,N_20188,N_20098);
and U21240 (N_21240,N_20177,N_20347);
nand U21241 (N_21241,N_20343,N_20754);
and U21242 (N_21242,N_20619,N_20383);
nor U21243 (N_21243,N_20389,N_20512);
or U21244 (N_21244,N_20519,N_20324);
nand U21245 (N_21245,N_20703,N_20563);
and U21246 (N_21246,N_20970,N_20199);
nand U21247 (N_21247,N_20477,N_20916);
xor U21248 (N_21248,N_20940,N_20140);
or U21249 (N_21249,N_20206,N_20003);
and U21250 (N_21250,N_20773,N_20126);
nand U21251 (N_21251,N_20129,N_20513);
nor U21252 (N_21252,N_20443,N_20366);
and U21253 (N_21253,N_20260,N_20762);
xor U21254 (N_21254,N_20757,N_20672);
xnor U21255 (N_21255,N_20749,N_20057);
or U21256 (N_21256,N_20011,N_20295);
nand U21257 (N_21257,N_20707,N_20701);
xnor U21258 (N_21258,N_20615,N_20493);
nand U21259 (N_21259,N_20334,N_20151);
nor U21260 (N_21260,N_20276,N_20210);
and U21261 (N_21261,N_20735,N_20075);
nand U21262 (N_21262,N_20047,N_20148);
and U21263 (N_21263,N_20687,N_20953);
xor U21264 (N_21264,N_20669,N_20061);
or U21265 (N_21265,N_20162,N_20163);
nor U21266 (N_21266,N_20587,N_20813);
nor U21267 (N_21267,N_20084,N_20453);
nor U21268 (N_21268,N_20539,N_20466);
nor U21269 (N_21269,N_20322,N_20517);
or U21270 (N_21270,N_20911,N_20568);
nand U21271 (N_21271,N_20883,N_20287);
nor U21272 (N_21272,N_20936,N_20954);
nor U21273 (N_21273,N_20190,N_20801);
xnor U21274 (N_21274,N_20349,N_20361);
and U21275 (N_21275,N_20926,N_20145);
or U21276 (N_21276,N_20984,N_20685);
or U21277 (N_21277,N_20520,N_20196);
nand U21278 (N_21278,N_20925,N_20156);
or U21279 (N_21279,N_20423,N_20378);
xnor U21280 (N_21280,N_20025,N_20000);
nand U21281 (N_21281,N_20273,N_20968);
xor U21282 (N_21282,N_20598,N_20152);
or U21283 (N_21283,N_20452,N_20424);
nor U21284 (N_21284,N_20437,N_20897);
nor U21285 (N_21285,N_20063,N_20618);
nand U21286 (N_21286,N_20982,N_20209);
or U21287 (N_21287,N_20623,N_20888);
nand U21288 (N_21288,N_20436,N_20675);
xor U21289 (N_21289,N_20933,N_20949);
or U21290 (N_21290,N_20099,N_20194);
xnor U21291 (N_21291,N_20160,N_20410);
nand U21292 (N_21292,N_20130,N_20589);
nor U21293 (N_21293,N_20558,N_20551);
nand U21294 (N_21294,N_20306,N_20479);
nand U21295 (N_21295,N_20009,N_20001);
nand U21296 (N_21296,N_20316,N_20231);
xnor U21297 (N_21297,N_20201,N_20794);
or U21298 (N_21298,N_20948,N_20311);
or U21299 (N_21299,N_20732,N_20693);
nand U21300 (N_21300,N_20106,N_20092);
nand U21301 (N_21301,N_20457,N_20365);
nand U21302 (N_21302,N_20193,N_20758);
or U21303 (N_21303,N_20605,N_20785);
and U21304 (N_21304,N_20947,N_20458);
or U21305 (N_21305,N_20635,N_20690);
xnor U21306 (N_21306,N_20072,N_20833);
xnor U21307 (N_21307,N_20733,N_20138);
nand U21308 (N_21308,N_20931,N_20387);
or U21309 (N_21309,N_20518,N_20293);
or U21310 (N_21310,N_20035,N_20235);
nor U21311 (N_21311,N_20014,N_20175);
nor U21312 (N_21312,N_20091,N_20403);
nand U21313 (N_21313,N_20471,N_20996);
or U21314 (N_21314,N_20029,N_20442);
and U21315 (N_21315,N_20537,N_20472);
or U21316 (N_21316,N_20224,N_20153);
nand U21317 (N_21317,N_20696,N_20049);
nor U21318 (N_21318,N_20088,N_20594);
and U21319 (N_21319,N_20019,N_20667);
nand U21320 (N_21320,N_20591,N_20637);
nor U21321 (N_21321,N_20485,N_20354);
and U21322 (N_21322,N_20565,N_20724);
or U21323 (N_21323,N_20713,N_20612);
or U21324 (N_21324,N_20112,N_20805);
xnor U21325 (N_21325,N_20412,N_20448);
nor U21326 (N_21326,N_20430,N_20269);
and U21327 (N_21327,N_20759,N_20262);
nand U21328 (N_21328,N_20767,N_20944);
xnor U21329 (N_21329,N_20967,N_20176);
nor U21330 (N_21330,N_20192,N_20761);
xor U21331 (N_21331,N_20904,N_20992);
or U21332 (N_21332,N_20398,N_20804);
or U21333 (N_21333,N_20574,N_20233);
nor U21334 (N_21334,N_20184,N_20634);
and U21335 (N_21335,N_20359,N_20553);
nand U21336 (N_21336,N_20041,N_20543);
or U21337 (N_21337,N_20358,N_20429);
nand U21338 (N_21338,N_20921,N_20985);
and U21339 (N_21339,N_20774,N_20571);
xor U21340 (N_21340,N_20421,N_20698);
xnor U21341 (N_21341,N_20274,N_20369);
nor U21342 (N_21342,N_20462,N_20815);
nor U21343 (N_21343,N_20511,N_20342);
xor U21344 (N_21344,N_20590,N_20245);
nor U21345 (N_21345,N_20946,N_20222);
xor U21346 (N_21346,N_20768,N_20974);
and U21347 (N_21347,N_20898,N_20503);
xor U21348 (N_21348,N_20086,N_20219);
and U21349 (N_21349,N_20730,N_20557);
nor U21350 (N_21350,N_20915,N_20008);
nand U21351 (N_21351,N_20841,N_20482);
nor U21352 (N_21352,N_20545,N_20087);
or U21353 (N_21353,N_20870,N_20636);
and U21354 (N_21354,N_20869,N_20379);
nor U21355 (N_21355,N_20340,N_20714);
or U21356 (N_21356,N_20613,N_20780);
or U21357 (N_21357,N_20728,N_20542);
or U21358 (N_21358,N_20045,N_20300);
and U21359 (N_21359,N_20237,N_20345);
nor U21360 (N_21360,N_20987,N_20015);
xor U21361 (N_21361,N_20042,N_20969);
and U21362 (N_21362,N_20536,N_20896);
nand U21363 (N_21363,N_20284,N_20094);
xnor U21364 (N_21364,N_20789,N_20344);
nand U21365 (N_21365,N_20973,N_20051);
nor U21366 (N_21366,N_20835,N_20807);
xor U21367 (N_21367,N_20375,N_20725);
nor U21368 (N_21368,N_20401,N_20022);
or U21369 (N_21369,N_20540,N_20928);
or U21370 (N_21370,N_20095,N_20610);
xor U21371 (N_21371,N_20878,N_20621);
nand U21372 (N_21372,N_20286,N_20195);
or U21373 (N_21373,N_20702,N_20164);
nor U21374 (N_21374,N_20010,N_20662);
nand U21375 (N_21375,N_20048,N_20828);
or U21376 (N_21376,N_20238,N_20515);
and U21377 (N_21377,N_20670,N_20120);
xnor U21378 (N_21378,N_20425,N_20840);
nor U21379 (N_21379,N_20573,N_20556);
nor U21380 (N_21380,N_20021,N_20872);
or U21381 (N_21381,N_20059,N_20744);
xor U21382 (N_21382,N_20454,N_20673);
xnor U21383 (N_21383,N_20544,N_20146);
nand U21384 (N_21384,N_20531,N_20351);
or U21385 (N_21385,N_20393,N_20489);
or U21386 (N_21386,N_20159,N_20376);
nor U21387 (N_21387,N_20700,N_20107);
xnor U21388 (N_21388,N_20756,N_20561);
or U21389 (N_21389,N_20606,N_20336);
and U21390 (N_21390,N_20871,N_20549);
nand U21391 (N_21391,N_20290,N_20082);
xor U21392 (N_21392,N_20302,N_20498);
xnor U21393 (N_21393,N_20043,N_20806);
xor U21394 (N_21394,N_20522,N_20991);
nor U21395 (N_21395,N_20469,N_20456);
and U21396 (N_21396,N_20624,N_20377);
or U21397 (N_21397,N_20811,N_20168);
xnor U21398 (N_21398,N_20333,N_20960);
nand U21399 (N_21399,N_20186,N_20432);
and U21400 (N_21400,N_20555,N_20899);
nor U21401 (N_21401,N_20971,N_20640);
xnor U21402 (N_21402,N_20717,N_20470);
and U21403 (N_21403,N_20779,N_20494);
or U21404 (N_21404,N_20297,N_20786);
xor U21405 (N_21405,N_20655,N_20627);
nand U21406 (N_21406,N_20829,N_20264);
xor U21407 (N_21407,N_20695,N_20170);
nand U21408 (N_21408,N_20149,N_20155);
and U21409 (N_21409,N_20962,N_20439);
nand U21410 (N_21410,N_20501,N_20895);
xnor U21411 (N_21411,N_20562,N_20956);
nor U21412 (N_21412,N_20792,N_20836);
or U21413 (N_21413,N_20119,N_20288);
nor U21414 (N_21414,N_20416,N_20839);
nor U21415 (N_21415,N_20018,N_20955);
and U21416 (N_21416,N_20308,N_20068);
xor U21417 (N_21417,N_20607,N_20242);
and U21418 (N_21418,N_20727,N_20461);
nor U21419 (N_21419,N_20321,N_20858);
or U21420 (N_21420,N_20122,N_20486);
and U21421 (N_21421,N_20776,N_20214);
or U21422 (N_21422,N_20328,N_20977);
nand U21423 (N_21423,N_20721,N_20261);
and U21424 (N_21424,N_20395,N_20599);
and U21425 (N_21425,N_20678,N_20339);
nor U21426 (N_21426,N_20979,N_20777);
and U21427 (N_21427,N_20134,N_20476);
or U21428 (N_21428,N_20923,N_20459);
xnor U21429 (N_21429,N_20312,N_20597);
and U21430 (N_21430,N_20575,N_20890);
and U21431 (N_21431,N_20699,N_20577);
and U21432 (N_21432,N_20746,N_20250);
nand U21433 (N_21433,N_20530,N_20859);
nand U21434 (N_21434,N_20415,N_20414);
xnor U21435 (N_21435,N_20200,N_20508);
xor U21436 (N_21436,N_20593,N_20054);
nand U21437 (N_21437,N_20256,N_20182);
or U21438 (N_21438,N_20110,N_20239);
nor U21439 (N_21439,N_20763,N_20660);
xnor U21440 (N_21440,N_20995,N_20720);
xor U21441 (N_21441,N_20834,N_20085);
nor U21442 (N_21442,N_20236,N_20291);
and U21443 (N_21443,N_20907,N_20674);
xnor U21444 (N_21444,N_20975,N_20418);
and U21445 (N_21445,N_20745,N_20031);
and U21446 (N_21446,N_20560,N_20500);
nor U21447 (N_21447,N_20873,N_20167);
or U21448 (N_21448,N_20892,N_20371);
or U21449 (N_21449,N_20620,N_20215);
nand U21450 (N_21450,N_20741,N_20509);
and U21451 (N_21451,N_20282,N_20999);
nand U21452 (N_21452,N_20370,N_20305);
or U21453 (N_21453,N_20006,N_20689);
nor U21454 (N_21454,N_20385,N_20812);
nor U21455 (N_21455,N_20737,N_20166);
nand U21456 (N_21456,N_20400,N_20319);
or U21457 (N_21457,N_20963,N_20002);
and U21458 (N_21458,N_20684,N_20692);
nor U21459 (N_21459,N_20504,N_20367);
xor U21460 (N_21460,N_20406,N_20903);
or U21461 (N_21461,N_20420,N_20629);
and U21462 (N_21462,N_20325,N_20020);
nor U21463 (N_21463,N_20934,N_20411);
nor U21464 (N_21464,N_20076,N_20254);
nand U21465 (N_21465,N_20117,N_20894);
xnor U21466 (N_21466,N_20800,N_20920);
nand U21467 (N_21467,N_20386,N_20067);
nor U21468 (N_21468,N_20676,N_20943);
or U21469 (N_21469,N_20433,N_20103);
nor U21470 (N_21470,N_20959,N_20664);
or U21471 (N_21471,N_20657,N_20141);
or U21472 (N_21472,N_20729,N_20150);
nor U21473 (N_21473,N_20346,N_20742);
nor U21474 (N_21474,N_20281,N_20644);
nor U21475 (N_21475,N_20189,N_20023);
nor U21476 (N_21476,N_20584,N_20275);
nand U21477 (N_21477,N_20827,N_20108);
and U21478 (N_21478,N_20362,N_20918);
or U21479 (N_21479,N_20181,N_20309);
xnor U21480 (N_21480,N_20595,N_20766);
and U21481 (N_21481,N_20111,N_20855);
or U21482 (N_21482,N_20259,N_20579);
or U21483 (N_21483,N_20039,N_20820);
or U21484 (N_21484,N_20718,N_20609);
or U21485 (N_21485,N_20307,N_20825);
nand U21486 (N_21486,N_20506,N_20363);
xor U21487 (N_21487,N_20220,N_20027);
and U21488 (N_21488,N_20538,N_20782);
or U21489 (N_21489,N_20451,N_20294);
nand U21490 (N_21490,N_20877,N_20368);
nand U21491 (N_21491,N_20753,N_20790);
nand U21492 (N_21492,N_20550,N_20100);
nor U21493 (N_21493,N_20036,N_20116);
or U21494 (N_21494,N_20682,N_20697);
or U21495 (N_21495,N_20548,N_20846);
xor U21496 (N_21496,N_20062,N_20671);
xnor U21497 (N_21497,N_20323,N_20608);
or U21498 (N_21498,N_20771,N_20625);
nor U21499 (N_21499,N_20158,N_20862);
nand U21500 (N_21500,N_20835,N_20792);
xnor U21501 (N_21501,N_20312,N_20625);
nand U21502 (N_21502,N_20409,N_20898);
xnor U21503 (N_21503,N_20988,N_20761);
nand U21504 (N_21504,N_20917,N_20129);
nor U21505 (N_21505,N_20132,N_20909);
nand U21506 (N_21506,N_20599,N_20041);
and U21507 (N_21507,N_20947,N_20906);
and U21508 (N_21508,N_20181,N_20566);
and U21509 (N_21509,N_20645,N_20750);
nor U21510 (N_21510,N_20735,N_20189);
and U21511 (N_21511,N_20749,N_20387);
and U21512 (N_21512,N_20772,N_20835);
xor U21513 (N_21513,N_20880,N_20447);
nand U21514 (N_21514,N_20646,N_20648);
or U21515 (N_21515,N_20934,N_20040);
and U21516 (N_21516,N_20017,N_20294);
and U21517 (N_21517,N_20037,N_20468);
and U21518 (N_21518,N_20480,N_20265);
nor U21519 (N_21519,N_20840,N_20889);
xor U21520 (N_21520,N_20519,N_20963);
xor U21521 (N_21521,N_20558,N_20067);
nand U21522 (N_21522,N_20680,N_20258);
nor U21523 (N_21523,N_20448,N_20881);
or U21524 (N_21524,N_20338,N_20828);
nor U21525 (N_21525,N_20613,N_20956);
or U21526 (N_21526,N_20379,N_20375);
nor U21527 (N_21527,N_20898,N_20628);
and U21528 (N_21528,N_20931,N_20485);
nor U21529 (N_21529,N_20299,N_20863);
and U21530 (N_21530,N_20484,N_20029);
nor U21531 (N_21531,N_20882,N_20918);
and U21532 (N_21532,N_20716,N_20112);
nand U21533 (N_21533,N_20287,N_20163);
or U21534 (N_21534,N_20692,N_20060);
xnor U21535 (N_21535,N_20901,N_20377);
nand U21536 (N_21536,N_20851,N_20996);
nand U21537 (N_21537,N_20646,N_20484);
and U21538 (N_21538,N_20373,N_20071);
nand U21539 (N_21539,N_20752,N_20109);
xor U21540 (N_21540,N_20792,N_20204);
or U21541 (N_21541,N_20279,N_20118);
nor U21542 (N_21542,N_20409,N_20850);
or U21543 (N_21543,N_20132,N_20742);
nand U21544 (N_21544,N_20683,N_20345);
nand U21545 (N_21545,N_20525,N_20375);
xor U21546 (N_21546,N_20040,N_20534);
and U21547 (N_21547,N_20557,N_20902);
and U21548 (N_21548,N_20656,N_20065);
nor U21549 (N_21549,N_20127,N_20922);
or U21550 (N_21550,N_20840,N_20634);
nor U21551 (N_21551,N_20476,N_20877);
xor U21552 (N_21552,N_20759,N_20930);
and U21553 (N_21553,N_20017,N_20171);
or U21554 (N_21554,N_20201,N_20728);
xnor U21555 (N_21555,N_20760,N_20231);
nand U21556 (N_21556,N_20780,N_20776);
nand U21557 (N_21557,N_20794,N_20820);
or U21558 (N_21558,N_20374,N_20806);
xnor U21559 (N_21559,N_20830,N_20136);
nand U21560 (N_21560,N_20236,N_20078);
or U21561 (N_21561,N_20236,N_20905);
and U21562 (N_21562,N_20517,N_20300);
or U21563 (N_21563,N_20633,N_20935);
nand U21564 (N_21564,N_20583,N_20850);
nand U21565 (N_21565,N_20448,N_20525);
or U21566 (N_21566,N_20308,N_20730);
or U21567 (N_21567,N_20461,N_20056);
nor U21568 (N_21568,N_20358,N_20447);
xnor U21569 (N_21569,N_20039,N_20941);
and U21570 (N_21570,N_20495,N_20329);
xnor U21571 (N_21571,N_20727,N_20652);
and U21572 (N_21572,N_20022,N_20838);
nor U21573 (N_21573,N_20179,N_20485);
nor U21574 (N_21574,N_20477,N_20218);
nand U21575 (N_21575,N_20738,N_20263);
xor U21576 (N_21576,N_20239,N_20380);
and U21577 (N_21577,N_20337,N_20670);
nand U21578 (N_21578,N_20118,N_20139);
or U21579 (N_21579,N_20153,N_20398);
and U21580 (N_21580,N_20209,N_20042);
xnor U21581 (N_21581,N_20424,N_20996);
or U21582 (N_21582,N_20615,N_20005);
and U21583 (N_21583,N_20287,N_20526);
and U21584 (N_21584,N_20540,N_20054);
and U21585 (N_21585,N_20897,N_20689);
nand U21586 (N_21586,N_20580,N_20205);
xor U21587 (N_21587,N_20764,N_20680);
or U21588 (N_21588,N_20508,N_20217);
nor U21589 (N_21589,N_20744,N_20807);
or U21590 (N_21590,N_20800,N_20338);
and U21591 (N_21591,N_20713,N_20019);
nor U21592 (N_21592,N_20807,N_20850);
nand U21593 (N_21593,N_20014,N_20792);
nor U21594 (N_21594,N_20724,N_20895);
xor U21595 (N_21595,N_20893,N_20161);
xor U21596 (N_21596,N_20718,N_20035);
xnor U21597 (N_21597,N_20486,N_20798);
or U21598 (N_21598,N_20300,N_20158);
or U21599 (N_21599,N_20794,N_20297);
or U21600 (N_21600,N_20000,N_20782);
nor U21601 (N_21601,N_20591,N_20095);
nor U21602 (N_21602,N_20847,N_20000);
nand U21603 (N_21603,N_20748,N_20352);
xor U21604 (N_21604,N_20427,N_20737);
or U21605 (N_21605,N_20018,N_20404);
or U21606 (N_21606,N_20568,N_20850);
and U21607 (N_21607,N_20915,N_20590);
and U21608 (N_21608,N_20971,N_20149);
or U21609 (N_21609,N_20652,N_20070);
nand U21610 (N_21610,N_20834,N_20399);
and U21611 (N_21611,N_20355,N_20822);
nor U21612 (N_21612,N_20404,N_20580);
nand U21613 (N_21613,N_20039,N_20116);
or U21614 (N_21614,N_20586,N_20053);
xor U21615 (N_21615,N_20359,N_20931);
xnor U21616 (N_21616,N_20596,N_20854);
or U21617 (N_21617,N_20361,N_20674);
nand U21618 (N_21618,N_20825,N_20357);
nand U21619 (N_21619,N_20066,N_20217);
and U21620 (N_21620,N_20075,N_20895);
and U21621 (N_21621,N_20234,N_20701);
xnor U21622 (N_21622,N_20883,N_20850);
or U21623 (N_21623,N_20505,N_20501);
nand U21624 (N_21624,N_20431,N_20657);
xor U21625 (N_21625,N_20665,N_20989);
nand U21626 (N_21626,N_20160,N_20255);
nand U21627 (N_21627,N_20708,N_20214);
and U21628 (N_21628,N_20331,N_20937);
nor U21629 (N_21629,N_20488,N_20803);
xor U21630 (N_21630,N_20676,N_20173);
and U21631 (N_21631,N_20076,N_20918);
or U21632 (N_21632,N_20825,N_20039);
nor U21633 (N_21633,N_20803,N_20477);
or U21634 (N_21634,N_20290,N_20889);
nand U21635 (N_21635,N_20744,N_20334);
and U21636 (N_21636,N_20824,N_20783);
nor U21637 (N_21637,N_20356,N_20419);
or U21638 (N_21638,N_20014,N_20618);
xnor U21639 (N_21639,N_20574,N_20542);
or U21640 (N_21640,N_20607,N_20449);
nand U21641 (N_21641,N_20756,N_20140);
nor U21642 (N_21642,N_20452,N_20105);
xnor U21643 (N_21643,N_20692,N_20506);
xor U21644 (N_21644,N_20148,N_20828);
or U21645 (N_21645,N_20142,N_20314);
nand U21646 (N_21646,N_20258,N_20793);
nor U21647 (N_21647,N_20272,N_20686);
xnor U21648 (N_21648,N_20300,N_20094);
nor U21649 (N_21649,N_20785,N_20682);
nor U21650 (N_21650,N_20311,N_20431);
xnor U21651 (N_21651,N_20533,N_20273);
or U21652 (N_21652,N_20223,N_20614);
nor U21653 (N_21653,N_20281,N_20354);
xor U21654 (N_21654,N_20786,N_20860);
nand U21655 (N_21655,N_20901,N_20863);
or U21656 (N_21656,N_20466,N_20337);
and U21657 (N_21657,N_20931,N_20112);
xnor U21658 (N_21658,N_20136,N_20834);
xor U21659 (N_21659,N_20187,N_20835);
and U21660 (N_21660,N_20386,N_20126);
nor U21661 (N_21661,N_20739,N_20815);
xnor U21662 (N_21662,N_20415,N_20516);
xnor U21663 (N_21663,N_20425,N_20737);
or U21664 (N_21664,N_20108,N_20433);
and U21665 (N_21665,N_20152,N_20256);
nor U21666 (N_21666,N_20103,N_20262);
nand U21667 (N_21667,N_20585,N_20920);
or U21668 (N_21668,N_20921,N_20837);
nor U21669 (N_21669,N_20517,N_20957);
or U21670 (N_21670,N_20894,N_20816);
xor U21671 (N_21671,N_20335,N_20074);
and U21672 (N_21672,N_20058,N_20435);
xnor U21673 (N_21673,N_20685,N_20928);
and U21674 (N_21674,N_20927,N_20064);
nor U21675 (N_21675,N_20624,N_20170);
nand U21676 (N_21676,N_20693,N_20199);
xnor U21677 (N_21677,N_20244,N_20015);
and U21678 (N_21678,N_20681,N_20882);
and U21679 (N_21679,N_20480,N_20807);
nor U21680 (N_21680,N_20861,N_20701);
xor U21681 (N_21681,N_20858,N_20466);
nand U21682 (N_21682,N_20819,N_20815);
xnor U21683 (N_21683,N_20515,N_20362);
xnor U21684 (N_21684,N_20095,N_20904);
and U21685 (N_21685,N_20539,N_20724);
and U21686 (N_21686,N_20959,N_20506);
or U21687 (N_21687,N_20298,N_20879);
xnor U21688 (N_21688,N_20761,N_20345);
nand U21689 (N_21689,N_20443,N_20967);
xor U21690 (N_21690,N_20232,N_20647);
nor U21691 (N_21691,N_20086,N_20311);
and U21692 (N_21692,N_20208,N_20917);
and U21693 (N_21693,N_20138,N_20918);
or U21694 (N_21694,N_20082,N_20863);
and U21695 (N_21695,N_20375,N_20705);
or U21696 (N_21696,N_20663,N_20467);
and U21697 (N_21697,N_20854,N_20896);
nand U21698 (N_21698,N_20775,N_20336);
xnor U21699 (N_21699,N_20481,N_20600);
or U21700 (N_21700,N_20114,N_20238);
nor U21701 (N_21701,N_20659,N_20020);
xor U21702 (N_21702,N_20623,N_20491);
and U21703 (N_21703,N_20516,N_20804);
and U21704 (N_21704,N_20549,N_20936);
nor U21705 (N_21705,N_20824,N_20867);
and U21706 (N_21706,N_20776,N_20972);
nand U21707 (N_21707,N_20824,N_20330);
nand U21708 (N_21708,N_20160,N_20295);
and U21709 (N_21709,N_20156,N_20732);
nand U21710 (N_21710,N_20011,N_20560);
nand U21711 (N_21711,N_20540,N_20747);
xor U21712 (N_21712,N_20668,N_20313);
xnor U21713 (N_21713,N_20620,N_20428);
nor U21714 (N_21714,N_20833,N_20770);
nor U21715 (N_21715,N_20942,N_20162);
or U21716 (N_21716,N_20492,N_20856);
nor U21717 (N_21717,N_20566,N_20220);
nand U21718 (N_21718,N_20744,N_20804);
nand U21719 (N_21719,N_20113,N_20364);
nor U21720 (N_21720,N_20090,N_20555);
nand U21721 (N_21721,N_20227,N_20543);
xor U21722 (N_21722,N_20891,N_20771);
and U21723 (N_21723,N_20328,N_20493);
nor U21724 (N_21724,N_20940,N_20820);
and U21725 (N_21725,N_20038,N_20458);
and U21726 (N_21726,N_20953,N_20955);
or U21727 (N_21727,N_20783,N_20025);
or U21728 (N_21728,N_20345,N_20903);
xor U21729 (N_21729,N_20510,N_20429);
nand U21730 (N_21730,N_20396,N_20277);
nand U21731 (N_21731,N_20681,N_20125);
and U21732 (N_21732,N_20631,N_20545);
or U21733 (N_21733,N_20681,N_20608);
xor U21734 (N_21734,N_20699,N_20731);
nor U21735 (N_21735,N_20265,N_20956);
and U21736 (N_21736,N_20313,N_20943);
and U21737 (N_21737,N_20540,N_20317);
nor U21738 (N_21738,N_20998,N_20883);
nor U21739 (N_21739,N_20410,N_20885);
xor U21740 (N_21740,N_20951,N_20909);
and U21741 (N_21741,N_20132,N_20896);
xnor U21742 (N_21742,N_20585,N_20592);
or U21743 (N_21743,N_20894,N_20134);
nand U21744 (N_21744,N_20249,N_20351);
nand U21745 (N_21745,N_20957,N_20018);
or U21746 (N_21746,N_20902,N_20237);
nor U21747 (N_21747,N_20681,N_20577);
xnor U21748 (N_21748,N_20099,N_20699);
and U21749 (N_21749,N_20052,N_20322);
and U21750 (N_21750,N_20166,N_20053);
nor U21751 (N_21751,N_20273,N_20389);
nor U21752 (N_21752,N_20196,N_20974);
nor U21753 (N_21753,N_20438,N_20521);
xnor U21754 (N_21754,N_20591,N_20189);
nand U21755 (N_21755,N_20723,N_20696);
and U21756 (N_21756,N_20134,N_20612);
or U21757 (N_21757,N_20993,N_20866);
xor U21758 (N_21758,N_20323,N_20855);
nand U21759 (N_21759,N_20292,N_20791);
nor U21760 (N_21760,N_20624,N_20773);
xor U21761 (N_21761,N_20995,N_20412);
or U21762 (N_21762,N_20236,N_20721);
or U21763 (N_21763,N_20975,N_20260);
nand U21764 (N_21764,N_20395,N_20503);
and U21765 (N_21765,N_20626,N_20305);
nor U21766 (N_21766,N_20045,N_20892);
xnor U21767 (N_21767,N_20432,N_20984);
xor U21768 (N_21768,N_20553,N_20290);
xnor U21769 (N_21769,N_20100,N_20058);
nand U21770 (N_21770,N_20355,N_20365);
xor U21771 (N_21771,N_20388,N_20231);
xnor U21772 (N_21772,N_20551,N_20168);
xnor U21773 (N_21773,N_20397,N_20799);
and U21774 (N_21774,N_20463,N_20047);
or U21775 (N_21775,N_20261,N_20883);
nand U21776 (N_21776,N_20219,N_20343);
nor U21777 (N_21777,N_20892,N_20258);
nand U21778 (N_21778,N_20899,N_20731);
nand U21779 (N_21779,N_20831,N_20009);
nand U21780 (N_21780,N_20989,N_20556);
nand U21781 (N_21781,N_20197,N_20657);
xnor U21782 (N_21782,N_20922,N_20049);
nor U21783 (N_21783,N_20339,N_20309);
xnor U21784 (N_21784,N_20613,N_20776);
and U21785 (N_21785,N_20855,N_20295);
and U21786 (N_21786,N_20558,N_20350);
nor U21787 (N_21787,N_20864,N_20600);
and U21788 (N_21788,N_20480,N_20244);
or U21789 (N_21789,N_20664,N_20910);
xor U21790 (N_21790,N_20191,N_20617);
nand U21791 (N_21791,N_20890,N_20431);
or U21792 (N_21792,N_20389,N_20230);
xor U21793 (N_21793,N_20871,N_20728);
nor U21794 (N_21794,N_20060,N_20929);
nor U21795 (N_21795,N_20487,N_20269);
or U21796 (N_21796,N_20325,N_20629);
xor U21797 (N_21797,N_20022,N_20567);
or U21798 (N_21798,N_20391,N_20427);
or U21799 (N_21799,N_20405,N_20059);
and U21800 (N_21800,N_20979,N_20485);
and U21801 (N_21801,N_20327,N_20248);
and U21802 (N_21802,N_20466,N_20424);
nor U21803 (N_21803,N_20146,N_20736);
nor U21804 (N_21804,N_20438,N_20728);
or U21805 (N_21805,N_20872,N_20859);
and U21806 (N_21806,N_20497,N_20545);
or U21807 (N_21807,N_20118,N_20238);
and U21808 (N_21808,N_20344,N_20838);
and U21809 (N_21809,N_20150,N_20272);
nand U21810 (N_21810,N_20153,N_20767);
nand U21811 (N_21811,N_20727,N_20990);
or U21812 (N_21812,N_20309,N_20657);
and U21813 (N_21813,N_20102,N_20498);
nor U21814 (N_21814,N_20888,N_20344);
xor U21815 (N_21815,N_20256,N_20236);
or U21816 (N_21816,N_20607,N_20903);
nand U21817 (N_21817,N_20299,N_20237);
nor U21818 (N_21818,N_20691,N_20819);
xnor U21819 (N_21819,N_20176,N_20307);
or U21820 (N_21820,N_20861,N_20816);
nand U21821 (N_21821,N_20267,N_20229);
or U21822 (N_21822,N_20442,N_20915);
or U21823 (N_21823,N_20305,N_20690);
nor U21824 (N_21824,N_20658,N_20792);
nor U21825 (N_21825,N_20896,N_20934);
or U21826 (N_21826,N_20774,N_20278);
xor U21827 (N_21827,N_20336,N_20745);
nand U21828 (N_21828,N_20628,N_20932);
or U21829 (N_21829,N_20430,N_20774);
and U21830 (N_21830,N_20480,N_20383);
xor U21831 (N_21831,N_20708,N_20473);
xor U21832 (N_21832,N_20453,N_20144);
or U21833 (N_21833,N_20956,N_20401);
xnor U21834 (N_21834,N_20788,N_20667);
xnor U21835 (N_21835,N_20135,N_20011);
nor U21836 (N_21836,N_20091,N_20975);
xor U21837 (N_21837,N_20880,N_20746);
or U21838 (N_21838,N_20810,N_20768);
xnor U21839 (N_21839,N_20333,N_20133);
nor U21840 (N_21840,N_20380,N_20214);
or U21841 (N_21841,N_20797,N_20830);
nor U21842 (N_21842,N_20239,N_20752);
or U21843 (N_21843,N_20373,N_20911);
nor U21844 (N_21844,N_20677,N_20473);
nand U21845 (N_21845,N_20259,N_20699);
nor U21846 (N_21846,N_20278,N_20397);
nand U21847 (N_21847,N_20726,N_20617);
or U21848 (N_21848,N_20278,N_20732);
and U21849 (N_21849,N_20481,N_20726);
nand U21850 (N_21850,N_20832,N_20108);
xor U21851 (N_21851,N_20902,N_20598);
nor U21852 (N_21852,N_20646,N_20777);
nor U21853 (N_21853,N_20369,N_20043);
nor U21854 (N_21854,N_20181,N_20992);
nor U21855 (N_21855,N_20985,N_20742);
nand U21856 (N_21856,N_20484,N_20345);
or U21857 (N_21857,N_20451,N_20742);
nand U21858 (N_21858,N_20494,N_20156);
nor U21859 (N_21859,N_20380,N_20589);
and U21860 (N_21860,N_20135,N_20763);
and U21861 (N_21861,N_20542,N_20592);
or U21862 (N_21862,N_20621,N_20097);
xnor U21863 (N_21863,N_20404,N_20459);
nor U21864 (N_21864,N_20898,N_20363);
or U21865 (N_21865,N_20898,N_20362);
nor U21866 (N_21866,N_20063,N_20043);
or U21867 (N_21867,N_20279,N_20393);
nand U21868 (N_21868,N_20167,N_20179);
and U21869 (N_21869,N_20237,N_20213);
nor U21870 (N_21870,N_20738,N_20879);
and U21871 (N_21871,N_20204,N_20794);
or U21872 (N_21872,N_20333,N_20821);
or U21873 (N_21873,N_20183,N_20882);
nand U21874 (N_21874,N_20021,N_20317);
and U21875 (N_21875,N_20475,N_20492);
nor U21876 (N_21876,N_20672,N_20405);
or U21877 (N_21877,N_20232,N_20059);
nand U21878 (N_21878,N_20771,N_20620);
nor U21879 (N_21879,N_20283,N_20573);
and U21880 (N_21880,N_20873,N_20465);
nor U21881 (N_21881,N_20488,N_20664);
nor U21882 (N_21882,N_20810,N_20162);
or U21883 (N_21883,N_20884,N_20134);
and U21884 (N_21884,N_20045,N_20333);
xnor U21885 (N_21885,N_20804,N_20058);
or U21886 (N_21886,N_20660,N_20665);
or U21887 (N_21887,N_20777,N_20370);
xor U21888 (N_21888,N_20761,N_20661);
and U21889 (N_21889,N_20978,N_20157);
xor U21890 (N_21890,N_20628,N_20493);
nand U21891 (N_21891,N_20157,N_20955);
nor U21892 (N_21892,N_20822,N_20037);
or U21893 (N_21893,N_20312,N_20623);
nand U21894 (N_21894,N_20507,N_20576);
xor U21895 (N_21895,N_20183,N_20902);
nor U21896 (N_21896,N_20154,N_20380);
nand U21897 (N_21897,N_20395,N_20731);
nand U21898 (N_21898,N_20956,N_20955);
nand U21899 (N_21899,N_20399,N_20256);
or U21900 (N_21900,N_20475,N_20208);
and U21901 (N_21901,N_20064,N_20272);
xnor U21902 (N_21902,N_20484,N_20948);
or U21903 (N_21903,N_20805,N_20308);
nor U21904 (N_21904,N_20693,N_20724);
xnor U21905 (N_21905,N_20185,N_20276);
nor U21906 (N_21906,N_20289,N_20023);
xor U21907 (N_21907,N_20284,N_20977);
nand U21908 (N_21908,N_20947,N_20589);
or U21909 (N_21909,N_20578,N_20862);
nand U21910 (N_21910,N_20563,N_20190);
nand U21911 (N_21911,N_20067,N_20625);
nand U21912 (N_21912,N_20497,N_20044);
nor U21913 (N_21913,N_20231,N_20918);
nor U21914 (N_21914,N_20186,N_20583);
nand U21915 (N_21915,N_20484,N_20693);
and U21916 (N_21916,N_20756,N_20037);
nor U21917 (N_21917,N_20683,N_20999);
nor U21918 (N_21918,N_20185,N_20216);
and U21919 (N_21919,N_20964,N_20780);
nor U21920 (N_21920,N_20115,N_20385);
and U21921 (N_21921,N_20125,N_20294);
nor U21922 (N_21922,N_20143,N_20538);
nand U21923 (N_21923,N_20460,N_20638);
nand U21924 (N_21924,N_20890,N_20393);
xnor U21925 (N_21925,N_20695,N_20883);
and U21926 (N_21926,N_20042,N_20479);
xnor U21927 (N_21927,N_20948,N_20782);
xor U21928 (N_21928,N_20044,N_20687);
and U21929 (N_21929,N_20393,N_20441);
xnor U21930 (N_21930,N_20715,N_20872);
and U21931 (N_21931,N_20777,N_20798);
or U21932 (N_21932,N_20452,N_20725);
nor U21933 (N_21933,N_20982,N_20276);
and U21934 (N_21934,N_20620,N_20892);
or U21935 (N_21935,N_20077,N_20245);
nor U21936 (N_21936,N_20837,N_20298);
and U21937 (N_21937,N_20007,N_20532);
and U21938 (N_21938,N_20667,N_20958);
nand U21939 (N_21939,N_20958,N_20695);
nand U21940 (N_21940,N_20873,N_20327);
and U21941 (N_21941,N_20953,N_20189);
or U21942 (N_21942,N_20549,N_20391);
xnor U21943 (N_21943,N_20809,N_20099);
nor U21944 (N_21944,N_20224,N_20064);
xor U21945 (N_21945,N_20054,N_20544);
nor U21946 (N_21946,N_20401,N_20164);
and U21947 (N_21947,N_20044,N_20785);
xor U21948 (N_21948,N_20622,N_20264);
and U21949 (N_21949,N_20814,N_20044);
nand U21950 (N_21950,N_20447,N_20129);
and U21951 (N_21951,N_20956,N_20901);
nor U21952 (N_21952,N_20443,N_20156);
xor U21953 (N_21953,N_20595,N_20952);
or U21954 (N_21954,N_20729,N_20781);
nor U21955 (N_21955,N_20147,N_20098);
and U21956 (N_21956,N_20737,N_20319);
xnor U21957 (N_21957,N_20088,N_20554);
and U21958 (N_21958,N_20697,N_20310);
and U21959 (N_21959,N_20073,N_20636);
and U21960 (N_21960,N_20817,N_20995);
and U21961 (N_21961,N_20797,N_20394);
or U21962 (N_21962,N_20640,N_20308);
or U21963 (N_21963,N_20900,N_20005);
xnor U21964 (N_21964,N_20287,N_20040);
nor U21965 (N_21965,N_20535,N_20411);
nand U21966 (N_21966,N_20364,N_20874);
xor U21967 (N_21967,N_20122,N_20453);
or U21968 (N_21968,N_20728,N_20509);
and U21969 (N_21969,N_20245,N_20279);
nor U21970 (N_21970,N_20726,N_20884);
nor U21971 (N_21971,N_20355,N_20402);
and U21972 (N_21972,N_20373,N_20057);
nor U21973 (N_21973,N_20179,N_20215);
and U21974 (N_21974,N_20358,N_20857);
xnor U21975 (N_21975,N_20270,N_20032);
or U21976 (N_21976,N_20091,N_20669);
xnor U21977 (N_21977,N_20386,N_20618);
nand U21978 (N_21978,N_20953,N_20783);
nand U21979 (N_21979,N_20939,N_20704);
nand U21980 (N_21980,N_20584,N_20529);
and U21981 (N_21981,N_20886,N_20497);
or U21982 (N_21982,N_20688,N_20677);
or U21983 (N_21983,N_20508,N_20760);
nand U21984 (N_21984,N_20075,N_20632);
nor U21985 (N_21985,N_20503,N_20609);
nand U21986 (N_21986,N_20987,N_20709);
and U21987 (N_21987,N_20762,N_20279);
xnor U21988 (N_21988,N_20285,N_20288);
and U21989 (N_21989,N_20837,N_20533);
and U21990 (N_21990,N_20841,N_20513);
xor U21991 (N_21991,N_20946,N_20667);
nor U21992 (N_21992,N_20806,N_20968);
nor U21993 (N_21993,N_20109,N_20065);
nand U21994 (N_21994,N_20316,N_20470);
or U21995 (N_21995,N_20238,N_20113);
nand U21996 (N_21996,N_20878,N_20690);
and U21997 (N_21997,N_20529,N_20864);
xnor U21998 (N_21998,N_20157,N_20004);
xnor U21999 (N_21999,N_20871,N_20672);
nand U22000 (N_22000,N_21586,N_21462);
xnor U22001 (N_22001,N_21339,N_21759);
xnor U22002 (N_22002,N_21865,N_21786);
and U22003 (N_22003,N_21286,N_21943);
xnor U22004 (N_22004,N_21141,N_21899);
nand U22005 (N_22005,N_21739,N_21548);
nor U22006 (N_22006,N_21640,N_21432);
or U22007 (N_22007,N_21061,N_21751);
and U22008 (N_22008,N_21258,N_21169);
or U22009 (N_22009,N_21316,N_21552);
or U22010 (N_22010,N_21594,N_21438);
and U22011 (N_22011,N_21585,N_21160);
xor U22012 (N_22012,N_21058,N_21372);
nand U22013 (N_22013,N_21748,N_21648);
xnor U22014 (N_22014,N_21939,N_21590);
nor U22015 (N_22015,N_21431,N_21181);
xnor U22016 (N_22016,N_21437,N_21935);
and U22017 (N_22017,N_21892,N_21091);
nor U22018 (N_22018,N_21234,N_21376);
and U22019 (N_22019,N_21832,N_21714);
nor U22020 (N_22020,N_21592,N_21205);
xor U22021 (N_22021,N_21427,N_21332);
nor U22022 (N_22022,N_21472,N_21127);
and U22023 (N_22023,N_21811,N_21595);
and U22024 (N_22024,N_21249,N_21496);
xnor U22025 (N_22025,N_21424,N_21840);
and U22026 (N_22026,N_21220,N_21947);
and U22027 (N_22027,N_21756,N_21370);
xor U22028 (N_22028,N_21508,N_21093);
or U22029 (N_22029,N_21991,N_21499);
nand U22030 (N_22030,N_21521,N_21494);
or U22031 (N_22031,N_21351,N_21192);
or U22032 (N_22032,N_21694,N_21107);
xor U22033 (N_22033,N_21771,N_21361);
or U22034 (N_22034,N_21932,N_21890);
nand U22035 (N_22035,N_21773,N_21902);
nand U22036 (N_22036,N_21262,N_21338);
nand U22037 (N_22037,N_21425,N_21356);
nor U22038 (N_22038,N_21214,N_21867);
or U22039 (N_22039,N_21426,N_21185);
and U22040 (N_22040,N_21956,N_21306);
nor U22041 (N_22041,N_21803,N_21682);
xor U22042 (N_22042,N_21394,N_21955);
or U22043 (N_22043,N_21466,N_21843);
or U22044 (N_22044,N_21422,N_21707);
nand U22045 (N_22045,N_21830,N_21129);
nor U22046 (N_22046,N_21657,N_21727);
or U22047 (N_22047,N_21551,N_21550);
nor U22048 (N_22048,N_21591,N_21568);
or U22049 (N_22049,N_21813,N_21664);
nor U22050 (N_22050,N_21027,N_21311);
or U22051 (N_22051,N_21400,N_21581);
and U22052 (N_22052,N_21645,N_21421);
nand U22053 (N_22053,N_21623,N_21252);
xor U22054 (N_22054,N_21742,N_21520);
and U22055 (N_22055,N_21495,N_21650);
xnor U22056 (N_22056,N_21024,N_21999);
nor U22057 (N_22057,N_21718,N_21194);
and U22058 (N_22058,N_21886,N_21760);
or U22059 (N_22059,N_21769,N_21284);
nand U22060 (N_22060,N_21383,N_21159);
xnor U22061 (N_22061,N_21534,N_21570);
nor U22062 (N_22062,N_21687,N_21195);
nand U22063 (N_22063,N_21621,N_21860);
xor U22064 (N_22064,N_21905,N_21131);
xor U22065 (N_22065,N_21271,N_21193);
and U22066 (N_22066,N_21066,N_21248);
or U22067 (N_22067,N_21894,N_21877);
or U22068 (N_22068,N_21084,N_21858);
or U22069 (N_22069,N_21602,N_21282);
and U22070 (N_22070,N_21580,N_21331);
and U22071 (N_22071,N_21766,N_21480);
nand U22072 (N_22072,N_21228,N_21683);
or U22073 (N_22073,N_21269,N_21299);
nor U22074 (N_22074,N_21785,N_21844);
nand U22075 (N_22075,N_21003,N_21671);
or U22076 (N_22076,N_21578,N_21676);
or U22077 (N_22077,N_21908,N_21665);
xor U22078 (N_22078,N_21577,N_21283);
and U22079 (N_22079,N_21133,N_21232);
and U22080 (N_22080,N_21642,N_21936);
or U22081 (N_22081,N_21746,N_21154);
or U22082 (N_22082,N_21673,N_21517);
nor U22083 (N_22083,N_21478,N_21810);
xor U22084 (N_22084,N_21243,N_21628);
or U22085 (N_22085,N_21966,N_21677);
and U22086 (N_22086,N_21375,N_21471);
nor U22087 (N_22087,N_21382,N_21168);
nor U22088 (N_22088,N_21691,N_21732);
and U22089 (N_22089,N_21149,N_21223);
nor U22090 (N_22090,N_21222,N_21402);
xor U22091 (N_22091,N_21651,N_21085);
or U22092 (N_22092,N_21365,N_21754);
nand U22093 (N_22093,N_21757,N_21977);
nor U22094 (N_22094,N_21950,N_21597);
or U22095 (N_22095,N_21562,N_21571);
xnor U22096 (N_22096,N_21068,N_21304);
or U22097 (N_22097,N_21788,N_21343);
nand U22098 (N_22098,N_21708,N_21393);
nand U22099 (N_22099,N_21000,N_21692);
or U22100 (N_22100,N_21423,N_21032);
nor U22101 (N_22101,N_21680,N_21914);
or U22102 (N_22102,N_21543,N_21138);
nor U22103 (N_22103,N_21741,N_21121);
nand U22104 (N_22104,N_21828,N_21044);
and U22105 (N_22105,N_21855,N_21006);
xnor U22106 (N_22106,N_21712,N_21142);
nor U22107 (N_22107,N_21120,N_21388);
nand U22108 (N_22108,N_21161,N_21864);
xor U22109 (N_22109,N_21895,N_21492);
or U22110 (N_22110,N_21328,N_21408);
or U22111 (N_22111,N_21418,N_21981);
xor U22112 (N_22112,N_21925,N_21720);
and U22113 (N_22113,N_21016,N_21430);
or U22114 (N_22114,N_21852,N_21104);
or U22115 (N_22115,N_21378,N_21226);
xor U22116 (N_22116,N_21716,N_21686);
or U22117 (N_22117,N_21689,N_21959);
nand U22118 (N_22118,N_21461,N_21790);
xnor U22119 (N_22119,N_21719,N_21506);
and U22120 (N_22120,N_21557,N_21774);
nor U22121 (N_22121,N_21389,N_21575);
xor U22122 (N_22122,N_21117,N_21130);
and U22123 (N_22123,N_21879,N_21170);
nor U22124 (N_22124,N_21611,N_21710);
nand U22125 (N_22125,N_21970,N_21979);
nor U22126 (N_22126,N_21025,N_21634);
or U22127 (N_22127,N_21037,N_21797);
nand U22128 (N_22128,N_21723,N_21164);
xnor U22129 (N_22129,N_21605,N_21176);
nand U22130 (N_22130,N_21020,N_21178);
nand U22131 (N_22131,N_21095,N_21949);
nand U22132 (N_22132,N_21435,N_21579);
and U22133 (N_22133,N_21005,N_21824);
xnor U22134 (N_22134,N_21404,N_21901);
or U22135 (N_22135,N_21148,N_21620);
and U22136 (N_22136,N_21919,N_21106);
or U22137 (N_22137,N_21730,N_21335);
xnor U22138 (N_22138,N_21017,N_21345);
nand U22139 (N_22139,N_21572,N_21028);
xnor U22140 (N_22140,N_21364,N_21770);
and U22141 (N_22141,N_21102,N_21745);
xnor U22142 (N_22142,N_21871,N_21729);
or U22143 (N_22143,N_21083,N_21653);
nand U22144 (N_22144,N_21878,N_21891);
xor U22145 (N_22145,N_21606,N_21661);
and U22146 (N_22146,N_21617,N_21491);
or U22147 (N_22147,N_21835,N_21538);
or U22148 (N_22148,N_21237,N_21583);
nor U22149 (N_22149,N_21416,N_21885);
or U22150 (N_22150,N_21474,N_21087);
or U22151 (N_22151,N_21359,N_21853);
xor U22152 (N_22152,N_21822,N_21030);
nor U22153 (N_22153,N_21450,N_21008);
nand U22154 (N_22154,N_21145,N_21726);
xor U22155 (N_22155,N_21446,N_21268);
nor U22156 (N_22156,N_21101,N_21374);
and U22157 (N_22157,N_21334,N_21463);
and U22158 (N_22158,N_21937,N_21569);
and U22159 (N_22159,N_21390,N_21696);
xor U22160 (N_22160,N_21532,N_21175);
and U22161 (N_22161,N_21941,N_21616);
and U22162 (N_22162,N_21330,N_21533);
or U22163 (N_22163,N_21218,N_21978);
and U22164 (N_22164,N_21272,N_21321);
nor U22165 (N_22165,N_21065,N_21433);
nand U22166 (N_22166,N_21307,N_21265);
nor U22167 (N_22167,N_21541,N_21350);
or U22168 (N_22168,N_21863,N_21371);
and U22169 (N_22169,N_21870,N_21267);
nand U22170 (N_22170,N_21787,N_21622);
or U22171 (N_22171,N_21927,N_21399);
or U22172 (N_22172,N_21553,N_21115);
or U22173 (N_22173,N_21080,N_21656);
nand U22174 (N_22174,N_21349,N_21781);
xnor U22175 (N_22175,N_21576,N_21281);
xor U22176 (N_22176,N_21625,N_21257);
or U22177 (N_22177,N_21618,N_21318);
nand U22178 (N_22178,N_21143,N_21315);
xor U22179 (N_22179,N_21889,N_21834);
nor U22180 (N_22180,N_21670,N_21197);
nor U22181 (N_22181,N_21051,N_21015);
nor U22182 (N_22182,N_21733,N_21549);
xor U22183 (N_22183,N_21225,N_21734);
nand U22184 (N_22184,N_21906,N_21573);
xor U22185 (N_22185,N_21998,N_21527);
xnor U22186 (N_22186,N_21439,N_21081);
xor U22187 (N_22187,N_21513,N_21264);
nor U22188 (N_22188,N_21124,N_21854);
or U22189 (N_22189,N_21109,N_21698);
xnor U22190 (N_22190,N_21445,N_21812);
xnor U22191 (N_22191,N_21352,N_21497);
and U22192 (N_22192,N_21132,N_21817);
nor U22193 (N_22193,N_21224,N_21638);
nor U22194 (N_22194,N_21007,N_21487);
nor U22195 (N_22195,N_21690,N_21486);
and U22196 (N_22196,N_21911,N_21184);
xnor U22197 (N_22197,N_21968,N_21410);
or U22198 (N_22198,N_21609,N_21391);
xor U22199 (N_22199,N_21458,N_21744);
nor U22200 (N_22200,N_21275,N_21011);
or U22201 (N_22201,N_21488,N_21512);
nand U22202 (N_22202,N_21910,N_21242);
nor U22203 (N_22203,N_21574,N_21397);
and U22204 (N_22204,N_21921,N_21535);
xnor U22205 (N_22205,N_21839,N_21094);
nand U22206 (N_22206,N_21403,N_21266);
nor U22207 (N_22207,N_21823,N_21381);
nand U22208 (N_22208,N_21479,N_21366);
nand U22209 (N_22209,N_21441,N_21483);
nor U22210 (N_22210,N_21826,N_21485);
xor U22211 (N_22211,N_21507,N_21920);
and U22212 (N_22212,N_21873,N_21146);
xor U22213 (N_22213,N_21200,N_21525);
nor U22214 (N_22214,N_21108,N_21152);
nor U22215 (N_22215,N_21587,N_21666);
nand U22216 (N_22216,N_21783,N_21711);
and U22217 (N_22217,N_21417,N_21260);
nand U22218 (N_22218,N_21155,N_21229);
nand U22219 (N_22219,N_21669,N_21147);
nor U22220 (N_22220,N_21026,N_21807);
nand U22221 (N_22221,N_21985,N_21357);
nor U22222 (N_22222,N_21019,N_21188);
or U22223 (N_22223,N_21704,N_21963);
or U22224 (N_22224,N_21747,N_21988);
or U22225 (N_22225,N_21777,N_21627);
nand U22226 (N_22226,N_21778,N_21624);
and U22227 (N_22227,N_21112,N_21821);
and U22228 (N_22228,N_21073,N_21455);
or U22229 (N_22229,N_21675,N_21457);
or U22230 (N_22230,N_21034,N_21559);
nor U22231 (N_22231,N_21452,N_21362);
nor U22232 (N_22232,N_21681,N_21392);
xnor U22233 (N_22233,N_21989,N_21615);
nand U22234 (N_22234,N_21764,N_21522);
xor U22235 (N_22235,N_21660,N_21516);
xor U22236 (N_22236,N_21961,N_21296);
nand U22237 (N_22237,N_21706,N_21872);
or U22238 (N_22238,N_21619,N_21277);
xor U22239 (N_22239,N_21244,N_21440);
and U22240 (N_22240,N_21255,N_21962);
nand U22241 (N_22241,N_21182,N_21274);
nand U22242 (N_22242,N_21217,N_21684);
or U22243 (N_22243,N_21526,N_21599);
and U22244 (N_22244,N_21097,N_21413);
and U22245 (N_22245,N_21815,N_21763);
nor U22246 (N_22246,N_21674,N_21428);
nor U22247 (N_22247,N_21114,N_21982);
or U22248 (N_22248,N_21449,N_21171);
nor U22249 (N_22249,N_21558,N_21113);
nor U22250 (N_22250,N_21158,N_21216);
or U22251 (N_22251,N_21049,N_21713);
nand U22252 (N_22252,N_21380,N_21056);
xor U22253 (N_22253,N_21111,N_21320);
xnor U22254 (N_22254,N_21603,N_21805);
or U22255 (N_22255,N_21808,N_21776);
xor U22256 (N_22256,N_21768,N_21273);
and U22257 (N_22257,N_21940,N_21276);
or U22258 (N_22258,N_21547,N_21793);
and U22259 (N_22259,N_21876,N_21310);
xnor U22260 (N_22260,N_21151,N_21725);
and U22261 (N_22261,N_21964,N_21088);
xnor U22262 (N_22262,N_21442,N_21183);
nor U22263 (N_22263,N_21031,N_21842);
nand U22264 (N_22264,N_21799,N_21233);
xnor U22265 (N_22265,N_21874,N_21062);
nor U22266 (N_22266,N_21126,N_21067);
or U22267 (N_22267,N_21510,N_21023);
nor U22268 (N_22268,N_21928,N_21705);
and U22269 (N_22269,N_21386,N_21098);
or U22270 (N_22270,N_21070,N_21014);
nand U22271 (N_22271,N_21162,N_21973);
nor U22272 (N_22272,N_21054,N_21633);
and U22273 (N_22273,N_21473,N_21614);
xor U22274 (N_22274,N_21325,N_21971);
nand U22275 (N_22275,N_21086,N_21658);
nor U22276 (N_22276,N_21213,N_21250);
nor U22277 (N_22277,N_21693,N_21379);
nor U22278 (N_22278,N_21827,N_21125);
nand U22279 (N_22279,N_21481,N_21884);
and U22280 (N_22280,N_21230,N_21912);
nor U22281 (N_22281,N_21672,N_21100);
nor U22282 (N_22282,N_21363,N_21795);
or U22283 (N_22283,N_21050,N_21253);
xor U22284 (N_22284,N_21134,N_21294);
nand U22285 (N_22285,N_21536,N_21280);
xnor U22286 (N_22286,N_21247,N_21415);
or U22287 (N_22287,N_21157,N_21857);
or U22288 (N_22288,N_21453,N_21075);
and U22289 (N_22289,N_21012,N_21780);
xor U22290 (N_22290,N_21293,N_21189);
nor U22291 (N_22291,N_21055,N_21122);
and U22292 (N_22292,N_21469,N_21092);
xor U22293 (N_22293,N_21644,N_21256);
and U22294 (N_22294,N_21493,N_21946);
or U22295 (N_22295,N_21849,N_21336);
nand U22296 (N_22296,N_21319,N_21323);
or U22297 (N_22297,N_21632,N_21322);
or U22298 (N_22298,N_21166,N_21983);
nand U22299 (N_22299,N_21235,N_21792);
xor U22300 (N_22300,N_21589,N_21150);
xnor U22301 (N_22301,N_21992,N_21700);
or U22302 (N_22302,N_21317,N_21287);
and U22303 (N_22303,N_21986,N_21245);
and U22304 (N_22304,N_21801,N_21679);
xnor U22305 (N_22305,N_21384,N_21721);
nor U22306 (N_22306,N_21414,N_21898);
nor U22307 (N_22307,N_21172,N_21360);
nor U22308 (N_22308,N_21021,N_21779);
and U22309 (N_22309,N_21459,N_21022);
or U22310 (N_22310,N_21598,N_21246);
and U22311 (N_22311,N_21072,N_21502);
nor U22312 (N_22312,N_21090,N_21156);
and U22313 (N_22313,N_21077,N_21782);
xor U22314 (N_22314,N_21637,N_21995);
or U22315 (N_22315,N_21530,N_21251);
nand U22316 (N_22316,N_21804,N_21649);
nand U22317 (N_22317,N_21903,N_21300);
nand U22318 (N_22318,N_21738,N_21043);
xor U22319 (N_22319,N_21663,N_21231);
nand U22320 (N_22320,N_21369,N_21994);
or U22321 (N_22321,N_21883,N_21717);
or U22322 (N_22322,N_21398,N_21668);
xor U22323 (N_22323,N_21960,N_21942);
or U22324 (N_22324,N_21059,N_21980);
nor U22325 (N_22325,N_21456,N_21238);
nor U22326 (N_22326,N_21975,N_21509);
or U22327 (N_22327,N_21118,N_21775);
or U22328 (N_22328,N_21796,N_21866);
and U22329 (N_22329,N_21869,N_21841);
xor U22330 (N_22330,N_21933,N_21144);
or U22331 (N_22331,N_21240,N_21825);
or U22332 (N_22332,N_21528,N_21953);
and U22333 (N_22333,N_21348,N_21476);
nor U22334 (N_22334,N_21604,N_21652);
and U22335 (N_22335,N_21137,N_21180);
or U22336 (N_22336,N_21875,N_21643);
xor U22337 (N_22337,N_21765,N_21554);
nand U22338 (N_22338,N_21654,N_21412);
or U22339 (N_22339,N_21846,N_21295);
xnor U22340 (N_22340,N_21053,N_21542);
nand U22341 (N_22341,N_21800,N_21009);
nand U22342 (N_22342,N_21116,N_21859);
and U22343 (N_22343,N_21646,N_21565);
nor U22344 (N_22344,N_21291,N_21703);
xor U22345 (N_22345,N_21444,N_21344);
or U22346 (N_22346,N_21210,N_21772);
nand U22347 (N_22347,N_21753,N_21341);
or U22348 (N_22348,N_21484,N_21454);
nor U22349 (N_22349,N_21206,N_21239);
nand U22350 (N_22350,N_21695,N_21353);
nand U22351 (N_22351,N_21909,N_21165);
or U22352 (N_22352,N_21794,N_21974);
and U22353 (N_22353,N_21896,N_21702);
nor U22354 (N_22354,N_21219,N_21018);
and U22355 (N_22355,N_21346,N_21967);
nand U22356 (N_22356,N_21954,N_21377);
nor U22357 (N_22357,N_21917,N_21136);
xnor U22358 (N_22358,N_21523,N_21153);
nand U22359 (N_22359,N_21593,N_21784);
nand U22360 (N_22360,N_21635,N_21736);
or U22361 (N_22361,N_21285,N_21179);
nor U22362 (N_22362,N_21545,N_21582);
nor U22363 (N_22363,N_21924,N_21965);
xnor U22364 (N_22364,N_21313,N_21951);
nand U22365 (N_22365,N_21737,N_21297);
nand U22366 (N_22366,N_21505,N_21685);
nor U22367 (N_22367,N_21071,N_21809);
nor U22368 (N_22368,N_21531,N_21724);
and U22369 (N_22369,N_21836,N_21036);
or U22370 (N_22370,N_21564,N_21972);
nor U22371 (N_22371,N_21990,N_21196);
nor U22372 (N_22372,N_21731,N_21040);
nand U22373 (N_22373,N_21140,N_21845);
or U22374 (N_22374,N_21261,N_21519);
xnor U22375 (N_22375,N_21096,N_21501);
or U22376 (N_22376,N_21607,N_21354);
xnor U22377 (N_22377,N_21177,N_21199);
or U22378 (N_22378,N_21128,N_21740);
nand U22379 (N_22379,N_21387,N_21987);
nor U22380 (N_22380,N_21907,N_21202);
or U22381 (N_22381,N_21791,N_21662);
or U22382 (N_22382,N_21221,N_21079);
nor U22383 (N_22383,N_21004,N_21046);
xor U22384 (N_22384,N_21798,N_21837);
xnor U22385 (N_22385,N_21838,N_21944);
xnor U22386 (N_22386,N_21047,N_21033);
and U22387 (N_22387,N_21831,N_21298);
xnor U22388 (N_22388,N_21588,N_21758);
xor U22389 (N_22389,N_21701,N_21082);
and U22390 (N_22390,N_21451,N_21750);
and U22391 (N_22391,N_21868,N_21326);
and U22392 (N_22392,N_21546,N_21013);
and U22393 (N_22393,N_21029,N_21187);
xor U22394 (N_22394,N_21659,N_21042);
nor U22395 (N_22395,N_21755,N_21814);
xnor U22396 (N_22396,N_21254,N_21918);
and U22397 (N_22397,N_21952,N_21103);
xnor U22398 (N_22398,N_21420,N_21342);
xor U22399 (N_22399,N_21861,N_21596);
nand U22400 (N_22400,N_21110,N_21856);
and U22401 (N_22401,N_21035,N_21305);
nor U22402 (N_22402,N_21893,N_21515);
xor U22403 (N_22403,N_21174,N_21888);
or U22404 (N_22404,N_21312,N_21529);
nor U22405 (N_22405,N_21511,N_21608);
or U22406 (N_22406,N_21540,N_21465);
or U22407 (N_22407,N_21052,N_21882);
xor U22408 (N_22408,N_21880,N_21897);
nand U22409 (N_22409,N_21816,N_21089);
xor U22410 (N_22410,N_21385,N_21847);
and U22411 (N_22411,N_21064,N_21309);
xor U22412 (N_22412,N_21409,N_21329);
xnor U22413 (N_22413,N_21105,N_21976);
nand U22414 (N_22414,N_21566,N_21957);
nand U22415 (N_22415,N_21099,N_21135);
nand U22416 (N_22416,N_21997,N_21405);
nor U22417 (N_22417,N_21010,N_21584);
or U22418 (N_22418,N_21802,N_21829);
xnor U22419 (N_22419,N_21367,N_21347);
or U22420 (N_22420,N_21767,N_21482);
nor U22421 (N_22421,N_21324,N_21722);
xor U22422 (N_22422,N_21612,N_21173);
nor U22423 (N_22423,N_21358,N_21567);
xor U22424 (N_22424,N_21862,N_21735);
xor U22425 (N_22425,N_21429,N_21984);
and U22426 (N_22426,N_21001,N_21926);
or U22427 (N_22427,N_21996,N_21373);
xor U22428 (N_22428,N_21806,N_21204);
or U22429 (N_22429,N_21163,N_21076);
nor U22430 (N_22430,N_21504,N_21048);
nor U22431 (N_22431,N_21211,N_21563);
or U22432 (N_22432,N_21655,N_21057);
and U22433 (N_22433,N_21209,N_21468);
nand U22434 (N_22434,N_21639,N_21288);
nand U22435 (N_22435,N_21560,N_21327);
or U22436 (N_22436,N_21544,N_21537);
and U22437 (N_22437,N_21833,N_21819);
nor U22438 (N_22438,N_21443,N_21601);
nor U22439 (N_22439,N_21292,N_21514);
nand U22440 (N_22440,N_21818,N_21851);
nand U22441 (N_22441,N_21489,N_21636);
and U22442 (N_22442,N_21167,N_21915);
nor U22443 (N_22443,N_21752,N_21850);
and U22444 (N_22444,N_21041,N_21555);
nand U22445 (N_22445,N_21789,N_21715);
and U22446 (N_22446,N_21667,N_21958);
nor U22447 (N_22447,N_21887,N_21930);
nor U22448 (N_22448,N_21436,N_21904);
xor U22449 (N_22449,N_21938,N_21401);
nor U22450 (N_22450,N_21923,N_21259);
nand U22451 (N_22451,N_21743,N_21208);
nand U22452 (N_22452,N_21629,N_21308);
nor U22453 (N_22453,N_21060,N_21518);
nor U22454 (N_22454,N_21697,N_21900);
or U22455 (N_22455,N_21600,N_21556);
nor U22456 (N_22456,N_21045,N_21434);
nor U22457 (N_22457,N_21477,N_21203);
nor U22458 (N_22458,N_21922,N_21227);
and U22459 (N_22459,N_21407,N_21709);
and U22460 (N_22460,N_21419,N_21278);
nor U22461 (N_22461,N_21470,N_21631);
or U22462 (N_22462,N_21699,N_21929);
or U22463 (N_22463,N_21123,N_21207);
and U22464 (N_22464,N_21303,N_21395);
nor U22465 (N_22465,N_21630,N_21215);
or U22466 (N_22466,N_21212,N_21969);
nand U22467 (N_22467,N_21333,N_21355);
nand U22468 (N_22468,N_21524,N_21467);
nor U22469 (N_22469,N_21993,N_21447);
or U22470 (N_22470,N_21190,N_21340);
or U22471 (N_22471,N_21241,N_21820);
or U22472 (N_22472,N_21236,N_21610);
and U22473 (N_22473,N_21074,N_21498);
nor U22474 (N_22474,N_21119,N_21201);
nor U22475 (N_22475,N_21289,N_21406);
nor U22476 (N_22476,N_21263,N_21881);
and U22477 (N_22477,N_21191,N_21368);
nand U22478 (N_22478,N_21561,N_21464);
nand U22479 (N_22479,N_21931,N_21500);
or U22480 (N_22480,N_21139,N_21490);
nand U22481 (N_22481,N_21290,N_21198);
xnor U22482 (N_22482,N_21761,N_21337);
or U22483 (N_22483,N_21688,N_21279);
nand U22484 (N_22484,N_21934,N_21301);
xnor U22485 (N_22485,N_21749,N_21460);
nor U22486 (N_22486,N_21063,N_21078);
nand U22487 (N_22487,N_21038,N_21647);
and U22488 (N_22488,N_21728,N_21913);
nor U22489 (N_22489,N_21762,N_21448);
and U22490 (N_22490,N_21475,N_21069);
nor U22491 (N_22491,N_21613,N_21396);
and U22492 (N_22492,N_21641,N_21314);
nand U22493 (N_22493,N_21539,N_21626);
nor U22494 (N_22494,N_21411,N_21916);
nor U22495 (N_22495,N_21002,N_21039);
and U22496 (N_22496,N_21186,N_21302);
or U22497 (N_22497,N_21948,N_21848);
or U22498 (N_22498,N_21270,N_21945);
nor U22499 (N_22499,N_21503,N_21678);
nor U22500 (N_22500,N_21342,N_21134);
and U22501 (N_22501,N_21023,N_21703);
nand U22502 (N_22502,N_21126,N_21156);
or U22503 (N_22503,N_21006,N_21703);
or U22504 (N_22504,N_21705,N_21717);
nor U22505 (N_22505,N_21766,N_21364);
nor U22506 (N_22506,N_21061,N_21469);
or U22507 (N_22507,N_21217,N_21817);
nand U22508 (N_22508,N_21744,N_21441);
or U22509 (N_22509,N_21914,N_21280);
xor U22510 (N_22510,N_21634,N_21645);
or U22511 (N_22511,N_21605,N_21394);
xnor U22512 (N_22512,N_21537,N_21353);
xor U22513 (N_22513,N_21429,N_21883);
nor U22514 (N_22514,N_21038,N_21251);
and U22515 (N_22515,N_21795,N_21465);
or U22516 (N_22516,N_21913,N_21827);
nor U22517 (N_22517,N_21171,N_21715);
nand U22518 (N_22518,N_21372,N_21020);
nor U22519 (N_22519,N_21999,N_21353);
or U22520 (N_22520,N_21202,N_21018);
nand U22521 (N_22521,N_21674,N_21205);
and U22522 (N_22522,N_21346,N_21778);
nand U22523 (N_22523,N_21366,N_21043);
and U22524 (N_22524,N_21490,N_21323);
or U22525 (N_22525,N_21587,N_21920);
nand U22526 (N_22526,N_21968,N_21574);
or U22527 (N_22527,N_21523,N_21837);
or U22528 (N_22528,N_21410,N_21311);
or U22529 (N_22529,N_21850,N_21576);
or U22530 (N_22530,N_21908,N_21094);
nor U22531 (N_22531,N_21833,N_21610);
and U22532 (N_22532,N_21041,N_21930);
xnor U22533 (N_22533,N_21059,N_21245);
or U22534 (N_22534,N_21459,N_21976);
or U22535 (N_22535,N_21236,N_21053);
or U22536 (N_22536,N_21768,N_21702);
nor U22537 (N_22537,N_21081,N_21730);
and U22538 (N_22538,N_21904,N_21607);
or U22539 (N_22539,N_21279,N_21881);
nand U22540 (N_22540,N_21102,N_21472);
and U22541 (N_22541,N_21089,N_21059);
or U22542 (N_22542,N_21754,N_21639);
xnor U22543 (N_22543,N_21648,N_21869);
nand U22544 (N_22544,N_21930,N_21817);
and U22545 (N_22545,N_21695,N_21588);
or U22546 (N_22546,N_21701,N_21073);
xnor U22547 (N_22547,N_21186,N_21963);
nor U22548 (N_22548,N_21984,N_21863);
nand U22549 (N_22549,N_21335,N_21574);
nand U22550 (N_22550,N_21008,N_21440);
nand U22551 (N_22551,N_21489,N_21618);
or U22552 (N_22552,N_21575,N_21431);
and U22553 (N_22553,N_21823,N_21880);
or U22554 (N_22554,N_21900,N_21842);
xnor U22555 (N_22555,N_21282,N_21310);
nor U22556 (N_22556,N_21472,N_21706);
nor U22557 (N_22557,N_21383,N_21930);
nand U22558 (N_22558,N_21028,N_21759);
xor U22559 (N_22559,N_21561,N_21130);
nand U22560 (N_22560,N_21633,N_21279);
nand U22561 (N_22561,N_21739,N_21336);
nand U22562 (N_22562,N_21802,N_21111);
and U22563 (N_22563,N_21423,N_21230);
and U22564 (N_22564,N_21962,N_21027);
nor U22565 (N_22565,N_21531,N_21791);
nor U22566 (N_22566,N_21409,N_21314);
and U22567 (N_22567,N_21826,N_21863);
xor U22568 (N_22568,N_21002,N_21375);
and U22569 (N_22569,N_21176,N_21046);
nor U22570 (N_22570,N_21068,N_21285);
or U22571 (N_22571,N_21461,N_21595);
or U22572 (N_22572,N_21376,N_21673);
nor U22573 (N_22573,N_21539,N_21637);
and U22574 (N_22574,N_21316,N_21358);
nor U22575 (N_22575,N_21854,N_21327);
xor U22576 (N_22576,N_21293,N_21388);
and U22577 (N_22577,N_21525,N_21238);
and U22578 (N_22578,N_21406,N_21503);
xnor U22579 (N_22579,N_21633,N_21188);
and U22580 (N_22580,N_21263,N_21562);
nor U22581 (N_22581,N_21762,N_21213);
and U22582 (N_22582,N_21796,N_21301);
nor U22583 (N_22583,N_21173,N_21511);
xnor U22584 (N_22584,N_21779,N_21249);
xor U22585 (N_22585,N_21744,N_21676);
or U22586 (N_22586,N_21746,N_21809);
or U22587 (N_22587,N_21853,N_21047);
or U22588 (N_22588,N_21662,N_21278);
nand U22589 (N_22589,N_21455,N_21156);
xnor U22590 (N_22590,N_21496,N_21996);
xor U22591 (N_22591,N_21695,N_21253);
nor U22592 (N_22592,N_21628,N_21271);
or U22593 (N_22593,N_21379,N_21060);
or U22594 (N_22594,N_21936,N_21298);
nor U22595 (N_22595,N_21455,N_21765);
nand U22596 (N_22596,N_21305,N_21091);
xor U22597 (N_22597,N_21610,N_21039);
or U22598 (N_22598,N_21047,N_21217);
xnor U22599 (N_22599,N_21908,N_21963);
and U22600 (N_22600,N_21762,N_21440);
nand U22601 (N_22601,N_21460,N_21103);
xnor U22602 (N_22602,N_21141,N_21159);
nor U22603 (N_22603,N_21506,N_21614);
nor U22604 (N_22604,N_21049,N_21977);
nor U22605 (N_22605,N_21386,N_21993);
or U22606 (N_22606,N_21047,N_21802);
nand U22607 (N_22607,N_21594,N_21670);
nand U22608 (N_22608,N_21822,N_21761);
xnor U22609 (N_22609,N_21586,N_21195);
nand U22610 (N_22610,N_21750,N_21073);
nand U22611 (N_22611,N_21340,N_21427);
and U22612 (N_22612,N_21443,N_21245);
nor U22613 (N_22613,N_21988,N_21236);
or U22614 (N_22614,N_21238,N_21214);
nor U22615 (N_22615,N_21793,N_21177);
xnor U22616 (N_22616,N_21288,N_21525);
or U22617 (N_22617,N_21090,N_21034);
nor U22618 (N_22618,N_21279,N_21617);
nor U22619 (N_22619,N_21478,N_21028);
xnor U22620 (N_22620,N_21251,N_21176);
and U22621 (N_22621,N_21041,N_21697);
nand U22622 (N_22622,N_21996,N_21310);
nand U22623 (N_22623,N_21221,N_21151);
or U22624 (N_22624,N_21195,N_21019);
and U22625 (N_22625,N_21526,N_21623);
or U22626 (N_22626,N_21598,N_21141);
or U22627 (N_22627,N_21340,N_21693);
and U22628 (N_22628,N_21449,N_21104);
and U22629 (N_22629,N_21277,N_21384);
xor U22630 (N_22630,N_21637,N_21697);
xnor U22631 (N_22631,N_21571,N_21422);
or U22632 (N_22632,N_21420,N_21144);
xnor U22633 (N_22633,N_21892,N_21603);
nor U22634 (N_22634,N_21305,N_21400);
or U22635 (N_22635,N_21773,N_21437);
xnor U22636 (N_22636,N_21923,N_21515);
nor U22637 (N_22637,N_21456,N_21399);
nor U22638 (N_22638,N_21882,N_21345);
or U22639 (N_22639,N_21959,N_21217);
or U22640 (N_22640,N_21422,N_21691);
xor U22641 (N_22641,N_21281,N_21660);
and U22642 (N_22642,N_21380,N_21774);
or U22643 (N_22643,N_21773,N_21592);
nor U22644 (N_22644,N_21420,N_21288);
xnor U22645 (N_22645,N_21059,N_21642);
nand U22646 (N_22646,N_21819,N_21611);
and U22647 (N_22647,N_21966,N_21538);
and U22648 (N_22648,N_21409,N_21550);
and U22649 (N_22649,N_21927,N_21086);
nand U22650 (N_22650,N_21048,N_21442);
or U22651 (N_22651,N_21963,N_21182);
nor U22652 (N_22652,N_21222,N_21374);
and U22653 (N_22653,N_21086,N_21321);
or U22654 (N_22654,N_21868,N_21498);
or U22655 (N_22655,N_21907,N_21284);
nor U22656 (N_22656,N_21967,N_21029);
or U22657 (N_22657,N_21885,N_21175);
nor U22658 (N_22658,N_21265,N_21791);
xnor U22659 (N_22659,N_21700,N_21497);
or U22660 (N_22660,N_21735,N_21572);
xor U22661 (N_22661,N_21855,N_21069);
nand U22662 (N_22662,N_21937,N_21097);
or U22663 (N_22663,N_21968,N_21132);
or U22664 (N_22664,N_21836,N_21724);
xnor U22665 (N_22665,N_21602,N_21214);
nor U22666 (N_22666,N_21340,N_21050);
nand U22667 (N_22667,N_21611,N_21297);
nor U22668 (N_22668,N_21869,N_21501);
nor U22669 (N_22669,N_21490,N_21497);
xor U22670 (N_22670,N_21959,N_21749);
or U22671 (N_22671,N_21755,N_21526);
nor U22672 (N_22672,N_21382,N_21391);
and U22673 (N_22673,N_21182,N_21407);
xnor U22674 (N_22674,N_21080,N_21727);
or U22675 (N_22675,N_21718,N_21609);
nor U22676 (N_22676,N_21807,N_21482);
xnor U22677 (N_22677,N_21016,N_21414);
xor U22678 (N_22678,N_21270,N_21653);
nor U22679 (N_22679,N_21574,N_21794);
or U22680 (N_22680,N_21803,N_21036);
nor U22681 (N_22681,N_21381,N_21318);
or U22682 (N_22682,N_21476,N_21964);
and U22683 (N_22683,N_21086,N_21270);
xor U22684 (N_22684,N_21805,N_21043);
nand U22685 (N_22685,N_21419,N_21235);
or U22686 (N_22686,N_21972,N_21639);
or U22687 (N_22687,N_21756,N_21985);
or U22688 (N_22688,N_21346,N_21763);
nor U22689 (N_22689,N_21744,N_21268);
xnor U22690 (N_22690,N_21154,N_21033);
and U22691 (N_22691,N_21877,N_21462);
and U22692 (N_22692,N_21670,N_21639);
and U22693 (N_22693,N_21195,N_21253);
and U22694 (N_22694,N_21604,N_21526);
nand U22695 (N_22695,N_21673,N_21314);
xnor U22696 (N_22696,N_21488,N_21011);
xor U22697 (N_22697,N_21703,N_21759);
nor U22698 (N_22698,N_21496,N_21269);
xor U22699 (N_22699,N_21192,N_21277);
and U22700 (N_22700,N_21651,N_21966);
xor U22701 (N_22701,N_21980,N_21908);
xnor U22702 (N_22702,N_21852,N_21363);
xor U22703 (N_22703,N_21643,N_21001);
or U22704 (N_22704,N_21755,N_21019);
nand U22705 (N_22705,N_21039,N_21673);
and U22706 (N_22706,N_21257,N_21455);
xor U22707 (N_22707,N_21135,N_21422);
or U22708 (N_22708,N_21023,N_21004);
nor U22709 (N_22709,N_21735,N_21340);
xnor U22710 (N_22710,N_21133,N_21325);
and U22711 (N_22711,N_21346,N_21880);
and U22712 (N_22712,N_21014,N_21737);
and U22713 (N_22713,N_21267,N_21989);
or U22714 (N_22714,N_21544,N_21660);
nor U22715 (N_22715,N_21453,N_21477);
xor U22716 (N_22716,N_21798,N_21149);
nand U22717 (N_22717,N_21406,N_21981);
xnor U22718 (N_22718,N_21383,N_21747);
nor U22719 (N_22719,N_21718,N_21540);
or U22720 (N_22720,N_21272,N_21927);
nand U22721 (N_22721,N_21525,N_21971);
nand U22722 (N_22722,N_21197,N_21499);
or U22723 (N_22723,N_21549,N_21421);
and U22724 (N_22724,N_21307,N_21622);
and U22725 (N_22725,N_21212,N_21220);
nand U22726 (N_22726,N_21568,N_21284);
nand U22727 (N_22727,N_21928,N_21731);
nor U22728 (N_22728,N_21908,N_21216);
and U22729 (N_22729,N_21598,N_21452);
and U22730 (N_22730,N_21443,N_21771);
and U22731 (N_22731,N_21269,N_21531);
xor U22732 (N_22732,N_21462,N_21781);
nor U22733 (N_22733,N_21397,N_21570);
or U22734 (N_22734,N_21910,N_21005);
nand U22735 (N_22735,N_21725,N_21271);
or U22736 (N_22736,N_21660,N_21018);
nand U22737 (N_22737,N_21063,N_21048);
or U22738 (N_22738,N_21121,N_21795);
or U22739 (N_22739,N_21174,N_21519);
or U22740 (N_22740,N_21645,N_21370);
nand U22741 (N_22741,N_21542,N_21952);
nor U22742 (N_22742,N_21039,N_21684);
xor U22743 (N_22743,N_21811,N_21499);
nor U22744 (N_22744,N_21566,N_21479);
xor U22745 (N_22745,N_21909,N_21275);
nand U22746 (N_22746,N_21687,N_21600);
or U22747 (N_22747,N_21667,N_21379);
nand U22748 (N_22748,N_21423,N_21623);
or U22749 (N_22749,N_21516,N_21700);
xnor U22750 (N_22750,N_21965,N_21423);
nor U22751 (N_22751,N_21931,N_21696);
xor U22752 (N_22752,N_21693,N_21945);
nand U22753 (N_22753,N_21896,N_21421);
or U22754 (N_22754,N_21224,N_21623);
nand U22755 (N_22755,N_21628,N_21248);
and U22756 (N_22756,N_21256,N_21204);
nor U22757 (N_22757,N_21892,N_21926);
nor U22758 (N_22758,N_21855,N_21180);
or U22759 (N_22759,N_21456,N_21020);
or U22760 (N_22760,N_21605,N_21029);
nor U22761 (N_22761,N_21690,N_21207);
or U22762 (N_22762,N_21154,N_21656);
and U22763 (N_22763,N_21247,N_21922);
and U22764 (N_22764,N_21605,N_21679);
nand U22765 (N_22765,N_21900,N_21714);
and U22766 (N_22766,N_21987,N_21272);
or U22767 (N_22767,N_21738,N_21290);
or U22768 (N_22768,N_21554,N_21342);
or U22769 (N_22769,N_21166,N_21262);
or U22770 (N_22770,N_21439,N_21537);
nand U22771 (N_22771,N_21786,N_21088);
nand U22772 (N_22772,N_21908,N_21264);
and U22773 (N_22773,N_21421,N_21126);
nor U22774 (N_22774,N_21877,N_21212);
xor U22775 (N_22775,N_21824,N_21506);
nor U22776 (N_22776,N_21364,N_21245);
nand U22777 (N_22777,N_21334,N_21298);
or U22778 (N_22778,N_21410,N_21997);
and U22779 (N_22779,N_21643,N_21239);
xnor U22780 (N_22780,N_21024,N_21133);
xor U22781 (N_22781,N_21596,N_21719);
or U22782 (N_22782,N_21454,N_21986);
xnor U22783 (N_22783,N_21328,N_21205);
and U22784 (N_22784,N_21852,N_21618);
xnor U22785 (N_22785,N_21138,N_21570);
nand U22786 (N_22786,N_21092,N_21330);
or U22787 (N_22787,N_21003,N_21521);
and U22788 (N_22788,N_21662,N_21467);
nand U22789 (N_22789,N_21213,N_21581);
nand U22790 (N_22790,N_21663,N_21149);
and U22791 (N_22791,N_21499,N_21128);
nand U22792 (N_22792,N_21331,N_21551);
xor U22793 (N_22793,N_21069,N_21343);
or U22794 (N_22794,N_21502,N_21399);
nand U22795 (N_22795,N_21311,N_21591);
or U22796 (N_22796,N_21011,N_21612);
nor U22797 (N_22797,N_21686,N_21118);
or U22798 (N_22798,N_21595,N_21389);
and U22799 (N_22799,N_21286,N_21637);
nand U22800 (N_22800,N_21344,N_21962);
nand U22801 (N_22801,N_21983,N_21413);
and U22802 (N_22802,N_21558,N_21767);
or U22803 (N_22803,N_21587,N_21506);
and U22804 (N_22804,N_21719,N_21498);
xnor U22805 (N_22805,N_21402,N_21535);
xor U22806 (N_22806,N_21992,N_21039);
xnor U22807 (N_22807,N_21419,N_21729);
or U22808 (N_22808,N_21611,N_21498);
and U22809 (N_22809,N_21783,N_21812);
nor U22810 (N_22810,N_21930,N_21757);
and U22811 (N_22811,N_21057,N_21302);
nand U22812 (N_22812,N_21671,N_21955);
nand U22813 (N_22813,N_21144,N_21779);
nor U22814 (N_22814,N_21775,N_21871);
nor U22815 (N_22815,N_21864,N_21924);
nor U22816 (N_22816,N_21900,N_21370);
xnor U22817 (N_22817,N_21393,N_21940);
nor U22818 (N_22818,N_21438,N_21605);
nand U22819 (N_22819,N_21898,N_21475);
xor U22820 (N_22820,N_21049,N_21012);
or U22821 (N_22821,N_21695,N_21511);
xnor U22822 (N_22822,N_21013,N_21515);
or U22823 (N_22823,N_21273,N_21628);
and U22824 (N_22824,N_21165,N_21276);
nor U22825 (N_22825,N_21955,N_21939);
nor U22826 (N_22826,N_21139,N_21718);
nand U22827 (N_22827,N_21697,N_21653);
xor U22828 (N_22828,N_21390,N_21179);
nand U22829 (N_22829,N_21877,N_21560);
nand U22830 (N_22830,N_21079,N_21608);
nor U22831 (N_22831,N_21893,N_21003);
or U22832 (N_22832,N_21369,N_21783);
or U22833 (N_22833,N_21636,N_21299);
xor U22834 (N_22834,N_21420,N_21681);
or U22835 (N_22835,N_21519,N_21234);
xor U22836 (N_22836,N_21608,N_21307);
and U22837 (N_22837,N_21238,N_21827);
xnor U22838 (N_22838,N_21241,N_21408);
nor U22839 (N_22839,N_21734,N_21162);
or U22840 (N_22840,N_21405,N_21863);
nand U22841 (N_22841,N_21270,N_21039);
xor U22842 (N_22842,N_21310,N_21345);
nand U22843 (N_22843,N_21563,N_21818);
xor U22844 (N_22844,N_21749,N_21655);
nand U22845 (N_22845,N_21168,N_21214);
nor U22846 (N_22846,N_21946,N_21161);
nand U22847 (N_22847,N_21876,N_21840);
nor U22848 (N_22848,N_21034,N_21256);
and U22849 (N_22849,N_21493,N_21318);
nor U22850 (N_22850,N_21650,N_21338);
and U22851 (N_22851,N_21905,N_21062);
and U22852 (N_22852,N_21424,N_21155);
or U22853 (N_22853,N_21541,N_21359);
nand U22854 (N_22854,N_21360,N_21027);
and U22855 (N_22855,N_21512,N_21601);
and U22856 (N_22856,N_21657,N_21838);
or U22857 (N_22857,N_21172,N_21488);
or U22858 (N_22858,N_21799,N_21477);
nor U22859 (N_22859,N_21635,N_21920);
nand U22860 (N_22860,N_21795,N_21329);
nand U22861 (N_22861,N_21617,N_21240);
xor U22862 (N_22862,N_21817,N_21006);
xnor U22863 (N_22863,N_21082,N_21542);
xor U22864 (N_22864,N_21179,N_21698);
and U22865 (N_22865,N_21129,N_21202);
nor U22866 (N_22866,N_21065,N_21522);
or U22867 (N_22867,N_21834,N_21484);
xnor U22868 (N_22868,N_21619,N_21740);
nand U22869 (N_22869,N_21661,N_21393);
nand U22870 (N_22870,N_21580,N_21713);
and U22871 (N_22871,N_21377,N_21173);
xnor U22872 (N_22872,N_21988,N_21170);
nor U22873 (N_22873,N_21047,N_21272);
and U22874 (N_22874,N_21188,N_21090);
nor U22875 (N_22875,N_21729,N_21063);
and U22876 (N_22876,N_21865,N_21072);
nand U22877 (N_22877,N_21884,N_21905);
and U22878 (N_22878,N_21923,N_21002);
nand U22879 (N_22879,N_21654,N_21899);
or U22880 (N_22880,N_21529,N_21742);
xor U22881 (N_22881,N_21379,N_21636);
xnor U22882 (N_22882,N_21705,N_21177);
nand U22883 (N_22883,N_21087,N_21979);
or U22884 (N_22884,N_21498,N_21340);
or U22885 (N_22885,N_21450,N_21682);
xnor U22886 (N_22886,N_21462,N_21637);
and U22887 (N_22887,N_21638,N_21346);
nand U22888 (N_22888,N_21302,N_21377);
or U22889 (N_22889,N_21632,N_21765);
and U22890 (N_22890,N_21090,N_21709);
and U22891 (N_22891,N_21336,N_21546);
or U22892 (N_22892,N_21508,N_21632);
and U22893 (N_22893,N_21491,N_21260);
or U22894 (N_22894,N_21586,N_21827);
and U22895 (N_22895,N_21657,N_21666);
and U22896 (N_22896,N_21540,N_21831);
and U22897 (N_22897,N_21070,N_21032);
or U22898 (N_22898,N_21430,N_21467);
nor U22899 (N_22899,N_21663,N_21988);
nor U22900 (N_22900,N_21782,N_21649);
and U22901 (N_22901,N_21184,N_21659);
xor U22902 (N_22902,N_21603,N_21965);
xor U22903 (N_22903,N_21073,N_21691);
nand U22904 (N_22904,N_21733,N_21569);
or U22905 (N_22905,N_21954,N_21190);
nor U22906 (N_22906,N_21678,N_21037);
xor U22907 (N_22907,N_21560,N_21379);
and U22908 (N_22908,N_21978,N_21364);
xor U22909 (N_22909,N_21423,N_21862);
xor U22910 (N_22910,N_21832,N_21180);
nor U22911 (N_22911,N_21900,N_21417);
nor U22912 (N_22912,N_21193,N_21594);
xnor U22913 (N_22913,N_21930,N_21040);
nor U22914 (N_22914,N_21056,N_21505);
xnor U22915 (N_22915,N_21556,N_21890);
and U22916 (N_22916,N_21258,N_21854);
nor U22917 (N_22917,N_21449,N_21713);
nor U22918 (N_22918,N_21141,N_21266);
and U22919 (N_22919,N_21845,N_21706);
or U22920 (N_22920,N_21199,N_21614);
nor U22921 (N_22921,N_21990,N_21360);
and U22922 (N_22922,N_21823,N_21461);
or U22923 (N_22923,N_21233,N_21870);
xnor U22924 (N_22924,N_21336,N_21753);
nand U22925 (N_22925,N_21559,N_21944);
or U22926 (N_22926,N_21875,N_21832);
xor U22927 (N_22927,N_21720,N_21251);
or U22928 (N_22928,N_21267,N_21353);
nand U22929 (N_22929,N_21383,N_21036);
nand U22930 (N_22930,N_21553,N_21311);
nand U22931 (N_22931,N_21904,N_21567);
nand U22932 (N_22932,N_21548,N_21471);
or U22933 (N_22933,N_21271,N_21793);
and U22934 (N_22934,N_21716,N_21042);
or U22935 (N_22935,N_21926,N_21515);
and U22936 (N_22936,N_21134,N_21743);
and U22937 (N_22937,N_21483,N_21803);
nor U22938 (N_22938,N_21695,N_21123);
or U22939 (N_22939,N_21685,N_21711);
nor U22940 (N_22940,N_21429,N_21160);
xnor U22941 (N_22941,N_21744,N_21516);
xor U22942 (N_22942,N_21007,N_21332);
or U22943 (N_22943,N_21083,N_21273);
or U22944 (N_22944,N_21032,N_21756);
nand U22945 (N_22945,N_21433,N_21817);
xor U22946 (N_22946,N_21727,N_21135);
and U22947 (N_22947,N_21424,N_21616);
nor U22948 (N_22948,N_21526,N_21780);
or U22949 (N_22949,N_21559,N_21569);
and U22950 (N_22950,N_21202,N_21320);
nand U22951 (N_22951,N_21911,N_21382);
xor U22952 (N_22952,N_21067,N_21304);
nand U22953 (N_22953,N_21651,N_21667);
or U22954 (N_22954,N_21003,N_21706);
xor U22955 (N_22955,N_21160,N_21603);
or U22956 (N_22956,N_21261,N_21252);
nand U22957 (N_22957,N_21017,N_21955);
nor U22958 (N_22958,N_21709,N_21328);
and U22959 (N_22959,N_21657,N_21689);
and U22960 (N_22960,N_21965,N_21908);
nor U22961 (N_22961,N_21668,N_21855);
nand U22962 (N_22962,N_21191,N_21661);
and U22963 (N_22963,N_21058,N_21334);
and U22964 (N_22964,N_21042,N_21807);
xnor U22965 (N_22965,N_21875,N_21595);
xnor U22966 (N_22966,N_21586,N_21839);
nor U22967 (N_22967,N_21221,N_21551);
nand U22968 (N_22968,N_21232,N_21717);
or U22969 (N_22969,N_21287,N_21730);
nor U22970 (N_22970,N_21199,N_21229);
nand U22971 (N_22971,N_21618,N_21722);
and U22972 (N_22972,N_21724,N_21043);
nand U22973 (N_22973,N_21417,N_21259);
or U22974 (N_22974,N_21514,N_21249);
nor U22975 (N_22975,N_21885,N_21499);
nand U22976 (N_22976,N_21700,N_21726);
xnor U22977 (N_22977,N_21599,N_21350);
nor U22978 (N_22978,N_21501,N_21789);
xnor U22979 (N_22979,N_21728,N_21499);
xnor U22980 (N_22980,N_21971,N_21367);
or U22981 (N_22981,N_21074,N_21797);
and U22982 (N_22982,N_21725,N_21688);
or U22983 (N_22983,N_21435,N_21899);
and U22984 (N_22984,N_21563,N_21533);
nor U22985 (N_22985,N_21030,N_21795);
and U22986 (N_22986,N_21210,N_21680);
xor U22987 (N_22987,N_21095,N_21418);
and U22988 (N_22988,N_21386,N_21684);
or U22989 (N_22989,N_21317,N_21978);
and U22990 (N_22990,N_21229,N_21448);
nand U22991 (N_22991,N_21463,N_21164);
and U22992 (N_22992,N_21721,N_21574);
or U22993 (N_22993,N_21386,N_21436);
and U22994 (N_22994,N_21548,N_21142);
or U22995 (N_22995,N_21543,N_21773);
and U22996 (N_22996,N_21319,N_21584);
and U22997 (N_22997,N_21649,N_21016);
and U22998 (N_22998,N_21103,N_21547);
or U22999 (N_22999,N_21290,N_21124);
nor U23000 (N_23000,N_22451,N_22707);
xnor U23001 (N_23001,N_22182,N_22852);
nand U23002 (N_23002,N_22299,N_22278);
or U23003 (N_23003,N_22519,N_22241);
xor U23004 (N_23004,N_22592,N_22317);
and U23005 (N_23005,N_22287,N_22889);
nor U23006 (N_23006,N_22552,N_22472);
xnor U23007 (N_23007,N_22234,N_22331);
or U23008 (N_23008,N_22784,N_22746);
xor U23009 (N_23009,N_22673,N_22365);
nor U23010 (N_23010,N_22450,N_22667);
or U23011 (N_23011,N_22052,N_22773);
nor U23012 (N_23012,N_22252,N_22334);
xor U23013 (N_23013,N_22992,N_22612);
and U23014 (N_23014,N_22143,N_22186);
nand U23015 (N_23015,N_22485,N_22113);
or U23016 (N_23016,N_22738,N_22525);
nand U23017 (N_23017,N_22933,N_22879);
xnor U23018 (N_23018,N_22548,N_22610);
nand U23019 (N_23019,N_22649,N_22940);
nor U23020 (N_23020,N_22863,N_22643);
and U23021 (N_23021,N_22513,N_22960);
nor U23022 (N_23022,N_22249,N_22590);
and U23023 (N_23023,N_22953,N_22936);
nand U23024 (N_23024,N_22417,N_22063);
nor U23025 (N_23025,N_22291,N_22016);
and U23026 (N_23026,N_22895,N_22545);
xnor U23027 (N_23027,N_22603,N_22445);
nand U23028 (N_23028,N_22396,N_22532);
xnor U23029 (N_23029,N_22920,N_22616);
xnor U23030 (N_23030,N_22251,N_22981);
and U23031 (N_23031,N_22039,N_22394);
or U23032 (N_23032,N_22235,N_22269);
or U23033 (N_23033,N_22921,N_22661);
and U23034 (N_23034,N_22861,N_22584);
and U23035 (N_23035,N_22801,N_22197);
and U23036 (N_23036,N_22289,N_22680);
or U23037 (N_23037,N_22491,N_22142);
xnor U23038 (N_23038,N_22869,N_22902);
and U23039 (N_23039,N_22218,N_22520);
nand U23040 (N_23040,N_22815,N_22273);
nor U23041 (N_23041,N_22414,N_22596);
nand U23042 (N_23042,N_22553,N_22957);
or U23043 (N_23043,N_22806,N_22792);
or U23044 (N_23044,N_22102,N_22298);
xnor U23045 (N_23045,N_22906,N_22478);
xnor U23046 (N_23046,N_22917,N_22389);
xnor U23047 (N_23047,N_22172,N_22715);
and U23048 (N_23048,N_22604,N_22517);
xnor U23049 (N_23049,N_22506,N_22140);
or U23050 (N_23050,N_22588,N_22132);
nor U23051 (N_23051,N_22338,N_22355);
xor U23052 (N_23052,N_22915,N_22372);
and U23053 (N_23053,N_22352,N_22856);
or U23054 (N_23054,N_22944,N_22217);
nor U23055 (N_23055,N_22483,N_22245);
xnor U23056 (N_23056,N_22911,N_22780);
nand U23057 (N_23057,N_22079,N_22498);
nor U23058 (N_23058,N_22275,N_22373);
nand U23059 (N_23059,N_22475,N_22432);
nor U23060 (N_23060,N_22288,N_22857);
and U23061 (N_23061,N_22510,N_22306);
nor U23062 (N_23062,N_22412,N_22573);
or U23063 (N_23063,N_22630,N_22037);
nor U23064 (N_23064,N_22579,N_22326);
nand U23065 (N_23065,N_22701,N_22810);
nand U23066 (N_23066,N_22121,N_22709);
xor U23067 (N_23067,N_22617,N_22176);
or U23068 (N_23068,N_22729,N_22134);
nand U23069 (N_23069,N_22246,N_22250);
nor U23070 (N_23070,N_22363,N_22758);
and U23071 (N_23071,N_22964,N_22939);
nor U23072 (N_23072,N_22435,N_22750);
and U23073 (N_23073,N_22332,N_22204);
or U23074 (N_23074,N_22319,N_22115);
xnor U23075 (N_23075,N_22832,N_22424);
xnor U23076 (N_23076,N_22350,N_22878);
or U23077 (N_23077,N_22265,N_22382);
xnor U23078 (N_23078,N_22523,N_22112);
and U23079 (N_23079,N_22401,N_22554);
xnor U23080 (N_23080,N_22711,N_22082);
or U23081 (N_23081,N_22117,N_22177);
nor U23082 (N_23082,N_22872,N_22200);
and U23083 (N_23083,N_22871,N_22670);
and U23084 (N_23084,N_22343,N_22515);
and U23085 (N_23085,N_22587,N_22873);
xor U23086 (N_23086,N_22640,N_22668);
nor U23087 (N_23087,N_22422,N_22018);
xor U23088 (N_23088,N_22452,N_22314);
and U23089 (N_23089,N_22034,N_22685);
xor U23090 (N_23090,N_22903,N_22625);
xor U23091 (N_23091,N_22844,N_22629);
or U23092 (N_23092,N_22081,N_22342);
nor U23093 (N_23093,N_22679,N_22221);
or U23094 (N_23094,N_22565,N_22387);
nand U23095 (N_23095,N_22511,N_22371);
xnor U23096 (N_23096,N_22682,N_22279);
nand U23097 (N_23097,N_22473,N_22004);
xor U23098 (N_23098,N_22244,N_22814);
nor U23099 (N_23099,N_22207,N_22222);
nor U23100 (N_23100,N_22173,N_22898);
and U23101 (N_23101,N_22571,N_22985);
nor U23102 (N_23102,N_22691,N_22188);
xor U23103 (N_23103,N_22540,N_22748);
nor U23104 (N_23104,N_22482,N_22829);
or U23105 (N_23105,N_22774,N_22615);
nand U23106 (N_23106,N_22977,N_22875);
or U23107 (N_23107,N_22448,N_22159);
and U23108 (N_23108,N_22533,N_22721);
nor U23109 (N_23109,N_22354,N_22664);
or U23110 (N_23110,N_22516,N_22892);
nand U23111 (N_23111,N_22767,N_22967);
nor U23112 (N_23112,N_22323,N_22837);
nand U23113 (N_23113,N_22083,N_22284);
or U23114 (N_23114,N_22644,N_22613);
nor U23115 (N_23115,N_22194,N_22267);
xor U23116 (N_23116,N_22595,N_22833);
nand U23117 (N_23117,N_22392,N_22524);
and U23118 (N_23118,N_22029,N_22305);
or U23119 (N_23119,N_22805,N_22061);
and U23120 (N_23120,N_22206,N_22700);
and U23121 (N_23121,N_22724,N_22794);
or U23122 (N_23122,N_22986,N_22051);
nor U23123 (N_23123,N_22348,N_22270);
nor U23124 (N_23124,N_22383,N_22202);
or U23125 (N_23125,N_22467,N_22044);
and U23126 (N_23126,N_22901,N_22942);
nand U23127 (N_23127,N_22203,N_22876);
xor U23128 (N_23128,N_22983,N_22544);
or U23129 (N_23129,N_22225,N_22243);
nor U23130 (N_23130,N_22990,N_22699);
xor U23131 (N_23131,N_22340,N_22038);
xnor U23132 (N_23132,N_22858,N_22577);
or U23133 (N_23133,N_22864,N_22555);
nand U23134 (N_23134,N_22219,N_22812);
nor U23135 (N_23135,N_22100,N_22716);
nor U23136 (N_23136,N_22458,N_22656);
xor U23137 (N_23137,N_22961,N_22862);
or U23138 (N_23138,N_22662,N_22349);
or U23139 (N_23139,N_22550,N_22247);
and U23140 (N_23140,N_22639,N_22675);
xnor U23141 (N_23141,N_22431,N_22995);
nor U23142 (N_23142,N_22022,N_22436);
and U23143 (N_23143,N_22786,N_22167);
and U23144 (N_23144,N_22357,N_22549);
and U23145 (N_23145,N_22522,N_22607);
xnor U23146 (N_23146,N_22881,N_22007);
and U23147 (N_23147,N_22280,N_22743);
and U23148 (N_23148,N_22487,N_22798);
or U23149 (N_23149,N_22740,N_22847);
nand U23150 (N_23150,N_22367,N_22120);
nor U23151 (N_23151,N_22341,N_22048);
and U23152 (N_23152,N_22313,N_22170);
nor U23153 (N_23153,N_22058,N_22916);
xor U23154 (N_23154,N_22315,N_22425);
and U23155 (N_23155,N_22228,N_22492);
and U23156 (N_23156,N_22253,N_22440);
nor U23157 (N_23157,N_22133,N_22413);
nor U23158 (N_23158,N_22771,N_22060);
xor U23159 (N_23159,N_22339,N_22518);
and U23160 (N_23160,N_22687,N_22777);
or U23161 (N_23161,N_22766,N_22541);
xnor U23162 (N_23162,N_22276,N_22931);
and U23163 (N_23163,N_22998,N_22379);
and U23164 (N_23164,N_22551,N_22529);
nand U23165 (N_23165,N_22465,N_22697);
or U23166 (N_23166,N_22442,N_22393);
nand U23167 (N_23167,N_22025,N_22226);
nand U23168 (N_23168,N_22975,N_22330);
and U23169 (N_23169,N_22578,N_22293);
and U23170 (N_23170,N_22376,N_22556);
nand U23171 (N_23171,N_22781,N_22528);
xnor U23172 (N_23172,N_22825,N_22180);
or U23173 (N_23173,N_22430,N_22240);
nand U23174 (N_23174,N_22599,N_22468);
nor U23175 (N_23175,N_22073,N_22867);
xnor U23176 (N_23176,N_22375,N_22271);
and U23177 (N_23177,N_22567,N_22659);
nand U23178 (N_23178,N_22110,N_22074);
and U23179 (N_23179,N_22024,N_22131);
nand U23180 (N_23180,N_22166,N_22645);
xnor U23181 (N_23181,N_22347,N_22290);
nor U23182 (N_23182,N_22984,N_22899);
nand U23183 (N_23183,N_22380,N_22793);
and U23184 (N_23184,N_22891,N_22078);
xnor U23185 (N_23185,N_22378,N_22236);
and U23186 (N_23186,N_22160,N_22259);
and U23187 (N_23187,N_22757,N_22500);
nor U23188 (N_23188,N_22502,N_22111);
nand U23189 (N_23189,N_22654,N_22789);
xnor U23190 (N_23190,N_22686,N_22486);
nor U23191 (N_23191,N_22714,N_22481);
or U23192 (N_23192,N_22437,N_22368);
nand U23193 (N_23193,N_22849,N_22614);
nand U23194 (N_23194,N_22185,N_22575);
nor U23195 (N_23195,N_22946,N_22105);
nor U23196 (N_23196,N_22521,N_22324);
xnor U23197 (N_23197,N_22318,N_22859);
nor U23198 (N_23198,N_22304,N_22381);
xor U23199 (N_23199,N_22154,N_22776);
xor U23200 (N_23200,N_22950,N_22606);
or U23201 (N_23201,N_22535,N_22817);
and U23202 (N_23202,N_22433,N_22224);
xor U23203 (N_23203,N_22416,N_22441);
nand U23204 (N_23204,N_22171,N_22333);
xnor U23205 (N_23205,N_22720,N_22469);
or U23206 (N_23206,N_22633,N_22157);
or U23207 (N_23207,N_22609,N_22955);
xor U23208 (N_23208,N_22736,N_22547);
and U23209 (N_23209,N_22734,N_22897);
or U23210 (N_23210,N_22164,N_22091);
and U23211 (N_23211,N_22050,N_22818);
xor U23212 (N_23212,N_22144,N_22890);
nand U23213 (N_23213,N_22665,N_22831);
nor U23214 (N_23214,N_22893,N_22201);
xor U23215 (N_23215,N_22749,N_22512);
or U23216 (N_23216,N_22641,N_22277);
xnor U23217 (N_23217,N_22453,N_22399);
xnor U23218 (N_23218,N_22108,N_22658);
nand U23219 (N_23219,N_22128,N_22621);
nor U23220 (N_23220,N_22395,N_22558);
nor U23221 (N_23221,N_22719,N_22894);
xor U23222 (N_23222,N_22619,N_22669);
xnor U23223 (N_23223,N_22427,N_22356);
or U23224 (N_23224,N_22261,N_22080);
and U23225 (N_23225,N_22796,N_22126);
xnor U23226 (N_23226,N_22183,N_22846);
or U23227 (N_23227,N_22137,N_22257);
nand U23228 (N_23228,N_22912,N_22761);
nand U23229 (N_23229,N_22103,N_22210);
or U23230 (N_23230,N_22148,N_22057);
or U23231 (N_23231,N_22900,N_22001);
nor U23232 (N_23232,N_22969,N_22403);
nand U23233 (N_23233,N_22145,N_22019);
nand U23234 (N_23234,N_22653,N_22098);
or U23235 (N_23235,N_22782,N_22227);
and U23236 (N_23236,N_22426,N_22650);
nand U23237 (N_23237,N_22642,N_22703);
or U23238 (N_23238,N_22747,N_22598);
or U23239 (N_23239,N_22211,N_22149);
and U23240 (N_23240,N_22464,N_22765);
xnor U23241 (N_23241,N_22843,N_22223);
or U23242 (N_23242,N_22914,N_22040);
or U23243 (N_23243,N_22484,N_22260);
or U23244 (N_23244,N_22353,N_22032);
xnor U23245 (N_23245,N_22820,N_22754);
nand U23246 (N_23246,N_22213,N_22772);
or U23247 (N_23247,N_22538,N_22769);
or U23248 (N_23248,N_22527,N_22497);
xnor U23249 (N_23249,N_22647,N_22708);
xnor U23250 (N_23250,N_22042,N_22605);
or U23251 (N_23251,N_22683,N_22735);
and U23252 (N_23252,N_22732,N_22360);
nand U23253 (N_23253,N_22344,N_22193);
nor U23254 (N_23254,N_22991,N_22581);
nor U23255 (N_23255,N_22231,N_22727);
nand U23256 (N_23256,N_22972,N_22646);
and U23257 (N_23257,N_22723,N_22301);
xor U23258 (N_23258,N_22994,N_22657);
nand U23259 (N_23259,N_22945,N_22865);
nor U23260 (N_23260,N_22196,N_22242);
nor U23261 (N_23261,N_22883,N_22043);
xor U23262 (N_23262,N_22281,N_22429);
nor U23263 (N_23263,N_22976,N_22067);
or U23264 (N_23264,N_22884,N_22993);
nand U23265 (N_23265,N_22826,N_22620);
xnor U23266 (N_23266,N_22824,N_22071);
xor U23267 (N_23267,N_22628,N_22263);
nand U23268 (N_23268,N_22119,N_22099);
xnor U23269 (N_23269,N_22704,N_22053);
or U23270 (N_23270,N_22239,N_22327);
nor U23271 (N_23271,N_22006,N_22161);
and U23272 (N_23272,N_22811,N_22070);
xor U23273 (N_23273,N_22493,N_22819);
nand U23274 (N_23274,N_22178,N_22813);
and U23275 (N_23275,N_22233,N_22768);
or U23276 (N_23276,N_22064,N_22123);
nor U23277 (N_23277,N_22854,N_22954);
and U23278 (N_23278,N_22086,N_22681);
or U23279 (N_23279,N_22919,N_22214);
xnor U23280 (N_23280,N_22020,N_22062);
nor U23281 (N_23281,N_22585,N_22479);
xnor U23282 (N_23282,N_22384,N_22733);
and U23283 (N_23283,N_22924,N_22104);
and U23284 (N_23284,N_22179,N_22205);
xnor U23285 (N_23285,N_22329,N_22966);
xnor U23286 (N_23286,N_22054,N_22005);
or U23287 (N_23287,N_22460,N_22335);
or U23288 (N_23288,N_22175,N_22256);
or U23289 (N_23289,N_22787,N_22385);
or U23290 (N_23290,N_22457,N_22778);
xnor U23291 (N_23291,N_22136,N_22415);
xnor U23292 (N_23292,N_22712,N_22096);
xnor U23293 (N_23293,N_22325,N_22965);
nand U23294 (N_23294,N_22952,N_22570);
nor U23295 (N_23295,N_22779,N_22611);
and U23296 (N_23296,N_22107,N_22302);
xnor U23297 (N_23297,N_22138,N_22254);
nor U23298 (N_23298,N_22909,N_22660);
xnor U23299 (N_23299,N_22821,N_22146);
and U23300 (N_23300,N_22866,N_22002);
and U23301 (N_23301,N_22232,N_22560);
xor U23302 (N_23302,N_22803,N_22695);
nand U23303 (N_23303,N_22737,N_22671);
nand U23304 (N_23304,N_22443,N_22122);
nor U23305 (N_23305,N_22359,N_22212);
xor U23306 (N_23306,N_22563,N_22209);
xnor U23307 (N_23307,N_22717,N_22808);
and U23308 (N_23308,N_22690,N_22677);
and U23309 (N_23309,N_22880,N_22021);
or U23310 (N_23310,N_22114,N_22274);
or U23311 (N_23311,N_22809,N_22594);
nand U23312 (N_23312,N_22125,N_22626);
or U23313 (N_23313,N_22853,N_22822);
nor U23314 (N_23314,N_22023,N_22576);
nor U23315 (N_23315,N_22836,N_22030);
nor U23316 (N_23316,N_22495,N_22935);
and U23317 (N_23317,N_22632,N_22835);
or U23318 (N_23318,N_22065,N_22090);
and U23319 (N_23319,N_22739,N_22237);
or U23320 (N_23320,N_22463,N_22461);
xor U23321 (N_23321,N_22566,N_22974);
nand U23322 (N_23322,N_22526,N_22586);
and U23323 (N_23323,N_22195,N_22471);
nor U23324 (N_23324,N_22568,N_22569);
xnor U23325 (N_23325,N_22151,N_22860);
nor U23326 (N_23326,N_22388,N_22168);
nor U23327 (N_23327,N_22141,N_22678);
xor U23328 (N_23328,N_22147,N_22480);
nand U23329 (N_23329,N_22896,N_22802);
nand U23330 (N_23330,N_22447,N_22589);
nor U23331 (N_23331,N_22913,N_22488);
xor U23332 (N_23332,N_22476,N_22593);
nand U23333 (N_23333,N_22085,N_22970);
and U23334 (N_23334,N_22877,N_22602);
nor U23335 (N_23335,N_22390,N_22583);
xnor U23336 (N_23336,N_22013,N_22208);
nand U23337 (N_23337,N_22345,N_22106);
or U23338 (N_23338,N_22907,N_22783);
xnor U23339 (N_23339,N_22351,N_22870);
and U23340 (N_23340,N_22718,N_22885);
nor U23341 (N_23341,N_22937,N_22949);
nand U23342 (N_23342,N_22572,N_22059);
and U23343 (N_23343,N_22742,N_22088);
and U23344 (N_23344,N_22618,N_22165);
nor U23345 (N_23345,N_22910,N_22838);
and U23346 (N_23346,N_22087,N_22189);
xor U23347 (N_23347,N_22655,N_22455);
or U23348 (N_23348,N_22509,N_22474);
nor U23349 (N_23349,N_22597,N_22294);
nor U23350 (N_23350,N_22705,N_22702);
or U23351 (N_23351,N_22676,N_22229);
nand U23352 (N_23352,N_22574,N_22215);
xnor U23353 (N_23353,N_22730,N_22499);
xor U23354 (N_23354,N_22187,N_22850);
or U23355 (N_23355,N_22255,N_22169);
nor U23356 (N_23356,N_22934,N_22109);
or U23357 (N_23357,N_22358,N_22968);
nor U23358 (N_23358,N_22636,N_22366);
nor U23359 (N_23359,N_22046,N_22346);
and U23360 (N_23360,N_22800,N_22364);
or U23361 (N_23361,N_22303,N_22409);
xnor U23362 (N_23362,N_22248,N_22580);
and U23363 (N_23363,N_22726,N_22069);
or U23364 (N_23364,N_22076,N_22423);
or U23365 (N_23365,N_22192,N_22258);
xor U23366 (N_23366,N_22987,N_22694);
and U23367 (N_23367,N_22663,N_22428);
or U23368 (N_23368,N_22674,N_22688);
or U23369 (N_23369,N_22963,N_22887);
nor U23370 (N_23370,N_22047,N_22292);
and U23371 (N_23371,N_22439,N_22421);
nor U23372 (N_23372,N_22198,N_22830);
xor U23373 (N_23373,N_22406,N_22084);
nand U23374 (N_23374,N_22400,N_22490);
xor U23375 (N_23375,N_22851,N_22397);
nand U23376 (N_23376,N_22444,N_22637);
nand U23377 (N_23377,N_22462,N_22028);
xor U23378 (N_23378,N_22066,N_22297);
and U23379 (N_23379,N_22904,N_22055);
xnor U23380 (N_23380,N_22958,N_22710);
and U23381 (N_23381,N_22841,N_22153);
and U23382 (N_23382,N_22300,N_22845);
nand U23383 (N_23383,N_22181,N_22537);
xor U23384 (N_23384,N_22072,N_22504);
nand U23385 (N_23385,N_22941,N_22882);
nand U23386 (N_23386,N_22296,N_22755);
xor U23387 (N_23387,N_22564,N_22932);
xnor U23388 (N_23388,N_22770,N_22557);
and U23389 (N_23389,N_22692,N_22014);
xor U23390 (N_23390,N_22652,N_22948);
and U23391 (N_23391,N_22477,N_22762);
and U23392 (N_23392,N_22316,N_22489);
xor U23393 (N_23393,N_22956,N_22842);
xnor U23394 (N_23394,N_22542,N_22174);
xor U23395 (N_23395,N_22097,N_22404);
or U23396 (N_23396,N_22285,N_22608);
xor U23397 (N_23397,N_22507,N_22622);
nand U23398 (N_23398,N_22698,N_22374);
and U23399 (N_23399,N_22000,N_22760);
or U23400 (N_23400,N_22238,N_22923);
or U23401 (N_23401,N_22418,N_22600);
or U23402 (N_23402,N_22124,N_22635);
nor U23403 (N_23403,N_22828,N_22925);
or U23404 (N_23404,N_22307,N_22264);
nand U23405 (N_23405,N_22756,N_22012);
nand U23406 (N_23406,N_22874,N_22947);
and U23407 (N_23407,N_22503,N_22689);
nor U23408 (N_23408,N_22135,N_22101);
and U23409 (N_23409,N_22158,N_22370);
and U23410 (N_23410,N_22311,N_22927);
nor U23411 (N_23411,N_22283,N_22938);
nor U23412 (N_23412,N_22449,N_22989);
or U23413 (N_23413,N_22731,N_22807);
or U23414 (N_23414,N_22693,N_22411);
and U23415 (N_23415,N_22980,N_22308);
nand U23416 (N_23416,N_22775,N_22713);
xnor U23417 (N_23417,N_22011,N_22268);
xor U23418 (N_23418,N_22790,N_22419);
or U23419 (N_23419,N_22009,N_22785);
nand U23420 (N_23420,N_22184,N_22216);
and U23421 (N_23421,N_22230,N_22591);
or U23422 (N_23422,N_22996,N_22266);
xor U23423 (N_23423,N_22799,N_22272);
nand U23424 (N_23424,N_22926,N_22868);
or U23425 (N_23425,N_22312,N_22156);
nor U23426 (N_23426,N_22118,N_22943);
or U23427 (N_23427,N_22530,N_22505);
nand U23428 (N_23428,N_22666,N_22336);
nand U23429 (N_23429,N_22908,N_22601);
nor U23430 (N_23430,N_22764,N_22139);
nor U23431 (N_23431,N_22706,N_22623);
nand U23432 (N_23432,N_22095,N_22410);
xnor U23433 (N_23433,N_22997,N_22722);
xnor U23434 (N_23434,N_22834,N_22262);
nor U23435 (N_23435,N_22027,N_22973);
nand U23436 (N_23436,N_22041,N_22362);
nor U23437 (N_23437,N_22496,N_22648);
or U23438 (N_23438,N_22797,N_22823);
and U23439 (N_23439,N_22651,N_22928);
and U23440 (N_23440,N_22408,N_22089);
or U23441 (N_23441,N_22988,N_22092);
xnor U23442 (N_23442,N_22446,N_22501);
xor U23443 (N_23443,N_22031,N_22982);
or U23444 (N_23444,N_22631,N_22369);
nor U23445 (N_23445,N_22035,N_22466);
xnor U23446 (N_23446,N_22026,N_22056);
and U23447 (N_23447,N_22816,N_22561);
or U23448 (N_23448,N_22420,N_22220);
and U23449 (N_23449,N_22015,N_22391);
xor U23450 (N_23450,N_22163,N_22150);
and U23451 (N_23451,N_22951,N_22638);
nand U23452 (N_23452,N_22398,N_22155);
or U23453 (N_23453,N_22068,N_22405);
xnor U23454 (N_23454,N_22930,N_22386);
nor U23455 (N_23455,N_22559,N_22546);
nor U23456 (N_23456,N_22978,N_22190);
or U23457 (N_23457,N_22127,N_22840);
or U23458 (N_23458,N_22839,N_22094);
and U23459 (N_23459,N_22804,N_22328);
nor U23460 (N_23460,N_22077,N_22627);
xor U23461 (N_23461,N_22886,N_22337);
xnor U23462 (N_23462,N_22008,N_22434);
nor U23463 (N_23463,N_22116,N_22322);
or U23464 (N_23464,N_22827,N_22959);
nand U23465 (N_23465,N_22045,N_22741);
nand U23466 (N_23466,N_22543,N_22725);
or U23467 (N_23467,N_22407,N_22438);
nand U23468 (N_23468,N_22684,N_22508);
nor U23469 (N_23469,N_22795,N_22017);
and U23470 (N_23470,N_22536,N_22282);
nand U23471 (N_23471,N_22531,N_22752);
nand U23472 (N_23472,N_22562,N_22162);
xnor U23473 (N_23473,N_22791,N_22093);
nand U23474 (N_23474,N_22539,N_22514);
nor U23475 (N_23475,N_22753,N_22494);
nand U23476 (N_23476,N_22075,N_22672);
and U23477 (N_23477,N_22922,N_22763);
and U23478 (N_23478,N_22459,N_22905);
and U23479 (N_23479,N_22788,N_22744);
nand U23480 (N_23480,N_22191,N_22999);
nor U23481 (N_23481,N_22454,N_22152);
nor U23482 (N_23482,N_22848,N_22129);
or U23483 (N_23483,N_22003,N_22010);
nand U23484 (N_23484,N_22130,N_22036);
and U23485 (N_23485,N_22049,N_22402);
or U23486 (N_23486,N_22751,N_22624);
nor U23487 (N_23487,N_22979,N_22310);
nor U23488 (N_23488,N_22470,N_22295);
and U23489 (N_23489,N_22199,N_22534);
nor U23490 (N_23490,N_22286,N_22456);
or U23491 (N_23491,N_22309,N_22759);
or U23492 (N_23492,N_22361,N_22962);
and U23493 (N_23493,N_22971,N_22377);
nand U23494 (N_23494,N_22320,N_22888);
and U23495 (N_23495,N_22634,N_22033);
nand U23496 (N_23496,N_22321,N_22745);
nor U23497 (N_23497,N_22918,N_22582);
nor U23498 (N_23498,N_22728,N_22696);
xor U23499 (N_23499,N_22929,N_22855);
or U23500 (N_23500,N_22850,N_22624);
nor U23501 (N_23501,N_22700,N_22636);
xor U23502 (N_23502,N_22518,N_22571);
and U23503 (N_23503,N_22093,N_22049);
nor U23504 (N_23504,N_22899,N_22544);
xor U23505 (N_23505,N_22672,N_22517);
nor U23506 (N_23506,N_22670,N_22238);
or U23507 (N_23507,N_22237,N_22719);
nand U23508 (N_23508,N_22206,N_22351);
xor U23509 (N_23509,N_22016,N_22784);
nand U23510 (N_23510,N_22731,N_22132);
and U23511 (N_23511,N_22723,N_22228);
nor U23512 (N_23512,N_22852,N_22396);
nand U23513 (N_23513,N_22522,N_22913);
nor U23514 (N_23514,N_22915,N_22483);
nand U23515 (N_23515,N_22343,N_22002);
nand U23516 (N_23516,N_22733,N_22364);
or U23517 (N_23517,N_22614,N_22762);
or U23518 (N_23518,N_22936,N_22512);
nor U23519 (N_23519,N_22471,N_22876);
or U23520 (N_23520,N_22245,N_22162);
nand U23521 (N_23521,N_22592,N_22787);
xnor U23522 (N_23522,N_22750,N_22181);
xor U23523 (N_23523,N_22807,N_22961);
and U23524 (N_23524,N_22031,N_22181);
and U23525 (N_23525,N_22123,N_22101);
xnor U23526 (N_23526,N_22184,N_22985);
nor U23527 (N_23527,N_22744,N_22724);
xor U23528 (N_23528,N_22033,N_22006);
or U23529 (N_23529,N_22532,N_22554);
xnor U23530 (N_23530,N_22083,N_22939);
nor U23531 (N_23531,N_22220,N_22817);
nor U23532 (N_23532,N_22000,N_22926);
xnor U23533 (N_23533,N_22063,N_22036);
and U23534 (N_23534,N_22742,N_22020);
nand U23535 (N_23535,N_22380,N_22915);
nand U23536 (N_23536,N_22176,N_22754);
nor U23537 (N_23537,N_22415,N_22285);
nand U23538 (N_23538,N_22883,N_22742);
or U23539 (N_23539,N_22785,N_22291);
or U23540 (N_23540,N_22698,N_22564);
or U23541 (N_23541,N_22423,N_22601);
or U23542 (N_23542,N_22912,N_22271);
nor U23543 (N_23543,N_22608,N_22647);
and U23544 (N_23544,N_22474,N_22320);
nor U23545 (N_23545,N_22451,N_22509);
nand U23546 (N_23546,N_22068,N_22936);
nor U23547 (N_23547,N_22611,N_22327);
nand U23548 (N_23548,N_22927,N_22118);
nand U23549 (N_23549,N_22622,N_22725);
nand U23550 (N_23550,N_22490,N_22638);
nand U23551 (N_23551,N_22103,N_22595);
and U23552 (N_23552,N_22027,N_22304);
or U23553 (N_23553,N_22504,N_22617);
or U23554 (N_23554,N_22426,N_22448);
nand U23555 (N_23555,N_22611,N_22431);
or U23556 (N_23556,N_22019,N_22685);
nand U23557 (N_23557,N_22054,N_22400);
xor U23558 (N_23558,N_22409,N_22176);
nor U23559 (N_23559,N_22533,N_22751);
and U23560 (N_23560,N_22815,N_22711);
and U23561 (N_23561,N_22130,N_22259);
and U23562 (N_23562,N_22540,N_22143);
and U23563 (N_23563,N_22932,N_22441);
or U23564 (N_23564,N_22291,N_22834);
and U23565 (N_23565,N_22890,N_22237);
nor U23566 (N_23566,N_22413,N_22303);
nand U23567 (N_23567,N_22184,N_22506);
xor U23568 (N_23568,N_22422,N_22712);
nand U23569 (N_23569,N_22051,N_22612);
nand U23570 (N_23570,N_22574,N_22405);
or U23571 (N_23571,N_22905,N_22033);
and U23572 (N_23572,N_22618,N_22084);
xor U23573 (N_23573,N_22580,N_22174);
nand U23574 (N_23574,N_22497,N_22942);
and U23575 (N_23575,N_22377,N_22072);
nor U23576 (N_23576,N_22964,N_22859);
nor U23577 (N_23577,N_22917,N_22299);
nand U23578 (N_23578,N_22298,N_22168);
nor U23579 (N_23579,N_22313,N_22269);
and U23580 (N_23580,N_22434,N_22700);
or U23581 (N_23581,N_22758,N_22656);
nor U23582 (N_23582,N_22779,N_22716);
and U23583 (N_23583,N_22225,N_22247);
or U23584 (N_23584,N_22413,N_22189);
nor U23585 (N_23585,N_22477,N_22741);
nand U23586 (N_23586,N_22428,N_22170);
nor U23587 (N_23587,N_22285,N_22863);
or U23588 (N_23588,N_22562,N_22038);
xnor U23589 (N_23589,N_22571,N_22617);
nand U23590 (N_23590,N_22692,N_22327);
and U23591 (N_23591,N_22530,N_22376);
and U23592 (N_23592,N_22634,N_22088);
nor U23593 (N_23593,N_22098,N_22732);
nand U23594 (N_23594,N_22171,N_22855);
nand U23595 (N_23595,N_22208,N_22188);
nand U23596 (N_23596,N_22899,N_22658);
nand U23597 (N_23597,N_22661,N_22940);
and U23598 (N_23598,N_22316,N_22235);
xor U23599 (N_23599,N_22063,N_22945);
xor U23600 (N_23600,N_22096,N_22947);
nand U23601 (N_23601,N_22465,N_22332);
nor U23602 (N_23602,N_22930,N_22238);
or U23603 (N_23603,N_22115,N_22934);
nor U23604 (N_23604,N_22345,N_22363);
or U23605 (N_23605,N_22331,N_22814);
nor U23606 (N_23606,N_22942,N_22074);
nor U23607 (N_23607,N_22634,N_22563);
nand U23608 (N_23608,N_22598,N_22118);
or U23609 (N_23609,N_22085,N_22095);
nand U23610 (N_23610,N_22165,N_22198);
xor U23611 (N_23611,N_22128,N_22115);
nor U23612 (N_23612,N_22137,N_22542);
and U23613 (N_23613,N_22622,N_22317);
nand U23614 (N_23614,N_22862,N_22037);
xnor U23615 (N_23615,N_22652,N_22939);
xor U23616 (N_23616,N_22100,N_22726);
or U23617 (N_23617,N_22809,N_22113);
xnor U23618 (N_23618,N_22820,N_22243);
nand U23619 (N_23619,N_22070,N_22258);
nand U23620 (N_23620,N_22975,N_22448);
and U23621 (N_23621,N_22035,N_22336);
xnor U23622 (N_23622,N_22823,N_22124);
and U23623 (N_23623,N_22532,N_22501);
nand U23624 (N_23624,N_22494,N_22465);
and U23625 (N_23625,N_22047,N_22615);
nand U23626 (N_23626,N_22521,N_22499);
or U23627 (N_23627,N_22795,N_22253);
and U23628 (N_23628,N_22717,N_22066);
nand U23629 (N_23629,N_22058,N_22078);
nor U23630 (N_23630,N_22716,N_22568);
or U23631 (N_23631,N_22735,N_22707);
nand U23632 (N_23632,N_22937,N_22440);
or U23633 (N_23633,N_22877,N_22366);
xor U23634 (N_23634,N_22819,N_22453);
nand U23635 (N_23635,N_22147,N_22626);
nor U23636 (N_23636,N_22108,N_22315);
nor U23637 (N_23637,N_22498,N_22887);
nand U23638 (N_23638,N_22878,N_22759);
and U23639 (N_23639,N_22254,N_22188);
xor U23640 (N_23640,N_22562,N_22541);
or U23641 (N_23641,N_22132,N_22737);
or U23642 (N_23642,N_22923,N_22585);
nor U23643 (N_23643,N_22137,N_22012);
and U23644 (N_23644,N_22491,N_22472);
nor U23645 (N_23645,N_22893,N_22034);
nor U23646 (N_23646,N_22745,N_22445);
nor U23647 (N_23647,N_22047,N_22298);
xor U23648 (N_23648,N_22452,N_22261);
or U23649 (N_23649,N_22553,N_22385);
and U23650 (N_23650,N_22754,N_22569);
and U23651 (N_23651,N_22902,N_22205);
and U23652 (N_23652,N_22734,N_22872);
xor U23653 (N_23653,N_22902,N_22697);
or U23654 (N_23654,N_22074,N_22430);
xor U23655 (N_23655,N_22734,N_22955);
nand U23656 (N_23656,N_22695,N_22737);
nand U23657 (N_23657,N_22180,N_22382);
nand U23658 (N_23658,N_22523,N_22294);
or U23659 (N_23659,N_22041,N_22782);
or U23660 (N_23660,N_22727,N_22425);
nand U23661 (N_23661,N_22504,N_22877);
nand U23662 (N_23662,N_22072,N_22170);
nand U23663 (N_23663,N_22517,N_22649);
and U23664 (N_23664,N_22833,N_22082);
and U23665 (N_23665,N_22421,N_22442);
and U23666 (N_23666,N_22207,N_22737);
nor U23667 (N_23667,N_22044,N_22025);
nand U23668 (N_23668,N_22299,N_22378);
nor U23669 (N_23669,N_22335,N_22542);
or U23670 (N_23670,N_22543,N_22567);
nand U23671 (N_23671,N_22250,N_22298);
nand U23672 (N_23672,N_22078,N_22497);
xnor U23673 (N_23673,N_22538,N_22724);
xor U23674 (N_23674,N_22893,N_22089);
or U23675 (N_23675,N_22954,N_22862);
nor U23676 (N_23676,N_22294,N_22459);
and U23677 (N_23677,N_22697,N_22481);
or U23678 (N_23678,N_22837,N_22737);
and U23679 (N_23679,N_22095,N_22760);
xnor U23680 (N_23680,N_22396,N_22518);
nor U23681 (N_23681,N_22455,N_22358);
nor U23682 (N_23682,N_22589,N_22010);
nand U23683 (N_23683,N_22836,N_22289);
nor U23684 (N_23684,N_22555,N_22611);
nor U23685 (N_23685,N_22460,N_22431);
nor U23686 (N_23686,N_22443,N_22156);
or U23687 (N_23687,N_22375,N_22627);
or U23688 (N_23688,N_22987,N_22312);
nor U23689 (N_23689,N_22400,N_22339);
or U23690 (N_23690,N_22789,N_22328);
xor U23691 (N_23691,N_22654,N_22772);
or U23692 (N_23692,N_22779,N_22980);
nand U23693 (N_23693,N_22191,N_22765);
or U23694 (N_23694,N_22924,N_22178);
xor U23695 (N_23695,N_22264,N_22256);
xor U23696 (N_23696,N_22434,N_22608);
xnor U23697 (N_23697,N_22694,N_22222);
xnor U23698 (N_23698,N_22437,N_22894);
nand U23699 (N_23699,N_22010,N_22077);
or U23700 (N_23700,N_22007,N_22661);
nand U23701 (N_23701,N_22714,N_22514);
and U23702 (N_23702,N_22858,N_22277);
nand U23703 (N_23703,N_22518,N_22419);
nor U23704 (N_23704,N_22017,N_22362);
xor U23705 (N_23705,N_22162,N_22422);
nand U23706 (N_23706,N_22467,N_22726);
nor U23707 (N_23707,N_22697,N_22991);
nor U23708 (N_23708,N_22471,N_22371);
and U23709 (N_23709,N_22520,N_22680);
and U23710 (N_23710,N_22355,N_22267);
and U23711 (N_23711,N_22961,N_22398);
and U23712 (N_23712,N_22339,N_22072);
xnor U23713 (N_23713,N_22776,N_22559);
or U23714 (N_23714,N_22834,N_22050);
nand U23715 (N_23715,N_22024,N_22629);
and U23716 (N_23716,N_22237,N_22335);
xor U23717 (N_23717,N_22528,N_22337);
xnor U23718 (N_23718,N_22333,N_22298);
or U23719 (N_23719,N_22228,N_22445);
nand U23720 (N_23720,N_22613,N_22481);
nor U23721 (N_23721,N_22305,N_22989);
nand U23722 (N_23722,N_22516,N_22398);
nor U23723 (N_23723,N_22824,N_22375);
and U23724 (N_23724,N_22273,N_22328);
and U23725 (N_23725,N_22820,N_22370);
nor U23726 (N_23726,N_22713,N_22491);
nand U23727 (N_23727,N_22306,N_22469);
or U23728 (N_23728,N_22733,N_22159);
xnor U23729 (N_23729,N_22799,N_22709);
xnor U23730 (N_23730,N_22679,N_22848);
nand U23731 (N_23731,N_22947,N_22076);
or U23732 (N_23732,N_22322,N_22911);
nor U23733 (N_23733,N_22933,N_22158);
nand U23734 (N_23734,N_22126,N_22025);
or U23735 (N_23735,N_22035,N_22371);
nand U23736 (N_23736,N_22888,N_22005);
nor U23737 (N_23737,N_22949,N_22288);
nor U23738 (N_23738,N_22377,N_22849);
and U23739 (N_23739,N_22784,N_22994);
xnor U23740 (N_23740,N_22405,N_22494);
or U23741 (N_23741,N_22083,N_22848);
nand U23742 (N_23742,N_22572,N_22429);
xor U23743 (N_23743,N_22787,N_22473);
xor U23744 (N_23744,N_22287,N_22280);
and U23745 (N_23745,N_22413,N_22851);
xnor U23746 (N_23746,N_22444,N_22552);
and U23747 (N_23747,N_22696,N_22318);
or U23748 (N_23748,N_22385,N_22393);
or U23749 (N_23749,N_22942,N_22713);
and U23750 (N_23750,N_22921,N_22417);
and U23751 (N_23751,N_22944,N_22090);
xnor U23752 (N_23752,N_22481,N_22006);
or U23753 (N_23753,N_22153,N_22688);
or U23754 (N_23754,N_22519,N_22540);
nor U23755 (N_23755,N_22134,N_22229);
xor U23756 (N_23756,N_22814,N_22135);
and U23757 (N_23757,N_22843,N_22821);
or U23758 (N_23758,N_22783,N_22855);
and U23759 (N_23759,N_22122,N_22881);
or U23760 (N_23760,N_22603,N_22486);
nand U23761 (N_23761,N_22306,N_22066);
or U23762 (N_23762,N_22767,N_22108);
and U23763 (N_23763,N_22771,N_22312);
xnor U23764 (N_23764,N_22975,N_22721);
nor U23765 (N_23765,N_22548,N_22191);
nand U23766 (N_23766,N_22830,N_22306);
or U23767 (N_23767,N_22241,N_22878);
nand U23768 (N_23768,N_22501,N_22893);
or U23769 (N_23769,N_22452,N_22372);
and U23770 (N_23770,N_22182,N_22539);
nand U23771 (N_23771,N_22031,N_22926);
nor U23772 (N_23772,N_22035,N_22734);
and U23773 (N_23773,N_22602,N_22939);
xnor U23774 (N_23774,N_22391,N_22217);
nand U23775 (N_23775,N_22169,N_22092);
nand U23776 (N_23776,N_22850,N_22675);
or U23777 (N_23777,N_22134,N_22904);
and U23778 (N_23778,N_22064,N_22054);
xor U23779 (N_23779,N_22972,N_22501);
and U23780 (N_23780,N_22720,N_22384);
or U23781 (N_23781,N_22644,N_22612);
nor U23782 (N_23782,N_22715,N_22122);
or U23783 (N_23783,N_22167,N_22947);
or U23784 (N_23784,N_22874,N_22000);
and U23785 (N_23785,N_22767,N_22549);
xor U23786 (N_23786,N_22698,N_22485);
xnor U23787 (N_23787,N_22968,N_22858);
and U23788 (N_23788,N_22654,N_22457);
xnor U23789 (N_23789,N_22022,N_22718);
and U23790 (N_23790,N_22037,N_22613);
nor U23791 (N_23791,N_22898,N_22294);
and U23792 (N_23792,N_22706,N_22725);
xnor U23793 (N_23793,N_22702,N_22611);
or U23794 (N_23794,N_22485,N_22734);
xor U23795 (N_23795,N_22374,N_22210);
nor U23796 (N_23796,N_22438,N_22685);
nor U23797 (N_23797,N_22599,N_22311);
or U23798 (N_23798,N_22118,N_22661);
nor U23799 (N_23799,N_22399,N_22999);
xnor U23800 (N_23800,N_22127,N_22204);
or U23801 (N_23801,N_22077,N_22822);
and U23802 (N_23802,N_22431,N_22548);
xor U23803 (N_23803,N_22152,N_22495);
and U23804 (N_23804,N_22075,N_22271);
and U23805 (N_23805,N_22568,N_22939);
or U23806 (N_23806,N_22832,N_22722);
xor U23807 (N_23807,N_22348,N_22066);
nand U23808 (N_23808,N_22824,N_22904);
and U23809 (N_23809,N_22190,N_22770);
nand U23810 (N_23810,N_22434,N_22064);
and U23811 (N_23811,N_22498,N_22038);
xnor U23812 (N_23812,N_22889,N_22597);
xor U23813 (N_23813,N_22614,N_22230);
xnor U23814 (N_23814,N_22047,N_22012);
nand U23815 (N_23815,N_22461,N_22636);
and U23816 (N_23816,N_22137,N_22237);
or U23817 (N_23817,N_22170,N_22761);
or U23818 (N_23818,N_22985,N_22781);
nand U23819 (N_23819,N_22644,N_22451);
and U23820 (N_23820,N_22148,N_22795);
and U23821 (N_23821,N_22366,N_22794);
or U23822 (N_23822,N_22274,N_22021);
or U23823 (N_23823,N_22988,N_22741);
nor U23824 (N_23824,N_22435,N_22504);
nand U23825 (N_23825,N_22900,N_22292);
and U23826 (N_23826,N_22121,N_22105);
or U23827 (N_23827,N_22203,N_22464);
or U23828 (N_23828,N_22561,N_22262);
nor U23829 (N_23829,N_22613,N_22264);
nor U23830 (N_23830,N_22183,N_22450);
nand U23831 (N_23831,N_22715,N_22757);
xnor U23832 (N_23832,N_22391,N_22333);
xor U23833 (N_23833,N_22468,N_22914);
nand U23834 (N_23834,N_22256,N_22199);
nand U23835 (N_23835,N_22878,N_22880);
xor U23836 (N_23836,N_22585,N_22073);
and U23837 (N_23837,N_22012,N_22782);
xor U23838 (N_23838,N_22946,N_22418);
or U23839 (N_23839,N_22083,N_22241);
or U23840 (N_23840,N_22253,N_22750);
or U23841 (N_23841,N_22927,N_22617);
nand U23842 (N_23842,N_22768,N_22720);
xor U23843 (N_23843,N_22760,N_22661);
and U23844 (N_23844,N_22380,N_22415);
nor U23845 (N_23845,N_22824,N_22976);
nor U23846 (N_23846,N_22715,N_22727);
xor U23847 (N_23847,N_22376,N_22754);
nor U23848 (N_23848,N_22179,N_22789);
nand U23849 (N_23849,N_22274,N_22850);
or U23850 (N_23850,N_22521,N_22932);
xnor U23851 (N_23851,N_22637,N_22238);
nor U23852 (N_23852,N_22498,N_22082);
or U23853 (N_23853,N_22606,N_22139);
xnor U23854 (N_23854,N_22419,N_22114);
and U23855 (N_23855,N_22078,N_22085);
or U23856 (N_23856,N_22067,N_22215);
and U23857 (N_23857,N_22794,N_22424);
or U23858 (N_23858,N_22547,N_22464);
and U23859 (N_23859,N_22705,N_22979);
or U23860 (N_23860,N_22836,N_22505);
nand U23861 (N_23861,N_22645,N_22210);
nand U23862 (N_23862,N_22567,N_22828);
nor U23863 (N_23863,N_22201,N_22608);
xor U23864 (N_23864,N_22041,N_22487);
and U23865 (N_23865,N_22427,N_22199);
and U23866 (N_23866,N_22533,N_22261);
nand U23867 (N_23867,N_22604,N_22713);
nand U23868 (N_23868,N_22210,N_22974);
xor U23869 (N_23869,N_22131,N_22142);
nor U23870 (N_23870,N_22747,N_22229);
or U23871 (N_23871,N_22565,N_22025);
and U23872 (N_23872,N_22172,N_22307);
nand U23873 (N_23873,N_22100,N_22934);
nor U23874 (N_23874,N_22183,N_22350);
xnor U23875 (N_23875,N_22920,N_22590);
nor U23876 (N_23876,N_22893,N_22314);
and U23877 (N_23877,N_22664,N_22431);
nor U23878 (N_23878,N_22552,N_22081);
nand U23879 (N_23879,N_22448,N_22780);
xor U23880 (N_23880,N_22898,N_22657);
nand U23881 (N_23881,N_22478,N_22473);
and U23882 (N_23882,N_22473,N_22098);
nand U23883 (N_23883,N_22813,N_22235);
or U23884 (N_23884,N_22425,N_22714);
nand U23885 (N_23885,N_22531,N_22116);
and U23886 (N_23886,N_22030,N_22207);
nor U23887 (N_23887,N_22308,N_22607);
or U23888 (N_23888,N_22494,N_22726);
xnor U23889 (N_23889,N_22725,N_22204);
or U23890 (N_23890,N_22347,N_22559);
nor U23891 (N_23891,N_22109,N_22523);
or U23892 (N_23892,N_22390,N_22290);
nand U23893 (N_23893,N_22853,N_22130);
xor U23894 (N_23894,N_22870,N_22480);
nor U23895 (N_23895,N_22923,N_22789);
and U23896 (N_23896,N_22930,N_22978);
or U23897 (N_23897,N_22778,N_22075);
or U23898 (N_23898,N_22231,N_22278);
nor U23899 (N_23899,N_22035,N_22984);
or U23900 (N_23900,N_22468,N_22947);
xnor U23901 (N_23901,N_22749,N_22651);
nand U23902 (N_23902,N_22881,N_22282);
or U23903 (N_23903,N_22648,N_22235);
nand U23904 (N_23904,N_22956,N_22322);
nand U23905 (N_23905,N_22142,N_22903);
xnor U23906 (N_23906,N_22704,N_22049);
nand U23907 (N_23907,N_22342,N_22614);
nor U23908 (N_23908,N_22537,N_22031);
or U23909 (N_23909,N_22241,N_22147);
nand U23910 (N_23910,N_22981,N_22740);
and U23911 (N_23911,N_22343,N_22863);
or U23912 (N_23912,N_22098,N_22812);
or U23913 (N_23913,N_22060,N_22844);
nand U23914 (N_23914,N_22642,N_22440);
or U23915 (N_23915,N_22766,N_22907);
xor U23916 (N_23916,N_22696,N_22028);
xor U23917 (N_23917,N_22320,N_22948);
nor U23918 (N_23918,N_22046,N_22503);
and U23919 (N_23919,N_22883,N_22268);
nor U23920 (N_23920,N_22900,N_22195);
nand U23921 (N_23921,N_22598,N_22066);
xnor U23922 (N_23922,N_22511,N_22875);
and U23923 (N_23923,N_22749,N_22562);
or U23924 (N_23924,N_22197,N_22257);
nand U23925 (N_23925,N_22963,N_22158);
xor U23926 (N_23926,N_22420,N_22783);
or U23927 (N_23927,N_22076,N_22387);
or U23928 (N_23928,N_22785,N_22077);
or U23929 (N_23929,N_22908,N_22857);
or U23930 (N_23930,N_22675,N_22024);
or U23931 (N_23931,N_22461,N_22774);
nand U23932 (N_23932,N_22687,N_22205);
xnor U23933 (N_23933,N_22866,N_22550);
xnor U23934 (N_23934,N_22208,N_22103);
or U23935 (N_23935,N_22205,N_22647);
or U23936 (N_23936,N_22174,N_22295);
xnor U23937 (N_23937,N_22169,N_22071);
xor U23938 (N_23938,N_22513,N_22402);
or U23939 (N_23939,N_22485,N_22740);
xor U23940 (N_23940,N_22073,N_22862);
nand U23941 (N_23941,N_22702,N_22737);
or U23942 (N_23942,N_22852,N_22567);
nand U23943 (N_23943,N_22944,N_22271);
and U23944 (N_23944,N_22135,N_22833);
and U23945 (N_23945,N_22509,N_22351);
or U23946 (N_23946,N_22303,N_22051);
nand U23947 (N_23947,N_22940,N_22079);
and U23948 (N_23948,N_22244,N_22985);
nor U23949 (N_23949,N_22275,N_22023);
xor U23950 (N_23950,N_22887,N_22113);
nand U23951 (N_23951,N_22280,N_22376);
and U23952 (N_23952,N_22211,N_22592);
nand U23953 (N_23953,N_22585,N_22217);
and U23954 (N_23954,N_22189,N_22076);
nor U23955 (N_23955,N_22949,N_22729);
or U23956 (N_23956,N_22800,N_22528);
nor U23957 (N_23957,N_22690,N_22591);
or U23958 (N_23958,N_22733,N_22782);
or U23959 (N_23959,N_22663,N_22445);
xnor U23960 (N_23960,N_22827,N_22635);
or U23961 (N_23961,N_22567,N_22386);
or U23962 (N_23962,N_22477,N_22545);
nor U23963 (N_23963,N_22874,N_22978);
nor U23964 (N_23964,N_22014,N_22288);
nor U23965 (N_23965,N_22164,N_22962);
nand U23966 (N_23966,N_22130,N_22093);
nor U23967 (N_23967,N_22353,N_22104);
nand U23968 (N_23968,N_22500,N_22524);
xnor U23969 (N_23969,N_22935,N_22672);
or U23970 (N_23970,N_22310,N_22788);
nand U23971 (N_23971,N_22964,N_22358);
nand U23972 (N_23972,N_22424,N_22967);
or U23973 (N_23973,N_22019,N_22175);
nand U23974 (N_23974,N_22093,N_22023);
nor U23975 (N_23975,N_22414,N_22171);
xnor U23976 (N_23976,N_22915,N_22263);
nand U23977 (N_23977,N_22382,N_22866);
nor U23978 (N_23978,N_22149,N_22441);
nand U23979 (N_23979,N_22113,N_22816);
nor U23980 (N_23980,N_22052,N_22574);
and U23981 (N_23981,N_22952,N_22004);
and U23982 (N_23982,N_22195,N_22627);
xnor U23983 (N_23983,N_22944,N_22049);
and U23984 (N_23984,N_22054,N_22188);
nand U23985 (N_23985,N_22418,N_22141);
nor U23986 (N_23986,N_22054,N_22607);
nor U23987 (N_23987,N_22433,N_22894);
and U23988 (N_23988,N_22736,N_22729);
nand U23989 (N_23989,N_22959,N_22126);
nor U23990 (N_23990,N_22143,N_22969);
nand U23991 (N_23991,N_22351,N_22750);
nor U23992 (N_23992,N_22598,N_22022);
and U23993 (N_23993,N_22129,N_22822);
nor U23994 (N_23994,N_22135,N_22085);
or U23995 (N_23995,N_22967,N_22630);
nor U23996 (N_23996,N_22275,N_22968);
nor U23997 (N_23997,N_22040,N_22860);
or U23998 (N_23998,N_22207,N_22660);
nand U23999 (N_23999,N_22931,N_22470);
nor U24000 (N_24000,N_23737,N_23118);
and U24001 (N_24001,N_23441,N_23784);
nand U24002 (N_24002,N_23738,N_23448);
and U24003 (N_24003,N_23342,N_23755);
xnor U24004 (N_24004,N_23111,N_23821);
nor U24005 (N_24005,N_23829,N_23485);
and U24006 (N_24006,N_23003,N_23418);
and U24007 (N_24007,N_23474,N_23202);
or U24008 (N_24008,N_23772,N_23084);
or U24009 (N_24009,N_23219,N_23692);
or U24010 (N_24010,N_23497,N_23181);
or U24011 (N_24011,N_23580,N_23892);
xor U24012 (N_24012,N_23421,N_23152);
nor U24013 (N_24013,N_23798,N_23088);
xnor U24014 (N_24014,N_23944,N_23843);
nand U24015 (N_24015,N_23036,N_23895);
xnor U24016 (N_24016,N_23354,N_23482);
and U24017 (N_24017,N_23980,N_23248);
and U24018 (N_24018,N_23365,N_23570);
and U24019 (N_24019,N_23067,N_23246);
nor U24020 (N_24020,N_23020,N_23536);
nand U24021 (N_24021,N_23483,N_23982);
and U24022 (N_24022,N_23484,N_23591);
nor U24023 (N_24023,N_23688,N_23573);
or U24024 (N_24024,N_23925,N_23142);
or U24025 (N_24025,N_23024,N_23263);
or U24026 (N_24026,N_23489,N_23782);
or U24027 (N_24027,N_23742,N_23693);
nor U24028 (N_24028,N_23956,N_23463);
nand U24029 (N_24029,N_23454,N_23333);
and U24030 (N_24030,N_23958,N_23222);
nor U24031 (N_24031,N_23093,N_23502);
nand U24032 (N_24032,N_23274,N_23596);
xnor U24033 (N_24033,N_23066,N_23861);
xnor U24034 (N_24034,N_23962,N_23227);
nor U24035 (N_24035,N_23240,N_23694);
xor U24036 (N_24036,N_23718,N_23286);
nor U24037 (N_24037,N_23432,N_23594);
xor U24038 (N_24038,N_23607,N_23823);
nand U24039 (N_24039,N_23252,N_23385);
nor U24040 (N_24040,N_23882,N_23458);
nor U24041 (N_24041,N_23178,N_23309);
and U24042 (N_24042,N_23667,N_23623);
nor U24043 (N_24043,N_23731,N_23068);
or U24044 (N_24044,N_23883,N_23700);
nand U24045 (N_24045,N_23087,N_23964);
nand U24046 (N_24046,N_23409,N_23563);
nor U24047 (N_24047,N_23059,N_23060);
or U24048 (N_24048,N_23120,N_23896);
xor U24049 (N_24049,N_23299,N_23705);
xnor U24050 (N_24050,N_23777,N_23691);
or U24051 (N_24051,N_23936,N_23771);
and U24052 (N_24052,N_23540,N_23824);
xor U24053 (N_24053,N_23906,N_23345);
or U24054 (N_24054,N_23983,N_23359);
nand U24055 (N_24055,N_23348,N_23986);
or U24056 (N_24056,N_23703,N_23650);
nand U24057 (N_24057,N_23113,N_23701);
and U24058 (N_24058,N_23099,N_23803);
nor U24059 (N_24059,N_23231,N_23201);
and U24060 (N_24060,N_23239,N_23213);
xnor U24061 (N_24061,N_23932,N_23704);
and U24062 (N_24062,N_23808,N_23229);
xor U24063 (N_24063,N_23075,N_23496);
and U24064 (N_24064,N_23297,N_23475);
or U24065 (N_24065,N_23002,N_23172);
or U24066 (N_24066,N_23480,N_23747);
nand U24067 (N_24067,N_23186,N_23853);
or U24068 (N_24068,N_23991,N_23245);
nor U24069 (N_24069,N_23726,N_23437);
nand U24070 (N_24070,N_23317,N_23907);
nor U24071 (N_24071,N_23207,N_23005);
xnor U24072 (N_24072,N_23452,N_23690);
xnor U24073 (N_24073,N_23813,N_23310);
and U24074 (N_24074,N_23080,N_23056);
or U24075 (N_24075,N_23757,N_23730);
nor U24076 (N_24076,N_23057,N_23038);
xor U24077 (N_24077,N_23405,N_23817);
xnor U24078 (N_24078,N_23426,N_23341);
xor U24079 (N_24079,N_23271,N_23927);
and U24080 (N_24080,N_23911,N_23714);
xnor U24081 (N_24081,N_23468,N_23761);
and U24082 (N_24082,N_23654,N_23871);
and U24083 (N_24083,N_23121,N_23040);
or U24084 (N_24084,N_23920,N_23600);
nand U24085 (N_24085,N_23007,N_23801);
or U24086 (N_24086,N_23361,N_23846);
nor U24087 (N_24087,N_23611,N_23177);
xor U24088 (N_24088,N_23104,N_23135);
nand U24089 (N_24089,N_23622,N_23678);
or U24090 (N_24090,N_23039,N_23505);
nand U24091 (N_24091,N_23306,N_23513);
xnor U24092 (N_24092,N_23526,N_23598);
and U24093 (N_24093,N_23786,N_23095);
and U24094 (N_24094,N_23762,N_23301);
nand U24095 (N_24095,N_23545,N_23429);
and U24096 (N_24096,N_23127,N_23880);
or U24097 (N_24097,N_23291,N_23388);
nand U24098 (N_24098,N_23233,N_23787);
nand U24099 (N_24099,N_23877,N_23320);
or U24100 (N_24100,N_23634,N_23656);
nor U24101 (N_24101,N_23620,N_23217);
and U24102 (N_24102,N_23063,N_23413);
or U24103 (N_24103,N_23126,N_23879);
xor U24104 (N_24104,N_23574,N_23122);
nand U24105 (N_24105,N_23220,N_23888);
and U24106 (N_24106,N_23613,N_23281);
nor U24107 (N_24107,N_23794,N_23903);
and U24108 (N_24108,N_23129,N_23499);
nor U24109 (N_24109,N_23032,N_23358);
nor U24110 (N_24110,N_23603,N_23529);
or U24111 (N_24111,N_23328,N_23585);
nand U24112 (N_24112,N_23994,N_23826);
xor U24113 (N_24113,N_23098,N_23710);
or U24114 (N_24114,N_23103,N_23716);
or U24115 (N_24115,N_23664,N_23472);
nand U24116 (N_24116,N_23939,N_23658);
and U24117 (N_24117,N_23732,N_23205);
or U24118 (N_24118,N_23973,N_23527);
nand U24119 (N_24119,N_23117,N_23128);
or U24120 (N_24120,N_23887,N_23391);
and U24121 (N_24121,N_23322,N_23356);
xnor U24122 (N_24122,N_23064,N_23516);
nor U24123 (N_24123,N_23914,N_23783);
xnor U24124 (N_24124,N_23107,N_23442);
nor U24125 (N_24125,N_23416,N_23072);
nor U24126 (N_24126,N_23438,N_23267);
and U24127 (N_24127,N_23456,N_23941);
nand U24128 (N_24128,N_23640,N_23865);
nor U24129 (N_24129,N_23957,N_23555);
nand U24130 (N_24130,N_23195,N_23885);
and U24131 (N_24131,N_23676,N_23715);
nor U24132 (N_24132,N_23828,N_23194);
or U24133 (N_24133,N_23006,N_23258);
and U24134 (N_24134,N_23054,N_23548);
xor U24135 (N_24135,N_23897,N_23709);
nand U24136 (N_24136,N_23711,N_23048);
or U24137 (N_24137,N_23773,N_23367);
or U24138 (N_24138,N_23999,N_23717);
or U24139 (N_24139,N_23133,N_23176);
and U24140 (N_24140,N_23139,N_23062);
or U24141 (N_24141,N_23164,N_23190);
or U24142 (N_24142,N_23140,N_23158);
xor U24143 (N_24143,N_23840,N_23930);
nand U24144 (N_24144,N_23410,N_23241);
xor U24145 (N_24145,N_23825,N_23867);
or U24146 (N_24146,N_23562,N_23073);
and U24147 (N_24147,N_23542,N_23566);
or U24148 (N_24148,N_23541,N_23235);
nor U24149 (N_24149,N_23768,N_23249);
or U24150 (N_24150,N_23276,N_23616);
nor U24151 (N_24151,N_23988,N_23017);
nor U24152 (N_24152,N_23807,N_23350);
nor U24153 (N_24153,N_23153,N_23856);
xor U24154 (N_24154,N_23950,N_23336);
nor U24155 (N_24155,N_23234,N_23295);
nand U24156 (N_24156,N_23028,N_23615);
nand U24157 (N_24157,N_23363,N_23269);
and U24158 (N_24158,N_23157,N_23841);
xor U24159 (N_24159,N_23800,N_23035);
or U24160 (N_24160,N_23124,N_23296);
or U24161 (N_24161,N_23904,N_23298);
and U24162 (N_24162,N_23180,N_23254);
nor U24163 (N_24163,N_23156,N_23144);
nand U24164 (N_24164,N_23764,N_23908);
and U24165 (N_24165,N_23642,N_23384);
or U24166 (N_24166,N_23225,N_23076);
or U24167 (N_24167,N_23192,N_23462);
nor U24168 (N_24168,N_23791,N_23943);
or U24169 (N_24169,N_23004,N_23009);
nor U24170 (N_24170,N_23754,N_23440);
nand U24171 (N_24171,N_23047,N_23137);
or U24172 (N_24172,N_23671,N_23457);
and U24173 (N_24173,N_23211,N_23668);
or U24174 (N_24174,N_23025,N_23770);
nor U24175 (N_24175,N_23387,N_23382);
xnor U24176 (N_24176,N_23366,N_23816);
xnor U24177 (N_24177,N_23101,N_23769);
nor U24178 (N_24178,N_23995,N_23488);
xnor U24179 (N_24179,N_23189,N_23696);
or U24180 (N_24180,N_23952,N_23935);
and U24181 (N_24181,N_23493,N_23406);
nand U24182 (N_24182,N_23109,N_23015);
nand U24183 (N_24183,N_23170,N_23461);
nand U24184 (N_24184,N_23455,N_23230);
nor U24185 (N_24185,N_23978,N_23961);
and U24186 (N_24186,N_23740,N_23444);
xor U24187 (N_24187,N_23265,N_23778);
nand U24188 (N_24188,N_23221,N_23138);
or U24189 (N_24189,N_23244,N_23556);
nor U24190 (N_24190,N_23878,N_23683);
nor U24191 (N_24191,N_23814,N_23197);
or U24192 (N_24192,N_23392,N_23069);
xor U24193 (N_24193,N_23974,N_23130);
xor U24194 (N_24194,N_23481,N_23796);
nand U24195 (N_24195,N_23237,N_23250);
nor U24196 (N_24196,N_23931,N_23268);
or U24197 (N_24197,N_23872,N_23191);
or U24198 (N_24198,N_23082,N_23605);
nor U24199 (N_24199,N_23682,N_23357);
xnor U24200 (N_24200,N_23013,N_23171);
xnor U24201 (N_24201,N_23323,N_23873);
nor U24202 (N_24202,N_23661,N_23599);
and U24203 (N_24203,N_23147,N_23335);
or U24204 (N_24204,N_23026,N_23987);
nor U24205 (N_24205,N_23094,N_23398);
nand U24206 (N_24206,N_23832,N_23123);
or U24207 (N_24207,N_23626,N_23108);
or U24208 (N_24208,N_23402,N_23728);
or U24209 (N_24209,N_23396,N_23624);
or U24210 (N_24210,N_23942,N_23305);
or U24211 (N_24211,N_23092,N_23970);
nand U24212 (N_24212,N_23251,N_23347);
xor U24213 (N_24213,N_23324,N_23012);
and U24214 (N_24214,N_23590,N_23627);
nand U24215 (N_24215,N_23788,N_23912);
xnor U24216 (N_24216,N_23053,N_23264);
nor U24217 (N_24217,N_23018,N_23355);
nand U24218 (N_24218,N_23262,N_23115);
or U24219 (N_24219,N_23173,N_23100);
nand U24220 (N_24220,N_23168,N_23765);
and U24221 (N_24221,N_23719,N_23415);
or U24222 (N_24222,N_23061,N_23698);
nand U24223 (N_24223,N_23504,N_23509);
or U24224 (N_24224,N_23604,N_23154);
nor U24225 (N_24225,N_23522,N_23460);
nand U24226 (N_24226,N_23334,N_23797);
or U24227 (N_24227,N_23326,N_23011);
or U24228 (N_24228,N_23558,N_23159);
nand U24229 (N_24229,N_23809,N_23758);
and U24230 (N_24230,N_23539,N_23739);
and U24231 (N_24231,N_23655,N_23597);
xor U24232 (N_24232,N_23951,N_23422);
and U24233 (N_24233,N_23175,N_23077);
nand U24234 (N_24234,N_23637,N_23318);
xor U24235 (N_24235,N_23967,N_23923);
nand U24236 (N_24236,N_23469,N_23776);
or U24237 (N_24237,N_23781,N_23439);
and U24238 (N_24238,N_23763,N_23198);
and U24239 (N_24239,N_23313,N_23282);
nand U24240 (N_24240,N_23304,N_23523);
nor U24241 (N_24241,N_23514,N_23148);
nand U24242 (N_24242,N_23855,N_23915);
or U24243 (N_24243,N_23352,N_23247);
nand U24244 (N_24244,N_23666,N_23780);
nand U24245 (N_24245,N_23836,N_23424);
and U24246 (N_24246,N_23652,N_23169);
nand U24247 (N_24247,N_23353,N_23097);
xnor U24248 (N_24248,N_23659,N_23495);
nor U24249 (N_24249,N_23632,N_23346);
xor U24250 (N_24250,N_23476,N_23820);
xor U24251 (N_24251,N_23532,N_23881);
and U24252 (N_24252,N_23465,N_23360);
nand U24253 (N_24253,N_23374,N_23584);
nand U24254 (N_24254,N_23969,N_23806);
nor U24255 (N_24255,N_23498,N_23021);
nand U24256 (N_24256,N_23606,N_23838);
nand U24257 (N_24257,N_23188,N_23378);
xor U24258 (N_24258,N_23071,N_23477);
nand U24259 (N_24259,N_23022,N_23567);
nand U24260 (N_24260,N_23815,N_23284);
xor U24261 (N_24261,N_23362,N_23102);
xor U24262 (N_24262,N_23381,N_23687);
and U24263 (N_24263,N_23512,N_23901);
or U24264 (N_24264,N_23232,N_23735);
xnor U24265 (N_24265,N_23766,N_23583);
xnor U24266 (N_24266,N_23894,N_23672);
xor U24267 (N_24267,N_23216,N_23638);
nor U24268 (N_24268,N_23775,N_23008);
nand U24269 (N_24269,N_23618,N_23280);
nand U24270 (N_24270,N_23131,N_23753);
xor U24271 (N_24271,N_23473,N_23275);
and U24272 (N_24272,N_23261,N_23517);
and U24273 (N_24273,N_23633,N_23091);
nand U24274 (N_24274,N_23308,N_23450);
nand U24275 (N_24275,N_23243,N_23023);
nand U24276 (N_24276,N_23926,N_23863);
or U24277 (N_24277,N_23707,N_23660);
or U24278 (N_24278,N_23534,N_23070);
xnor U24279 (N_24279,N_23149,N_23434);
and U24280 (N_24280,N_23435,N_23528);
or U24281 (N_24281,N_23641,N_23720);
nand U24282 (N_24282,N_23551,N_23500);
xor U24283 (N_24283,N_23743,N_23893);
xnor U24284 (N_24284,N_23218,N_23582);
nand U24285 (N_24285,N_23966,N_23373);
nor U24286 (N_24286,N_23960,N_23253);
xnor U24287 (N_24287,N_23431,N_23287);
and U24288 (N_24288,N_23850,N_23212);
nor U24289 (N_24289,N_23546,N_23050);
nor U24290 (N_24290,N_23270,N_23215);
and U24291 (N_24291,N_23371,N_23602);
and U24292 (N_24292,N_23617,N_23016);
and U24293 (N_24293,N_23533,N_23937);
and U24294 (N_24294,N_23827,N_23343);
or U24295 (N_24295,N_23575,N_23272);
nor U24296 (N_24296,N_23674,N_23182);
nand U24297 (N_24297,N_23226,N_23459);
nand U24298 (N_24298,N_23518,N_23610);
nor U24299 (N_24299,N_23859,N_23277);
xor U24300 (N_24300,N_23079,N_23266);
or U24301 (N_24301,N_23403,N_23756);
xnor U24302 (N_24302,N_23552,N_23689);
or U24303 (N_24303,N_23507,N_23849);
xor U24304 (N_24304,N_23464,N_23206);
xor U24305 (N_24305,N_23535,N_23725);
or U24306 (N_24306,N_23630,N_23364);
xor U24307 (N_24307,N_23662,N_23125);
and U24308 (N_24308,N_23785,N_23290);
xor U24309 (N_24309,N_23412,N_23578);
xor U24310 (N_24310,N_23116,N_23145);
xor U24311 (N_24311,N_23315,N_23921);
and U24312 (N_24312,N_23046,N_23185);
xor U24313 (N_24313,N_23549,N_23034);
or U24314 (N_24314,N_23645,N_23058);
nand U24315 (N_24315,N_23947,N_23390);
nand U24316 (N_24316,N_23579,N_23204);
or U24317 (N_24317,N_23407,N_23723);
and U24318 (N_24318,N_23030,N_23996);
xnor U24319 (N_24319,N_23644,N_23411);
xnor U24320 (N_24320,N_23478,N_23494);
and U24321 (N_24321,N_23319,N_23490);
and U24322 (N_24322,N_23033,N_23955);
nor U24323 (N_24323,N_23621,N_23848);
nor U24324 (N_24324,N_23303,N_23394);
nor U24325 (N_24325,N_23933,N_23560);
xor U24326 (N_24326,N_23327,N_23344);
and U24327 (N_24327,N_23889,N_23760);
nand U24328 (N_24328,N_23420,N_23379);
nand U24329 (N_24329,N_23647,N_23913);
nand U24330 (N_24330,N_23238,N_23027);
nor U24331 (N_24331,N_23677,N_23759);
nand U24332 (N_24332,N_23041,N_23184);
nand U24333 (N_24333,N_23792,N_23953);
nand U24334 (N_24334,N_23257,N_23708);
nor U24335 (N_24335,N_23553,N_23981);
xnor U24336 (N_24336,N_23819,N_23537);
or U24337 (N_24337,N_23854,N_23372);
nand U24338 (N_24338,N_23467,N_23368);
or U24339 (N_24339,N_23721,N_23179);
and U24340 (N_24340,N_23802,N_23530);
or U24341 (N_24341,N_23805,N_23110);
nand U24342 (N_24342,N_23279,N_23589);
xnor U24343 (N_24343,N_23886,N_23083);
nand U24344 (N_24344,N_23569,N_23712);
nor U24345 (N_24345,N_23612,N_23608);
or U24346 (N_24346,N_23857,N_23090);
nand U24347 (N_24347,N_23491,N_23874);
nand U24348 (N_24348,N_23492,N_23744);
nor U24349 (N_24349,N_23330,N_23695);
or U24350 (N_24350,N_23985,N_23918);
nand U24351 (N_24351,N_23400,N_23001);
and U24352 (N_24352,N_23968,N_23614);
xor U24353 (N_24353,N_23163,N_23065);
xnor U24354 (N_24354,N_23134,N_23669);
or U24355 (N_24355,N_23414,N_23224);
nand U24356 (N_24356,N_23375,N_23587);
xor U24357 (N_24357,N_23547,N_23568);
xnor U24358 (N_24358,N_23884,N_23000);
xnor U24359 (N_24359,N_23052,N_23486);
and U24360 (N_24360,N_23833,N_23055);
nand U24361 (N_24361,N_23161,N_23515);
or U24362 (N_24362,N_23259,N_23868);
and U24363 (N_24363,N_23449,N_23288);
nand U24364 (N_24364,N_23564,N_23971);
or U24365 (N_24365,N_23165,N_23453);
or U24366 (N_24366,N_23559,N_23869);
nand U24367 (N_24367,N_23593,N_23214);
xnor U24368 (N_24368,N_23900,N_23899);
nand U24369 (N_24369,N_23369,N_23588);
and U24370 (N_24370,N_23818,N_23155);
xnor U24371 (N_24371,N_23501,N_23273);
nand U24372 (N_24372,N_23997,N_23713);
and U24373 (N_24373,N_23289,N_23636);
nand U24374 (N_24374,N_23089,N_23675);
and U24375 (N_24375,N_23255,N_23702);
xor U24376 (N_24376,N_23625,N_23917);
xor U24377 (N_24377,N_23685,N_23860);
xor U24378 (N_24378,N_23433,N_23037);
and U24379 (N_24379,N_23525,N_23699);
xnor U24380 (N_24380,N_23977,N_23031);
xor U24381 (N_24381,N_23436,N_23830);
nand U24382 (N_24382,N_23684,N_23876);
nand U24383 (N_24383,N_23581,N_23954);
xor U24384 (N_24384,N_23294,N_23260);
or U24385 (N_24385,N_23293,N_23831);
and U24386 (N_24386,N_23844,N_23653);
nand U24387 (N_24387,N_23870,N_23086);
nand U24388 (N_24388,N_23576,N_23834);
or U24389 (N_24389,N_23822,N_23752);
and U24390 (N_24390,N_23990,N_23601);
or U24391 (N_24391,N_23670,N_23916);
or U24392 (N_24392,N_23141,N_23078);
nand U24393 (N_24393,N_23922,N_23285);
and U24394 (N_24394,N_23619,N_23487);
or U24395 (N_24395,N_23934,N_23042);
nand U24396 (N_24396,N_23851,N_23949);
and U24397 (N_24397,N_23919,N_23680);
and U24398 (N_24398,N_23554,N_23858);
xor U24399 (N_24399,N_23767,N_23114);
nand U24400 (N_24400,N_23875,N_23506);
nand U24401 (N_24401,N_23146,N_23793);
and U24402 (N_24402,N_23998,N_23804);
nand U24403 (N_24403,N_23187,N_23561);
and U24404 (N_24404,N_23150,N_23423);
nor U24405 (N_24405,N_23314,N_23852);
nor U24406 (N_24406,N_23902,N_23393);
and U24407 (N_24407,N_23651,N_23325);
xnor U24408 (N_24408,N_23430,N_23408);
or U24409 (N_24409,N_23928,N_23938);
nor U24410 (N_24410,N_23043,N_23779);
and U24411 (N_24411,N_23521,N_23445);
or U24412 (N_24412,N_23193,N_23479);
xnor U24413 (N_24413,N_23948,N_23377);
and U24414 (N_24414,N_23891,N_23029);
nand U24415 (N_24415,N_23543,N_23044);
nor U24416 (N_24416,N_23136,N_23466);
xor U24417 (N_24417,N_23639,N_23209);
and U24418 (N_24418,N_23331,N_23631);
nor U24419 (N_24419,N_23338,N_23727);
or U24420 (N_24420,N_23510,N_23741);
or U24421 (N_24421,N_23697,N_23160);
nand U24422 (N_24422,N_23242,N_23706);
and U24423 (N_24423,N_23105,N_23085);
and U24424 (N_24424,N_23081,N_23965);
nand U24425 (N_24425,N_23538,N_23837);
and U24426 (N_24426,N_23300,N_23471);
nand U24427 (N_24427,N_23643,N_23096);
nor U24428 (N_24428,N_23112,N_23196);
xor U24429 (N_24429,N_23746,N_23993);
xnor U24430 (N_24430,N_23508,N_23734);
nand U24431 (N_24431,N_23470,N_23223);
xnor U24432 (N_24432,N_23419,N_23370);
or U24433 (N_24433,N_23751,N_23199);
or U24434 (N_24434,N_23586,N_23203);
xor U24435 (N_24435,N_23686,N_23311);
xnor U24436 (N_24436,N_23745,N_23945);
or U24437 (N_24437,N_23045,N_23845);
or U24438 (N_24438,N_23511,N_23749);
or U24439 (N_24439,N_23989,N_23389);
and U24440 (N_24440,N_23166,N_23811);
and U24441 (N_24441,N_23399,N_23307);
or U24442 (N_24442,N_23657,N_23864);
nand U24443 (N_24443,N_23898,N_23427);
nand U24444 (N_24444,N_23940,N_23302);
or U24445 (N_24445,N_23417,N_23283);
or U24446 (N_24446,N_23629,N_23924);
and U24447 (N_24447,N_23386,N_23842);
xnor U24448 (N_24448,N_23349,N_23774);
and U24449 (N_24449,N_23524,N_23862);
nand U24450 (N_24450,N_23278,N_23151);
or U24451 (N_24451,N_23019,N_23228);
or U24452 (N_24452,N_23649,N_23014);
or U24453 (N_24453,N_23167,N_23074);
nor U24454 (N_24454,N_23648,N_23992);
xnor U24455 (N_24455,N_23984,N_23210);
and U24456 (N_24456,N_23635,N_23132);
or U24457 (N_24457,N_23572,N_23397);
or U24458 (N_24458,N_23446,N_23256);
nor U24459 (N_24459,N_23592,N_23425);
xor U24460 (N_24460,N_23733,N_23401);
nand U24461 (N_24461,N_23946,N_23380);
xor U24462 (N_24462,N_23332,N_23106);
nor U24463 (N_24463,N_23329,N_23795);
nand U24464 (N_24464,N_23963,N_23810);
nor U24465 (N_24465,N_23519,N_23351);
nand U24466 (N_24466,N_23565,N_23292);
nand U24467 (N_24467,N_23839,N_23910);
or U24468 (N_24468,N_23890,N_23531);
and U24469 (N_24469,N_23679,N_23395);
xor U24470 (N_24470,N_23628,N_23010);
xnor U24471 (N_24471,N_23979,N_23557);
or U24472 (N_24472,N_23404,N_23383);
nor U24473 (N_24473,N_23835,N_23321);
or U24474 (N_24474,N_23905,N_23183);
or U24475 (N_24475,N_23339,N_23976);
or U24476 (N_24476,N_23503,N_23681);
nor U24477 (N_24477,N_23051,N_23609);
nand U24478 (N_24478,N_23544,N_23312);
nor U24479 (N_24479,N_23673,N_23790);
nor U24480 (N_24480,N_23975,N_23119);
nor U24481 (N_24481,N_23736,N_23162);
and U24482 (N_24482,N_23722,N_23929);
nor U24483 (N_24483,N_23595,N_23143);
or U24484 (N_24484,N_23812,N_23208);
nand U24485 (N_24485,N_23577,N_23376);
and U24486 (N_24486,N_23174,N_23337);
xor U24487 (N_24487,N_23316,N_23443);
nand U24488 (N_24488,N_23236,N_23520);
nor U24489 (N_24489,N_23866,N_23750);
and U24490 (N_24490,N_23847,N_23724);
nor U24491 (N_24491,N_23550,N_23799);
xnor U24492 (N_24492,N_23972,N_23200);
nand U24493 (N_24493,N_23729,N_23909);
nand U24494 (N_24494,N_23049,N_23959);
nor U24495 (N_24495,N_23665,N_23571);
or U24496 (N_24496,N_23789,N_23646);
nor U24497 (N_24497,N_23748,N_23447);
nor U24498 (N_24498,N_23340,N_23663);
or U24499 (N_24499,N_23451,N_23428);
xor U24500 (N_24500,N_23464,N_23921);
nand U24501 (N_24501,N_23511,N_23254);
xor U24502 (N_24502,N_23977,N_23273);
xor U24503 (N_24503,N_23442,N_23155);
nor U24504 (N_24504,N_23028,N_23692);
or U24505 (N_24505,N_23409,N_23782);
and U24506 (N_24506,N_23040,N_23656);
or U24507 (N_24507,N_23803,N_23107);
and U24508 (N_24508,N_23269,N_23628);
xor U24509 (N_24509,N_23373,N_23217);
nor U24510 (N_24510,N_23119,N_23252);
nor U24511 (N_24511,N_23844,N_23961);
nand U24512 (N_24512,N_23853,N_23088);
or U24513 (N_24513,N_23969,N_23417);
nand U24514 (N_24514,N_23311,N_23419);
or U24515 (N_24515,N_23921,N_23051);
xor U24516 (N_24516,N_23757,N_23271);
nor U24517 (N_24517,N_23106,N_23680);
nor U24518 (N_24518,N_23993,N_23504);
or U24519 (N_24519,N_23885,N_23661);
and U24520 (N_24520,N_23018,N_23131);
xor U24521 (N_24521,N_23043,N_23130);
and U24522 (N_24522,N_23589,N_23018);
or U24523 (N_24523,N_23917,N_23614);
nor U24524 (N_24524,N_23635,N_23528);
and U24525 (N_24525,N_23988,N_23744);
xnor U24526 (N_24526,N_23949,N_23184);
xnor U24527 (N_24527,N_23466,N_23603);
or U24528 (N_24528,N_23654,N_23299);
xor U24529 (N_24529,N_23788,N_23680);
or U24530 (N_24530,N_23045,N_23572);
nand U24531 (N_24531,N_23633,N_23270);
nand U24532 (N_24532,N_23283,N_23522);
or U24533 (N_24533,N_23867,N_23977);
and U24534 (N_24534,N_23133,N_23138);
and U24535 (N_24535,N_23640,N_23641);
nor U24536 (N_24536,N_23630,N_23269);
or U24537 (N_24537,N_23092,N_23430);
and U24538 (N_24538,N_23508,N_23986);
nor U24539 (N_24539,N_23309,N_23520);
and U24540 (N_24540,N_23339,N_23669);
xnor U24541 (N_24541,N_23682,N_23642);
or U24542 (N_24542,N_23659,N_23110);
xnor U24543 (N_24543,N_23813,N_23884);
and U24544 (N_24544,N_23281,N_23584);
xor U24545 (N_24545,N_23122,N_23845);
xor U24546 (N_24546,N_23938,N_23976);
or U24547 (N_24547,N_23186,N_23740);
or U24548 (N_24548,N_23189,N_23018);
and U24549 (N_24549,N_23066,N_23971);
or U24550 (N_24550,N_23754,N_23971);
and U24551 (N_24551,N_23396,N_23135);
nand U24552 (N_24552,N_23918,N_23302);
xor U24553 (N_24553,N_23196,N_23381);
and U24554 (N_24554,N_23132,N_23555);
nor U24555 (N_24555,N_23274,N_23095);
and U24556 (N_24556,N_23023,N_23796);
nor U24557 (N_24557,N_23280,N_23760);
or U24558 (N_24558,N_23737,N_23796);
and U24559 (N_24559,N_23992,N_23447);
nand U24560 (N_24560,N_23530,N_23210);
nor U24561 (N_24561,N_23582,N_23158);
or U24562 (N_24562,N_23183,N_23935);
or U24563 (N_24563,N_23693,N_23860);
and U24564 (N_24564,N_23461,N_23248);
and U24565 (N_24565,N_23615,N_23284);
and U24566 (N_24566,N_23421,N_23044);
and U24567 (N_24567,N_23642,N_23167);
nor U24568 (N_24568,N_23740,N_23917);
and U24569 (N_24569,N_23402,N_23417);
nand U24570 (N_24570,N_23646,N_23233);
or U24571 (N_24571,N_23612,N_23390);
and U24572 (N_24572,N_23225,N_23958);
xor U24573 (N_24573,N_23976,N_23317);
nand U24574 (N_24574,N_23029,N_23613);
or U24575 (N_24575,N_23321,N_23052);
nand U24576 (N_24576,N_23824,N_23208);
and U24577 (N_24577,N_23410,N_23357);
xor U24578 (N_24578,N_23679,N_23050);
nor U24579 (N_24579,N_23706,N_23842);
nor U24580 (N_24580,N_23916,N_23157);
nand U24581 (N_24581,N_23569,N_23404);
nor U24582 (N_24582,N_23374,N_23642);
or U24583 (N_24583,N_23102,N_23415);
xnor U24584 (N_24584,N_23072,N_23130);
nor U24585 (N_24585,N_23161,N_23417);
nand U24586 (N_24586,N_23683,N_23434);
and U24587 (N_24587,N_23382,N_23625);
and U24588 (N_24588,N_23296,N_23705);
nor U24589 (N_24589,N_23599,N_23842);
nand U24590 (N_24590,N_23191,N_23422);
xnor U24591 (N_24591,N_23343,N_23971);
or U24592 (N_24592,N_23401,N_23867);
or U24593 (N_24593,N_23434,N_23590);
xor U24594 (N_24594,N_23413,N_23695);
nand U24595 (N_24595,N_23917,N_23084);
xor U24596 (N_24596,N_23072,N_23791);
xor U24597 (N_24597,N_23973,N_23122);
nor U24598 (N_24598,N_23875,N_23002);
and U24599 (N_24599,N_23041,N_23364);
nor U24600 (N_24600,N_23098,N_23354);
nand U24601 (N_24601,N_23903,N_23302);
or U24602 (N_24602,N_23466,N_23193);
xor U24603 (N_24603,N_23154,N_23563);
or U24604 (N_24604,N_23114,N_23103);
nand U24605 (N_24605,N_23510,N_23520);
and U24606 (N_24606,N_23750,N_23577);
and U24607 (N_24607,N_23725,N_23448);
nand U24608 (N_24608,N_23529,N_23122);
nor U24609 (N_24609,N_23360,N_23055);
or U24610 (N_24610,N_23143,N_23400);
nor U24611 (N_24611,N_23781,N_23098);
xor U24612 (N_24612,N_23080,N_23027);
nor U24613 (N_24613,N_23639,N_23051);
and U24614 (N_24614,N_23622,N_23398);
nand U24615 (N_24615,N_23313,N_23770);
nand U24616 (N_24616,N_23551,N_23187);
or U24617 (N_24617,N_23135,N_23497);
nor U24618 (N_24618,N_23385,N_23214);
nor U24619 (N_24619,N_23759,N_23891);
nand U24620 (N_24620,N_23081,N_23326);
xor U24621 (N_24621,N_23425,N_23871);
and U24622 (N_24622,N_23393,N_23033);
nor U24623 (N_24623,N_23845,N_23320);
xor U24624 (N_24624,N_23735,N_23952);
or U24625 (N_24625,N_23035,N_23359);
and U24626 (N_24626,N_23966,N_23605);
and U24627 (N_24627,N_23518,N_23541);
and U24628 (N_24628,N_23337,N_23419);
nor U24629 (N_24629,N_23554,N_23101);
nand U24630 (N_24630,N_23993,N_23950);
xnor U24631 (N_24631,N_23008,N_23646);
xnor U24632 (N_24632,N_23213,N_23877);
nand U24633 (N_24633,N_23538,N_23500);
xor U24634 (N_24634,N_23615,N_23191);
nor U24635 (N_24635,N_23640,N_23169);
nor U24636 (N_24636,N_23394,N_23065);
nand U24637 (N_24637,N_23692,N_23215);
nor U24638 (N_24638,N_23718,N_23594);
xor U24639 (N_24639,N_23934,N_23560);
or U24640 (N_24640,N_23508,N_23587);
xor U24641 (N_24641,N_23140,N_23922);
or U24642 (N_24642,N_23457,N_23092);
and U24643 (N_24643,N_23411,N_23337);
nand U24644 (N_24644,N_23092,N_23223);
xor U24645 (N_24645,N_23008,N_23840);
xor U24646 (N_24646,N_23139,N_23937);
nand U24647 (N_24647,N_23926,N_23462);
nand U24648 (N_24648,N_23972,N_23270);
and U24649 (N_24649,N_23387,N_23001);
nand U24650 (N_24650,N_23355,N_23918);
or U24651 (N_24651,N_23780,N_23528);
or U24652 (N_24652,N_23262,N_23592);
and U24653 (N_24653,N_23891,N_23066);
nor U24654 (N_24654,N_23822,N_23609);
nor U24655 (N_24655,N_23248,N_23660);
xnor U24656 (N_24656,N_23519,N_23317);
and U24657 (N_24657,N_23282,N_23895);
or U24658 (N_24658,N_23645,N_23208);
and U24659 (N_24659,N_23341,N_23706);
nand U24660 (N_24660,N_23144,N_23605);
or U24661 (N_24661,N_23696,N_23060);
xnor U24662 (N_24662,N_23378,N_23511);
or U24663 (N_24663,N_23735,N_23927);
and U24664 (N_24664,N_23540,N_23033);
and U24665 (N_24665,N_23031,N_23396);
and U24666 (N_24666,N_23405,N_23280);
xnor U24667 (N_24667,N_23139,N_23512);
and U24668 (N_24668,N_23975,N_23086);
nor U24669 (N_24669,N_23363,N_23729);
or U24670 (N_24670,N_23121,N_23506);
nand U24671 (N_24671,N_23113,N_23633);
nand U24672 (N_24672,N_23597,N_23018);
nand U24673 (N_24673,N_23871,N_23452);
nor U24674 (N_24674,N_23372,N_23691);
and U24675 (N_24675,N_23581,N_23338);
or U24676 (N_24676,N_23478,N_23628);
nor U24677 (N_24677,N_23453,N_23475);
nand U24678 (N_24678,N_23661,N_23893);
or U24679 (N_24679,N_23149,N_23239);
and U24680 (N_24680,N_23706,N_23620);
or U24681 (N_24681,N_23242,N_23726);
and U24682 (N_24682,N_23491,N_23864);
or U24683 (N_24683,N_23800,N_23339);
nor U24684 (N_24684,N_23824,N_23065);
xnor U24685 (N_24685,N_23585,N_23293);
or U24686 (N_24686,N_23491,N_23743);
nand U24687 (N_24687,N_23356,N_23900);
or U24688 (N_24688,N_23715,N_23342);
and U24689 (N_24689,N_23275,N_23875);
or U24690 (N_24690,N_23422,N_23622);
and U24691 (N_24691,N_23206,N_23893);
or U24692 (N_24692,N_23953,N_23172);
nand U24693 (N_24693,N_23793,N_23483);
nor U24694 (N_24694,N_23987,N_23057);
and U24695 (N_24695,N_23132,N_23881);
nand U24696 (N_24696,N_23578,N_23236);
or U24697 (N_24697,N_23587,N_23226);
xnor U24698 (N_24698,N_23056,N_23564);
nor U24699 (N_24699,N_23640,N_23729);
xor U24700 (N_24700,N_23481,N_23077);
or U24701 (N_24701,N_23919,N_23447);
xor U24702 (N_24702,N_23416,N_23574);
and U24703 (N_24703,N_23461,N_23300);
and U24704 (N_24704,N_23696,N_23014);
and U24705 (N_24705,N_23824,N_23546);
or U24706 (N_24706,N_23728,N_23562);
nand U24707 (N_24707,N_23884,N_23867);
nor U24708 (N_24708,N_23176,N_23924);
or U24709 (N_24709,N_23279,N_23684);
nor U24710 (N_24710,N_23089,N_23195);
nand U24711 (N_24711,N_23922,N_23933);
nand U24712 (N_24712,N_23127,N_23684);
nand U24713 (N_24713,N_23576,N_23302);
or U24714 (N_24714,N_23884,N_23588);
xor U24715 (N_24715,N_23231,N_23961);
nand U24716 (N_24716,N_23397,N_23498);
and U24717 (N_24717,N_23498,N_23719);
nand U24718 (N_24718,N_23942,N_23719);
and U24719 (N_24719,N_23579,N_23519);
or U24720 (N_24720,N_23428,N_23802);
or U24721 (N_24721,N_23254,N_23734);
xor U24722 (N_24722,N_23647,N_23673);
or U24723 (N_24723,N_23640,N_23069);
nor U24724 (N_24724,N_23857,N_23019);
xor U24725 (N_24725,N_23605,N_23408);
nor U24726 (N_24726,N_23199,N_23476);
xor U24727 (N_24727,N_23610,N_23113);
nor U24728 (N_24728,N_23840,N_23430);
or U24729 (N_24729,N_23276,N_23740);
xor U24730 (N_24730,N_23384,N_23420);
and U24731 (N_24731,N_23836,N_23447);
nand U24732 (N_24732,N_23805,N_23722);
or U24733 (N_24733,N_23097,N_23051);
nand U24734 (N_24734,N_23883,N_23677);
and U24735 (N_24735,N_23096,N_23844);
nand U24736 (N_24736,N_23507,N_23093);
nand U24737 (N_24737,N_23295,N_23237);
or U24738 (N_24738,N_23263,N_23831);
or U24739 (N_24739,N_23909,N_23662);
nand U24740 (N_24740,N_23744,N_23443);
xor U24741 (N_24741,N_23016,N_23262);
nor U24742 (N_24742,N_23431,N_23854);
and U24743 (N_24743,N_23764,N_23771);
nor U24744 (N_24744,N_23693,N_23859);
nand U24745 (N_24745,N_23751,N_23329);
nor U24746 (N_24746,N_23448,N_23632);
xnor U24747 (N_24747,N_23326,N_23541);
nand U24748 (N_24748,N_23296,N_23743);
nand U24749 (N_24749,N_23585,N_23458);
nor U24750 (N_24750,N_23820,N_23328);
and U24751 (N_24751,N_23482,N_23445);
nand U24752 (N_24752,N_23747,N_23119);
nor U24753 (N_24753,N_23636,N_23129);
xnor U24754 (N_24754,N_23438,N_23182);
or U24755 (N_24755,N_23540,N_23037);
and U24756 (N_24756,N_23019,N_23551);
nand U24757 (N_24757,N_23446,N_23371);
and U24758 (N_24758,N_23319,N_23148);
nand U24759 (N_24759,N_23125,N_23437);
and U24760 (N_24760,N_23662,N_23693);
nor U24761 (N_24761,N_23776,N_23681);
nor U24762 (N_24762,N_23526,N_23548);
or U24763 (N_24763,N_23190,N_23388);
and U24764 (N_24764,N_23689,N_23103);
nand U24765 (N_24765,N_23768,N_23742);
and U24766 (N_24766,N_23920,N_23924);
xnor U24767 (N_24767,N_23928,N_23561);
or U24768 (N_24768,N_23927,N_23864);
xnor U24769 (N_24769,N_23164,N_23576);
and U24770 (N_24770,N_23130,N_23938);
nand U24771 (N_24771,N_23703,N_23792);
nor U24772 (N_24772,N_23586,N_23666);
xor U24773 (N_24773,N_23323,N_23872);
nor U24774 (N_24774,N_23243,N_23656);
and U24775 (N_24775,N_23273,N_23165);
nand U24776 (N_24776,N_23835,N_23109);
nand U24777 (N_24777,N_23989,N_23496);
or U24778 (N_24778,N_23481,N_23633);
nor U24779 (N_24779,N_23078,N_23184);
or U24780 (N_24780,N_23181,N_23625);
or U24781 (N_24781,N_23844,N_23983);
xor U24782 (N_24782,N_23157,N_23184);
nand U24783 (N_24783,N_23804,N_23410);
or U24784 (N_24784,N_23657,N_23786);
or U24785 (N_24785,N_23509,N_23392);
nand U24786 (N_24786,N_23933,N_23832);
nor U24787 (N_24787,N_23916,N_23080);
or U24788 (N_24788,N_23127,N_23787);
and U24789 (N_24789,N_23365,N_23214);
and U24790 (N_24790,N_23680,N_23408);
nor U24791 (N_24791,N_23415,N_23762);
nor U24792 (N_24792,N_23367,N_23208);
nand U24793 (N_24793,N_23415,N_23909);
and U24794 (N_24794,N_23023,N_23196);
and U24795 (N_24795,N_23781,N_23932);
or U24796 (N_24796,N_23359,N_23570);
or U24797 (N_24797,N_23485,N_23566);
nor U24798 (N_24798,N_23146,N_23499);
and U24799 (N_24799,N_23887,N_23009);
and U24800 (N_24800,N_23650,N_23208);
or U24801 (N_24801,N_23146,N_23101);
xor U24802 (N_24802,N_23594,N_23901);
and U24803 (N_24803,N_23372,N_23937);
nor U24804 (N_24804,N_23884,N_23497);
and U24805 (N_24805,N_23294,N_23853);
or U24806 (N_24806,N_23017,N_23531);
or U24807 (N_24807,N_23824,N_23552);
nor U24808 (N_24808,N_23906,N_23782);
and U24809 (N_24809,N_23608,N_23772);
or U24810 (N_24810,N_23635,N_23021);
xnor U24811 (N_24811,N_23575,N_23654);
xor U24812 (N_24812,N_23220,N_23369);
or U24813 (N_24813,N_23624,N_23114);
nor U24814 (N_24814,N_23636,N_23488);
xnor U24815 (N_24815,N_23710,N_23658);
nand U24816 (N_24816,N_23951,N_23425);
nand U24817 (N_24817,N_23591,N_23239);
nand U24818 (N_24818,N_23874,N_23617);
nand U24819 (N_24819,N_23534,N_23844);
nor U24820 (N_24820,N_23046,N_23405);
nor U24821 (N_24821,N_23571,N_23535);
and U24822 (N_24822,N_23824,N_23245);
nand U24823 (N_24823,N_23954,N_23147);
xor U24824 (N_24824,N_23667,N_23807);
nor U24825 (N_24825,N_23211,N_23428);
and U24826 (N_24826,N_23156,N_23570);
xnor U24827 (N_24827,N_23613,N_23466);
nor U24828 (N_24828,N_23162,N_23757);
and U24829 (N_24829,N_23722,N_23667);
or U24830 (N_24830,N_23667,N_23922);
xnor U24831 (N_24831,N_23998,N_23815);
nor U24832 (N_24832,N_23664,N_23207);
and U24833 (N_24833,N_23461,N_23692);
nor U24834 (N_24834,N_23186,N_23240);
xnor U24835 (N_24835,N_23539,N_23048);
xor U24836 (N_24836,N_23098,N_23603);
or U24837 (N_24837,N_23934,N_23073);
or U24838 (N_24838,N_23505,N_23234);
or U24839 (N_24839,N_23538,N_23772);
or U24840 (N_24840,N_23467,N_23385);
nand U24841 (N_24841,N_23698,N_23761);
nand U24842 (N_24842,N_23701,N_23637);
nor U24843 (N_24843,N_23573,N_23375);
or U24844 (N_24844,N_23336,N_23309);
nand U24845 (N_24845,N_23832,N_23507);
or U24846 (N_24846,N_23341,N_23473);
or U24847 (N_24847,N_23945,N_23139);
nand U24848 (N_24848,N_23556,N_23780);
xnor U24849 (N_24849,N_23339,N_23602);
nor U24850 (N_24850,N_23063,N_23616);
nor U24851 (N_24851,N_23025,N_23620);
and U24852 (N_24852,N_23103,N_23854);
xnor U24853 (N_24853,N_23316,N_23436);
xor U24854 (N_24854,N_23973,N_23427);
nor U24855 (N_24855,N_23975,N_23008);
or U24856 (N_24856,N_23202,N_23839);
or U24857 (N_24857,N_23771,N_23667);
nor U24858 (N_24858,N_23943,N_23079);
xor U24859 (N_24859,N_23707,N_23454);
or U24860 (N_24860,N_23575,N_23404);
or U24861 (N_24861,N_23483,N_23760);
or U24862 (N_24862,N_23644,N_23720);
nor U24863 (N_24863,N_23132,N_23685);
xnor U24864 (N_24864,N_23366,N_23149);
nand U24865 (N_24865,N_23678,N_23639);
and U24866 (N_24866,N_23372,N_23293);
nor U24867 (N_24867,N_23044,N_23426);
or U24868 (N_24868,N_23477,N_23861);
nor U24869 (N_24869,N_23810,N_23895);
xor U24870 (N_24870,N_23008,N_23125);
nor U24871 (N_24871,N_23771,N_23479);
nand U24872 (N_24872,N_23669,N_23612);
xnor U24873 (N_24873,N_23188,N_23859);
or U24874 (N_24874,N_23272,N_23140);
xor U24875 (N_24875,N_23586,N_23164);
nand U24876 (N_24876,N_23680,N_23155);
xor U24877 (N_24877,N_23392,N_23942);
and U24878 (N_24878,N_23571,N_23711);
xnor U24879 (N_24879,N_23262,N_23401);
nand U24880 (N_24880,N_23710,N_23791);
nor U24881 (N_24881,N_23465,N_23100);
nor U24882 (N_24882,N_23582,N_23760);
nor U24883 (N_24883,N_23805,N_23358);
nor U24884 (N_24884,N_23509,N_23121);
or U24885 (N_24885,N_23847,N_23285);
or U24886 (N_24886,N_23200,N_23501);
or U24887 (N_24887,N_23846,N_23859);
or U24888 (N_24888,N_23327,N_23940);
or U24889 (N_24889,N_23239,N_23478);
xor U24890 (N_24890,N_23935,N_23546);
or U24891 (N_24891,N_23624,N_23776);
and U24892 (N_24892,N_23780,N_23430);
nand U24893 (N_24893,N_23192,N_23980);
xnor U24894 (N_24894,N_23166,N_23056);
and U24895 (N_24895,N_23033,N_23870);
xor U24896 (N_24896,N_23460,N_23121);
or U24897 (N_24897,N_23583,N_23701);
or U24898 (N_24898,N_23084,N_23455);
nand U24899 (N_24899,N_23960,N_23033);
and U24900 (N_24900,N_23900,N_23067);
or U24901 (N_24901,N_23581,N_23330);
nand U24902 (N_24902,N_23920,N_23687);
and U24903 (N_24903,N_23880,N_23628);
nor U24904 (N_24904,N_23174,N_23254);
nor U24905 (N_24905,N_23023,N_23290);
nor U24906 (N_24906,N_23806,N_23918);
nand U24907 (N_24907,N_23425,N_23183);
or U24908 (N_24908,N_23847,N_23601);
nor U24909 (N_24909,N_23315,N_23347);
nor U24910 (N_24910,N_23103,N_23098);
nand U24911 (N_24911,N_23356,N_23483);
xnor U24912 (N_24912,N_23413,N_23144);
or U24913 (N_24913,N_23529,N_23719);
xor U24914 (N_24914,N_23454,N_23908);
xor U24915 (N_24915,N_23187,N_23607);
xnor U24916 (N_24916,N_23545,N_23446);
nand U24917 (N_24917,N_23437,N_23305);
and U24918 (N_24918,N_23446,N_23086);
and U24919 (N_24919,N_23118,N_23182);
or U24920 (N_24920,N_23669,N_23989);
xnor U24921 (N_24921,N_23859,N_23372);
nand U24922 (N_24922,N_23664,N_23237);
nand U24923 (N_24923,N_23527,N_23998);
and U24924 (N_24924,N_23157,N_23108);
and U24925 (N_24925,N_23279,N_23353);
or U24926 (N_24926,N_23485,N_23834);
and U24927 (N_24927,N_23766,N_23566);
nand U24928 (N_24928,N_23988,N_23985);
nand U24929 (N_24929,N_23602,N_23894);
or U24930 (N_24930,N_23840,N_23139);
and U24931 (N_24931,N_23624,N_23298);
nor U24932 (N_24932,N_23080,N_23277);
or U24933 (N_24933,N_23751,N_23299);
xnor U24934 (N_24934,N_23763,N_23833);
xnor U24935 (N_24935,N_23927,N_23027);
nand U24936 (N_24936,N_23764,N_23436);
nand U24937 (N_24937,N_23132,N_23436);
xnor U24938 (N_24938,N_23605,N_23467);
xor U24939 (N_24939,N_23721,N_23259);
or U24940 (N_24940,N_23945,N_23627);
or U24941 (N_24941,N_23467,N_23148);
and U24942 (N_24942,N_23933,N_23257);
or U24943 (N_24943,N_23157,N_23992);
xnor U24944 (N_24944,N_23402,N_23865);
or U24945 (N_24945,N_23729,N_23535);
or U24946 (N_24946,N_23760,N_23865);
xnor U24947 (N_24947,N_23479,N_23434);
and U24948 (N_24948,N_23562,N_23134);
nor U24949 (N_24949,N_23902,N_23575);
nand U24950 (N_24950,N_23075,N_23232);
xnor U24951 (N_24951,N_23260,N_23076);
xor U24952 (N_24952,N_23478,N_23043);
nor U24953 (N_24953,N_23317,N_23069);
and U24954 (N_24954,N_23853,N_23396);
nand U24955 (N_24955,N_23792,N_23023);
nand U24956 (N_24956,N_23809,N_23051);
or U24957 (N_24957,N_23658,N_23279);
nand U24958 (N_24958,N_23447,N_23955);
nor U24959 (N_24959,N_23303,N_23412);
and U24960 (N_24960,N_23253,N_23527);
xnor U24961 (N_24961,N_23672,N_23795);
xnor U24962 (N_24962,N_23799,N_23819);
or U24963 (N_24963,N_23528,N_23745);
nor U24964 (N_24964,N_23841,N_23949);
and U24965 (N_24965,N_23375,N_23602);
nand U24966 (N_24966,N_23818,N_23545);
and U24967 (N_24967,N_23913,N_23491);
xnor U24968 (N_24968,N_23680,N_23016);
and U24969 (N_24969,N_23650,N_23699);
xor U24970 (N_24970,N_23497,N_23822);
or U24971 (N_24971,N_23043,N_23388);
nor U24972 (N_24972,N_23274,N_23633);
nor U24973 (N_24973,N_23993,N_23150);
nand U24974 (N_24974,N_23908,N_23635);
and U24975 (N_24975,N_23480,N_23312);
nand U24976 (N_24976,N_23663,N_23852);
nor U24977 (N_24977,N_23792,N_23255);
or U24978 (N_24978,N_23058,N_23770);
and U24979 (N_24979,N_23457,N_23932);
nor U24980 (N_24980,N_23086,N_23571);
nor U24981 (N_24981,N_23063,N_23604);
nor U24982 (N_24982,N_23655,N_23683);
nand U24983 (N_24983,N_23828,N_23700);
nand U24984 (N_24984,N_23994,N_23728);
or U24985 (N_24985,N_23049,N_23127);
or U24986 (N_24986,N_23284,N_23312);
or U24987 (N_24987,N_23745,N_23093);
nand U24988 (N_24988,N_23306,N_23280);
nor U24989 (N_24989,N_23231,N_23799);
nand U24990 (N_24990,N_23388,N_23098);
nor U24991 (N_24991,N_23552,N_23625);
nand U24992 (N_24992,N_23137,N_23943);
xnor U24993 (N_24993,N_23928,N_23458);
or U24994 (N_24994,N_23688,N_23711);
nand U24995 (N_24995,N_23756,N_23622);
or U24996 (N_24996,N_23675,N_23822);
xor U24997 (N_24997,N_23202,N_23179);
xnor U24998 (N_24998,N_23584,N_23142);
xor U24999 (N_24999,N_23070,N_23038);
and UO_0 (O_0,N_24979,N_24845);
and UO_1 (O_1,N_24082,N_24169);
or UO_2 (O_2,N_24801,N_24482);
and UO_3 (O_3,N_24199,N_24194);
and UO_4 (O_4,N_24192,N_24548);
nor UO_5 (O_5,N_24704,N_24505);
and UO_6 (O_6,N_24654,N_24069);
nand UO_7 (O_7,N_24418,N_24003);
nand UO_8 (O_8,N_24464,N_24282);
and UO_9 (O_9,N_24636,N_24989);
nand UO_10 (O_10,N_24036,N_24817);
nand UO_11 (O_11,N_24029,N_24735);
or UO_12 (O_12,N_24998,N_24869);
nand UO_13 (O_13,N_24070,N_24853);
nor UO_14 (O_14,N_24965,N_24374);
xnor UO_15 (O_15,N_24190,N_24369);
xor UO_16 (O_16,N_24818,N_24838);
or UO_17 (O_17,N_24427,N_24837);
nand UO_18 (O_18,N_24034,N_24090);
or UO_19 (O_19,N_24014,N_24479);
xor UO_20 (O_20,N_24571,N_24132);
nor UO_21 (O_21,N_24920,N_24432);
nor UO_22 (O_22,N_24330,N_24612);
xnor UO_23 (O_23,N_24906,N_24545);
or UO_24 (O_24,N_24809,N_24327);
nor UO_25 (O_25,N_24737,N_24325);
or UO_26 (O_26,N_24902,N_24883);
or UO_27 (O_27,N_24272,N_24512);
xnor UO_28 (O_28,N_24580,N_24791);
nor UO_29 (O_29,N_24614,N_24072);
and UO_30 (O_30,N_24573,N_24969);
nand UO_31 (O_31,N_24716,N_24581);
xor UO_32 (O_32,N_24147,N_24298);
or UO_33 (O_33,N_24059,N_24910);
xnor UO_34 (O_34,N_24492,N_24160);
or UO_35 (O_35,N_24008,N_24865);
xor UO_36 (O_36,N_24745,N_24814);
and UO_37 (O_37,N_24625,N_24359);
nand UO_38 (O_38,N_24100,N_24113);
xnor UO_39 (O_39,N_24261,N_24894);
nand UO_40 (O_40,N_24855,N_24110);
nor UO_41 (O_41,N_24225,N_24280);
nand UO_42 (O_42,N_24134,N_24552);
or UO_43 (O_43,N_24551,N_24347);
nand UO_44 (O_44,N_24019,N_24970);
nor UO_45 (O_45,N_24229,N_24044);
or UO_46 (O_46,N_24243,N_24462);
nor UO_47 (O_47,N_24365,N_24972);
xor UO_48 (O_48,N_24043,N_24651);
and UO_49 (O_49,N_24688,N_24286);
and UO_50 (O_50,N_24690,N_24712);
xor UO_51 (O_51,N_24670,N_24893);
nand UO_52 (O_52,N_24924,N_24143);
nor UO_53 (O_53,N_24981,N_24460);
nand UO_54 (O_54,N_24540,N_24398);
xor UO_55 (O_55,N_24278,N_24815);
nor UO_56 (O_56,N_24089,N_24615);
and UO_57 (O_57,N_24084,N_24351);
and UO_58 (O_58,N_24717,N_24494);
or UO_59 (O_59,N_24425,N_24810);
nand UO_60 (O_60,N_24237,N_24471);
nand UO_61 (O_61,N_24643,N_24589);
xor UO_62 (O_62,N_24976,N_24481);
nand UO_63 (O_63,N_24634,N_24267);
nor UO_64 (O_64,N_24642,N_24586);
xor UO_65 (O_65,N_24364,N_24146);
and UO_66 (O_66,N_24005,N_24181);
nor UO_67 (O_67,N_24734,N_24459);
or UO_68 (O_68,N_24748,N_24394);
nor UO_69 (O_69,N_24547,N_24054);
nand UO_70 (O_70,N_24456,N_24977);
or UO_71 (O_71,N_24684,N_24104);
xor UO_72 (O_72,N_24909,N_24385);
nor UO_73 (O_73,N_24379,N_24193);
xor UO_74 (O_74,N_24326,N_24944);
or UO_75 (O_75,N_24052,N_24081);
or UO_76 (O_76,N_24974,N_24322);
and UO_77 (O_77,N_24532,N_24824);
nor UO_78 (O_78,N_24339,N_24640);
nor UO_79 (O_79,N_24495,N_24496);
nor UO_80 (O_80,N_24045,N_24442);
nor UO_81 (O_81,N_24564,N_24161);
nor UO_82 (O_82,N_24117,N_24268);
nor UO_83 (O_83,N_24443,N_24644);
nand UO_84 (O_84,N_24918,N_24355);
or UO_85 (O_85,N_24046,N_24493);
and UO_86 (O_86,N_24483,N_24851);
xor UO_87 (O_87,N_24119,N_24277);
xnor UO_88 (O_88,N_24429,N_24395);
nor UO_89 (O_89,N_24303,N_24676);
nand UO_90 (O_90,N_24658,N_24451);
xnor UO_91 (O_91,N_24032,N_24685);
nor UO_92 (O_92,N_24795,N_24811);
nand UO_93 (O_93,N_24775,N_24677);
nor UO_94 (O_94,N_24919,N_24596);
nor UO_95 (O_95,N_24291,N_24118);
xnor UO_96 (O_96,N_24889,N_24997);
xor UO_97 (O_97,N_24234,N_24733);
xor UO_98 (O_98,N_24312,N_24189);
and UO_99 (O_99,N_24531,N_24057);
or UO_100 (O_100,N_24083,N_24230);
and UO_101 (O_101,N_24696,N_24021);
and UO_102 (O_102,N_24139,N_24254);
and UO_103 (O_103,N_24252,N_24561);
xor UO_104 (O_104,N_24660,N_24892);
nand UO_105 (O_105,N_24749,N_24144);
xnor UO_106 (O_106,N_24516,N_24341);
nand UO_107 (O_107,N_24773,N_24804);
and UO_108 (O_108,N_24752,N_24635);
nor UO_109 (O_109,N_24334,N_24458);
xor UO_110 (O_110,N_24687,N_24746);
xor UO_111 (O_111,N_24004,N_24202);
and UO_112 (O_112,N_24633,N_24060);
nor UO_113 (O_113,N_24832,N_24543);
nand UO_114 (O_114,N_24820,N_24714);
nand UO_115 (O_115,N_24890,N_24410);
nor UO_116 (O_116,N_24954,N_24539);
and UO_117 (O_117,N_24366,N_24904);
or UO_118 (O_118,N_24725,N_24433);
xnor UO_119 (O_119,N_24841,N_24629);
xor UO_120 (O_120,N_24628,N_24352);
or UO_121 (O_121,N_24928,N_24020);
and UO_122 (O_122,N_24662,N_24509);
nand UO_123 (O_123,N_24541,N_24363);
nor UO_124 (O_124,N_24127,N_24565);
xnor UO_125 (O_125,N_24729,N_24595);
nor UO_126 (O_126,N_24211,N_24111);
xnor UO_127 (O_127,N_24120,N_24793);
nor UO_128 (O_128,N_24491,N_24900);
or UO_129 (O_129,N_24416,N_24637);
or UO_130 (O_130,N_24231,N_24338);
or UO_131 (O_131,N_24171,N_24064);
nor UO_132 (O_132,N_24276,N_24835);
xor UO_133 (O_133,N_24472,N_24942);
and UO_134 (O_134,N_24137,N_24674);
xor UO_135 (O_135,N_24689,N_24393);
and UO_136 (O_136,N_24769,N_24881);
nor UO_137 (O_137,N_24450,N_24723);
and UO_138 (O_138,N_24345,N_24705);
and UO_139 (O_139,N_24220,N_24186);
or UO_140 (O_140,N_24309,N_24630);
or UO_141 (O_141,N_24321,N_24150);
nor UO_142 (O_142,N_24130,N_24774);
nor UO_143 (O_143,N_24441,N_24513);
nand UO_144 (O_144,N_24049,N_24927);
or UO_145 (O_145,N_24535,N_24026);
or UO_146 (O_146,N_24131,N_24736);
nand UO_147 (O_147,N_24911,N_24715);
xnor UO_148 (O_148,N_24408,N_24116);
nand UO_149 (O_149,N_24626,N_24686);
nor UO_150 (O_150,N_24031,N_24324);
or UO_151 (O_151,N_24527,N_24732);
xor UO_152 (O_152,N_24417,N_24183);
nand UO_153 (O_153,N_24740,N_24899);
nor UO_154 (O_154,N_24536,N_24444);
xor UO_155 (O_155,N_24062,N_24647);
xnor UO_156 (O_156,N_24649,N_24078);
nor UO_157 (O_157,N_24788,N_24343);
or UO_158 (O_158,N_24389,N_24165);
and UO_159 (O_159,N_24667,N_24681);
and UO_160 (O_160,N_24554,N_24148);
xor UO_161 (O_161,N_24831,N_24269);
xor UO_162 (O_162,N_24214,N_24528);
xnor UO_163 (O_163,N_24510,N_24203);
nand UO_164 (O_164,N_24999,N_24933);
or UO_165 (O_165,N_24271,N_24390);
or UO_166 (O_166,N_24848,N_24027);
nor UO_167 (O_167,N_24102,N_24273);
and UO_168 (O_168,N_24648,N_24164);
nand UO_169 (O_169,N_24163,N_24713);
nand UO_170 (O_170,N_24987,N_24097);
nand UO_171 (O_171,N_24124,N_24295);
nor UO_172 (O_172,N_24123,N_24145);
nor UO_173 (O_173,N_24270,N_24567);
and UO_174 (O_174,N_24958,N_24984);
nand UO_175 (O_175,N_24159,N_24784);
nand UO_176 (O_176,N_24995,N_24632);
or UO_177 (O_177,N_24091,N_24446);
nor UO_178 (O_178,N_24287,N_24138);
nor UO_179 (O_179,N_24764,N_24655);
or UO_180 (O_180,N_24711,N_24297);
and UO_181 (O_181,N_24317,N_24833);
nor UO_182 (O_182,N_24498,N_24821);
and UO_183 (O_183,N_24122,N_24357);
nand UO_184 (O_184,N_24665,N_24400);
xnor UO_185 (O_185,N_24682,N_24013);
xnor UO_186 (O_186,N_24420,N_24411);
and UO_187 (O_187,N_24973,N_24386);
or UO_188 (O_188,N_24358,N_24743);
or UO_189 (O_189,N_24010,N_24604);
nand UO_190 (O_190,N_24176,N_24434);
nand UO_191 (O_191,N_24659,N_24299);
and UO_192 (O_192,N_24870,N_24422);
xor UO_193 (O_193,N_24125,N_24405);
xnor UO_194 (O_194,N_24871,N_24264);
nor UO_195 (O_195,N_24945,N_24631);
nand UO_196 (O_196,N_24787,N_24772);
nor UO_197 (O_197,N_24938,N_24524);
nand UO_198 (O_198,N_24912,N_24867);
xnor UO_199 (O_199,N_24223,N_24862);
xor UO_200 (O_200,N_24693,N_24786);
or UO_201 (O_201,N_24075,N_24412);
and UO_202 (O_202,N_24467,N_24040);
nor UO_203 (O_203,N_24315,N_24609);
nand UO_204 (O_204,N_24461,N_24490);
xor UO_205 (O_205,N_24486,N_24766);
xnor UO_206 (O_206,N_24285,N_24426);
nor UO_207 (O_207,N_24511,N_24093);
and UO_208 (O_208,N_24988,N_24372);
nor UO_209 (O_209,N_24779,N_24799);
xor UO_210 (O_210,N_24859,N_24507);
xnor UO_211 (O_211,N_24092,N_24095);
nor UO_212 (O_212,N_24594,N_24088);
nand UO_213 (O_213,N_24328,N_24975);
or UO_214 (O_214,N_24308,N_24392);
and UO_215 (O_215,N_24797,N_24789);
nor UO_216 (O_216,N_24584,N_24863);
nor UO_217 (O_217,N_24048,N_24603);
xnor UO_218 (O_218,N_24200,N_24396);
or UO_219 (O_219,N_24218,N_24421);
and UO_220 (O_220,N_24323,N_24866);
nor UO_221 (O_221,N_24065,N_24949);
nand UO_222 (O_222,N_24167,N_24248);
or UO_223 (O_223,N_24534,N_24213);
or UO_224 (O_224,N_24114,N_24476);
or UO_225 (O_225,N_24279,N_24262);
and UO_226 (O_226,N_24915,N_24292);
xor UO_227 (O_227,N_24850,N_24652);
nand UO_228 (O_228,N_24166,N_24591);
xnor UO_229 (O_229,N_24336,N_24011);
xnor UO_230 (O_230,N_24439,N_24128);
nor UO_231 (O_231,N_24042,N_24205);
nor UO_232 (O_232,N_24738,N_24399);
xnor UO_233 (O_233,N_24101,N_24868);
xor UO_234 (O_234,N_24886,N_24239);
or UO_235 (O_235,N_24613,N_24575);
and UO_236 (O_236,N_24739,N_24963);
and UO_237 (O_237,N_24638,N_24699);
nand UO_238 (O_238,N_24402,N_24066);
or UO_239 (O_239,N_24695,N_24255);
nor UO_240 (O_240,N_24542,N_24506);
or UO_241 (O_241,N_24812,N_24103);
and UO_242 (O_242,N_24700,N_24593);
nor UO_243 (O_243,N_24901,N_24897);
nor UO_244 (O_244,N_24457,N_24721);
or UO_245 (O_245,N_24073,N_24950);
or UO_246 (O_246,N_24415,N_24071);
nor UO_247 (O_247,N_24521,N_24990);
nor UO_248 (O_248,N_24035,N_24844);
or UO_249 (O_249,N_24608,N_24503);
nor UO_250 (O_250,N_24546,N_24265);
nand UO_251 (O_251,N_24378,N_24468);
and UO_252 (O_252,N_24115,N_24196);
nand UO_253 (O_253,N_24435,N_24294);
nor UO_254 (O_254,N_24227,N_24217);
nor UO_255 (O_255,N_24597,N_24437);
nor UO_256 (O_256,N_24477,N_24618);
and UO_257 (O_257,N_24246,N_24522);
and UO_258 (O_258,N_24489,N_24023);
xor UO_259 (O_259,N_24611,N_24484);
xnor UO_260 (O_260,N_24041,N_24993);
xor UO_261 (O_261,N_24653,N_24570);
xor UO_262 (O_262,N_24179,N_24300);
xnor UO_263 (O_263,N_24932,N_24941);
or UO_264 (O_264,N_24807,N_24627);
or UO_265 (O_265,N_24133,N_24236);
and UO_266 (O_266,N_24056,N_24947);
nor UO_267 (O_267,N_24184,N_24290);
nand UO_268 (O_268,N_24852,N_24228);
xnor UO_269 (O_269,N_24606,N_24404);
xor UO_270 (O_270,N_24816,N_24639);
and UO_271 (O_271,N_24782,N_24302);
nand UO_272 (O_272,N_24158,N_24348);
xnor UO_273 (O_273,N_24770,N_24952);
or UO_274 (O_274,N_24533,N_24553);
or UO_275 (O_275,N_24079,N_24387);
nor UO_276 (O_276,N_24307,N_24985);
or UO_277 (O_277,N_24112,N_24657);
nand UO_278 (O_278,N_24210,N_24129);
or UO_279 (O_279,N_24051,N_24304);
and UO_280 (O_280,N_24473,N_24238);
nand UO_281 (O_281,N_24880,N_24908);
and UO_282 (O_282,N_24759,N_24525);
xor UO_283 (O_283,N_24602,N_24623);
xor UO_284 (O_284,N_24409,N_24961);
and UO_285 (O_285,N_24391,N_24560);
xor UO_286 (O_286,N_24703,N_24680);
xnor UO_287 (O_287,N_24275,N_24962);
nor UO_288 (O_288,N_24940,N_24215);
xnor UO_289 (O_289,N_24226,N_24666);
and UO_290 (O_290,N_24038,N_24331);
xnor UO_291 (O_291,N_24025,N_24724);
or UO_292 (O_292,N_24898,N_24397);
and UO_293 (O_293,N_24982,N_24173);
and UO_294 (O_294,N_24755,N_24563);
nor UO_295 (O_295,N_24293,N_24679);
nor UO_296 (O_296,N_24356,N_24247);
and UO_297 (O_297,N_24673,N_24605);
nand UO_298 (O_298,N_24731,N_24288);
nor UO_299 (O_299,N_24475,N_24376);
nor UO_300 (O_300,N_24747,N_24361);
or UO_301 (O_301,N_24424,N_24825);
or UO_302 (O_302,N_24861,N_24951);
or UO_303 (O_303,N_24469,N_24966);
and UO_304 (O_304,N_24926,N_24449);
nand UO_305 (O_305,N_24968,N_24790);
nor UO_306 (O_306,N_24502,N_24087);
or UO_307 (O_307,N_24562,N_24805);
nor UO_308 (O_308,N_24916,N_24796);
xnor UO_309 (O_309,N_24216,N_24518);
xnor UO_310 (O_310,N_24340,N_24140);
xnor UO_311 (O_311,N_24407,N_24156);
nor UO_312 (O_312,N_24346,N_24175);
and UO_313 (O_313,N_24669,N_24758);
and UO_314 (O_314,N_24577,N_24953);
nand UO_315 (O_315,N_24697,N_24109);
xnor UO_316 (O_316,N_24012,N_24403);
and UO_317 (O_317,N_24701,N_24879);
nor UO_318 (O_318,N_24702,N_24232);
and UO_319 (O_319,N_24470,N_24517);
or UO_320 (O_320,N_24624,N_24438);
and UO_321 (O_321,N_24619,N_24204);
nor UO_322 (O_322,N_24077,N_24878);
xnor UO_323 (O_323,N_24827,N_24730);
nand UO_324 (O_324,N_24576,N_24994);
nand UO_325 (O_325,N_24258,N_24126);
nor UO_326 (O_326,N_24305,N_24767);
or UO_327 (O_327,N_24971,N_24349);
nor UO_328 (O_328,N_24678,N_24206);
nand UO_329 (O_329,N_24182,N_24719);
or UO_330 (O_330,N_24251,N_24447);
and UO_331 (O_331,N_24884,N_24224);
or UO_332 (O_332,N_24319,N_24250);
or UO_333 (O_333,N_24936,N_24854);
or UO_334 (O_334,N_24785,N_24826);
or UO_335 (O_335,N_24930,N_24263);
and UO_336 (O_336,N_24980,N_24431);
nand UO_337 (O_337,N_24955,N_24537);
or UO_338 (O_338,N_24096,N_24530);
or UO_339 (O_339,N_24846,N_24007);
xnor UO_340 (O_340,N_24086,N_24550);
nand UO_341 (O_341,N_24440,N_24708);
nand UO_342 (O_342,N_24763,N_24592);
xor UO_343 (O_343,N_24006,N_24921);
nand UO_344 (O_344,N_24610,N_24157);
xor UO_345 (O_345,N_24937,N_24948);
nor UO_346 (O_346,N_24501,N_24320);
or UO_347 (O_347,N_24413,N_24939);
or UO_348 (O_348,N_24430,N_24474);
and UO_349 (O_349,N_24960,N_24284);
and UO_350 (O_350,N_24557,N_24368);
or UO_351 (O_351,N_24497,N_24842);
xor UO_352 (O_352,N_24555,N_24500);
xor UO_353 (O_353,N_24741,N_24519);
and UO_354 (O_354,N_24778,N_24212);
and UO_355 (O_355,N_24946,N_24423);
nor UO_356 (O_356,N_24621,N_24381);
nand UO_357 (O_357,N_24478,N_24219);
nor UO_358 (O_358,N_24362,N_24568);
and UO_359 (O_359,N_24872,N_24903);
and UO_360 (O_360,N_24105,N_24992);
xnor UO_361 (O_361,N_24983,N_24664);
nor UO_362 (O_362,N_24600,N_24843);
nand UO_363 (O_363,N_24463,N_24514);
nor UO_364 (O_364,N_24661,N_24860);
xor UO_365 (O_365,N_24485,N_24757);
xnor UO_366 (O_366,N_24722,N_24813);
and UO_367 (O_367,N_24380,N_24344);
nand UO_368 (O_368,N_24620,N_24819);
nor UO_369 (O_369,N_24149,N_24499);
and UO_370 (O_370,N_24245,N_24360);
or UO_371 (O_371,N_24375,N_24885);
nand UO_372 (O_372,N_24419,N_24201);
or UO_373 (O_373,N_24242,N_24296);
or UO_374 (O_374,N_24777,N_24726);
xnor UO_375 (O_375,N_24388,N_24780);
xor UO_376 (O_376,N_24266,N_24207);
nor UO_377 (O_377,N_24776,N_24698);
or UO_378 (O_378,N_24033,N_24771);
or UO_379 (O_379,N_24706,N_24174);
nand UO_380 (O_380,N_24488,N_24830);
or UO_381 (O_381,N_24221,N_24311);
xor UO_382 (O_382,N_24047,N_24922);
xor UO_383 (O_383,N_24466,N_24382);
or UO_384 (O_384,N_24935,N_24751);
nor UO_385 (O_385,N_24762,N_24259);
nor UO_386 (O_386,N_24847,N_24121);
or UO_387 (O_387,N_24544,N_24646);
and UO_388 (O_388,N_24142,N_24896);
nor UO_389 (O_389,N_24017,N_24170);
nor UO_390 (O_390,N_24016,N_24750);
nor UO_391 (O_391,N_24792,N_24768);
nor UO_392 (O_392,N_24337,N_24151);
nor UO_393 (O_393,N_24742,N_24335);
nand UO_394 (O_394,N_24281,N_24377);
nand UO_395 (O_395,N_24692,N_24350);
nand UO_396 (O_396,N_24967,N_24022);
nor UO_397 (O_397,N_24187,N_24480);
nand UO_398 (O_398,N_24914,N_24289);
or UO_399 (O_399,N_24015,N_24508);
xor UO_400 (O_400,N_24875,N_24839);
nand UO_401 (O_401,N_24858,N_24233);
or UO_402 (O_402,N_24188,N_24822);
nand UO_403 (O_403,N_24329,N_24578);
and UO_404 (O_404,N_24141,N_24197);
nand UO_405 (O_405,N_24249,N_24094);
nor UO_406 (O_406,N_24549,N_24943);
nor UO_407 (O_407,N_24931,N_24178);
or UO_408 (O_408,N_24063,N_24802);
nand UO_409 (O_409,N_24913,N_24882);
and UO_410 (O_410,N_24001,N_24556);
or UO_411 (O_411,N_24956,N_24857);
nor UO_412 (O_412,N_24760,N_24002);
nor UO_413 (O_413,N_24333,N_24452);
or UO_414 (O_414,N_24874,N_24195);
xnor UO_415 (O_415,N_24098,N_24876);
nand UO_416 (O_416,N_24616,N_24332);
or UO_417 (O_417,N_24436,N_24465);
nor UO_418 (O_418,N_24709,N_24907);
and UO_419 (O_419,N_24401,N_24316);
nand UO_420 (O_420,N_24691,N_24024);
and UO_421 (O_421,N_24753,N_24765);
and UO_422 (O_422,N_24917,N_24558);
nor UO_423 (O_423,N_24301,N_24836);
xnor UO_424 (O_424,N_24353,N_24783);
nor UO_425 (O_425,N_24198,N_24849);
nand UO_426 (O_426,N_24707,N_24136);
xnor UO_427 (O_427,N_24834,N_24099);
and UO_428 (O_428,N_24454,N_24504);
nand UO_429 (O_429,N_24959,N_24068);
xnor UO_430 (O_430,N_24318,N_24108);
nor UO_431 (O_431,N_24445,N_24185);
xor UO_432 (O_432,N_24756,N_24000);
and UO_433 (O_433,N_24342,N_24155);
nor UO_434 (O_434,N_24617,N_24283);
nor UO_435 (O_435,N_24168,N_24583);
nor UO_436 (O_436,N_24453,N_24253);
or UO_437 (O_437,N_24663,N_24240);
or UO_438 (O_438,N_24515,N_24055);
xor UO_439 (O_439,N_24569,N_24037);
nand UO_440 (O_440,N_24028,N_24566);
nor UO_441 (O_441,N_24367,N_24744);
or UO_442 (O_442,N_24106,N_24996);
xor UO_443 (O_443,N_24260,N_24856);
nand UO_444 (O_444,N_24803,N_24672);
and UO_445 (O_445,N_24683,N_24829);
xor UO_446 (O_446,N_24957,N_24823);
nand UO_447 (O_447,N_24671,N_24590);
xnor UO_448 (O_448,N_24828,N_24373);
and UO_449 (O_449,N_24162,N_24754);
xnor UO_450 (O_450,N_24053,N_24964);
and UO_451 (O_451,N_24622,N_24370);
and UO_452 (O_452,N_24306,N_24929);
or UO_453 (O_453,N_24180,N_24085);
nor UO_454 (O_454,N_24645,N_24191);
nand UO_455 (O_455,N_24076,N_24641);
and UO_456 (O_456,N_24154,N_24428);
nor UO_457 (O_457,N_24520,N_24067);
nor UO_458 (O_458,N_24840,N_24107);
and UO_459 (O_459,N_24761,N_24018);
or UO_460 (O_460,N_24009,N_24172);
and UO_461 (O_461,N_24274,N_24794);
or UO_462 (O_462,N_24383,N_24588);
nor UO_463 (O_463,N_24209,N_24864);
nor UO_464 (O_464,N_24986,N_24607);
nor UO_465 (O_465,N_24529,N_24177);
xnor UO_466 (O_466,N_24406,N_24257);
xnor UO_467 (O_467,N_24135,N_24256);
xnor UO_468 (O_468,N_24727,N_24222);
xor UO_469 (O_469,N_24934,N_24800);
xor UO_470 (O_470,N_24808,N_24030);
nand UO_471 (O_471,N_24244,N_24235);
xnor UO_472 (O_472,N_24877,N_24991);
nor UO_473 (O_473,N_24582,N_24559);
nand UO_474 (O_474,N_24873,N_24887);
nor UO_475 (O_475,N_24601,N_24978);
xnor UO_476 (O_476,N_24585,N_24905);
nor UO_477 (O_477,N_24058,N_24487);
nor UO_478 (O_478,N_24598,N_24574);
or UO_479 (O_479,N_24448,N_24538);
nand UO_480 (O_480,N_24523,N_24599);
and UO_481 (O_481,N_24241,N_24310);
nor UO_482 (O_482,N_24923,N_24080);
xor UO_483 (O_483,N_24039,N_24710);
or UO_484 (O_484,N_24152,N_24153);
nand UO_485 (O_485,N_24650,N_24384);
or UO_486 (O_486,N_24925,N_24781);
or UO_487 (O_487,N_24728,N_24414);
nand UO_488 (O_488,N_24720,N_24587);
xnor UO_489 (O_489,N_24656,N_24371);
nor UO_490 (O_490,N_24455,N_24572);
xor UO_491 (O_491,N_24354,N_24888);
or UO_492 (O_492,N_24694,N_24579);
nor UO_493 (O_493,N_24718,N_24675);
nor UO_494 (O_494,N_24208,N_24050);
or UO_495 (O_495,N_24798,N_24895);
or UO_496 (O_496,N_24313,N_24526);
or UO_497 (O_497,N_24074,N_24314);
nor UO_498 (O_498,N_24668,N_24061);
xor UO_499 (O_499,N_24891,N_24806);
nand UO_500 (O_500,N_24624,N_24417);
nand UO_501 (O_501,N_24860,N_24136);
nand UO_502 (O_502,N_24049,N_24501);
nand UO_503 (O_503,N_24856,N_24292);
nand UO_504 (O_504,N_24691,N_24861);
nor UO_505 (O_505,N_24137,N_24516);
or UO_506 (O_506,N_24839,N_24205);
xor UO_507 (O_507,N_24745,N_24093);
xnor UO_508 (O_508,N_24641,N_24060);
nand UO_509 (O_509,N_24251,N_24299);
or UO_510 (O_510,N_24820,N_24919);
nand UO_511 (O_511,N_24473,N_24391);
or UO_512 (O_512,N_24927,N_24268);
xnor UO_513 (O_513,N_24242,N_24790);
or UO_514 (O_514,N_24280,N_24130);
xnor UO_515 (O_515,N_24021,N_24425);
nand UO_516 (O_516,N_24799,N_24622);
and UO_517 (O_517,N_24333,N_24453);
nor UO_518 (O_518,N_24087,N_24363);
nand UO_519 (O_519,N_24554,N_24749);
xor UO_520 (O_520,N_24430,N_24573);
or UO_521 (O_521,N_24995,N_24912);
and UO_522 (O_522,N_24256,N_24396);
nor UO_523 (O_523,N_24175,N_24121);
nand UO_524 (O_524,N_24366,N_24961);
or UO_525 (O_525,N_24988,N_24882);
xor UO_526 (O_526,N_24639,N_24264);
and UO_527 (O_527,N_24055,N_24198);
and UO_528 (O_528,N_24458,N_24798);
nor UO_529 (O_529,N_24595,N_24750);
or UO_530 (O_530,N_24840,N_24630);
nor UO_531 (O_531,N_24444,N_24331);
xor UO_532 (O_532,N_24712,N_24182);
and UO_533 (O_533,N_24846,N_24981);
or UO_534 (O_534,N_24042,N_24214);
xor UO_535 (O_535,N_24941,N_24879);
xor UO_536 (O_536,N_24749,N_24377);
or UO_537 (O_537,N_24041,N_24243);
xnor UO_538 (O_538,N_24373,N_24151);
or UO_539 (O_539,N_24270,N_24524);
xor UO_540 (O_540,N_24740,N_24207);
xor UO_541 (O_541,N_24933,N_24400);
xnor UO_542 (O_542,N_24824,N_24992);
xnor UO_543 (O_543,N_24631,N_24508);
nor UO_544 (O_544,N_24128,N_24341);
or UO_545 (O_545,N_24748,N_24785);
nor UO_546 (O_546,N_24370,N_24114);
nand UO_547 (O_547,N_24706,N_24089);
and UO_548 (O_548,N_24880,N_24279);
or UO_549 (O_549,N_24258,N_24576);
xor UO_550 (O_550,N_24847,N_24380);
or UO_551 (O_551,N_24891,N_24871);
xor UO_552 (O_552,N_24981,N_24741);
nor UO_553 (O_553,N_24453,N_24522);
and UO_554 (O_554,N_24107,N_24858);
nor UO_555 (O_555,N_24437,N_24389);
or UO_556 (O_556,N_24272,N_24428);
nor UO_557 (O_557,N_24340,N_24143);
nand UO_558 (O_558,N_24658,N_24754);
and UO_559 (O_559,N_24045,N_24272);
nor UO_560 (O_560,N_24765,N_24560);
nor UO_561 (O_561,N_24050,N_24948);
or UO_562 (O_562,N_24434,N_24365);
nand UO_563 (O_563,N_24538,N_24145);
or UO_564 (O_564,N_24170,N_24382);
and UO_565 (O_565,N_24960,N_24800);
xnor UO_566 (O_566,N_24517,N_24153);
nand UO_567 (O_567,N_24223,N_24373);
or UO_568 (O_568,N_24403,N_24067);
nand UO_569 (O_569,N_24801,N_24117);
or UO_570 (O_570,N_24757,N_24094);
and UO_571 (O_571,N_24848,N_24983);
and UO_572 (O_572,N_24420,N_24000);
and UO_573 (O_573,N_24865,N_24770);
or UO_574 (O_574,N_24464,N_24317);
or UO_575 (O_575,N_24252,N_24550);
nor UO_576 (O_576,N_24658,N_24645);
xor UO_577 (O_577,N_24861,N_24820);
nor UO_578 (O_578,N_24114,N_24019);
nand UO_579 (O_579,N_24359,N_24008);
or UO_580 (O_580,N_24872,N_24831);
and UO_581 (O_581,N_24028,N_24586);
and UO_582 (O_582,N_24397,N_24970);
and UO_583 (O_583,N_24569,N_24560);
nand UO_584 (O_584,N_24212,N_24530);
and UO_585 (O_585,N_24446,N_24028);
nor UO_586 (O_586,N_24554,N_24638);
xnor UO_587 (O_587,N_24856,N_24136);
xor UO_588 (O_588,N_24682,N_24634);
nor UO_589 (O_589,N_24633,N_24359);
and UO_590 (O_590,N_24650,N_24969);
or UO_591 (O_591,N_24200,N_24495);
and UO_592 (O_592,N_24250,N_24172);
and UO_593 (O_593,N_24742,N_24553);
nand UO_594 (O_594,N_24064,N_24536);
nor UO_595 (O_595,N_24830,N_24606);
nand UO_596 (O_596,N_24459,N_24064);
and UO_597 (O_597,N_24288,N_24645);
or UO_598 (O_598,N_24752,N_24822);
and UO_599 (O_599,N_24305,N_24669);
nand UO_600 (O_600,N_24576,N_24134);
nor UO_601 (O_601,N_24020,N_24772);
xor UO_602 (O_602,N_24554,N_24409);
nor UO_603 (O_603,N_24695,N_24294);
or UO_604 (O_604,N_24749,N_24235);
nor UO_605 (O_605,N_24653,N_24405);
nand UO_606 (O_606,N_24480,N_24827);
xor UO_607 (O_607,N_24045,N_24041);
nand UO_608 (O_608,N_24717,N_24859);
and UO_609 (O_609,N_24145,N_24334);
nor UO_610 (O_610,N_24014,N_24130);
nor UO_611 (O_611,N_24313,N_24547);
nor UO_612 (O_612,N_24827,N_24749);
nor UO_613 (O_613,N_24143,N_24460);
or UO_614 (O_614,N_24271,N_24915);
xnor UO_615 (O_615,N_24899,N_24149);
or UO_616 (O_616,N_24591,N_24545);
or UO_617 (O_617,N_24110,N_24123);
nand UO_618 (O_618,N_24280,N_24730);
and UO_619 (O_619,N_24486,N_24615);
nor UO_620 (O_620,N_24481,N_24454);
nand UO_621 (O_621,N_24593,N_24414);
and UO_622 (O_622,N_24761,N_24330);
or UO_623 (O_623,N_24873,N_24177);
nand UO_624 (O_624,N_24131,N_24339);
or UO_625 (O_625,N_24135,N_24943);
nor UO_626 (O_626,N_24032,N_24339);
and UO_627 (O_627,N_24852,N_24232);
nand UO_628 (O_628,N_24994,N_24403);
or UO_629 (O_629,N_24500,N_24296);
nor UO_630 (O_630,N_24034,N_24462);
xnor UO_631 (O_631,N_24253,N_24877);
xor UO_632 (O_632,N_24620,N_24447);
xnor UO_633 (O_633,N_24206,N_24456);
nor UO_634 (O_634,N_24148,N_24793);
xnor UO_635 (O_635,N_24993,N_24525);
xor UO_636 (O_636,N_24253,N_24865);
nor UO_637 (O_637,N_24792,N_24695);
nor UO_638 (O_638,N_24729,N_24455);
and UO_639 (O_639,N_24247,N_24292);
nor UO_640 (O_640,N_24604,N_24167);
nand UO_641 (O_641,N_24852,N_24362);
nor UO_642 (O_642,N_24857,N_24519);
and UO_643 (O_643,N_24921,N_24029);
and UO_644 (O_644,N_24507,N_24529);
nand UO_645 (O_645,N_24023,N_24367);
or UO_646 (O_646,N_24832,N_24902);
nor UO_647 (O_647,N_24058,N_24231);
and UO_648 (O_648,N_24575,N_24386);
xor UO_649 (O_649,N_24723,N_24043);
or UO_650 (O_650,N_24219,N_24489);
nand UO_651 (O_651,N_24204,N_24557);
and UO_652 (O_652,N_24900,N_24526);
nor UO_653 (O_653,N_24036,N_24040);
and UO_654 (O_654,N_24866,N_24213);
and UO_655 (O_655,N_24169,N_24096);
xnor UO_656 (O_656,N_24157,N_24645);
xor UO_657 (O_657,N_24093,N_24399);
nand UO_658 (O_658,N_24938,N_24780);
nand UO_659 (O_659,N_24500,N_24617);
and UO_660 (O_660,N_24388,N_24190);
or UO_661 (O_661,N_24060,N_24293);
nor UO_662 (O_662,N_24513,N_24795);
nand UO_663 (O_663,N_24389,N_24052);
nand UO_664 (O_664,N_24387,N_24425);
or UO_665 (O_665,N_24653,N_24295);
nor UO_666 (O_666,N_24550,N_24228);
nor UO_667 (O_667,N_24443,N_24244);
and UO_668 (O_668,N_24935,N_24673);
or UO_669 (O_669,N_24945,N_24058);
xnor UO_670 (O_670,N_24022,N_24754);
nor UO_671 (O_671,N_24166,N_24037);
or UO_672 (O_672,N_24221,N_24775);
nor UO_673 (O_673,N_24138,N_24270);
and UO_674 (O_674,N_24995,N_24778);
and UO_675 (O_675,N_24463,N_24628);
nand UO_676 (O_676,N_24755,N_24120);
nand UO_677 (O_677,N_24915,N_24446);
and UO_678 (O_678,N_24475,N_24884);
nor UO_679 (O_679,N_24171,N_24198);
and UO_680 (O_680,N_24781,N_24001);
and UO_681 (O_681,N_24156,N_24412);
nor UO_682 (O_682,N_24719,N_24247);
xor UO_683 (O_683,N_24413,N_24030);
xnor UO_684 (O_684,N_24171,N_24164);
and UO_685 (O_685,N_24318,N_24908);
nand UO_686 (O_686,N_24416,N_24127);
and UO_687 (O_687,N_24557,N_24751);
or UO_688 (O_688,N_24528,N_24183);
xor UO_689 (O_689,N_24182,N_24550);
xor UO_690 (O_690,N_24660,N_24992);
nand UO_691 (O_691,N_24699,N_24289);
xor UO_692 (O_692,N_24606,N_24124);
xor UO_693 (O_693,N_24889,N_24563);
nand UO_694 (O_694,N_24517,N_24222);
or UO_695 (O_695,N_24318,N_24870);
nand UO_696 (O_696,N_24592,N_24834);
nand UO_697 (O_697,N_24381,N_24530);
and UO_698 (O_698,N_24317,N_24357);
xnor UO_699 (O_699,N_24868,N_24200);
xnor UO_700 (O_700,N_24216,N_24267);
or UO_701 (O_701,N_24534,N_24435);
xor UO_702 (O_702,N_24132,N_24411);
and UO_703 (O_703,N_24528,N_24953);
nor UO_704 (O_704,N_24152,N_24916);
and UO_705 (O_705,N_24088,N_24865);
nor UO_706 (O_706,N_24338,N_24853);
or UO_707 (O_707,N_24476,N_24388);
nand UO_708 (O_708,N_24662,N_24367);
and UO_709 (O_709,N_24662,N_24708);
xor UO_710 (O_710,N_24572,N_24359);
xor UO_711 (O_711,N_24639,N_24770);
and UO_712 (O_712,N_24622,N_24474);
nand UO_713 (O_713,N_24703,N_24035);
nand UO_714 (O_714,N_24741,N_24329);
nand UO_715 (O_715,N_24446,N_24110);
nand UO_716 (O_716,N_24118,N_24038);
nand UO_717 (O_717,N_24336,N_24408);
nor UO_718 (O_718,N_24041,N_24225);
xor UO_719 (O_719,N_24382,N_24080);
nor UO_720 (O_720,N_24330,N_24261);
and UO_721 (O_721,N_24876,N_24460);
or UO_722 (O_722,N_24355,N_24715);
nor UO_723 (O_723,N_24278,N_24240);
xor UO_724 (O_724,N_24684,N_24782);
xor UO_725 (O_725,N_24311,N_24907);
or UO_726 (O_726,N_24231,N_24317);
or UO_727 (O_727,N_24290,N_24356);
nand UO_728 (O_728,N_24166,N_24762);
nand UO_729 (O_729,N_24527,N_24430);
or UO_730 (O_730,N_24954,N_24853);
and UO_731 (O_731,N_24878,N_24046);
nand UO_732 (O_732,N_24362,N_24329);
xor UO_733 (O_733,N_24499,N_24746);
and UO_734 (O_734,N_24750,N_24794);
nand UO_735 (O_735,N_24261,N_24756);
nor UO_736 (O_736,N_24850,N_24588);
or UO_737 (O_737,N_24532,N_24061);
nor UO_738 (O_738,N_24900,N_24324);
nor UO_739 (O_739,N_24427,N_24155);
nand UO_740 (O_740,N_24249,N_24308);
nor UO_741 (O_741,N_24245,N_24220);
xnor UO_742 (O_742,N_24959,N_24105);
and UO_743 (O_743,N_24550,N_24425);
xor UO_744 (O_744,N_24035,N_24646);
or UO_745 (O_745,N_24959,N_24635);
or UO_746 (O_746,N_24987,N_24420);
or UO_747 (O_747,N_24127,N_24710);
xnor UO_748 (O_748,N_24534,N_24565);
xor UO_749 (O_749,N_24711,N_24840);
nor UO_750 (O_750,N_24670,N_24514);
xor UO_751 (O_751,N_24937,N_24955);
xor UO_752 (O_752,N_24848,N_24094);
or UO_753 (O_753,N_24164,N_24158);
nand UO_754 (O_754,N_24370,N_24658);
nand UO_755 (O_755,N_24071,N_24383);
or UO_756 (O_756,N_24598,N_24086);
xnor UO_757 (O_757,N_24152,N_24597);
and UO_758 (O_758,N_24419,N_24730);
and UO_759 (O_759,N_24494,N_24088);
nand UO_760 (O_760,N_24559,N_24977);
and UO_761 (O_761,N_24010,N_24313);
nor UO_762 (O_762,N_24819,N_24057);
and UO_763 (O_763,N_24467,N_24512);
or UO_764 (O_764,N_24563,N_24990);
nor UO_765 (O_765,N_24771,N_24686);
or UO_766 (O_766,N_24766,N_24506);
nor UO_767 (O_767,N_24864,N_24196);
or UO_768 (O_768,N_24324,N_24730);
xnor UO_769 (O_769,N_24883,N_24918);
or UO_770 (O_770,N_24275,N_24805);
or UO_771 (O_771,N_24359,N_24988);
and UO_772 (O_772,N_24674,N_24092);
nor UO_773 (O_773,N_24190,N_24486);
and UO_774 (O_774,N_24068,N_24585);
nor UO_775 (O_775,N_24721,N_24226);
xor UO_776 (O_776,N_24378,N_24066);
and UO_777 (O_777,N_24171,N_24676);
xnor UO_778 (O_778,N_24739,N_24924);
or UO_779 (O_779,N_24270,N_24536);
and UO_780 (O_780,N_24342,N_24513);
nand UO_781 (O_781,N_24805,N_24680);
or UO_782 (O_782,N_24465,N_24141);
nand UO_783 (O_783,N_24972,N_24168);
or UO_784 (O_784,N_24062,N_24488);
xnor UO_785 (O_785,N_24919,N_24184);
or UO_786 (O_786,N_24026,N_24187);
and UO_787 (O_787,N_24094,N_24307);
nand UO_788 (O_788,N_24909,N_24462);
xnor UO_789 (O_789,N_24023,N_24814);
and UO_790 (O_790,N_24345,N_24669);
nand UO_791 (O_791,N_24018,N_24424);
xnor UO_792 (O_792,N_24613,N_24428);
or UO_793 (O_793,N_24673,N_24034);
and UO_794 (O_794,N_24952,N_24789);
nor UO_795 (O_795,N_24951,N_24451);
nor UO_796 (O_796,N_24657,N_24940);
xor UO_797 (O_797,N_24814,N_24908);
nand UO_798 (O_798,N_24480,N_24108);
nor UO_799 (O_799,N_24786,N_24043);
xor UO_800 (O_800,N_24813,N_24519);
nand UO_801 (O_801,N_24178,N_24626);
nand UO_802 (O_802,N_24234,N_24541);
xnor UO_803 (O_803,N_24983,N_24642);
or UO_804 (O_804,N_24037,N_24233);
or UO_805 (O_805,N_24447,N_24464);
nor UO_806 (O_806,N_24390,N_24660);
nand UO_807 (O_807,N_24344,N_24959);
xnor UO_808 (O_808,N_24852,N_24073);
and UO_809 (O_809,N_24688,N_24160);
nor UO_810 (O_810,N_24306,N_24103);
and UO_811 (O_811,N_24475,N_24752);
nand UO_812 (O_812,N_24934,N_24388);
nor UO_813 (O_813,N_24910,N_24647);
and UO_814 (O_814,N_24829,N_24672);
nor UO_815 (O_815,N_24212,N_24382);
and UO_816 (O_816,N_24160,N_24716);
xor UO_817 (O_817,N_24308,N_24767);
xnor UO_818 (O_818,N_24388,N_24203);
xor UO_819 (O_819,N_24058,N_24950);
or UO_820 (O_820,N_24398,N_24231);
or UO_821 (O_821,N_24533,N_24912);
nand UO_822 (O_822,N_24035,N_24753);
xor UO_823 (O_823,N_24420,N_24553);
nor UO_824 (O_824,N_24821,N_24496);
or UO_825 (O_825,N_24985,N_24515);
and UO_826 (O_826,N_24824,N_24794);
nor UO_827 (O_827,N_24740,N_24121);
or UO_828 (O_828,N_24192,N_24867);
and UO_829 (O_829,N_24840,N_24950);
xnor UO_830 (O_830,N_24968,N_24197);
nor UO_831 (O_831,N_24939,N_24760);
xnor UO_832 (O_832,N_24635,N_24618);
nand UO_833 (O_833,N_24416,N_24883);
or UO_834 (O_834,N_24834,N_24703);
xor UO_835 (O_835,N_24758,N_24908);
and UO_836 (O_836,N_24184,N_24340);
or UO_837 (O_837,N_24422,N_24089);
nand UO_838 (O_838,N_24304,N_24876);
and UO_839 (O_839,N_24933,N_24131);
or UO_840 (O_840,N_24062,N_24206);
or UO_841 (O_841,N_24189,N_24474);
nor UO_842 (O_842,N_24764,N_24858);
xor UO_843 (O_843,N_24213,N_24005);
or UO_844 (O_844,N_24636,N_24185);
nor UO_845 (O_845,N_24025,N_24838);
or UO_846 (O_846,N_24330,N_24023);
or UO_847 (O_847,N_24436,N_24717);
or UO_848 (O_848,N_24540,N_24567);
xnor UO_849 (O_849,N_24522,N_24262);
or UO_850 (O_850,N_24257,N_24748);
nor UO_851 (O_851,N_24019,N_24827);
xor UO_852 (O_852,N_24914,N_24224);
and UO_853 (O_853,N_24925,N_24495);
nor UO_854 (O_854,N_24340,N_24718);
xor UO_855 (O_855,N_24362,N_24234);
xnor UO_856 (O_856,N_24855,N_24854);
or UO_857 (O_857,N_24980,N_24938);
xnor UO_858 (O_858,N_24106,N_24943);
and UO_859 (O_859,N_24042,N_24443);
nand UO_860 (O_860,N_24573,N_24252);
nor UO_861 (O_861,N_24517,N_24866);
nor UO_862 (O_862,N_24586,N_24249);
xor UO_863 (O_863,N_24500,N_24434);
and UO_864 (O_864,N_24739,N_24244);
and UO_865 (O_865,N_24903,N_24727);
nor UO_866 (O_866,N_24332,N_24179);
and UO_867 (O_867,N_24909,N_24262);
and UO_868 (O_868,N_24007,N_24888);
and UO_869 (O_869,N_24332,N_24449);
nand UO_870 (O_870,N_24840,N_24823);
xnor UO_871 (O_871,N_24920,N_24004);
xnor UO_872 (O_872,N_24137,N_24812);
or UO_873 (O_873,N_24397,N_24196);
nand UO_874 (O_874,N_24783,N_24127);
and UO_875 (O_875,N_24993,N_24369);
nand UO_876 (O_876,N_24584,N_24353);
nand UO_877 (O_877,N_24853,N_24274);
nand UO_878 (O_878,N_24507,N_24412);
and UO_879 (O_879,N_24288,N_24469);
or UO_880 (O_880,N_24114,N_24105);
or UO_881 (O_881,N_24599,N_24250);
and UO_882 (O_882,N_24280,N_24911);
and UO_883 (O_883,N_24482,N_24922);
and UO_884 (O_884,N_24423,N_24007);
and UO_885 (O_885,N_24727,N_24040);
and UO_886 (O_886,N_24764,N_24830);
and UO_887 (O_887,N_24408,N_24251);
xor UO_888 (O_888,N_24554,N_24923);
nand UO_889 (O_889,N_24252,N_24464);
and UO_890 (O_890,N_24638,N_24788);
and UO_891 (O_891,N_24286,N_24796);
or UO_892 (O_892,N_24757,N_24421);
xnor UO_893 (O_893,N_24008,N_24831);
or UO_894 (O_894,N_24450,N_24417);
or UO_895 (O_895,N_24569,N_24730);
nand UO_896 (O_896,N_24354,N_24362);
nor UO_897 (O_897,N_24590,N_24930);
and UO_898 (O_898,N_24138,N_24715);
or UO_899 (O_899,N_24430,N_24941);
and UO_900 (O_900,N_24199,N_24661);
xnor UO_901 (O_901,N_24292,N_24116);
xnor UO_902 (O_902,N_24999,N_24242);
or UO_903 (O_903,N_24275,N_24378);
xnor UO_904 (O_904,N_24490,N_24295);
or UO_905 (O_905,N_24260,N_24889);
nand UO_906 (O_906,N_24983,N_24924);
xor UO_907 (O_907,N_24706,N_24517);
and UO_908 (O_908,N_24210,N_24086);
or UO_909 (O_909,N_24594,N_24960);
xor UO_910 (O_910,N_24664,N_24752);
nand UO_911 (O_911,N_24613,N_24722);
or UO_912 (O_912,N_24795,N_24529);
xnor UO_913 (O_913,N_24454,N_24386);
nor UO_914 (O_914,N_24873,N_24545);
nor UO_915 (O_915,N_24913,N_24074);
nor UO_916 (O_916,N_24762,N_24872);
xor UO_917 (O_917,N_24116,N_24030);
nand UO_918 (O_918,N_24526,N_24221);
xor UO_919 (O_919,N_24445,N_24229);
or UO_920 (O_920,N_24951,N_24681);
and UO_921 (O_921,N_24422,N_24508);
nor UO_922 (O_922,N_24929,N_24051);
and UO_923 (O_923,N_24236,N_24337);
xnor UO_924 (O_924,N_24457,N_24820);
and UO_925 (O_925,N_24693,N_24800);
or UO_926 (O_926,N_24221,N_24918);
xnor UO_927 (O_927,N_24923,N_24796);
and UO_928 (O_928,N_24425,N_24250);
nor UO_929 (O_929,N_24153,N_24068);
xnor UO_930 (O_930,N_24450,N_24670);
and UO_931 (O_931,N_24601,N_24241);
nand UO_932 (O_932,N_24452,N_24324);
xnor UO_933 (O_933,N_24187,N_24297);
and UO_934 (O_934,N_24451,N_24313);
nand UO_935 (O_935,N_24774,N_24726);
xor UO_936 (O_936,N_24175,N_24280);
or UO_937 (O_937,N_24242,N_24036);
nand UO_938 (O_938,N_24713,N_24149);
nor UO_939 (O_939,N_24401,N_24942);
and UO_940 (O_940,N_24326,N_24218);
nor UO_941 (O_941,N_24041,N_24024);
xnor UO_942 (O_942,N_24490,N_24074);
nand UO_943 (O_943,N_24343,N_24034);
and UO_944 (O_944,N_24837,N_24233);
nor UO_945 (O_945,N_24133,N_24267);
nand UO_946 (O_946,N_24911,N_24178);
xnor UO_947 (O_947,N_24846,N_24132);
or UO_948 (O_948,N_24360,N_24556);
or UO_949 (O_949,N_24671,N_24663);
or UO_950 (O_950,N_24791,N_24606);
nand UO_951 (O_951,N_24559,N_24153);
or UO_952 (O_952,N_24780,N_24072);
or UO_953 (O_953,N_24857,N_24731);
or UO_954 (O_954,N_24623,N_24782);
or UO_955 (O_955,N_24897,N_24648);
and UO_956 (O_956,N_24761,N_24027);
and UO_957 (O_957,N_24120,N_24987);
nand UO_958 (O_958,N_24208,N_24172);
nand UO_959 (O_959,N_24241,N_24439);
or UO_960 (O_960,N_24124,N_24343);
xor UO_961 (O_961,N_24926,N_24346);
nor UO_962 (O_962,N_24024,N_24187);
or UO_963 (O_963,N_24760,N_24032);
or UO_964 (O_964,N_24016,N_24615);
and UO_965 (O_965,N_24500,N_24683);
xnor UO_966 (O_966,N_24268,N_24462);
and UO_967 (O_967,N_24341,N_24130);
nand UO_968 (O_968,N_24176,N_24592);
nor UO_969 (O_969,N_24841,N_24590);
and UO_970 (O_970,N_24479,N_24676);
nand UO_971 (O_971,N_24077,N_24286);
nand UO_972 (O_972,N_24725,N_24453);
and UO_973 (O_973,N_24692,N_24826);
nor UO_974 (O_974,N_24077,N_24791);
nor UO_975 (O_975,N_24548,N_24682);
and UO_976 (O_976,N_24056,N_24411);
nor UO_977 (O_977,N_24425,N_24685);
nor UO_978 (O_978,N_24863,N_24625);
and UO_979 (O_979,N_24563,N_24242);
xnor UO_980 (O_980,N_24691,N_24763);
xor UO_981 (O_981,N_24117,N_24870);
nand UO_982 (O_982,N_24951,N_24029);
nor UO_983 (O_983,N_24765,N_24464);
nor UO_984 (O_984,N_24910,N_24921);
or UO_985 (O_985,N_24931,N_24341);
nand UO_986 (O_986,N_24660,N_24656);
nor UO_987 (O_987,N_24175,N_24600);
or UO_988 (O_988,N_24402,N_24355);
and UO_989 (O_989,N_24034,N_24499);
nor UO_990 (O_990,N_24810,N_24457);
and UO_991 (O_991,N_24457,N_24428);
or UO_992 (O_992,N_24889,N_24455);
nor UO_993 (O_993,N_24249,N_24651);
xnor UO_994 (O_994,N_24998,N_24598);
and UO_995 (O_995,N_24004,N_24147);
nor UO_996 (O_996,N_24287,N_24001);
nor UO_997 (O_997,N_24350,N_24169);
xnor UO_998 (O_998,N_24488,N_24277);
nand UO_999 (O_999,N_24065,N_24618);
nand UO_1000 (O_1000,N_24352,N_24300);
nor UO_1001 (O_1001,N_24398,N_24471);
and UO_1002 (O_1002,N_24561,N_24352);
and UO_1003 (O_1003,N_24547,N_24137);
nor UO_1004 (O_1004,N_24831,N_24474);
or UO_1005 (O_1005,N_24897,N_24507);
nand UO_1006 (O_1006,N_24591,N_24158);
or UO_1007 (O_1007,N_24336,N_24938);
nor UO_1008 (O_1008,N_24154,N_24034);
and UO_1009 (O_1009,N_24244,N_24738);
and UO_1010 (O_1010,N_24485,N_24170);
nand UO_1011 (O_1011,N_24556,N_24528);
and UO_1012 (O_1012,N_24623,N_24418);
or UO_1013 (O_1013,N_24830,N_24070);
nand UO_1014 (O_1014,N_24683,N_24543);
and UO_1015 (O_1015,N_24720,N_24193);
and UO_1016 (O_1016,N_24480,N_24821);
nor UO_1017 (O_1017,N_24829,N_24947);
xor UO_1018 (O_1018,N_24747,N_24449);
nor UO_1019 (O_1019,N_24314,N_24477);
or UO_1020 (O_1020,N_24849,N_24981);
or UO_1021 (O_1021,N_24028,N_24104);
xor UO_1022 (O_1022,N_24320,N_24704);
xnor UO_1023 (O_1023,N_24060,N_24993);
and UO_1024 (O_1024,N_24891,N_24028);
xor UO_1025 (O_1025,N_24330,N_24704);
nand UO_1026 (O_1026,N_24838,N_24811);
and UO_1027 (O_1027,N_24778,N_24426);
and UO_1028 (O_1028,N_24635,N_24395);
or UO_1029 (O_1029,N_24278,N_24093);
nor UO_1030 (O_1030,N_24093,N_24662);
nand UO_1031 (O_1031,N_24504,N_24054);
nand UO_1032 (O_1032,N_24423,N_24950);
and UO_1033 (O_1033,N_24419,N_24120);
nand UO_1034 (O_1034,N_24174,N_24858);
xor UO_1035 (O_1035,N_24228,N_24235);
nor UO_1036 (O_1036,N_24292,N_24368);
xnor UO_1037 (O_1037,N_24329,N_24443);
nor UO_1038 (O_1038,N_24212,N_24117);
xor UO_1039 (O_1039,N_24304,N_24111);
nand UO_1040 (O_1040,N_24272,N_24867);
nand UO_1041 (O_1041,N_24995,N_24647);
xnor UO_1042 (O_1042,N_24813,N_24214);
or UO_1043 (O_1043,N_24455,N_24451);
or UO_1044 (O_1044,N_24012,N_24067);
nand UO_1045 (O_1045,N_24619,N_24262);
nor UO_1046 (O_1046,N_24148,N_24338);
nor UO_1047 (O_1047,N_24969,N_24122);
xnor UO_1048 (O_1048,N_24916,N_24213);
nand UO_1049 (O_1049,N_24057,N_24031);
and UO_1050 (O_1050,N_24549,N_24021);
nand UO_1051 (O_1051,N_24834,N_24210);
xnor UO_1052 (O_1052,N_24550,N_24628);
and UO_1053 (O_1053,N_24898,N_24979);
and UO_1054 (O_1054,N_24974,N_24846);
nor UO_1055 (O_1055,N_24735,N_24086);
or UO_1056 (O_1056,N_24575,N_24168);
xnor UO_1057 (O_1057,N_24874,N_24093);
xnor UO_1058 (O_1058,N_24168,N_24516);
nor UO_1059 (O_1059,N_24046,N_24460);
and UO_1060 (O_1060,N_24722,N_24593);
xor UO_1061 (O_1061,N_24127,N_24002);
xnor UO_1062 (O_1062,N_24103,N_24973);
and UO_1063 (O_1063,N_24236,N_24092);
or UO_1064 (O_1064,N_24868,N_24447);
nor UO_1065 (O_1065,N_24518,N_24185);
nor UO_1066 (O_1066,N_24065,N_24337);
and UO_1067 (O_1067,N_24184,N_24156);
and UO_1068 (O_1068,N_24392,N_24127);
and UO_1069 (O_1069,N_24209,N_24747);
or UO_1070 (O_1070,N_24769,N_24297);
nor UO_1071 (O_1071,N_24776,N_24612);
and UO_1072 (O_1072,N_24293,N_24953);
and UO_1073 (O_1073,N_24010,N_24504);
nor UO_1074 (O_1074,N_24910,N_24384);
or UO_1075 (O_1075,N_24622,N_24659);
nand UO_1076 (O_1076,N_24120,N_24055);
and UO_1077 (O_1077,N_24687,N_24084);
nor UO_1078 (O_1078,N_24351,N_24205);
xnor UO_1079 (O_1079,N_24247,N_24254);
or UO_1080 (O_1080,N_24920,N_24441);
nor UO_1081 (O_1081,N_24661,N_24105);
or UO_1082 (O_1082,N_24935,N_24667);
and UO_1083 (O_1083,N_24378,N_24402);
and UO_1084 (O_1084,N_24725,N_24143);
xor UO_1085 (O_1085,N_24784,N_24382);
or UO_1086 (O_1086,N_24108,N_24571);
or UO_1087 (O_1087,N_24473,N_24127);
xnor UO_1088 (O_1088,N_24649,N_24705);
and UO_1089 (O_1089,N_24143,N_24516);
nor UO_1090 (O_1090,N_24489,N_24720);
and UO_1091 (O_1091,N_24332,N_24491);
nand UO_1092 (O_1092,N_24449,N_24342);
xnor UO_1093 (O_1093,N_24993,N_24972);
xor UO_1094 (O_1094,N_24401,N_24126);
or UO_1095 (O_1095,N_24110,N_24063);
nand UO_1096 (O_1096,N_24097,N_24984);
and UO_1097 (O_1097,N_24220,N_24584);
xor UO_1098 (O_1098,N_24017,N_24359);
nand UO_1099 (O_1099,N_24542,N_24031);
or UO_1100 (O_1100,N_24197,N_24561);
nor UO_1101 (O_1101,N_24808,N_24886);
and UO_1102 (O_1102,N_24159,N_24423);
or UO_1103 (O_1103,N_24522,N_24813);
nand UO_1104 (O_1104,N_24953,N_24617);
xnor UO_1105 (O_1105,N_24810,N_24684);
or UO_1106 (O_1106,N_24507,N_24154);
xor UO_1107 (O_1107,N_24357,N_24065);
and UO_1108 (O_1108,N_24047,N_24667);
and UO_1109 (O_1109,N_24496,N_24671);
or UO_1110 (O_1110,N_24935,N_24312);
nand UO_1111 (O_1111,N_24771,N_24569);
and UO_1112 (O_1112,N_24425,N_24552);
nor UO_1113 (O_1113,N_24870,N_24910);
or UO_1114 (O_1114,N_24455,N_24840);
nand UO_1115 (O_1115,N_24254,N_24064);
or UO_1116 (O_1116,N_24552,N_24518);
and UO_1117 (O_1117,N_24109,N_24002);
xor UO_1118 (O_1118,N_24976,N_24974);
nor UO_1119 (O_1119,N_24406,N_24374);
xnor UO_1120 (O_1120,N_24261,N_24092);
nand UO_1121 (O_1121,N_24440,N_24083);
or UO_1122 (O_1122,N_24783,N_24646);
and UO_1123 (O_1123,N_24951,N_24397);
nand UO_1124 (O_1124,N_24999,N_24338);
nor UO_1125 (O_1125,N_24792,N_24298);
nor UO_1126 (O_1126,N_24664,N_24055);
or UO_1127 (O_1127,N_24074,N_24401);
xnor UO_1128 (O_1128,N_24813,N_24142);
xor UO_1129 (O_1129,N_24330,N_24260);
or UO_1130 (O_1130,N_24865,N_24342);
nand UO_1131 (O_1131,N_24069,N_24017);
or UO_1132 (O_1132,N_24391,N_24737);
nor UO_1133 (O_1133,N_24812,N_24848);
or UO_1134 (O_1134,N_24050,N_24739);
or UO_1135 (O_1135,N_24139,N_24090);
and UO_1136 (O_1136,N_24047,N_24737);
nor UO_1137 (O_1137,N_24997,N_24532);
nor UO_1138 (O_1138,N_24944,N_24366);
and UO_1139 (O_1139,N_24816,N_24844);
nor UO_1140 (O_1140,N_24849,N_24421);
xnor UO_1141 (O_1141,N_24958,N_24145);
or UO_1142 (O_1142,N_24049,N_24314);
nand UO_1143 (O_1143,N_24103,N_24304);
nor UO_1144 (O_1144,N_24248,N_24762);
nor UO_1145 (O_1145,N_24365,N_24984);
xnor UO_1146 (O_1146,N_24525,N_24960);
and UO_1147 (O_1147,N_24226,N_24151);
nand UO_1148 (O_1148,N_24183,N_24512);
and UO_1149 (O_1149,N_24251,N_24939);
nand UO_1150 (O_1150,N_24072,N_24286);
or UO_1151 (O_1151,N_24383,N_24459);
nor UO_1152 (O_1152,N_24099,N_24343);
and UO_1153 (O_1153,N_24335,N_24306);
nand UO_1154 (O_1154,N_24209,N_24517);
nand UO_1155 (O_1155,N_24852,N_24240);
and UO_1156 (O_1156,N_24921,N_24180);
or UO_1157 (O_1157,N_24061,N_24305);
nand UO_1158 (O_1158,N_24279,N_24306);
and UO_1159 (O_1159,N_24618,N_24093);
nor UO_1160 (O_1160,N_24363,N_24493);
and UO_1161 (O_1161,N_24839,N_24257);
nand UO_1162 (O_1162,N_24391,N_24638);
or UO_1163 (O_1163,N_24701,N_24413);
and UO_1164 (O_1164,N_24188,N_24573);
nor UO_1165 (O_1165,N_24542,N_24955);
nor UO_1166 (O_1166,N_24083,N_24939);
xor UO_1167 (O_1167,N_24742,N_24174);
and UO_1168 (O_1168,N_24091,N_24142);
xnor UO_1169 (O_1169,N_24340,N_24156);
xor UO_1170 (O_1170,N_24033,N_24166);
xnor UO_1171 (O_1171,N_24273,N_24326);
or UO_1172 (O_1172,N_24751,N_24957);
or UO_1173 (O_1173,N_24501,N_24445);
xor UO_1174 (O_1174,N_24538,N_24321);
xor UO_1175 (O_1175,N_24130,N_24672);
nand UO_1176 (O_1176,N_24506,N_24990);
nand UO_1177 (O_1177,N_24234,N_24383);
or UO_1178 (O_1178,N_24290,N_24150);
nand UO_1179 (O_1179,N_24117,N_24561);
or UO_1180 (O_1180,N_24691,N_24203);
or UO_1181 (O_1181,N_24068,N_24703);
nor UO_1182 (O_1182,N_24757,N_24808);
xnor UO_1183 (O_1183,N_24357,N_24425);
nand UO_1184 (O_1184,N_24332,N_24117);
or UO_1185 (O_1185,N_24501,N_24010);
or UO_1186 (O_1186,N_24916,N_24541);
nand UO_1187 (O_1187,N_24325,N_24558);
nor UO_1188 (O_1188,N_24973,N_24799);
nor UO_1189 (O_1189,N_24878,N_24483);
and UO_1190 (O_1190,N_24430,N_24850);
and UO_1191 (O_1191,N_24087,N_24055);
nor UO_1192 (O_1192,N_24789,N_24520);
and UO_1193 (O_1193,N_24315,N_24039);
xor UO_1194 (O_1194,N_24961,N_24499);
nor UO_1195 (O_1195,N_24359,N_24546);
and UO_1196 (O_1196,N_24927,N_24274);
or UO_1197 (O_1197,N_24065,N_24945);
and UO_1198 (O_1198,N_24748,N_24187);
and UO_1199 (O_1199,N_24889,N_24363);
xnor UO_1200 (O_1200,N_24915,N_24803);
and UO_1201 (O_1201,N_24530,N_24902);
nand UO_1202 (O_1202,N_24278,N_24921);
xor UO_1203 (O_1203,N_24867,N_24321);
nand UO_1204 (O_1204,N_24459,N_24429);
xor UO_1205 (O_1205,N_24753,N_24532);
xor UO_1206 (O_1206,N_24918,N_24364);
and UO_1207 (O_1207,N_24893,N_24975);
or UO_1208 (O_1208,N_24679,N_24988);
xnor UO_1209 (O_1209,N_24563,N_24100);
or UO_1210 (O_1210,N_24751,N_24041);
and UO_1211 (O_1211,N_24984,N_24945);
nand UO_1212 (O_1212,N_24436,N_24323);
nand UO_1213 (O_1213,N_24447,N_24580);
nand UO_1214 (O_1214,N_24513,N_24171);
nor UO_1215 (O_1215,N_24645,N_24188);
nand UO_1216 (O_1216,N_24440,N_24374);
or UO_1217 (O_1217,N_24271,N_24423);
and UO_1218 (O_1218,N_24248,N_24730);
and UO_1219 (O_1219,N_24230,N_24580);
xnor UO_1220 (O_1220,N_24289,N_24084);
xnor UO_1221 (O_1221,N_24129,N_24233);
xnor UO_1222 (O_1222,N_24517,N_24851);
xor UO_1223 (O_1223,N_24897,N_24183);
or UO_1224 (O_1224,N_24575,N_24056);
and UO_1225 (O_1225,N_24781,N_24095);
and UO_1226 (O_1226,N_24407,N_24185);
nand UO_1227 (O_1227,N_24769,N_24761);
xnor UO_1228 (O_1228,N_24036,N_24240);
xnor UO_1229 (O_1229,N_24635,N_24271);
nand UO_1230 (O_1230,N_24847,N_24169);
nand UO_1231 (O_1231,N_24253,N_24354);
nor UO_1232 (O_1232,N_24318,N_24113);
or UO_1233 (O_1233,N_24986,N_24034);
and UO_1234 (O_1234,N_24166,N_24693);
nand UO_1235 (O_1235,N_24799,N_24929);
or UO_1236 (O_1236,N_24313,N_24858);
xnor UO_1237 (O_1237,N_24178,N_24756);
nand UO_1238 (O_1238,N_24260,N_24796);
and UO_1239 (O_1239,N_24513,N_24328);
nor UO_1240 (O_1240,N_24305,N_24092);
nand UO_1241 (O_1241,N_24660,N_24969);
or UO_1242 (O_1242,N_24413,N_24698);
nand UO_1243 (O_1243,N_24494,N_24318);
nand UO_1244 (O_1244,N_24389,N_24906);
nor UO_1245 (O_1245,N_24311,N_24879);
nand UO_1246 (O_1246,N_24170,N_24841);
nand UO_1247 (O_1247,N_24532,N_24739);
xor UO_1248 (O_1248,N_24232,N_24425);
xor UO_1249 (O_1249,N_24671,N_24168);
and UO_1250 (O_1250,N_24433,N_24510);
or UO_1251 (O_1251,N_24875,N_24880);
and UO_1252 (O_1252,N_24285,N_24640);
or UO_1253 (O_1253,N_24734,N_24195);
xor UO_1254 (O_1254,N_24548,N_24670);
nand UO_1255 (O_1255,N_24919,N_24961);
and UO_1256 (O_1256,N_24483,N_24280);
or UO_1257 (O_1257,N_24147,N_24998);
or UO_1258 (O_1258,N_24279,N_24398);
or UO_1259 (O_1259,N_24939,N_24181);
and UO_1260 (O_1260,N_24084,N_24209);
and UO_1261 (O_1261,N_24354,N_24964);
and UO_1262 (O_1262,N_24375,N_24941);
nand UO_1263 (O_1263,N_24621,N_24727);
xor UO_1264 (O_1264,N_24250,N_24232);
nor UO_1265 (O_1265,N_24275,N_24532);
nor UO_1266 (O_1266,N_24496,N_24873);
and UO_1267 (O_1267,N_24743,N_24293);
and UO_1268 (O_1268,N_24096,N_24208);
nor UO_1269 (O_1269,N_24602,N_24475);
xnor UO_1270 (O_1270,N_24765,N_24367);
nand UO_1271 (O_1271,N_24831,N_24434);
xnor UO_1272 (O_1272,N_24751,N_24184);
and UO_1273 (O_1273,N_24859,N_24783);
nor UO_1274 (O_1274,N_24321,N_24897);
nand UO_1275 (O_1275,N_24263,N_24965);
xor UO_1276 (O_1276,N_24586,N_24922);
and UO_1277 (O_1277,N_24646,N_24548);
nand UO_1278 (O_1278,N_24823,N_24378);
xnor UO_1279 (O_1279,N_24261,N_24751);
or UO_1280 (O_1280,N_24790,N_24821);
or UO_1281 (O_1281,N_24402,N_24263);
nand UO_1282 (O_1282,N_24960,N_24422);
xor UO_1283 (O_1283,N_24735,N_24573);
nor UO_1284 (O_1284,N_24945,N_24272);
xnor UO_1285 (O_1285,N_24234,N_24354);
xor UO_1286 (O_1286,N_24386,N_24241);
or UO_1287 (O_1287,N_24124,N_24330);
or UO_1288 (O_1288,N_24532,N_24545);
nand UO_1289 (O_1289,N_24344,N_24696);
nor UO_1290 (O_1290,N_24098,N_24147);
and UO_1291 (O_1291,N_24926,N_24064);
or UO_1292 (O_1292,N_24951,N_24055);
xor UO_1293 (O_1293,N_24910,N_24138);
xnor UO_1294 (O_1294,N_24726,N_24491);
nand UO_1295 (O_1295,N_24182,N_24202);
xor UO_1296 (O_1296,N_24984,N_24990);
nor UO_1297 (O_1297,N_24047,N_24153);
nor UO_1298 (O_1298,N_24542,N_24194);
and UO_1299 (O_1299,N_24479,N_24860);
nor UO_1300 (O_1300,N_24586,N_24324);
xnor UO_1301 (O_1301,N_24649,N_24479);
and UO_1302 (O_1302,N_24708,N_24717);
xnor UO_1303 (O_1303,N_24992,N_24421);
nor UO_1304 (O_1304,N_24561,N_24113);
and UO_1305 (O_1305,N_24987,N_24620);
nor UO_1306 (O_1306,N_24339,N_24894);
or UO_1307 (O_1307,N_24244,N_24420);
xor UO_1308 (O_1308,N_24443,N_24524);
nand UO_1309 (O_1309,N_24254,N_24840);
or UO_1310 (O_1310,N_24498,N_24305);
and UO_1311 (O_1311,N_24810,N_24923);
and UO_1312 (O_1312,N_24441,N_24759);
nand UO_1313 (O_1313,N_24452,N_24129);
xor UO_1314 (O_1314,N_24678,N_24374);
nand UO_1315 (O_1315,N_24913,N_24779);
or UO_1316 (O_1316,N_24069,N_24828);
nand UO_1317 (O_1317,N_24978,N_24998);
xnor UO_1318 (O_1318,N_24033,N_24866);
and UO_1319 (O_1319,N_24905,N_24989);
or UO_1320 (O_1320,N_24026,N_24822);
nand UO_1321 (O_1321,N_24245,N_24174);
xor UO_1322 (O_1322,N_24200,N_24166);
nand UO_1323 (O_1323,N_24387,N_24802);
or UO_1324 (O_1324,N_24362,N_24702);
nand UO_1325 (O_1325,N_24713,N_24668);
xor UO_1326 (O_1326,N_24124,N_24967);
or UO_1327 (O_1327,N_24346,N_24256);
xor UO_1328 (O_1328,N_24530,N_24410);
nor UO_1329 (O_1329,N_24647,N_24654);
nand UO_1330 (O_1330,N_24366,N_24672);
nand UO_1331 (O_1331,N_24694,N_24587);
nor UO_1332 (O_1332,N_24835,N_24432);
xnor UO_1333 (O_1333,N_24884,N_24236);
or UO_1334 (O_1334,N_24859,N_24842);
nor UO_1335 (O_1335,N_24589,N_24680);
nand UO_1336 (O_1336,N_24632,N_24723);
or UO_1337 (O_1337,N_24602,N_24420);
nand UO_1338 (O_1338,N_24944,N_24578);
nand UO_1339 (O_1339,N_24672,N_24288);
nand UO_1340 (O_1340,N_24533,N_24435);
or UO_1341 (O_1341,N_24479,N_24478);
xnor UO_1342 (O_1342,N_24849,N_24977);
nor UO_1343 (O_1343,N_24354,N_24921);
or UO_1344 (O_1344,N_24495,N_24984);
or UO_1345 (O_1345,N_24891,N_24401);
nand UO_1346 (O_1346,N_24196,N_24446);
and UO_1347 (O_1347,N_24482,N_24612);
or UO_1348 (O_1348,N_24831,N_24535);
and UO_1349 (O_1349,N_24107,N_24625);
nand UO_1350 (O_1350,N_24330,N_24650);
or UO_1351 (O_1351,N_24205,N_24462);
and UO_1352 (O_1352,N_24465,N_24482);
nor UO_1353 (O_1353,N_24931,N_24675);
nor UO_1354 (O_1354,N_24459,N_24394);
and UO_1355 (O_1355,N_24871,N_24417);
nand UO_1356 (O_1356,N_24201,N_24750);
xor UO_1357 (O_1357,N_24854,N_24738);
or UO_1358 (O_1358,N_24115,N_24312);
and UO_1359 (O_1359,N_24605,N_24462);
nor UO_1360 (O_1360,N_24538,N_24147);
and UO_1361 (O_1361,N_24596,N_24084);
xor UO_1362 (O_1362,N_24624,N_24497);
xnor UO_1363 (O_1363,N_24386,N_24127);
xor UO_1364 (O_1364,N_24822,N_24581);
xor UO_1365 (O_1365,N_24622,N_24354);
xnor UO_1366 (O_1366,N_24268,N_24545);
and UO_1367 (O_1367,N_24756,N_24943);
or UO_1368 (O_1368,N_24140,N_24028);
or UO_1369 (O_1369,N_24931,N_24162);
xor UO_1370 (O_1370,N_24640,N_24664);
or UO_1371 (O_1371,N_24843,N_24803);
nand UO_1372 (O_1372,N_24316,N_24749);
nand UO_1373 (O_1373,N_24221,N_24983);
or UO_1374 (O_1374,N_24555,N_24820);
and UO_1375 (O_1375,N_24216,N_24991);
nor UO_1376 (O_1376,N_24502,N_24078);
and UO_1377 (O_1377,N_24218,N_24006);
and UO_1378 (O_1378,N_24626,N_24489);
or UO_1379 (O_1379,N_24373,N_24188);
or UO_1380 (O_1380,N_24520,N_24048);
nand UO_1381 (O_1381,N_24637,N_24495);
nor UO_1382 (O_1382,N_24493,N_24592);
xor UO_1383 (O_1383,N_24077,N_24533);
nand UO_1384 (O_1384,N_24930,N_24057);
and UO_1385 (O_1385,N_24020,N_24110);
nand UO_1386 (O_1386,N_24188,N_24490);
and UO_1387 (O_1387,N_24768,N_24243);
nand UO_1388 (O_1388,N_24527,N_24415);
and UO_1389 (O_1389,N_24562,N_24968);
nand UO_1390 (O_1390,N_24039,N_24725);
nor UO_1391 (O_1391,N_24851,N_24809);
xnor UO_1392 (O_1392,N_24316,N_24158);
nor UO_1393 (O_1393,N_24335,N_24087);
nand UO_1394 (O_1394,N_24906,N_24752);
or UO_1395 (O_1395,N_24839,N_24602);
nand UO_1396 (O_1396,N_24478,N_24661);
xor UO_1397 (O_1397,N_24374,N_24821);
nand UO_1398 (O_1398,N_24697,N_24920);
or UO_1399 (O_1399,N_24140,N_24532);
or UO_1400 (O_1400,N_24965,N_24101);
nor UO_1401 (O_1401,N_24692,N_24897);
xnor UO_1402 (O_1402,N_24607,N_24205);
nand UO_1403 (O_1403,N_24188,N_24315);
and UO_1404 (O_1404,N_24823,N_24949);
nand UO_1405 (O_1405,N_24189,N_24374);
nand UO_1406 (O_1406,N_24548,N_24838);
nor UO_1407 (O_1407,N_24329,N_24492);
nor UO_1408 (O_1408,N_24403,N_24791);
and UO_1409 (O_1409,N_24803,N_24481);
and UO_1410 (O_1410,N_24347,N_24265);
nor UO_1411 (O_1411,N_24783,N_24416);
xnor UO_1412 (O_1412,N_24005,N_24616);
nand UO_1413 (O_1413,N_24204,N_24382);
nand UO_1414 (O_1414,N_24507,N_24438);
or UO_1415 (O_1415,N_24832,N_24168);
or UO_1416 (O_1416,N_24109,N_24621);
nand UO_1417 (O_1417,N_24215,N_24030);
xnor UO_1418 (O_1418,N_24063,N_24860);
nor UO_1419 (O_1419,N_24078,N_24568);
and UO_1420 (O_1420,N_24228,N_24388);
and UO_1421 (O_1421,N_24378,N_24988);
nand UO_1422 (O_1422,N_24221,N_24231);
nor UO_1423 (O_1423,N_24342,N_24579);
xor UO_1424 (O_1424,N_24922,N_24177);
xnor UO_1425 (O_1425,N_24096,N_24461);
nor UO_1426 (O_1426,N_24918,N_24874);
or UO_1427 (O_1427,N_24519,N_24551);
nand UO_1428 (O_1428,N_24442,N_24988);
nand UO_1429 (O_1429,N_24984,N_24302);
xnor UO_1430 (O_1430,N_24770,N_24290);
xnor UO_1431 (O_1431,N_24775,N_24156);
nand UO_1432 (O_1432,N_24353,N_24145);
and UO_1433 (O_1433,N_24237,N_24071);
nor UO_1434 (O_1434,N_24759,N_24597);
or UO_1435 (O_1435,N_24249,N_24830);
nand UO_1436 (O_1436,N_24543,N_24050);
nor UO_1437 (O_1437,N_24824,N_24131);
nor UO_1438 (O_1438,N_24579,N_24850);
and UO_1439 (O_1439,N_24739,N_24149);
or UO_1440 (O_1440,N_24849,N_24640);
nor UO_1441 (O_1441,N_24321,N_24281);
or UO_1442 (O_1442,N_24646,N_24171);
and UO_1443 (O_1443,N_24645,N_24918);
or UO_1444 (O_1444,N_24662,N_24855);
and UO_1445 (O_1445,N_24977,N_24152);
xor UO_1446 (O_1446,N_24007,N_24800);
and UO_1447 (O_1447,N_24249,N_24742);
nor UO_1448 (O_1448,N_24377,N_24732);
and UO_1449 (O_1449,N_24120,N_24410);
and UO_1450 (O_1450,N_24604,N_24637);
nor UO_1451 (O_1451,N_24972,N_24873);
or UO_1452 (O_1452,N_24588,N_24513);
or UO_1453 (O_1453,N_24528,N_24406);
nor UO_1454 (O_1454,N_24816,N_24911);
nand UO_1455 (O_1455,N_24407,N_24831);
or UO_1456 (O_1456,N_24264,N_24322);
or UO_1457 (O_1457,N_24160,N_24090);
xnor UO_1458 (O_1458,N_24857,N_24059);
xor UO_1459 (O_1459,N_24309,N_24869);
and UO_1460 (O_1460,N_24451,N_24883);
or UO_1461 (O_1461,N_24721,N_24322);
xor UO_1462 (O_1462,N_24746,N_24647);
xnor UO_1463 (O_1463,N_24751,N_24538);
xnor UO_1464 (O_1464,N_24509,N_24182);
or UO_1465 (O_1465,N_24827,N_24921);
and UO_1466 (O_1466,N_24683,N_24898);
and UO_1467 (O_1467,N_24159,N_24357);
nand UO_1468 (O_1468,N_24848,N_24003);
nor UO_1469 (O_1469,N_24843,N_24155);
xnor UO_1470 (O_1470,N_24685,N_24802);
nor UO_1471 (O_1471,N_24393,N_24737);
xor UO_1472 (O_1472,N_24105,N_24281);
nor UO_1473 (O_1473,N_24983,N_24864);
and UO_1474 (O_1474,N_24315,N_24266);
and UO_1475 (O_1475,N_24587,N_24989);
nand UO_1476 (O_1476,N_24315,N_24947);
nand UO_1477 (O_1477,N_24729,N_24155);
and UO_1478 (O_1478,N_24569,N_24235);
or UO_1479 (O_1479,N_24538,N_24189);
and UO_1480 (O_1480,N_24981,N_24004);
xor UO_1481 (O_1481,N_24148,N_24831);
nand UO_1482 (O_1482,N_24346,N_24852);
or UO_1483 (O_1483,N_24896,N_24866);
nand UO_1484 (O_1484,N_24611,N_24099);
nor UO_1485 (O_1485,N_24926,N_24491);
xnor UO_1486 (O_1486,N_24895,N_24282);
xor UO_1487 (O_1487,N_24723,N_24131);
nor UO_1488 (O_1488,N_24385,N_24710);
nor UO_1489 (O_1489,N_24612,N_24554);
or UO_1490 (O_1490,N_24427,N_24326);
nand UO_1491 (O_1491,N_24673,N_24772);
xnor UO_1492 (O_1492,N_24036,N_24509);
and UO_1493 (O_1493,N_24249,N_24592);
xnor UO_1494 (O_1494,N_24498,N_24053);
nor UO_1495 (O_1495,N_24639,N_24882);
nor UO_1496 (O_1496,N_24982,N_24467);
nor UO_1497 (O_1497,N_24041,N_24574);
nand UO_1498 (O_1498,N_24044,N_24697);
xor UO_1499 (O_1499,N_24969,N_24675);
nor UO_1500 (O_1500,N_24617,N_24213);
or UO_1501 (O_1501,N_24798,N_24763);
nor UO_1502 (O_1502,N_24289,N_24838);
nand UO_1503 (O_1503,N_24938,N_24423);
and UO_1504 (O_1504,N_24174,N_24305);
nand UO_1505 (O_1505,N_24568,N_24721);
xor UO_1506 (O_1506,N_24399,N_24580);
and UO_1507 (O_1507,N_24860,N_24327);
nand UO_1508 (O_1508,N_24304,N_24337);
xor UO_1509 (O_1509,N_24705,N_24499);
and UO_1510 (O_1510,N_24559,N_24567);
nor UO_1511 (O_1511,N_24163,N_24807);
xnor UO_1512 (O_1512,N_24772,N_24918);
or UO_1513 (O_1513,N_24491,N_24732);
and UO_1514 (O_1514,N_24436,N_24958);
nor UO_1515 (O_1515,N_24709,N_24641);
nand UO_1516 (O_1516,N_24865,N_24013);
nor UO_1517 (O_1517,N_24140,N_24232);
xnor UO_1518 (O_1518,N_24372,N_24588);
xor UO_1519 (O_1519,N_24552,N_24991);
and UO_1520 (O_1520,N_24291,N_24866);
nor UO_1521 (O_1521,N_24135,N_24277);
xnor UO_1522 (O_1522,N_24153,N_24755);
nand UO_1523 (O_1523,N_24373,N_24722);
nand UO_1524 (O_1524,N_24436,N_24897);
and UO_1525 (O_1525,N_24168,N_24555);
and UO_1526 (O_1526,N_24293,N_24396);
xnor UO_1527 (O_1527,N_24562,N_24444);
nor UO_1528 (O_1528,N_24165,N_24794);
or UO_1529 (O_1529,N_24051,N_24605);
nor UO_1530 (O_1530,N_24296,N_24583);
and UO_1531 (O_1531,N_24746,N_24015);
xnor UO_1532 (O_1532,N_24747,N_24939);
or UO_1533 (O_1533,N_24553,N_24120);
or UO_1534 (O_1534,N_24673,N_24587);
nor UO_1535 (O_1535,N_24659,N_24615);
or UO_1536 (O_1536,N_24928,N_24040);
and UO_1537 (O_1537,N_24717,N_24279);
or UO_1538 (O_1538,N_24306,N_24979);
and UO_1539 (O_1539,N_24002,N_24375);
or UO_1540 (O_1540,N_24951,N_24670);
or UO_1541 (O_1541,N_24153,N_24021);
or UO_1542 (O_1542,N_24857,N_24042);
nor UO_1543 (O_1543,N_24049,N_24866);
and UO_1544 (O_1544,N_24001,N_24390);
xor UO_1545 (O_1545,N_24010,N_24020);
and UO_1546 (O_1546,N_24237,N_24162);
nor UO_1547 (O_1547,N_24059,N_24919);
and UO_1548 (O_1548,N_24620,N_24671);
nor UO_1549 (O_1549,N_24042,N_24943);
nand UO_1550 (O_1550,N_24312,N_24198);
or UO_1551 (O_1551,N_24781,N_24761);
nor UO_1552 (O_1552,N_24686,N_24329);
nor UO_1553 (O_1553,N_24866,N_24598);
xor UO_1554 (O_1554,N_24779,N_24172);
nor UO_1555 (O_1555,N_24713,N_24848);
nor UO_1556 (O_1556,N_24904,N_24035);
and UO_1557 (O_1557,N_24313,N_24583);
nand UO_1558 (O_1558,N_24475,N_24356);
and UO_1559 (O_1559,N_24088,N_24842);
and UO_1560 (O_1560,N_24146,N_24376);
nor UO_1561 (O_1561,N_24151,N_24084);
and UO_1562 (O_1562,N_24369,N_24187);
and UO_1563 (O_1563,N_24115,N_24862);
or UO_1564 (O_1564,N_24049,N_24689);
or UO_1565 (O_1565,N_24357,N_24854);
and UO_1566 (O_1566,N_24120,N_24836);
nor UO_1567 (O_1567,N_24395,N_24159);
nand UO_1568 (O_1568,N_24211,N_24133);
xnor UO_1569 (O_1569,N_24936,N_24680);
and UO_1570 (O_1570,N_24016,N_24513);
and UO_1571 (O_1571,N_24291,N_24393);
and UO_1572 (O_1572,N_24865,N_24841);
nor UO_1573 (O_1573,N_24927,N_24925);
or UO_1574 (O_1574,N_24152,N_24576);
or UO_1575 (O_1575,N_24134,N_24597);
or UO_1576 (O_1576,N_24853,N_24212);
nor UO_1577 (O_1577,N_24004,N_24144);
or UO_1578 (O_1578,N_24678,N_24610);
and UO_1579 (O_1579,N_24904,N_24986);
nor UO_1580 (O_1580,N_24014,N_24311);
nand UO_1581 (O_1581,N_24300,N_24274);
xnor UO_1582 (O_1582,N_24515,N_24812);
and UO_1583 (O_1583,N_24577,N_24350);
nand UO_1584 (O_1584,N_24877,N_24067);
and UO_1585 (O_1585,N_24460,N_24730);
and UO_1586 (O_1586,N_24555,N_24873);
nor UO_1587 (O_1587,N_24307,N_24627);
nand UO_1588 (O_1588,N_24411,N_24533);
nor UO_1589 (O_1589,N_24966,N_24827);
and UO_1590 (O_1590,N_24796,N_24337);
or UO_1591 (O_1591,N_24881,N_24676);
or UO_1592 (O_1592,N_24296,N_24630);
xor UO_1593 (O_1593,N_24019,N_24463);
xor UO_1594 (O_1594,N_24637,N_24857);
or UO_1595 (O_1595,N_24066,N_24536);
nor UO_1596 (O_1596,N_24822,N_24187);
xnor UO_1597 (O_1597,N_24772,N_24723);
and UO_1598 (O_1598,N_24686,N_24502);
or UO_1599 (O_1599,N_24034,N_24655);
and UO_1600 (O_1600,N_24951,N_24495);
nand UO_1601 (O_1601,N_24378,N_24357);
nand UO_1602 (O_1602,N_24298,N_24830);
and UO_1603 (O_1603,N_24200,N_24611);
xor UO_1604 (O_1604,N_24753,N_24736);
nor UO_1605 (O_1605,N_24300,N_24899);
or UO_1606 (O_1606,N_24072,N_24800);
xnor UO_1607 (O_1607,N_24667,N_24390);
and UO_1608 (O_1608,N_24347,N_24652);
and UO_1609 (O_1609,N_24653,N_24584);
nand UO_1610 (O_1610,N_24158,N_24861);
nor UO_1611 (O_1611,N_24275,N_24671);
xnor UO_1612 (O_1612,N_24809,N_24099);
or UO_1613 (O_1613,N_24421,N_24560);
or UO_1614 (O_1614,N_24334,N_24379);
nor UO_1615 (O_1615,N_24684,N_24617);
xor UO_1616 (O_1616,N_24545,N_24370);
nand UO_1617 (O_1617,N_24999,N_24110);
xor UO_1618 (O_1618,N_24857,N_24272);
xor UO_1619 (O_1619,N_24303,N_24907);
or UO_1620 (O_1620,N_24829,N_24021);
nor UO_1621 (O_1621,N_24966,N_24889);
and UO_1622 (O_1622,N_24169,N_24277);
and UO_1623 (O_1623,N_24033,N_24006);
nand UO_1624 (O_1624,N_24134,N_24160);
nand UO_1625 (O_1625,N_24118,N_24459);
and UO_1626 (O_1626,N_24025,N_24179);
or UO_1627 (O_1627,N_24595,N_24805);
nand UO_1628 (O_1628,N_24124,N_24401);
and UO_1629 (O_1629,N_24466,N_24824);
and UO_1630 (O_1630,N_24441,N_24693);
nand UO_1631 (O_1631,N_24060,N_24980);
xnor UO_1632 (O_1632,N_24563,N_24736);
nand UO_1633 (O_1633,N_24237,N_24963);
and UO_1634 (O_1634,N_24833,N_24608);
xor UO_1635 (O_1635,N_24086,N_24286);
nand UO_1636 (O_1636,N_24183,N_24964);
xor UO_1637 (O_1637,N_24876,N_24836);
xor UO_1638 (O_1638,N_24767,N_24043);
nand UO_1639 (O_1639,N_24712,N_24808);
nor UO_1640 (O_1640,N_24032,N_24260);
or UO_1641 (O_1641,N_24024,N_24370);
nor UO_1642 (O_1642,N_24527,N_24891);
nand UO_1643 (O_1643,N_24110,N_24374);
and UO_1644 (O_1644,N_24044,N_24880);
or UO_1645 (O_1645,N_24784,N_24630);
xor UO_1646 (O_1646,N_24046,N_24754);
nor UO_1647 (O_1647,N_24516,N_24002);
or UO_1648 (O_1648,N_24067,N_24183);
and UO_1649 (O_1649,N_24131,N_24731);
nor UO_1650 (O_1650,N_24355,N_24197);
xor UO_1651 (O_1651,N_24474,N_24942);
or UO_1652 (O_1652,N_24616,N_24264);
nor UO_1653 (O_1653,N_24634,N_24945);
nand UO_1654 (O_1654,N_24619,N_24011);
xnor UO_1655 (O_1655,N_24657,N_24960);
xnor UO_1656 (O_1656,N_24841,N_24555);
nand UO_1657 (O_1657,N_24481,N_24483);
or UO_1658 (O_1658,N_24057,N_24906);
and UO_1659 (O_1659,N_24591,N_24662);
xor UO_1660 (O_1660,N_24964,N_24825);
or UO_1661 (O_1661,N_24115,N_24145);
and UO_1662 (O_1662,N_24213,N_24105);
or UO_1663 (O_1663,N_24524,N_24153);
nand UO_1664 (O_1664,N_24460,N_24288);
xor UO_1665 (O_1665,N_24748,N_24841);
nand UO_1666 (O_1666,N_24692,N_24688);
xnor UO_1667 (O_1667,N_24503,N_24069);
or UO_1668 (O_1668,N_24585,N_24051);
or UO_1669 (O_1669,N_24580,N_24967);
or UO_1670 (O_1670,N_24535,N_24902);
and UO_1671 (O_1671,N_24924,N_24370);
nor UO_1672 (O_1672,N_24633,N_24378);
nor UO_1673 (O_1673,N_24249,N_24205);
and UO_1674 (O_1674,N_24177,N_24399);
or UO_1675 (O_1675,N_24417,N_24496);
nor UO_1676 (O_1676,N_24500,N_24958);
nor UO_1677 (O_1677,N_24001,N_24921);
nor UO_1678 (O_1678,N_24532,N_24930);
and UO_1679 (O_1679,N_24180,N_24688);
nand UO_1680 (O_1680,N_24542,N_24368);
nand UO_1681 (O_1681,N_24725,N_24936);
and UO_1682 (O_1682,N_24355,N_24037);
nand UO_1683 (O_1683,N_24150,N_24349);
xor UO_1684 (O_1684,N_24492,N_24687);
and UO_1685 (O_1685,N_24291,N_24801);
xor UO_1686 (O_1686,N_24773,N_24551);
nand UO_1687 (O_1687,N_24019,N_24961);
or UO_1688 (O_1688,N_24983,N_24822);
and UO_1689 (O_1689,N_24081,N_24129);
nor UO_1690 (O_1690,N_24340,N_24308);
and UO_1691 (O_1691,N_24966,N_24428);
or UO_1692 (O_1692,N_24704,N_24854);
and UO_1693 (O_1693,N_24668,N_24931);
and UO_1694 (O_1694,N_24334,N_24719);
and UO_1695 (O_1695,N_24951,N_24548);
nor UO_1696 (O_1696,N_24136,N_24684);
nand UO_1697 (O_1697,N_24477,N_24565);
or UO_1698 (O_1698,N_24759,N_24140);
and UO_1699 (O_1699,N_24990,N_24389);
or UO_1700 (O_1700,N_24390,N_24285);
or UO_1701 (O_1701,N_24784,N_24801);
and UO_1702 (O_1702,N_24738,N_24897);
nand UO_1703 (O_1703,N_24301,N_24718);
and UO_1704 (O_1704,N_24472,N_24916);
nand UO_1705 (O_1705,N_24136,N_24290);
nand UO_1706 (O_1706,N_24088,N_24540);
nand UO_1707 (O_1707,N_24131,N_24072);
nor UO_1708 (O_1708,N_24949,N_24416);
and UO_1709 (O_1709,N_24666,N_24082);
xnor UO_1710 (O_1710,N_24182,N_24686);
or UO_1711 (O_1711,N_24725,N_24168);
xnor UO_1712 (O_1712,N_24988,N_24876);
nand UO_1713 (O_1713,N_24484,N_24648);
and UO_1714 (O_1714,N_24005,N_24664);
or UO_1715 (O_1715,N_24629,N_24200);
or UO_1716 (O_1716,N_24257,N_24442);
or UO_1717 (O_1717,N_24838,N_24404);
xnor UO_1718 (O_1718,N_24755,N_24455);
nand UO_1719 (O_1719,N_24156,N_24822);
nor UO_1720 (O_1720,N_24772,N_24760);
nor UO_1721 (O_1721,N_24911,N_24805);
or UO_1722 (O_1722,N_24670,N_24141);
or UO_1723 (O_1723,N_24520,N_24076);
nor UO_1724 (O_1724,N_24567,N_24370);
nor UO_1725 (O_1725,N_24919,N_24023);
nor UO_1726 (O_1726,N_24756,N_24506);
nor UO_1727 (O_1727,N_24082,N_24120);
and UO_1728 (O_1728,N_24042,N_24117);
and UO_1729 (O_1729,N_24238,N_24560);
nand UO_1730 (O_1730,N_24252,N_24208);
xnor UO_1731 (O_1731,N_24631,N_24431);
xnor UO_1732 (O_1732,N_24970,N_24620);
xnor UO_1733 (O_1733,N_24750,N_24773);
xor UO_1734 (O_1734,N_24768,N_24769);
and UO_1735 (O_1735,N_24649,N_24458);
xor UO_1736 (O_1736,N_24934,N_24106);
nor UO_1737 (O_1737,N_24186,N_24104);
or UO_1738 (O_1738,N_24501,N_24894);
or UO_1739 (O_1739,N_24856,N_24303);
nor UO_1740 (O_1740,N_24164,N_24983);
xor UO_1741 (O_1741,N_24939,N_24951);
and UO_1742 (O_1742,N_24236,N_24776);
or UO_1743 (O_1743,N_24677,N_24623);
nand UO_1744 (O_1744,N_24886,N_24820);
or UO_1745 (O_1745,N_24332,N_24649);
xor UO_1746 (O_1746,N_24730,N_24781);
or UO_1747 (O_1747,N_24152,N_24858);
xnor UO_1748 (O_1748,N_24651,N_24470);
xor UO_1749 (O_1749,N_24509,N_24297);
nor UO_1750 (O_1750,N_24603,N_24541);
nand UO_1751 (O_1751,N_24698,N_24206);
nand UO_1752 (O_1752,N_24630,N_24080);
and UO_1753 (O_1753,N_24954,N_24682);
xor UO_1754 (O_1754,N_24451,N_24755);
nand UO_1755 (O_1755,N_24038,N_24665);
or UO_1756 (O_1756,N_24654,N_24131);
xor UO_1757 (O_1757,N_24332,N_24801);
xor UO_1758 (O_1758,N_24191,N_24508);
and UO_1759 (O_1759,N_24302,N_24107);
nor UO_1760 (O_1760,N_24921,N_24582);
nand UO_1761 (O_1761,N_24452,N_24918);
nor UO_1762 (O_1762,N_24557,N_24621);
nand UO_1763 (O_1763,N_24415,N_24061);
nand UO_1764 (O_1764,N_24978,N_24101);
and UO_1765 (O_1765,N_24141,N_24194);
nand UO_1766 (O_1766,N_24903,N_24642);
xor UO_1767 (O_1767,N_24765,N_24453);
nor UO_1768 (O_1768,N_24897,N_24776);
xor UO_1769 (O_1769,N_24692,N_24013);
or UO_1770 (O_1770,N_24707,N_24970);
xnor UO_1771 (O_1771,N_24911,N_24799);
nand UO_1772 (O_1772,N_24154,N_24402);
nand UO_1773 (O_1773,N_24697,N_24686);
xor UO_1774 (O_1774,N_24998,N_24634);
or UO_1775 (O_1775,N_24199,N_24105);
or UO_1776 (O_1776,N_24757,N_24279);
nand UO_1777 (O_1777,N_24118,N_24842);
nor UO_1778 (O_1778,N_24646,N_24386);
or UO_1779 (O_1779,N_24853,N_24558);
nor UO_1780 (O_1780,N_24967,N_24404);
or UO_1781 (O_1781,N_24721,N_24012);
and UO_1782 (O_1782,N_24877,N_24314);
and UO_1783 (O_1783,N_24364,N_24160);
xor UO_1784 (O_1784,N_24544,N_24409);
nand UO_1785 (O_1785,N_24440,N_24489);
nand UO_1786 (O_1786,N_24753,N_24497);
nand UO_1787 (O_1787,N_24560,N_24928);
or UO_1788 (O_1788,N_24084,N_24949);
nor UO_1789 (O_1789,N_24796,N_24027);
xnor UO_1790 (O_1790,N_24922,N_24534);
xor UO_1791 (O_1791,N_24360,N_24294);
and UO_1792 (O_1792,N_24016,N_24608);
and UO_1793 (O_1793,N_24736,N_24172);
or UO_1794 (O_1794,N_24020,N_24537);
xnor UO_1795 (O_1795,N_24325,N_24191);
xnor UO_1796 (O_1796,N_24010,N_24816);
or UO_1797 (O_1797,N_24444,N_24443);
or UO_1798 (O_1798,N_24214,N_24099);
nor UO_1799 (O_1799,N_24162,N_24397);
nand UO_1800 (O_1800,N_24531,N_24403);
or UO_1801 (O_1801,N_24513,N_24202);
xor UO_1802 (O_1802,N_24117,N_24322);
xnor UO_1803 (O_1803,N_24145,N_24304);
xor UO_1804 (O_1804,N_24982,N_24489);
xor UO_1805 (O_1805,N_24012,N_24671);
nor UO_1806 (O_1806,N_24448,N_24982);
xor UO_1807 (O_1807,N_24071,N_24972);
and UO_1808 (O_1808,N_24154,N_24990);
xnor UO_1809 (O_1809,N_24326,N_24413);
or UO_1810 (O_1810,N_24812,N_24008);
and UO_1811 (O_1811,N_24514,N_24970);
xor UO_1812 (O_1812,N_24368,N_24323);
nor UO_1813 (O_1813,N_24299,N_24118);
xor UO_1814 (O_1814,N_24483,N_24805);
nand UO_1815 (O_1815,N_24269,N_24356);
xnor UO_1816 (O_1816,N_24313,N_24528);
nor UO_1817 (O_1817,N_24340,N_24775);
or UO_1818 (O_1818,N_24629,N_24569);
nand UO_1819 (O_1819,N_24225,N_24606);
nand UO_1820 (O_1820,N_24335,N_24116);
or UO_1821 (O_1821,N_24169,N_24070);
xnor UO_1822 (O_1822,N_24783,N_24515);
nand UO_1823 (O_1823,N_24797,N_24724);
nand UO_1824 (O_1824,N_24612,N_24152);
xor UO_1825 (O_1825,N_24506,N_24875);
nor UO_1826 (O_1826,N_24578,N_24263);
or UO_1827 (O_1827,N_24178,N_24946);
and UO_1828 (O_1828,N_24862,N_24575);
and UO_1829 (O_1829,N_24281,N_24429);
nor UO_1830 (O_1830,N_24601,N_24157);
nor UO_1831 (O_1831,N_24568,N_24608);
xnor UO_1832 (O_1832,N_24535,N_24324);
and UO_1833 (O_1833,N_24792,N_24567);
nand UO_1834 (O_1834,N_24758,N_24689);
nand UO_1835 (O_1835,N_24800,N_24992);
xor UO_1836 (O_1836,N_24220,N_24501);
and UO_1837 (O_1837,N_24491,N_24350);
nor UO_1838 (O_1838,N_24789,N_24050);
and UO_1839 (O_1839,N_24990,N_24541);
and UO_1840 (O_1840,N_24875,N_24357);
or UO_1841 (O_1841,N_24084,N_24653);
and UO_1842 (O_1842,N_24776,N_24207);
and UO_1843 (O_1843,N_24112,N_24630);
or UO_1844 (O_1844,N_24676,N_24510);
xor UO_1845 (O_1845,N_24673,N_24522);
nand UO_1846 (O_1846,N_24502,N_24000);
nand UO_1847 (O_1847,N_24790,N_24470);
nor UO_1848 (O_1848,N_24017,N_24318);
and UO_1849 (O_1849,N_24665,N_24487);
nand UO_1850 (O_1850,N_24964,N_24159);
nand UO_1851 (O_1851,N_24125,N_24843);
or UO_1852 (O_1852,N_24025,N_24791);
xor UO_1853 (O_1853,N_24976,N_24404);
nand UO_1854 (O_1854,N_24231,N_24673);
and UO_1855 (O_1855,N_24568,N_24391);
nor UO_1856 (O_1856,N_24909,N_24393);
xnor UO_1857 (O_1857,N_24543,N_24845);
xnor UO_1858 (O_1858,N_24785,N_24335);
xor UO_1859 (O_1859,N_24455,N_24312);
nand UO_1860 (O_1860,N_24208,N_24162);
nand UO_1861 (O_1861,N_24829,N_24783);
nand UO_1862 (O_1862,N_24510,N_24316);
or UO_1863 (O_1863,N_24239,N_24132);
and UO_1864 (O_1864,N_24986,N_24176);
or UO_1865 (O_1865,N_24854,N_24886);
or UO_1866 (O_1866,N_24238,N_24659);
xnor UO_1867 (O_1867,N_24657,N_24671);
and UO_1868 (O_1868,N_24130,N_24515);
and UO_1869 (O_1869,N_24934,N_24913);
and UO_1870 (O_1870,N_24783,N_24249);
or UO_1871 (O_1871,N_24062,N_24400);
nand UO_1872 (O_1872,N_24006,N_24339);
or UO_1873 (O_1873,N_24883,N_24034);
xnor UO_1874 (O_1874,N_24470,N_24904);
nand UO_1875 (O_1875,N_24021,N_24820);
nand UO_1876 (O_1876,N_24236,N_24844);
or UO_1877 (O_1877,N_24631,N_24462);
xnor UO_1878 (O_1878,N_24092,N_24775);
xor UO_1879 (O_1879,N_24515,N_24456);
or UO_1880 (O_1880,N_24045,N_24921);
or UO_1881 (O_1881,N_24293,N_24171);
nand UO_1882 (O_1882,N_24834,N_24964);
and UO_1883 (O_1883,N_24736,N_24972);
nand UO_1884 (O_1884,N_24874,N_24473);
nor UO_1885 (O_1885,N_24989,N_24005);
and UO_1886 (O_1886,N_24510,N_24896);
and UO_1887 (O_1887,N_24549,N_24772);
nor UO_1888 (O_1888,N_24727,N_24800);
and UO_1889 (O_1889,N_24236,N_24407);
or UO_1890 (O_1890,N_24974,N_24255);
and UO_1891 (O_1891,N_24146,N_24497);
or UO_1892 (O_1892,N_24032,N_24402);
or UO_1893 (O_1893,N_24265,N_24963);
or UO_1894 (O_1894,N_24352,N_24319);
or UO_1895 (O_1895,N_24700,N_24287);
and UO_1896 (O_1896,N_24324,N_24476);
nor UO_1897 (O_1897,N_24080,N_24594);
nand UO_1898 (O_1898,N_24028,N_24647);
or UO_1899 (O_1899,N_24603,N_24542);
xnor UO_1900 (O_1900,N_24211,N_24815);
or UO_1901 (O_1901,N_24863,N_24868);
or UO_1902 (O_1902,N_24372,N_24218);
xnor UO_1903 (O_1903,N_24001,N_24928);
nand UO_1904 (O_1904,N_24569,N_24217);
xor UO_1905 (O_1905,N_24478,N_24743);
nand UO_1906 (O_1906,N_24424,N_24152);
nor UO_1907 (O_1907,N_24449,N_24155);
nand UO_1908 (O_1908,N_24576,N_24777);
and UO_1909 (O_1909,N_24874,N_24340);
xor UO_1910 (O_1910,N_24160,N_24203);
xor UO_1911 (O_1911,N_24631,N_24258);
xnor UO_1912 (O_1912,N_24228,N_24365);
nand UO_1913 (O_1913,N_24149,N_24718);
or UO_1914 (O_1914,N_24218,N_24191);
nor UO_1915 (O_1915,N_24446,N_24437);
nor UO_1916 (O_1916,N_24170,N_24399);
nor UO_1917 (O_1917,N_24794,N_24369);
nor UO_1918 (O_1918,N_24389,N_24619);
nand UO_1919 (O_1919,N_24400,N_24300);
or UO_1920 (O_1920,N_24704,N_24054);
and UO_1921 (O_1921,N_24462,N_24372);
or UO_1922 (O_1922,N_24662,N_24325);
nand UO_1923 (O_1923,N_24860,N_24722);
or UO_1924 (O_1924,N_24511,N_24648);
xor UO_1925 (O_1925,N_24831,N_24120);
nand UO_1926 (O_1926,N_24551,N_24941);
or UO_1927 (O_1927,N_24912,N_24624);
nand UO_1928 (O_1928,N_24757,N_24139);
nor UO_1929 (O_1929,N_24839,N_24728);
and UO_1930 (O_1930,N_24305,N_24750);
nand UO_1931 (O_1931,N_24513,N_24117);
nand UO_1932 (O_1932,N_24744,N_24028);
xor UO_1933 (O_1933,N_24628,N_24607);
xnor UO_1934 (O_1934,N_24053,N_24342);
xnor UO_1935 (O_1935,N_24052,N_24837);
or UO_1936 (O_1936,N_24056,N_24124);
nand UO_1937 (O_1937,N_24044,N_24517);
or UO_1938 (O_1938,N_24493,N_24202);
nor UO_1939 (O_1939,N_24235,N_24874);
nor UO_1940 (O_1940,N_24431,N_24119);
and UO_1941 (O_1941,N_24699,N_24688);
and UO_1942 (O_1942,N_24160,N_24861);
nand UO_1943 (O_1943,N_24058,N_24881);
and UO_1944 (O_1944,N_24996,N_24453);
or UO_1945 (O_1945,N_24889,N_24217);
nand UO_1946 (O_1946,N_24420,N_24662);
nor UO_1947 (O_1947,N_24700,N_24040);
nand UO_1948 (O_1948,N_24414,N_24452);
nand UO_1949 (O_1949,N_24020,N_24934);
nor UO_1950 (O_1950,N_24022,N_24107);
or UO_1951 (O_1951,N_24632,N_24888);
or UO_1952 (O_1952,N_24872,N_24087);
xor UO_1953 (O_1953,N_24590,N_24346);
nand UO_1954 (O_1954,N_24684,N_24462);
nor UO_1955 (O_1955,N_24926,N_24723);
xor UO_1956 (O_1956,N_24539,N_24560);
nor UO_1957 (O_1957,N_24410,N_24074);
nor UO_1958 (O_1958,N_24769,N_24023);
nand UO_1959 (O_1959,N_24733,N_24640);
nand UO_1960 (O_1960,N_24073,N_24101);
or UO_1961 (O_1961,N_24316,N_24707);
nand UO_1962 (O_1962,N_24679,N_24761);
nor UO_1963 (O_1963,N_24116,N_24540);
nand UO_1964 (O_1964,N_24455,N_24226);
and UO_1965 (O_1965,N_24226,N_24294);
or UO_1966 (O_1966,N_24477,N_24494);
or UO_1967 (O_1967,N_24852,N_24335);
xor UO_1968 (O_1968,N_24787,N_24368);
nand UO_1969 (O_1969,N_24884,N_24842);
and UO_1970 (O_1970,N_24844,N_24247);
nand UO_1971 (O_1971,N_24811,N_24905);
xor UO_1972 (O_1972,N_24455,N_24641);
and UO_1973 (O_1973,N_24073,N_24902);
nand UO_1974 (O_1974,N_24269,N_24494);
nor UO_1975 (O_1975,N_24259,N_24171);
or UO_1976 (O_1976,N_24964,N_24256);
and UO_1977 (O_1977,N_24944,N_24935);
nor UO_1978 (O_1978,N_24542,N_24521);
and UO_1979 (O_1979,N_24696,N_24684);
xnor UO_1980 (O_1980,N_24592,N_24059);
nand UO_1981 (O_1981,N_24834,N_24432);
nor UO_1982 (O_1982,N_24383,N_24506);
nor UO_1983 (O_1983,N_24876,N_24573);
or UO_1984 (O_1984,N_24989,N_24380);
nand UO_1985 (O_1985,N_24141,N_24263);
or UO_1986 (O_1986,N_24010,N_24110);
and UO_1987 (O_1987,N_24081,N_24971);
nand UO_1988 (O_1988,N_24673,N_24206);
nand UO_1989 (O_1989,N_24456,N_24882);
nand UO_1990 (O_1990,N_24655,N_24928);
and UO_1991 (O_1991,N_24049,N_24816);
or UO_1992 (O_1992,N_24751,N_24071);
and UO_1993 (O_1993,N_24737,N_24143);
xor UO_1994 (O_1994,N_24854,N_24320);
or UO_1995 (O_1995,N_24824,N_24523);
xor UO_1996 (O_1996,N_24101,N_24231);
xnor UO_1997 (O_1997,N_24964,N_24766);
nand UO_1998 (O_1998,N_24345,N_24072);
or UO_1999 (O_1999,N_24509,N_24172);
xnor UO_2000 (O_2000,N_24087,N_24070);
xor UO_2001 (O_2001,N_24439,N_24249);
nand UO_2002 (O_2002,N_24037,N_24542);
nand UO_2003 (O_2003,N_24878,N_24367);
and UO_2004 (O_2004,N_24694,N_24576);
and UO_2005 (O_2005,N_24138,N_24071);
nor UO_2006 (O_2006,N_24984,N_24077);
nor UO_2007 (O_2007,N_24060,N_24403);
or UO_2008 (O_2008,N_24032,N_24116);
nand UO_2009 (O_2009,N_24328,N_24715);
or UO_2010 (O_2010,N_24723,N_24482);
nor UO_2011 (O_2011,N_24178,N_24711);
xnor UO_2012 (O_2012,N_24270,N_24462);
nor UO_2013 (O_2013,N_24402,N_24059);
and UO_2014 (O_2014,N_24278,N_24403);
or UO_2015 (O_2015,N_24881,N_24334);
and UO_2016 (O_2016,N_24815,N_24742);
or UO_2017 (O_2017,N_24750,N_24006);
xor UO_2018 (O_2018,N_24943,N_24316);
nand UO_2019 (O_2019,N_24592,N_24580);
xor UO_2020 (O_2020,N_24132,N_24683);
or UO_2021 (O_2021,N_24923,N_24890);
or UO_2022 (O_2022,N_24272,N_24845);
xnor UO_2023 (O_2023,N_24030,N_24820);
xor UO_2024 (O_2024,N_24448,N_24102);
or UO_2025 (O_2025,N_24187,N_24572);
xnor UO_2026 (O_2026,N_24249,N_24920);
xor UO_2027 (O_2027,N_24056,N_24254);
nor UO_2028 (O_2028,N_24481,N_24451);
nand UO_2029 (O_2029,N_24732,N_24846);
and UO_2030 (O_2030,N_24929,N_24860);
nor UO_2031 (O_2031,N_24941,N_24028);
nand UO_2032 (O_2032,N_24014,N_24902);
and UO_2033 (O_2033,N_24737,N_24031);
nor UO_2034 (O_2034,N_24039,N_24025);
xnor UO_2035 (O_2035,N_24718,N_24998);
nand UO_2036 (O_2036,N_24777,N_24816);
nand UO_2037 (O_2037,N_24405,N_24851);
xor UO_2038 (O_2038,N_24332,N_24302);
or UO_2039 (O_2039,N_24708,N_24503);
nand UO_2040 (O_2040,N_24154,N_24552);
nor UO_2041 (O_2041,N_24106,N_24795);
xor UO_2042 (O_2042,N_24119,N_24650);
and UO_2043 (O_2043,N_24129,N_24828);
and UO_2044 (O_2044,N_24508,N_24439);
and UO_2045 (O_2045,N_24071,N_24025);
nor UO_2046 (O_2046,N_24924,N_24090);
xnor UO_2047 (O_2047,N_24801,N_24047);
xor UO_2048 (O_2048,N_24431,N_24163);
nand UO_2049 (O_2049,N_24726,N_24844);
and UO_2050 (O_2050,N_24810,N_24167);
xnor UO_2051 (O_2051,N_24057,N_24170);
xnor UO_2052 (O_2052,N_24723,N_24680);
nand UO_2053 (O_2053,N_24270,N_24550);
xnor UO_2054 (O_2054,N_24921,N_24409);
or UO_2055 (O_2055,N_24697,N_24197);
xnor UO_2056 (O_2056,N_24080,N_24165);
nand UO_2057 (O_2057,N_24011,N_24093);
nor UO_2058 (O_2058,N_24594,N_24666);
nor UO_2059 (O_2059,N_24846,N_24346);
nor UO_2060 (O_2060,N_24662,N_24875);
and UO_2061 (O_2061,N_24801,N_24778);
and UO_2062 (O_2062,N_24714,N_24254);
and UO_2063 (O_2063,N_24067,N_24970);
nand UO_2064 (O_2064,N_24279,N_24649);
nor UO_2065 (O_2065,N_24373,N_24652);
xnor UO_2066 (O_2066,N_24681,N_24216);
or UO_2067 (O_2067,N_24137,N_24085);
or UO_2068 (O_2068,N_24685,N_24125);
xor UO_2069 (O_2069,N_24644,N_24753);
xor UO_2070 (O_2070,N_24284,N_24909);
nor UO_2071 (O_2071,N_24158,N_24054);
nand UO_2072 (O_2072,N_24591,N_24849);
nor UO_2073 (O_2073,N_24098,N_24130);
or UO_2074 (O_2074,N_24843,N_24805);
nor UO_2075 (O_2075,N_24911,N_24085);
xnor UO_2076 (O_2076,N_24863,N_24272);
xor UO_2077 (O_2077,N_24761,N_24953);
xnor UO_2078 (O_2078,N_24018,N_24466);
nand UO_2079 (O_2079,N_24039,N_24377);
or UO_2080 (O_2080,N_24358,N_24723);
xor UO_2081 (O_2081,N_24764,N_24518);
or UO_2082 (O_2082,N_24001,N_24565);
xor UO_2083 (O_2083,N_24407,N_24507);
and UO_2084 (O_2084,N_24757,N_24123);
xor UO_2085 (O_2085,N_24339,N_24245);
and UO_2086 (O_2086,N_24396,N_24804);
xor UO_2087 (O_2087,N_24259,N_24146);
nand UO_2088 (O_2088,N_24552,N_24799);
nor UO_2089 (O_2089,N_24752,N_24838);
nor UO_2090 (O_2090,N_24014,N_24042);
nand UO_2091 (O_2091,N_24026,N_24537);
and UO_2092 (O_2092,N_24615,N_24421);
xor UO_2093 (O_2093,N_24251,N_24525);
and UO_2094 (O_2094,N_24929,N_24525);
xnor UO_2095 (O_2095,N_24844,N_24435);
nor UO_2096 (O_2096,N_24823,N_24951);
and UO_2097 (O_2097,N_24589,N_24874);
xor UO_2098 (O_2098,N_24764,N_24976);
nor UO_2099 (O_2099,N_24476,N_24717);
xor UO_2100 (O_2100,N_24028,N_24506);
and UO_2101 (O_2101,N_24456,N_24092);
nand UO_2102 (O_2102,N_24155,N_24578);
xor UO_2103 (O_2103,N_24532,N_24295);
and UO_2104 (O_2104,N_24759,N_24267);
xor UO_2105 (O_2105,N_24511,N_24058);
nand UO_2106 (O_2106,N_24320,N_24985);
and UO_2107 (O_2107,N_24033,N_24273);
or UO_2108 (O_2108,N_24243,N_24353);
xnor UO_2109 (O_2109,N_24778,N_24314);
and UO_2110 (O_2110,N_24322,N_24061);
nor UO_2111 (O_2111,N_24872,N_24665);
or UO_2112 (O_2112,N_24648,N_24851);
xnor UO_2113 (O_2113,N_24018,N_24822);
xnor UO_2114 (O_2114,N_24049,N_24926);
nand UO_2115 (O_2115,N_24043,N_24073);
and UO_2116 (O_2116,N_24703,N_24179);
and UO_2117 (O_2117,N_24116,N_24542);
xor UO_2118 (O_2118,N_24868,N_24962);
and UO_2119 (O_2119,N_24768,N_24336);
xnor UO_2120 (O_2120,N_24859,N_24350);
xnor UO_2121 (O_2121,N_24333,N_24080);
or UO_2122 (O_2122,N_24960,N_24957);
nand UO_2123 (O_2123,N_24864,N_24498);
nand UO_2124 (O_2124,N_24104,N_24099);
and UO_2125 (O_2125,N_24769,N_24035);
nor UO_2126 (O_2126,N_24862,N_24520);
and UO_2127 (O_2127,N_24743,N_24790);
and UO_2128 (O_2128,N_24722,N_24780);
nor UO_2129 (O_2129,N_24399,N_24920);
and UO_2130 (O_2130,N_24962,N_24919);
nor UO_2131 (O_2131,N_24362,N_24006);
or UO_2132 (O_2132,N_24217,N_24634);
nand UO_2133 (O_2133,N_24638,N_24115);
and UO_2134 (O_2134,N_24157,N_24464);
xnor UO_2135 (O_2135,N_24034,N_24133);
xnor UO_2136 (O_2136,N_24111,N_24718);
nand UO_2137 (O_2137,N_24199,N_24261);
nand UO_2138 (O_2138,N_24437,N_24398);
nor UO_2139 (O_2139,N_24869,N_24509);
or UO_2140 (O_2140,N_24582,N_24931);
xnor UO_2141 (O_2141,N_24279,N_24458);
nor UO_2142 (O_2142,N_24340,N_24636);
nand UO_2143 (O_2143,N_24821,N_24244);
nor UO_2144 (O_2144,N_24778,N_24205);
or UO_2145 (O_2145,N_24028,N_24248);
or UO_2146 (O_2146,N_24705,N_24253);
or UO_2147 (O_2147,N_24236,N_24508);
nand UO_2148 (O_2148,N_24164,N_24694);
or UO_2149 (O_2149,N_24955,N_24267);
and UO_2150 (O_2150,N_24596,N_24207);
and UO_2151 (O_2151,N_24198,N_24509);
or UO_2152 (O_2152,N_24531,N_24613);
nand UO_2153 (O_2153,N_24534,N_24277);
xor UO_2154 (O_2154,N_24177,N_24538);
nor UO_2155 (O_2155,N_24183,N_24849);
nor UO_2156 (O_2156,N_24835,N_24021);
xor UO_2157 (O_2157,N_24206,N_24495);
or UO_2158 (O_2158,N_24975,N_24566);
and UO_2159 (O_2159,N_24221,N_24329);
xnor UO_2160 (O_2160,N_24580,N_24261);
xnor UO_2161 (O_2161,N_24128,N_24853);
xor UO_2162 (O_2162,N_24801,N_24708);
xnor UO_2163 (O_2163,N_24206,N_24888);
nand UO_2164 (O_2164,N_24256,N_24903);
or UO_2165 (O_2165,N_24559,N_24611);
or UO_2166 (O_2166,N_24829,N_24026);
and UO_2167 (O_2167,N_24984,N_24279);
or UO_2168 (O_2168,N_24887,N_24831);
or UO_2169 (O_2169,N_24223,N_24000);
and UO_2170 (O_2170,N_24295,N_24526);
nor UO_2171 (O_2171,N_24556,N_24632);
and UO_2172 (O_2172,N_24383,N_24009);
and UO_2173 (O_2173,N_24836,N_24662);
nor UO_2174 (O_2174,N_24723,N_24992);
nand UO_2175 (O_2175,N_24493,N_24864);
and UO_2176 (O_2176,N_24094,N_24493);
or UO_2177 (O_2177,N_24208,N_24324);
or UO_2178 (O_2178,N_24334,N_24179);
and UO_2179 (O_2179,N_24106,N_24097);
xor UO_2180 (O_2180,N_24062,N_24477);
nor UO_2181 (O_2181,N_24410,N_24857);
nor UO_2182 (O_2182,N_24415,N_24977);
nand UO_2183 (O_2183,N_24128,N_24735);
nand UO_2184 (O_2184,N_24395,N_24829);
xor UO_2185 (O_2185,N_24754,N_24633);
or UO_2186 (O_2186,N_24569,N_24348);
or UO_2187 (O_2187,N_24800,N_24482);
or UO_2188 (O_2188,N_24969,N_24080);
xor UO_2189 (O_2189,N_24052,N_24292);
and UO_2190 (O_2190,N_24367,N_24572);
xnor UO_2191 (O_2191,N_24000,N_24771);
nand UO_2192 (O_2192,N_24440,N_24218);
nand UO_2193 (O_2193,N_24882,N_24737);
xor UO_2194 (O_2194,N_24377,N_24843);
nor UO_2195 (O_2195,N_24246,N_24169);
and UO_2196 (O_2196,N_24617,N_24826);
and UO_2197 (O_2197,N_24212,N_24216);
and UO_2198 (O_2198,N_24773,N_24731);
nor UO_2199 (O_2199,N_24696,N_24873);
and UO_2200 (O_2200,N_24645,N_24535);
or UO_2201 (O_2201,N_24887,N_24323);
or UO_2202 (O_2202,N_24225,N_24326);
or UO_2203 (O_2203,N_24207,N_24116);
or UO_2204 (O_2204,N_24159,N_24714);
xnor UO_2205 (O_2205,N_24936,N_24783);
xor UO_2206 (O_2206,N_24970,N_24399);
nor UO_2207 (O_2207,N_24264,N_24853);
nand UO_2208 (O_2208,N_24006,N_24409);
nor UO_2209 (O_2209,N_24157,N_24749);
or UO_2210 (O_2210,N_24493,N_24174);
and UO_2211 (O_2211,N_24161,N_24473);
nand UO_2212 (O_2212,N_24655,N_24205);
nor UO_2213 (O_2213,N_24068,N_24074);
and UO_2214 (O_2214,N_24881,N_24900);
and UO_2215 (O_2215,N_24783,N_24007);
and UO_2216 (O_2216,N_24758,N_24544);
and UO_2217 (O_2217,N_24184,N_24412);
xor UO_2218 (O_2218,N_24742,N_24927);
or UO_2219 (O_2219,N_24513,N_24652);
nand UO_2220 (O_2220,N_24612,N_24880);
xor UO_2221 (O_2221,N_24848,N_24504);
and UO_2222 (O_2222,N_24833,N_24788);
nand UO_2223 (O_2223,N_24327,N_24386);
nand UO_2224 (O_2224,N_24326,N_24101);
and UO_2225 (O_2225,N_24235,N_24288);
or UO_2226 (O_2226,N_24689,N_24561);
or UO_2227 (O_2227,N_24375,N_24213);
or UO_2228 (O_2228,N_24674,N_24221);
nand UO_2229 (O_2229,N_24790,N_24596);
or UO_2230 (O_2230,N_24367,N_24578);
xor UO_2231 (O_2231,N_24099,N_24517);
and UO_2232 (O_2232,N_24414,N_24442);
or UO_2233 (O_2233,N_24837,N_24284);
or UO_2234 (O_2234,N_24954,N_24434);
or UO_2235 (O_2235,N_24839,N_24466);
nand UO_2236 (O_2236,N_24802,N_24129);
nand UO_2237 (O_2237,N_24294,N_24580);
xor UO_2238 (O_2238,N_24037,N_24563);
and UO_2239 (O_2239,N_24290,N_24633);
nand UO_2240 (O_2240,N_24465,N_24612);
and UO_2241 (O_2241,N_24211,N_24803);
nand UO_2242 (O_2242,N_24303,N_24643);
and UO_2243 (O_2243,N_24124,N_24413);
or UO_2244 (O_2244,N_24897,N_24853);
xor UO_2245 (O_2245,N_24450,N_24715);
nor UO_2246 (O_2246,N_24142,N_24361);
or UO_2247 (O_2247,N_24193,N_24209);
nand UO_2248 (O_2248,N_24942,N_24994);
and UO_2249 (O_2249,N_24286,N_24015);
or UO_2250 (O_2250,N_24405,N_24610);
nand UO_2251 (O_2251,N_24747,N_24087);
and UO_2252 (O_2252,N_24795,N_24066);
or UO_2253 (O_2253,N_24104,N_24492);
or UO_2254 (O_2254,N_24314,N_24218);
nand UO_2255 (O_2255,N_24853,N_24644);
nand UO_2256 (O_2256,N_24251,N_24465);
and UO_2257 (O_2257,N_24134,N_24853);
xor UO_2258 (O_2258,N_24107,N_24475);
xor UO_2259 (O_2259,N_24060,N_24482);
nor UO_2260 (O_2260,N_24792,N_24041);
or UO_2261 (O_2261,N_24873,N_24852);
nand UO_2262 (O_2262,N_24150,N_24715);
and UO_2263 (O_2263,N_24111,N_24339);
xor UO_2264 (O_2264,N_24694,N_24392);
nand UO_2265 (O_2265,N_24946,N_24430);
xor UO_2266 (O_2266,N_24071,N_24390);
and UO_2267 (O_2267,N_24842,N_24887);
nand UO_2268 (O_2268,N_24509,N_24124);
xnor UO_2269 (O_2269,N_24834,N_24263);
or UO_2270 (O_2270,N_24334,N_24852);
nand UO_2271 (O_2271,N_24074,N_24260);
nand UO_2272 (O_2272,N_24565,N_24289);
or UO_2273 (O_2273,N_24089,N_24841);
nand UO_2274 (O_2274,N_24611,N_24865);
nand UO_2275 (O_2275,N_24703,N_24393);
nor UO_2276 (O_2276,N_24614,N_24464);
xor UO_2277 (O_2277,N_24369,N_24008);
and UO_2278 (O_2278,N_24054,N_24920);
xor UO_2279 (O_2279,N_24948,N_24143);
nand UO_2280 (O_2280,N_24734,N_24923);
nor UO_2281 (O_2281,N_24795,N_24056);
nand UO_2282 (O_2282,N_24074,N_24245);
or UO_2283 (O_2283,N_24026,N_24448);
nor UO_2284 (O_2284,N_24439,N_24412);
xnor UO_2285 (O_2285,N_24561,N_24160);
nand UO_2286 (O_2286,N_24933,N_24182);
xnor UO_2287 (O_2287,N_24091,N_24658);
nor UO_2288 (O_2288,N_24665,N_24769);
xnor UO_2289 (O_2289,N_24364,N_24561);
or UO_2290 (O_2290,N_24644,N_24524);
nand UO_2291 (O_2291,N_24113,N_24323);
and UO_2292 (O_2292,N_24457,N_24795);
xor UO_2293 (O_2293,N_24856,N_24185);
xor UO_2294 (O_2294,N_24041,N_24350);
xor UO_2295 (O_2295,N_24979,N_24272);
nand UO_2296 (O_2296,N_24331,N_24513);
or UO_2297 (O_2297,N_24088,N_24064);
nand UO_2298 (O_2298,N_24734,N_24086);
and UO_2299 (O_2299,N_24639,N_24349);
nor UO_2300 (O_2300,N_24406,N_24069);
and UO_2301 (O_2301,N_24858,N_24300);
or UO_2302 (O_2302,N_24118,N_24881);
nor UO_2303 (O_2303,N_24300,N_24176);
and UO_2304 (O_2304,N_24007,N_24753);
or UO_2305 (O_2305,N_24401,N_24271);
and UO_2306 (O_2306,N_24654,N_24454);
nand UO_2307 (O_2307,N_24331,N_24107);
or UO_2308 (O_2308,N_24731,N_24931);
and UO_2309 (O_2309,N_24530,N_24971);
and UO_2310 (O_2310,N_24056,N_24592);
or UO_2311 (O_2311,N_24169,N_24166);
nand UO_2312 (O_2312,N_24261,N_24353);
nand UO_2313 (O_2313,N_24431,N_24495);
xor UO_2314 (O_2314,N_24048,N_24104);
and UO_2315 (O_2315,N_24288,N_24777);
nand UO_2316 (O_2316,N_24881,N_24574);
nor UO_2317 (O_2317,N_24775,N_24977);
nor UO_2318 (O_2318,N_24112,N_24979);
nor UO_2319 (O_2319,N_24137,N_24243);
nand UO_2320 (O_2320,N_24392,N_24561);
xor UO_2321 (O_2321,N_24056,N_24650);
and UO_2322 (O_2322,N_24470,N_24971);
or UO_2323 (O_2323,N_24840,N_24244);
nand UO_2324 (O_2324,N_24932,N_24764);
nand UO_2325 (O_2325,N_24175,N_24231);
or UO_2326 (O_2326,N_24090,N_24243);
and UO_2327 (O_2327,N_24217,N_24034);
and UO_2328 (O_2328,N_24297,N_24470);
nor UO_2329 (O_2329,N_24984,N_24943);
nand UO_2330 (O_2330,N_24164,N_24560);
nor UO_2331 (O_2331,N_24420,N_24402);
nor UO_2332 (O_2332,N_24823,N_24409);
nand UO_2333 (O_2333,N_24770,N_24240);
nor UO_2334 (O_2334,N_24171,N_24501);
and UO_2335 (O_2335,N_24318,N_24119);
and UO_2336 (O_2336,N_24051,N_24457);
xnor UO_2337 (O_2337,N_24646,N_24423);
nor UO_2338 (O_2338,N_24970,N_24537);
xor UO_2339 (O_2339,N_24633,N_24550);
xnor UO_2340 (O_2340,N_24337,N_24067);
xnor UO_2341 (O_2341,N_24944,N_24634);
or UO_2342 (O_2342,N_24702,N_24426);
or UO_2343 (O_2343,N_24781,N_24516);
nand UO_2344 (O_2344,N_24366,N_24792);
or UO_2345 (O_2345,N_24220,N_24172);
xnor UO_2346 (O_2346,N_24122,N_24478);
and UO_2347 (O_2347,N_24832,N_24767);
or UO_2348 (O_2348,N_24671,N_24690);
xnor UO_2349 (O_2349,N_24007,N_24341);
or UO_2350 (O_2350,N_24723,N_24631);
xnor UO_2351 (O_2351,N_24399,N_24708);
xor UO_2352 (O_2352,N_24813,N_24646);
nand UO_2353 (O_2353,N_24560,N_24618);
and UO_2354 (O_2354,N_24125,N_24630);
xnor UO_2355 (O_2355,N_24693,N_24389);
xor UO_2356 (O_2356,N_24991,N_24692);
and UO_2357 (O_2357,N_24658,N_24510);
xnor UO_2358 (O_2358,N_24331,N_24065);
or UO_2359 (O_2359,N_24404,N_24875);
or UO_2360 (O_2360,N_24693,N_24881);
xnor UO_2361 (O_2361,N_24443,N_24700);
and UO_2362 (O_2362,N_24588,N_24219);
xnor UO_2363 (O_2363,N_24490,N_24540);
or UO_2364 (O_2364,N_24299,N_24687);
or UO_2365 (O_2365,N_24666,N_24643);
and UO_2366 (O_2366,N_24178,N_24797);
nor UO_2367 (O_2367,N_24125,N_24475);
xnor UO_2368 (O_2368,N_24804,N_24125);
nand UO_2369 (O_2369,N_24643,N_24737);
nor UO_2370 (O_2370,N_24975,N_24704);
nor UO_2371 (O_2371,N_24549,N_24670);
or UO_2372 (O_2372,N_24891,N_24634);
nand UO_2373 (O_2373,N_24219,N_24566);
or UO_2374 (O_2374,N_24752,N_24954);
xor UO_2375 (O_2375,N_24388,N_24317);
nor UO_2376 (O_2376,N_24734,N_24752);
and UO_2377 (O_2377,N_24747,N_24311);
or UO_2378 (O_2378,N_24796,N_24813);
nand UO_2379 (O_2379,N_24211,N_24973);
or UO_2380 (O_2380,N_24978,N_24216);
xor UO_2381 (O_2381,N_24175,N_24122);
or UO_2382 (O_2382,N_24659,N_24807);
nand UO_2383 (O_2383,N_24990,N_24777);
xnor UO_2384 (O_2384,N_24100,N_24281);
nor UO_2385 (O_2385,N_24755,N_24270);
nand UO_2386 (O_2386,N_24403,N_24553);
xnor UO_2387 (O_2387,N_24430,N_24831);
xor UO_2388 (O_2388,N_24073,N_24363);
and UO_2389 (O_2389,N_24437,N_24591);
xnor UO_2390 (O_2390,N_24588,N_24117);
nor UO_2391 (O_2391,N_24814,N_24944);
nand UO_2392 (O_2392,N_24736,N_24370);
nand UO_2393 (O_2393,N_24566,N_24138);
nor UO_2394 (O_2394,N_24531,N_24773);
nand UO_2395 (O_2395,N_24028,N_24547);
xor UO_2396 (O_2396,N_24095,N_24324);
xor UO_2397 (O_2397,N_24710,N_24501);
and UO_2398 (O_2398,N_24516,N_24363);
xor UO_2399 (O_2399,N_24371,N_24215);
and UO_2400 (O_2400,N_24850,N_24947);
xnor UO_2401 (O_2401,N_24089,N_24368);
or UO_2402 (O_2402,N_24607,N_24523);
nand UO_2403 (O_2403,N_24644,N_24078);
xor UO_2404 (O_2404,N_24049,N_24265);
or UO_2405 (O_2405,N_24340,N_24113);
xor UO_2406 (O_2406,N_24183,N_24797);
xor UO_2407 (O_2407,N_24129,N_24518);
or UO_2408 (O_2408,N_24223,N_24841);
xnor UO_2409 (O_2409,N_24512,N_24642);
or UO_2410 (O_2410,N_24515,N_24479);
nand UO_2411 (O_2411,N_24443,N_24111);
nand UO_2412 (O_2412,N_24265,N_24291);
nor UO_2413 (O_2413,N_24916,N_24841);
nor UO_2414 (O_2414,N_24843,N_24916);
and UO_2415 (O_2415,N_24798,N_24307);
and UO_2416 (O_2416,N_24354,N_24092);
and UO_2417 (O_2417,N_24966,N_24474);
and UO_2418 (O_2418,N_24290,N_24486);
nand UO_2419 (O_2419,N_24588,N_24166);
nand UO_2420 (O_2420,N_24951,N_24125);
and UO_2421 (O_2421,N_24594,N_24826);
nor UO_2422 (O_2422,N_24141,N_24261);
nor UO_2423 (O_2423,N_24245,N_24051);
nand UO_2424 (O_2424,N_24776,N_24330);
xor UO_2425 (O_2425,N_24326,N_24652);
nor UO_2426 (O_2426,N_24161,N_24468);
and UO_2427 (O_2427,N_24635,N_24893);
and UO_2428 (O_2428,N_24565,N_24311);
and UO_2429 (O_2429,N_24634,N_24117);
or UO_2430 (O_2430,N_24339,N_24390);
xnor UO_2431 (O_2431,N_24598,N_24347);
and UO_2432 (O_2432,N_24816,N_24370);
xor UO_2433 (O_2433,N_24662,N_24630);
and UO_2434 (O_2434,N_24081,N_24018);
and UO_2435 (O_2435,N_24268,N_24076);
and UO_2436 (O_2436,N_24527,N_24607);
nand UO_2437 (O_2437,N_24036,N_24842);
or UO_2438 (O_2438,N_24586,N_24222);
nand UO_2439 (O_2439,N_24226,N_24727);
nand UO_2440 (O_2440,N_24322,N_24686);
nor UO_2441 (O_2441,N_24291,N_24120);
nor UO_2442 (O_2442,N_24780,N_24591);
and UO_2443 (O_2443,N_24246,N_24365);
xnor UO_2444 (O_2444,N_24375,N_24457);
xor UO_2445 (O_2445,N_24612,N_24561);
or UO_2446 (O_2446,N_24240,N_24114);
nand UO_2447 (O_2447,N_24061,N_24576);
nand UO_2448 (O_2448,N_24782,N_24239);
and UO_2449 (O_2449,N_24683,N_24043);
and UO_2450 (O_2450,N_24474,N_24718);
and UO_2451 (O_2451,N_24595,N_24949);
nand UO_2452 (O_2452,N_24367,N_24525);
or UO_2453 (O_2453,N_24254,N_24385);
nor UO_2454 (O_2454,N_24941,N_24657);
xor UO_2455 (O_2455,N_24440,N_24583);
nor UO_2456 (O_2456,N_24919,N_24601);
or UO_2457 (O_2457,N_24521,N_24716);
and UO_2458 (O_2458,N_24793,N_24985);
nor UO_2459 (O_2459,N_24322,N_24477);
or UO_2460 (O_2460,N_24982,N_24052);
or UO_2461 (O_2461,N_24238,N_24140);
or UO_2462 (O_2462,N_24704,N_24105);
or UO_2463 (O_2463,N_24112,N_24366);
xor UO_2464 (O_2464,N_24933,N_24358);
nor UO_2465 (O_2465,N_24289,N_24493);
nand UO_2466 (O_2466,N_24551,N_24758);
xor UO_2467 (O_2467,N_24276,N_24616);
or UO_2468 (O_2468,N_24259,N_24779);
xor UO_2469 (O_2469,N_24518,N_24781);
xor UO_2470 (O_2470,N_24504,N_24817);
xor UO_2471 (O_2471,N_24577,N_24380);
or UO_2472 (O_2472,N_24695,N_24786);
nand UO_2473 (O_2473,N_24970,N_24335);
and UO_2474 (O_2474,N_24262,N_24682);
and UO_2475 (O_2475,N_24983,N_24168);
nor UO_2476 (O_2476,N_24369,N_24958);
xnor UO_2477 (O_2477,N_24208,N_24868);
or UO_2478 (O_2478,N_24778,N_24246);
nand UO_2479 (O_2479,N_24526,N_24335);
nand UO_2480 (O_2480,N_24684,N_24765);
nand UO_2481 (O_2481,N_24573,N_24349);
or UO_2482 (O_2482,N_24627,N_24068);
xor UO_2483 (O_2483,N_24186,N_24601);
nor UO_2484 (O_2484,N_24825,N_24154);
nor UO_2485 (O_2485,N_24127,N_24556);
nand UO_2486 (O_2486,N_24912,N_24787);
nand UO_2487 (O_2487,N_24019,N_24695);
or UO_2488 (O_2488,N_24333,N_24923);
or UO_2489 (O_2489,N_24231,N_24834);
xnor UO_2490 (O_2490,N_24425,N_24103);
or UO_2491 (O_2491,N_24422,N_24164);
and UO_2492 (O_2492,N_24457,N_24750);
xor UO_2493 (O_2493,N_24481,N_24938);
nor UO_2494 (O_2494,N_24387,N_24384);
or UO_2495 (O_2495,N_24954,N_24808);
and UO_2496 (O_2496,N_24302,N_24403);
or UO_2497 (O_2497,N_24977,N_24195);
nand UO_2498 (O_2498,N_24211,N_24391);
nor UO_2499 (O_2499,N_24020,N_24478);
nand UO_2500 (O_2500,N_24760,N_24577);
and UO_2501 (O_2501,N_24096,N_24099);
or UO_2502 (O_2502,N_24928,N_24934);
and UO_2503 (O_2503,N_24814,N_24986);
nor UO_2504 (O_2504,N_24889,N_24308);
nand UO_2505 (O_2505,N_24720,N_24179);
or UO_2506 (O_2506,N_24710,N_24778);
nand UO_2507 (O_2507,N_24642,N_24493);
nand UO_2508 (O_2508,N_24644,N_24866);
nand UO_2509 (O_2509,N_24540,N_24234);
nand UO_2510 (O_2510,N_24809,N_24993);
and UO_2511 (O_2511,N_24349,N_24649);
or UO_2512 (O_2512,N_24907,N_24417);
or UO_2513 (O_2513,N_24363,N_24618);
xnor UO_2514 (O_2514,N_24839,N_24597);
and UO_2515 (O_2515,N_24182,N_24108);
or UO_2516 (O_2516,N_24324,N_24649);
nor UO_2517 (O_2517,N_24429,N_24325);
or UO_2518 (O_2518,N_24710,N_24927);
and UO_2519 (O_2519,N_24407,N_24479);
nand UO_2520 (O_2520,N_24791,N_24341);
or UO_2521 (O_2521,N_24416,N_24059);
and UO_2522 (O_2522,N_24323,N_24513);
and UO_2523 (O_2523,N_24218,N_24937);
nand UO_2524 (O_2524,N_24225,N_24164);
xor UO_2525 (O_2525,N_24994,N_24473);
nor UO_2526 (O_2526,N_24603,N_24520);
xnor UO_2527 (O_2527,N_24452,N_24517);
or UO_2528 (O_2528,N_24876,N_24992);
xor UO_2529 (O_2529,N_24099,N_24628);
nand UO_2530 (O_2530,N_24505,N_24693);
or UO_2531 (O_2531,N_24770,N_24291);
or UO_2532 (O_2532,N_24064,N_24458);
xor UO_2533 (O_2533,N_24490,N_24890);
nand UO_2534 (O_2534,N_24028,N_24238);
or UO_2535 (O_2535,N_24694,N_24785);
xor UO_2536 (O_2536,N_24405,N_24959);
xnor UO_2537 (O_2537,N_24012,N_24887);
nor UO_2538 (O_2538,N_24546,N_24444);
nor UO_2539 (O_2539,N_24240,N_24053);
nand UO_2540 (O_2540,N_24457,N_24971);
and UO_2541 (O_2541,N_24559,N_24309);
xor UO_2542 (O_2542,N_24663,N_24808);
or UO_2543 (O_2543,N_24499,N_24295);
xor UO_2544 (O_2544,N_24341,N_24945);
and UO_2545 (O_2545,N_24278,N_24876);
nor UO_2546 (O_2546,N_24007,N_24711);
nand UO_2547 (O_2547,N_24283,N_24279);
or UO_2548 (O_2548,N_24069,N_24497);
xnor UO_2549 (O_2549,N_24794,N_24337);
nand UO_2550 (O_2550,N_24317,N_24260);
xor UO_2551 (O_2551,N_24778,N_24497);
nor UO_2552 (O_2552,N_24883,N_24385);
nand UO_2553 (O_2553,N_24350,N_24362);
nand UO_2554 (O_2554,N_24197,N_24723);
nor UO_2555 (O_2555,N_24849,N_24817);
or UO_2556 (O_2556,N_24222,N_24228);
xor UO_2557 (O_2557,N_24238,N_24799);
nor UO_2558 (O_2558,N_24947,N_24224);
nor UO_2559 (O_2559,N_24897,N_24444);
and UO_2560 (O_2560,N_24711,N_24830);
or UO_2561 (O_2561,N_24164,N_24256);
xnor UO_2562 (O_2562,N_24373,N_24778);
and UO_2563 (O_2563,N_24213,N_24777);
or UO_2564 (O_2564,N_24548,N_24671);
xor UO_2565 (O_2565,N_24331,N_24320);
nand UO_2566 (O_2566,N_24029,N_24635);
or UO_2567 (O_2567,N_24248,N_24235);
and UO_2568 (O_2568,N_24369,N_24955);
or UO_2569 (O_2569,N_24154,N_24437);
nand UO_2570 (O_2570,N_24409,N_24710);
xnor UO_2571 (O_2571,N_24395,N_24248);
xnor UO_2572 (O_2572,N_24077,N_24751);
nand UO_2573 (O_2573,N_24143,N_24936);
and UO_2574 (O_2574,N_24629,N_24821);
nor UO_2575 (O_2575,N_24985,N_24317);
nor UO_2576 (O_2576,N_24570,N_24244);
nor UO_2577 (O_2577,N_24383,N_24134);
nor UO_2578 (O_2578,N_24220,N_24847);
or UO_2579 (O_2579,N_24514,N_24190);
and UO_2580 (O_2580,N_24169,N_24155);
or UO_2581 (O_2581,N_24908,N_24777);
and UO_2582 (O_2582,N_24566,N_24984);
or UO_2583 (O_2583,N_24908,N_24885);
nand UO_2584 (O_2584,N_24950,N_24821);
nor UO_2585 (O_2585,N_24413,N_24811);
and UO_2586 (O_2586,N_24936,N_24697);
and UO_2587 (O_2587,N_24641,N_24668);
xor UO_2588 (O_2588,N_24980,N_24434);
or UO_2589 (O_2589,N_24063,N_24711);
nand UO_2590 (O_2590,N_24626,N_24292);
or UO_2591 (O_2591,N_24602,N_24501);
nor UO_2592 (O_2592,N_24720,N_24454);
nand UO_2593 (O_2593,N_24773,N_24181);
or UO_2594 (O_2594,N_24247,N_24737);
or UO_2595 (O_2595,N_24807,N_24980);
or UO_2596 (O_2596,N_24570,N_24387);
nand UO_2597 (O_2597,N_24231,N_24210);
nor UO_2598 (O_2598,N_24021,N_24813);
or UO_2599 (O_2599,N_24581,N_24434);
xor UO_2600 (O_2600,N_24526,N_24031);
and UO_2601 (O_2601,N_24870,N_24875);
and UO_2602 (O_2602,N_24433,N_24143);
nor UO_2603 (O_2603,N_24055,N_24543);
xnor UO_2604 (O_2604,N_24260,N_24398);
nand UO_2605 (O_2605,N_24570,N_24527);
and UO_2606 (O_2606,N_24796,N_24438);
or UO_2607 (O_2607,N_24118,N_24729);
nor UO_2608 (O_2608,N_24009,N_24481);
nand UO_2609 (O_2609,N_24471,N_24818);
nor UO_2610 (O_2610,N_24869,N_24816);
nand UO_2611 (O_2611,N_24758,N_24108);
or UO_2612 (O_2612,N_24484,N_24107);
or UO_2613 (O_2613,N_24774,N_24572);
nor UO_2614 (O_2614,N_24350,N_24699);
xnor UO_2615 (O_2615,N_24592,N_24270);
or UO_2616 (O_2616,N_24264,N_24549);
and UO_2617 (O_2617,N_24828,N_24261);
and UO_2618 (O_2618,N_24955,N_24126);
and UO_2619 (O_2619,N_24252,N_24503);
xor UO_2620 (O_2620,N_24934,N_24497);
nor UO_2621 (O_2621,N_24946,N_24345);
and UO_2622 (O_2622,N_24497,N_24743);
and UO_2623 (O_2623,N_24676,N_24857);
xor UO_2624 (O_2624,N_24171,N_24713);
nor UO_2625 (O_2625,N_24521,N_24175);
or UO_2626 (O_2626,N_24384,N_24662);
nand UO_2627 (O_2627,N_24786,N_24561);
xnor UO_2628 (O_2628,N_24965,N_24294);
nor UO_2629 (O_2629,N_24916,N_24041);
or UO_2630 (O_2630,N_24849,N_24291);
and UO_2631 (O_2631,N_24948,N_24119);
nand UO_2632 (O_2632,N_24462,N_24902);
or UO_2633 (O_2633,N_24880,N_24197);
xor UO_2634 (O_2634,N_24108,N_24775);
xor UO_2635 (O_2635,N_24086,N_24646);
nor UO_2636 (O_2636,N_24026,N_24746);
xnor UO_2637 (O_2637,N_24232,N_24438);
xnor UO_2638 (O_2638,N_24904,N_24415);
or UO_2639 (O_2639,N_24881,N_24323);
nand UO_2640 (O_2640,N_24325,N_24915);
nand UO_2641 (O_2641,N_24302,N_24530);
xor UO_2642 (O_2642,N_24523,N_24195);
or UO_2643 (O_2643,N_24679,N_24193);
xor UO_2644 (O_2644,N_24768,N_24104);
or UO_2645 (O_2645,N_24010,N_24361);
nand UO_2646 (O_2646,N_24757,N_24425);
xnor UO_2647 (O_2647,N_24961,N_24018);
or UO_2648 (O_2648,N_24946,N_24473);
xnor UO_2649 (O_2649,N_24982,N_24980);
nand UO_2650 (O_2650,N_24908,N_24051);
nor UO_2651 (O_2651,N_24334,N_24223);
xnor UO_2652 (O_2652,N_24931,N_24600);
and UO_2653 (O_2653,N_24432,N_24390);
and UO_2654 (O_2654,N_24244,N_24957);
nand UO_2655 (O_2655,N_24608,N_24396);
xor UO_2656 (O_2656,N_24363,N_24925);
nor UO_2657 (O_2657,N_24721,N_24183);
xor UO_2658 (O_2658,N_24308,N_24059);
nor UO_2659 (O_2659,N_24516,N_24957);
xor UO_2660 (O_2660,N_24099,N_24387);
and UO_2661 (O_2661,N_24668,N_24828);
or UO_2662 (O_2662,N_24364,N_24558);
or UO_2663 (O_2663,N_24753,N_24962);
nand UO_2664 (O_2664,N_24000,N_24243);
nor UO_2665 (O_2665,N_24812,N_24071);
nor UO_2666 (O_2666,N_24983,N_24636);
nor UO_2667 (O_2667,N_24967,N_24279);
nand UO_2668 (O_2668,N_24014,N_24695);
nor UO_2669 (O_2669,N_24317,N_24106);
or UO_2670 (O_2670,N_24813,N_24235);
and UO_2671 (O_2671,N_24755,N_24228);
or UO_2672 (O_2672,N_24564,N_24338);
and UO_2673 (O_2673,N_24338,N_24942);
nor UO_2674 (O_2674,N_24074,N_24749);
or UO_2675 (O_2675,N_24155,N_24824);
or UO_2676 (O_2676,N_24817,N_24054);
and UO_2677 (O_2677,N_24284,N_24193);
and UO_2678 (O_2678,N_24268,N_24074);
nor UO_2679 (O_2679,N_24942,N_24867);
and UO_2680 (O_2680,N_24161,N_24288);
nor UO_2681 (O_2681,N_24423,N_24796);
or UO_2682 (O_2682,N_24799,N_24714);
nor UO_2683 (O_2683,N_24815,N_24501);
nor UO_2684 (O_2684,N_24298,N_24801);
nor UO_2685 (O_2685,N_24387,N_24652);
nor UO_2686 (O_2686,N_24285,N_24143);
nor UO_2687 (O_2687,N_24167,N_24132);
and UO_2688 (O_2688,N_24276,N_24748);
nor UO_2689 (O_2689,N_24133,N_24892);
xor UO_2690 (O_2690,N_24685,N_24597);
nand UO_2691 (O_2691,N_24744,N_24617);
or UO_2692 (O_2692,N_24713,N_24374);
or UO_2693 (O_2693,N_24473,N_24018);
and UO_2694 (O_2694,N_24466,N_24001);
nand UO_2695 (O_2695,N_24333,N_24291);
nand UO_2696 (O_2696,N_24408,N_24988);
xor UO_2697 (O_2697,N_24140,N_24945);
xnor UO_2698 (O_2698,N_24220,N_24095);
nand UO_2699 (O_2699,N_24600,N_24078);
or UO_2700 (O_2700,N_24510,N_24957);
xnor UO_2701 (O_2701,N_24459,N_24665);
xor UO_2702 (O_2702,N_24481,N_24550);
or UO_2703 (O_2703,N_24726,N_24482);
nand UO_2704 (O_2704,N_24067,N_24219);
xor UO_2705 (O_2705,N_24001,N_24605);
nand UO_2706 (O_2706,N_24715,N_24839);
or UO_2707 (O_2707,N_24688,N_24617);
xor UO_2708 (O_2708,N_24647,N_24246);
xnor UO_2709 (O_2709,N_24853,N_24044);
nor UO_2710 (O_2710,N_24039,N_24362);
nand UO_2711 (O_2711,N_24527,N_24295);
and UO_2712 (O_2712,N_24252,N_24249);
xnor UO_2713 (O_2713,N_24325,N_24251);
xor UO_2714 (O_2714,N_24301,N_24433);
nor UO_2715 (O_2715,N_24460,N_24977);
and UO_2716 (O_2716,N_24496,N_24659);
xor UO_2717 (O_2717,N_24023,N_24237);
nand UO_2718 (O_2718,N_24419,N_24244);
nor UO_2719 (O_2719,N_24268,N_24100);
or UO_2720 (O_2720,N_24566,N_24725);
nand UO_2721 (O_2721,N_24187,N_24500);
nor UO_2722 (O_2722,N_24326,N_24293);
or UO_2723 (O_2723,N_24629,N_24955);
nand UO_2724 (O_2724,N_24939,N_24680);
nand UO_2725 (O_2725,N_24797,N_24184);
nand UO_2726 (O_2726,N_24042,N_24322);
and UO_2727 (O_2727,N_24181,N_24278);
or UO_2728 (O_2728,N_24191,N_24158);
xnor UO_2729 (O_2729,N_24618,N_24592);
and UO_2730 (O_2730,N_24879,N_24887);
nand UO_2731 (O_2731,N_24284,N_24922);
nand UO_2732 (O_2732,N_24710,N_24363);
and UO_2733 (O_2733,N_24737,N_24991);
and UO_2734 (O_2734,N_24538,N_24994);
nor UO_2735 (O_2735,N_24681,N_24771);
and UO_2736 (O_2736,N_24740,N_24504);
xor UO_2737 (O_2737,N_24426,N_24813);
and UO_2738 (O_2738,N_24754,N_24844);
or UO_2739 (O_2739,N_24740,N_24144);
and UO_2740 (O_2740,N_24648,N_24759);
nor UO_2741 (O_2741,N_24073,N_24918);
or UO_2742 (O_2742,N_24037,N_24648);
and UO_2743 (O_2743,N_24424,N_24995);
or UO_2744 (O_2744,N_24082,N_24626);
or UO_2745 (O_2745,N_24589,N_24702);
xnor UO_2746 (O_2746,N_24428,N_24802);
or UO_2747 (O_2747,N_24942,N_24153);
and UO_2748 (O_2748,N_24796,N_24790);
nand UO_2749 (O_2749,N_24918,N_24739);
xor UO_2750 (O_2750,N_24931,N_24645);
nor UO_2751 (O_2751,N_24302,N_24099);
nor UO_2752 (O_2752,N_24850,N_24396);
nor UO_2753 (O_2753,N_24807,N_24739);
and UO_2754 (O_2754,N_24755,N_24187);
nor UO_2755 (O_2755,N_24911,N_24057);
nor UO_2756 (O_2756,N_24135,N_24064);
or UO_2757 (O_2757,N_24397,N_24438);
nor UO_2758 (O_2758,N_24619,N_24530);
xor UO_2759 (O_2759,N_24473,N_24119);
xor UO_2760 (O_2760,N_24804,N_24363);
nand UO_2761 (O_2761,N_24614,N_24671);
nor UO_2762 (O_2762,N_24007,N_24901);
nor UO_2763 (O_2763,N_24134,N_24115);
or UO_2764 (O_2764,N_24942,N_24502);
nor UO_2765 (O_2765,N_24266,N_24452);
nor UO_2766 (O_2766,N_24904,N_24850);
nor UO_2767 (O_2767,N_24141,N_24545);
nand UO_2768 (O_2768,N_24174,N_24554);
and UO_2769 (O_2769,N_24743,N_24691);
nor UO_2770 (O_2770,N_24561,N_24579);
nor UO_2771 (O_2771,N_24488,N_24777);
or UO_2772 (O_2772,N_24332,N_24739);
nor UO_2773 (O_2773,N_24154,N_24183);
nand UO_2774 (O_2774,N_24385,N_24220);
xor UO_2775 (O_2775,N_24618,N_24111);
or UO_2776 (O_2776,N_24493,N_24954);
or UO_2777 (O_2777,N_24181,N_24035);
nor UO_2778 (O_2778,N_24683,N_24918);
xor UO_2779 (O_2779,N_24015,N_24211);
xnor UO_2780 (O_2780,N_24030,N_24925);
nand UO_2781 (O_2781,N_24565,N_24286);
xnor UO_2782 (O_2782,N_24914,N_24080);
nor UO_2783 (O_2783,N_24690,N_24185);
nand UO_2784 (O_2784,N_24047,N_24936);
or UO_2785 (O_2785,N_24590,N_24939);
nand UO_2786 (O_2786,N_24257,N_24437);
and UO_2787 (O_2787,N_24029,N_24134);
or UO_2788 (O_2788,N_24458,N_24275);
nor UO_2789 (O_2789,N_24819,N_24844);
xnor UO_2790 (O_2790,N_24948,N_24205);
nor UO_2791 (O_2791,N_24501,N_24755);
nand UO_2792 (O_2792,N_24184,N_24266);
nor UO_2793 (O_2793,N_24711,N_24089);
nand UO_2794 (O_2794,N_24095,N_24629);
and UO_2795 (O_2795,N_24114,N_24438);
nor UO_2796 (O_2796,N_24921,N_24930);
or UO_2797 (O_2797,N_24484,N_24941);
nor UO_2798 (O_2798,N_24830,N_24639);
or UO_2799 (O_2799,N_24172,N_24157);
nor UO_2800 (O_2800,N_24844,N_24508);
nor UO_2801 (O_2801,N_24448,N_24833);
and UO_2802 (O_2802,N_24780,N_24752);
or UO_2803 (O_2803,N_24830,N_24453);
and UO_2804 (O_2804,N_24892,N_24269);
and UO_2805 (O_2805,N_24783,N_24136);
xor UO_2806 (O_2806,N_24524,N_24968);
nor UO_2807 (O_2807,N_24776,N_24260);
nand UO_2808 (O_2808,N_24374,N_24591);
nand UO_2809 (O_2809,N_24520,N_24857);
nand UO_2810 (O_2810,N_24283,N_24407);
nor UO_2811 (O_2811,N_24946,N_24433);
nor UO_2812 (O_2812,N_24219,N_24554);
and UO_2813 (O_2813,N_24167,N_24479);
and UO_2814 (O_2814,N_24015,N_24071);
nand UO_2815 (O_2815,N_24156,N_24995);
nand UO_2816 (O_2816,N_24609,N_24929);
and UO_2817 (O_2817,N_24295,N_24517);
nand UO_2818 (O_2818,N_24438,N_24069);
and UO_2819 (O_2819,N_24348,N_24002);
and UO_2820 (O_2820,N_24482,N_24539);
or UO_2821 (O_2821,N_24627,N_24685);
xor UO_2822 (O_2822,N_24565,N_24549);
or UO_2823 (O_2823,N_24676,N_24725);
nor UO_2824 (O_2824,N_24043,N_24715);
xnor UO_2825 (O_2825,N_24094,N_24058);
nor UO_2826 (O_2826,N_24841,N_24028);
nand UO_2827 (O_2827,N_24004,N_24130);
and UO_2828 (O_2828,N_24323,N_24950);
nand UO_2829 (O_2829,N_24641,N_24899);
and UO_2830 (O_2830,N_24364,N_24112);
or UO_2831 (O_2831,N_24077,N_24838);
xor UO_2832 (O_2832,N_24855,N_24516);
nor UO_2833 (O_2833,N_24497,N_24723);
and UO_2834 (O_2834,N_24082,N_24089);
nand UO_2835 (O_2835,N_24351,N_24935);
or UO_2836 (O_2836,N_24060,N_24897);
and UO_2837 (O_2837,N_24840,N_24145);
nor UO_2838 (O_2838,N_24789,N_24317);
nor UO_2839 (O_2839,N_24984,N_24681);
nor UO_2840 (O_2840,N_24387,N_24950);
xnor UO_2841 (O_2841,N_24602,N_24481);
nand UO_2842 (O_2842,N_24216,N_24895);
or UO_2843 (O_2843,N_24232,N_24077);
xnor UO_2844 (O_2844,N_24374,N_24718);
or UO_2845 (O_2845,N_24061,N_24479);
nand UO_2846 (O_2846,N_24459,N_24960);
nand UO_2847 (O_2847,N_24057,N_24269);
nor UO_2848 (O_2848,N_24219,N_24969);
or UO_2849 (O_2849,N_24668,N_24394);
or UO_2850 (O_2850,N_24983,N_24932);
and UO_2851 (O_2851,N_24131,N_24163);
nor UO_2852 (O_2852,N_24117,N_24350);
and UO_2853 (O_2853,N_24630,N_24394);
and UO_2854 (O_2854,N_24174,N_24271);
nor UO_2855 (O_2855,N_24641,N_24494);
and UO_2856 (O_2856,N_24258,N_24290);
or UO_2857 (O_2857,N_24178,N_24966);
nor UO_2858 (O_2858,N_24100,N_24209);
or UO_2859 (O_2859,N_24036,N_24308);
xor UO_2860 (O_2860,N_24283,N_24960);
or UO_2861 (O_2861,N_24856,N_24896);
nor UO_2862 (O_2862,N_24834,N_24639);
nand UO_2863 (O_2863,N_24511,N_24313);
nand UO_2864 (O_2864,N_24881,N_24221);
nand UO_2865 (O_2865,N_24808,N_24613);
and UO_2866 (O_2866,N_24372,N_24641);
nand UO_2867 (O_2867,N_24914,N_24015);
or UO_2868 (O_2868,N_24108,N_24617);
or UO_2869 (O_2869,N_24196,N_24953);
nor UO_2870 (O_2870,N_24727,N_24899);
xnor UO_2871 (O_2871,N_24404,N_24708);
nand UO_2872 (O_2872,N_24518,N_24341);
and UO_2873 (O_2873,N_24817,N_24226);
xor UO_2874 (O_2874,N_24556,N_24403);
xor UO_2875 (O_2875,N_24909,N_24089);
nor UO_2876 (O_2876,N_24204,N_24011);
and UO_2877 (O_2877,N_24779,N_24676);
nand UO_2878 (O_2878,N_24715,N_24534);
or UO_2879 (O_2879,N_24468,N_24517);
xnor UO_2880 (O_2880,N_24837,N_24743);
nand UO_2881 (O_2881,N_24281,N_24605);
nand UO_2882 (O_2882,N_24266,N_24893);
nor UO_2883 (O_2883,N_24654,N_24373);
or UO_2884 (O_2884,N_24597,N_24757);
or UO_2885 (O_2885,N_24792,N_24832);
or UO_2886 (O_2886,N_24130,N_24701);
xor UO_2887 (O_2887,N_24645,N_24731);
or UO_2888 (O_2888,N_24862,N_24942);
nor UO_2889 (O_2889,N_24517,N_24742);
nand UO_2890 (O_2890,N_24934,N_24430);
xor UO_2891 (O_2891,N_24231,N_24847);
nand UO_2892 (O_2892,N_24736,N_24654);
nand UO_2893 (O_2893,N_24150,N_24528);
nor UO_2894 (O_2894,N_24436,N_24301);
and UO_2895 (O_2895,N_24375,N_24922);
nand UO_2896 (O_2896,N_24302,N_24486);
and UO_2897 (O_2897,N_24588,N_24779);
xnor UO_2898 (O_2898,N_24228,N_24138);
xor UO_2899 (O_2899,N_24442,N_24393);
or UO_2900 (O_2900,N_24454,N_24485);
or UO_2901 (O_2901,N_24832,N_24664);
nand UO_2902 (O_2902,N_24740,N_24171);
xor UO_2903 (O_2903,N_24525,N_24708);
xor UO_2904 (O_2904,N_24715,N_24551);
or UO_2905 (O_2905,N_24563,N_24559);
nor UO_2906 (O_2906,N_24677,N_24799);
nand UO_2907 (O_2907,N_24871,N_24608);
nand UO_2908 (O_2908,N_24458,N_24933);
nor UO_2909 (O_2909,N_24512,N_24529);
nor UO_2910 (O_2910,N_24297,N_24789);
nand UO_2911 (O_2911,N_24125,N_24092);
nand UO_2912 (O_2912,N_24169,N_24815);
xor UO_2913 (O_2913,N_24543,N_24327);
nand UO_2914 (O_2914,N_24653,N_24792);
nand UO_2915 (O_2915,N_24039,N_24473);
or UO_2916 (O_2916,N_24952,N_24773);
nand UO_2917 (O_2917,N_24601,N_24081);
xor UO_2918 (O_2918,N_24670,N_24612);
xor UO_2919 (O_2919,N_24782,N_24211);
or UO_2920 (O_2920,N_24166,N_24448);
or UO_2921 (O_2921,N_24040,N_24805);
xor UO_2922 (O_2922,N_24955,N_24005);
xor UO_2923 (O_2923,N_24861,N_24258);
nor UO_2924 (O_2924,N_24215,N_24633);
nand UO_2925 (O_2925,N_24059,N_24686);
xor UO_2926 (O_2926,N_24986,N_24948);
nand UO_2927 (O_2927,N_24030,N_24743);
xnor UO_2928 (O_2928,N_24786,N_24206);
nand UO_2929 (O_2929,N_24902,N_24044);
nand UO_2930 (O_2930,N_24896,N_24105);
nand UO_2931 (O_2931,N_24002,N_24459);
nand UO_2932 (O_2932,N_24505,N_24770);
nor UO_2933 (O_2933,N_24997,N_24065);
or UO_2934 (O_2934,N_24368,N_24833);
or UO_2935 (O_2935,N_24760,N_24309);
and UO_2936 (O_2936,N_24425,N_24530);
or UO_2937 (O_2937,N_24196,N_24211);
xnor UO_2938 (O_2938,N_24583,N_24864);
xnor UO_2939 (O_2939,N_24692,N_24127);
xnor UO_2940 (O_2940,N_24135,N_24804);
nand UO_2941 (O_2941,N_24180,N_24801);
and UO_2942 (O_2942,N_24441,N_24413);
and UO_2943 (O_2943,N_24420,N_24086);
and UO_2944 (O_2944,N_24526,N_24702);
nand UO_2945 (O_2945,N_24206,N_24957);
or UO_2946 (O_2946,N_24527,N_24585);
nand UO_2947 (O_2947,N_24198,N_24673);
and UO_2948 (O_2948,N_24943,N_24418);
nor UO_2949 (O_2949,N_24022,N_24497);
or UO_2950 (O_2950,N_24691,N_24902);
nand UO_2951 (O_2951,N_24011,N_24703);
or UO_2952 (O_2952,N_24472,N_24848);
nand UO_2953 (O_2953,N_24757,N_24729);
xnor UO_2954 (O_2954,N_24444,N_24376);
and UO_2955 (O_2955,N_24465,N_24615);
nand UO_2956 (O_2956,N_24711,N_24207);
xor UO_2957 (O_2957,N_24045,N_24786);
xor UO_2958 (O_2958,N_24778,N_24738);
and UO_2959 (O_2959,N_24510,N_24945);
and UO_2960 (O_2960,N_24516,N_24458);
xnor UO_2961 (O_2961,N_24822,N_24881);
and UO_2962 (O_2962,N_24686,N_24814);
xnor UO_2963 (O_2963,N_24162,N_24927);
nor UO_2964 (O_2964,N_24347,N_24817);
and UO_2965 (O_2965,N_24419,N_24537);
nand UO_2966 (O_2966,N_24681,N_24838);
and UO_2967 (O_2967,N_24554,N_24560);
or UO_2968 (O_2968,N_24642,N_24786);
nor UO_2969 (O_2969,N_24285,N_24200);
and UO_2970 (O_2970,N_24722,N_24236);
nand UO_2971 (O_2971,N_24468,N_24865);
and UO_2972 (O_2972,N_24309,N_24494);
xor UO_2973 (O_2973,N_24300,N_24475);
nand UO_2974 (O_2974,N_24749,N_24582);
nand UO_2975 (O_2975,N_24895,N_24002);
and UO_2976 (O_2976,N_24404,N_24943);
xnor UO_2977 (O_2977,N_24411,N_24949);
xnor UO_2978 (O_2978,N_24237,N_24710);
xnor UO_2979 (O_2979,N_24632,N_24090);
or UO_2980 (O_2980,N_24202,N_24822);
or UO_2981 (O_2981,N_24190,N_24666);
xor UO_2982 (O_2982,N_24613,N_24292);
and UO_2983 (O_2983,N_24014,N_24455);
nor UO_2984 (O_2984,N_24902,N_24089);
nand UO_2985 (O_2985,N_24777,N_24211);
nor UO_2986 (O_2986,N_24175,N_24622);
nand UO_2987 (O_2987,N_24845,N_24367);
or UO_2988 (O_2988,N_24779,N_24033);
xor UO_2989 (O_2989,N_24572,N_24378);
xnor UO_2990 (O_2990,N_24937,N_24890);
xor UO_2991 (O_2991,N_24916,N_24496);
or UO_2992 (O_2992,N_24972,N_24528);
and UO_2993 (O_2993,N_24417,N_24138);
and UO_2994 (O_2994,N_24339,N_24209);
and UO_2995 (O_2995,N_24672,N_24010);
and UO_2996 (O_2996,N_24828,N_24590);
xor UO_2997 (O_2997,N_24868,N_24135);
nand UO_2998 (O_2998,N_24513,N_24312);
nor UO_2999 (O_2999,N_24889,N_24413);
endmodule