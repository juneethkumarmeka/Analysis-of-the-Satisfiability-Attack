module basic_500_3000_500_30_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_251,In_481);
xor U1 (N_1,In_165,In_443);
or U2 (N_2,In_321,In_489);
or U3 (N_3,In_381,In_497);
or U4 (N_4,In_88,In_263);
or U5 (N_5,In_142,In_341);
and U6 (N_6,In_22,In_300);
and U7 (N_7,In_477,In_408);
xor U8 (N_8,In_417,In_322);
xor U9 (N_9,In_178,In_224);
nor U10 (N_10,In_91,In_284);
and U11 (N_11,In_77,In_375);
or U12 (N_12,In_498,In_236);
and U13 (N_13,In_266,In_84);
nand U14 (N_14,In_406,In_370);
nor U15 (N_15,In_256,In_76);
and U16 (N_16,In_439,In_136);
xnor U17 (N_17,In_237,In_380);
or U18 (N_18,In_289,In_253);
nor U19 (N_19,In_315,In_60);
and U20 (N_20,In_94,In_350);
or U21 (N_21,In_86,In_271);
and U22 (N_22,In_106,In_59);
nand U23 (N_23,In_97,In_391);
or U24 (N_24,In_376,In_234);
nand U25 (N_25,In_435,In_105);
xor U26 (N_26,In_199,In_451);
or U27 (N_27,In_27,In_495);
nand U28 (N_28,In_385,In_50);
xnor U29 (N_29,In_14,In_378);
xor U30 (N_30,In_265,In_482);
nand U31 (N_31,In_144,In_389);
nand U32 (N_32,In_467,In_273);
nor U33 (N_33,In_145,In_334);
xnor U34 (N_34,In_67,In_302);
nor U35 (N_35,In_281,In_64);
nand U36 (N_36,In_261,In_311);
nand U37 (N_37,In_112,In_171);
nand U38 (N_38,In_411,In_173);
and U39 (N_39,In_398,In_195);
and U40 (N_40,In_15,In_9);
nor U41 (N_41,In_221,In_464);
or U42 (N_42,In_348,In_137);
and U43 (N_43,In_146,In_351);
and U44 (N_44,In_201,In_213);
nand U45 (N_45,In_222,In_499);
nand U46 (N_46,In_286,In_107);
or U47 (N_47,In_329,In_190);
and U48 (N_48,In_231,In_241);
and U49 (N_49,In_465,In_421);
xnor U50 (N_50,In_364,In_245);
or U51 (N_51,In_38,In_353);
xor U52 (N_52,In_139,In_78);
and U53 (N_53,In_330,In_423);
xnor U54 (N_54,In_327,In_373);
nand U55 (N_55,In_480,In_39);
xnor U56 (N_56,In_17,In_43);
nand U57 (N_57,In_243,In_57);
nor U58 (N_58,In_155,In_83);
nor U59 (N_59,In_470,In_153);
or U60 (N_60,In_238,In_156);
xnor U61 (N_61,In_340,In_187);
nor U62 (N_62,In_130,In_129);
or U63 (N_63,In_184,In_242);
nor U64 (N_64,In_328,In_276);
xor U65 (N_65,In_349,In_100);
xnor U66 (N_66,In_157,In_210);
nand U67 (N_67,In_432,In_298);
and U68 (N_68,In_401,In_407);
or U69 (N_69,In_384,In_475);
or U70 (N_70,In_186,In_388);
xor U71 (N_71,In_62,In_496);
xnor U72 (N_72,In_49,In_240);
nand U73 (N_73,In_175,In_205);
or U74 (N_74,In_471,In_312);
and U75 (N_75,In_377,In_249);
nor U76 (N_76,In_361,In_197);
nand U77 (N_77,In_454,In_424);
nor U78 (N_78,In_1,In_202);
and U79 (N_79,In_40,In_152);
nand U80 (N_80,In_441,In_147);
nor U81 (N_81,In_434,In_345);
or U82 (N_82,In_126,In_306);
and U83 (N_83,In_32,In_396);
xor U84 (N_84,In_230,In_487);
and U85 (N_85,In_93,In_272);
nor U86 (N_86,In_232,In_10);
and U87 (N_87,In_324,In_490);
nand U88 (N_88,In_70,In_397);
xor U89 (N_89,In_422,In_73);
and U90 (N_90,In_419,In_358);
or U91 (N_91,In_71,In_102);
or U92 (N_92,In_404,In_479);
or U93 (N_93,In_19,In_274);
or U94 (N_94,In_218,In_257);
nand U95 (N_95,In_176,In_214);
and U96 (N_96,In_239,In_399);
xnor U97 (N_97,In_437,In_293);
and U98 (N_98,In_275,In_65);
nor U99 (N_99,In_34,In_486);
or U100 (N_100,N_84,In_191);
or U101 (N_101,N_57,In_430);
nand U102 (N_102,In_162,In_356);
or U103 (N_103,In_121,N_78);
xor U104 (N_104,In_248,In_25);
nor U105 (N_105,In_29,N_1);
nand U106 (N_106,In_81,In_414);
nor U107 (N_107,In_82,N_35);
nor U108 (N_108,In_41,In_143);
or U109 (N_109,In_267,N_31);
xor U110 (N_110,In_89,N_12);
xor U111 (N_111,In_123,N_0);
nand U112 (N_112,N_6,In_270);
and U113 (N_113,In_444,In_336);
nand U114 (N_114,In_402,In_24);
nor U115 (N_115,N_89,In_51);
nand U116 (N_116,N_90,N_55);
nand U117 (N_117,In_357,In_135);
and U118 (N_118,N_41,N_98);
or U119 (N_119,In_13,In_409);
nand U120 (N_120,In_198,N_24);
and U121 (N_121,In_87,In_374);
and U122 (N_122,N_66,In_48);
nand U123 (N_123,In_288,In_203);
nor U124 (N_124,In_285,In_448);
and U125 (N_125,In_117,In_119);
xnor U126 (N_126,In_254,In_235);
xnor U127 (N_127,N_5,In_193);
and U128 (N_128,In_220,N_21);
nor U129 (N_129,N_86,In_352);
nor U130 (N_130,In_339,In_154);
nor U131 (N_131,N_11,In_20);
nor U132 (N_132,In_368,N_65);
nand U133 (N_133,In_438,In_447);
nor U134 (N_134,N_75,In_194);
xnor U135 (N_135,N_16,N_58);
xnor U136 (N_136,In_440,N_17);
and U137 (N_137,In_168,In_363);
or U138 (N_138,In_283,N_64);
and U139 (N_139,In_305,N_15);
nor U140 (N_140,In_11,N_74);
nor U141 (N_141,In_308,In_114);
nand U142 (N_142,N_18,In_69);
or U143 (N_143,In_200,N_29);
nor U144 (N_144,In_468,N_30);
nand U145 (N_145,In_189,In_75);
nand U146 (N_146,In_405,In_113);
or U147 (N_147,N_62,In_244);
or U148 (N_148,N_25,In_295);
and U149 (N_149,In_208,In_54);
nand U150 (N_150,In_463,In_268);
nand U151 (N_151,In_460,N_37);
nor U152 (N_152,N_69,N_96);
nor U153 (N_153,N_4,In_160);
and U154 (N_154,In_4,N_95);
xor U155 (N_155,N_99,In_151);
and U156 (N_156,In_138,In_412);
nand U157 (N_157,In_46,In_456);
and U158 (N_158,In_92,In_120);
nor U159 (N_159,In_252,In_56);
or U160 (N_160,In_204,In_403);
nor U161 (N_161,In_260,In_333);
nor U162 (N_162,In_418,In_37);
nor U163 (N_163,N_26,In_354);
and U164 (N_164,In_280,In_453);
nand U165 (N_165,In_346,In_335);
or U166 (N_166,N_94,In_318);
and U167 (N_167,N_48,In_85);
xnor U168 (N_168,In_278,In_258);
nor U169 (N_169,In_316,N_44);
nor U170 (N_170,In_294,In_392);
nor U171 (N_171,In_18,In_416);
xor U172 (N_172,In_192,In_35);
nor U173 (N_173,In_183,In_469);
and U174 (N_174,N_47,In_33);
and U175 (N_175,In_319,In_299);
xor U176 (N_176,In_371,In_359);
nor U177 (N_177,In_28,In_413);
or U178 (N_178,In_6,In_255);
xnor U179 (N_179,In_449,In_8);
xnor U180 (N_180,N_27,N_14);
or U181 (N_181,In_95,In_90);
nor U182 (N_182,In_338,N_2);
or U183 (N_183,In_303,In_337);
nand U184 (N_184,In_233,N_56);
xnor U185 (N_185,N_49,N_67);
nor U186 (N_186,In_317,In_291);
xnor U187 (N_187,In_229,In_124);
xnor U188 (N_188,In_492,N_63);
nand U189 (N_189,In_149,In_410);
xor U190 (N_190,In_109,N_13);
and U191 (N_191,In_219,In_279);
or U192 (N_192,N_28,In_30);
and U193 (N_193,In_206,In_2);
nor U194 (N_194,N_34,In_360);
and U195 (N_195,N_88,N_7);
and U196 (N_196,In_7,In_172);
nand U197 (N_197,In_159,In_287);
nor U198 (N_198,N_81,In_188);
xnor U199 (N_199,In_494,In_72);
xor U200 (N_200,In_478,In_170);
nand U201 (N_201,N_124,In_400);
nand U202 (N_202,In_382,In_128);
nand U203 (N_203,N_137,In_132);
nand U204 (N_204,In_31,N_167);
and U205 (N_205,In_420,N_150);
and U206 (N_206,In_223,N_120);
and U207 (N_207,N_9,In_45);
or U208 (N_208,N_52,In_290);
or U209 (N_209,N_106,N_103);
nor U210 (N_210,N_146,In_55);
nand U211 (N_211,N_130,N_59);
or U212 (N_212,In_394,N_197);
nand U213 (N_213,N_113,N_85);
or U214 (N_214,N_195,N_165);
xnor U215 (N_215,N_36,N_40);
xor U216 (N_216,N_184,In_379);
nand U217 (N_217,N_193,N_73);
xor U218 (N_218,In_466,In_169);
and U219 (N_219,N_169,In_433);
nor U220 (N_220,In_247,In_446);
nand U221 (N_221,N_91,In_5);
or U222 (N_222,In_68,In_127);
and U223 (N_223,In_125,N_178);
nand U224 (N_224,N_163,In_63);
or U225 (N_225,In_344,N_155);
or U226 (N_226,N_140,In_429);
xor U227 (N_227,In_485,In_313);
nor U228 (N_228,N_187,N_61);
or U229 (N_229,In_342,In_179);
and U230 (N_230,In_326,N_151);
or U231 (N_231,N_46,In_150);
nor U232 (N_232,In_462,N_186);
or U233 (N_233,In_366,In_415);
and U234 (N_234,N_134,N_158);
nand U235 (N_235,In_161,In_343);
and U236 (N_236,In_185,In_457);
xor U237 (N_237,N_143,N_45);
and U238 (N_238,N_133,In_79);
nand U239 (N_239,In_450,N_147);
nand U240 (N_240,N_111,N_157);
nand U241 (N_241,N_182,N_180);
nand U242 (N_242,N_118,In_472);
or U243 (N_243,N_159,In_166);
nand U244 (N_244,In_292,In_111);
nor U245 (N_245,In_365,N_176);
nand U246 (N_246,N_183,N_132);
and U247 (N_247,N_50,In_332);
xnor U248 (N_248,N_177,In_80);
xor U249 (N_249,In_104,N_60);
or U250 (N_250,In_367,In_44);
or U251 (N_251,In_461,In_369);
nor U252 (N_252,In_174,N_68);
and U253 (N_253,In_211,In_386);
or U254 (N_254,In_331,N_114);
or U255 (N_255,N_54,In_0);
or U256 (N_256,N_142,N_79);
and U257 (N_257,N_80,N_102);
xor U258 (N_258,In_225,N_194);
nand U259 (N_259,In_395,In_428);
nor U260 (N_260,In_148,In_99);
and U261 (N_261,N_192,N_129);
and U262 (N_262,In_131,In_21);
nor U263 (N_263,In_309,N_119);
or U264 (N_264,In_42,In_262);
and U265 (N_265,N_110,In_431);
xor U266 (N_266,N_93,In_52);
nand U267 (N_267,In_53,N_76);
xor U268 (N_268,N_175,In_212);
or U269 (N_269,In_259,N_170);
nand U270 (N_270,In_133,N_168);
or U271 (N_271,In_488,In_296);
and U272 (N_272,In_476,In_304);
and U273 (N_273,N_190,In_250);
or U274 (N_274,In_181,In_297);
and U275 (N_275,N_181,N_107);
and U276 (N_276,In_459,In_96);
xnor U277 (N_277,In_158,In_246);
xor U278 (N_278,In_116,N_123);
and U279 (N_279,N_43,N_116);
xor U280 (N_280,In_445,N_138);
xnor U281 (N_281,In_310,In_427);
or U282 (N_282,N_188,In_167);
nor U283 (N_283,N_104,N_172);
xnor U284 (N_284,N_166,N_131);
and U285 (N_285,In_314,In_3);
nor U286 (N_286,N_185,In_36);
or U287 (N_287,In_458,N_8);
xnor U288 (N_288,N_112,In_118);
nand U289 (N_289,N_128,N_101);
nand U290 (N_290,N_83,N_160);
xnor U291 (N_291,In_307,In_301);
nor U292 (N_292,In_226,N_82);
or U293 (N_293,N_144,N_141);
nor U294 (N_294,N_117,N_198);
and U295 (N_295,N_174,N_38);
or U296 (N_296,N_20,In_436);
nor U297 (N_297,N_173,In_180);
nor U298 (N_298,N_23,In_141);
and U299 (N_299,N_191,In_493);
xor U300 (N_300,In_452,In_207);
or U301 (N_301,N_298,N_105);
or U302 (N_302,In_103,In_269);
xor U303 (N_303,N_256,N_115);
nand U304 (N_304,N_125,N_283);
xnor U305 (N_305,N_148,In_140);
nand U306 (N_306,In_163,N_145);
nor U307 (N_307,N_196,In_282);
or U308 (N_308,N_238,In_455);
nor U309 (N_309,In_209,In_47);
nor U310 (N_310,N_241,N_149);
nand U311 (N_311,N_275,N_126);
nand U312 (N_312,N_32,In_215);
nand U313 (N_313,N_214,In_227);
nor U314 (N_314,In_58,N_297);
nor U315 (N_315,N_289,N_276);
or U316 (N_316,N_156,N_154);
xor U317 (N_317,N_263,N_229);
or U318 (N_318,N_299,N_261);
and U319 (N_319,N_282,N_273);
xor U320 (N_320,In_491,N_72);
xnor U321 (N_321,N_219,N_162);
or U322 (N_322,N_260,N_230);
nor U323 (N_323,N_136,N_258);
or U324 (N_324,N_294,N_239);
nand U325 (N_325,N_262,N_100);
or U326 (N_326,N_237,N_267);
xor U327 (N_327,N_268,N_274);
and U328 (N_328,N_292,N_269);
or U329 (N_329,N_272,N_245);
nor U330 (N_330,N_242,N_221);
nor U331 (N_331,In_393,In_182);
nor U332 (N_332,N_135,In_355);
nor U333 (N_333,In_61,N_266);
nor U334 (N_334,In_347,N_71);
or U335 (N_335,N_209,N_220);
xnor U336 (N_336,N_291,N_202);
nand U337 (N_337,N_211,N_152);
and U338 (N_338,In_101,N_287);
nor U339 (N_339,N_207,N_252);
nand U340 (N_340,N_231,N_240);
nand U341 (N_341,N_253,N_246);
nor U342 (N_342,N_216,N_247);
and U343 (N_343,In_177,N_22);
or U344 (N_344,N_97,In_108);
nor U345 (N_345,N_127,In_277);
or U346 (N_346,In_66,N_277);
or U347 (N_347,In_383,N_121);
or U348 (N_348,N_53,N_248);
nor U349 (N_349,In_26,N_228);
or U350 (N_350,N_249,N_171);
xnor U351 (N_351,N_257,In_372);
xnor U352 (N_352,N_232,N_226);
nand U353 (N_353,N_224,N_285);
nand U354 (N_354,In_164,In_483);
xor U355 (N_355,N_244,N_109);
nand U356 (N_356,N_19,N_42);
and U357 (N_357,N_200,N_255);
nand U358 (N_358,N_233,N_278);
nand U359 (N_359,In_362,N_208);
or U360 (N_360,N_243,N_280);
and U361 (N_361,N_270,N_236);
or U362 (N_362,N_235,N_3);
xnor U363 (N_363,N_288,N_223);
nor U364 (N_364,In_74,N_203);
xor U365 (N_365,N_215,N_222);
xnor U366 (N_366,N_251,N_295);
and U367 (N_367,In_390,N_179);
nor U368 (N_368,N_279,N_108);
xor U369 (N_369,N_250,N_77);
or U370 (N_370,N_122,N_70);
or U371 (N_371,In_484,N_51);
xor U372 (N_372,In_473,N_212);
or U373 (N_373,In_228,In_98);
and U374 (N_374,N_33,N_210);
and U375 (N_375,In_323,In_196);
and U376 (N_376,N_92,N_254);
or U377 (N_377,N_87,In_115);
and U378 (N_378,In_12,N_264);
nand U379 (N_379,N_204,N_39);
nand U380 (N_380,N_259,N_234);
xor U381 (N_381,N_161,In_217);
or U382 (N_382,In_23,N_271);
xor U383 (N_383,N_201,N_218);
and U384 (N_384,In_264,N_225);
xor U385 (N_385,N_265,N_164);
and U386 (N_386,In_320,In_325);
nand U387 (N_387,N_284,In_110);
xor U388 (N_388,N_293,N_10);
or U389 (N_389,In_442,In_426);
nand U390 (N_390,N_227,N_205);
xnor U391 (N_391,N_189,In_425);
xnor U392 (N_392,In_134,N_281);
xnor U393 (N_393,In_216,In_387);
nand U394 (N_394,N_213,N_290);
nand U395 (N_395,In_16,In_474);
or U396 (N_396,N_217,N_199);
xor U397 (N_397,N_286,In_122);
nand U398 (N_398,N_296,N_153);
nand U399 (N_399,N_206,N_139);
and U400 (N_400,N_387,N_345);
and U401 (N_401,N_355,N_346);
and U402 (N_402,N_367,N_396);
xnor U403 (N_403,N_374,N_372);
xnor U404 (N_404,N_365,N_315);
nor U405 (N_405,N_389,N_373);
or U406 (N_406,N_301,N_302);
or U407 (N_407,N_384,N_340);
or U408 (N_408,N_344,N_349);
xnor U409 (N_409,N_379,N_341);
nand U410 (N_410,N_331,N_337);
nand U411 (N_411,N_332,N_390);
or U412 (N_412,N_324,N_378);
xor U413 (N_413,N_397,N_347);
nand U414 (N_414,N_392,N_317);
and U415 (N_415,N_391,N_307);
xnor U416 (N_416,N_358,N_382);
xor U417 (N_417,N_386,N_350);
and U418 (N_418,N_395,N_368);
nand U419 (N_419,N_359,N_383);
or U420 (N_420,N_353,N_325);
nand U421 (N_421,N_375,N_369);
or U422 (N_422,N_380,N_356);
xnor U423 (N_423,N_304,N_388);
and U424 (N_424,N_376,N_312);
and U425 (N_425,N_327,N_338);
xnor U426 (N_426,N_399,N_371);
and U427 (N_427,N_318,N_343);
or U428 (N_428,N_328,N_314);
or U429 (N_429,N_334,N_393);
nand U430 (N_430,N_330,N_352);
nand U431 (N_431,N_342,N_322);
or U432 (N_432,N_320,N_329);
or U433 (N_433,N_323,N_316);
nand U434 (N_434,N_363,N_310);
nor U435 (N_435,N_326,N_348);
and U436 (N_436,N_351,N_333);
and U437 (N_437,N_394,N_354);
nand U438 (N_438,N_357,N_305);
and U439 (N_439,N_311,N_398);
xnor U440 (N_440,N_385,N_309);
xor U441 (N_441,N_364,N_306);
and U442 (N_442,N_366,N_370);
and U443 (N_443,N_362,N_321);
xnor U444 (N_444,N_303,N_361);
nor U445 (N_445,N_381,N_313);
nand U446 (N_446,N_339,N_360);
nand U447 (N_447,N_336,N_319);
xor U448 (N_448,N_300,N_335);
or U449 (N_449,N_377,N_308);
nor U450 (N_450,N_344,N_300);
or U451 (N_451,N_366,N_332);
and U452 (N_452,N_316,N_382);
nor U453 (N_453,N_387,N_358);
or U454 (N_454,N_337,N_352);
and U455 (N_455,N_361,N_352);
xnor U456 (N_456,N_360,N_304);
nand U457 (N_457,N_342,N_357);
nor U458 (N_458,N_355,N_327);
or U459 (N_459,N_338,N_320);
nor U460 (N_460,N_334,N_379);
nor U461 (N_461,N_387,N_385);
or U462 (N_462,N_398,N_387);
nor U463 (N_463,N_393,N_315);
and U464 (N_464,N_356,N_378);
nand U465 (N_465,N_322,N_313);
xor U466 (N_466,N_356,N_343);
nor U467 (N_467,N_389,N_333);
nand U468 (N_468,N_369,N_323);
nand U469 (N_469,N_398,N_368);
or U470 (N_470,N_365,N_339);
xnor U471 (N_471,N_396,N_363);
nand U472 (N_472,N_377,N_358);
or U473 (N_473,N_308,N_301);
nand U474 (N_474,N_351,N_387);
and U475 (N_475,N_321,N_328);
nor U476 (N_476,N_368,N_370);
or U477 (N_477,N_373,N_357);
and U478 (N_478,N_310,N_371);
nand U479 (N_479,N_300,N_394);
and U480 (N_480,N_332,N_371);
nor U481 (N_481,N_336,N_330);
nand U482 (N_482,N_381,N_375);
xnor U483 (N_483,N_387,N_367);
and U484 (N_484,N_344,N_372);
nand U485 (N_485,N_369,N_388);
nand U486 (N_486,N_344,N_395);
xor U487 (N_487,N_392,N_322);
or U488 (N_488,N_399,N_330);
or U489 (N_489,N_321,N_336);
or U490 (N_490,N_325,N_301);
and U491 (N_491,N_307,N_332);
or U492 (N_492,N_348,N_301);
nor U493 (N_493,N_302,N_319);
and U494 (N_494,N_318,N_372);
and U495 (N_495,N_354,N_321);
nor U496 (N_496,N_304,N_340);
and U497 (N_497,N_313,N_356);
and U498 (N_498,N_384,N_373);
and U499 (N_499,N_381,N_333);
nand U500 (N_500,N_473,N_494);
nand U501 (N_501,N_406,N_420);
nand U502 (N_502,N_447,N_402);
xor U503 (N_503,N_476,N_481);
nor U504 (N_504,N_443,N_444);
or U505 (N_505,N_489,N_449);
xor U506 (N_506,N_429,N_432);
nor U507 (N_507,N_487,N_475);
nand U508 (N_508,N_416,N_472);
nor U509 (N_509,N_462,N_461);
or U510 (N_510,N_497,N_404);
and U511 (N_511,N_435,N_423);
nor U512 (N_512,N_468,N_496);
nor U513 (N_513,N_457,N_438);
or U514 (N_514,N_433,N_418);
or U515 (N_515,N_426,N_466);
xor U516 (N_516,N_456,N_480);
xnor U517 (N_517,N_460,N_439);
and U518 (N_518,N_408,N_440);
nand U519 (N_519,N_446,N_464);
or U520 (N_520,N_492,N_483);
xnor U521 (N_521,N_415,N_422);
or U522 (N_522,N_458,N_430);
nand U523 (N_523,N_488,N_465);
nand U524 (N_524,N_427,N_482);
nor U525 (N_525,N_486,N_431);
or U526 (N_526,N_436,N_428);
or U527 (N_527,N_453,N_441);
nand U528 (N_528,N_407,N_467);
xor U529 (N_529,N_417,N_490);
and U530 (N_530,N_412,N_401);
and U531 (N_531,N_493,N_442);
nand U532 (N_532,N_491,N_484);
or U533 (N_533,N_424,N_445);
and U534 (N_534,N_463,N_437);
xor U535 (N_535,N_495,N_474);
xnor U536 (N_536,N_411,N_409);
and U537 (N_537,N_454,N_452);
and U538 (N_538,N_485,N_499);
or U539 (N_539,N_459,N_450);
nor U540 (N_540,N_414,N_403);
and U541 (N_541,N_470,N_448);
nand U542 (N_542,N_425,N_405);
xnor U543 (N_543,N_419,N_479);
nand U544 (N_544,N_410,N_498);
and U545 (N_545,N_455,N_434);
or U546 (N_546,N_471,N_451);
xor U547 (N_547,N_478,N_413);
or U548 (N_548,N_477,N_469);
or U549 (N_549,N_421,N_400);
xor U550 (N_550,N_417,N_489);
and U551 (N_551,N_492,N_491);
and U552 (N_552,N_464,N_487);
and U553 (N_553,N_427,N_464);
nor U554 (N_554,N_470,N_456);
xnor U555 (N_555,N_411,N_485);
or U556 (N_556,N_421,N_417);
and U557 (N_557,N_408,N_495);
and U558 (N_558,N_439,N_496);
xor U559 (N_559,N_415,N_409);
nand U560 (N_560,N_443,N_491);
nor U561 (N_561,N_478,N_457);
xnor U562 (N_562,N_477,N_499);
nor U563 (N_563,N_457,N_435);
nand U564 (N_564,N_472,N_424);
nor U565 (N_565,N_499,N_439);
and U566 (N_566,N_428,N_491);
nor U567 (N_567,N_424,N_449);
nand U568 (N_568,N_402,N_407);
nor U569 (N_569,N_411,N_473);
xnor U570 (N_570,N_415,N_446);
and U571 (N_571,N_454,N_446);
or U572 (N_572,N_437,N_486);
nor U573 (N_573,N_446,N_401);
xnor U574 (N_574,N_409,N_433);
and U575 (N_575,N_477,N_450);
xnor U576 (N_576,N_448,N_428);
nor U577 (N_577,N_477,N_489);
xor U578 (N_578,N_468,N_431);
xnor U579 (N_579,N_484,N_430);
xor U580 (N_580,N_491,N_458);
and U581 (N_581,N_430,N_436);
nor U582 (N_582,N_472,N_464);
xor U583 (N_583,N_427,N_445);
nand U584 (N_584,N_482,N_498);
xor U585 (N_585,N_428,N_447);
nor U586 (N_586,N_415,N_474);
nor U587 (N_587,N_460,N_403);
nor U588 (N_588,N_469,N_484);
xor U589 (N_589,N_429,N_493);
and U590 (N_590,N_402,N_473);
nor U591 (N_591,N_425,N_484);
xor U592 (N_592,N_455,N_478);
or U593 (N_593,N_435,N_407);
nor U594 (N_594,N_464,N_430);
nand U595 (N_595,N_485,N_473);
nand U596 (N_596,N_469,N_444);
or U597 (N_597,N_454,N_464);
or U598 (N_598,N_429,N_450);
nand U599 (N_599,N_421,N_442);
nor U600 (N_600,N_506,N_592);
nand U601 (N_601,N_585,N_507);
or U602 (N_602,N_505,N_503);
xor U603 (N_603,N_501,N_558);
and U604 (N_604,N_575,N_533);
xor U605 (N_605,N_566,N_532);
nor U606 (N_606,N_510,N_567);
nand U607 (N_607,N_526,N_598);
nand U608 (N_608,N_548,N_513);
and U609 (N_609,N_564,N_595);
and U610 (N_610,N_597,N_518);
and U611 (N_611,N_508,N_552);
xnor U612 (N_612,N_569,N_563);
nor U613 (N_613,N_584,N_500);
nand U614 (N_614,N_511,N_524);
or U615 (N_615,N_562,N_588);
nand U616 (N_616,N_516,N_568);
and U617 (N_617,N_529,N_547);
nor U618 (N_618,N_554,N_539);
and U619 (N_619,N_556,N_594);
xor U620 (N_620,N_538,N_545);
nand U621 (N_621,N_519,N_561);
and U622 (N_622,N_504,N_530);
xnor U623 (N_623,N_573,N_576);
and U624 (N_624,N_502,N_535);
nand U625 (N_625,N_596,N_591);
or U626 (N_626,N_583,N_525);
xnor U627 (N_627,N_514,N_599);
nand U628 (N_628,N_559,N_590);
or U629 (N_629,N_580,N_565);
or U630 (N_630,N_572,N_586);
xor U631 (N_631,N_549,N_541);
nand U632 (N_632,N_557,N_523);
and U633 (N_633,N_536,N_550);
nor U634 (N_634,N_579,N_582);
or U635 (N_635,N_542,N_521);
and U636 (N_636,N_560,N_522);
nor U637 (N_637,N_543,N_534);
and U638 (N_638,N_589,N_528);
nand U639 (N_639,N_544,N_509);
nor U640 (N_640,N_577,N_571);
nor U641 (N_641,N_578,N_537);
and U642 (N_642,N_546,N_570);
nand U643 (N_643,N_520,N_540);
xor U644 (N_644,N_551,N_587);
nor U645 (N_645,N_593,N_517);
and U646 (N_646,N_512,N_515);
nor U647 (N_647,N_527,N_574);
or U648 (N_648,N_531,N_555);
nor U649 (N_649,N_581,N_553);
nand U650 (N_650,N_525,N_556);
xnor U651 (N_651,N_576,N_510);
nand U652 (N_652,N_559,N_518);
and U653 (N_653,N_548,N_585);
or U654 (N_654,N_584,N_582);
nand U655 (N_655,N_529,N_512);
and U656 (N_656,N_568,N_523);
xor U657 (N_657,N_580,N_525);
and U658 (N_658,N_530,N_587);
xor U659 (N_659,N_574,N_553);
or U660 (N_660,N_594,N_585);
nand U661 (N_661,N_513,N_545);
and U662 (N_662,N_576,N_505);
nor U663 (N_663,N_539,N_524);
and U664 (N_664,N_525,N_529);
and U665 (N_665,N_502,N_506);
and U666 (N_666,N_512,N_534);
nor U667 (N_667,N_538,N_511);
nand U668 (N_668,N_548,N_506);
or U669 (N_669,N_576,N_569);
or U670 (N_670,N_586,N_517);
nand U671 (N_671,N_531,N_582);
nor U672 (N_672,N_538,N_591);
and U673 (N_673,N_599,N_525);
nand U674 (N_674,N_553,N_554);
or U675 (N_675,N_580,N_596);
nand U676 (N_676,N_505,N_565);
nand U677 (N_677,N_553,N_538);
nand U678 (N_678,N_536,N_565);
xor U679 (N_679,N_549,N_551);
and U680 (N_680,N_580,N_570);
xor U681 (N_681,N_525,N_595);
nand U682 (N_682,N_578,N_584);
xor U683 (N_683,N_505,N_567);
nand U684 (N_684,N_599,N_590);
or U685 (N_685,N_547,N_510);
nor U686 (N_686,N_509,N_555);
nand U687 (N_687,N_516,N_555);
or U688 (N_688,N_564,N_562);
and U689 (N_689,N_571,N_553);
nor U690 (N_690,N_555,N_580);
nor U691 (N_691,N_526,N_571);
and U692 (N_692,N_510,N_514);
nor U693 (N_693,N_599,N_534);
and U694 (N_694,N_589,N_559);
nor U695 (N_695,N_572,N_512);
nand U696 (N_696,N_561,N_554);
or U697 (N_697,N_598,N_596);
nand U698 (N_698,N_523,N_594);
nand U699 (N_699,N_560,N_504);
or U700 (N_700,N_637,N_679);
or U701 (N_701,N_638,N_675);
or U702 (N_702,N_663,N_694);
and U703 (N_703,N_645,N_658);
and U704 (N_704,N_633,N_695);
nor U705 (N_705,N_652,N_636);
xor U706 (N_706,N_676,N_626);
nor U707 (N_707,N_672,N_641);
or U708 (N_708,N_691,N_610);
xnor U709 (N_709,N_603,N_648);
xnor U710 (N_710,N_609,N_662);
nor U711 (N_711,N_602,N_696);
and U712 (N_712,N_689,N_659);
xor U713 (N_713,N_688,N_680);
nand U714 (N_714,N_670,N_622);
xor U715 (N_715,N_692,N_605);
nor U716 (N_716,N_617,N_686);
and U717 (N_717,N_608,N_625);
nor U718 (N_718,N_621,N_671);
nand U719 (N_719,N_650,N_600);
and U720 (N_720,N_668,N_601);
or U721 (N_721,N_643,N_655);
nand U722 (N_722,N_674,N_697);
nor U723 (N_723,N_660,N_635);
or U724 (N_724,N_644,N_634);
and U725 (N_725,N_604,N_639);
nand U726 (N_726,N_654,N_656);
and U727 (N_727,N_677,N_651);
or U728 (N_728,N_619,N_653);
or U729 (N_729,N_630,N_607);
nand U730 (N_730,N_665,N_646);
and U731 (N_731,N_669,N_693);
xor U732 (N_732,N_690,N_627);
and U733 (N_733,N_684,N_682);
xnor U734 (N_734,N_657,N_647);
or U735 (N_735,N_661,N_624);
xor U736 (N_736,N_642,N_664);
xor U737 (N_737,N_616,N_698);
xor U738 (N_738,N_631,N_667);
xnor U739 (N_739,N_649,N_673);
nor U740 (N_740,N_615,N_623);
nor U741 (N_741,N_611,N_632);
xor U742 (N_742,N_683,N_606);
nor U743 (N_743,N_613,N_666);
xnor U744 (N_744,N_640,N_699);
nor U745 (N_745,N_678,N_620);
or U746 (N_746,N_685,N_681);
nor U747 (N_747,N_629,N_628);
nor U748 (N_748,N_618,N_614);
nand U749 (N_749,N_687,N_612);
nor U750 (N_750,N_652,N_612);
or U751 (N_751,N_625,N_670);
and U752 (N_752,N_623,N_653);
nor U753 (N_753,N_608,N_684);
xor U754 (N_754,N_624,N_665);
nand U755 (N_755,N_635,N_621);
nor U756 (N_756,N_616,N_682);
xnor U757 (N_757,N_606,N_607);
and U758 (N_758,N_683,N_637);
or U759 (N_759,N_607,N_657);
xnor U760 (N_760,N_661,N_696);
or U761 (N_761,N_674,N_677);
nor U762 (N_762,N_644,N_639);
xnor U763 (N_763,N_675,N_604);
xor U764 (N_764,N_659,N_688);
nand U765 (N_765,N_680,N_687);
xnor U766 (N_766,N_601,N_655);
or U767 (N_767,N_657,N_677);
nand U768 (N_768,N_684,N_645);
xor U769 (N_769,N_681,N_693);
and U770 (N_770,N_624,N_663);
xnor U771 (N_771,N_631,N_666);
or U772 (N_772,N_630,N_689);
xnor U773 (N_773,N_694,N_624);
or U774 (N_774,N_665,N_668);
nor U775 (N_775,N_681,N_664);
and U776 (N_776,N_686,N_688);
xnor U777 (N_777,N_635,N_658);
xnor U778 (N_778,N_640,N_601);
nor U779 (N_779,N_601,N_693);
xnor U780 (N_780,N_647,N_694);
nand U781 (N_781,N_640,N_631);
xor U782 (N_782,N_692,N_606);
and U783 (N_783,N_659,N_684);
and U784 (N_784,N_616,N_693);
nand U785 (N_785,N_688,N_663);
nand U786 (N_786,N_694,N_695);
xor U787 (N_787,N_632,N_621);
and U788 (N_788,N_697,N_685);
nor U789 (N_789,N_661,N_649);
nor U790 (N_790,N_620,N_677);
or U791 (N_791,N_695,N_624);
xnor U792 (N_792,N_648,N_635);
nand U793 (N_793,N_603,N_658);
and U794 (N_794,N_622,N_679);
nor U795 (N_795,N_622,N_619);
and U796 (N_796,N_681,N_616);
nor U797 (N_797,N_697,N_613);
or U798 (N_798,N_657,N_686);
and U799 (N_799,N_644,N_671);
nand U800 (N_800,N_701,N_738);
nor U801 (N_801,N_743,N_797);
and U802 (N_802,N_722,N_741);
nor U803 (N_803,N_746,N_771);
nand U804 (N_804,N_798,N_726);
xnor U805 (N_805,N_791,N_788);
nor U806 (N_806,N_734,N_703);
nand U807 (N_807,N_761,N_710);
or U808 (N_808,N_702,N_728);
xor U809 (N_809,N_778,N_744);
or U810 (N_810,N_708,N_795);
or U811 (N_811,N_760,N_775);
and U812 (N_812,N_794,N_732);
nand U813 (N_813,N_768,N_712);
or U814 (N_814,N_745,N_709);
and U815 (N_815,N_749,N_756);
nor U816 (N_816,N_792,N_776);
nor U817 (N_817,N_777,N_765);
xnor U818 (N_818,N_714,N_796);
xnor U819 (N_819,N_721,N_713);
nor U820 (N_820,N_707,N_784);
nor U821 (N_821,N_757,N_758);
nor U822 (N_822,N_705,N_782);
xnor U823 (N_823,N_737,N_731);
and U824 (N_824,N_729,N_717);
xor U825 (N_825,N_720,N_766);
xor U826 (N_826,N_735,N_785);
nor U827 (N_827,N_762,N_753);
or U828 (N_828,N_793,N_774);
nor U829 (N_829,N_719,N_790);
nand U830 (N_830,N_723,N_715);
nor U831 (N_831,N_770,N_724);
xnor U832 (N_832,N_740,N_711);
nand U833 (N_833,N_751,N_763);
or U834 (N_834,N_773,N_779);
or U835 (N_835,N_750,N_727);
or U836 (N_836,N_739,N_789);
xor U837 (N_837,N_725,N_718);
xor U838 (N_838,N_767,N_706);
and U839 (N_839,N_704,N_759);
and U840 (N_840,N_730,N_772);
nor U841 (N_841,N_781,N_769);
or U842 (N_842,N_783,N_755);
xor U843 (N_843,N_780,N_787);
nor U844 (N_844,N_752,N_700);
nor U845 (N_845,N_764,N_754);
nand U846 (N_846,N_736,N_786);
xor U847 (N_847,N_799,N_742);
nor U848 (N_848,N_733,N_716);
nor U849 (N_849,N_747,N_748);
and U850 (N_850,N_790,N_727);
and U851 (N_851,N_727,N_712);
and U852 (N_852,N_729,N_700);
nor U853 (N_853,N_789,N_705);
xor U854 (N_854,N_715,N_713);
or U855 (N_855,N_792,N_728);
or U856 (N_856,N_722,N_702);
or U857 (N_857,N_750,N_703);
and U858 (N_858,N_792,N_734);
or U859 (N_859,N_737,N_727);
xor U860 (N_860,N_702,N_720);
or U861 (N_861,N_752,N_787);
xor U862 (N_862,N_732,N_703);
xor U863 (N_863,N_734,N_708);
nor U864 (N_864,N_724,N_799);
nand U865 (N_865,N_792,N_756);
and U866 (N_866,N_711,N_793);
nand U867 (N_867,N_792,N_738);
or U868 (N_868,N_798,N_730);
or U869 (N_869,N_757,N_766);
and U870 (N_870,N_731,N_708);
nand U871 (N_871,N_723,N_756);
nand U872 (N_872,N_701,N_781);
or U873 (N_873,N_788,N_792);
nor U874 (N_874,N_782,N_766);
nor U875 (N_875,N_741,N_736);
xnor U876 (N_876,N_769,N_734);
and U877 (N_877,N_785,N_720);
and U878 (N_878,N_758,N_760);
nand U879 (N_879,N_793,N_754);
nor U880 (N_880,N_763,N_703);
and U881 (N_881,N_733,N_793);
xor U882 (N_882,N_752,N_781);
and U883 (N_883,N_749,N_722);
and U884 (N_884,N_710,N_705);
nand U885 (N_885,N_765,N_768);
nor U886 (N_886,N_759,N_736);
nand U887 (N_887,N_757,N_726);
or U888 (N_888,N_711,N_784);
nor U889 (N_889,N_706,N_780);
or U890 (N_890,N_740,N_781);
xor U891 (N_891,N_717,N_741);
nand U892 (N_892,N_741,N_732);
and U893 (N_893,N_763,N_752);
nor U894 (N_894,N_706,N_778);
nor U895 (N_895,N_751,N_705);
nand U896 (N_896,N_703,N_719);
and U897 (N_897,N_745,N_704);
nor U898 (N_898,N_777,N_773);
or U899 (N_899,N_740,N_761);
nand U900 (N_900,N_888,N_805);
xnor U901 (N_901,N_831,N_814);
nand U902 (N_902,N_873,N_898);
xor U903 (N_903,N_891,N_865);
nor U904 (N_904,N_877,N_866);
and U905 (N_905,N_813,N_846);
xor U906 (N_906,N_840,N_867);
nand U907 (N_907,N_882,N_848);
nand U908 (N_908,N_836,N_801);
and U909 (N_909,N_857,N_828);
nand U910 (N_910,N_842,N_810);
xor U911 (N_911,N_817,N_897);
and U912 (N_912,N_870,N_802);
xor U913 (N_913,N_824,N_821);
or U914 (N_914,N_869,N_851);
xor U915 (N_915,N_880,N_886);
nor U916 (N_916,N_800,N_809);
nor U917 (N_917,N_838,N_825);
nand U918 (N_918,N_843,N_826);
nand U919 (N_919,N_875,N_890);
nor U920 (N_920,N_849,N_823);
nor U921 (N_921,N_896,N_859);
nor U922 (N_922,N_899,N_804);
nor U923 (N_923,N_858,N_894);
nor U924 (N_924,N_820,N_807);
nor U925 (N_925,N_860,N_874);
nand U926 (N_926,N_887,N_893);
or U927 (N_927,N_806,N_883);
nor U928 (N_928,N_863,N_829);
nor U929 (N_929,N_879,N_856);
and U930 (N_930,N_853,N_811);
or U931 (N_931,N_839,N_847);
and U932 (N_932,N_868,N_832);
nor U933 (N_933,N_889,N_812);
xnor U934 (N_934,N_895,N_884);
or U935 (N_935,N_881,N_871);
and U936 (N_936,N_885,N_864);
nor U937 (N_937,N_852,N_815);
nor U938 (N_938,N_872,N_854);
nand U939 (N_939,N_878,N_862);
nand U940 (N_940,N_855,N_861);
nand U941 (N_941,N_850,N_892);
xor U942 (N_942,N_827,N_833);
nand U943 (N_943,N_830,N_822);
nor U944 (N_944,N_816,N_835);
nand U945 (N_945,N_841,N_803);
nand U946 (N_946,N_845,N_876);
or U947 (N_947,N_837,N_834);
and U948 (N_948,N_818,N_808);
and U949 (N_949,N_819,N_844);
nand U950 (N_950,N_843,N_810);
nor U951 (N_951,N_886,N_878);
xnor U952 (N_952,N_878,N_871);
xor U953 (N_953,N_858,N_842);
nand U954 (N_954,N_829,N_861);
or U955 (N_955,N_843,N_836);
nor U956 (N_956,N_872,N_887);
nor U957 (N_957,N_880,N_814);
or U958 (N_958,N_808,N_850);
nor U959 (N_959,N_868,N_882);
nor U960 (N_960,N_812,N_819);
or U961 (N_961,N_828,N_814);
nand U962 (N_962,N_813,N_862);
or U963 (N_963,N_880,N_894);
or U964 (N_964,N_882,N_843);
or U965 (N_965,N_873,N_882);
or U966 (N_966,N_882,N_811);
nand U967 (N_967,N_879,N_840);
or U968 (N_968,N_814,N_889);
nand U969 (N_969,N_886,N_879);
xor U970 (N_970,N_852,N_835);
nand U971 (N_971,N_853,N_867);
nor U972 (N_972,N_818,N_893);
xnor U973 (N_973,N_876,N_818);
nand U974 (N_974,N_842,N_880);
nor U975 (N_975,N_896,N_885);
or U976 (N_976,N_897,N_843);
nand U977 (N_977,N_849,N_830);
xor U978 (N_978,N_889,N_869);
nand U979 (N_979,N_889,N_893);
or U980 (N_980,N_854,N_874);
xnor U981 (N_981,N_813,N_844);
nand U982 (N_982,N_891,N_835);
and U983 (N_983,N_858,N_881);
or U984 (N_984,N_822,N_876);
or U985 (N_985,N_848,N_872);
or U986 (N_986,N_809,N_872);
nand U987 (N_987,N_874,N_836);
nor U988 (N_988,N_811,N_885);
and U989 (N_989,N_866,N_850);
nand U990 (N_990,N_867,N_897);
and U991 (N_991,N_807,N_895);
nor U992 (N_992,N_829,N_899);
and U993 (N_993,N_865,N_837);
or U994 (N_994,N_817,N_808);
nand U995 (N_995,N_807,N_812);
xor U996 (N_996,N_853,N_817);
and U997 (N_997,N_833,N_881);
or U998 (N_998,N_846,N_886);
nor U999 (N_999,N_887,N_861);
xnor U1000 (N_1000,N_912,N_941);
xnor U1001 (N_1001,N_942,N_931);
or U1002 (N_1002,N_921,N_940);
nand U1003 (N_1003,N_967,N_966);
nand U1004 (N_1004,N_968,N_916);
and U1005 (N_1005,N_969,N_907);
or U1006 (N_1006,N_996,N_913);
and U1007 (N_1007,N_908,N_918);
or U1008 (N_1008,N_985,N_989);
or U1009 (N_1009,N_959,N_994);
nand U1010 (N_1010,N_998,N_932);
nand U1011 (N_1011,N_934,N_999);
and U1012 (N_1012,N_950,N_992);
nand U1013 (N_1013,N_903,N_958);
xnor U1014 (N_1014,N_963,N_919);
xor U1015 (N_1015,N_964,N_970);
nand U1016 (N_1016,N_984,N_917);
and U1017 (N_1017,N_957,N_925);
nor U1018 (N_1018,N_981,N_955);
nand U1019 (N_1019,N_930,N_920);
nand U1020 (N_1020,N_926,N_929);
xor U1021 (N_1021,N_924,N_904);
xnor U1022 (N_1022,N_906,N_988);
nor U1023 (N_1023,N_923,N_972);
nand U1024 (N_1024,N_922,N_995);
nand U1025 (N_1025,N_953,N_976);
nand U1026 (N_1026,N_978,N_944);
and U1027 (N_1027,N_935,N_997);
nand U1028 (N_1028,N_951,N_952);
nor U1029 (N_1029,N_915,N_943);
nand U1030 (N_1030,N_901,N_991);
and U1031 (N_1031,N_977,N_945);
xnor U1032 (N_1032,N_948,N_911);
and U1033 (N_1033,N_983,N_937);
and U1034 (N_1034,N_949,N_982);
and U1035 (N_1035,N_936,N_914);
nand U1036 (N_1036,N_905,N_960);
or U1037 (N_1037,N_962,N_979);
nand U1038 (N_1038,N_965,N_954);
and U1039 (N_1039,N_902,N_980);
and U1040 (N_1040,N_909,N_928);
and U1041 (N_1041,N_974,N_993);
xor U1042 (N_1042,N_947,N_971);
and U1043 (N_1043,N_939,N_938);
nor U1044 (N_1044,N_910,N_927);
xor U1045 (N_1045,N_990,N_987);
nand U1046 (N_1046,N_961,N_975);
xnor U1047 (N_1047,N_956,N_986);
nor U1048 (N_1048,N_946,N_933);
nand U1049 (N_1049,N_900,N_973);
or U1050 (N_1050,N_915,N_933);
or U1051 (N_1051,N_943,N_905);
or U1052 (N_1052,N_903,N_933);
or U1053 (N_1053,N_977,N_920);
or U1054 (N_1054,N_961,N_909);
nor U1055 (N_1055,N_953,N_929);
xor U1056 (N_1056,N_947,N_902);
and U1057 (N_1057,N_986,N_929);
and U1058 (N_1058,N_918,N_931);
and U1059 (N_1059,N_945,N_967);
nand U1060 (N_1060,N_978,N_909);
nand U1061 (N_1061,N_910,N_917);
and U1062 (N_1062,N_956,N_920);
nand U1063 (N_1063,N_955,N_972);
and U1064 (N_1064,N_936,N_989);
or U1065 (N_1065,N_940,N_954);
nand U1066 (N_1066,N_917,N_993);
xor U1067 (N_1067,N_967,N_935);
nand U1068 (N_1068,N_916,N_926);
and U1069 (N_1069,N_955,N_922);
nand U1070 (N_1070,N_965,N_973);
xnor U1071 (N_1071,N_973,N_915);
or U1072 (N_1072,N_950,N_967);
xor U1073 (N_1073,N_909,N_921);
nor U1074 (N_1074,N_942,N_982);
or U1075 (N_1075,N_929,N_903);
or U1076 (N_1076,N_919,N_941);
xor U1077 (N_1077,N_957,N_948);
xnor U1078 (N_1078,N_996,N_911);
xor U1079 (N_1079,N_999,N_931);
and U1080 (N_1080,N_983,N_966);
nand U1081 (N_1081,N_935,N_927);
and U1082 (N_1082,N_967,N_925);
nand U1083 (N_1083,N_991,N_928);
and U1084 (N_1084,N_945,N_947);
nor U1085 (N_1085,N_984,N_926);
or U1086 (N_1086,N_954,N_910);
or U1087 (N_1087,N_982,N_970);
nand U1088 (N_1088,N_939,N_902);
or U1089 (N_1089,N_988,N_917);
nand U1090 (N_1090,N_917,N_974);
or U1091 (N_1091,N_986,N_907);
and U1092 (N_1092,N_984,N_910);
and U1093 (N_1093,N_947,N_954);
nand U1094 (N_1094,N_914,N_939);
or U1095 (N_1095,N_979,N_901);
nand U1096 (N_1096,N_941,N_937);
or U1097 (N_1097,N_965,N_950);
xor U1098 (N_1098,N_987,N_909);
nand U1099 (N_1099,N_953,N_930);
and U1100 (N_1100,N_1095,N_1048);
xnor U1101 (N_1101,N_1046,N_1069);
nor U1102 (N_1102,N_1006,N_1093);
or U1103 (N_1103,N_1049,N_1027);
or U1104 (N_1104,N_1003,N_1087);
nand U1105 (N_1105,N_1081,N_1089);
and U1106 (N_1106,N_1033,N_1067);
xor U1107 (N_1107,N_1007,N_1038);
xor U1108 (N_1108,N_1013,N_1073);
or U1109 (N_1109,N_1000,N_1051);
nand U1110 (N_1110,N_1011,N_1024);
nor U1111 (N_1111,N_1017,N_1078);
nor U1112 (N_1112,N_1020,N_1012);
xor U1113 (N_1113,N_1061,N_1099);
or U1114 (N_1114,N_1008,N_1056);
xnor U1115 (N_1115,N_1097,N_1077);
xnor U1116 (N_1116,N_1045,N_1018);
nor U1117 (N_1117,N_1086,N_1080);
and U1118 (N_1118,N_1055,N_1092);
xor U1119 (N_1119,N_1005,N_1062);
nand U1120 (N_1120,N_1009,N_1064);
nor U1121 (N_1121,N_1019,N_1029);
nor U1122 (N_1122,N_1026,N_1032);
nand U1123 (N_1123,N_1053,N_1010);
xor U1124 (N_1124,N_1060,N_1035);
and U1125 (N_1125,N_1098,N_1057);
nand U1126 (N_1126,N_1025,N_1030);
nor U1127 (N_1127,N_1052,N_1075);
nor U1128 (N_1128,N_1058,N_1091);
xor U1129 (N_1129,N_1050,N_1063);
xor U1130 (N_1130,N_1059,N_1039);
and U1131 (N_1131,N_1066,N_1088);
xor U1132 (N_1132,N_1028,N_1014);
nor U1133 (N_1133,N_1044,N_1036);
xnor U1134 (N_1134,N_1083,N_1074);
nand U1135 (N_1135,N_1001,N_1047);
nand U1136 (N_1136,N_1082,N_1023);
nand U1137 (N_1137,N_1085,N_1076);
nor U1138 (N_1138,N_1070,N_1004);
or U1139 (N_1139,N_1072,N_1054);
nand U1140 (N_1140,N_1068,N_1037);
or U1141 (N_1141,N_1016,N_1065);
nand U1142 (N_1142,N_1042,N_1031);
and U1143 (N_1143,N_1090,N_1043);
nor U1144 (N_1144,N_1071,N_1079);
nand U1145 (N_1145,N_1022,N_1034);
xnor U1146 (N_1146,N_1041,N_1002);
nand U1147 (N_1147,N_1015,N_1021);
nor U1148 (N_1148,N_1096,N_1094);
or U1149 (N_1149,N_1084,N_1040);
xnor U1150 (N_1150,N_1031,N_1080);
and U1151 (N_1151,N_1088,N_1016);
and U1152 (N_1152,N_1054,N_1075);
or U1153 (N_1153,N_1080,N_1001);
or U1154 (N_1154,N_1073,N_1041);
nor U1155 (N_1155,N_1019,N_1031);
xnor U1156 (N_1156,N_1071,N_1096);
or U1157 (N_1157,N_1000,N_1037);
xor U1158 (N_1158,N_1093,N_1099);
nand U1159 (N_1159,N_1071,N_1091);
xnor U1160 (N_1160,N_1095,N_1093);
nor U1161 (N_1161,N_1004,N_1095);
or U1162 (N_1162,N_1008,N_1066);
or U1163 (N_1163,N_1088,N_1017);
or U1164 (N_1164,N_1005,N_1075);
or U1165 (N_1165,N_1098,N_1021);
or U1166 (N_1166,N_1091,N_1036);
nor U1167 (N_1167,N_1096,N_1029);
nor U1168 (N_1168,N_1025,N_1084);
or U1169 (N_1169,N_1065,N_1047);
and U1170 (N_1170,N_1077,N_1013);
nor U1171 (N_1171,N_1053,N_1037);
nand U1172 (N_1172,N_1099,N_1015);
and U1173 (N_1173,N_1058,N_1008);
nor U1174 (N_1174,N_1027,N_1002);
nor U1175 (N_1175,N_1072,N_1095);
nor U1176 (N_1176,N_1027,N_1089);
and U1177 (N_1177,N_1096,N_1087);
nand U1178 (N_1178,N_1029,N_1050);
nand U1179 (N_1179,N_1063,N_1035);
and U1180 (N_1180,N_1024,N_1091);
nor U1181 (N_1181,N_1066,N_1072);
or U1182 (N_1182,N_1045,N_1042);
and U1183 (N_1183,N_1039,N_1049);
and U1184 (N_1184,N_1006,N_1095);
nand U1185 (N_1185,N_1056,N_1094);
nand U1186 (N_1186,N_1093,N_1098);
or U1187 (N_1187,N_1073,N_1014);
nand U1188 (N_1188,N_1064,N_1066);
and U1189 (N_1189,N_1072,N_1009);
nor U1190 (N_1190,N_1004,N_1024);
and U1191 (N_1191,N_1088,N_1000);
xor U1192 (N_1192,N_1091,N_1087);
nor U1193 (N_1193,N_1039,N_1053);
or U1194 (N_1194,N_1026,N_1006);
and U1195 (N_1195,N_1055,N_1058);
and U1196 (N_1196,N_1053,N_1059);
or U1197 (N_1197,N_1053,N_1049);
or U1198 (N_1198,N_1054,N_1035);
nor U1199 (N_1199,N_1032,N_1075);
xor U1200 (N_1200,N_1174,N_1190);
and U1201 (N_1201,N_1150,N_1193);
and U1202 (N_1202,N_1155,N_1153);
nand U1203 (N_1203,N_1123,N_1189);
or U1204 (N_1204,N_1101,N_1143);
or U1205 (N_1205,N_1148,N_1186);
and U1206 (N_1206,N_1184,N_1121);
nand U1207 (N_1207,N_1111,N_1118);
and U1208 (N_1208,N_1108,N_1199);
nor U1209 (N_1209,N_1178,N_1198);
xnor U1210 (N_1210,N_1149,N_1158);
nand U1211 (N_1211,N_1183,N_1115);
nor U1212 (N_1212,N_1191,N_1125);
nand U1213 (N_1213,N_1179,N_1120);
and U1214 (N_1214,N_1131,N_1133);
nand U1215 (N_1215,N_1154,N_1127);
nand U1216 (N_1216,N_1117,N_1100);
nor U1217 (N_1217,N_1156,N_1135);
nor U1218 (N_1218,N_1182,N_1170);
or U1219 (N_1219,N_1128,N_1107);
nor U1220 (N_1220,N_1173,N_1192);
nor U1221 (N_1221,N_1160,N_1163);
or U1222 (N_1222,N_1114,N_1171);
nor U1223 (N_1223,N_1188,N_1110);
xor U1224 (N_1224,N_1167,N_1161);
nand U1225 (N_1225,N_1136,N_1106);
nor U1226 (N_1226,N_1139,N_1176);
or U1227 (N_1227,N_1142,N_1146);
nor U1228 (N_1228,N_1109,N_1151);
and U1229 (N_1229,N_1165,N_1187);
or U1230 (N_1230,N_1104,N_1113);
and U1231 (N_1231,N_1175,N_1137);
or U1232 (N_1232,N_1129,N_1138);
and U1233 (N_1233,N_1196,N_1147);
or U1234 (N_1234,N_1194,N_1119);
nor U1235 (N_1235,N_1124,N_1102);
nor U1236 (N_1236,N_1144,N_1162);
xor U1237 (N_1237,N_1181,N_1112);
or U1238 (N_1238,N_1152,N_1122);
xnor U1239 (N_1239,N_1169,N_1197);
nor U1240 (N_1240,N_1105,N_1103);
and U1241 (N_1241,N_1172,N_1168);
nor U1242 (N_1242,N_1166,N_1185);
nand U1243 (N_1243,N_1177,N_1164);
nor U1244 (N_1244,N_1145,N_1116);
xnor U1245 (N_1245,N_1141,N_1195);
xor U1246 (N_1246,N_1157,N_1132);
and U1247 (N_1247,N_1180,N_1126);
or U1248 (N_1248,N_1159,N_1140);
nand U1249 (N_1249,N_1134,N_1130);
nand U1250 (N_1250,N_1184,N_1180);
and U1251 (N_1251,N_1199,N_1181);
xor U1252 (N_1252,N_1130,N_1152);
and U1253 (N_1253,N_1103,N_1144);
nand U1254 (N_1254,N_1166,N_1153);
xnor U1255 (N_1255,N_1134,N_1199);
or U1256 (N_1256,N_1126,N_1189);
nand U1257 (N_1257,N_1174,N_1109);
nor U1258 (N_1258,N_1146,N_1136);
and U1259 (N_1259,N_1143,N_1115);
nand U1260 (N_1260,N_1107,N_1115);
nor U1261 (N_1261,N_1149,N_1179);
xor U1262 (N_1262,N_1195,N_1108);
xor U1263 (N_1263,N_1185,N_1188);
and U1264 (N_1264,N_1127,N_1142);
xor U1265 (N_1265,N_1188,N_1160);
xor U1266 (N_1266,N_1165,N_1119);
or U1267 (N_1267,N_1141,N_1112);
xor U1268 (N_1268,N_1171,N_1151);
nand U1269 (N_1269,N_1180,N_1162);
and U1270 (N_1270,N_1177,N_1128);
and U1271 (N_1271,N_1196,N_1186);
or U1272 (N_1272,N_1114,N_1193);
xnor U1273 (N_1273,N_1139,N_1130);
xor U1274 (N_1274,N_1125,N_1151);
and U1275 (N_1275,N_1169,N_1135);
nor U1276 (N_1276,N_1182,N_1181);
xor U1277 (N_1277,N_1136,N_1126);
nor U1278 (N_1278,N_1199,N_1115);
xor U1279 (N_1279,N_1189,N_1168);
nor U1280 (N_1280,N_1102,N_1198);
or U1281 (N_1281,N_1118,N_1192);
xor U1282 (N_1282,N_1107,N_1172);
nor U1283 (N_1283,N_1118,N_1152);
nand U1284 (N_1284,N_1131,N_1166);
nor U1285 (N_1285,N_1183,N_1134);
or U1286 (N_1286,N_1170,N_1172);
and U1287 (N_1287,N_1197,N_1180);
nand U1288 (N_1288,N_1166,N_1172);
xor U1289 (N_1289,N_1104,N_1179);
xor U1290 (N_1290,N_1135,N_1109);
nand U1291 (N_1291,N_1109,N_1164);
xnor U1292 (N_1292,N_1138,N_1115);
or U1293 (N_1293,N_1176,N_1115);
and U1294 (N_1294,N_1110,N_1140);
and U1295 (N_1295,N_1173,N_1188);
and U1296 (N_1296,N_1140,N_1119);
and U1297 (N_1297,N_1117,N_1110);
nor U1298 (N_1298,N_1135,N_1115);
xor U1299 (N_1299,N_1141,N_1184);
nand U1300 (N_1300,N_1236,N_1272);
and U1301 (N_1301,N_1299,N_1264);
nor U1302 (N_1302,N_1221,N_1243);
xor U1303 (N_1303,N_1238,N_1275);
nor U1304 (N_1304,N_1234,N_1281);
or U1305 (N_1305,N_1290,N_1255);
nor U1306 (N_1306,N_1284,N_1267);
nand U1307 (N_1307,N_1223,N_1231);
or U1308 (N_1308,N_1293,N_1204);
nand U1309 (N_1309,N_1210,N_1273);
or U1310 (N_1310,N_1297,N_1282);
and U1311 (N_1311,N_1246,N_1277);
xor U1312 (N_1312,N_1205,N_1263);
and U1313 (N_1313,N_1237,N_1228);
nand U1314 (N_1314,N_1276,N_1295);
xnor U1315 (N_1315,N_1209,N_1203);
or U1316 (N_1316,N_1250,N_1292);
or U1317 (N_1317,N_1253,N_1240);
or U1318 (N_1318,N_1287,N_1283);
nand U1319 (N_1319,N_1259,N_1268);
xnor U1320 (N_1320,N_1206,N_1242);
xnor U1321 (N_1321,N_1251,N_1226);
or U1322 (N_1322,N_1212,N_1269);
nor U1323 (N_1323,N_1220,N_1211);
nand U1324 (N_1324,N_1245,N_1271);
nor U1325 (N_1325,N_1285,N_1254);
nor U1326 (N_1326,N_1215,N_1286);
xor U1327 (N_1327,N_1233,N_1288);
and U1328 (N_1328,N_1225,N_1218);
or U1329 (N_1329,N_1274,N_1232);
xnor U1330 (N_1330,N_1265,N_1280);
xor U1331 (N_1331,N_1270,N_1291);
or U1332 (N_1332,N_1229,N_1241);
nand U1333 (N_1333,N_1258,N_1266);
or U1334 (N_1334,N_1222,N_1260);
or U1335 (N_1335,N_1257,N_1296);
xnor U1336 (N_1336,N_1298,N_1249);
or U1337 (N_1337,N_1248,N_1217);
and U1338 (N_1338,N_1252,N_1262);
and U1339 (N_1339,N_1200,N_1247);
and U1340 (N_1340,N_1244,N_1256);
and U1341 (N_1341,N_1235,N_1261);
or U1342 (N_1342,N_1227,N_1294);
nand U1343 (N_1343,N_1201,N_1216);
or U1344 (N_1344,N_1289,N_1219);
xor U1345 (N_1345,N_1214,N_1279);
and U1346 (N_1346,N_1208,N_1207);
xor U1347 (N_1347,N_1224,N_1239);
nand U1348 (N_1348,N_1230,N_1202);
nand U1349 (N_1349,N_1278,N_1213);
nand U1350 (N_1350,N_1273,N_1209);
nand U1351 (N_1351,N_1227,N_1210);
and U1352 (N_1352,N_1297,N_1218);
and U1353 (N_1353,N_1277,N_1200);
and U1354 (N_1354,N_1281,N_1251);
nand U1355 (N_1355,N_1222,N_1256);
nand U1356 (N_1356,N_1264,N_1284);
xor U1357 (N_1357,N_1283,N_1262);
nor U1358 (N_1358,N_1279,N_1246);
xor U1359 (N_1359,N_1204,N_1266);
xnor U1360 (N_1360,N_1246,N_1269);
or U1361 (N_1361,N_1250,N_1277);
nor U1362 (N_1362,N_1231,N_1260);
xnor U1363 (N_1363,N_1213,N_1248);
or U1364 (N_1364,N_1280,N_1279);
xor U1365 (N_1365,N_1208,N_1289);
and U1366 (N_1366,N_1231,N_1253);
and U1367 (N_1367,N_1247,N_1249);
or U1368 (N_1368,N_1290,N_1206);
or U1369 (N_1369,N_1291,N_1263);
or U1370 (N_1370,N_1276,N_1218);
nand U1371 (N_1371,N_1253,N_1279);
xnor U1372 (N_1372,N_1272,N_1283);
nor U1373 (N_1373,N_1255,N_1292);
and U1374 (N_1374,N_1202,N_1291);
nor U1375 (N_1375,N_1291,N_1276);
nor U1376 (N_1376,N_1265,N_1229);
or U1377 (N_1377,N_1224,N_1259);
nor U1378 (N_1378,N_1226,N_1298);
nor U1379 (N_1379,N_1228,N_1247);
nand U1380 (N_1380,N_1210,N_1278);
xor U1381 (N_1381,N_1255,N_1241);
xor U1382 (N_1382,N_1234,N_1238);
nand U1383 (N_1383,N_1259,N_1247);
xor U1384 (N_1384,N_1221,N_1229);
xor U1385 (N_1385,N_1258,N_1220);
nand U1386 (N_1386,N_1237,N_1283);
and U1387 (N_1387,N_1229,N_1256);
nor U1388 (N_1388,N_1283,N_1208);
and U1389 (N_1389,N_1270,N_1257);
and U1390 (N_1390,N_1242,N_1207);
nand U1391 (N_1391,N_1238,N_1239);
nor U1392 (N_1392,N_1230,N_1247);
nand U1393 (N_1393,N_1204,N_1287);
xnor U1394 (N_1394,N_1295,N_1233);
and U1395 (N_1395,N_1216,N_1205);
nor U1396 (N_1396,N_1215,N_1221);
nand U1397 (N_1397,N_1244,N_1259);
or U1398 (N_1398,N_1278,N_1227);
nand U1399 (N_1399,N_1221,N_1281);
and U1400 (N_1400,N_1335,N_1339);
and U1401 (N_1401,N_1380,N_1390);
nor U1402 (N_1402,N_1372,N_1320);
xnor U1403 (N_1403,N_1316,N_1342);
nand U1404 (N_1404,N_1394,N_1389);
and U1405 (N_1405,N_1304,N_1350);
nor U1406 (N_1406,N_1351,N_1327);
nand U1407 (N_1407,N_1382,N_1319);
nor U1408 (N_1408,N_1318,N_1321);
nand U1409 (N_1409,N_1308,N_1363);
nor U1410 (N_1410,N_1313,N_1399);
nor U1411 (N_1411,N_1305,N_1395);
or U1412 (N_1412,N_1322,N_1386);
nor U1413 (N_1413,N_1328,N_1314);
nand U1414 (N_1414,N_1344,N_1310);
xor U1415 (N_1415,N_1326,N_1354);
nor U1416 (N_1416,N_1315,N_1329);
or U1417 (N_1417,N_1323,N_1355);
and U1418 (N_1418,N_1341,N_1365);
and U1419 (N_1419,N_1374,N_1309);
nand U1420 (N_1420,N_1387,N_1336);
or U1421 (N_1421,N_1303,N_1369);
or U1422 (N_1422,N_1384,N_1360);
nor U1423 (N_1423,N_1371,N_1357);
nor U1424 (N_1424,N_1337,N_1332);
and U1425 (N_1425,N_1343,N_1391);
nand U1426 (N_1426,N_1385,N_1333);
xnor U1427 (N_1427,N_1381,N_1334);
and U1428 (N_1428,N_1388,N_1368);
and U1429 (N_1429,N_1358,N_1311);
nand U1430 (N_1430,N_1373,N_1393);
and U1431 (N_1431,N_1392,N_1362);
nor U1432 (N_1432,N_1398,N_1325);
nor U1433 (N_1433,N_1396,N_1349);
or U1434 (N_1434,N_1300,N_1383);
nor U1435 (N_1435,N_1338,N_1306);
xor U1436 (N_1436,N_1378,N_1345);
nand U1437 (N_1437,N_1307,N_1347);
and U1438 (N_1438,N_1348,N_1352);
nor U1439 (N_1439,N_1359,N_1364);
or U1440 (N_1440,N_1377,N_1397);
nand U1441 (N_1441,N_1317,N_1324);
and U1442 (N_1442,N_1331,N_1367);
or U1443 (N_1443,N_1366,N_1330);
nor U1444 (N_1444,N_1356,N_1376);
and U1445 (N_1445,N_1370,N_1361);
xor U1446 (N_1446,N_1346,N_1353);
or U1447 (N_1447,N_1302,N_1340);
xor U1448 (N_1448,N_1375,N_1301);
nor U1449 (N_1449,N_1379,N_1312);
xnor U1450 (N_1450,N_1341,N_1398);
nand U1451 (N_1451,N_1371,N_1332);
or U1452 (N_1452,N_1348,N_1337);
or U1453 (N_1453,N_1331,N_1383);
and U1454 (N_1454,N_1357,N_1335);
xnor U1455 (N_1455,N_1373,N_1399);
nor U1456 (N_1456,N_1372,N_1392);
and U1457 (N_1457,N_1306,N_1337);
or U1458 (N_1458,N_1380,N_1360);
nand U1459 (N_1459,N_1375,N_1306);
or U1460 (N_1460,N_1326,N_1396);
or U1461 (N_1461,N_1397,N_1322);
or U1462 (N_1462,N_1328,N_1347);
nor U1463 (N_1463,N_1381,N_1325);
and U1464 (N_1464,N_1358,N_1357);
and U1465 (N_1465,N_1345,N_1399);
nand U1466 (N_1466,N_1355,N_1398);
xnor U1467 (N_1467,N_1335,N_1358);
or U1468 (N_1468,N_1318,N_1371);
xnor U1469 (N_1469,N_1335,N_1397);
nand U1470 (N_1470,N_1370,N_1319);
and U1471 (N_1471,N_1391,N_1305);
and U1472 (N_1472,N_1361,N_1303);
nor U1473 (N_1473,N_1363,N_1377);
nor U1474 (N_1474,N_1303,N_1353);
or U1475 (N_1475,N_1377,N_1331);
xnor U1476 (N_1476,N_1300,N_1382);
and U1477 (N_1477,N_1362,N_1329);
nor U1478 (N_1478,N_1314,N_1350);
nand U1479 (N_1479,N_1339,N_1367);
nor U1480 (N_1480,N_1378,N_1326);
nor U1481 (N_1481,N_1311,N_1347);
nor U1482 (N_1482,N_1331,N_1362);
and U1483 (N_1483,N_1378,N_1336);
nand U1484 (N_1484,N_1313,N_1343);
xor U1485 (N_1485,N_1351,N_1357);
or U1486 (N_1486,N_1318,N_1325);
xnor U1487 (N_1487,N_1399,N_1336);
and U1488 (N_1488,N_1301,N_1379);
nor U1489 (N_1489,N_1373,N_1377);
nand U1490 (N_1490,N_1316,N_1373);
and U1491 (N_1491,N_1321,N_1337);
nand U1492 (N_1492,N_1373,N_1313);
nand U1493 (N_1493,N_1361,N_1328);
and U1494 (N_1494,N_1385,N_1396);
nand U1495 (N_1495,N_1308,N_1336);
nor U1496 (N_1496,N_1378,N_1347);
or U1497 (N_1497,N_1352,N_1349);
nor U1498 (N_1498,N_1301,N_1346);
or U1499 (N_1499,N_1323,N_1344);
xor U1500 (N_1500,N_1436,N_1408);
nor U1501 (N_1501,N_1460,N_1446);
nor U1502 (N_1502,N_1493,N_1448);
xor U1503 (N_1503,N_1445,N_1440);
nand U1504 (N_1504,N_1427,N_1438);
or U1505 (N_1505,N_1443,N_1451);
and U1506 (N_1506,N_1498,N_1455);
nand U1507 (N_1507,N_1424,N_1491);
nor U1508 (N_1508,N_1441,N_1456);
nand U1509 (N_1509,N_1442,N_1494);
or U1510 (N_1510,N_1471,N_1492);
and U1511 (N_1511,N_1466,N_1458);
nor U1512 (N_1512,N_1417,N_1483);
or U1513 (N_1513,N_1422,N_1444);
and U1514 (N_1514,N_1468,N_1453);
nand U1515 (N_1515,N_1499,N_1418);
nand U1516 (N_1516,N_1426,N_1425);
xnor U1517 (N_1517,N_1409,N_1488);
xnor U1518 (N_1518,N_1497,N_1431);
xor U1519 (N_1519,N_1454,N_1472);
nand U1520 (N_1520,N_1421,N_1478);
or U1521 (N_1521,N_1481,N_1490);
nor U1522 (N_1522,N_1473,N_1439);
and U1523 (N_1523,N_1475,N_1415);
nor U1524 (N_1524,N_1428,N_1484);
nand U1525 (N_1525,N_1467,N_1405);
xnor U1526 (N_1526,N_1462,N_1470);
nor U1527 (N_1527,N_1450,N_1433);
and U1528 (N_1528,N_1452,N_1435);
xor U1529 (N_1529,N_1465,N_1486);
and U1530 (N_1530,N_1461,N_1411);
and U1531 (N_1531,N_1432,N_1419);
xnor U1532 (N_1532,N_1496,N_1464);
xor U1533 (N_1533,N_1477,N_1410);
xnor U1534 (N_1534,N_1459,N_1485);
and U1535 (N_1535,N_1403,N_1437);
and U1536 (N_1536,N_1430,N_1429);
and U1537 (N_1537,N_1423,N_1420);
nand U1538 (N_1538,N_1407,N_1434);
nand U1539 (N_1539,N_1404,N_1412);
nor U1540 (N_1540,N_1401,N_1479);
and U1541 (N_1541,N_1447,N_1487);
xnor U1542 (N_1542,N_1480,N_1482);
xnor U1543 (N_1543,N_1495,N_1402);
xor U1544 (N_1544,N_1463,N_1406);
xnor U1545 (N_1545,N_1414,N_1469);
xnor U1546 (N_1546,N_1457,N_1476);
or U1547 (N_1547,N_1416,N_1449);
xor U1548 (N_1548,N_1400,N_1413);
nor U1549 (N_1549,N_1474,N_1489);
nor U1550 (N_1550,N_1488,N_1416);
xor U1551 (N_1551,N_1428,N_1450);
and U1552 (N_1552,N_1495,N_1440);
xor U1553 (N_1553,N_1426,N_1471);
and U1554 (N_1554,N_1405,N_1454);
or U1555 (N_1555,N_1491,N_1470);
xor U1556 (N_1556,N_1448,N_1496);
nand U1557 (N_1557,N_1455,N_1446);
nor U1558 (N_1558,N_1413,N_1455);
and U1559 (N_1559,N_1468,N_1471);
xnor U1560 (N_1560,N_1472,N_1401);
and U1561 (N_1561,N_1494,N_1480);
and U1562 (N_1562,N_1495,N_1417);
or U1563 (N_1563,N_1498,N_1408);
xnor U1564 (N_1564,N_1476,N_1437);
nor U1565 (N_1565,N_1481,N_1430);
xnor U1566 (N_1566,N_1433,N_1400);
and U1567 (N_1567,N_1459,N_1472);
nand U1568 (N_1568,N_1488,N_1423);
nor U1569 (N_1569,N_1461,N_1456);
and U1570 (N_1570,N_1473,N_1469);
or U1571 (N_1571,N_1446,N_1450);
nor U1572 (N_1572,N_1453,N_1443);
or U1573 (N_1573,N_1470,N_1468);
xnor U1574 (N_1574,N_1453,N_1438);
xor U1575 (N_1575,N_1459,N_1499);
or U1576 (N_1576,N_1497,N_1482);
xnor U1577 (N_1577,N_1478,N_1420);
xor U1578 (N_1578,N_1455,N_1423);
or U1579 (N_1579,N_1453,N_1408);
nor U1580 (N_1580,N_1485,N_1466);
and U1581 (N_1581,N_1456,N_1429);
or U1582 (N_1582,N_1487,N_1479);
nand U1583 (N_1583,N_1431,N_1457);
or U1584 (N_1584,N_1477,N_1476);
nor U1585 (N_1585,N_1417,N_1497);
and U1586 (N_1586,N_1455,N_1482);
and U1587 (N_1587,N_1409,N_1415);
nand U1588 (N_1588,N_1463,N_1489);
and U1589 (N_1589,N_1458,N_1495);
and U1590 (N_1590,N_1404,N_1405);
nand U1591 (N_1591,N_1437,N_1425);
and U1592 (N_1592,N_1462,N_1417);
nand U1593 (N_1593,N_1448,N_1425);
or U1594 (N_1594,N_1497,N_1407);
and U1595 (N_1595,N_1430,N_1424);
nand U1596 (N_1596,N_1483,N_1426);
xor U1597 (N_1597,N_1451,N_1415);
xnor U1598 (N_1598,N_1448,N_1432);
xnor U1599 (N_1599,N_1430,N_1432);
or U1600 (N_1600,N_1572,N_1510);
xnor U1601 (N_1601,N_1537,N_1587);
nor U1602 (N_1602,N_1590,N_1564);
nand U1603 (N_1603,N_1595,N_1550);
nand U1604 (N_1604,N_1586,N_1535);
xnor U1605 (N_1605,N_1511,N_1566);
nand U1606 (N_1606,N_1515,N_1505);
xnor U1607 (N_1607,N_1597,N_1528);
or U1608 (N_1608,N_1589,N_1571);
or U1609 (N_1609,N_1512,N_1516);
nand U1610 (N_1610,N_1568,N_1517);
nor U1611 (N_1611,N_1541,N_1534);
xnor U1612 (N_1612,N_1520,N_1581);
nor U1613 (N_1613,N_1563,N_1561);
nor U1614 (N_1614,N_1567,N_1579);
and U1615 (N_1615,N_1542,N_1555);
or U1616 (N_1616,N_1558,N_1538);
nor U1617 (N_1617,N_1594,N_1530);
nand U1618 (N_1618,N_1588,N_1506);
xnor U1619 (N_1619,N_1514,N_1519);
nand U1620 (N_1620,N_1560,N_1500);
or U1621 (N_1621,N_1591,N_1546);
or U1622 (N_1622,N_1559,N_1583);
xor U1623 (N_1623,N_1584,N_1504);
or U1624 (N_1624,N_1562,N_1565);
nand U1625 (N_1625,N_1508,N_1522);
and U1626 (N_1626,N_1526,N_1547);
nor U1627 (N_1627,N_1575,N_1552);
nand U1628 (N_1628,N_1540,N_1525);
and U1629 (N_1629,N_1502,N_1574);
xor U1630 (N_1630,N_1556,N_1569);
nor U1631 (N_1631,N_1532,N_1531);
xor U1632 (N_1632,N_1549,N_1585);
or U1633 (N_1633,N_1557,N_1553);
nor U1634 (N_1634,N_1529,N_1578);
nor U1635 (N_1635,N_1501,N_1507);
or U1636 (N_1636,N_1554,N_1548);
or U1637 (N_1637,N_1570,N_1524);
nand U1638 (N_1638,N_1523,N_1582);
nand U1639 (N_1639,N_1518,N_1573);
or U1640 (N_1640,N_1544,N_1593);
nand U1641 (N_1641,N_1580,N_1527);
xnor U1642 (N_1642,N_1598,N_1599);
or U1643 (N_1643,N_1576,N_1545);
or U1644 (N_1644,N_1596,N_1509);
nor U1645 (N_1645,N_1577,N_1536);
or U1646 (N_1646,N_1551,N_1539);
xnor U1647 (N_1647,N_1592,N_1503);
nor U1648 (N_1648,N_1521,N_1533);
and U1649 (N_1649,N_1513,N_1543);
xor U1650 (N_1650,N_1575,N_1518);
nand U1651 (N_1651,N_1556,N_1519);
or U1652 (N_1652,N_1541,N_1579);
xor U1653 (N_1653,N_1597,N_1578);
or U1654 (N_1654,N_1599,N_1596);
or U1655 (N_1655,N_1593,N_1566);
xor U1656 (N_1656,N_1540,N_1510);
nand U1657 (N_1657,N_1534,N_1592);
nand U1658 (N_1658,N_1504,N_1553);
nand U1659 (N_1659,N_1514,N_1597);
and U1660 (N_1660,N_1548,N_1553);
nor U1661 (N_1661,N_1531,N_1595);
nand U1662 (N_1662,N_1588,N_1570);
or U1663 (N_1663,N_1588,N_1504);
xnor U1664 (N_1664,N_1527,N_1514);
or U1665 (N_1665,N_1508,N_1591);
nand U1666 (N_1666,N_1534,N_1553);
nand U1667 (N_1667,N_1515,N_1587);
and U1668 (N_1668,N_1538,N_1592);
nor U1669 (N_1669,N_1540,N_1533);
nor U1670 (N_1670,N_1563,N_1575);
xor U1671 (N_1671,N_1592,N_1520);
xnor U1672 (N_1672,N_1529,N_1560);
nand U1673 (N_1673,N_1579,N_1559);
nand U1674 (N_1674,N_1500,N_1531);
nor U1675 (N_1675,N_1513,N_1556);
and U1676 (N_1676,N_1529,N_1563);
xor U1677 (N_1677,N_1566,N_1515);
nor U1678 (N_1678,N_1596,N_1593);
xnor U1679 (N_1679,N_1500,N_1525);
or U1680 (N_1680,N_1549,N_1588);
and U1681 (N_1681,N_1522,N_1568);
and U1682 (N_1682,N_1545,N_1583);
nand U1683 (N_1683,N_1538,N_1559);
xor U1684 (N_1684,N_1595,N_1556);
nand U1685 (N_1685,N_1555,N_1557);
or U1686 (N_1686,N_1592,N_1516);
nor U1687 (N_1687,N_1542,N_1590);
nand U1688 (N_1688,N_1518,N_1535);
nand U1689 (N_1689,N_1567,N_1569);
xor U1690 (N_1690,N_1552,N_1541);
xor U1691 (N_1691,N_1517,N_1509);
and U1692 (N_1692,N_1573,N_1528);
xnor U1693 (N_1693,N_1511,N_1571);
xor U1694 (N_1694,N_1543,N_1515);
or U1695 (N_1695,N_1570,N_1533);
nor U1696 (N_1696,N_1568,N_1581);
nand U1697 (N_1697,N_1559,N_1589);
and U1698 (N_1698,N_1591,N_1512);
nor U1699 (N_1699,N_1510,N_1504);
nand U1700 (N_1700,N_1644,N_1665);
nor U1701 (N_1701,N_1647,N_1651);
nor U1702 (N_1702,N_1609,N_1640);
and U1703 (N_1703,N_1611,N_1666);
nor U1704 (N_1704,N_1663,N_1691);
nand U1705 (N_1705,N_1690,N_1637);
nor U1706 (N_1706,N_1671,N_1689);
nor U1707 (N_1707,N_1607,N_1688);
xnor U1708 (N_1708,N_1606,N_1603);
nor U1709 (N_1709,N_1675,N_1653);
nor U1710 (N_1710,N_1601,N_1669);
xor U1711 (N_1711,N_1655,N_1652);
nor U1712 (N_1712,N_1623,N_1670);
nor U1713 (N_1713,N_1639,N_1679);
and U1714 (N_1714,N_1682,N_1698);
xnor U1715 (N_1715,N_1614,N_1605);
nand U1716 (N_1716,N_1622,N_1642);
xor U1717 (N_1717,N_1648,N_1677);
nand U1718 (N_1718,N_1624,N_1631);
xor U1719 (N_1719,N_1613,N_1649);
xnor U1720 (N_1720,N_1683,N_1617);
and U1721 (N_1721,N_1636,N_1621);
xnor U1722 (N_1722,N_1630,N_1654);
and U1723 (N_1723,N_1638,N_1626);
and U1724 (N_1724,N_1645,N_1650);
xnor U1725 (N_1725,N_1604,N_1673);
nor U1726 (N_1726,N_1608,N_1668);
nand U1727 (N_1727,N_1612,N_1667);
nor U1728 (N_1728,N_1684,N_1643);
and U1729 (N_1729,N_1672,N_1662);
and U1730 (N_1730,N_1619,N_1687);
nor U1731 (N_1731,N_1680,N_1674);
nor U1732 (N_1732,N_1678,N_1676);
and U1733 (N_1733,N_1646,N_1685);
xor U1734 (N_1734,N_1656,N_1697);
nor U1735 (N_1735,N_1694,N_1686);
xor U1736 (N_1736,N_1699,N_1600);
and U1737 (N_1737,N_1661,N_1658);
xnor U1738 (N_1738,N_1664,N_1620);
and U1739 (N_1739,N_1695,N_1632);
or U1740 (N_1740,N_1628,N_1634);
nor U1741 (N_1741,N_1660,N_1641);
nand U1742 (N_1742,N_1610,N_1616);
nor U1743 (N_1743,N_1602,N_1618);
xnor U1744 (N_1744,N_1692,N_1657);
nor U1745 (N_1745,N_1693,N_1625);
xor U1746 (N_1746,N_1635,N_1627);
xor U1747 (N_1747,N_1681,N_1615);
and U1748 (N_1748,N_1629,N_1633);
and U1749 (N_1749,N_1659,N_1696);
or U1750 (N_1750,N_1643,N_1644);
nand U1751 (N_1751,N_1692,N_1628);
nor U1752 (N_1752,N_1620,N_1683);
nor U1753 (N_1753,N_1681,N_1687);
and U1754 (N_1754,N_1665,N_1624);
nand U1755 (N_1755,N_1699,N_1658);
and U1756 (N_1756,N_1692,N_1671);
xor U1757 (N_1757,N_1693,N_1618);
nor U1758 (N_1758,N_1692,N_1661);
nor U1759 (N_1759,N_1611,N_1672);
nand U1760 (N_1760,N_1647,N_1646);
and U1761 (N_1761,N_1694,N_1645);
and U1762 (N_1762,N_1609,N_1643);
and U1763 (N_1763,N_1635,N_1691);
and U1764 (N_1764,N_1619,N_1607);
and U1765 (N_1765,N_1693,N_1691);
nor U1766 (N_1766,N_1622,N_1660);
or U1767 (N_1767,N_1636,N_1673);
xor U1768 (N_1768,N_1672,N_1607);
nor U1769 (N_1769,N_1624,N_1637);
nor U1770 (N_1770,N_1678,N_1697);
nor U1771 (N_1771,N_1692,N_1646);
xor U1772 (N_1772,N_1648,N_1617);
and U1773 (N_1773,N_1678,N_1686);
nand U1774 (N_1774,N_1633,N_1635);
nand U1775 (N_1775,N_1673,N_1669);
and U1776 (N_1776,N_1669,N_1687);
nand U1777 (N_1777,N_1641,N_1638);
nor U1778 (N_1778,N_1606,N_1611);
xnor U1779 (N_1779,N_1662,N_1654);
or U1780 (N_1780,N_1687,N_1629);
and U1781 (N_1781,N_1673,N_1642);
or U1782 (N_1782,N_1647,N_1639);
xor U1783 (N_1783,N_1651,N_1657);
or U1784 (N_1784,N_1629,N_1606);
or U1785 (N_1785,N_1669,N_1644);
nor U1786 (N_1786,N_1647,N_1652);
and U1787 (N_1787,N_1609,N_1654);
and U1788 (N_1788,N_1620,N_1661);
nand U1789 (N_1789,N_1667,N_1607);
xnor U1790 (N_1790,N_1633,N_1600);
xor U1791 (N_1791,N_1672,N_1610);
xnor U1792 (N_1792,N_1648,N_1659);
nand U1793 (N_1793,N_1656,N_1682);
and U1794 (N_1794,N_1611,N_1657);
and U1795 (N_1795,N_1611,N_1625);
or U1796 (N_1796,N_1630,N_1626);
and U1797 (N_1797,N_1657,N_1602);
xor U1798 (N_1798,N_1633,N_1667);
nand U1799 (N_1799,N_1674,N_1624);
or U1800 (N_1800,N_1729,N_1719);
or U1801 (N_1801,N_1773,N_1758);
nor U1802 (N_1802,N_1731,N_1754);
or U1803 (N_1803,N_1718,N_1743);
xnor U1804 (N_1804,N_1797,N_1732);
xor U1805 (N_1805,N_1733,N_1791);
xnor U1806 (N_1806,N_1761,N_1728);
nor U1807 (N_1807,N_1755,N_1711);
xnor U1808 (N_1808,N_1749,N_1796);
xor U1809 (N_1809,N_1766,N_1715);
and U1810 (N_1810,N_1785,N_1787);
nand U1811 (N_1811,N_1792,N_1793);
xnor U1812 (N_1812,N_1710,N_1717);
or U1813 (N_1813,N_1708,N_1751);
and U1814 (N_1814,N_1722,N_1744);
nand U1815 (N_1815,N_1701,N_1727);
nor U1816 (N_1816,N_1794,N_1712);
nand U1817 (N_1817,N_1740,N_1720);
xor U1818 (N_1818,N_1770,N_1788);
and U1819 (N_1819,N_1704,N_1735);
and U1820 (N_1820,N_1772,N_1769);
nor U1821 (N_1821,N_1777,N_1762);
nor U1822 (N_1822,N_1768,N_1783);
xnor U1823 (N_1823,N_1790,N_1778);
nor U1824 (N_1824,N_1747,N_1725);
xor U1825 (N_1825,N_1784,N_1700);
nand U1826 (N_1826,N_1764,N_1746);
nor U1827 (N_1827,N_1702,N_1709);
nand U1828 (N_1828,N_1734,N_1713);
or U1829 (N_1829,N_1737,N_1706);
or U1830 (N_1830,N_1767,N_1741);
or U1831 (N_1831,N_1799,N_1745);
or U1832 (N_1832,N_1795,N_1765);
and U1833 (N_1833,N_1757,N_1748);
or U1834 (N_1834,N_1782,N_1730);
or U1835 (N_1835,N_1739,N_1775);
xnor U1836 (N_1836,N_1716,N_1752);
xor U1837 (N_1837,N_1724,N_1726);
xor U1838 (N_1838,N_1736,N_1798);
nand U1839 (N_1839,N_1781,N_1753);
xnor U1840 (N_1840,N_1789,N_1771);
and U1841 (N_1841,N_1756,N_1742);
nand U1842 (N_1842,N_1763,N_1776);
nand U1843 (N_1843,N_1721,N_1786);
or U1844 (N_1844,N_1723,N_1779);
nor U1845 (N_1845,N_1750,N_1714);
xor U1846 (N_1846,N_1774,N_1703);
nand U1847 (N_1847,N_1760,N_1759);
and U1848 (N_1848,N_1738,N_1705);
and U1849 (N_1849,N_1707,N_1780);
nor U1850 (N_1850,N_1742,N_1722);
and U1851 (N_1851,N_1798,N_1782);
or U1852 (N_1852,N_1758,N_1705);
or U1853 (N_1853,N_1786,N_1702);
xnor U1854 (N_1854,N_1795,N_1711);
nor U1855 (N_1855,N_1714,N_1793);
nor U1856 (N_1856,N_1797,N_1751);
or U1857 (N_1857,N_1791,N_1712);
or U1858 (N_1858,N_1735,N_1702);
nor U1859 (N_1859,N_1752,N_1794);
or U1860 (N_1860,N_1706,N_1726);
xnor U1861 (N_1861,N_1773,N_1775);
nor U1862 (N_1862,N_1722,N_1743);
or U1863 (N_1863,N_1729,N_1782);
or U1864 (N_1864,N_1747,N_1756);
nor U1865 (N_1865,N_1753,N_1789);
nor U1866 (N_1866,N_1778,N_1744);
xnor U1867 (N_1867,N_1744,N_1749);
xor U1868 (N_1868,N_1706,N_1727);
and U1869 (N_1869,N_1786,N_1771);
nor U1870 (N_1870,N_1794,N_1709);
or U1871 (N_1871,N_1753,N_1702);
nand U1872 (N_1872,N_1754,N_1718);
nor U1873 (N_1873,N_1719,N_1734);
nand U1874 (N_1874,N_1709,N_1712);
nor U1875 (N_1875,N_1771,N_1755);
or U1876 (N_1876,N_1781,N_1756);
nand U1877 (N_1877,N_1753,N_1773);
nand U1878 (N_1878,N_1701,N_1729);
and U1879 (N_1879,N_1799,N_1752);
xor U1880 (N_1880,N_1714,N_1704);
and U1881 (N_1881,N_1778,N_1767);
and U1882 (N_1882,N_1725,N_1787);
and U1883 (N_1883,N_1744,N_1792);
or U1884 (N_1884,N_1769,N_1722);
and U1885 (N_1885,N_1730,N_1781);
nand U1886 (N_1886,N_1747,N_1745);
nor U1887 (N_1887,N_1724,N_1722);
nand U1888 (N_1888,N_1741,N_1735);
nand U1889 (N_1889,N_1766,N_1769);
nand U1890 (N_1890,N_1701,N_1771);
and U1891 (N_1891,N_1786,N_1794);
nor U1892 (N_1892,N_1703,N_1755);
xor U1893 (N_1893,N_1710,N_1798);
nor U1894 (N_1894,N_1719,N_1716);
xor U1895 (N_1895,N_1774,N_1755);
or U1896 (N_1896,N_1709,N_1781);
xnor U1897 (N_1897,N_1751,N_1768);
nand U1898 (N_1898,N_1769,N_1795);
and U1899 (N_1899,N_1716,N_1751);
xnor U1900 (N_1900,N_1894,N_1851);
nand U1901 (N_1901,N_1841,N_1878);
and U1902 (N_1902,N_1867,N_1882);
xnor U1903 (N_1903,N_1835,N_1818);
xor U1904 (N_1904,N_1808,N_1825);
and U1905 (N_1905,N_1837,N_1862);
and U1906 (N_1906,N_1896,N_1870);
xor U1907 (N_1907,N_1840,N_1801);
or U1908 (N_1908,N_1871,N_1852);
and U1909 (N_1909,N_1856,N_1872);
nand U1910 (N_1910,N_1832,N_1849);
xor U1911 (N_1911,N_1884,N_1891);
or U1912 (N_1912,N_1826,N_1815);
nand U1913 (N_1913,N_1888,N_1893);
nand U1914 (N_1914,N_1853,N_1863);
nand U1915 (N_1915,N_1864,N_1881);
or U1916 (N_1916,N_1885,N_1820);
and U1917 (N_1917,N_1824,N_1821);
or U1918 (N_1918,N_1813,N_1836);
and U1919 (N_1919,N_1897,N_1828);
or U1920 (N_1920,N_1810,N_1869);
and U1921 (N_1921,N_1843,N_1857);
or U1922 (N_1922,N_1822,N_1833);
nor U1923 (N_1923,N_1859,N_1834);
or U1924 (N_1924,N_1887,N_1819);
xnor U1925 (N_1925,N_1814,N_1877);
nor U1926 (N_1926,N_1831,N_1874);
xnor U1927 (N_1927,N_1899,N_1865);
xor U1928 (N_1928,N_1812,N_1875);
nor U1929 (N_1929,N_1847,N_1873);
nand U1930 (N_1930,N_1800,N_1889);
xnor U1931 (N_1931,N_1850,N_1890);
nor U1932 (N_1932,N_1838,N_1829);
and U1933 (N_1933,N_1892,N_1809);
or U1934 (N_1934,N_1846,N_1886);
and U1935 (N_1935,N_1844,N_1830);
xor U1936 (N_1936,N_1861,N_1855);
nor U1937 (N_1937,N_1879,N_1805);
nor U1938 (N_1938,N_1845,N_1802);
or U1939 (N_1939,N_1868,N_1817);
or U1940 (N_1940,N_1880,N_1807);
nand U1941 (N_1941,N_1839,N_1806);
and U1942 (N_1942,N_1804,N_1898);
nor U1943 (N_1943,N_1858,N_1876);
nand U1944 (N_1944,N_1883,N_1895);
or U1945 (N_1945,N_1866,N_1811);
xor U1946 (N_1946,N_1823,N_1860);
nor U1947 (N_1947,N_1848,N_1803);
or U1948 (N_1948,N_1854,N_1816);
and U1949 (N_1949,N_1842,N_1827);
or U1950 (N_1950,N_1891,N_1819);
or U1951 (N_1951,N_1863,N_1809);
nand U1952 (N_1952,N_1882,N_1859);
xor U1953 (N_1953,N_1823,N_1837);
nand U1954 (N_1954,N_1826,N_1856);
nand U1955 (N_1955,N_1829,N_1821);
nor U1956 (N_1956,N_1867,N_1842);
nor U1957 (N_1957,N_1881,N_1834);
xor U1958 (N_1958,N_1842,N_1815);
nor U1959 (N_1959,N_1825,N_1877);
and U1960 (N_1960,N_1805,N_1862);
xnor U1961 (N_1961,N_1857,N_1884);
nand U1962 (N_1962,N_1833,N_1816);
and U1963 (N_1963,N_1867,N_1824);
or U1964 (N_1964,N_1833,N_1837);
xor U1965 (N_1965,N_1810,N_1843);
xor U1966 (N_1966,N_1804,N_1832);
and U1967 (N_1967,N_1850,N_1818);
or U1968 (N_1968,N_1868,N_1802);
nand U1969 (N_1969,N_1866,N_1869);
xnor U1970 (N_1970,N_1826,N_1868);
xnor U1971 (N_1971,N_1866,N_1830);
nor U1972 (N_1972,N_1827,N_1889);
xor U1973 (N_1973,N_1812,N_1805);
or U1974 (N_1974,N_1826,N_1820);
and U1975 (N_1975,N_1819,N_1822);
and U1976 (N_1976,N_1834,N_1846);
or U1977 (N_1977,N_1880,N_1824);
xnor U1978 (N_1978,N_1808,N_1850);
xor U1979 (N_1979,N_1844,N_1835);
xor U1980 (N_1980,N_1874,N_1858);
nand U1981 (N_1981,N_1826,N_1831);
xor U1982 (N_1982,N_1833,N_1861);
and U1983 (N_1983,N_1846,N_1843);
or U1984 (N_1984,N_1819,N_1865);
and U1985 (N_1985,N_1858,N_1856);
and U1986 (N_1986,N_1823,N_1869);
nor U1987 (N_1987,N_1891,N_1857);
nand U1988 (N_1988,N_1864,N_1892);
nor U1989 (N_1989,N_1859,N_1815);
xor U1990 (N_1990,N_1802,N_1862);
nand U1991 (N_1991,N_1859,N_1844);
xor U1992 (N_1992,N_1891,N_1823);
and U1993 (N_1993,N_1863,N_1825);
nor U1994 (N_1994,N_1821,N_1828);
or U1995 (N_1995,N_1877,N_1899);
nand U1996 (N_1996,N_1803,N_1872);
nor U1997 (N_1997,N_1886,N_1880);
xor U1998 (N_1998,N_1840,N_1894);
or U1999 (N_1999,N_1855,N_1879);
xor U2000 (N_2000,N_1939,N_1957);
or U2001 (N_2001,N_1992,N_1906);
nand U2002 (N_2002,N_1932,N_1991);
or U2003 (N_2003,N_1931,N_1901);
nor U2004 (N_2004,N_1994,N_1973);
or U2005 (N_2005,N_1928,N_1974);
nor U2006 (N_2006,N_1929,N_1937);
nand U2007 (N_2007,N_1981,N_1976);
nand U2008 (N_2008,N_1987,N_1988);
or U2009 (N_2009,N_1911,N_1977);
and U2010 (N_2010,N_1923,N_1920);
nand U2011 (N_2011,N_1979,N_1902);
and U2012 (N_2012,N_1946,N_1936);
xnor U2013 (N_2013,N_1971,N_1975);
and U2014 (N_2014,N_1954,N_1955);
or U2015 (N_2015,N_1953,N_1986);
and U2016 (N_2016,N_1980,N_1900);
nor U2017 (N_2017,N_1938,N_1903);
nor U2018 (N_2018,N_1927,N_1904);
and U2019 (N_2019,N_1913,N_1941);
or U2020 (N_2020,N_1907,N_1995);
or U2021 (N_2021,N_1969,N_1989);
or U2022 (N_2022,N_1912,N_1965);
nand U2023 (N_2023,N_1984,N_1966);
or U2024 (N_2024,N_1997,N_1999);
or U2025 (N_2025,N_1959,N_1905);
nand U2026 (N_2026,N_1909,N_1910);
or U2027 (N_2027,N_1948,N_1944);
nand U2028 (N_2028,N_1982,N_1908);
xor U2029 (N_2029,N_1915,N_1947);
or U2030 (N_2030,N_1962,N_1935);
nand U2031 (N_2031,N_1993,N_1925);
xor U2032 (N_2032,N_1996,N_1921);
or U2033 (N_2033,N_1926,N_1918);
xor U2034 (N_2034,N_1934,N_1919);
nand U2035 (N_2035,N_1943,N_1968);
nor U2036 (N_2036,N_1952,N_1940);
nor U2037 (N_2037,N_1978,N_1964);
xnor U2038 (N_2038,N_1924,N_1960);
nor U2039 (N_2039,N_1922,N_1917);
nor U2040 (N_2040,N_1950,N_1983);
nor U2041 (N_2041,N_1956,N_1949);
or U2042 (N_2042,N_1930,N_1933);
or U2043 (N_2043,N_1951,N_1945);
or U2044 (N_2044,N_1972,N_1985);
nor U2045 (N_2045,N_1967,N_1970);
nand U2046 (N_2046,N_1990,N_1961);
or U2047 (N_2047,N_1914,N_1916);
nor U2048 (N_2048,N_1963,N_1942);
or U2049 (N_2049,N_1998,N_1958);
nand U2050 (N_2050,N_1921,N_1940);
or U2051 (N_2051,N_1923,N_1925);
and U2052 (N_2052,N_1940,N_1933);
and U2053 (N_2053,N_1924,N_1933);
nand U2054 (N_2054,N_1929,N_1940);
xor U2055 (N_2055,N_1983,N_1901);
and U2056 (N_2056,N_1933,N_1922);
and U2057 (N_2057,N_1982,N_1921);
nor U2058 (N_2058,N_1965,N_1918);
and U2059 (N_2059,N_1948,N_1940);
and U2060 (N_2060,N_1989,N_1943);
nand U2061 (N_2061,N_1971,N_1963);
and U2062 (N_2062,N_1952,N_1949);
nand U2063 (N_2063,N_1985,N_1926);
and U2064 (N_2064,N_1975,N_1985);
xor U2065 (N_2065,N_1908,N_1960);
and U2066 (N_2066,N_1990,N_1935);
and U2067 (N_2067,N_1964,N_1938);
and U2068 (N_2068,N_1980,N_1975);
nand U2069 (N_2069,N_1928,N_1983);
and U2070 (N_2070,N_1942,N_1924);
nand U2071 (N_2071,N_1926,N_1920);
or U2072 (N_2072,N_1910,N_1970);
xnor U2073 (N_2073,N_1942,N_1990);
nand U2074 (N_2074,N_1941,N_1964);
nor U2075 (N_2075,N_1969,N_1910);
or U2076 (N_2076,N_1973,N_1974);
xnor U2077 (N_2077,N_1944,N_1900);
nand U2078 (N_2078,N_1939,N_1906);
xor U2079 (N_2079,N_1954,N_1972);
xor U2080 (N_2080,N_1938,N_1901);
xor U2081 (N_2081,N_1920,N_1995);
and U2082 (N_2082,N_1913,N_1926);
or U2083 (N_2083,N_1959,N_1902);
nand U2084 (N_2084,N_1951,N_1987);
xnor U2085 (N_2085,N_1930,N_1944);
or U2086 (N_2086,N_1950,N_1902);
or U2087 (N_2087,N_1994,N_1916);
nor U2088 (N_2088,N_1960,N_1915);
nand U2089 (N_2089,N_1966,N_1958);
and U2090 (N_2090,N_1919,N_1996);
xor U2091 (N_2091,N_1986,N_1983);
nand U2092 (N_2092,N_1952,N_1931);
and U2093 (N_2093,N_1962,N_1938);
xor U2094 (N_2094,N_1900,N_1920);
nor U2095 (N_2095,N_1921,N_1933);
nor U2096 (N_2096,N_1992,N_1943);
and U2097 (N_2097,N_1991,N_1987);
and U2098 (N_2098,N_1928,N_1994);
xor U2099 (N_2099,N_1934,N_1943);
xnor U2100 (N_2100,N_2015,N_2078);
xnor U2101 (N_2101,N_2096,N_2067);
nor U2102 (N_2102,N_2050,N_2033);
xor U2103 (N_2103,N_2093,N_2017);
and U2104 (N_2104,N_2046,N_2084);
xnor U2105 (N_2105,N_2064,N_2082);
xnor U2106 (N_2106,N_2020,N_2010);
nand U2107 (N_2107,N_2094,N_2034);
xnor U2108 (N_2108,N_2024,N_2081);
nand U2109 (N_2109,N_2023,N_2025);
and U2110 (N_2110,N_2095,N_2083);
nand U2111 (N_2111,N_2035,N_2047);
and U2112 (N_2112,N_2055,N_2089);
nand U2113 (N_2113,N_2085,N_2063);
xor U2114 (N_2114,N_2036,N_2026);
and U2115 (N_2115,N_2099,N_2006);
nand U2116 (N_2116,N_2057,N_2054);
xnor U2117 (N_2117,N_2028,N_2002);
nand U2118 (N_2118,N_2011,N_2073);
or U2119 (N_2119,N_2021,N_2042);
nand U2120 (N_2120,N_2014,N_2071);
nor U2121 (N_2121,N_2045,N_2030);
and U2122 (N_2122,N_2003,N_2065);
xnor U2123 (N_2123,N_2049,N_2075);
xor U2124 (N_2124,N_2088,N_2019);
and U2125 (N_2125,N_2016,N_2087);
xnor U2126 (N_2126,N_2097,N_2041);
xor U2127 (N_2127,N_2005,N_2008);
nor U2128 (N_2128,N_2076,N_2051);
or U2129 (N_2129,N_2080,N_2068);
xnor U2130 (N_2130,N_2069,N_2052);
or U2131 (N_2131,N_2038,N_2091);
xnor U2132 (N_2132,N_2031,N_2059);
or U2133 (N_2133,N_2060,N_2098);
xor U2134 (N_2134,N_2044,N_2048);
and U2135 (N_2135,N_2037,N_2032);
nand U2136 (N_2136,N_2022,N_2039);
and U2137 (N_2137,N_2070,N_2062);
xnor U2138 (N_2138,N_2029,N_2013);
xor U2139 (N_2139,N_2074,N_2027);
xnor U2140 (N_2140,N_2092,N_2000);
and U2141 (N_2141,N_2086,N_2090);
nand U2142 (N_2142,N_2053,N_2043);
and U2143 (N_2143,N_2072,N_2079);
nor U2144 (N_2144,N_2077,N_2009);
xor U2145 (N_2145,N_2066,N_2007);
xnor U2146 (N_2146,N_2040,N_2058);
nand U2147 (N_2147,N_2018,N_2056);
xnor U2148 (N_2148,N_2061,N_2004);
nor U2149 (N_2149,N_2012,N_2001);
xor U2150 (N_2150,N_2013,N_2020);
and U2151 (N_2151,N_2033,N_2047);
or U2152 (N_2152,N_2062,N_2068);
nand U2153 (N_2153,N_2046,N_2051);
or U2154 (N_2154,N_2055,N_2067);
nand U2155 (N_2155,N_2010,N_2083);
nand U2156 (N_2156,N_2053,N_2057);
nor U2157 (N_2157,N_2099,N_2090);
nor U2158 (N_2158,N_2046,N_2049);
nand U2159 (N_2159,N_2090,N_2094);
xor U2160 (N_2160,N_2014,N_2088);
or U2161 (N_2161,N_2014,N_2007);
xnor U2162 (N_2162,N_2053,N_2004);
nor U2163 (N_2163,N_2062,N_2061);
xor U2164 (N_2164,N_2055,N_2033);
or U2165 (N_2165,N_2008,N_2099);
nor U2166 (N_2166,N_2051,N_2019);
nor U2167 (N_2167,N_2073,N_2042);
nor U2168 (N_2168,N_2050,N_2091);
or U2169 (N_2169,N_2013,N_2072);
and U2170 (N_2170,N_2098,N_2022);
or U2171 (N_2171,N_2010,N_2026);
xor U2172 (N_2172,N_2088,N_2039);
xor U2173 (N_2173,N_2069,N_2033);
or U2174 (N_2174,N_2083,N_2053);
or U2175 (N_2175,N_2031,N_2045);
nand U2176 (N_2176,N_2024,N_2032);
xor U2177 (N_2177,N_2008,N_2053);
nand U2178 (N_2178,N_2002,N_2016);
nand U2179 (N_2179,N_2056,N_2013);
nor U2180 (N_2180,N_2022,N_2081);
nor U2181 (N_2181,N_2050,N_2049);
and U2182 (N_2182,N_2032,N_2096);
xnor U2183 (N_2183,N_2026,N_2028);
nor U2184 (N_2184,N_2079,N_2000);
nand U2185 (N_2185,N_2031,N_2044);
nor U2186 (N_2186,N_2040,N_2050);
and U2187 (N_2187,N_2051,N_2026);
nor U2188 (N_2188,N_2055,N_2034);
or U2189 (N_2189,N_2023,N_2031);
nor U2190 (N_2190,N_2090,N_2029);
xor U2191 (N_2191,N_2040,N_2020);
and U2192 (N_2192,N_2028,N_2063);
or U2193 (N_2193,N_2077,N_2066);
nand U2194 (N_2194,N_2012,N_2089);
or U2195 (N_2195,N_2083,N_2058);
nor U2196 (N_2196,N_2090,N_2000);
nand U2197 (N_2197,N_2012,N_2088);
xnor U2198 (N_2198,N_2017,N_2097);
nand U2199 (N_2199,N_2027,N_2009);
nor U2200 (N_2200,N_2183,N_2144);
xor U2201 (N_2201,N_2185,N_2103);
or U2202 (N_2202,N_2121,N_2184);
or U2203 (N_2203,N_2142,N_2131);
nand U2204 (N_2204,N_2186,N_2165);
and U2205 (N_2205,N_2106,N_2126);
xnor U2206 (N_2206,N_2161,N_2176);
or U2207 (N_2207,N_2115,N_2174);
xnor U2208 (N_2208,N_2110,N_2141);
nor U2209 (N_2209,N_2128,N_2164);
and U2210 (N_2210,N_2145,N_2118);
and U2211 (N_2211,N_2112,N_2133);
nor U2212 (N_2212,N_2170,N_2187);
nor U2213 (N_2213,N_2125,N_2175);
nand U2214 (N_2214,N_2138,N_2114);
nand U2215 (N_2215,N_2116,N_2182);
nand U2216 (N_2216,N_2166,N_2129);
or U2217 (N_2217,N_2196,N_2140);
nor U2218 (N_2218,N_2151,N_2163);
nand U2219 (N_2219,N_2194,N_2190);
nor U2220 (N_2220,N_2159,N_2152);
nor U2221 (N_2221,N_2100,N_2168);
nand U2222 (N_2222,N_2188,N_2177);
xnor U2223 (N_2223,N_2146,N_2179);
nand U2224 (N_2224,N_2192,N_2117);
or U2225 (N_2225,N_2173,N_2111);
or U2226 (N_2226,N_2137,N_2139);
xnor U2227 (N_2227,N_2154,N_2149);
or U2228 (N_2228,N_2135,N_2119);
nand U2229 (N_2229,N_2171,N_2143);
or U2230 (N_2230,N_2156,N_2122);
nor U2231 (N_2231,N_2157,N_2123);
or U2232 (N_2232,N_2199,N_2162);
nand U2233 (N_2233,N_2191,N_2181);
xnor U2234 (N_2234,N_2178,N_2198);
xor U2235 (N_2235,N_2172,N_2113);
nand U2236 (N_2236,N_2101,N_2153);
and U2237 (N_2237,N_2155,N_2147);
nor U2238 (N_2238,N_2132,N_2150);
nand U2239 (N_2239,N_2104,N_2124);
and U2240 (N_2240,N_2148,N_2108);
and U2241 (N_2241,N_2180,N_2169);
nand U2242 (N_2242,N_2197,N_2160);
nand U2243 (N_2243,N_2167,N_2136);
xnor U2244 (N_2244,N_2109,N_2102);
nand U2245 (N_2245,N_2134,N_2120);
nand U2246 (N_2246,N_2127,N_2130);
nand U2247 (N_2247,N_2195,N_2105);
nor U2248 (N_2248,N_2158,N_2193);
or U2249 (N_2249,N_2107,N_2189);
nand U2250 (N_2250,N_2125,N_2139);
nand U2251 (N_2251,N_2167,N_2148);
xnor U2252 (N_2252,N_2182,N_2184);
nor U2253 (N_2253,N_2199,N_2133);
nand U2254 (N_2254,N_2190,N_2185);
and U2255 (N_2255,N_2126,N_2124);
or U2256 (N_2256,N_2133,N_2141);
nor U2257 (N_2257,N_2166,N_2151);
xnor U2258 (N_2258,N_2189,N_2171);
nor U2259 (N_2259,N_2198,N_2126);
or U2260 (N_2260,N_2175,N_2139);
nand U2261 (N_2261,N_2139,N_2124);
or U2262 (N_2262,N_2185,N_2174);
or U2263 (N_2263,N_2140,N_2159);
nand U2264 (N_2264,N_2150,N_2142);
nor U2265 (N_2265,N_2168,N_2117);
nand U2266 (N_2266,N_2181,N_2124);
xor U2267 (N_2267,N_2118,N_2155);
or U2268 (N_2268,N_2156,N_2143);
or U2269 (N_2269,N_2107,N_2147);
or U2270 (N_2270,N_2148,N_2168);
nor U2271 (N_2271,N_2120,N_2114);
nor U2272 (N_2272,N_2132,N_2195);
nand U2273 (N_2273,N_2169,N_2177);
nor U2274 (N_2274,N_2152,N_2187);
and U2275 (N_2275,N_2122,N_2184);
and U2276 (N_2276,N_2106,N_2140);
xnor U2277 (N_2277,N_2131,N_2114);
and U2278 (N_2278,N_2110,N_2176);
and U2279 (N_2279,N_2159,N_2147);
or U2280 (N_2280,N_2168,N_2176);
or U2281 (N_2281,N_2144,N_2109);
and U2282 (N_2282,N_2166,N_2132);
xnor U2283 (N_2283,N_2139,N_2131);
nor U2284 (N_2284,N_2171,N_2128);
and U2285 (N_2285,N_2100,N_2105);
nand U2286 (N_2286,N_2115,N_2192);
nand U2287 (N_2287,N_2149,N_2106);
or U2288 (N_2288,N_2119,N_2141);
nor U2289 (N_2289,N_2142,N_2143);
nor U2290 (N_2290,N_2150,N_2178);
nand U2291 (N_2291,N_2137,N_2129);
and U2292 (N_2292,N_2185,N_2142);
nand U2293 (N_2293,N_2197,N_2188);
and U2294 (N_2294,N_2112,N_2138);
nor U2295 (N_2295,N_2185,N_2111);
nand U2296 (N_2296,N_2149,N_2193);
xor U2297 (N_2297,N_2179,N_2108);
nand U2298 (N_2298,N_2130,N_2109);
or U2299 (N_2299,N_2163,N_2108);
and U2300 (N_2300,N_2286,N_2220);
or U2301 (N_2301,N_2211,N_2247);
nand U2302 (N_2302,N_2232,N_2219);
nand U2303 (N_2303,N_2237,N_2267);
xnor U2304 (N_2304,N_2207,N_2288);
and U2305 (N_2305,N_2203,N_2298);
and U2306 (N_2306,N_2238,N_2208);
or U2307 (N_2307,N_2221,N_2278);
nor U2308 (N_2308,N_2281,N_2218);
or U2309 (N_2309,N_2293,N_2276);
or U2310 (N_2310,N_2223,N_2215);
nor U2311 (N_2311,N_2204,N_2240);
and U2312 (N_2312,N_2290,N_2214);
and U2313 (N_2313,N_2212,N_2255);
xnor U2314 (N_2314,N_2277,N_2206);
nand U2315 (N_2315,N_2231,N_2258);
and U2316 (N_2316,N_2254,N_2263);
nor U2317 (N_2317,N_2269,N_2248);
or U2318 (N_2318,N_2279,N_2268);
and U2319 (N_2319,N_2274,N_2210);
or U2320 (N_2320,N_2201,N_2245);
and U2321 (N_2321,N_2285,N_2236);
and U2322 (N_2322,N_2283,N_2234);
and U2323 (N_2323,N_2249,N_2256);
xor U2324 (N_2324,N_2239,N_2202);
nand U2325 (N_2325,N_2227,N_2297);
and U2326 (N_2326,N_2250,N_2216);
or U2327 (N_2327,N_2270,N_2222);
and U2328 (N_2328,N_2253,N_2252);
xor U2329 (N_2329,N_2233,N_2244);
or U2330 (N_2330,N_2229,N_2224);
xnor U2331 (N_2331,N_2226,N_2296);
or U2332 (N_2332,N_2299,N_2213);
and U2333 (N_2333,N_2260,N_2217);
nor U2334 (N_2334,N_2225,N_2265);
nor U2335 (N_2335,N_2266,N_2264);
and U2336 (N_2336,N_2228,N_2284);
xor U2337 (N_2337,N_2261,N_2205);
and U2338 (N_2338,N_2251,N_2295);
or U2339 (N_2339,N_2292,N_2271);
xnor U2340 (N_2340,N_2243,N_2280);
nor U2341 (N_2341,N_2259,N_2282);
nand U2342 (N_2342,N_2262,N_2209);
and U2343 (N_2343,N_2272,N_2294);
nand U2344 (N_2344,N_2242,N_2287);
nor U2345 (N_2345,N_2235,N_2291);
nand U2346 (N_2346,N_2246,N_2241);
nor U2347 (N_2347,N_2289,N_2257);
nor U2348 (N_2348,N_2275,N_2200);
xnor U2349 (N_2349,N_2273,N_2230);
xnor U2350 (N_2350,N_2295,N_2238);
and U2351 (N_2351,N_2278,N_2232);
xnor U2352 (N_2352,N_2233,N_2222);
nor U2353 (N_2353,N_2292,N_2201);
and U2354 (N_2354,N_2241,N_2214);
nand U2355 (N_2355,N_2249,N_2273);
xor U2356 (N_2356,N_2244,N_2265);
nor U2357 (N_2357,N_2288,N_2273);
or U2358 (N_2358,N_2259,N_2237);
or U2359 (N_2359,N_2241,N_2213);
and U2360 (N_2360,N_2265,N_2241);
or U2361 (N_2361,N_2206,N_2224);
nand U2362 (N_2362,N_2277,N_2280);
xor U2363 (N_2363,N_2220,N_2244);
nor U2364 (N_2364,N_2295,N_2269);
or U2365 (N_2365,N_2264,N_2205);
and U2366 (N_2366,N_2229,N_2285);
or U2367 (N_2367,N_2259,N_2249);
or U2368 (N_2368,N_2280,N_2203);
nand U2369 (N_2369,N_2244,N_2286);
nor U2370 (N_2370,N_2261,N_2245);
or U2371 (N_2371,N_2234,N_2233);
nor U2372 (N_2372,N_2216,N_2284);
xnor U2373 (N_2373,N_2236,N_2227);
nor U2374 (N_2374,N_2271,N_2232);
xnor U2375 (N_2375,N_2294,N_2247);
and U2376 (N_2376,N_2254,N_2266);
nor U2377 (N_2377,N_2260,N_2259);
and U2378 (N_2378,N_2299,N_2252);
xnor U2379 (N_2379,N_2200,N_2204);
and U2380 (N_2380,N_2269,N_2215);
nor U2381 (N_2381,N_2250,N_2220);
nor U2382 (N_2382,N_2251,N_2293);
and U2383 (N_2383,N_2282,N_2251);
nand U2384 (N_2384,N_2205,N_2242);
nor U2385 (N_2385,N_2220,N_2248);
and U2386 (N_2386,N_2296,N_2202);
or U2387 (N_2387,N_2235,N_2259);
xnor U2388 (N_2388,N_2255,N_2202);
nand U2389 (N_2389,N_2291,N_2257);
or U2390 (N_2390,N_2233,N_2257);
xnor U2391 (N_2391,N_2244,N_2263);
nor U2392 (N_2392,N_2241,N_2201);
nand U2393 (N_2393,N_2220,N_2283);
nor U2394 (N_2394,N_2297,N_2268);
nor U2395 (N_2395,N_2215,N_2276);
or U2396 (N_2396,N_2214,N_2234);
nand U2397 (N_2397,N_2201,N_2298);
or U2398 (N_2398,N_2262,N_2299);
or U2399 (N_2399,N_2246,N_2292);
and U2400 (N_2400,N_2348,N_2385);
nand U2401 (N_2401,N_2388,N_2387);
nand U2402 (N_2402,N_2391,N_2315);
nand U2403 (N_2403,N_2333,N_2358);
xnor U2404 (N_2404,N_2313,N_2331);
xor U2405 (N_2405,N_2354,N_2304);
or U2406 (N_2406,N_2395,N_2397);
nor U2407 (N_2407,N_2335,N_2320);
nand U2408 (N_2408,N_2334,N_2323);
xor U2409 (N_2409,N_2373,N_2317);
or U2410 (N_2410,N_2303,N_2351);
xor U2411 (N_2411,N_2357,N_2355);
xnor U2412 (N_2412,N_2396,N_2377);
nor U2413 (N_2413,N_2347,N_2393);
nor U2414 (N_2414,N_2306,N_2360);
or U2415 (N_2415,N_2375,N_2380);
nand U2416 (N_2416,N_2302,N_2364);
xor U2417 (N_2417,N_2367,N_2362);
or U2418 (N_2418,N_2341,N_2311);
xor U2419 (N_2419,N_2350,N_2349);
nand U2420 (N_2420,N_2308,N_2370);
nor U2421 (N_2421,N_2369,N_2305);
nand U2422 (N_2422,N_2389,N_2386);
nand U2423 (N_2423,N_2300,N_2316);
nor U2424 (N_2424,N_2314,N_2365);
nor U2425 (N_2425,N_2329,N_2378);
nand U2426 (N_2426,N_2322,N_2366);
or U2427 (N_2427,N_2399,N_2327);
xor U2428 (N_2428,N_2394,N_2346);
xor U2429 (N_2429,N_2336,N_2301);
nor U2430 (N_2430,N_2356,N_2345);
nand U2431 (N_2431,N_2321,N_2309);
nand U2432 (N_2432,N_2374,N_2381);
nand U2433 (N_2433,N_2328,N_2307);
or U2434 (N_2434,N_2332,N_2344);
nor U2435 (N_2435,N_2326,N_2382);
xnor U2436 (N_2436,N_2338,N_2352);
or U2437 (N_2437,N_2379,N_2343);
xnor U2438 (N_2438,N_2376,N_2383);
and U2439 (N_2439,N_2384,N_2325);
nand U2440 (N_2440,N_2319,N_2318);
xnor U2441 (N_2441,N_2392,N_2339);
nand U2442 (N_2442,N_2353,N_2361);
xor U2443 (N_2443,N_2371,N_2372);
xnor U2444 (N_2444,N_2324,N_2337);
and U2445 (N_2445,N_2390,N_2312);
and U2446 (N_2446,N_2368,N_2310);
nand U2447 (N_2447,N_2359,N_2342);
or U2448 (N_2448,N_2330,N_2340);
nor U2449 (N_2449,N_2363,N_2398);
nor U2450 (N_2450,N_2300,N_2384);
or U2451 (N_2451,N_2308,N_2319);
xnor U2452 (N_2452,N_2311,N_2303);
and U2453 (N_2453,N_2374,N_2363);
nand U2454 (N_2454,N_2354,N_2325);
xnor U2455 (N_2455,N_2335,N_2390);
nor U2456 (N_2456,N_2352,N_2331);
or U2457 (N_2457,N_2305,N_2340);
or U2458 (N_2458,N_2305,N_2330);
nor U2459 (N_2459,N_2345,N_2391);
nor U2460 (N_2460,N_2396,N_2384);
and U2461 (N_2461,N_2356,N_2336);
nand U2462 (N_2462,N_2374,N_2349);
nor U2463 (N_2463,N_2332,N_2334);
and U2464 (N_2464,N_2342,N_2324);
and U2465 (N_2465,N_2399,N_2329);
xor U2466 (N_2466,N_2353,N_2351);
nand U2467 (N_2467,N_2356,N_2305);
nor U2468 (N_2468,N_2398,N_2399);
and U2469 (N_2469,N_2381,N_2321);
or U2470 (N_2470,N_2312,N_2388);
xnor U2471 (N_2471,N_2371,N_2336);
or U2472 (N_2472,N_2335,N_2365);
xor U2473 (N_2473,N_2399,N_2392);
nor U2474 (N_2474,N_2391,N_2301);
xor U2475 (N_2475,N_2335,N_2337);
nand U2476 (N_2476,N_2330,N_2379);
and U2477 (N_2477,N_2370,N_2323);
nor U2478 (N_2478,N_2301,N_2321);
or U2479 (N_2479,N_2390,N_2363);
and U2480 (N_2480,N_2366,N_2333);
or U2481 (N_2481,N_2318,N_2300);
nor U2482 (N_2482,N_2390,N_2394);
or U2483 (N_2483,N_2375,N_2302);
or U2484 (N_2484,N_2342,N_2374);
xor U2485 (N_2485,N_2380,N_2346);
nand U2486 (N_2486,N_2388,N_2378);
and U2487 (N_2487,N_2380,N_2317);
and U2488 (N_2488,N_2308,N_2337);
and U2489 (N_2489,N_2386,N_2329);
nor U2490 (N_2490,N_2377,N_2397);
nor U2491 (N_2491,N_2343,N_2381);
and U2492 (N_2492,N_2360,N_2394);
or U2493 (N_2493,N_2310,N_2325);
and U2494 (N_2494,N_2332,N_2315);
nand U2495 (N_2495,N_2372,N_2301);
and U2496 (N_2496,N_2338,N_2355);
and U2497 (N_2497,N_2384,N_2310);
and U2498 (N_2498,N_2358,N_2359);
xor U2499 (N_2499,N_2350,N_2391);
xnor U2500 (N_2500,N_2441,N_2437);
xnor U2501 (N_2501,N_2480,N_2421);
xor U2502 (N_2502,N_2414,N_2450);
or U2503 (N_2503,N_2452,N_2406);
nand U2504 (N_2504,N_2447,N_2422);
nor U2505 (N_2505,N_2412,N_2479);
xor U2506 (N_2506,N_2464,N_2456);
or U2507 (N_2507,N_2433,N_2478);
or U2508 (N_2508,N_2477,N_2492);
nand U2509 (N_2509,N_2411,N_2461);
xnor U2510 (N_2510,N_2484,N_2428);
xor U2511 (N_2511,N_2454,N_2420);
and U2512 (N_2512,N_2405,N_2434);
nand U2513 (N_2513,N_2415,N_2449);
or U2514 (N_2514,N_2486,N_2408);
nor U2515 (N_2515,N_2426,N_2489);
or U2516 (N_2516,N_2400,N_2417);
nand U2517 (N_2517,N_2475,N_2459);
nand U2518 (N_2518,N_2460,N_2407);
nand U2519 (N_2519,N_2443,N_2482);
and U2520 (N_2520,N_2485,N_2453);
nand U2521 (N_2521,N_2465,N_2472);
nand U2522 (N_2522,N_2483,N_2451);
nand U2523 (N_2523,N_2488,N_2413);
nand U2524 (N_2524,N_2455,N_2487);
nand U2525 (N_2525,N_2424,N_2499);
nor U2526 (N_2526,N_2427,N_2444);
nor U2527 (N_2527,N_2419,N_2468);
nor U2528 (N_2528,N_2471,N_2469);
and U2529 (N_2529,N_2463,N_2496);
xor U2530 (N_2530,N_2473,N_2416);
xor U2531 (N_2531,N_2495,N_2448);
and U2532 (N_2532,N_2445,N_2476);
nor U2533 (N_2533,N_2402,N_2493);
nand U2534 (N_2534,N_2401,N_2491);
or U2535 (N_2535,N_2410,N_2497);
and U2536 (N_2536,N_2494,N_2442);
and U2537 (N_2537,N_2462,N_2404);
nor U2538 (N_2538,N_2409,N_2481);
nand U2539 (N_2539,N_2436,N_2490);
xnor U2540 (N_2540,N_2438,N_2425);
nand U2541 (N_2541,N_2440,N_2498);
nor U2542 (N_2542,N_2457,N_2432);
nor U2543 (N_2543,N_2474,N_2466);
nand U2544 (N_2544,N_2430,N_2470);
nor U2545 (N_2545,N_2429,N_2403);
and U2546 (N_2546,N_2446,N_2458);
xnor U2547 (N_2547,N_2435,N_2439);
or U2548 (N_2548,N_2431,N_2423);
xnor U2549 (N_2549,N_2467,N_2418);
or U2550 (N_2550,N_2436,N_2477);
or U2551 (N_2551,N_2437,N_2471);
xnor U2552 (N_2552,N_2425,N_2410);
and U2553 (N_2553,N_2414,N_2436);
nand U2554 (N_2554,N_2436,N_2423);
nor U2555 (N_2555,N_2498,N_2431);
nor U2556 (N_2556,N_2450,N_2415);
or U2557 (N_2557,N_2412,N_2467);
xnor U2558 (N_2558,N_2432,N_2476);
and U2559 (N_2559,N_2421,N_2417);
nand U2560 (N_2560,N_2437,N_2438);
and U2561 (N_2561,N_2446,N_2456);
nor U2562 (N_2562,N_2438,N_2485);
nand U2563 (N_2563,N_2441,N_2498);
xnor U2564 (N_2564,N_2429,N_2460);
nor U2565 (N_2565,N_2479,N_2438);
nand U2566 (N_2566,N_2408,N_2456);
nand U2567 (N_2567,N_2488,N_2437);
or U2568 (N_2568,N_2410,N_2471);
and U2569 (N_2569,N_2466,N_2437);
nor U2570 (N_2570,N_2483,N_2475);
nor U2571 (N_2571,N_2464,N_2470);
nand U2572 (N_2572,N_2432,N_2407);
or U2573 (N_2573,N_2442,N_2438);
nor U2574 (N_2574,N_2408,N_2448);
nor U2575 (N_2575,N_2421,N_2431);
and U2576 (N_2576,N_2440,N_2458);
or U2577 (N_2577,N_2401,N_2418);
nor U2578 (N_2578,N_2450,N_2444);
xnor U2579 (N_2579,N_2425,N_2409);
or U2580 (N_2580,N_2434,N_2429);
and U2581 (N_2581,N_2407,N_2437);
xnor U2582 (N_2582,N_2403,N_2432);
nand U2583 (N_2583,N_2484,N_2446);
nor U2584 (N_2584,N_2408,N_2437);
and U2585 (N_2585,N_2439,N_2418);
and U2586 (N_2586,N_2461,N_2418);
nand U2587 (N_2587,N_2486,N_2446);
nor U2588 (N_2588,N_2466,N_2403);
or U2589 (N_2589,N_2454,N_2449);
xor U2590 (N_2590,N_2429,N_2401);
and U2591 (N_2591,N_2452,N_2454);
or U2592 (N_2592,N_2448,N_2436);
xor U2593 (N_2593,N_2446,N_2427);
nor U2594 (N_2594,N_2459,N_2427);
and U2595 (N_2595,N_2429,N_2464);
and U2596 (N_2596,N_2404,N_2434);
xor U2597 (N_2597,N_2469,N_2441);
nand U2598 (N_2598,N_2426,N_2403);
xnor U2599 (N_2599,N_2483,N_2463);
nand U2600 (N_2600,N_2565,N_2524);
and U2601 (N_2601,N_2589,N_2507);
nand U2602 (N_2602,N_2512,N_2564);
xor U2603 (N_2603,N_2548,N_2595);
nor U2604 (N_2604,N_2581,N_2515);
nand U2605 (N_2605,N_2547,N_2500);
and U2606 (N_2606,N_2527,N_2592);
and U2607 (N_2607,N_2552,N_2528);
xnor U2608 (N_2608,N_2517,N_2522);
xnor U2609 (N_2609,N_2573,N_2519);
or U2610 (N_2610,N_2577,N_2584);
xnor U2611 (N_2611,N_2599,N_2541);
nor U2612 (N_2612,N_2516,N_2562);
nor U2613 (N_2613,N_2591,N_2555);
xnor U2614 (N_2614,N_2576,N_2505);
xor U2615 (N_2615,N_2590,N_2597);
and U2616 (N_2616,N_2575,N_2570);
or U2617 (N_2617,N_2518,N_2574);
and U2618 (N_2618,N_2523,N_2593);
or U2619 (N_2619,N_2556,N_2543);
and U2620 (N_2620,N_2532,N_2572);
xor U2621 (N_2621,N_2582,N_2549);
and U2622 (N_2622,N_2509,N_2558);
or U2623 (N_2623,N_2506,N_2571);
and U2624 (N_2624,N_2537,N_2540);
xor U2625 (N_2625,N_2554,N_2568);
xnor U2626 (N_2626,N_2508,N_2533);
and U2627 (N_2627,N_2578,N_2586);
nand U2628 (N_2628,N_2531,N_2596);
or U2629 (N_2629,N_2553,N_2526);
nor U2630 (N_2630,N_2587,N_2594);
nor U2631 (N_2631,N_2567,N_2513);
nor U2632 (N_2632,N_2538,N_2511);
and U2633 (N_2633,N_2520,N_2550);
nor U2634 (N_2634,N_2566,N_2545);
or U2635 (N_2635,N_2504,N_2534);
nor U2636 (N_2636,N_2560,N_2563);
and U2637 (N_2637,N_2535,N_2510);
nand U2638 (N_2638,N_2546,N_2536);
nand U2639 (N_2639,N_2502,N_2501);
and U2640 (N_2640,N_2588,N_2529);
nor U2641 (N_2641,N_2539,N_2525);
nor U2642 (N_2642,N_2561,N_2542);
and U2643 (N_2643,N_2559,N_2598);
nand U2644 (N_2644,N_2521,N_2580);
nand U2645 (N_2645,N_2551,N_2544);
xnor U2646 (N_2646,N_2503,N_2583);
xnor U2647 (N_2647,N_2514,N_2579);
and U2648 (N_2648,N_2557,N_2530);
and U2649 (N_2649,N_2569,N_2585);
nor U2650 (N_2650,N_2501,N_2507);
xnor U2651 (N_2651,N_2582,N_2523);
and U2652 (N_2652,N_2508,N_2567);
or U2653 (N_2653,N_2510,N_2552);
or U2654 (N_2654,N_2509,N_2559);
and U2655 (N_2655,N_2569,N_2553);
nor U2656 (N_2656,N_2594,N_2517);
nand U2657 (N_2657,N_2597,N_2522);
and U2658 (N_2658,N_2530,N_2598);
xor U2659 (N_2659,N_2508,N_2575);
nor U2660 (N_2660,N_2527,N_2545);
and U2661 (N_2661,N_2536,N_2532);
nor U2662 (N_2662,N_2544,N_2511);
nor U2663 (N_2663,N_2549,N_2578);
xor U2664 (N_2664,N_2526,N_2524);
and U2665 (N_2665,N_2569,N_2502);
or U2666 (N_2666,N_2515,N_2564);
or U2667 (N_2667,N_2540,N_2512);
nand U2668 (N_2668,N_2502,N_2566);
and U2669 (N_2669,N_2560,N_2595);
nor U2670 (N_2670,N_2547,N_2596);
xor U2671 (N_2671,N_2503,N_2501);
nand U2672 (N_2672,N_2590,N_2576);
and U2673 (N_2673,N_2534,N_2550);
nor U2674 (N_2674,N_2572,N_2598);
xor U2675 (N_2675,N_2583,N_2590);
and U2676 (N_2676,N_2529,N_2542);
nand U2677 (N_2677,N_2524,N_2541);
or U2678 (N_2678,N_2555,N_2522);
and U2679 (N_2679,N_2568,N_2500);
xor U2680 (N_2680,N_2564,N_2502);
and U2681 (N_2681,N_2500,N_2588);
or U2682 (N_2682,N_2531,N_2514);
nor U2683 (N_2683,N_2571,N_2534);
or U2684 (N_2684,N_2599,N_2576);
nor U2685 (N_2685,N_2511,N_2518);
xnor U2686 (N_2686,N_2582,N_2500);
or U2687 (N_2687,N_2595,N_2551);
xnor U2688 (N_2688,N_2523,N_2511);
and U2689 (N_2689,N_2561,N_2504);
nand U2690 (N_2690,N_2579,N_2542);
or U2691 (N_2691,N_2571,N_2565);
xnor U2692 (N_2692,N_2572,N_2534);
or U2693 (N_2693,N_2544,N_2539);
and U2694 (N_2694,N_2535,N_2565);
xnor U2695 (N_2695,N_2596,N_2564);
nor U2696 (N_2696,N_2525,N_2591);
nand U2697 (N_2697,N_2516,N_2500);
or U2698 (N_2698,N_2504,N_2598);
nor U2699 (N_2699,N_2513,N_2509);
nor U2700 (N_2700,N_2603,N_2618);
nor U2701 (N_2701,N_2653,N_2691);
nor U2702 (N_2702,N_2664,N_2666);
nand U2703 (N_2703,N_2607,N_2629);
or U2704 (N_2704,N_2628,N_2606);
and U2705 (N_2705,N_2646,N_2651);
nor U2706 (N_2706,N_2695,N_2613);
xor U2707 (N_2707,N_2620,N_2612);
nand U2708 (N_2708,N_2677,N_2640);
xnor U2709 (N_2709,N_2625,N_2604);
nor U2710 (N_2710,N_2616,N_2662);
nand U2711 (N_2711,N_2643,N_2657);
and U2712 (N_2712,N_2619,N_2659);
and U2713 (N_2713,N_2667,N_2661);
nor U2714 (N_2714,N_2631,N_2621);
or U2715 (N_2715,N_2650,N_2673);
nand U2716 (N_2716,N_2637,N_2698);
or U2717 (N_2717,N_2641,N_2647);
xnor U2718 (N_2718,N_2697,N_2622);
nor U2719 (N_2719,N_2670,N_2627);
xor U2720 (N_2720,N_2635,N_2686);
nor U2721 (N_2721,N_2692,N_2672);
nand U2722 (N_2722,N_2674,N_2602);
and U2723 (N_2723,N_2644,N_2699);
nor U2724 (N_2724,N_2648,N_2665);
xnor U2725 (N_2725,N_2668,N_2610);
nor U2726 (N_2726,N_2694,N_2611);
xnor U2727 (N_2727,N_2669,N_2681);
or U2728 (N_2728,N_2636,N_2634);
or U2729 (N_2729,N_2658,N_2601);
nor U2730 (N_2730,N_2671,N_2638);
nand U2731 (N_2731,N_2630,N_2609);
nand U2732 (N_2732,N_2683,N_2688);
nand U2733 (N_2733,N_2687,N_2624);
and U2734 (N_2734,N_2642,N_2684);
nor U2735 (N_2735,N_2614,N_2639);
and U2736 (N_2736,N_2626,N_2645);
nand U2737 (N_2737,N_2690,N_2663);
xor U2738 (N_2738,N_2615,N_2654);
nand U2739 (N_2739,N_2680,N_2682);
xnor U2740 (N_2740,N_2656,N_2679);
or U2741 (N_2741,N_2632,N_2605);
xor U2742 (N_2742,N_2600,N_2693);
nor U2743 (N_2743,N_2649,N_2696);
nand U2744 (N_2744,N_2617,N_2676);
nor U2745 (N_2745,N_2623,N_2655);
or U2746 (N_2746,N_2608,N_2675);
and U2747 (N_2747,N_2678,N_2652);
and U2748 (N_2748,N_2660,N_2689);
xnor U2749 (N_2749,N_2685,N_2633);
nor U2750 (N_2750,N_2640,N_2693);
nor U2751 (N_2751,N_2624,N_2657);
xnor U2752 (N_2752,N_2692,N_2620);
xnor U2753 (N_2753,N_2680,N_2611);
xor U2754 (N_2754,N_2689,N_2670);
nand U2755 (N_2755,N_2606,N_2657);
or U2756 (N_2756,N_2680,N_2642);
nand U2757 (N_2757,N_2688,N_2602);
nor U2758 (N_2758,N_2600,N_2610);
nand U2759 (N_2759,N_2640,N_2656);
xor U2760 (N_2760,N_2643,N_2646);
nand U2761 (N_2761,N_2662,N_2629);
nor U2762 (N_2762,N_2697,N_2673);
or U2763 (N_2763,N_2668,N_2673);
nand U2764 (N_2764,N_2677,N_2610);
nor U2765 (N_2765,N_2645,N_2623);
xnor U2766 (N_2766,N_2634,N_2640);
and U2767 (N_2767,N_2669,N_2646);
or U2768 (N_2768,N_2629,N_2696);
or U2769 (N_2769,N_2680,N_2685);
or U2770 (N_2770,N_2607,N_2699);
xnor U2771 (N_2771,N_2677,N_2603);
or U2772 (N_2772,N_2675,N_2683);
xor U2773 (N_2773,N_2634,N_2661);
xnor U2774 (N_2774,N_2620,N_2652);
or U2775 (N_2775,N_2627,N_2626);
and U2776 (N_2776,N_2660,N_2644);
nand U2777 (N_2777,N_2619,N_2688);
xor U2778 (N_2778,N_2634,N_2695);
nand U2779 (N_2779,N_2627,N_2686);
nor U2780 (N_2780,N_2675,N_2654);
xnor U2781 (N_2781,N_2616,N_2602);
xor U2782 (N_2782,N_2655,N_2645);
nand U2783 (N_2783,N_2602,N_2691);
nand U2784 (N_2784,N_2605,N_2609);
nand U2785 (N_2785,N_2678,N_2672);
and U2786 (N_2786,N_2697,N_2603);
xor U2787 (N_2787,N_2654,N_2646);
nand U2788 (N_2788,N_2696,N_2681);
nor U2789 (N_2789,N_2633,N_2617);
or U2790 (N_2790,N_2621,N_2654);
nor U2791 (N_2791,N_2656,N_2644);
xor U2792 (N_2792,N_2607,N_2614);
and U2793 (N_2793,N_2621,N_2694);
or U2794 (N_2794,N_2667,N_2645);
or U2795 (N_2795,N_2601,N_2647);
xnor U2796 (N_2796,N_2643,N_2651);
xor U2797 (N_2797,N_2615,N_2652);
or U2798 (N_2798,N_2642,N_2696);
and U2799 (N_2799,N_2698,N_2639);
xor U2800 (N_2800,N_2783,N_2799);
and U2801 (N_2801,N_2780,N_2795);
or U2802 (N_2802,N_2786,N_2743);
nor U2803 (N_2803,N_2791,N_2784);
and U2804 (N_2804,N_2765,N_2773);
nor U2805 (N_2805,N_2782,N_2712);
nor U2806 (N_2806,N_2719,N_2710);
xnor U2807 (N_2807,N_2798,N_2749);
nor U2808 (N_2808,N_2767,N_2769);
nand U2809 (N_2809,N_2716,N_2755);
xnor U2810 (N_2810,N_2771,N_2731);
nand U2811 (N_2811,N_2779,N_2790);
nand U2812 (N_2812,N_2747,N_2729);
and U2813 (N_2813,N_2788,N_2733);
nand U2814 (N_2814,N_2754,N_2726);
and U2815 (N_2815,N_2761,N_2722);
nor U2816 (N_2816,N_2715,N_2759);
or U2817 (N_2817,N_2796,N_2713);
nand U2818 (N_2818,N_2725,N_2775);
xor U2819 (N_2819,N_2708,N_2762);
nor U2820 (N_2820,N_2736,N_2777);
nor U2821 (N_2821,N_2739,N_2723);
nand U2822 (N_2822,N_2728,N_2707);
nand U2823 (N_2823,N_2721,N_2787);
or U2824 (N_2824,N_2756,N_2700);
nor U2825 (N_2825,N_2738,N_2770);
or U2826 (N_2826,N_2752,N_2793);
xnor U2827 (N_2827,N_2744,N_2742);
nor U2828 (N_2828,N_2732,N_2704);
nand U2829 (N_2829,N_2717,N_2760);
and U2830 (N_2830,N_2711,N_2737);
xor U2831 (N_2831,N_2718,N_2789);
and U2832 (N_2832,N_2776,N_2785);
nand U2833 (N_2833,N_2764,N_2763);
or U2834 (N_2834,N_2706,N_2781);
xor U2835 (N_2835,N_2757,N_2772);
xnor U2836 (N_2836,N_2746,N_2797);
nand U2837 (N_2837,N_2745,N_2766);
nand U2838 (N_2838,N_2774,N_2778);
nand U2839 (N_2839,N_2703,N_2702);
nor U2840 (N_2840,N_2720,N_2724);
nor U2841 (N_2841,N_2701,N_2714);
or U2842 (N_2842,N_2705,N_2751);
and U2843 (N_2843,N_2750,N_2741);
or U2844 (N_2844,N_2735,N_2748);
nand U2845 (N_2845,N_2709,N_2792);
or U2846 (N_2846,N_2753,N_2794);
nor U2847 (N_2847,N_2730,N_2727);
nand U2848 (N_2848,N_2734,N_2768);
nand U2849 (N_2849,N_2740,N_2758);
nor U2850 (N_2850,N_2713,N_2737);
or U2851 (N_2851,N_2716,N_2743);
nand U2852 (N_2852,N_2709,N_2719);
or U2853 (N_2853,N_2706,N_2767);
or U2854 (N_2854,N_2795,N_2728);
nand U2855 (N_2855,N_2707,N_2790);
or U2856 (N_2856,N_2791,N_2703);
or U2857 (N_2857,N_2733,N_2722);
or U2858 (N_2858,N_2741,N_2749);
nor U2859 (N_2859,N_2794,N_2780);
nand U2860 (N_2860,N_2726,N_2779);
xor U2861 (N_2861,N_2701,N_2700);
nor U2862 (N_2862,N_2749,N_2721);
and U2863 (N_2863,N_2774,N_2794);
or U2864 (N_2864,N_2702,N_2776);
and U2865 (N_2865,N_2781,N_2744);
and U2866 (N_2866,N_2746,N_2780);
nand U2867 (N_2867,N_2748,N_2796);
and U2868 (N_2868,N_2756,N_2733);
xor U2869 (N_2869,N_2720,N_2751);
or U2870 (N_2870,N_2742,N_2772);
and U2871 (N_2871,N_2786,N_2748);
and U2872 (N_2872,N_2745,N_2728);
or U2873 (N_2873,N_2757,N_2767);
or U2874 (N_2874,N_2771,N_2782);
nand U2875 (N_2875,N_2789,N_2761);
or U2876 (N_2876,N_2714,N_2790);
nand U2877 (N_2877,N_2762,N_2723);
nor U2878 (N_2878,N_2763,N_2782);
xnor U2879 (N_2879,N_2757,N_2737);
and U2880 (N_2880,N_2729,N_2745);
xnor U2881 (N_2881,N_2737,N_2729);
or U2882 (N_2882,N_2792,N_2798);
and U2883 (N_2883,N_2725,N_2755);
xor U2884 (N_2884,N_2784,N_2770);
xor U2885 (N_2885,N_2716,N_2764);
nand U2886 (N_2886,N_2750,N_2746);
xor U2887 (N_2887,N_2725,N_2736);
and U2888 (N_2888,N_2732,N_2711);
xnor U2889 (N_2889,N_2774,N_2782);
xnor U2890 (N_2890,N_2710,N_2740);
nor U2891 (N_2891,N_2796,N_2712);
and U2892 (N_2892,N_2725,N_2781);
xnor U2893 (N_2893,N_2783,N_2725);
and U2894 (N_2894,N_2729,N_2785);
or U2895 (N_2895,N_2741,N_2723);
xnor U2896 (N_2896,N_2779,N_2738);
xnor U2897 (N_2897,N_2789,N_2705);
xor U2898 (N_2898,N_2747,N_2762);
and U2899 (N_2899,N_2788,N_2765);
nand U2900 (N_2900,N_2883,N_2811);
nor U2901 (N_2901,N_2837,N_2830);
and U2902 (N_2902,N_2893,N_2880);
and U2903 (N_2903,N_2876,N_2864);
nor U2904 (N_2904,N_2873,N_2871);
xnor U2905 (N_2905,N_2890,N_2808);
nand U2906 (N_2906,N_2833,N_2882);
or U2907 (N_2907,N_2848,N_2889);
and U2908 (N_2908,N_2807,N_2828);
nor U2909 (N_2909,N_2835,N_2817);
xor U2910 (N_2910,N_2868,N_2847);
xor U2911 (N_2911,N_2809,N_2822);
and U2912 (N_2912,N_2821,N_2800);
and U2913 (N_2913,N_2852,N_2874);
xnor U2914 (N_2914,N_2849,N_2899);
and U2915 (N_2915,N_2801,N_2856);
nor U2916 (N_2916,N_2854,N_2881);
or U2917 (N_2917,N_2832,N_2831);
or U2918 (N_2918,N_2841,N_2869);
nor U2919 (N_2919,N_2812,N_2887);
nor U2920 (N_2920,N_2898,N_2804);
and U2921 (N_2921,N_2894,N_2838);
xnor U2922 (N_2922,N_2820,N_2884);
nor U2923 (N_2923,N_2862,N_2863);
nand U2924 (N_2924,N_2860,N_2896);
nand U2925 (N_2925,N_2813,N_2844);
xnor U2926 (N_2926,N_2853,N_2840);
xor U2927 (N_2927,N_2845,N_2810);
and U2928 (N_2928,N_2875,N_2805);
and U2929 (N_2929,N_2826,N_2892);
and U2930 (N_2930,N_2859,N_2865);
xor U2931 (N_2931,N_2867,N_2885);
nor U2932 (N_2932,N_2877,N_2866);
or U2933 (N_2933,N_2836,N_2897);
nand U2934 (N_2934,N_2803,N_2823);
nor U2935 (N_2935,N_2814,N_2886);
xnor U2936 (N_2936,N_2829,N_2846);
xor U2937 (N_2937,N_2855,N_2818);
and U2938 (N_2938,N_2870,N_2861);
nor U2939 (N_2939,N_2843,N_2872);
nor U2940 (N_2940,N_2827,N_2825);
xnor U2941 (N_2941,N_2850,N_2857);
and U2942 (N_2942,N_2824,N_2839);
xnor U2943 (N_2943,N_2816,N_2842);
and U2944 (N_2944,N_2806,N_2815);
xnor U2945 (N_2945,N_2802,N_2891);
or U2946 (N_2946,N_2895,N_2851);
nor U2947 (N_2947,N_2858,N_2834);
nor U2948 (N_2948,N_2879,N_2888);
xnor U2949 (N_2949,N_2878,N_2819);
xor U2950 (N_2950,N_2847,N_2887);
and U2951 (N_2951,N_2857,N_2845);
nor U2952 (N_2952,N_2819,N_2887);
xor U2953 (N_2953,N_2894,N_2859);
nor U2954 (N_2954,N_2861,N_2855);
or U2955 (N_2955,N_2873,N_2819);
nor U2956 (N_2956,N_2899,N_2840);
nor U2957 (N_2957,N_2869,N_2826);
nor U2958 (N_2958,N_2812,N_2822);
nor U2959 (N_2959,N_2880,N_2881);
or U2960 (N_2960,N_2891,N_2878);
xor U2961 (N_2961,N_2889,N_2870);
nor U2962 (N_2962,N_2823,N_2862);
xnor U2963 (N_2963,N_2887,N_2852);
nand U2964 (N_2964,N_2882,N_2819);
or U2965 (N_2965,N_2807,N_2806);
nand U2966 (N_2966,N_2861,N_2865);
nor U2967 (N_2967,N_2890,N_2831);
or U2968 (N_2968,N_2879,N_2873);
nand U2969 (N_2969,N_2829,N_2813);
or U2970 (N_2970,N_2867,N_2815);
nand U2971 (N_2971,N_2841,N_2826);
nand U2972 (N_2972,N_2832,N_2809);
nand U2973 (N_2973,N_2810,N_2878);
and U2974 (N_2974,N_2810,N_2887);
or U2975 (N_2975,N_2841,N_2853);
or U2976 (N_2976,N_2884,N_2841);
nor U2977 (N_2977,N_2877,N_2870);
nand U2978 (N_2978,N_2884,N_2816);
nor U2979 (N_2979,N_2800,N_2869);
xnor U2980 (N_2980,N_2823,N_2822);
or U2981 (N_2981,N_2835,N_2877);
and U2982 (N_2982,N_2873,N_2899);
or U2983 (N_2983,N_2812,N_2813);
xor U2984 (N_2984,N_2896,N_2841);
or U2985 (N_2985,N_2857,N_2802);
and U2986 (N_2986,N_2832,N_2883);
xnor U2987 (N_2987,N_2882,N_2806);
and U2988 (N_2988,N_2867,N_2835);
nand U2989 (N_2989,N_2821,N_2820);
nand U2990 (N_2990,N_2857,N_2800);
nand U2991 (N_2991,N_2883,N_2880);
xnor U2992 (N_2992,N_2887,N_2873);
and U2993 (N_2993,N_2815,N_2860);
nand U2994 (N_2994,N_2895,N_2847);
nor U2995 (N_2995,N_2810,N_2803);
or U2996 (N_2996,N_2874,N_2846);
nor U2997 (N_2997,N_2851,N_2845);
and U2998 (N_2998,N_2851,N_2814);
xor U2999 (N_2999,N_2856,N_2823);
or UO_0 (O_0,N_2905,N_2929);
xnor UO_1 (O_1,N_2901,N_2909);
nand UO_2 (O_2,N_2975,N_2996);
nand UO_3 (O_3,N_2959,N_2930);
xnor UO_4 (O_4,N_2917,N_2907);
nor UO_5 (O_5,N_2953,N_2919);
and UO_6 (O_6,N_2967,N_2983);
and UO_7 (O_7,N_2979,N_2960);
or UO_8 (O_8,N_2922,N_2977);
and UO_9 (O_9,N_2927,N_2980);
and UO_10 (O_10,N_2902,N_2926);
xnor UO_11 (O_11,N_2954,N_2969);
nand UO_12 (O_12,N_2987,N_2921);
and UO_13 (O_13,N_2956,N_2971);
nand UO_14 (O_14,N_2952,N_2940);
nand UO_15 (O_15,N_2900,N_2994);
nand UO_16 (O_16,N_2986,N_2957);
and UO_17 (O_17,N_2992,N_2949);
xnor UO_18 (O_18,N_2928,N_2906);
xnor UO_19 (O_19,N_2934,N_2976);
xor UO_20 (O_20,N_2963,N_2989);
nand UO_21 (O_21,N_2942,N_2965);
and UO_22 (O_22,N_2908,N_2974);
and UO_23 (O_23,N_2933,N_2970);
or UO_24 (O_24,N_2903,N_2951);
nor UO_25 (O_25,N_2925,N_2972);
nor UO_26 (O_26,N_2932,N_2950);
nor UO_27 (O_27,N_2973,N_2945);
nand UO_28 (O_28,N_2944,N_2998);
and UO_29 (O_29,N_2937,N_2948);
or UO_30 (O_30,N_2914,N_2985);
or UO_31 (O_31,N_2913,N_2924);
or UO_32 (O_32,N_2964,N_2968);
xor UO_33 (O_33,N_2993,N_2910);
nand UO_34 (O_34,N_2946,N_2911);
xnor UO_35 (O_35,N_2904,N_2938);
nand UO_36 (O_36,N_2931,N_2936);
nor UO_37 (O_37,N_2995,N_2982);
nor UO_38 (O_38,N_2939,N_2981);
nand UO_39 (O_39,N_2958,N_2961);
or UO_40 (O_40,N_2935,N_2966);
nor UO_41 (O_41,N_2988,N_2990);
xor UO_42 (O_42,N_2912,N_2920);
and UO_43 (O_43,N_2943,N_2941);
nand UO_44 (O_44,N_2991,N_2955);
or UO_45 (O_45,N_2947,N_2978);
nor UO_46 (O_46,N_2915,N_2999);
and UO_47 (O_47,N_2916,N_2997);
nor UO_48 (O_48,N_2984,N_2918);
xnor UO_49 (O_49,N_2962,N_2923);
xor UO_50 (O_50,N_2966,N_2939);
nor UO_51 (O_51,N_2989,N_2974);
or UO_52 (O_52,N_2946,N_2957);
nor UO_53 (O_53,N_2994,N_2965);
xnor UO_54 (O_54,N_2920,N_2900);
and UO_55 (O_55,N_2936,N_2995);
nand UO_56 (O_56,N_2932,N_2951);
xor UO_57 (O_57,N_2943,N_2989);
nand UO_58 (O_58,N_2905,N_2972);
xnor UO_59 (O_59,N_2957,N_2926);
nand UO_60 (O_60,N_2967,N_2978);
nor UO_61 (O_61,N_2940,N_2900);
xor UO_62 (O_62,N_2930,N_2922);
and UO_63 (O_63,N_2909,N_2932);
nor UO_64 (O_64,N_2949,N_2979);
and UO_65 (O_65,N_2997,N_2976);
nor UO_66 (O_66,N_2972,N_2998);
or UO_67 (O_67,N_2908,N_2914);
nor UO_68 (O_68,N_2993,N_2949);
nand UO_69 (O_69,N_2939,N_2940);
or UO_70 (O_70,N_2966,N_2924);
and UO_71 (O_71,N_2995,N_2905);
and UO_72 (O_72,N_2948,N_2970);
xnor UO_73 (O_73,N_2951,N_2980);
and UO_74 (O_74,N_2919,N_2932);
or UO_75 (O_75,N_2984,N_2971);
nor UO_76 (O_76,N_2949,N_2990);
and UO_77 (O_77,N_2904,N_2902);
nor UO_78 (O_78,N_2990,N_2937);
and UO_79 (O_79,N_2975,N_2911);
nor UO_80 (O_80,N_2999,N_2913);
xnor UO_81 (O_81,N_2958,N_2993);
xnor UO_82 (O_82,N_2994,N_2991);
and UO_83 (O_83,N_2961,N_2983);
nor UO_84 (O_84,N_2967,N_2972);
xor UO_85 (O_85,N_2909,N_2941);
nand UO_86 (O_86,N_2920,N_2926);
nand UO_87 (O_87,N_2949,N_2930);
or UO_88 (O_88,N_2935,N_2995);
and UO_89 (O_89,N_2900,N_2943);
xor UO_90 (O_90,N_2954,N_2914);
or UO_91 (O_91,N_2961,N_2930);
and UO_92 (O_92,N_2951,N_2985);
or UO_93 (O_93,N_2916,N_2933);
nor UO_94 (O_94,N_2929,N_2961);
or UO_95 (O_95,N_2944,N_2937);
nand UO_96 (O_96,N_2905,N_2998);
nand UO_97 (O_97,N_2943,N_2909);
xor UO_98 (O_98,N_2916,N_2968);
nand UO_99 (O_99,N_2919,N_2978);
or UO_100 (O_100,N_2908,N_2941);
and UO_101 (O_101,N_2973,N_2971);
and UO_102 (O_102,N_2977,N_2995);
xnor UO_103 (O_103,N_2920,N_2966);
nand UO_104 (O_104,N_2932,N_2961);
or UO_105 (O_105,N_2919,N_2926);
or UO_106 (O_106,N_2909,N_2949);
and UO_107 (O_107,N_2919,N_2992);
nor UO_108 (O_108,N_2918,N_2917);
or UO_109 (O_109,N_2989,N_2970);
xnor UO_110 (O_110,N_2976,N_2950);
nor UO_111 (O_111,N_2928,N_2997);
xnor UO_112 (O_112,N_2904,N_2909);
nor UO_113 (O_113,N_2905,N_2979);
and UO_114 (O_114,N_2955,N_2906);
and UO_115 (O_115,N_2932,N_2980);
nor UO_116 (O_116,N_2980,N_2941);
nand UO_117 (O_117,N_2972,N_2933);
and UO_118 (O_118,N_2938,N_2962);
or UO_119 (O_119,N_2941,N_2976);
or UO_120 (O_120,N_2981,N_2962);
xnor UO_121 (O_121,N_2956,N_2901);
nand UO_122 (O_122,N_2992,N_2915);
and UO_123 (O_123,N_2971,N_2920);
nand UO_124 (O_124,N_2995,N_2943);
xnor UO_125 (O_125,N_2957,N_2976);
xnor UO_126 (O_126,N_2957,N_2960);
nor UO_127 (O_127,N_2917,N_2915);
or UO_128 (O_128,N_2935,N_2938);
nand UO_129 (O_129,N_2918,N_2994);
xor UO_130 (O_130,N_2926,N_2996);
xor UO_131 (O_131,N_2948,N_2935);
and UO_132 (O_132,N_2967,N_2935);
nor UO_133 (O_133,N_2951,N_2983);
nor UO_134 (O_134,N_2910,N_2926);
nand UO_135 (O_135,N_2908,N_2910);
nand UO_136 (O_136,N_2965,N_2944);
or UO_137 (O_137,N_2911,N_2945);
nand UO_138 (O_138,N_2995,N_2918);
and UO_139 (O_139,N_2986,N_2947);
xnor UO_140 (O_140,N_2928,N_2969);
nor UO_141 (O_141,N_2964,N_2905);
and UO_142 (O_142,N_2948,N_2946);
nand UO_143 (O_143,N_2930,N_2982);
and UO_144 (O_144,N_2963,N_2996);
xor UO_145 (O_145,N_2952,N_2917);
nand UO_146 (O_146,N_2916,N_2905);
nand UO_147 (O_147,N_2912,N_2932);
nor UO_148 (O_148,N_2979,N_2986);
nand UO_149 (O_149,N_2993,N_2934);
or UO_150 (O_150,N_2913,N_2939);
xor UO_151 (O_151,N_2911,N_2996);
and UO_152 (O_152,N_2991,N_2907);
and UO_153 (O_153,N_2959,N_2911);
and UO_154 (O_154,N_2906,N_2915);
xnor UO_155 (O_155,N_2970,N_2936);
nand UO_156 (O_156,N_2923,N_2998);
xnor UO_157 (O_157,N_2977,N_2946);
xor UO_158 (O_158,N_2970,N_2952);
nor UO_159 (O_159,N_2927,N_2944);
nor UO_160 (O_160,N_2900,N_2908);
nor UO_161 (O_161,N_2907,N_2955);
nor UO_162 (O_162,N_2996,N_2995);
or UO_163 (O_163,N_2933,N_2923);
nand UO_164 (O_164,N_2991,N_2903);
nor UO_165 (O_165,N_2973,N_2988);
and UO_166 (O_166,N_2992,N_2972);
and UO_167 (O_167,N_2988,N_2984);
nor UO_168 (O_168,N_2973,N_2920);
nor UO_169 (O_169,N_2935,N_2922);
xnor UO_170 (O_170,N_2976,N_2998);
nand UO_171 (O_171,N_2958,N_2926);
xor UO_172 (O_172,N_2969,N_2943);
nand UO_173 (O_173,N_2907,N_2982);
xnor UO_174 (O_174,N_2970,N_2969);
xnor UO_175 (O_175,N_2923,N_2903);
xor UO_176 (O_176,N_2950,N_2931);
nand UO_177 (O_177,N_2992,N_2954);
xor UO_178 (O_178,N_2999,N_2974);
and UO_179 (O_179,N_2975,N_2943);
or UO_180 (O_180,N_2997,N_2922);
xnor UO_181 (O_181,N_2994,N_2975);
or UO_182 (O_182,N_2932,N_2963);
xnor UO_183 (O_183,N_2944,N_2915);
xnor UO_184 (O_184,N_2958,N_2904);
or UO_185 (O_185,N_2926,N_2929);
or UO_186 (O_186,N_2941,N_2985);
xor UO_187 (O_187,N_2974,N_2914);
nand UO_188 (O_188,N_2976,N_2937);
nand UO_189 (O_189,N_2972,N_2955);
xnor UO_190 (O_190,N_2956,N_2907);
nor UO_191 (O_191,N_2942,N_2979);
and UO_192 (O_192,N_2961,N_2939);
and UO_193 (O_193,N_2966,N_2952);
or UO_194 (O_194,N_2916,N_2975);
xnor UO_195 (O_195,N_2909,N_2953);
nand UO_196 (O_196,N_2991,N_2962);
and UO_197 (O_197,N_2990,N_2992);
or UO_198 (O_198,N_2990,N_2923);
and UO_199 (O_199,N_2953,N_2963);
or UO_200 (O_200,N_2957,N_2936);
or UO_201 (O_201,N_2970,N_2991);
and UO_202 (O_202,N_2979,N_2946);
nor UO_203 (O_203,N_2926,N_2977);
xnor UO_204 (O_204,N_2966,N_2979);
and UO_205 (O_205,N_2935,N_2973);
or UO_206 (O_206,N_2949,N_2939);
xor UO_207 (O_207,N_2913,N_2992);
nand UO_208 (O_208,N_2939,N_2921);
xor UO_209 (O_209,N_2933,N_2993);
nand UO_210 (O_210,N_2912,N_2911);
or UO_211 (O_211,N_2921,N_2961);
nor UO_212 (O_212,N_2982,N_2921);
or UO_213 (O_213,N_2937,N_2908);
and UO_214 (O_214,N_2986,N_2919);
nand UO_215 (O_215,N_2987,N_2991);
nor UO_216 (O_216,N_2936,N_2952);
or UO_217 (O_217,N_2950,N_2974);
nor UO_218 (O_218,N_2996,N_2964);
or UO_219 (O_219,N_2965,N_2941);
nor UO_220 (O_220,N_2935,N_2961);
xor UO_221 (O_221,N_2910,N_2918);
xnor UO_222 (O_222,N_2907,N_2962);
nand UO_223 (O_223,N_2905,N_2944);
nand UO_224 (O_224,N_2986,N_2933);
nor UO_225 (O_225,N_2976,N_2940);
and UO_226 (O_226,N_2917,N_2930);
nand UO_227 (O_227,N_2905,N_2974);
xor UO_228 (O_228,N_2978,N_2949);
nand UO_229 (O_229,N_2959,N_2919);
nor UO_230 (O_230,N_2989,N_2956);
nand UO_231 (O_231,N_2948,N_2920);
and UO_232 (O_232,N_2930,N_2957);
and UO_233 (O_233,N_2938,N_2983);
nor UO_234 (O_234,N_2948,N_2996);
and UO_235 (O_235,N_2975,N_2959);
xor UO_236 (O_236,N_2923,N_2996);
nor UO_237 (O_237,N_2911,N_2954);
or UO_238 (O_238,N_2968,N_2908);
nand UO_239 (O_239,N_2923,N_2939);
nand UO_240 (O_240,N_2906,N_2975);
or UO_241 (O_241,N_2952,N_2912);
and UO_242 (O_242,N_2959,N_2944);
xor UO_243 (O_243,N_2903,N_2947);
xnor UO_244 (O_244,N_2954,N_2958);
nand UO_245 (O_245,N_2928,N_2908);
nand UO_246 (O_246,N_2993,N_2928);
nor UO_247 (O_247,N_2917,N_2953);
xor UO_248 (O_248,N_2972,N_2923);
and UO_249 (O_249,N_2945,N_2944);
nand UO_250 (O_250,N_2976,N_2902);
nand UO_251 (O_251,N_2937,N_2974);
xnor UO_252 (O_252,N_2900,N_2975);
nor UO_253 (O_253,N_2980,N_2949);
or UO_254 (O_254,N_2994,N_2908);
or UO_255 (O_255,N_2954,N_2967);
and UO_256 (O_256,N_2954,N_2937);
nand UO_257 (O_257,N_2926,N_2965);
nand UO_258 (O_258,N_2927,N_2983);
xnor UO_259 (O_259,N_2962,N_2975);
xor UO_260 (O_260,N_2992,N_2973);
nor UO_261 (O_261,N_2957,N_2968);
nor UO_262 (O_262,N_2940,N_2922);
or UO_263 (O_263,N_2972,N_2929);
xor UO_264 (O_264,N_2907,N_2943);
and UO_265 (O_265,N_2974,N_2941);
and UO_266 (O_266,N_2920,N_2908);
and UO_267 (O_267,N_2933,N_2940);
nand UO_268 (O_268,N_2928,N_2903);
xnor UO_269 (O_269,N_2916,N_2993);
nor UO_270 (O_270,N_2906,N_2963);
and UO_271 (O_271,N_2986,N_2914);
nor UO_272 (O_272,N_2914,N_2915);
xor UO_273 (O_273,N_2936,N_2942);
or UO_274 (O_274,N_2907,N_2933);
and UO_275 (O_275,N_2921,N_2927);
nand UO_276 (O_276,N_2996,N_2931);
nor UO_277 (O_277,N_2915,N_2975);
and UO_278 (O_278,N_2959,N_2963);
nand UO_279 (O_279,N_2908,N_2956);
nor UO_280 (O_280,N_2986,N_2928);
or UO_281 (O_281,N_2949,N_2920);
and UO_282 (O_282,N_2999,N_2927);
xnor UO_283 (O_283,N_2915,N_2983);
or UO_284 (O_284,N_2988,N_2906);
nand UO_285 (O_285,N_2913,N_2975);
and UO_286 (O_286,N_2939,N_2978);
xnor UO_287 (O_287,N_2977,N_2912);
and UO_288 (O_288,N_2953,N_2991);
xor UO_289 (O_289,N_2969,N_2989);
or UO_290 (O_290,N_2930,N_2956);
nor UO_291 (O_291,N_2928,N_2999);
xnor UO_292 (O_292,N_2931,N_2956);
or UO_293 (O_293,N_2981,N_2960);
xor UO_294 (O_294,N_2973,N_2982);
or UO_295 (O_295,N_2973,N_2991);
xnor UO_296 (O_296,N_2928,N_2937);
nand UO_297 (O_297,N_2940,N_2960);
nor UO_298 (O_298,N_2904,N_2999);
nor UO_299 (O_299,N_2942,N_2957);
xor UO_300 (O_300,N_2965,N_2902);
nor UO_301 (O_301,N_2907,N_2912);
or UO_302 (O_302,N_2983,N_2931);
and UO_303 (O_303,N_2964,N_2929);
nand UO_304 (O_304,N_2945,N_2910);
nand UO_305 (O_305,N_2939,N_2970);
xor UO_306 (O_306,N_2903,N_2956);
nand UO_307 (O_307,N_2994,N_2974);
nor UO_308 (O_308,N_2907,N_2971);
or UO_309 (O_309,N_2910,N_2930);
or UO_310 (O_310,N_2959,N_2949);
and UO_311 (O_311,N_2971,N_2948);
and UO_312 (O_312,N_2977,N_2998);
nand UO_313 (O_313,N_2905,N_2984);
nor UO_314 (O_314,N_2958,N_2919);
nand UO_315 (O_315,N_2996,N_2935);
nand UO_316 (O_316,N_2984,N_2968);
xor UO_317 (O_317,N_2982,N_2962);
and UO_318 (O_318,N_2953,N_2935);
nor UO_319 (O_319,N_2975,N_2926);
nand UO_320 (O_320,N_2904,N_2995);
xnor UO_321 (O_321,N_2930,N_2989);
or UO_322 (O_322,N_2991,N_2983);
and UO_323 (O_323,N_2957,N_2901);
and UO_324 (O_324,N_2903,N_2996);
or UO_325 (O_325,N_2902,N_2949);
or UO_326 (O_326,N_2967,N_2925);
or UO_327 (O_327,N_2937,N_2900);
xor UO_328 (O_328,N_2914,N_2924);
xor UO_329 (O_329,N_2910,N_2923);
or UO_330 (O_330,N_2939,N_2955);
nand UO_331 (O_331,N_2922,N_2923);
xor UO_332 (O_332,N_2954,N_2999);
or UO_333 (O_333,N_2911,N_2918);
nor UO_334 (O_334,N_2954,N_2924);
nand UO_335 (O_335,N_2997,N_2996);
and UO_336 (O_336,N_2941,N_2900);
xnor UO_337 (O_337,N_2944,N_2948);
or UO_338 (O_338,N_2991,N_2948);
and UO_339 (O_339,N_2955,N_2979);
or UO_340 (O_340,N_2973,N_2925);
nor UO_341 (O_341,N_2984,N_2976);
or UO_342 (O_342,N_2940,N_2953);
nor UO_343 (O_343,N_2990,N_2910);
nor UO_344 (O_344,N_2947,N_2990);
nand UO_345 (O_345,N_2912,N_2988);
xor UO_346 (O_346,N_2980,N_2989);
and UO_347 (O_347,N_2986,N_2943);
nand UO_348 (O_348,N_2918,N_2947);
nand UO_349 (O_349,N_2985,N_2946);
nor UO_350 (O_350,N_2990,N_2979);
xor UO_351 (O_351,N_2975,N_2968);
xnor UO_352 (O_352,N_2907,N_2986);
and UO_353 (O_353,N_2906,N_2965);
or UO_354 (O_354,N_2926,N_2915);
and UO_355 (O_355,N_2968,N_2976);
xnor UO_356 (O_356,N_2962,N_2955);
or UO_357 (O_357,N_2923,N_2955);
and UO_358 (O_358,N_2974,N_2971);
nor UO_359 (O_359,N_2982,N_2999);
and UO_360 (O_360,N_2939,N_2931);
nor UO_361 (O_361,N_2916,N_2917);
nand UO_362 (O_362,N_2921,N_2963);
xor UO_363 (O_363,N_2989,N_2944);
and UO_364 (O_364,N_2962,N_2946);
or UO_365 (O_365,N_2966,N_2932);
nand UO_366 (O_366,N_2977,N_2909);
nand UO_367 (O_367,N_2992,N_2993);
nor UO_368 (O_368,N_2995,N_2975);
or UO_369 (O_369,N_2939,N_2914);
and UO_370 (O_370,N_2984,N_2983);
nor UO_371 (O_371,N_2903,N_2981);
xor UO_372 (O_372,N_2939,N_2936);
xnor UO_373 (O_373,N_2992,N_2938);
or UO_374 (O_374,N_2953,N_2913);
nand UO_375 (O_375,N_2927,N_2905);
nor UO_376 (O_376,N_2945,N_2962);
nand UO_377 (O_377,N_2905,N_2923);
nand UO_378 (O_378,N_2990,N_2939);
nand UO_379 (O_379,N_2997,N_2927);
xnor UO_380 (O_380,N_2922,N_2951);
nand UO_381 (O_381,N_2901,N_2986);
or UO_382 (O_382,N_2942,N_2953);
or UO_383 (O_383,N_2923,N_2924);
nand UO_384 (O_384,N_2995,N_2979);
and UO_385 (O_385,N_2996,N_2927);
and UO_386 (O_386,N_2918,N_2921);
or UO_387 (O_387,N_2964,N_2998);
or UO_388 (O_388,N_2995,N_2903);
nand UO_389 (O_389,N_2948,N_2951);
nor UO_390 (O_390,N_2968,N_2982);
nor UO_391 (O_391,N_2996,N_2970);
nor UO_392 (O_392,N_2914,N_2988);
nor UO_393 (O_393,N_2998,N_2914);
nand UO_394 (O_394,N_2908,N_2921);
xnor UO_395 (O_395,N_2925,N_2928);
xor UO_396 (O_396,N_2952,N_2923);
or UO_397 (O_397,N_2987,N_2940);
and UO_398 (O_398,N_2995,N_2990);
or UO_399 (O_399,N_2989,N_2934);
xor UO_400 (O_400,N_2942,N_2981);
or UO_401 (O_401,N_2998,N_2963);
or UO_402 (O_402,N_2993,N_2923);
xnor UO_403 (O_403,N_2973,N_2977);
xor UO_404 (O_404,N_2959,N_2953);
and UO_405 (O_405,N_2994,N_2972);
xnor UO_406 (O_406,N_2968,N_2921);
nor UO_407 (O_407,N_2996,N_2934);
and UO_408 (O_408,N_2964,N_2937);
and UO_409 (O_409,N_2933,N_2908);
nand UO_410 (O_410,N_2988,N_2962);
nand UO_411 (O_411,N_2968,N_2972);
or UO_412 (O_412,N_2904,N_2990);
xor UO_413 (O_413,N_2918,N_2932);
nand UO_414 (O_414,N_2981,N_2922);
nor UO_415 (O_415,N_2956,N_2934);
xnor UO_416 (O_416,N_2983,N_2977);
xnor UO_417 (O_417,N_2944,N_2951);
xor UO_418 (O_418,N_2948,N_2997);
xor UO_419 (O_419,N_2921,N_2957);
or UO_420 (O_420,N_2938,N_2916);
nor UO_421 (O_421,N_2967,N_2975);
nand UO_422 (O_422,N_2970,N_2906);
nand UO_423 (O_423,N_2993,N_2924);
or UO_424 (O_424,N_2941,N_2945);
xnor UO_425 (O_425,N_2985,N_2938);
and UO_426 (O_426,N_2926,N_2993);
or UO_427 (O_427,N_2992,N_2965);
nand UO_428 (O_428,N_2948,N_2968);
xnor UO_429 (O_429,N_2991,N_2922);
nand UO_430 (O_430,N_2931,N_2972);
nor UO_431 (O_431,N_2912,N_2931);
nor UO_432 (O_432,N_2940,N_2928);
and UO_433 (O_433,N_2928,N_2943);
nand UO_434 (O_434,N_2920,N_2997);
nor UO_435 (O_435,N_2974,N_2903);
and UO_436 (O_436,N_2933,N_2942);
and UO_437 (O_437,N_2946,N_2968);
or UO_438 (O_438,N_2928,N_2995);
and UO_439 (O_439,N_2984,N_2904);
nor UO_440 (O_440,N_2955,N_2965);
or UO_441 (O_441,N_2999,N_2977);
nor UO_442 (O_442,N_2928,N_2952);
nand UO_443 (O_443,N_2907,N_2904);
xnor UO_444 (O_444,N_2935,N_2903);
or UO_445 (O_445,N_2990,N_2927);
xor UO_446 (O_446,N_2925,N_2905);
and UO_447 (O_447,N_2930,N_2945);
and UO_448 (O_448,N_2977,N_2957);
nor UO_449 (O_449,N_2909,N_2908);
xor UO_450 (O_450,N_2934,N_2929);
xnor UO_451 (O_451,N_2982,N_2983);
nor UO_452 (O_452,N_2923,N_2986);
xor UO_453 (O_453,N_2986,N_2977);
xnor UO_454 (O_454,N_2908,N_2943);
nor UO_455 (O_455,N_2938,N_2973);
or UO_456 (O_456,N_2943,N_2982);
and UO_457 (O_457,N_2993,N_2904);
nor UO_458 (O_458,N_2934,N_2901);
nor UO_459 (O_459,N_2929,N_2986);
nand UO_460 (O_460,N_2901,N_2984);
or UO_461 (O_461,N_2932,N_2983);
nand UO_462 (O_462,N_2961,N_2986);
nor UO_463 (O_463,N_2942,N_2996);
nand UO_464 (O_464,N_2954,N_2951);
nor UO_465 (O_465,N_2943,N_2971);
and UO_466 (O_466,N_2982,N_2960);
xor UO_467 (O_467,N_2925,N_2982);
xnor UO_468 (O_468,N_2947,N_2987);
nand UO_469 (O_469,N_2983,N_2917);
nand UO_470 (O_470,N_2929,N_2953);
or UO_471 (O_471,N_2970,N_2965);
or UO_472 (O_472,N_2911,N_2933);
xnor UO_473 (O_473,N_2932,N_2946);
and UO_474 (O_474,N_2909,N_2994);
nor UO_475 (O_475,N_2981,N_2907);
xnor UO_476 (O_476,N_2927,N_2918);
nor UO_477 (O_477,N_2928,N_2950);
nand UO_478 (O_478,N_2910,N_2946);
xnor UO_479 (O_479,N_2922,N_2988);
and UO_480 (O_480,N_2906,N_2949);
nand UO_481 (O_481,N_2987,N_2949);
xor UO_482 (O_482,N_2909,N_2933);
nor UO_483 (O_483,N_2921,N_2997);
nand UO_484 (O_484,N_2920,N_2911);
or UO_485 (O_485,N_2919,N_2968);
and UO_486 (O_486,N_2992,N_2966);
xor UO_487 (O_487,N_2972,N_2981);
nand UO_488 (O_488,N_2974,N_2930);
or UO_489 (O_489,N_2934,N_2940);
or UO_490 (O_490,N_2939,N_2906);
xnor UO_491 (O_491,N_2966,N_2923);
xor UO_492 (O_492,N_2919,N_2924);
nand UO_493 (O_493,N_2999,N_2963);
or UO_494 (O_494,N_2994,N_2962);
and UO_495 (O_495,N_2927,N_2956);
nor UO_496 (O_496,N_2963,N_2949);
xor UO_497 (O_497,N_2927,N_2945);
and UO_498 (O_498,N_2911,N_2902);
nor UO_499 (O_499,N_2951,N_2969);
endmodule