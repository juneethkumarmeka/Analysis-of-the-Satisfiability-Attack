module basic_1000_10000_1500_4_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
xor U0 (N_0,In_427,In_840);
or U1 (N_1,In_58,In_692);
nand U2 (N_2,In_272,In_144);
nand U3 (N_3,In_901,In_621);
or U4 (N_4,In_639,In_242);
xor U5 (N_5,In_228,In_369);
nor U6 (N_6,In_653,In_512);
or U7 (N_7,In_865,In_185);
nor U8 (N_8,In_588,In_345);
or U9 (N_9,In_173,In_633);
nor U10 (N_10,In_294,In_978);
xor U11 (N_11,In_608,In_233);
nor U12 (N_12,In_642,In_816);
and U13 (N_13,In_758,In_883);
nor U14 (N_14,In_81,In_352);
and U15 (N_15,In_542,In_763);
nor U16 (N_16,In_553,In_159);
nor U17 (N_17,In_806,In_734);
or U18 (N_18,In_85,In_699);
nor U19 (N_19,In_197,In_833);
nand U20 (N_20,In_18,In_537);
nor U21 (N_21,In_885,In_141);
xor U22 (N_22,In_899,In_567);
nor U23 (N_23,In_855,In_726);
or U24 (N_24,In_112,In_577);
nand U25 (N_25,In_264,In_86);
or U26 (N_26,In_7,In_679);
nor U27 (N_27,In_501,In_492);
or U28 (N_28,In_234,In_889);
nor U29 (N_29,In_519,In_593);
and U30 (N_30,In_171,In_839);
nor U31 (N_31,In_829,In_617);
or U32 (N_32,In_143,In_516);
nor U33 (N_33,In_504,In_64);
xor U34 (N_34,In_353,In_192);
nor U35 (N_35,In_483,In_971);
and U36 (N_36,In_456,In_569);
and U37 (N_37,In_227,In_999);
xnor U38 (N_38,In_939,In_761);
or U39 (N_39,In_582,In_206);
and U40 (N_40,In_757,In_290);
and U41 (N_41,In_321,In_663);
or U42 (N_42,In_163,In_802);
or U43 (N_43,In_405,In_302);
xnor U44 (N_44,In_273,In_98);
or U45 (N_45,In_138,In_993);
and U46 (N_46,In_475,In_662);
or U47 (N_47,In_732,In_74);
nand U48 (N_48,In_271,In_853);
nor U49 (N_49,In_245,In_380);
nor U50 (N_50,In_152,In_32);
nand U51 (N_51,In_884,In_913);
or U52 (N_52,In_818,In_694);
nor U53 (N_53,In_781,In_896);
nor U54 (N_54,In_47,In_991);
nand U55 (N_55,In_624,In_389);
and U56 (N_56,In_421,In_296);
or U57 (N_57,In_626,In_960);
and U58 (N_58,In_348,In_727);
nand U59 (N_59,In_876,In_390);
and U60 (N_60,In_386,In_246);
and U61 (N_61,In_35,In_480);
nand U62 (N_62,In_869,In_297);
xor U63 (N_63,In_441,In_4);
nor U64 (N_64,In_814,In_933);
nor U65 (N_65,In_465,In_160);
nor U66 (N_66,In_422,In_515);
xnor U67 (N_67,In_332,In_924);
or U68 (N_68,In_27,In_344);
and U69 (N_69,In_837,In_986);
or U70 (N_70,In_44,In_410);
xnor U71 (N_71,In_387,In_607);
xnor U72 (N_72,In_282,In_276);
or U73 (N_73,In_691,In_366);
nand U74 (N_74,In_555,In_716);
and U75 (N_75,In_964,In_956);
and U76 (N_76,In_605,In_499);
nand U77 (N_77,In_852,In_807);
nand U78 (N_78,In_832,In_48);
nand U79 (N_79,In_771,In_628);
nand U80 (N_80,In_908,In_927);
nor U81 (N_81,In_510,In_306);
nor U82 (N_82,In_14,In_643);
and U83 (N_83,In_697,In_307);
and U84 (N_84,In_376,In_768);
and U85 (N_85,In_792,In_647);
or U86 (N_86,In_961,In_725);
nand U87 (N_87,In_992,In_821);
and U88 (N_88,In_293,In_857);
or U89 (N_89,In_911,In_550);
or U90 (N_90,In_436,In_120);
nor U91 (N_91,In_110,In_904);
nand U92 (N_92,In_798,In_230);
nor U93 (N_93,In_938,In_985);
nand U94 (N_94,In_533,In_162);
and U95 (N_95,In_258,In_459);
nor U96 (N_96,In_72,In_998);
nor U97 (N_97,In_256,In_255);
or U98 (N_98,In_133,In_252);
nor U99 (N_99,In_146,In_278);
nand U100 (N_100,In_406,In_949);
and U101 (N_101,In_619,In_905);
nor U102 (N_102,In_817,In_616);
nand U103 (N_103,In_240,In_864);
or U104 (N_104,In_161,In_695);
and U105 (N_105,In_489,In_664);
nor U106 (N_106,In_75,In_164);
nor U107 (N_107,In_77,In_990);
nand U108 (N_108,In_898,In_473);
nand U109 (N_109,In_528,In_648);
or U110 (N_110,In_870,In_303);
and U111 (N_111,In_708,In_600);
and U112 (N_112,In_801,In_450);
or U113 (N_113,In_804,In_950);
nor U114 (N_114,In_474,In_45);
xnor U115 (N_115,In_432,In_326);
xor U116 (N_116,In_718,In_559);
or U117 (N_117,In_92,In_844);
and U118 (N_118,In_56,In_360);
and U119 (N_119,In_638,In_523);
and U120 (N_120,In_661,In_733);
nor U121 (N_121,In_765,In_862);
and U122 (N_122,In_683,In_836);
nand U123 (N_123,In_611,In_413);
nand U124 (N_124,In_87,In_738);
nor U125 (N_125,In_31,In_481);
xor U126 (N_126,In_851,In_590);
and U127 (N_127,In_931,In_828);
nand U128 (N_128,In_320,In_269);
or U129 (N_129,In_544,In_29);
or U130 (N_130,In_214,In_113);
or U131 (N_131,In_457,In_579);
or U132 (N_132,In_356,In_170);
nor U133 (N_133,In_742,In_793);
nand U134 (N_134,In_751,In_583);
nor U135 (N_135,In_637,In_116);
or U136 (N_136,In_522,In_540);
nand U137 (N_137,In_552,In_903);
nor U138 (N_138,In_127,In_415);
nor U139 (N_139,In_6,In_923);
nor U140 (N_140,In_872,In_224);
and U141 (N_141,In_351,In_10);
nor U142 (N_142,In_244,In_79);
nor U143 (N_143,In_155,In_169);
and U144 (N_144,In_641,In_919);
nand U145 (N_145,In_129,In_279);
nor U146 (N_146,In_397,In_330);
nor U147 (N_147,In_682,In_759);
or U148 (N_148,In_20,In_104);
and U149 (N_149,In_894,In_724);
or U150 (N_150,In_684,In_222);
nor U151 (N_151,In_313,In_40);
nand U152 (N_152,In_310,In_28);
nand U153 (N_153,In_575,In_36);
xor U154 (N_154,In_811,In_767);
and U155 (N_155,In_478,In_462);
nand U156 (N_156,In_399,In_741);
nor U157 (N_157,In_597,In_594);
and U158 (N_158,In_414,In_188);
xor U159 (N_159,In_791,In_176);
nor U160 (N_160,In_591,In_674);
nor U161 (N_161,In_139,In_437);
or U162 (N_162,In_654,In_805);
and U163 (N_163,In_825,In_630);
or U164 (N_164,In_953,In_447);
and U165 (N_165,In_912,In_518);
nor U166 (N_166,In_711,In_976);
or U167 (N_167,In_150,In_43);
nand U168 (N_168,In_744,In_917);
nor U169 (N_169,In_444,In_543);
nand U170 (N_170,In_167,In_565);
or U171 (N_171,In_225,In_687);
xor U172 (N_172,In_723,In_808);
nor U173 (N_173,In_729,In_983);
or U174 (N_174,In_880,In_122);
and U175 (N_175,In_442,In_706);
nand U176 (N_176,In_788,In_774);
nand U177 (N_177,In_586,In_49);
nand U178 (N_178,In_854,In_668);
or U179 (N_179,In_347,In_393);
or U180 (N_180,In_261,In_17);
nor U181 (N_181,In_612,In_34);
or U182 (N_182,In_941,In_823);
and U183 (N_183,In_204,In_66);
xnor U184 (N_184,In_215,In_90);
and U185 (N_185,In_117,In_810);
or U186 (N_186,In_997,In_267);
nand U187 (N_187,In_673,In_93);
and U188 (N_188,In_308,In_468);
and U189 (N_189,In_789,In_461);
and U190 (N_190,In_241,In_482);
or U191 (N_191,In_531,In_698);
nand U192 (N_192,In_766,In_400);
nand U193 (N_193,In_498,In_598);
or U194 (N_194,In_384,In_314);
xnor U195 (N_195,In_424,In_764);
nand U196 (N_196,In_819,In_3);
nor U197 (N_197,In_721,In_790);
nor U198 (N_198,In_70,In_707);
nand U199 (N_199,In_128,In_249);
nand U200 (N_200,In_355,In_604);
nor U201 (N_201,In_95,In_322);
xor U202 (N_202,In_454,In_878);
and U203 (N_203,In_100,In_275);
nor U204 (N_204,In_403,In_262);
nor U205 (N_205,In_728,In_189);
xnor U206 (N_206,In_336,In_538);
nor U207 (N_207,In_982,In_115);
or U208 (N_208,In_319,In_316);
nand U209 (N_209,In_809,In_902);
and U210 (N_210,In_218,In_378);
or U211 (N_211,In_486,In_300);
xnor U212 (N_212,In_21,In_370);
or U213 (N_213,In_97,In_105);
or U214 (N_214,In_312,In_860);
or U215 (N_215,In_346,In_560);
or U216 (N_216,In_84,In_41);
nor U217 (N_217,In_507,In_720);
nor U218 (N_218,In_895,In_815);
nand U219 (N_219,In_301,In_539);
nand U220 (N_220,In_268,In_676);
nand U221 (N_221,In_921,In_596);
nand U222 (N_222,In_419,In_700);
and U223 (N_223,In_752,In_988);
nor U224 (N_224,In_970,In_715);
and U225 (N_225,In_505,In_859);
or U226 (N_226,In_38,In_603);
or U227 (N_227,In_886,In_123);
nor U228 (N_228,In_257,In_137);
nand U229 (N_229,In_392,In_614);
and U230 (N_230,In_304,In_142);
xor U231 (N_231,In_566,In_179);
and U232 (N_232,In_796,In_194);
and U233 (N_233,In_73,In_750);
and U234 (N_234,In_1,In_417);
nor U235 (N_235,In_713,In_401);
nand U236 (N_236,In_357,In_263);
nor U237 (N_237,In_359,In_527);
and U238 (N_238,In_497,In_915);
and U239 (N_239,In_340,In_443);
nor U240 (N_240,In_205,In_782);
nand U241 (N_241,In_182,In_794);
and U242 (N_242,In_193,In_265);
and U243 (N_243,In_253,In_900);
nand U244 (N_244,In_223,In_13);
xnor U245 (N_245,In_584,In_660);
or U246 (N_246,In_944,In_918);
nor U247 (N_247,In_946,In_735);
and U248 (N_248,In_65,In_650);
and U249 (N_249,In_165,In_78);
and U250 (N_250,In_756,In_61);
nand U251 (N_251,In_503,In_856);
nor U252 (N_252,In_53,In_250);
or U253 (N_253,In_592,In_502);
nor U254 (N_254,In_63,In_777);
and U255 (N_255,In_776,In_89);
nor U256 (N_256,In_595,In_799);
nand U257 (N_257,In_820,In_848);
nand U258 (N_258,In_266,In_636);
nor U259 (N_259,In_281,In_822);
nor U260 (N_260,In_396,In_824);
nand U261 (N_261,In_495,In_198);
nand U262 (N_262,In_158,In_868);
nor U263 (N_263,In_574,In_963);
nor U264 (N_264,In_168,In_237);
nor U265 (N_265,In_76,In_930);
xnor U266 (N_266,In_358,In_132);
nand U267 (N_267,In_813,In_954);
or U268 (N_268,In_199,In_745);
nand U269 (N_269,In_845,In_299);
and U270 (N_270,In_463,In_644);
nor U271 (N_271,In_831,In_609);
nor U272 (N_272,In_342,In_94);
nand U273 (N_273,In_907,In_554);
xor U274 (N_274,In_364,In_585);
or U275 (N_275,In_610,In_381);
nand U276 (N_276,In_175,In_243);
or U277 (N_277,In_259,In_339);
or U278 (N_278,In_787,In_874);
and U279 (N_279,In_680,In_826);
and U280 (N_280,In_925,In_841);
or U281 (N_281,In_153,In_371);
and U282 (N_282,In_208,In_656);
xnor U283 (N_283,In_827,In_909);
xnor U284 (N_284,In_103,In_797);
nor U285 (N_285,In_375,In_157);
and U286 (N_286,In_529,In_893);
or U287 (N_287,In_471,In_305);
nand U288 (N_288,In_866,In_629);
and U289 (N_289,In_573,In_106);
and U290 (N_290,In_966,In_251);
and U291 (N_291,In_846,In_270);
nor U292 (N_292,In_62,In_379);
or U293 (N_293,In_172,In_689);
and U294 (N_294,In_755,In_317);
nor U295 (N_295,In_408,In_51);
and U296 (N_296,In_335,In_477);
or U297 (N_297,In_328,In_920);
and U298 (N_298,In_362,In_260);
nand U299 (N_299,In_108,In_433);
nor U300 (N_300,In_388,In_337);
xnor U301 (N_301,In_753,In_635);
or U302 (N_302,In_452,In_446);
and U303 (N_303,In_88,In_995);
nand U304 (N_304,In_140,In_196);
xor U305 (N_305,In_121,In_549);
or U306 (N_306,In_16,In_341);
nor U307 (N_307,In_526,In_570);
and U308 (N_308,In_331,In_277);
nor U309 (N_309,In_942,In_508);
nor U310 (N_310,In_119,In_54);
and U311 (N_311,In_5,In_690);
xor U312 (N_312,In_704,In_631);
or U313 (N_313,In_315,In_928);
or U314 (N_314,In_666,In_67);
and U315 (N_315,In_778,In_373);
xnor U316 (N_316,In_186,In_430);
or U317 (N_317,In_385,In_535);
nand U318 (N_318,In_145,In_25);
or U319 (N_319,In_82,In_323);
and U320 (N_320,In_365,In_216);
and U321 (N_321,In_760,In_625);
and U322 (N_322,In_311,In_835);
and U323 (N_323,In_407,In_219);
or U324 (N_324,In_968,In_298);
nand U325 (N_325,In_572,In_935);
and U326 (N_326,In_685,In_382);
nor U327 (N_327,In_779,In_398);
nand U328 (N_328,In_428,In_520);
nor U329 (N_329,In_717,In_236);
nand U330 (N_330,In_295,In_484);
nand U331 (N_331,In_910,In_99);
and U332 (N_332,In_453,In_368);
nor U333 (N_333,In_181,In_843);
and U334 (N_334,In_975,In_632);
nor U335 (N_335,In_479,In_563);
nor U336 (N_336,In_247,In_291);
or U337 (N_337,In_361,In_965);
and U338 (N_338,In_979,In_367);
or U339 (N_339,In_775,In_532);
nor U340 (N_340,In_50,In_800);
nand U341 (N_341,In_769,In_688);
and U342 (N_342,In_525,In_449);
and U343 (N_343,In_994,In_937);
nand U344 (N_344,In_602,In_850);
nor U345 (N_345,In_80,In_534);
or U346 (N_346,In_576,In_669);
nand U347 (N_347,In_488,In_945);
or U348 (N_348,In_803,In_890);
nand U349 (N_349,In_12,In_812);
nor U350 (N_350,In_551,In_363);
or U351 (N_351,In_101,In_22);
nand U352 (N_352,In_135,In_517);
nand U353 (N_353,In_784,In_786);
nand U354 (N_354,In_286,In_622);
xor U355 (N_355,In_743,In_232);
nor U356 (N_356,In_672,In_747);
and U357 (N_357,In_606,In_649);
nor U358 (N_358,In_701,In_309);
nor U359 (N_359,In_420,In_111);
nand U360 (N_360,In_37,In_102);
nor U361 (N_361,In_425,In_887);
nor U362 (N_362,In_615,In_235);
nand U363 (N_363,In_536,In_974);
or U364 (N_364,In_984,In_96);
or U365 (N_365,In_26,In_458);
nand U366 (N_366,In_429,In_125);
nor U367 (N_367,In_545,In_435);
nand U368 (N_368,In_418,In_785);
nor U369 (N_369,In_184,In_736);
nand U370 (N_370,In_220,In_338);
and U371 (N_371,In_740,In_254);
nor U372 (N_372,In_147,In_634);
and U373 (N_373,In_318,In_334);
or U374 (N_374,In_178,In_548);
or U375 (N_375,In_730,In_148);
nor U376 (N_376,In_847,In_423);
nor U377 (N_377,In_472,In_434);
nor U378 (N_378,In_292,In_705);
and U379 (N_379,In_731,In_118);
or U380 (N_380,In_659,In_213);
nand U381 (N_381,In_987,In_487);
or U382 (N_382,In_861,In_238);
or U383 (N_383,In_71,In_24);
or U384 (N_384,In_466,In_571);
nor U385 (N_385,In_558,In_922);
nand U386 (N_386,In_151,In_191);
nand U387 (N_387,In_748,In_412);
and U388 (N_388,In_969,In_329);
and U389 (N_389,In_858,In_248);
or U390 (N_390,In_947,In_934);
nand U391 (N_391,In_52,In_156);
nor U392 (N_392,In_324,In_211);
nand U393 (N_393,In_59,In_906);
xor U394 (N_394,In_957,In_842);
nor U395 (N_395,In_327,In_212);
nor U396 (N_396,In_209,In_469);
nand U397 (N_397,In_601,In_391);
xor U398 (N_398,In_546,In_183);
nor U399 (N_399,In_195,In_940);
nand U400 (N_400,In_349,In_411);
or U401 (N_401,In_404,In_667);
or U402 (N_402,In_556,In_174);
nor U403 (N_403,In_620,In_564);
nand U404 (N_404,In_521,In_287);
nor U405 (N_405,In_562,In_402);
nor U406 (N_406,In_943,In_675);
nand U407 (N_407,In_618,In_409);
nor U408 (N_408,In_383,In_149);
and U409 (N_409,In_696,In_274);
nand U410 (N_410,In_737,In_958);
nand U411 (N_411,In_166,In_581);
nor U412 (N_412,In_439,In_863);
nor U413 (N_413,In_60,In_873);
or U414 (N_414,In_686,In_15);
nand U415 (N_415,In_914,In_877);
nand U416 (N_416,In_980,In_107);
and U417 (N_417,In_514,In_681);
nor U418 (N_418,In_485,In_200);
and U419 (N_419,In_490,In_30);
or U420 (N_420,In_952,In_114);
nor U421 (N_421,In_702,In_530);
nand U422 (N_422,In_541,In_580);
nand U423 (N_423,In_445,In_283);
nor U424 (N_424,In_395,In_640);
nand U425 (N_425,In_221,In_892);
nor U426 (N_426,In_709,In_714);
nor U427 (N_427,In_8,In_426);
and U428 (N_428,In_494,In_416);
nor U429 (N_429,In_929,In_9);
and U430 (N_430,In_967,In_977);
and U431 (N_431,In_879,In_448);
nand U432 (N_432,In_126,In_867);
or U433 (N_433,In_394,In_746);
nor U434 (N_434,In_834,In_109);
nor U435 (N_435,In_849,In_627);
nor U436 (N_436,In_981,In_926);
or U437 (N_437,In_136,In_948);
nor U438 (N_438,In_451,In_202);
or U439 (N_439,In_68,In_578);
nor U440 (N_440,In_749,In_284);
xnor U441 (N_441,In_671,In_973);
nand U442 (N_442,In_374,In_280);
nor U443 (N_443,In_897,In_226);
and U444 (N_444,In_440,In_470);
and U445 (N_445,In_131,In_722);
or U446 (N_446,In_180,In_783);
nand U447 (N_447,In_210,In_773);
or U448 (N_448,In_464,In_561);
and U449 (N_449,In_506,In_936);
nand U450 (N_450,In_496,In_932);
nor U451 (N_451,In_589,In_438);
xor U452 (N_452,In_455,In_646);
nand U453 (N_453,In_325,In_69);
or U454 (N_454,In_55,In_288);
and U455 (N_455,In_652,In_693);
nand U456 (N_456,In_795,In_670);
and U457 (N_457,In_623,In_962);
nand U458 (N_458,In_770,In_124);
or U459 (N_459,In_710,In_996);
or U460 (N_460,In_217,In_951);
nor U461 (N_461,In_959,In_888);
and U462 (N_462,In_881,In_754);
or U463 (N_463,In_891,In_91);
xnor U464 (N_464,In_677,In_130);
nor U465 (N_465,In_289,In_231);
or U466 (N_466,In_739,In_229);
nor U467 (N_467,In_350,In_882);
nand U468 (N_468,In_207,In_989);
nor U469 (N_469,In_524,In_154);
and U470 (N_470,In_780,In_658);
nor U471 (N_471,In_500,In_871);
nand U472 (N_472,In_372,In_719);
nor U473 (N_473,In_875,In_343);
or U474 (N_474,In_645,In_916);
xor U475 (N_475,In_460,In_613);
nand U476 (N_476,In_46,In_703);
and U477 (N_477,In_11,In_19);
nor U478 (N_478,In_42,In_651);
nand U479 (N_479,In_678,In_187);
or U480 (N_480,In_830,In_587);
nand U481 (N_481,In_33,In_2);
or U482 (N_482,In_201,In_83);
and U483 (N_483,In_190,In_354);
nor U484 (N_484,In_655,In_177);
and U485 (N_485,In_431,In_333);
nor U486 (N_486,In_377,In_491);
nor U487 (N_487,In_493,In_547);
xor U488 (N_488,In_568,In_972);
nor U489 (N_489,In_513,In_557);
nor U490 (N_490,In_762,In_467);
xor U491 (N_491,In_23,In_39);
nor U492 (N_492,In_955,In_657);
nor U493 (N_493,In_203,In_599);
and U494 (N_494,In_838,In_476);
nand U495 (N_495,In_57,In_712);
and U496 (N_496,In_511,In_772);
nand U497 (N_497,In_665,In_509);
nor U498 (N_498,In_0,In_285);
and U499 (N_499,In_134,In_239);
nand U500 (N_500,In_651,In_25);
nor U501 (N_501,In_817,In_71);
nand U502 (N_502,In_522,In_148);
or U503 (N_503,In_602,In_384);
or U504 (N_504,In_422,In_753);
nor U505 (N_505,In_213,In_256);
and U506 (N_506,In_359,In_640);
or U507 (N_507,In_461,In_924);
xnor U508 (N_508,In_597,In_662);
nand U509 (N_509,In_447,In_258);
nor U510 (N_510,In_157,In_427);
and U511 (N_511,In_35,In_37);
xnor U512 (N_512,In_56,In_28);
nor U513 (N_513,In_442,In_475);
nor U514 (N_514,In_69,In_262);
or U515 (N_515,In_736,In_443);
and U516 (N_516,In_566,In_347);
nor U517 (N_517,In_931,In_269);
or U518 (N_518,In_669,In_158);
and U519 (N_519,In_481,In_690);
and U520 (N_520,In_642,In_972);
and U521 (N_521,In_650,In_732);
nor U522 (N_522,In_110,In_634);
or U523 (N_523,In_574,In_841);
nor U524 (N_524,In_180,In_635);
nand U525 (N_525,In_861,In_92);
nor U526 (N_526,In_48,In_809);
or U527 (N_527,In_341,In_69);
and U528 (N_528,In_668,In_856);
or U529 (N_529,In_262,In_310);
nand U530 (N_530,In_59,In_949);
and U531 (N_531,In_648,In_376);
and U532 (N_532,In_453,In_831);
or U533 (N_533,In_106,In_815);
nor U534 (N_534,In_559,In_66);
nand U535 (N_535,In_891,In_505);
and U536 (N_536,In_712,In_845);
xnor U537 (N_537,In_272,In_725);
or U538 (N_538,In_366,In_3);
and U539 (N_539,In_371,In_764);
nor U540 (N_540,In_172,In_850);
nor U541 (N_541,In_457,In_45);
and U542 (N_542,In_630,In_434);
xnor U543 (N_543,In_527,In_818);
nand U544 (N_544,In_183,In_912);
and U545 (N_545,In_336,In_855);
or U546 (N_546,In_15,In_886);
and U547 (N_547,In_870,In_104);
and U548 (N_548,In_191,In_954);
nand U549 (N_549,In_251,In_888);
or U550 (N_550,In_681,In_932);
nand U551 (N_551,In_962,In_96);
xnor U552 (N_552,In_756,In_979);
and U553 (N_553,In_522,In_866);
or U554 (N_554,In_310,In_129);
nor U555 (N_555,In_21,In_367);
nor U556 (N_556,In_320,In_237);
and U557 (N_557,In_685,In_307);
nor U558 (N_558,In_106,In_654);
nor U559 (N_559,In_950,In_679);
nand U560 (N_560,In_458,In_108);
nand U561 (N_561,In_433,In_186);
nand U562 (N_562,In_80,In_222);
nor U563 (N_563,In_910,In_757);
nand U564 (N_564,In_921,In_250);
nand U565 (N_565,In_312,In_185);
nor U566 (N_566,In_684,In_135);
and U567 (N_567,In_218,In_899);
and U568 (N_568,In_220,In_831);
or U569 (N_569,In_244,In_962);
or U570 (N_570,In_483,In_715);
and U571 (N_571,In_386,In_584);
or U572 (N_572,In_83,In_711);
nand U573 (N_573,In_699,In_453);
nand U574 (N_574,In_489,In_181);
nor U575 (N_575,In_298,In_437);
and U576 (N_576,In_422,In_788);
nor U577 (N_577,In_206,In_238);
nand U578 (N_578,In_230,In_214);
nand U579 (N_579,In_654,In_850);
nand U580 (N_580,In_781,In_526);
nand U581 (N_581,In_284,In_825);
or U582 (N_582,In_501,In_279);
nand U583 (N_583,In_829,In_400);
nand U584 (N_584,In_46,In_348);
nand U585 (N_585,In_165,In_144);
nand U586 (N_586,In_36,In_631);
nand U587 (N_587,In_263,In_184);
nand U588 (N_588,In_80,In_23);
or U589 (N_589,In_790,In_638);
or U590 (N_590,In_891,In_986);
nor U591 (N_591,In_503,In_262);
nand U592 (N_592,In_395,In_243);
nand U593 (N_593,In_712,In_926);
or U594 (N_594,In_635,In_52);
nand U595 (N_595,In_757,In_614);
xnor U596 (N_596,In_729,In_922);
nor U597 (N_597,In_979,In_4);
or U598 (N_598,In_403,In_799);
and U599 (N_599,In_685,In_560);
nor U600 (N_600,In_970,In_920);
or U601 (N_601,In_462,In_793);
nand U602 (N_602,In_886,In_491);
and U603 (N_603,In_57,In_831);
nand U604 (N_604,In_387,In_671);
or U605 (N_605,In_244,In_113);
and U606 (N_606,In_611,In_922);
xnor U607 (N_607,In_319,In_683);
or U608 (N_608,In_215,In_745);
nand U609 (N_609,In_825,In_89);
or U610 (N_610,In_364,In_826);
and U611 (N_611,In_801,In_964);
nand U612 (N_612,In_380,In_522);
or U613 (N_613,In_356,In_154);
nor U614 (N_614,In_514,In_574);
xor U615 (N_615,In_750,In_620);
nand U616 (N_616,In_671,In_720);
and U617 (N_617,In_747,In_728);
nor U618 (N_618,In_552,In_887);
or U619 (N_619,In_997,In_544);
nor U620 (N_620,In_834,In_89);
nor U621 (N_621,In_568,In_312);
and U622 (N_622,In_79,In_325);
or U623 (N_623,In_825,In_616);
or U624 (N_624,In_608,In_647);
and U625 (N_625,In_412,In_76);
nand U626 (N_626,In_516,In_824);
xnor U627 (N_627,In_584,In_764);
or U628 (N_628,In_721,In_484);
nand U629 (N_629,In_205,In_617);
nor U630 (N_630,In_225,In_544);
and U631 (N_631,In_833,In_291);
nand U632 (N_632,In_93,In_395);
nand U633 (N_633,In_624,In_247);
xnor U634 (N_634,In_511,In_199);
nor U635 (N_635,In_730,In_150);
nor U636 (N_636,In_515,In_686);
xor U637 (N_637,In_543,In_996);
nand U638 (N_638,In_603,In_570);
or U639 (N_639,In_530,In_692);
and U640 (N_640,In_809,In_270);
and U641 (N_641,In_790,In_297);
nand U642 (N_642,In_989,In_427);
nor U643 (N_643,In_769,In_886);
or U644 (N_644,In_425,In_817);
and U645 (N_645,In_528,In_184);
or U646 (N_646,In_460,In_738);
nand U647 (N_647,In_564,In_667);
or U648 (N_648,In_205,In_825);
or U649 (N_649,In_724,In_487);
or U650 (N_650,In_756,In_978);
or U651 (N_651,In_733,In_822);
xor U652 (N_652,In_893,In_577);
nor U653 (N_653,In_670,In_874);
nor U654 (N_654,In_718,In_284);
or U655 (N_655,In_46,In_716);
nor U656 (N_656,In_639,In_288);
and U657 (N_657,In_4,In_851);
nor U658 (N_658,In_280,In_491);
nor U659 (N_659,In_268,In_846);
nand U660 (N_660,In_925,In_739);
nor U661 (N_661,In_547,In_380);
nand U662 (N_662,In_107,In_967);
nand U663 (N_663,In_1,In_713);
or U664 (N_664,In_106,In_952);
xnor U665 (N_665,In_968,In_258);
and U666 (N_666,In_94,In_162);
nand U667 (N_667,In_269,In_668);
or U668 (N_668,In_866,In_180);
or U669 (N_669,In_855,In_590);
or U670 (N_670,In_145,In_607);
or U671 (N_671,In_97,In_74);
nor U672 (N_672,In_929,In_21);
or U673 (N_673,In_777,In_46);
nor U674 (N_674,In_679,In_921);
nor U675 (N_675,In_875,In_491);
nand U676 (N_676,In_140,In_536);
and U677 (N_677,In_87,In_704);
nor U678 (N_678,In_348,In_145);
and U679 (N_679,In_972,In_471);
or U680 (N_680,In_573,In_68);
nand U681 (N_681,In_352,In_331);
and U682 (N_682,In_399,In_894);
and U683 (N_683,In_759,In_514);
or U684 (N_684,In_673,In_897);
xnor U685 (N_685,In_400,In_969);
nor U686 (N_686,In_281,In_120);
and U687 (N_687,In_103,In_967);
nor U688 (N_688,In_61,In_483);
or U689 (N_689,In_569,In_331);
and U690 (N_690,In_6,In_761);
and U691 (N_691,In_995,In_594);
nand U692 (N_692,In_526,In_169);
nand U693 (N_693,In_630,In_301);
xnor U694 (N_694,In_462,In_770);
nor U695 (N_695,In_493,In_16);
or U696 (N_696,In_852,In_962);
and U697 (N_697,In_357,In_565);
nor U698 (N_698,In_197,In_56);
nor U699 (N_699,In_860,In_980);
and U700 (N_700,In_987,In_123);
nor U701 (N_701,In_286,In_191);
nor U702 (N_702,In_269,In_282);
and U703 (N_703,In_552,In_988);
xor U704 (N_704,In_493,In_451);
nor U705 (N_705,In_182,In_923);
nand U706 (N_706,In_738,In_381);
nand U707 (N_707,In_189,In_780);
nor U708 (N_708,In_915,In_650);
xor U709 (N_709,In_217,In_677);
nand U710 (N_710,In_785,In_631);
or U711 (N_711,In_885,In_351);
nand U712 (N_712,In_585,In_574);
nand U713 (N_713,In_728,In_554);
xor U714 (N_714,In_379,In_857);
nand U715 (N_715,In_584,In_885);
nor U716 (N_716,In_524,In_899);
nand U717 (N_717,In_623,In_460);
nand U718 (N_718,In_776,In_903);
nand U719 (N_719,In_97,In_977);
and U720 (N_720,In_95,In_450);
nand U721 (N_721,In_190,In_603);
or U722 (N_722,In_900,In_314);
xor U723 (N_723,In_445,In_227);
xor U724 (N_724,In_763,In_425);
and U725 (N_725,In_253,In_170);
nand U726 (N_726,In_232,In_802);
and U727 (N_727,In_263,In_215);
nand U728 (N_728,In_704,In_594);
xnor U729 (N_729,In_765,In_775);
or U730 (N_730,In_960,In_163);
and U731 (N_731,In_753,In_161);
and U732 (N_732,In_555,In_784);
or U733 (N_733,In_135,In_500);
nand U734 (N_734,In_740,In_931);
xnor U735 (N_735,In_234,In_411);
nand U736 (N_736,In_784,In_449);
or U737 (N_737,In_928,In_233);
and U738 (N_738,In_217,In_368);
and U739 (N_739,In_384,In_668);
or U740 (N_740,In_527,In_28);
nor U741 (N_741,In_403,In_867);
nand U742 (N_742,In_36,In_605);
and U743 (N_743,In_922,In_300);
and U744 (N_744,In_407,In_764);
or U745 (N_745,In_947,In_938);
nor U746 (N_746,In_110,In_470);
xnor U747 (N_747,In_529,In_194);
nand U748 (N_748,In_343,In_607);
and U749 (N_749,In_362,In_423);
and U750 (N_750,In_380,In_696);
or U751 (N_751,In_49,In_584);
nand U752 (N_752,In_221,In_219);
nand U753 (N_753,In_19,In_994);
nand U754 (N_754,In_270,In_701);
xnor U755 (N_755,In_780,In_662);
and U756 (N_756,In_263,In_141);
xor U757 (N_757,In_682,In_638);
and U758 (N_758,In_639,In_254);
nand U759 (N_759,In_383,In_909);
nand U760 (N_760,In_409,In_513);
and U761 (N_761,In_792,In_539);
nand U762 (N_762,In_22,In_619);
or U763 (N_763,In_719,In_484);
nand U764 (N_764,In_586,In_551);
nor U765 (N_765,In_650,In_529);
nand U766 (N_766,In_658,In_16);
xnor U767 (N_767,In_92,In_453);
nor U768 (N_768,In_439,In_206);
xnor U769 (N_769,In_963,In_629);
and U770 (N_770,In_357,In_127);
nor U771 (N_771,In_177,In_434);
nor U772 (N_772,In_396,In_376);
or U773 (N_773,In_121,In_67);
and U774 (N_774,In_927,In_400);
nor U775 (N_775,In_303,In_688);
and U776 (N_776,In_498,In_130);
and U777 (N_777,In_320,In_817);
nor U778 (N_778,In_350,In_512);
and U779 (N_779,In_863,In_698);
xnor U780 (N_780,In_918,In_832);
nor U781 (N_781,In_954,In_388);
or U782 (N_782,In_241,In_6);
nand U783 (N_783,In_884,In_848);
nor U784 (N_784,In_384,In_621);
nor U785 (N_785,In_25,In_906);
nor U786 (N_786,In_891,In_565);
nor U787 (N_787,In_403,In_976);
and U788 (N_788,In_451,In_4);
nand U789 (N_789,In_339,In_905);
or U790 (N_790,In_371,In_753);
or U791 (N_791,In_218,In_510);
and U792 (N_792,In_212,In_309);
or U793 (N_793,In_298,In_704);
or U794 (N_794,In_689,In_641);
or U795 (N_795,In_945,In_660);
nand U796 (N_796,In_444,In_715);
nand U797 (N_797,In_893,In_649);
or U798 (N_798,In_453,In_674);
or U799 (N_799,In_923,In_753);
or U800 (N_800,In_345,In_542);
nor U801 (N_801,In_54,In_730);
and U802 (N_802,In_570,In_188);
nor U803 (N_803,In_972,In_736);
and U804 (N_804,In_161,In_490);
nor U805 (N_805,In_956,In_23);
nor U806 (N_806,In_345,In_308);
nand U807 (N_807,In_387,In_597);
or U808 (N_808,In_567,In_771);
and U809 (N_809,In_260,In_290);
nor U810 (N_810,In_160,In_331);
and U811 (N_811,In_234,In_445);
nand U812 (N_812,In_762,In_549);
or U813 (N_813,In_572,In_643);
and U814 (N_814,In_185,In_733);
and U815 (N_815,In_889,In_372);
nor U816 (N_816,In_861,In_590);
and U817 (N_817,In_953,In_583);
nor U818 (N_818,In_962,In_542);
nand U819 (N_819,In_109,In_36);
nor U820 (N_820,In_200,In_339);
nor U821 (N_821,In_355,In_752);
and U822 (N_822,In_505,In_572);
nand U823 (N_823,In_558,In_878);
nor U824 (N_824,In_434,In_845);
or U825 (N_825,In_278,In_269);
xor U826 (N_826,In_273,In_874);
and U827 (N_827,In_664,In_702);
xor U828 (N_828,In_977,In_486);
and U829 (N_829,In_511,In_448);
nand U830 (N_830,In_600,In_442);
nand U831 (N_831,In_6,In_89);
nand U832 (N_832,In_4,In_768);
and U833 (N_833,In_477,In_864);
nand U834 (N_834,In_304,In_955);
xor U835 (N_835,In_376,In_221);
or U836 (N_836,In_176,In_932);
nand U837 (N_837,In_632,In_182);
nor U838 (N_838,In_383,In_67);
nand U839 (N_839,In_895,In_594);
xnor U840 (N_840,In_829,In_696);
and U841 (N_841,In_471,In_444);
nand U842 (N_842,In_611,In_444);
nand U843 (N_843,In_728,In_762);
and U844 (N_844,In_1,In_946);
or U845 (N_845,In_47,In_163);
or U846 (N_846,In_438,In_738);
nand U847 (N_847,In_122,In_200);
nand U848 (N_848,In_679,In_779);
nor U849 (N_849,In_473,In_46);
or U850 (N_850,In_223,In_175);
or U851 (N_851,In_936,In_691);
and U852 (N_852,In_724,In_148);
nand U853 (N_853,In_309,In_590);
nand U854 (N_854,In_788,In_188);
or U855 (N_855,In_178,In_256);
nor U856 (N_856,In_883,In_648);
nand U857 (N_857,In_338,In_395);
or U858 (N_858,In_464,In_64);
or U859 (N_859,In_922,In_120);
or U860 (N_860,In_296,In_377);
and U861 (N_861,In_946,In_179);
and U862 (N_862,In_442,In_955);
or U863 (N_863,In_363,In_509);
nand U864 (N_864,In_371,In_292);
and U865 (N_865,In_439,In_886);
nand U866 (N_866,In_883,In_756);
and U867 (N_867,In_561,In_839);
nor U868 (N_868,In_632,In_604);
or U869 (N_869,In_460,In_605);
or U870 (N_870,In_701,In_188);
nand U871 (N_871,In_316,In_649);
and U872 (N_872,In_737,In_751);
and U873 (N_873,In_423,In_725);
nor U874 (N_874,In_798,In_399);
and U875 (N_875,In_851,In_310);
nor U876 (N_876,In_254,In_421);
nand U877 (N_877,In_830,In_826);
or U878 (N_878,In_538,In_1);
nor U879 (N_879,In_262,In_792);
or U880 (N_880,In_407,In_722);
and U881 (N_881,In_164,In_385);
nand U882 (N_882,In_617,In_430);
nand U883 (N_883,In_768,In_74);
and U884 (N_884,In_334,In_229);
and U885 (N_885,In_755,In_82);
and U886 (N_886,In_146,In_625);
nor U887 (N_887,In_630,In_257);
nor U888 (N_888,In_317,In_221);
or U889 (N_889,In_60,In_293);
or U890 (N_890,In_824,In_856);
or U891 (N_891,In_279,In_732);
or U892 (N_892,In_418,In_85);
or U893 (N_893,In_403,In_569);
and U894 (N_894,In_790,In_606);
nand U895 (N_895,In_880,In_932);
and U896 (N_896,In_195,In_491);
nand U897 (N_897,In_649,In_306);
or U898 (N_898,In_781,In_335);
nor U899 (N_899,In_860,In_923);
or U900 (N_900,In_329,In_826);
nor U901 (N_901,In_782,In_196);
and U902 (N_902,In_333,In_539);
nor U903 (N_903,In_223,In_366);
and U904 (N_904,In_708,In_354);
and U905 (N_905,In_684,In_137);
and U906 (N_906,In_186,In_850);
or U907 (N_907,In_680,In_277);
nor U908 (N_908,In_100,In_791);
and U909 (N_909,In_767,In_943);
and U910 (N_910,In_418,In_374);
and U911 (N_911,In_299,In_242);
or U912 (N_912,In_546,In_395);
nor U913 (N_913,In_766,In_244);
xnor U914 (N_914,In_229,In_348);
or U915 (N_915,In_961,In_877);
nor U916 (N_916,In_226,In_271);
xnor U917 (N_917,In_695,In_878);
xnor U918 (N_918,In_180,In_232);
nor U919 (N_919,In_599,In_736);
xor U920 (N_920,In_780,In_50);
or U921 (N_921,In_831,In_173);
nand U922 (N_922,In_859,In_476);
and U923 (N_923,In_603,In_752);
nor U924 (N_924,In_547,In_482);
nor U925 (N_925,In_48,In_714);
and U926 (N_926,In_66,In_703);
xor U927 (N_927,In_508,In_619);
and U928 (N_928,In_75,In_527);
or U929 (N_929,In_946,In_809);
nand U930 (N_930,In_374,In_522);
nand U931 (N_931,In_82,In_623);
and U932 (N_932,In_264,In_322);
nor U933 (N_933,In_557,In_841);
nor U934 (N_934,In_428,In_377);
nand U935 (N_935,In_138,In_852);
and U936 (N_936,In_727,In_480);
or U937 (N_937,In_898,In_486);
nor U938 (N_938,In_536,In_279);
xnor U939 (N_939,In_196,In_929);
or U940 (N_940,In_544,In_259);
nor U941 (N_941,In_593,In_353);
and U942 (N_942,In_705,In_508);
and U943 (N_943,In_366,In_781);
nor U944 (N_944,In_932,In_368);
and U945 (N_945,In_536,In_390);
nor U946 (N_946,In_273,In_619);
or U947 (N_947,In_150,In_308);
or U948 (N_948,In_726,In_740);
nand U949 (N_949,In_601,In_936);
xnor U950 (N_950,In_435,In_593);
or U951 (N_951,In_546,In_181);
nor U952 (N_952,In_914,In_55);
and U953 (N_953,In_252,In_819);
nand U954 (N_954,In_821,In_123);
and U955 (N_955,In_411,In_625);
or U956 (N_956,In_271,In_710);
xnor U957 (N_957,In_892,In_467);
or U958 (N_958,In_806,In_349);
or U959 (N_959,In_890,In_922);
nor U960 (N_960,In_835,In_752);
and U961 (N_961,In_500,In_730);
xnor U962 (N_962,In_749,In_598);
or U963 (N_963,In_892,In_406);
or U964 (N_964,In_430,In_301);
nand U965 (N_965,In_180,In_776);
nand U966 (N_966,In_983,In_544);
or U967 (N_967,In_860,In_174);
nand U968 (N_968,In_529,In_450);
xnor U969 (N_969,In_954,In_268);
and U970 (N_970,In_650,In_874);
or U971 (N_971,In_447,In_409);
nor U972 (N_972,In_650,In_97);
nand U973 (N_973,In_856,In_430);
nand U974 (N_974,In_623,In_286);
nand U975 (N_975,In_582,In_572);
xor U976 (N_976,In_147,In_173);
nand U977 (N_977,In_638,In_227);
and U978 (N_978,In_489,In_889);
and U979 (N_979,In_605,In_975);
nor U980 (N_980,In_712,In_461);
nand U981 (N_981,In_52,In_757);
or U982 (N_982,In_518,In_969);
and U983 (N_983,In_491,In_805);
or U984 (N_984,In_501,In_380);
and U985 (N_985,In_19,In_867);
and U986 (N_986,In_907,In_781);
xnor U987 (N_987,In_474,In_541);
nor U988 (N_988,In_929,In_597);
or U989 (N_989,In_277,In_125);
xor U990 (N_990,In_692,In_290);
or U991 (N_991,In_600,In_720);
and U992 (N_992,In_835,In_181);
or U993 (N_993,In_847,In_97);
and U994 (N_994,In_643,In_158);
nand U995 (N_995,In_461,In_85);
and U996 (N_996,In_767,In_190);
or U997 (N_997,In_422,In_818);
nand U998 (N_998,In_560,In_797);
or U999 (N_999,In_142,In_662);
and U1000 (N_1000,In_874,In_724);
and U1001 (N_1001,In_525,In_764);
and U1002 (N_1002,In_891,In_381);
nor U1003 (N_1003,In_585,In_270);
xor U1004 (N_1004,In_47,In_450);
and U1005 (N_1005,In_724,In_903);
nand U1006 (N_1006,In_854,In_33);
xnor U1007 (N_1007,In_220,In_340);
or U1008 (N_1008,In_860,In_10);
nor U1009 (N_1009,In_48,In_249);
and U1010 (N_1010,In_325,In_749);
or U1011 (N_1011,In_253,In_914);
or U1012 (N_1012,In_984,In_246);
xnor U1013 (N_1013,In_941,In_359);
and U1014 (N_1014,In_684,In_444);
nor U1015 (N_1015,In_214,In_254);
xor U1016 (N_1016,In_70,In_937);
or U1017 (N_1017,In_817,In_63);
or U1018 (N_1018,In_465,In_459);
and U1019 (N_1019,In_981,In_99);
and U1020 (N_1020,In_835,In_567);
nor U1021 (N_1021,In_830,In_46);
xor U1022 (N_1022,In_476,In_364);
nor U1023 (N_1023,In_344,In_535);
nand U1024 (N_1024,In_838,In_154);
nor U1025 (N_1025,In_135,In_211);
and U1026 (N_1026,In_381,In_667);
nor U1027 (N_1027,In_187,In_426);
or U1028 (N_1028,In_254,In_781);
or U1029 (N_1029,In_949,In_576);
xnor U1030 (N_1030,In_163,In_422);
or U1031 (N_1031,In_748,In_925);
and U1032 (N_1032,In_72,In_692);
and U1033 (N_1033,In_309,In_24);
nand U1034 (N_1034,In_844,In_161);
and U1035 (N_1035,In_339,In_410);
and U1036 (N_1036,In_641,In_574);
nor U1037 (N_1037,In_35,In_399);
or U1038 (N_1038,In_256,In_300);
and U1039 (N_1039,In_157,In_244);
xnor U1040 (N_1040,In_843,In_846);
or U1041 (N_1041,In_83,In_759);
or U1042 (N_1042,In_205,In_973);
nor U1043 (N_1043,In_117,In_954);
or U1044 (N_1044,In_673,In_553);
and U1045 (N_1045,In_162,In_51);
or U1046 (N_1046,In_520,In_427);
nand U1047 (N_1047,In_112,In_878);
and U1048 (N_1048,In_945,In_584);
and U1049 (N_1049,In_9,In_387);
xnor U1050 (N_1050,In_632,In_696);
nand U1051 (N_1051,In_348,In_381);
or U1052 (N_1052,In_193,In_19);
and U1053 (N_1053,In_891,In_36);
or U1054 (N_1054,In_544,In_617);
or U1055 (N_1055,In_887,In_901);
nor U1056 (N_1056,In_556,In_955);
and U1057 (N_1057,In_775,In_1);
or U1058 (N_1058,In_639,In_358);
nand U1059 (N_1059,In_737,In_656);
nand U1060 (N_1060,In_30,In_929);
or U1061 (N_1061,In_764,In_832);
and U1062 (N_1062,In_483,In_984);
nand U1063 (N_1063,In_185,In_295);
or U1064 (N_1064,In_314,In_543);
xnor U1065 (N_1065,In_877,In_884);
nand U1066 (N_1066,In_342,In_172);
nor U1067 (N_1067,In_310,In_645);
nand U1068 (N_1068,In_531,In_231);
nor U1069 (N_1069,In_376,In_607);
nand U1070 (N_1070,In_316,In_970);
nor U1071 (N_1071,In_559,In_862);
and U1072 (N_1072,In_686,In_239);
nor U1073 (N_1073,In_609,In_528);
xor U1074 (N_1074,In_660,In_533);
or U1075 (N_1075,In_114,In_390);
nor U1076 (N_1076,In_327,In_760);
or U1077 (N_1077,In_827,In_512);
or U1078 (N_1078,In_585,In_847);
and U1079 (N_1079,In_883,In_712);
and U1080 (N_1080,In_885,In_132);
nor U1081 (N_1081,In_182,In_995);
and U1082 (N_1082,In_37,In_3);
and U1083 (N_1083,In_405,In_86);
and U1084 (N_1084,In_998,In_847);
and U1085 (N_1085,In_395,In_267);
nand U1086 (N_1086,In_968,In_937);
xor U1087 (N_1087,In_977,In_41);
nor U1088 (N_1088,In_727,In_240);
and U1089 (N_1089,In_815,In_853);
nand U1090 (N_1090,In_105,In_293);
and U1091 (N_1091,In_998,In_127);
nand U1092 (N_1092,In_338,In_714);
nor U1093 (N_1093,In_831,In_270);
nand U1094 (N_1094,In_673,In_316);
nand U1095 (N_1095,In_765,In_80);
or U1096 (N_1096,In_113,In_683);
xor U1097 (N_1097,In_545,In_976);
and U1098 (N_1098,In_336,In_34);
and U1099 (N_1099,In_853,In_107);
nor U1100 (N_1100,In_872,In_622);
nor U1101 (N_1101,In_411,In_33);
nor U1102 (N_1102,In_545,In_568);
and U1103 (N_1103,In_699,In_336);
and U1104 (N_1104,In_250,In_124);
or U1105 (N_1105,In_791,In_887);
nand U1106 (N_1106,In_353,In_340);
and U1107 (N_1107,In_183,In_675);
xnor U1108 (N_1108,In_608,In_197);
or U1109 (N_1109,In_690,In_439);
nand U1110 (N_1110,In_714,In_535);
xor U1111 (N_1111,In_76,In_968);
or U1112 (N_1112,In_446,In_409);
nor U1113 (N_1113,In_297,In_24);
nand U1114 (N_1114,In_511,In_657);
nand U1115 (N_1115,In_558,In_160);
nand U1116 (N_1116,In_975,In_196);
and U1117 (N_1117,In_220,In_684);
nand U1118 (N_1118,In_5,In_517);
nand U1119 (N_1119,In_129,In_741);
nand U1120 (N_1120,In_805,In_619);
nand U1121 (N_1121,In_850,In_324);
xor U1122 (N_1122,In_145,In_840);
nor U1123 (N_1123,In_375,In_747);
xor U1124 (N_1124,In_152,In_861);
and U1125 (N_1125,In_168,In_950);
or U1126 (N_1126,In_709,In_905);
and U1127 (N_1127,In_769,In_82);
nor U1128 (N_1128,In_831,In_73);
nor U1129 (N_1129,In_949,In_412);
nand U1130 (N_1130,In_115,In_738);
nand U1131 (N_1131,In_892,In_10);
xor U1132 (N_1132,In_878,In_955);
xor U1133 (N_1133,In_671,In_517);
nor U1134 (N_1134,In_311,In_587);
nor U1135 (N_1135,In_546,In_6);
nand U1136 (N_1136,In_524,In_512);
or U1137 (N_1137,In_240,In_497);
nor U1138 (N_1138,In_882,In_917);
or U1139 (N_1139,In_640,In_316);
nand U1140 (N_1140,In_368,In_854);
nand U1141 (N_1141,In_121,In_29);
or U1142 (N_1142,In_696,In_289);
nor U1143 (N_1143,In_28,In_562);
or U1144 (N_1144,In_862,In_130);
or U1145 (N_1145,In_904,In_832);
nand U1146 (N_1146,In_674,In_575);
or U1147 (N_1147,In_495,In_696);
or U1148 (N_1148,In_598,In_771);
nor U1149 (N_1149,In_792,In_205);
nand U1150 (N_1150,In_958,In_767);
or U1151 (N_1151,In_221,In_460);
nor U1152 (N_1152,In_62,In_567);
nor U1153 (N_1153,In_987,In_295);
nand U1154 (N_1154,In_561,In_283);
nor U1155 (N_1155,In_558,In_886);
nor U1156 (N_1156,In_790,In_467);
and U1157 (N_1157,In_531,In_404);
nor U1158 (N_1158,In_931,In_860);
nor U1159 (N_1159,In_234,In_633);
and U1160 (N_1160,In_186,In_21);
nor U1161 (N_1161,In_869,In_782);
and U1162 (N_1162,In_87,In_987);
nor U1163 (N_1163,In_252,In_791);
and U1164 (N_1164,In_82,In_348);
xor U1165 (N_1165,In_683,In_280);
nor U1166 (N_1166,In_295,In_7);
or U1167 (N_1167,In_711,In_404);
or U1168 (N_1168,In_303,In_57);
and U1169 (N_1169,In_301,In_348);
nor U1170 (N_1170,In_633,In_554);
and U1171 (N_1171,In_780,In_57);
nand U1172 (N_1172,In_547,In_133);
nor U1173 (N_1173,In_823,In_958);
and U1174 (N_1174,In_138,In_914);
or U1175 (N_1175,In_379,In_116);
and U1176 (N_1176,In_216,In_330);
or U1177 (N_1177,In_486,In_512);
nor U1178 (N_1178,In_920,In_533);
and U1179 (N_1179,In_869,In_22);
and U1180 (N_1180,In_171,In_408);
nand U1181 (N_1181,In_915,In_154);
xnor U1182 (N_1182,In_376,In_405);
xnor U1183 (N_1183,In_310,In_97);
nand U1184 (N_1184,In_320,In_553);
and U1185 (N_1185,In_607,In_998);
or U1186 (N_1186,In_439,In_461);
or U1187 (N_1187,In_516,In_26);
or U1188 (N_1188,In_176,In_72);
nor U1189 (N_1189,In_947,In_281);
and U1190 (N_1190,In_914,In_64);
or U1191 (N_1191,In_679,In_170);
or U1192 (N_1192,In_31,In_693);
and U1193 (N_1193,In_925,In_326);
or U1194 (N_1194,In_547,In_89);
nor U1195 (N_1195,In_348,In_711);
or U1196 (N_1196,In_963,In_54);
and U1197 (N_1197,In_169,In_976);
or U1198 (N_1198,In_874,In_236);
and U1199 (N_1199,In_123,In_789);
or U1200 (N_1200,In_115,In_908);
or U1201 (N_1201,In_903,In_425);
xnor U1202 (N_1202,In_697,In_505);
xnor U1203 (N_1203,In_531,In_220);
nor U1204 (N_1204,In_504,In_517);
nor U1205 (N_1205,In_573,In_319);
nor U1206 (N_1206,In_452,In_174);
and U1207 (N_1207,In_792,In_630);
nand U1208 (N_1208,In_462,In_61);
nand U1209 (N_1209,In_513,In_717);
and U1210 (N_1210,In_305,In_545);
and U1211 (N_1211,In_715,In_890);
and U1212 (N_1212,In_215,In_329);
xnor U1213 (N_1213,In_211,In_271);
or U1214 (N_1214,In_463,In_710);
and U1215 (N_1215,In_171,In_528);
and U1216 (N_1216,In_495,In_77);
nand U1217 (N_1217,In_400,In_481);
nand U1218 (N_1218,In_93,In_553);
nor U1219 (N_1219,In_85,In_977);
or U1220 (N_1220,In_804,In_877);
and U1221 (N_1221,In_637,In_168);
or U1222 (N_1222,In_471,In_887);
and U1223 (N_1223,In_519,In_864);
or U1224 (N_1224,In_124,In_89);
and U1225 (N_1225,In_909,In_727);
nor U1226 (N_1226,In_990,In_987);
nor U1227 (N_1227,In_476,In_817);
and U1228 (N_1228,In_198,In_118);
or U1229 (N_1229,In_605,In_739);
and U1230 (N_1230,In_2,In_367);
and U1231 (N_1231,In_424,In_841);
and U1232 (N_1232,In_63,In_945);
and U1233 (N_1233,In_570,In_990);
nor U1234 (N_1234,In_872,In_466);
nor U1235 (N_1235,In_48,In_937);
nand U1236 (N_1236,In_686,In_614);
nor U1237 (N_1237,In_176,In_215);
and U1238 (N_1238,In_737,In_908);
nor U1239 (N_1239,In_660,In_502);
or U1240 (N_1240,In_703,In_933);
nor U1241 (N_1241,In_422,In_282);
and U1242 (N_1242,In_607,In_135);
or U1243 (N_1243,In_44,In_51);
nand U1244 (N_1244,In_753,In_466);
and U1245 (N_1245,In_442,In_277);
nor U1246 (N_1246,In_215,In_437);
nand U1247 (N_1247,In_980,In_0);
and U1248 (N_1248,In_986,In_508);
nor U1249 (N_1249,In_961,In_200);
and U1250 (N_1250,In_386,In_902);
or U1251 (N_1251,In_718,In_452);
nor U1252 (N_1252,In_662,In_775);
and U1253 (N_1253,In_392,In_225);
nor U1254 (N_1254,In_663,In_678);
xor U1255 (N_1255,In_463,In_818);
or U1256 (N_1256,In_594,In_13);
or U1257 (N_1257,In_483,In_100);
nor U1258 (N_1258,In_748,In_446);
nor U1259 (N_1259,In_568,In_180);
or U1260 (N_1260,In_973,In_722);
xor U1261 (N_1261,In_571,In_498);
or U1262 (N_1262,In_441,In_296);
nor U1263 (N_1263,In_161,In_771);
and U1264 (N_1264,In_127,In_805);
and U1265 (N_1265,In_986,In_899);
or U1266 (N_1266,In_858,In_741);
nand U1267 (N_1267,In_402,In_544);
and U1268 (N_1268,In_615,In_849);
or U1269 (N_1269,In_694,In_634);
or U1270 (N_1270,In_292,In_551);
or U1271 (N_1271,In_170,In_940);
nor U1272 (N_1272,In_386,In_72);
nand U1273 (N_1273,In_587,In_239);
and U1274 (N_1274,In_526,In_537);
nor U1275 (N_1275,In_445,In_12);
xnor U1276 (N_1276,In_576,In_259);
or U1277 (N_1277,In_697,In_331);
xnor U1278 (N_1278,In_289,In_21);
nor U1279 (N_1279,In_720,In_616);
nor U1280 (N_1280,In_229,In_369);
nand U1281 (N_1281,In_556,In_378);
nand U1282 (N_1282,In_281,In_663);
or U1283 (N_1283,In_25,In_467);
and U1284 (N_1284,In_969,In_565);
nor U1285 (N_1285,In_843,In_679);
or U1286 (N_1286,In_227,In_236);
nor U1287 (N_1287,In_660,In_102);
nand U1288 (N_1288,In_587,In_640);
or U1289 (N_1289,In_399,In_728);
nor U1290 (N_1290,In_51,In_669);
and U1291 (N_1291,In_787,In_502);
or U1292 (N_1292,In_377,In_138);
nor U1293 (N_1293,In_455,In_556);
nor U1294 (N_1294,In_559,In_535);
nand U1295 (N_1295,In_151,In_240);
xor U1296 (N_1296,In_322,In_525);
or U1297 (N_1297,In_362,In_600);
xor U1298 (N_1298,In_782,In_60);
nor U1299 (N_1299,In_978,In_739);
or U1300 (N_1300,In_678,In_271);
nor U1301 (N_1301,In_473,In_408);
and U1302 (N_1302,In_149,In_742);
nor U1303 (N_1303,In_902,In_399);
or U1304 (N_1304,In_112,In_806);
nand U1305 (N_1305,In_240,In_724);
or U1306 (N_1306,In_475,In_708);
or U1307 (N_1307,In_127,In_119);
and U1308 (N_1308,In_855,In_270);
nor U1309 (N_1309,In_268,In_856);
or U1310 (N_1310,In_233,In_277);
nand U1311 (N_1311,In_328,In_691);
xor U1312 (N_1312,In_28,In_725);
xor U1313 (N_1313,In_329,In_205);
or U1314 (N_1314,In_550,In_800);
nand U1315 (N_1315,In_218,In_976);
and U1316 (N_1316,In_516,In_578);
nor U1317 (N_1317,In_496,In_443);
or U1318 (N_1318,In_844,In_746);
and U1319 (N_1319,In_309,In_80);
and U1320 (N_1320,In_685,In_924);
nor U1321 (N_1321,In_167,In_806);
and U1322 (N_1322,In_249,In_522);
nand U1323 (N_1323,In_762,In_45);
and U1324 (N_1324,In_246,In_299);
nand U1325 (N_1325,In_533,In_644);
nor U1326 (N_1326,In_278,In_893);
and U1327 (N_1327,In_420,In_2);
xnor U1328 (N_1328,In_737,In_701);
nor U1329 (N_1329,In_855,In_768);
nand U1330 (N_1330,In_936,In_703);
nor U1331 (N_1331,In_495,In_15);
nand U1332 (N_1332,In_146,In_327);
nand U1333 (N_1333,In_189,In_657);
xor U1334 (N_1334,In_685,In_398);
nand U1335 (N_1335,In_475,In_52);
nand U1336 (N_1336,In_559,In_164);
xor U1337 (N_1337,In_427,In_632);
nand U1338 (N_1338,In_850,In_167);
and U1339 (N_1339,In_434,In_481);
nand U1340 (N_1340,In_869,In_390);
nor U1341 (N_1341,In_904,In_537);
nor U1342 (N_1342,In_727,In_904);
xnor U1343 (N_1343,In_649,In_506);
nand U1344 (N_1344,In_289,In_852);
nor U1345 (N_1345,In_709,In_669);
nor U1346 (N_1346,In_921,In_370);
xnor U1347 (N_1347,In_298,In_784);
and U1348 (N_1348,In_972,In_233);
or U1349 (N_1349,In_446,In_238);
or U1350 (N_1350,In_862,In_998);
nor U1351 (N_1351,In_302,In_477);
or U1352 (N_1352,In_10,In_20);
nor U1353 (N_1353,In_717,In_901);
or U1354 (N_1354,In_619,In_587);
nand U1355 (N_1355,In_70,In_340);
nand U1356 (N_1356,In_762,In_547);
nand U1357 (N_1357,In_406,In_953);
nor U1358 (N_1358,In_333,In_252);
or U1359 (N_1359,In_702,In_461);
nor U1360 (N_1360,In_246,In_451);
nor U1361 (N_1361,In_769,In_956);
xnor U1362 (N_1362,In_868,In_306);
nand U1363 (N_1363,In_899,In_665);
nor U1364 (N_1364,In_695,In_62);
nand U1365 (N_1365,In_687,In_879);
xor U1366 (N_1366,In_369,In_384);
and U1367 (N_1367,In_96,In_625);
nor U1368 (N_1368,In_95,In_766);
xor U1369 (N_1369,In_439,In_849);
or U1370 (N_1370,In_240,In_986);
nand U1371 (N_1371,In_818,In_786);
or U1372 (N_1372,In_85,In_539);
nand U1373 (N_1373,In_600,In_775);
or U1374 (N_1374,In_439,In_360);
nand U1375 (N_1375,In_113,In_795);
or U1376 (N_1376,In_584,In_703);
nor U1377 (N_1377,In_299,In_418);
nand U1378 (N_1378,In_910,In_893);
nand U1379 (N_1379,In_253,In_85);
nand U1380 (N_1380,In_566,In_928);
or U1381 (N_1381,In_317,In_942);
nand U1382 (N_1382,In_168,In_4);
nor U1383 (N_1383,In_700,In_164);
and U1384 (N_1384,In_303,In_825);
and U1385 (N_1385,In_296,In_171);
nor U1386 (N_1386,In_727,In_580);
or U1387 (N_1387,In_124,In_440);
or U1388 (N_1388,In_875,In_994);
or U1389 (N_1389,In_720,In_946);
or U1390 (N_1390,In_377,In_234);
nor U1391 (N_1391,In_704,In_358);
nor U1392 (N_1392,In_909,In_959);
and U1393 (N_1393,In_970,In_947);
nand U1394 (N_1394,In_807,In_979);
or U1395 (N_1395,In_996,In_504);
nand U1396 (N_1396,In_116,In_186);
nor U1397 (N_1397,In_305,In_380);
nand U1398 (N_1398,In_525,In_795);
or U1399 (N_1399,In_783,In_758);
or U1400 (N_1400,In_443,In_799);
nand U1401 (N_1401,In_711,In_294);
nor U1402 (N_1402,In_741,In_337);
or U1403 (N_1403,In_355,In_328);
and U1404 (N_1404,In_993,In_938);
xor U1405 (N_1405,In_102,In_300);
or U1406 (N_1406,In_532,In_479);
and U1407 (N_1407,In_873,In_142);
or U1408 (N_1408,In_995,In_928);
nand U1409 (N_1409,In_816,In_233);
or U1410 (N_1410,In_626,In_16);
and U1411 (N_1411,In_863,In_844);
and U1412 (N_1412,In_578,In_658);
nor U1413 (N_1413,In_201,In_30);
nor U1414 (N_1414,In_940,In_555);
nor U1415 (N_1415,In_483,In_124);
nor U1416 (N_1416,In_779,In_160);
and U1417 (N_1417,In_833,In_283);
nor U1418 (N_1418,In_215,In_403);
and U1419 (N_1419,In_213,In_982);
and U1420 (N_1420,In_663,In_215);
nand U1421 (N_1421,In_778,In_116);
and U1422 (N_1422,In_951,In_418);
nor U1423 (N_1423,In_836,In_776);
and U1424 (N_1424,In_644,In_879);
or U1425 (N_1425,In_215,In_414);
or U1426 (N_1426,In_282,In_853);
xnor U1427 (N_1427,In_65,In_659);
nand U1428 (N_1428,In_419,In_479);
and U1429 (N_1429,In_324,In_446);
or U1430 (N_1430,In_707,In_580);
nand U1431 (N_1431,In_494,In_714);
nand U1432 (N_1432,In_355,In_466);
xnor U1433 (N_1433,In_210,In_514);
and U1434 (N_1434,In_508,In_361);
xnor U1435 (N_1435,In_783,In_147);
nor U1436 (N_1436,In_864,In_717);
or U1437 (N_1437,In_448,In_443);
nor U1438 (N_1438,In_254,In_343);
xnor U1439 (N_1439,In_461,In_233);
nand U1440 (N_1440,In_947,In_329);
nor U1441 (N_1441,In_193,In_739);
xor U1442 (N_1442,In_769,In_995);
and U1443 (N_1443,In_44,In_225);
or U1444 (N_1444,In_926,In_380);
and U1445 (N_1445,In_826,In_495);
nor U1446 (N_1446,In_443,In_908);
or U1447 (N_1447,In_428,In_635);
nor U1448 (N_1448,In_195,In_631);
and U1449 (N_1449,In_559,In_78);
nor U1450 (N_1450,In_390,In_848);
and U1451 (N_1451,In_207,In_77);
nor U1452 (N_1452,In_522,In_645);
nand U1453 (N_1453,In_433,In_764);
nor U1454 (N_1454,In_412,In_525);
or U1455 (N_1455,In_214,In_738);
or U1456 (N_1456,In_515,In_750);
and U1457 (N_1457,In_783,In_381);
or U1458 (N_1458,In_55,In_407);
or U1459 (N_1459,In_661,In_299);
nor U1460 (N_1460,In_384,In_345);
nand U1461 (N_1461,In_81,In_487);
and U1462 (N_1462,In_863,In_724);
nor U1463 (N_1463,In_11,In_398);
and U1464 (N_1464,In_31,In_30);
nand U1465 (N_1465,In_227,In_216);
and U1466 (N_1466,In_369,In_550);
or U1467 (N_1467,In_335,In_600);
or U1468 (N_1468,In_270,In_65);
nor U1469 (N_1469,In_648,In_414);
or U1470 (N_1470,In_481,In_732);
or U1471 (N_1471,In_919,In_9);
nand U1472 (N_1472,In_564,In_749);
or U1473 (N_1473,In_874,In_117);
nand U1474 (N_1474,In_693,In_467);
nor U1475 (N_1475,In_913,In_75);
and U1476 (N_1476,In_403,In_136);
nor U1477 (N_1477,In_215,In_590);
nand U1478 (N_1478,In_813,In_572);
and U1479 (N_1479,In_974,In_751);
and U1480 (N_1480,In_614,In_809);
or U1481 (N_1481,In_596,In_639);
or U1482 (N_1482,In_872,In_201);
xnor U1483 (N_1483,In_176,In_408);
nor U1484 (N_1484,In_107,In_240);
and U1485 (N_1485,In_389,In_736);
and U1486 (N_1486,In_361,In_335);
nor U1487 (N_1487,In_123,In_639);
or U1488 (N_1488,In_607,In_367);
nand U1489 (N_1489,In_970,In_338);
and U1490 (N_1490,In_982,In_822);
nand U1491 (N_1491,In_731,In_824);
xnor U1492 (N_1492,In_663,In_942);
nand U1493 (N_1493,In_575,In_56);
nor U1494 (N_1494,In_674,In_547);
xnor U1495 (N_1495,In_384,In_674);
nor U1496 (N_1496,In_987,In_29);
or U1497 (N_1497,In_169,In_233);
nand U1498 (N_1498,In_28,In_933);
and U1499 (N_1499,In_417,In_67);
and U1500 (N_1500,In_659,In_751);
or U1501 (N_1501,In_149,In_587);
and U1502 (N_1502,In_203,In_104);
and U1503 (N_1503,In_310,In_969);
nand U1504 (N_1504,In_319,In_729);
and U1505 (N_1505,In_933,In_186);
xor U1506 (N_1506,In_420,In_936);
xnor U1507 (N_1507,In_300,In_296);
nand U1508 (N_1508,In_514,In_533);
nor U1509 (N_1509,In_800,In_391);
nor U1510 (N_1510,In_951,In_98);
or U1511 (N_1511,In_170,In_276);
xor U1512 (N_1512,In_98,In_917);
xor U1513 (N_1513,In_534,In_535);
nand U1514 (N_1514,In_317,In_560);
xor U1515 (N_1515,In_879,In_90);
nand U1516 (N_1516,In_71,In_637);
nand U1517 (N_1517,In_635,In_382);
nand U1518 (N_1518,In_581,In_476);
and U1519 (N_1519,In_812,In_197);
or U1520 (N_1520,In_118,In_688);
nand U1521 (N_1521,In_744,In_202);
and U1522 (N_1522,In_830,In_733);
or U1523 (N_1523,In_784,In_753);
or U1524 (N_1524,In_312,In_18);
xor U1525 (N_1525,In_908,In_493);
or U1526 (N_1526,In_9,In_546);
and U1527 (N_1527,In_288,In_689);
nor U1528 (N_1528,In_69,In_443);
nor U1529 (N_1529,In_283,In_97);
nand U1530 (N_1530,In_850,In_262);
nand U1531 (N_1531,In_858,In_814);
nor U1532 (N_1532,In_81,In_103);
and U1533 (N_1533,In_714,In_843);
and U1534 (N_1534,In_41,In_263);
or U1535 (N_1535,In_619,In_633);
and U1536 (N_1536,In_742,In_48);
nor U1537 (N_1537,In_291,In_955);
nand U1538 (N_1538,In_592,In_6);
nand U1539 (N_1539,In_20,In_913);
and U1540 (N_1540,In_106,In_986);
nor U1541 (N_1541,In_380,In_572);
or U1542 (N_1542,In_171,In_606);
and U1543 (N_1543,In_967,In_399);
or U1544 (N_1544,In_227,In_994);
and U1545 (N_1545,In_492,In_433);
nor U1546 (N_1546,In_696,In_66);
and U1547 (N_1547,In_546,In_768);
and U1548 (N_1548,In_529,In_159);
or U1549 (N_1549,In_631,In_262);
and U1550 (N_1550,In_739,In_534);
or U1551 (N_1551,In_867,In_578);
nor U1552 (N_1552,In_162,In_538);
nor U1553 (N_1553,In_84,In_40);
and U1554 (N_1554,In_548,In_438);
nor U1555 (N_1555,In_575,In_855);
and U1556 (N_1556,In_75,In_565);
nand U1557 (N_1557,In_143,In_469);
nand U1558 (N_1558,In_634,In_898);
nor U1559 (N_1559,In_908,In_792);
nor U1560 (N_1560,In_254,In_667);
nor U1561 (N_1561,In_892,In_331);
nand U1562 (N_1562,In_7,In_308);
and U1563 (N_1563,In_912,In_346);
nor U1564 (N_1564,In_790,In_637);
nand U1565 (N_1565,In_681,In_86);
and U1566 (N_1566,In_51,In_510);
nand U1567 (N_1567,In_614,In_138);
and U1568 (N_1568,In_321,In_83);
or U1569 (N_1569,In_413,In_96);
and U1570 (N_1570,In_940,In_212);
or U1571 (N_1571,In_763,In_930);
and U1572 (N_1572,In_408,In_447);
xnor U1573 (N_1573,In_257,In_869);
nor U1574 (N_1574,In_581,In_913);
or U1575 (N_1575,In_203,In_844);
nor U1576 (N_1576,In_756,In_477);
nor U1577 (N_1577,In_242,In_491);
nor U1578 (N_1578,In_229,In_476);
xnor U1579 (N_1579,In_615,In_12);
and U1580 (N_1580,In_745,In_708);
or U1581 (N_1581,In_123,In_42);
or U1582 (N_1582,In_795,In_489);
nand U1583 (N_1583,In_315,In_464);
xor U1584 (N_1584,In_530,In_205);
or U1585 (N_1585,In_490,In_812);
nor U1586 (N_1586,In_597,In_255);
or U1587 (N_1587,In_441,In_913);
or U1588 (N_1588,In_26,In_604);
nand U1589 (N_1589,In_692,In_718);
and U1590 (N_1590,In_891,In_808);
nor U1591 (N_1591,In_848,In_157);
xor U1592 (N_1592,In_758,In_699);
nand U1593 (N_1593,In_319,In_119);
nand U1594 (N_1594,In_417,In_712);
xnor U1595 (N_1595,In_477,In_911);
nand U1596 (N_1596,In_813,In_716);
nand U1597 (N_1597,In_732,In_137);
nand U1598 (N_1598,In_579,In_801);
nand U1599 (N_1599,In_388,In_600);
nand U1600 (N_1600,In_414,In_105);
xor U1601 (N_1601,In_967,In_445);
and U1602 (N_1602,In_28,In_307);
and U1603 (N_1603,In_753,In_513);
or U1604 (N_1604,In_320,In_655);
nand U1605 (N_1605,In_183,In_311);
or U1606 (N_1606,In_911,In_518);
nand U1607 (N_1607,In_577,In_262);
nor U1608 (N_1608,In_123,In_780);
nand U1609 (N_1609,In_375,In_581);
nand U1610 (N_1610,In_844,In_655);
and U1611 (N_1611,In_952,In_563);
nor U1612 (N_1612,In_60,In_893);
nor U1613 (N_1613,In_391,In_979);
or U1614 (N_1614,In_820,In_667);
nand U1615 (N_1615,In_178,In_301);
nand U1616 (N_1616,In_216,In_927);
nor U1617 (N_1617,In_12,In_141);
nor U1618 (N_1618,In_334,In_827);
or U1619 (N_1619,In_563,In_118);
or U1620 (N_1620,In_880,In_750);
nor U1621 (N_1621,In_265,In_596);
xnor U1622 (N_1622,In_883,In_406);
or U1623 (N_1623,In_713,In_274);
xnor U1624 (N_1624,In_935,In_156);
nor U1625 (N_1625,In_723,In_623);
nand U1626 (N_1626,In_455,In_325);
nand U1627 (N_1627,In_174,In_850);
or U1628 (N_1628,In_407,In_768);
nand U1629 (N_1629,In_577,In_911);
and U1630 (N_1630,In_518,In_238);
nand U1631 (N_1631,In_795,In_832);
xor U1632 (N_1632,In_632,In_808);
and U1633 (N_1633,In_756,In_177);
or U1634 (N_1634,In_594,In_298);
and U1635 (N_1635,In_665,In_939);
nor U1636 (N_1636,In_150,In_620);
nor U1637 (N_1637,In_449,In_808);
and U1638 (N_1638,In_582,In_916);
or U1639 (N_1639,In_767,In_186);
and U1640 (N_1640,In_237,In_620);
nand U1641 (N_1641,In_978,In_586);
nand U1642 (N_1642,In_469,In_265);
nor U1643 (N_1643,In_959,In_502);
nand U1644 (N_1644,In_216,In_437);
and U1645 (N_1645,In_872,In_820);
and U1646 (N_1646,In_726,In_446);
nor U1647 (N_1647,In_359,In_675);
or U1648 (N_1648,In_727,In_535);
xnor U1649 (N_1649,In_565,In_551);
nand U1650 (N_1650,In_571,In_755);
and U1651 (N_1651,In_112,In_762);
and U1652 (N_1652,In_399,In_521);
or U1653 (N_1653,In_287,In_959);
or U1654 (N_1654,In_545,In_596);
nor U1655 (N_1655,In_603,In_794);
nand U1656 (N_1656,In_724,In_451);
or U1657 (N_1657,In_815,In_182);
or U1658 (N_1658,In_263,In_219);
nand U1659 (N_1659,In_827,In_176);
nand U1660 (N_1660,In_318,In_216);
and U1661 (N_1661,In_313,In_18);
or U1662 (N_1662,In_71,In_171);
xnor U1663 (N_1663,In_435,In_350);
nor U1664 (N_1664,In_750,In_513);
nor U1665 (N_1665,In_489,In_962);
xor U1666 (N_1666,In_720,In_615);
xor U1667 (N_1667,In_573,In_871);
xnor U1668 (N_1668,In_234,In_351);
or U1669 (N_1669,In_215,In_464);
and U1670 (N_1670,In_648,In_893);
nor U1671 (N_1671,In_694,In_922);
xnor U1672 (N_1672,In_768,In_221);
nand U1673 (N_1673,In_553,In_494);
or U1674 (N_1674,In_80,In_440);
xnor U1675 (N_1675,In_982,In_170);
or U1676 (N_1676,In_40,In_162);
nand U1677 (N_1677,In_377,In_449);
or U1678 (N_1678,In_3,In_988);
nand U1679 (N_1679,In_686,In_85);
xnor U1680 (N_1680,In_509,In_689);
nor U1681 (N_1681,In_27,In_415);
xor U1682 (N_1682,In_597,In_480);
nor U1683 (N_1683,In_467,In_785);
or U1684 (N_1684,In_127,In_221);
nand U1685 (N_1685,In_30,In_709);
nand U1686 (N_1686,In_799,In_327);
or U1687 (N_1687,In_905,In_920);
xnor U1688 (N_1688,In_996,In_806);
or U1689 (N_1689,In_389,In_489);
nand U1690 (N_1690,In_315,In_140);
nand U1691 (N_1691,In_955,In_454);
nand U1692 (N_1692,In_332,In_975);
and U1693 (N_1693,In_516,In_388);
nand U1694 (N_1694,In_163,In_322);
nand U1695 (N_1695,In_486,In_106);
xnor U1696 (N_1696,In_90,In_592);
nor U1697 (N_1697,In_927,In_31);
nand U1698 (N_1698,In_747,In_374);
nand U1699 (N_1699,In_948,In_628);
nor U1700 (N_1700,In_504,In_803);
or U1701 (N_1701,In_973,In_958);
and U1702 (N_1702,In_658,In_535);
or U1703 (N_1703,In_51,In_728);
or U1704 (N_1704,In_636,In_232);
or U1705 (N_1705,In_290,In_610);
or U1706 (N_1706,In_424,In_713);
and U1707 (N_1707,In_28,In_184);
xnor U1708 (N_1708,In_850,In_742);
nor U1709 (N_1709,In_306,In_495);
or U1710 (N_1710,In_578,In_44);
and U1711 (N_1711,In_922,In_203);
nand U1712 (N_1712,In_472,In_110);
and U1713 (N_1713,In_33,In_305);
nand U1714 (N_1714,In_487,In_200);
nand U1715 (N_1715,In_408,In_975);
and U1716 (N_1716,In_389,In_921);
or U1717 (N_1717,In_8,In_784);
xnor U1718 (N_1718,In_489,In_867);
or U1719 (N_1719,In_185,In_904);
and U1720 (N_1720,In_745,In_827);
or U1721 (N_1721,In_234,In_805);
nor U1722 (N_1722,In_953,In_420);
nor U1723 (N_1723,In_352,In_68);
or U1724 (N_1724,In_862,In_632);
nand U1725 (N_1725,In_976,In_409);
and U1726 (N_1726,In_485,In_724);
or U1727 (N_1727,In_607,In_890);
and U1728 (N_1728,In_293,In_661);
or U1729 (N_1729,In_964,In_59);
or U1730 (N_1730,In_985,In_380);
nor U1731 (N_1731,In_378,In_611);
xor U1732 (N_1732,In_644,In_630);
nor U1733 (N_1733,In_448,In_74);
or U1734 (N_1734,In_464,In_390);
or U1735 (N_1735,In_559,In_655);
or U1736 (N_1736,In_57,In_76);
or U1737 (N_1737,In_715,In_922);
nand U1738 (N_1738,In_444,In_368);
and U1739 (N_1739,In_749,In_559);
nor U1740 (N_1740,In_381,In_270);
nor U1741 (N_1741,In_545,In_426);
and U1742 (N_1742,In_92,In_519);
or U1743 (N_1743,In_197,In_294);
and U1744 (N_1744,In_367,In_40);
or U1745 (N_1745,In_185,In_397);
or U1746 (N_1746,In_4,In_135);
nor U1747 (N_1747,In_905,In_47);
nand U1748 (N_1748,In_411,In_884);
nand U1749 (N_1749,In_433,In_680);
and U1750 (N_1750,In_616,In_591);
nor U1751 (N_1751,In_707,In_605);
nand U1752 (N_1752,In_715,In_779);
nor U1753 (N_1753,In_200,In_25);
nor U1754 (N_1754,In_558,In_94);
and U1755 (N_1755,In_495,In_231);
or U1756 (N_1756,In_358,In_44);
nand U1757 (N_1757,In_822,In_248);
nand U1758 (N_1758,In_23,In_316);
or U1759 (N_1759,In_570,In_770);
or U1760 (N_1760,In_378,In_405);
nand U1761 (N_1761,In_61,In_424);
nor U1762 (N_1762,In_477,In_504);
and U1763 (N_1763,In_576,In_625);
nand U1764 (N_1764,In_18,In_652);
or U1765 (N_1765,In_232,In_7);
or U1766 (N_1766,In_559,In_301);
and U1767 (N_1767,In_379,In_483);
nor U1768 (N_1768,In_373,In_33);
and U1769 (N_1769,In_796,In_517);
xnor U1770 (N_1770,In_927,In_619);
or U1771 (N_1771,In_137,In_884);
and U1772 (N_1772,In_863,In_946);
xor U1773 (N_1773,In_229,In_864);
nor U1774 (N_1774,In_909,In_966);
xnor U1775 (N_1775,In_335,In_947);
nand U1776 (N_1776,In_8,In_519);
or U1777 (N_1777,In_352,In_931);
and U1778 (N_1778,In_589,In_974);
nand U1779 (N_1779,In_413,In_565);
nand U1780 (N_1780,In_34,In_460);
or U1781 (N_1781,In_64,In_153);
or U1782 (N_1782,In_614,In_79);
and U1783 (N_1783,In_282,In_288);
nor U1784 (N_1784,In_238,In_311);
nand U1785 (N_1785,In_851,In_615);
and U1786 (N_1786,In_450,In_855);
nand U1787 (N_1787,In_151,In_682);
nor U1788 (N_1788,In_677,In_848);
or U1789 (N_1789,In_214,In_351);
nor U1790 (N_1790,In_596,In_801);
or U1791 (N_1791,In_696,In_840);
nor U1792 (N_1792,In_364,In_707);
and U1793 (N_1793,In_531,In_829);
nor U1794 (N_1794,In_276,In_399);
nor U1795 (N_1795,In_276,In_701);
nor U1796 (N_1796,In_55,In_392);
and U1797 (N_1797,In_727,In_714);
and U1798 (N_1798,In_241,In_9);
or U1799 (N_1799,In_159,In_844);
or U1800 (N_1800,In_619,In_955);
or U1801 (N_1801,In_645,In_193);
nor U1802 (N_1802,In_970,In_181);
and U1803 (N_1803,In_201,In_153);
and U1804 (N_1804,In_975,In_443);
nand U1805 (N_1805,In_180,In_104);
and U1806 (N_1806,In_514,In_264);
xor U1807 (N_1807,In_857,In_536);
or U1808 (N_1808,In_152,In_105);
and U1809 (N_1809,In_270,In_768);
and U1810 (N_1810,In_99,In_192);
or U1811 (N_1811,In_104,In_310);
and U1812 (N_1812,In_440,In_586);
or U1813 (N_1813,In_250,In_634);
nor U1814 (N_1814,In_849,In_245);
xor U1815 (N_1815,In_904,In_839);
xor U1816 (N_1816,In_860,In_278);
nand U1817 (N_1817,In_450,In_850);
and U1818 (N_1818,In_394,In_928);
xor U1819 (N_1819,In_281,In_113);
xor U1820 (N_1820,In_434,In_541);
and U1821 (N_1821,In_714,In_9);
and U1822 (N_1822,In_731,In_977);
and U1823 (N_1823,In_41,In_383);
or U1824 (N_1824,In_588,In_286);
or U1825 (N_1825,In_916,In_842);
or U1826 (N_1826,In_683,In_815);
nor U1827 (N_1827,In_491,In_728);
or U1828 (N_1828,In_748,In_203);
and U1829 (N_1829,In_211,In_907);
nand U1830 (N_1830,In_114,In_597);
nor U1831 (N_1831,In_909,In_166);
nor U1832 (N_1832,In_207,In_93);
and U1833 (N_1833,In_697,In_322);
nand U1834 (N_1834,In_269,In_332);
or U1835 (N_1835,In_839,In_303);
nand U1836 (N_1836,In_138,In_125);
or U1837 (N_1837,In_655,In_52);
nand U1838 (N_1838,In_519,In_100);
or U1839 (N_1839,In_422,In_736);
nand U1840 (N_1840,In_501,In_365);
nand U1841 (N_1841,In_989,In_981);
xor U1842 (N_1842,In_269,In_899);
or U1843 (N_1843,In_832,In_323);
and U1844 (N_1844,In_930,In_332);
nand U1845 (N_1845,In_356,In_264);
and U1846 (N_1846,In_182,In_888);
nor U1847 (N_1847,In_794,In_534);
or U1848 (N_1848,In_378,In_903);
and U1849 (N_1849,In_93,In_715);
and U1850 (N_1850,In_384,In_14);
nor U1851 (N_1851,In_20,In_667);
and U1852 (N_1852,In_47,In_66);
nand U1853 (N_1853,In_282,In_909);
and U1854 (N_1854,In_387,In_101);
nor U1855 (N_1855,In_137,In_805);
nor U1856 (N_1856,In_931,In_713);
xnor U1857 (N_1857,In_554,In_680);
and U1858 (N_1858,In_652,In_730);
nor U1859 (N_1859,In_245,In_972);
xor U1860 (N_1860,In_17,In_268);
and U1861 (N_1861,In_490,In_557);
or U1862 (N_1862,In_584,In_531);
and U1863 (N_1863,In_296,In_156);
nand U1864 (N_1864,In_366,In_809);
nor U1865 (N_1865,In_350,In_469);
and U1866 (N_1866,In_671,In_113);
nand U1867 (N_1867,In_625,In_515);
nor U1868 (N_1868,In_192,In_956);
nand U1869 (N_1869,In_271,In_932);
nor U1870 (N_1870,In_44,In_206);
xor U1871 (N_1871,In_831,In_827);
nand U1872 (N_1872,In_366,In_113);
nor U1873 (N_1873,In_834,In_508);
nand U1874 (N_1874,In_738,In_163);
nand U1875 (N_1875,In_465,In_329);
and U1876 (N_1876,In_418,In_559);
xnor U1877 (N_1877,In_884,In_286);
or U1878 (N_1878,In_337,In_135);
nand U1879 (N_1879,In_723,In_98);
xor U1880 (N_1880,In_29,In_131);
nor U1881 (N_1881,In_683,In_375);
and U1882 (N_1882,In_787,In_340);
nand U1883 (N_1883,In_745,In_468);
or U1884 (N_1884,In_243,In_296);
nor U1885 (N_1885,In_717,In_134);
or U1886 (N_1886,In_15,In_548);
or U1887 (N_1887,In_572,In_130);
nand U1888 (N_1888,In_956,In_710);
nand U1889 (N_1889,In_961,In_834);
or U1890 (N_1890,In_609,In_432);
xor U1891 (N_1891,In_267,In_71);
nand U1892 (N_1892,In_38,In_247);
nand U1893 (N_1893,In_694,In_333);
nand U1894 (N_1894,In_7,In_570);
nand U1895 (N_1895,In_475,In_918);
and U1896 (N_1896,In_531,In_711);
nand U1897 (N_1897,In_987,In_519);
and U1898 (N_1898,In_266,In_12);
or U1899 (N_1899,In_872,In_326);
nor U1900 (N_1900,In_224,In_169);
or U1901 (N_1901,In_693,In_598);
or U1902 (N_1902,In_422,In_376);
nor U1903 (N_1903,In_961,In_438);
or U1904 (N_1904,In_603,In_809);
nor U1905 (N_1905,In_377,In_481);
nand U1906 (N_1906,In_766,In_430);
or U1907 (N_1907,In_549,In_833);
xnor U1908 (N_1908,In_401,In_985);
xor U1909 (N_1909,In_166,In_634);
nand U1910 (N_1910,In_150,In_74);
nand U1911 (N_1911,In_906,In_561);
nor U1912 (N_1912,In_663,In_648);
and U1913 (N_1913,In_447,In_200);
nand U1914 (N_1914,In_383,In_559);
or U1915 (N_1915,In_848,In_56);
nor U1916 (N_1916,In_268,In_331);
xor U1917 (N_1917,In_353,In_580);
nor U1918 (N_1918,In_974,In_81);
and U1919 (N_1919,In_223,In_426);
and U1920 (N_1920,In_466,In_248);
nor U1921 (N_1921,In_924,In_485);
or U1922 (N_1922,In_976,In_707);
nand U1923 (N_1923,In_193,In_310);
or U1924 (N_1924,In_169,In_164);
and U1925 (N_1925,In_17,In_789);
nor U1926 (N_1926,In_215,In_479);
and U1927 (N_1927,In_14,In_5);
nand U1928 (N_1928,In_59,In_87);
nand U1929 (N_1929,In_968,In_49);
nand U1930 (N_1930,In_311,In_749);
or U1931 (N_1931,In_405,In_520);
and U1932 (N_1932,In_37,In_316);
or U1933 (N_1933,In_358,In_278);
nand U1934 (N_1934,In_922,In_369);
or U1935 (N_1935,In_372,In_706);
or U1936 (N_1936,In_929,In_255);
xor U1937 (N_1937,In_691,In_663);
nand U1938 (N_1938,In_207,In_108);
and U1939 (N_1939,In_231,In_765);
or U1940 (N_1940,In_281,In_338);
or U1941 (N_1941,In_39,In_294);
nor U1942 (N_1942,In_154,In_133);
and U1943 (N_1943,In_675,In_947);
or U1944 (N_1944,In_515,In_521);
xnor U1945 (N_1945,In_599,In_692);
nand U1946 (N_1946,In_445,In_830);
nand U1947 (N_1947,In_166,In_127);
nor U1948 (N_1948,In_659,In_396);
xor U1949 (N_1949,In_171,In_869);
nand U1950 (N_1950,In_466,In_798);
or U1951 (N_1951,In_538,In_771);
or U1952 (N_1952,In_30,In_435);
nor U1953 (N_1953,In_815,In_484);
or U1954 (N_1954,In_358,In_866);
or U1955 (N_1955,In_825,In_86);
and U1956 (N_1956,In_825,In_652);
or U1957 (N_1957,In_209,In_518);
nor U1958 (N_1958,In_610,In_136);
nor U1959 (N_1959,In_390,In_260);
or U1960 (N_1960,In_801,In_686);
and U1961 (N_1961,In_150,In_159);
nand U1962 (N_1962,In_925,In_863);
nand U1963 (N_1963,In_634,In_408);
or U1964 (N_1964,In_104,In_421);
or U1965 (N_1965,In_798,In_750);
and U1966 (N_1966,In_305,In_399);
and U1967 (N_1967,In_675,In_700);
and U1968 (N_1968,In_412,In_400);
nor U1969 (N_1969,In_194,In_749);
nor U1970 (N_1970,In_716,In_80);
nor U1971 (N_1971,In_765,In_104);
nor U1972 (N_1972,In_866,In_468);
and U1973 (N_1973,In_702,In_989);
xnor U1974 (N_1974,In_675,In_545);
xor U1975 (N_1975,In_869,In_446);
nand U1976 (N_1976,In_525,In_254);
and U1977 (N_1977,In_44,In_726);
nand U1978 (N_1978,In_201,In_290);
nor U1979 (N_1979,In_530,In_519);
nand U1980 (N_1980,In_432,In_747);
or U1981 (N_1981,In_586,In_675);
or U1982 (N_1982,In_303,In_349);
nor U1983 (N_1983,In_877,In_678);
or U1984 (N_1984,In_640,In_525);
nor U1985 (N_1985,In_117,In_362);
xor U1986 (N_1986,In_680,In_854);
nor U1987 (N_1987,In_868,In_281);
nor U1988 (N_1988,In_798,In_541);
nor U1989 (N_1989,In_945,In_740);
nor U1990 (N_1990,In_839,In_342);
nand U1991 (N_1991,In_507,In_298);
nor U1992 (N_1992,In_363,In_731);
xor U1993 (N_1993,In_515,In_80);
nor U1994 (N_1994,In_503,In_796);
and U1995 (N_1995,In_549,In_4);
nor U1996 (N_1996,In_740,In_882);
nor U1997 (N_1997,In_741,In_41);
nand U1998 (N_1998,In_87,In_450);
or U1999 (N_1999,In_537,In_244);
and U2000 (N_2000,In_121,In_915);
nand U2001 (N_2001,In_237,In_365);
nor U2002 (N_2002,In_957,In_660);
nand U2003 (N_2003,In_397,In_540);
or U2004 (N_2004,In_273,In_174);
or U2005 (N_2005,In_795,In_345);
or U2006 (N_2006,In_424,In_135);
nand U2007 (N_2007,In_940,In_326);
or U2008 (N_2008,In_803,In_482);
nor U2009 (N_2009,In_877,In_114);
nor U2010 (N_2010,In_995,In_386);
nand U2011 (N_2011,In_110,In_466);
nor U2012 (N_2012,In_370,In_358);
or U2013 (N_2013,In_620,In_690);
xnor U2014 (N_2014,In_298,In_196);
and U2015 (N_2015,In_999,In_708);
nor U2016 (N_2016,In_204,In_584);
and U2017 (N_2017,In_738,In_523);
nor U2018 (N_2018,In_879,In_552);
or U2019 (N_2019,In_412,In_703);
or U2020 (N_2020,In_294,In_369);
and U2021 (N_2021,In_259,In_289);
nand U2022 (N_2022,In_804,In_549);
and U2023 (N_2023,In_336,In_545);
and U2024 (N_2024,In_905,In_362);
nand U2025 (N_2025,In_20,In_369);
or U2026 (N_2026,In_119,In_314);
or U2027 (N_2027,In_76,In_715);
xor U2028 (N_2028,In_346,In_91);
and U2029 (N_2029,In_137,In_871);
nor U2030 (N_2030,In_111,In_957);
and U2031 (N_2031,In_529,In_842);
or U2032 (N_2032,In_917,In_423);
nor U2033 (N_2033,In_794,In_545);
nor U2034 (N_2034,In_633,In_822);
and U2035 (N_2035,In_200,In_616);
or U2036 (N_2036,In_842,In_634);
or U2037 (N_2037,In_577,In_374);
and U2038 (N_2038,In_264,In_787);
nor U2039 (N_2039,In_830,In_492);
nand U2040 (N_2040,In_891,In_371);
or U2041 (N_2041,In_882,In_572);
xor U2042 (N_2042,In_659,In_23);
nand U2043 (N_2043,In_445,In_41);
and U2044 (N_2044,In_793,In_622);
xnor U2045 (N_2045,In_500,In_973);
or U2046 (N_2046,In_706,In_798);
nand U2047 (N_2047,In_836,In_96);
nor U2048 (N_2048,In_672,In_216);
nand U2049 (N_2049,In_714,In_259);
and U2050 (N_2050,In_806,In_993);
and U2051 (N_2051,In_737,In_943);
and U2052 (N_2052,In_7,In_911);
or U2053 (N_2053,In_190,In_769);
and U2054 (N_2054,In_845,In_460);
or U2055 (N_2055,In_689,In_159);
nor U2056 (N_2056,In_625,In_151);
nor U2057 (N_2057,In_69,In_871);
nor U2058 (N_2058,In_592,In_812);
and U2059 (N_2059,In_235,In_1);
nor U2060 (N_2060,In_227,In_720);
nand U2061 (N_2061,In_738,In_989);
nand U2062 (N_2062,In_392,In_880);
or U2063 (N_2063,In_649,In_869);
nand U2064 (N_2064,In_796,In_30);
nor U2065 (N_2065,In_641,In_984);
nand U2066 (N_2066,In_603,In_465);
or U2067 (N_2067,In_182,In_742);
and U2068 (N_2068,In_638,In_461);
xnor U2069 (N_2069,In_502,In_379);
nand U2070 (N_2070,In_928,In_869);
and U2071 (N_2071,In_928,In_271);
and U2072 (N_2072,In_959,In_580);
nor U2073 (N_2073,In_474,In_774);
xnor U2074 (N_2074,In_175,In_757);
nand U2075 (N_2075,In_126,In_754);
nand U2076 (N_2076,In_668,In_867);
xnor U2077 (N_2077,In_340,In_487);
or U2078 (N_2078,In_101,In_628);
and U2079 (N_2079,In_966,In_475);
and U2080 (N_2080,In_250,In_595);
nor U2081 (N_2081,In_242,In_87);
xnor U2082 (N_2082,In_532,In_437);
or U2083 (N_2083,In_822,In_440);
nor U2084 (N_2084,In_611,In_696);
nand U2085 (N_2085,In_147,In_212);
and U2086 (N_2086,In_239,In_423);
xor U2087 (N_2087,In_842,In_34);
and U2088 (N_2088,In_23,In_356);
and U2089 (N_2089,In_530,In_473);
nor U2090 (N_2090,In_674,In_912);
or U2091 (N_2091,In_424,In_917);
nor U2092 (N_2092,In_798,In_205);
or U2093 (N_2093,In_692,In_560);
xor U2094 (N_2094,In_151,In_586);
nor U2095 (N_2095,In_558,In_835);
nor U2096 (N_2096,In_806,In_987);
nor U2097 (N_2097,In_711,In_953);
nor U2098 (N_2098,In_848,In_854);
nand U2099 (N_2099,In_104,In_603);
nor U2100 (N_2100,In_343,In_372);
or U2101 (N_2101,In_473,In_317);
nand U2102 (N_2102,In_196,In_244);
nor U2103 (N_2103,In_15,In_480);
or U2104 (N_2104,In_122,In_260);
nor U2105 (N_2105,In_619,In_634);
nand U2106 (N_2106,In_106,In_467);
nor U2107 (N_2107,In_544,In_690);
nand U2108 (N_2108,In_815,In_173);
or U2109 (N_2109,In_137,In_968);
or U2110 (N_2110,In_15,In_481);
xor U2111 (N_2111,In_712,In_328);
xnor U2112 (N_2112,In_60,In_148);
nor U2113 (N_2113,In_103,In_362);
nor U2114 (N_2114,In_928,In_178);
or U2115 (N_2115,In_938,In_560);
nand U2116 (N_2116,In_428,In_19);
or U2117 (N_2117,In_655,In_995);
and U2118 (N_2118,In_393,In_959);
nor U2119 (N_2119,In_9,In_521);
nor U2120 (N_2120,In_835,In_787);
or U2121 (N_2121,In_787,In_890);
or U2122 (N_2122,In_191,In_542);
xor U2123 (N_2123,In_509,In_982);
or U2124 (N_2124,In_201,In_887);
nor U2125 (N_2125,In_20,In_534);
and U2126 (N_2126,In_434,In_944);
nand U2127 (N_2127,In_372,In_941);
or U2128 (N_2128,In_323,In_450);
or U2129 (N_2129,In_72,In_770);
and U2130 (N_2130,In_883,In_95);
nand U2131 (N_2131,In_851,In_667);
nand U2132 (N_2132,In_66,In_23);
nor U2133 (N_2133,In_680,In_804);
and U2134 (N_2134,In_308,In_518);
nor U2135 (N_2135,In_607,In_522);
nor U2136 (N_2136,In_413,In_629);
or U2137 (N_2137,In_428,In_420);
nor U2138 (N_2138,In_372,In_53);
and U2139 (N_2139,In_218,In_892);
and U2140 (N_2140,In_962,In_275);
or U2141 (N_2141,In_550,In_728);
or U2142 (N_2142,In_897,In_737);
or U2143 (N_2143,In_18,In_298);
nand U2144 (N_2144,In_974,In_929);
and U2145 (N_2145,In_629,In_783);
nand U2146 (N_2146,In_638,In_520);
nor U2147 (N_2147,In_84,In_640);
nor U2148 (N_2148,In_47,In_607);
nor U2149 (N_2149,In_486,In_874);
nand U2150 (N_2150,In_41,In_797);
or U2151 (N_2151,In_32,In_553);
and U2152 (N_2152,In_89,In_799);
and U2153 (N_2153,In_584,In_346);
and U2154 (N_2154,In_842,In_719);
nand U2155 (N_2155,In_171,In_947);
or U2156 (N_2156,In_182,In_214);
nand U2157 (N_2157,In_176,In_375);
and U2158 (N_2158,In_575,In_453);
nor U2159 (N_2159,In_635,In_53);
and U2160 (N_2160,In_399,In_816);
nand U2161 (N_2161,In_313,In_994);
xnor U2162 (N_2162,In_37,In_280);
nor U2163 (N_2163,In_941,In_796);
and U2164 (N_2164,In_630,In_459);
and U2165 (N_2165,In_632,In_733);
and U2166 (N_2166,In_112,In_45);
or U2167 (N_2167,In_735,In_777);
and U2168 (N_2168,In_412,In_519);
nor U2169 (N_2169,In_299,In_380);
nor U2170 (N_2170,In_29,In_683);
nand U2171 (N_2171,In_330,In_455);
or U2172 (N_2172,In_579,In_661);
and U2173 (N_2173,In_545,In_159);
nor U2174 (N_2174,In_897,In_242);
xnor U2175 (N_2175,In_147,In_13);
nor U2176 (N_2176,In_239,In_652);
nand U2177 (N_2177,In_330,In_533);
or U2178 (N_2178,In_652,In_126);
xor U2179 (N_2179,In_635,In_292);
xor U2180 (N_2180,In_355,In_935);
nand U2181 (N_2181,In_549,In_65);
nand U2182 (N_2182,In_252,In_746);
nand U2183 (N_2183,In_498,In_98);
nand U2184 (N_2184,In_39,In_314);
or U2185 (N_2185,In_875,In_459);
nor U2186 (N_2186,In_383,In_826);
and U2187 (N_2187,In_641,In_686);
or U2188 (N_2188,In_745,In_726);
or U2189 (N_2189,In_438,In_716);
or U2190 (N_2190,In_433,In_353);
nor U2191 (N_2191,In_168,In_710);
or U2192 (N_2192,In_328,In_430);
and U2193 (N_2193,In_550,In_814);
nand U2194 (N_2194,In_502,In_956);
and U2195 (N_2195,In_369,In_30);
nor U2196 (N_2196,In_620,In_898);
nand U2197 (N_2197,In_602,In_421);
nand U2198 (N_2198,In_6,In_718);
and U2199 (N_2199,In_220,In_969);
and U2200 (N_2200,In_323,In_276);
or U2201 (N_2201,In_346,In_658);
or U2202 (N_2202,In_734,In_425);
nand U2203 (N_2203,In_86,In_816);
or U2204 (N_2204,In_165,In_580);
nand U2205 (N_2205,In_465,In_719);
nand U2206 (N_2206,In_992,In_401);
or U2207 (N_2207,In_419,In_847);
nor U2208 (N_2208,In_141,In_340);
nand U2209 (N_2209,In_89,In_370);
nand U2210 (N_2210,In_466,In_65);
nand U2211 (N_2211,In_188,In_792);
nand U2212 (N_2212,In_405,In_486);
nor U2213 (N_2213,In_150,In_998);
nor U2214 (N_2214,In_673,In_7);
nand U2215 (N_2215,In_308,In_123);
and U2216 (N_2216,In_507,In_691);
or U2217 (N_2217,In_771,In_275);
and U2218 (N_2218,In_887,In_228);
and U2219 (N_2219,In_710,In_240);
xor U2220 (N_2220,In_870,In_674);
nor U2221 (N_2221,In_664,In_29);
nand U2222 (N_2222,In_558,In_908);
nor U2223 (N_2223,In_897,In_404);
and U2224 (N_2224,In_958,In_380);
and U2225 (N_2225,In_33,In_265);
nand U2226 (N_2226,In_772,In_454);
nand U2227 (N_2227,In_945,In_592);
nand U2228 (N_2228,In_601,In_523);
nand U2229 (N_2229,In_714,In_558);
xnor U2230 (N_2230,In_754,In_303);
nor U2231 (N_2231,In_624,In_159);
and U2232 (N_2232,In_56,In_373);
and U2233 (N_2233,In_445,In_490);
and U2234 (N_2234,In_536,In_549);
xnor U2235 (N_2235,In_374,In_566);
nand U2236 (N_2236,In_748,In_872);
or U2237 (N_2237,In_962,In_246);
xor U2238 (N_2238,In_943,In_28);
xor U2239 (N_2239,In_770,In_271);
xnor U2240 (N_2240,In_261,In_825);
and U2241 (N_2241,In_639,In_882);
or U2242 (N_2242,In_351,In_901);
or U2243 (N_2243,In_864,In_148);
and U2244 (N_2244,In_877,In_0);
or U2245 (N_2245,In_717,In_471);
nand U2246 (N_2246,In_961,In_981);
nor U2247 (N_2247,In_266,In_584);
nand U2248 (N_2248,In_515,In_484);
nand U2249 (N_2249,In_874,In_87);
nor U2250 (N_2250,In_463,In_769);
nor U2251 (N_2251,In_141,In_424);
or U2252 (N_2252,In_41,In_387);
xnor U2253 (N_2253,In_970,In_913);
or U2254 (N_2254,In_38,In_895);
nor U2255 (N_2255,In_677,In_880);
nand U2256 (N_2256,In_502,In_852);
and U2257 (N_2257,In_507,In_434);
or U2258 (N_2258,In_522,In_842);
nand U2259 (N_2259,In_962,In_169);
nor U2260 (N_2260,In_335,In_172);
and U2261 (N_2261,In_804,In_987);
or U2262 (N_2262,In_682,In_138);
and U2263 (N_2263,In_776,In_673);
xnor U2264 (N_2264,In_478,In_857);
nand U2265 (N_2265,In_787,In_5);
nor U2266 (N_2266,In_808,In_488);
nand U2267 (N_2267,In_73,In_713);
nand U2268 (N_2268,In_78,In_377);
xor U2269 (N_2269,In_594,In_728);
nor U2270 (N_2270,In_892,In_711);
nor U2271 (N_2271,In_199,In_657);
or U2272 (N_2272,In_207,In_904);
and U2273 (N_2273,In_629,In_620);
and U2274 (N_2274,In_741,In_29);
nand U2275 (N_2275,In_160,In_480);
nor U2276 (N_2276,In_588,In_877);
and U2277 (N_2277,In_78,In_815);
nand U2278 (N_2278,In_338,In_389);
nand U2279 (N_2279,In_238,In_329);
nand U2280 (N_2280,In_123,In_904);
or U2281 (N_2281,In_762,In_989);
nor U2282 (N_2282,In_890,In_433);
nor U2283 (N_2283,In_947,In_378);
nor U2284 (N_2284,In_50,In_253);
nand U2285 (N_2285,In_826,In_715);
xnor U2286 (N_2286,In_768,In_890);
nor U2287 (N_2287,In_700,In_960);
nand U2288 (N_2288,In_307,In_299);
or U2289 (N_2289,In_145,In_993);
and U2290 (N_2290,In_814,In_450);
nand U2291 (N_2291,In_287,In_116);
nand U2292 (N_2292,In_546,In_633);
or U2293 (N_2293,In_816,In_240);
or U2294 (N_2294,In_261,In_913);
and U2295 (N_2295,In_298,In_249);
nand U2296 (N_2296,In_308,In_310);
or U2297 (N_2297,In_37,In_869);
nor U2298 (N_2298,In_809,In_625);
and U2299 (N_2299,In_254,In_314);
and U2300 (N_2300,In_623,In_534);
nor U2301 (N_2301,In_478,In_795);
or U2302 (N_2302,In_289,In_609);
nand U2303 (N_2303,In_372,In_895);
nand U2304 (N_2304,In_531,In_930);
and U2305 (N_2305,In_467,In_431);
nor U2306 (N_2306,In_45,In_367);
nor U2307 (N_2307,In_612,In_500);
and U2308 (N_2308,In_257,In_442);
nor U2309 (N_2309,In_170,In_905);
nor U2310 (N_2310,In_454,In_981);
nand U2311 (N_2311,In_181,In_349);
nor U2312 (N_2312,In_791,In_785);
and U2313 (N_2313,In_715,In_34);
nor U2314 (N_2314,In_16,In_828);
nand U2315 (N_2315,In_159,In_216);
or U2316 (N_2316,In_334,In_127);
or U2317 (N_2317,In_800,In_212);
and U2318 (N_2318,In_973,In_855);
xnor U2319 (N_2319,In_774,In_65);
or U2320 (N_2320,In_388,In_935);
and U2321 (N_2321,In_733,In_980);
nand U2322 (N_2322,In_476,In_637);
and U2323 (N_2323,In_168,In_194);
nand U2324 (N_2324,In_712,In_151);
or U2325 (N_2325,In_780,In_595);
or U2326 (N_2326,In_292,In_288);
nor U2327 (N_2327,In_582,In_309);
and U2328 (N_2328,In_590,In_745);
nand U2329 (N_2329,In_772,In_555);
nor U2330 (N_2330,In_903,In_34);
or U2331 (N_2331,In_552,In_299);
nand U2332 (N_2332,In_288,In_814);
nand U2333 (N_2333,In_822,In_716);
nor U2334 (N_2334,In_973,In_46);
nand U2335 (N_2335,In_266,In_300);
and U2336 (N_2336,In_66,In_910);
xnor U2337 (N_2337,In_429,In_333);
or U2338 (N_2338,In_975,In_983);
nand U2339 (N_2339,In_92,In_986);
nand U2340 (N_2340,In_485,In_257);
nor U2341 (N_2341,In_849,In_563);
xor U2342 (N_2342,In_997,In_388);
nor U2343 (N_2343,In_980,In_208);
and U2344 (N_2344,In_168,In_907);
or U2345 (N_2345,In_104,In_79);
or U2346 (N_2346,In_749,In_601);
xnor U2347 (N_2347,In_986,In_47);
and U2348 (N_2348,In_568,In_584);
or U2349 (N_2349,In_820,In_898);
or U2350 (N_2350,In_346,In_200);
nand U2351 (N_2351,In_416,In_544);
or U2352 (N_2352,In_249,In_840);
nand U2353 (N_2353,In_857,In_506);
nor U2354 (N_2354,In_854,In_257);
and U2355 (N_2355,In_435,In_272);
and U2356 (N_2356,In_851,In_525);
and U2357 (N_2357,In_317,In_398);
nor U2358 (N_2358,In_944,In_9);
and U2359 (N_2359,In_57,In_14);
nand U2360 (N_2360,In_104,In_706);
nand U2361 (N_2361,In_191,In_388);
or U2362 (N_2362,In_380,In_263);
and U2363 (N_2363,In_200,In_202);
and U2364 (N_2364,In_209,In_483);
or U2365 (N_2365,In_898,In_601);
or U2366 (N_2366,In_670,In_32);
xor U2367 (N_2367,In_927,In_996);
and U2368 (N_2368,In_124,In_826);
nor U2369 (N_2369,In_264,In_5);
or U2370 (N_2370,In_853,In_186);
nand U2371 (N_2371,In_936,In_216);
and U2372 (N_2372,In_348,In_506);
nand U2373 (N_2373,In_464,In_735);
or U2374 (N_2374,In_235,In_47);
nand U2375 (N_2375,In_266,In_579);
nor U2376 (N_2376,In_561,In_378);
and U2377 (N_2377,In_437,In_504);
nand U2378 (N_2378,In_896,In_691);
or U2379 (N_2379,In_40,In_827);
and U2380 (N_2380,In_682,In_196);
xor U2381 (N_2381,In_875,In_330);
nand U2382 (N_2382,In_604,In_523);
nand U2383 (N_2383,In_821,In_159);
nand U2384 (N_2384,In_800,In_565);
nor U2385 (N_2385,In_167,In_972);
nand U2386 (N_2386,In_857,In_147);
nand U2387 (N_2387,In_102,In_290);
xor U2388 (N_2388,In_433,In_573);
nor U2389 (N_2389,In_554,In_905);
and U2390 (N_2390,In_858,In_674);
nand U2391 (N_2391,In_178,In_825);
or U2392 (N_2392,In_930,In_855);
nand U2393 (N_2393,In_413,In_414);
and U2394 (N_2394,In_600,In_668);
nor U2395 (N_2395,In_731,In_923);
nand U2396 (N_2396,In_348,In_143);
nor U2397 (N_2397,In_380,In_151);
or U2398 (N_2398,In_95,In_816);
and U2399 (N_2399,In_26,In_259);
or U2400 (N_2400,In_157,In_125);
nor U2401 (N_2401,In_928,In_205);
or U2402 (N_2402,In_567,In_766);
nand U2403 (N_2403,In_847,In_166);
nand U2404 (N_2404,In_507,In_100);
or U2405 (N_2405,In_504,In_355);
xor U2406 (N_2406,In_708,In_371);
and U2407 (N_2407,In_369,In_157);
nor U2408 (N_2408,In_107,In_200);
nand U2409 (N_2409,In_438,In_481);
nand U2410 (N_2410,In_739,In_389);
xnor U2411 (N_2411,In_525,In_49);
and U2412 (N_2412,In_749,In_228);
nor U2413 (N_2413,In_19,In_787);
nand U2414 (N_2414,In_230,In_865);
nand U2415 (N_2415,In_123,In_332);
or U2416 (N_2416,In_245,In_113);
or U2417 (N_2417,In_772,In_883);
nor U2418 (N_2418,In_280,In_917);
and U2419 (N_2419,In_477,In_587);
nor U2420 (N_2420,In_94,In_941);
nand U2421 (N_2421,In_947,In_905);
and U2422 (N_2422,In_151,In_55);
nor U2423 (N_2423,In_490,In_108);
nor U2424 (N_2424,In_2,In_41);
nand U2425 (N_2425,In_160,In_658);
nor U2426 (N_2426,In_367,In_292);
xnor U2427 (N_2427,In_450,In_270);
nor U2428 (N_2428,In_872,In_640);
nand U2429 (N_2429,In_350,In_434);
or U2430 (N_2430,In_115,In_773);
xnor U2431 (N_2431,In_730,In_240);
and U2432 (N_2432,In_654,In_72);
nor U2433 (N_2433,In_424,In_808);
nand U2434 (N_2434,In_298,In_138);
and U2435 (N_2435,In_910,In_987);
nand U2436 (N_2436,In_180,In_749);
nand U2437 (N_2437,In_611,In_700);
and U2438 (N_2438,In_936,In_874);
or U2439 (N_2439,In_638,In_969);
or U2440 (N_2440,In_178,In_9);
nand U2441 (N_2441,In_404,In_20);
and U2442 (N_2442,In_113,In_66);
nand U2443 (N_2443,In_191,In_760);
nand U2444 (N_2444,In_962,In_226);
or U2445 (N_2445,In_480,In_204);
and U2446 (N_2446,In_660,In_875);
nor U2447 (N_2447,In_682,In_5);
or U2448 (N_2448,In_893,In_372);
and U2449 (N_2449,In_389,In_1);
nor U2450 (N_2450,In_331,In_49);
xor U2451 (N_2451,In_63,In_239);
xnor U2452 (N_2452,In_183,In_657);
xnor U2453 (N_2453,In_599,In_144);
nor U2454 (N_2454,In_606,In_27);
nand U2455 (N_2455,In_531,In_867);
and U2456 (N_2456,In_134,In_493);
or U2457 (N_2457,In_113,In_42);
nor U2458 (N_2458,In_955,In_994);
nand U2459 (N_2459,In_852,In_914);
nor U2460 (N_2460,In_493,In_522);
nor U2461 (N_2461,In_607,In_654);
and U2462 (N_2462,In_775,In_877);
nor U2463 (N_2463,In_179,In_957);
and U2464 (N_2464,In_589,In_937);
nand U2465 (N_2465,In_41,In_282);
nand U2466 (N_2466,In_118,In_476);
nand U2467 (N_2467,In_448,In_246);
and U2468 (N_2468,In_341,In_842);
nor U2469 (N_2469,In_334,In_715);
or U2470 (N_2470,In_746,In_268);
or U2471 (N_2471,In_911,In_640);
or U2472 (N_2472,In_817,In_377);
and U2473 (N_2473,In_903,In_7);
nand U2474 (N_2474,In_401,In_265);
xor U2475 (N_2475,In_590,In_633);
nand U2476 (N_2476,In_474,In_309);
or U2477 (N_2477,In_962,In_398);
or U2478 (N_2478,In_943,In_833);
nor U2479 (N_2479,In_688,In_530);
xor U2480 (N_2480,In_32,In_909);
or U2481 (N_2481,In_522,In_906);
nand U2482 (N_2482,In_93,In_863);
or U2483 (N_2483,In_615,In_135);
nor U2484 (N_2484,In_640,In_408);
nor U2485 (N_2485,In_522,In_415);
nand U2486 (N_2486,In_614,In_777);
nand U2487 (N_2487,In_573,In_468);
and U2488 (N_2488,In_710,In_872);
or U2489 (N_2489,In_628,In_725);
and U2490 (N_2490,In_6,In_117);
nand U2491 (N_2491,In_225,In_236);
or U2492 (N_2492,In_211,In_372);
or U2493 (N_2493,In_108,In_603);
and U2494 (N_2494,In_665,In_817);
nand U2495 (N_2495,In_163,In_654);
and U2496 (N_2496,In_242,In_806);
xor U2497 (N_2497,In_694,In_219);
and U2498 (N_2498,In_667,In_835);
nand U2499 (N_2499,In_594,In_378);
and U2500 (N_2500,N_1380,N_1528);
or U2501 (N_2501,N_2250,N_1044);
nor U2502 (N_2502,N_1319,N_421);
nor U2503 (N_2503,N_1767,N_2307);
and U2504 (N_2504,N_471,N_1702);
xnor U2505 (N_2505,N_2458,N_899);
nand U2506 (N_2506,N_1155,N_857);
and U2507 (N_2507,N_1193,N_93);
or U2508 (N_2508,N_1845,N_3);
nor U2509 (N_2509,N_1101,N_2262);
nor U2510 (N_2510,N_1343,N_55);
or U2511 (N_2511,N_2409,N_2478);
or U2512 (N_2512,N_1909,N_218);
xor U2513 (N_2513,N_2203,N_1456);
nand U2514 (N_2514,N_2328,N_1653);
nand U2515 (N_2515,N_1925,N_306);
nand U2516 (N_2516,N_952,N_169);
nand U2517 (N_2517,N_1102,N_1640);
or U2518 (N_2518,N_476,N_1849);
or U2519 (N_2519,N_2047,N_791);
nand U2520 (N_2520,N_1360,N_2255);
nand U2521 (N_2521,N_1546,N_2287);
or U2522 (N_2522,N_1554,N_567);
or U2523 (N_2523,N_51,N_189);
nand U2524 (N_2524,N_372,N_1932);
nor U2525 (N_2525,N_959,N_2393);
nand U2526 (N_2526,N_2322,N_950);
and U2527 (N_2527,N_2156,N_1612);
xor U2528 (N_2528,N_124,N_1074);
nand U2529 (N_2529,N_2312,N_406);
and U2530 (N_2530,N_788,N_1938);
or U2531 (N_2531,N_1591,N_1782);
nand U2532 (N_2532,N_580,N_1210);
and U2533 (N_2533,N_1561,N_2043);
nand U2534 (N_2534,N_991,N_1841);
nor U2535 (N_2535,N_804,N_40);
and U2536 (N_2536,N_1179,N_2069);
and U2537 (N_2537,N_2329,N_840);
and U2538 (N_2538,N_1971,N_1658);
xor U2539 (N_2539,N_947,N_2389);
nand U2540 (N_2540,N_2179,N_2023);
xnor U2541 (N_2541,N_828,N_2057);
and U2542 (N_2542,N_818,N_311);
or U2543 (N_2543,N_2116,N_996);
nand U2544 (N_2544,N_2463,N_803);
and U2545 (N_2545,N_258,N_1355);
and U2546 (N_2546,N_1792,N_909);
nand U2547 (N_2547,N_533,N_822);
nand U2548 (N_2548,N_1933,N_446);
xnor U2549 (N_2549,N_934,N_1391);
or U2550 (N_2550,N_271,N_482);
and U2551 (N_2551,N_700,N_1454);
and U2552 (N_2552,N_958,N_1259);
and U2553 (N_2553,N_1347,N_1182);
nand U2554 (N_2554,N_326,N_1085);
and U2555 (N_2555,N_1489,N_2239);
or U2556 (N_2556,N_1007,N_1382);
nor U2557 (N_2557,N_1296,N_2192);
nand U2558 (N_2558,N_2146,N_727);
or U2559 (N_2559,N_1698,N_1649);
nand U2560 (N_2560,N_585,N_1378);
or U2561 (N_2561,N_252,N_2451);
or U2562 (N_2562,N_759,N_154);
or U2563 (N_2563,N_535,N_1293);
xor U2564 (N_2564,N_2141,N_1566);
and U2565 (N_2565,N_962,N_355);
or U2566 (N_2566,N_1225,N_1395);
and U2567 (N_2567,N_1599,N_612);
xnor U2568 (N_2568,N_2035,N_2194);
or U2569 (N_2569,N_1854,N_2034);
nand U2570 (N_2570,N_2437,N_763);
nor U2571 (N_2571,N_1969,N_1756);
and U2572 (N_2572,N_356,N_809);
or U2573 (N_2573,N_1681,N_88);
nor U2574 (N_2574,N_590,N_855);
nor U2575 (N_2575,N_1470,N_1757);
and U2576 (N_2576,N_1864,N_1384);
nand U2577 (N_2577,N_1537,N_1967);
and U2578 (N_2578,N_2177,N_96);
or U2579 (N_2579,N_1831,N_1688);
nand U2580 (N_2580,N_1582,N_1577);
xor U2581 (N_2581,N_1981,N_1132);
and U2582 (N_2582,N_308,N_911);
nor U2583 (N_2583,N_1066,N_1423);
or U2584 (N_2584,N_1677,N_1705);
nand U2585 (N_2585,N_2219,N_550);
or U2586 (N_2586,N_2425,N_2433);
nor U2587 (N_2587,N_2176,N_2137);
nor U2588 (N_2588,N_552,N_466);
xnor U2589 (N_2589,N_1374,N_1247);
and U2590 (N_2590,N_2446,N_536);
and U2591 (N_2591,N_41,N_2016);
nor U2592 (N_2592,N_2324,N_2435);
and U2593 (N_2593,N_725,N_1533);
and U2594 (N_2594,N_1913,N_181);
and U2595 (N_2595,N_1338,N_350);
nor U2596 (N_2596,N_1467,N_891);
and U2597 (N_2597,N_92,N_2229);
or U2598 (N_2598,N_383,N_2046);
nand U2599 (N_2599,N_2481,N_2450);
or U2600 (N_2600,N_1987,N_1885);
xor U2601 (N_2601,N_1742,N_1991);
or U2602 (N_2602,N_1960,N_1890);
or U2603 (N_2603,N_1755,N_916);
nor U2604 (N_2604,N_1483,N_246);
or U2605 (N_2605,N_1594,N_2222);
or U2606 (N_2606,N_2292,N_1112);
nand U2607 (N_2607,N_2431,N_904);
or U2608 (N_2608,N_754,N_1156);
or U2609 (N_2609,N_301,N_1200);
or U2610 (N_2610,N_1766,N_1060);
nand U2611 (N_2611,N_1027,N_1258);
xnor U2612 (N_2612,N_1696,N_1006);
nor U2613 (N_2613,N_2368,N_474);
nor U2614 (N_2614,N_87,N_858);
or U2615 (N_2615,N_213,N_2007);
nor U2616 (N_2616,N_1114,N_640);
xor U2617 (N_2617,N_1525,N_2215);
and U2618 (N_2618,N_1813,N_795);
or U2619 (N_2619,N_173,N_478);
and U2620 (N_2620,N_2358,N_1486);
and U2621 (N_2621,N_1254,N_2012);
nor U2622 (N_2622,N_2126,N_297);
nor U2623 (N_2623,N_2140,N_691);
or U2624 (N_2624,N_522,N_842);
nand U2625 (N_2625,N_902,N_706);
and U2626 (N_2626,N_1405,N_2442);
or U2627 (N_2627,N_1096,N_2441);
xnor U2628 (N_2628,N_978,N_453);
nor U2629 (N_2629,N_2074,N_1117);
nand U2630 (N_2630,N_465,N_2482);
xnor U2631 (N_2631,N_2273,N_1772);
or U2632 (N_2632,N_2489,N_101);
nor U2633 (N_2633,N_1059,N_582);
nand U2634 (N_2634,N_267,N_658);
nand U2635 (N_2635,N_382,N_562);
and U2636 (N_2636,N_1219,N_2171);
or U2637 (N_2637,N_86,N_1778);
and U2638 (N_2638,N_2211,N_666);
and U2639 (N_2639,N_643,N_994);
xor U2640 (N_2640,N_678,N_1671);
and U2641 (N_2641,N_2336,N_313);
nor U2642 (N_2642,N_1553,N_2295);
nor U2643 (N_2643,N_1260,N_58);
or U2644 (N_2644,N_821,N_519);
or U2645 (N_2645,N_2420,N_2495);
nand U2646 (N_2646,N_1387,N_456);
nand U2647 (N_2647,N_829,N_1003);
xnor U2648 (N_2648,N_1680,N_1793);
nor U2649 (N_2649,N_264,N_1507);
nand U2650 (N_2650,N_128,N_1125);
nor U2651 (N_2651,N_1383,N_1004);
nor U2652 (N_2652,N_2131,N_506);
nand U2653 (N_2653,N_990,N_2468);
and U2654 (N_2654,N_1603,N_2319);
and U2655 (N_2655,N_1359,N_1522);
xnor U2656 (N_2656,N_1307,N_45);
nand U2657 (N_2657,N_427,N_1021);
nor U2658 (N_2658,N_2004,N_284);
nand U2659 (N_2659,N_789,N_2053);
and U2660 (N_2660,N_2209,N_2108);
and U2661 (N_2661,N_1945,N_2300);
and U2662 (N_2662,N_376,N_420);
nand U2663 (N_2663,N_867,N_229);
and U2664 (N_2664,N_749,N_896);
or U2665 (N_2665,N_1737,N_273);
nor U2666 (N_2666,N_1284,N_254);
nand U2667 (N_2667,N_1833,N_238);
or U2668 (N_2668,N_1840,N_2228);
or U2669 (N_2669,N_1328,N_2129);
nor U2670 (N_2670,N_1189,N_660);
or U2671 (N_2671,N_1823,N_1278);
nor U2672 (N_2672,N_2284,N_508);
or U2673 (N_2673,N_275,N_2357);
nor U2674 (N_2674,N_1245,N_1542);
nand U2675 (N_2675,N_1076,N_1419);
nand U2676 (N_2676,N_647,N_1207);
nand U2677 (N_2677,N_2460,N_1272);
nand U2678 (N_2678,N_1973,N_1334);
nand U2679 (N_2679,N_1398,N_665);
or U2680 (N_2680,N_1955,N_1131);
and U2681 (N_2681,N_1053,N_620);
nand U2682 (N_2682,N_2,N_94);
or U2683 (N_2683,N_852,N_115);
nand U2684 (N_2684,N_1738,N_982);
nor U2685 (N_2685,N_1313,N_462);
and U2686 (N_2686,N_831,N_433);
nor U2687 (N_2687,N_1999,N_1265);
nor U2688 (N_2688,N_27,N_2380);
nor U2689 (N_2689,N_1493,N_1013);
nor U2690 (N_2690,N_1220,N_1298);
nor U2691 (N_2691,N_1113,N_2052);
nor U2692 (N_2692,N_425,N_1320);
xnor U2693 (N_2693,N_1572,N_20);
nor U2694 (N_2694,N_227,N_1828);
or U2695 (N_2695,N_1867,N_1838);
or U2696 (N_2696,N_1351,N_2220);
nand U2697 (N_2697,N_339,N_89);
nand U2698 (N_2698,N_419,N_980);
nand U2699 (N_2699,N_680,N_143);
nand U2700 (N_2700,N_48,N_1993);
nor U2701 (N_2701,N_460,N_2280);
or U2702 (N_2702,N_1550,N_2373);
nand U2703 (N_2703,N_1455,N_2354);
and U2704 (N_2704,N_1379,N_1409);
nor U2705 (N_2705,N_1396,N_2275);
xor U2706 (N_2706,N_1226,N_1954);
xor U2707 (N_2707,N_610,N_956);
nand U2708 (N_2708,N_895,N_1115);
and U2709 (N_2709,N_1237,N_695);
or U2710 (N_2710,N_1267,N_1883);
nand U2711 (N_2711,N_1228,N_613);
or U2712 (N_2712,N_2241,N_25);
or U2713 (N_2713,N_2498,N_2430);
nor U2714 (N_2714,N_1604,N_2288);
xor U2715 (N_2715,N_1055,N_677);
or U2716 (N_2716,N_1301,N_158);
nor U2717 (N_2717,N_540,N_2163);
and U2718 (N_2718,N_817,N_200);
xor U2719 (N_2719,N_2318,N_1326);
nor U2720 (N_2720,N_6,N_927);
or U2721 (N_2721,N_2417,N_1386);
nand U2722 (N_2722,N_1090,N_1161);
nor U2723 (N_2723,N_1305,N_1795);
nor U2724 (N_2724,N_558,N_1961);
nor U2725 (N_2725,N_2419,N_1408);
and U2726 (N_2726,N_1562,N_2279);
nor U2727 (N_2727,N_1997,N_312);
and U2728 (N_2728,N_1468,N_679);
nor U2729 (N_2729,N_1708,N_2310);
nor U2730 (N_2730,N_467,N_127);
nand U2731 (N_2731,N_987,N_629);
and U2732 (N_2732,N_2369,N_703);
or U2733 (N_2733,N_1729,N_2118);
nor U2734 (N_2734,N_168,N_1884);
nor U2735 (N_2735,N_464,N_1116);
nor U2736 (N_2736,N_514,N_192);
nor U2737 (N_2737,N_215,N_2344);
xnor U2738 (N_2738,N_1484,N_1643);
and U2739 (N_2739,N_2413,N_1881);
nand U2740 (N_2740,N_166,N_65);
or U2741 (N_2741,N_1299,N_515);
nor U2742 (N_2742,N_1682,N_1903);
and U2743 (N_2743,N_918,N_1679);
or U2744 (N_2744,N_1229,N_131);
nand U2745 (N_2745,N_716,N_929);
nand U2746 (N_2746,N_1356,N_2302);
nand U2747 (N_2747,N_872,N_1184);
nand U2748 (N_2748,N_1816,N_396);
or U2749 (N_2749,N_2375,N_2038);
or U2750 (N_2750,N_1518,N_177);
xnor U2751 (N_2751,N_2355,N_882);
nand U2752 (N_2752,N_1928,N_413);
nand U2753 (N_2753,N_577,N_1151);
xor U2754 (N_2754,N_979,N_2119);
nor U2755 (N_2755,N_1201,N_2236);
and U2756 (N_2756,N_757,N_1404);
or U2757 (N_2757,N_72,N_1835);
xnor U2758 (N_2758,N_747,N_1982);
and U2759 (N_2759,N_901,N_925);
and U2760 (N_2760,N_2376,N_365);
or U2761 (N_2761,N_1972,N_2338);
nand U2762 (N_2762,N_1690,N_1370);
nand U2763 (N_2763,N_224,N_2252);
nand U2764 (N_2764,N_995,N_1771);
nand U2765 (N_2765,N_167,N_750);
nor U2766 (N_2766,N_729,N_1316);
nor U2767 (N_2767,N_2415,N_894);
nor U2768 (N_2768,N_1930,N_2234);
and U2769 (N_2769,N_1709,N_1803);
nor U2770 (N_2770,N_240,N_2031);
nor U2771 (N_2771,N_1610,N_1631);
or U2772 (N_2772,N_1908,N_863);
and U2773 (N_2773,N_1722,N_1819);
xor U2774 (N_2774,N_2165,N_1744);
nor U2775 (N_2775,N_208,N_1695);
nand U2776 (N_2776,N_854,N_2400);
xnor U2777 (N_2777,N_330,N_1887);
xnor U2778 (N_2778,N_1984,N_2121);
nand U2779 (N_2779,N_178,N_1820);
nand U2780 (N_2780,N_2408,N_305);
nand U2781 (N_2781,N_2251,N_216);
and U2782 (N_2782,N_371,N_718);
and U2783 (N_2783,N_1980,N_575);
nand U2784 (N_2784,N_307,N_323);
and U2785 (N_2785,N_1432,N_2485);
and U2786 (N_2786,N_2340,N_2390);
or U2787 (N_2787,N_2080,N_837);
or U2788 (N_2788,N_1691,N_1148);
and U2789 (N_2789,N_2225,N_1595);
and U2790 (N_2790,N_1894,N_1907);
and U2791 (N_2791,N_283,N_1152);
nand U2792 (N_2792,N_1145,N_555);
nor U2793 (N_2793,N_2257,N_2217);
and U2794 (N_2794,N_1882,N_1635);
nand U2795 (N_2795,N_199,N_602);
xor U2796 (N_2796,N_162,N_2351);
nor U2797 (N_2797,N_928,N_887);
or U2798 (N_2798,N_1246,N_1661);
or U2799 (N_2799,N_1327,N_1936);
xnor U2800 (N_2800,N_1585,N_1989);
nor U2801 (N_2801,N_457,N_607);
and U2802 (N_2802,N_1271,N_2378);
or U2803 (N_2803,N_1964,N_251);
or U2804 (N_2804,N_874,N_211);
and U2805 (N_2805,N_1567,N_1812);
nor U2806 (N_2806,N_1336,N_2127);
or U2807 (N_2807,N_1652,N_1983);
nor U2808 (N_2808,N_1593,N_416);
nand U2809 (N_2809,N_1811,N_487);
or U2810 (N_2810,N_1922,N_2055);
nand U2811 (N_2811,N_1367,N_391);
xnor U2812 (N_2812,N_2411,N_2144);
nor U2813 (N_2813,N_2049,N_1762);
and U2814 (N_2814,N_185,N_1769);
nand U2815 (N_2815,N_654,N_614);
nor U2816 (N_2816,N_304,N_1285);
and U2817 (N_2817,N_29,N_1233);
nand U2818 (N_2818,N_2469,N_1977);
nor U2819 (N_2819,N_2175,N_2405);
or U2820 (N_2820,N_1552,N_960);
nand U2821 (N_2821,N_2439,N_1634);
or U2822 (N_2822,N_1269,N_1150);
nand U2823 (N_2823,N_1712,N_1439);
nor U2824 (N_2824,N_2073,N_1166);
nor U2825 (N_2825,N_1037,N_1821);
nand U2826 (N_2826,N_2346,N_2032);
and U2827 (N_2827,N_286,N_770);
and U2828 (N_2828,N_864,N_2095);
or U2829 (N_2829,N_572,N_1477);
nand U2830 (N_2830,N_799,N_75);
nand U2831 (N_2831,N_1213,N_34);
nor U2832 (N_2832,N_983,N_2014);
nor U2833 (N_2833,N_46,N_2083);
nor U2834 (N_2834,N_1401,N_1734);
and U2835 (N_2835,N_944,N_182);
or U2836 (N_2836,N_1354,N_2153);
nor U2837 (N_2837,N_21,N_2470);
xnor U2838 (N_2838,N_611,N_1944);
nand U2839 (N_2839,N_2428,N_1753);
and U2840 (N_2840,N_1789,N_2051);
or U2841 (N_2841,N_1222,N_1672);
nor U2842 (N_2842,N_792,N_111);
or U2843 (N_2843,N_191,N_2311);
or U2844 (N_2844,N_1720,N_400);
or U2845 (N_2845,N_1082,N_1797);
nand U2846 (N_2846,N_986,N_1199);
and U2847 (N_2847,N_2396,N_2407);
nand U2848 (N_2848,N_624,N_714);
nand U2849 (N_2849,N_917,N_1331);
and U2850 (N_2850,N_123,N_2476);
and U2851 (N_2851,N_1375,N_1776);
nor U2852 (N_2852,N_1045,N_1586);
xor U2853 (N_2853,N_1279,N_1503);
and U2854 (N_2854,N_935,N_1346);
nand U2855 (N_2855,N_84,N_2399);
xnor U2856 (N_2856,N_1363,N_1565);
nand U2857 (N_2857,N_1646,N_249);
nor U2858 (N_2858,N_395,N_890);
and U2859 (N_2859,N_2427,N_367);
nor U2860 (N_2860,N_847,N_2436);
nand U2861 (N_2861,N_1312,N_593);
nor U2862 (N_2862,N_912,N_507);
and U2863 (N_2863,N_539,N_2459);
nand U2864 (N_2864,N_1399,N_1995);
or U2865 (N_2865,N_1668,N_2005);
nor U2866 (N_2866,N_1948,N_317);
nand U2867 (N_2867,N_1574,N_1073);
and U2868 (N_2868,N_988,N_970);
nand U2869 (N_2869,N_31,N_2044);
nand U2870 (N_2870,N_2210,N_1711);
nand U2871 (N_2871,N_1119,N_2105);
or U2872 (N_2872,N_188,N_1715);
nor U2873 (N_2873,N_2013,N_1422);
nor U2874 (N_2874,N_352,N_2356);
nor U2875 (N_2875,N_1424,N_2199);
xor U2876 (N_2876,N_739,N_941);
or U2877 (N_2877,N_79,N_1524);
nand U2878 (N_2878,N_2438,N_878);
or U2879 (N_2879,N_1025,N_2193);
nor U2880 (N_2880,N_741,N_497);
nand U2881 (N_2881,N_1790,N_2246);
nor U2882 (N_2882,N_99,N_717);
and U2883 (N_2883,N_1875,N_2198);
and U2884 (N_2884,N_209,N_963);
nor U2885 (N_2885,N_541,N_2196);
nand U2886 (N_2886,N_1311,N_576);
nor U2887 (N_2887,N_600,N_2001);
xnor U2888 (N_2888,N_2342,N_566);
nand U2889 (N_2889,N_2135,N_1230);
or U2890 (N_2890,N_2464,N_922);
and U2891 (N_2891,N_2362,N_1569);
nand U2892 (N_2892,N_2041,N_1089);
or U2893 (N_2893,N_135,N_528);
or U2894 (N_2894,N_953,N_898);
nor U2895 (N_2895,N_752,N_573);
nand U2896 (N_2896,N_2071,N_2332);
or U2897 (N_2897,N_2191,N_274);
or U2898 (N_2898,N_850,N_150);
and U2899 (N_2899,N_2372,N_1622);
or U2900 (N_2900,N_2101,N_905);
and U2901 (N_2901,N_97,N_560);
or U2902 (N_2902,N_1613,N_2448);
nand U2903 (N_2903,N_2125,N_325);
and U2904 (N_2904,N_1321,N_268);
nand U2905 (N_2905,N_203,N_1262);
nand U2906 (N_2906,N_961,N_424);
and U2907 (N_2907,N_1041,N_870);
nor U2908 (N_2908,N_33,N_684);
nor U2909 (N_2909,N_1372,N_219);
nand U2910 (N_2910,N_315,N_239);
nor U2911 (N_2911,N_1694,N_2202);
nand U2912 (N_2912,N_1748,N_1557);
nor U2913 (N_2913,N_1763,N_969);
and U2914 (N_2914,N_1825,N_1801);
and U2915 (N_2915,N_2265,N_2124);
and U2916 (N_2916,N_473,N_1487);
and U2917 (N_2917,N_1368,N_1494);
and U2918 (N_2918,N_998,N_2237);
xnor U2919 (N_2919,N_2060,N_2480);
nand U2920 (N_2920,N_1590,N_1261);
xor U2921 (N_2921,N_1764,N_1431);
and U2922 (N_2922,N_1842,N_1086);
nand U2923 (N_2923,N_62,N_556);
xor U2924 (N_2924,N_914,N_1618);
and U2925 (N_2925,N_1440,N_321);
nand U2926 (N_2926,N_800,N_2185);
nor U2927 (N_2927,N_295,N_234);
xor U2928 (N_2928,N_1879,N_2235);
nor U2929 (N_2929,N_2472,N_1015);
or U2930 (N_2930,N_627,N_450);
and U2931 (N_2931,N_888,N_2320);
nor U2932 (N_2932,N_410,N_441);
and U2933 (N_2933,N_2114,N_1685);
nor U2934 (N_2934,N_737,N_631);
nand U2935 (N_2935,N_1335,N_1892);
and U2936 (N_2936,N_699,N_596);
or U2937 (N_2937,N_1527,N_348);
nor U2938 (N_2938,N_592,N_1804);
or U2939 (N_2939,N_155,N_1214);
xnor U2940 (N_2940,N_1072,N_697);
xnor U2941 (N_2941,N_920,N_1880);
and U2942 (N_2942,N_1416,N_28);
and U2943 (N_2943,N_1459,N_2461);
nand U2944 (N_2944,N_938,N_319);
xor U2945 (N_2945,N_784,N_604);
and U2946 (N_2946,N_109,N_2216);
or U2947 (N_2947,N_2024,N_430);
nor U2948 (N_2948,N_1723,N_2084);
and U2949 (N_2949,N_1765,N_309);
xor U2950 (N_2950,N_1923,N_2189);
or U2951 (N_2951,N_1693,N_1);
nor U2952 (N_2952,N_2326,N_1188);
or U2953 (N_2953,N_2155,N_17);
or U2954 (N_2954,N_869,N_136);
nand U2955 (N_2955,N_1515,N_1071);
and U2956 (N_2956,N_586,N_744);
xor U2957 (N_2957,N_1517,N_2077);
nand U2958 (N_2958,N_2264,N_256);
and U2959 (N_2959,N_426,N_357);
xor U2960 (N_2960,N_2113,N_394);
nand U2961 (N_2961,N_1340,N_838);
nor U2962 (N_2962,N_1031,N_2444);
nor U2963 (N_2963,N_1918,N_1232);
nand U2964 (N_2964,N_636,N_906);
and U2965 (N_2965,N_1600,N_1498);
nor U2966 (N_2966,N_1202,N_1787);
nor U2967 (N_2967,N_664,N_2282);
nand U2968 (N_2968,N_1425,N_1822);
or U2969 (N_2969,N_187,N_1240);
or U2970 (N_2970,N_1505,N_322);
xor U2971 (N_2971,N_361,N_1276);
xor U2972 (N_2972,N_1502,N_1290);
nand U2973 (N_2973,N_61,N_10);
or U2974 (N_2974,N_374,N_599);
nor U2975 (N_2975,N_708,N_1413);
nand U2976 (N_2976,N_2467,N_1727);
nand U2977 (N_2977,N_1836,N_1029);
nand U2978 (N_2978,N_1302,N_205);
and U2979 (N_2979,N_1626,N_2120);
nor U2980 (N_2980,N_1236,N_1196);
nor U2981 (N_2981,N_387,N_2314);
nand U2982 (N_2982,N_1065,N_1619);
nand U2983 (N_2983,N_13,N_1728);
or U2984 (N_2984,N_2379,N_530);
or U2985 (N_2985,N_1392,N_14);
nand U2986 (N_2986,N_1531,N_1994);
or U2987 (N_2987,N_183,N_1052);
or U2988 (N_2988,N_1376,N_1942);
or U2989 (N_2989,N_2160,N_1442);
nor U2990 (N_2990,N_1558,N_1446);
nor U2991 (N_2991,N_2187,N_1579);
xnor U2992 (N_2992,N_1627,N_1862);
nand U2993 (N_2993,N_735,N_2245);
and U2994 (N_2994,N_2339,N_1427);
nand U2995 (N_2995,N_704,N_1120);
and U2996 (N_2996,N_2395,N_412);
nand U2997 (N_2997,N_1851,N_1988);
xnor U2998 (N_2998,N_1163,N_242);
nand U2999 (N_2999,N_711,N_1647);
nand U3000 (N_3000,N_226,N_723);
or U3001 (N_3001,N_1480,N_2208);
nand U3002 (N_3002,N_1203,N_1147);
and U3003 (N_3003,N_1926,N_810);
xnor U3004 (N_3004,N_1968,N_1929);
nor U3005 (N_3005,N_1244,N_1443);
nor U3006 (N_3006,N_52,N_223);
xnor U3007 (N_3007,N_1017,N_1775);
or U3008 (N_3008,N_245,N_1655);
nand U3009 (N_3009,N_1578,N_2253);
nand U3010 (N_3010,N_832,N_2152);
and U3011 (N_3011,N_1287,N_2333);
xnor U3012 (N_3012,N_1042,N_674);
and U3013 (N_3013,N_118,N_559);
xor U3014 (N_3014,N_957,N_1807);
nor U3015 (N_3015,N_715,N_2274);
or U3016 (N_3016,N_1718,N_843);
and U3017 (N_3017,N_68,N_534);
and U3018 (N_3018,N_2059,N_2406);
and U3019 (N_3019,N_649,N_2183);
and U3020 (N_3020,N_946,N_434);
and U3021 (N_3021,N_331,N_786);
xnor U3022 (N_3022,N_2094,N_746);
nor U3023 (N_3023,N_919,N_232);
xor U3024 (N_3024,N_477,N_1056);
and U3025 (N_3025,N_1084,N_778);
and U3026 (N_3026,N_1779,N_1539);
or U3027 (N_3027,N_2087,N_2258);
or U3028 (N_3028,N_1630,N_1314);
nor U3029 (N_3029,N_2412,N_1601);
and U3030 (N_3030,N_774,N_2088);
or U3031 (N_3031,N_1014,N_1075);
xor U3032 (N_3032,N_618,N_2487);
and U3033 (N_3033,N_2267,N_2337);
nand U3034 (N_3034,N_2207,N_2254);
xor U3035 (N_3035,N_1817,N_2096);
and U3036 (N_3036,N_1149,N_316);
and U3037 (N_3037,N_1176,N_1448);
or U3038 (N_3038,N_900,N_1496);
xnor U3039 (N_3039,N_1217,N_1270);
nor U3040 (N_3040,N_1221,N_2188);
and U3041 (N_3041,N_1026,N_853);
or U3042 (N_3042,N_145,N_653);
nand U3043 (N_3043,N_548,N_1141);
and U3044 (N_3044,N_504,N_364);
nand U3045 (N_3045,N_2232,N_1280);
nand U3046 (N_3046,N_1212,N_1597);
or U3047 (N_3047,N_351,N_2304);
and U3048 (N_3048,N_243,N_1009);
and U3049 (N_3049,N_1917,N_133);
nand U3050 (N_3050,N_2161,N_1122);
nor U3051 (N_3051,N_411,N_1654);
xor U3052 (N_3052,N_671,N_1592);
xnor U3053 (N_3053,N_2299,N_1450);
nand U3054 (N_3054,N_2499,N_1966);
and U3055 (N_3055,N_939,N_2091);
nand U3056 (N_3056,N_551,N_1295);
nor U3057 (N_3057,N_2082,N_808);
nor U3058 (N_3058,N_363,N_839);
xnor U3059 (N_3059,N_529,N_2491);
nand U3060 (N_3060,N_82,N_1780);
or U3061 (N_3061,N_71,N_965);
and U3062 (N_3062,N_1511,N_2098);
and U3063 (N_3063,N_165,N_543);
nor U3064 (N_3064,N_626,N_1098);
or U3065 (N_3065,N_587,N_2230);
and U3066 (N_3066,N_1128,N_937);
nand U3067 (N_3067,N_104,N_1371);
xnor U3068 (N_3068,N_1645,N_175);
nor U3069 (N_3069,N_332,N_738);
nand U3070 (N_3070,N_1568,N_967);
nor U3071 (N_3071,N_2213,N_1692);
nand U3072 (N_3072,N_1160,N_2382);
or U3073 (N_3073,N_722,N_1436);
or U3074 (N_3074,N_399,N_579);
or U3075 (N_3075,N_972,N_335);
nor U3076 (N_3076,N_1726,N_1407);
nand U3077 (N_3077,N_1426,N_2477);
nand U3078 (N_3078,N_193,N_1008);
or U3079 (N_3079,N_948,N_1167);
nor U3080 (N_3080,N_1717,N_1412);
xor U3081 (N_3081,N_1673,N_1274);
nor U3082 (N_3082,N_1342,N_2449);
nand U3083 (N_3083,N_255,N_334);
xnor U3084 (N_3084,N_404,N_1023);
and U3085 (N_3085,N_1914,N_1636);
or U3086 (N_3086,N_1598,N_1965);
or U3087 (N_3087,N_1081,N_1308);
or U3088 (N_3088,N_1033,N_1956);
and U3089 (N_3089,N_1069,N_2401);
nor U3090 (N_3090,N_1083,N_76);
or U3091 (N_3091,N_105,N_1700);
and U3092 (N_3092,N_381,N_1350);
or U3093 (N_3093,N_1428,N_2037);
nand U3094 (N_3094,N_384,N_1802);
nor U3095 (N_3095,N_1872,N_1277);
xor U3096 (N_3096,N_542,N_1099);
nor U3097 (N_3097,N_897,N_1998);
or U3098 (N_3098,N_921,N_2466);
and U3099 (N_3099,N_1637,N_1135);
nor U3100 (N_3100,N_1941,N_1488);
and U3101 (N_3101,N_1475,N_1154);
nand U3102 (N_3102,N_2190,N_1310);
and U3103 (N_3103,N_270,N_1024);
and U3104 (N_3104,N_1641,N_2045);
nor U3105 (N_3105,N_1747,N_940);
or U3106 (N_3106,N_2475,N_2456);
or U3107 (N_3107,N_646,N_1786);
nand U3108 (N_3108,N_2154,N_1606);
or U3109 (N_3109,N_860,N_2309);
or U3110 (N_3110,N_2117,N_91);
nor U3111 (N_3111,N_873,N_686);
nor U3112 (N_3112,N_1478,N_231);
nor U3113 (N_3113,N_1457,N_1241);
and U3114 (N_3114,N_1286,N_1758);
and U3115 (N_3115,N_802,N_1874);
or U3116 (N_3116,N_617,N_222);
nor U3117 (N_3117,N_1444,N_945);
nand U3118 (N_3118,N_1068,N_1759);
or U3119 (N_3119,N_1251,N_2200);
nand U3120 (N_3120,N_2316,N_2128);
nor U3121 (N_3121,N_2266,N_1902);
nand U3122 (N_3122,N_1019,N_1011);
or U3123 (N_3123,N_1548,N_2164);
and U3124 (N_3124,N_1571,N_23);
nand U3125 (N_3125,N_1741,N_1341);
nand U3126 (N_3126,N_1106,N_632);
nor U3127 (N_3127,N_1855,N_1458);
nand U3128 (N_3128,N_1050,N_510);
or U3129 (N_3129,N_1940,N_1364);
or U3130 (N_3130,N_140,N_824);
nor U3131 (N_3131,N_493,N_236);
nand U3132 (N_3132,N_2350,N_2133);
nand U3133 (N_3133,N_2454,N_2367);
and U3134 (N_3134,N_152,N_1893);
nand U3135 (N_3135,N_2112,N_2102);
nor U3136 (N_3136,N_369,N_418);
nor U3137 (N_3137,N_2138,N_2147);
xor U3138 (N_3138,N_1877,N_221);
or U3139 (N_3139,N_1224,N_1231);
nand U3140 (N_3140,N_574,N_877);
or U3141 (N_3141,N_2040,N_2042);
and U3142 (N_3142,N_324,N_176);
nand U3143 (N_3143,N_210,N_414);
nand U3144 (N_3144,N_380,N_661);
nor U3145 (N_3145,N_100,N_125);
nand U3146 (N_3146,N_688,N_915);
nand U3147 (N_3147,N_1949,N_112);
and U3148 (N_3148,N_1876,N_1197);
and U3149 (N_3149,N_2157,N_1891);
nor U3150 (N_3150,N_830,N_1519);
nand U3151 (N_3151,N_2374,N_942);
nand U3152 (N_3152,N_120,N_327);
and U3153 (N_3153,N_1777,N_1317);
nand U3154 (N_3154,N_2093,N_681);
and U3155 (N_3155,N_1818,N_1173);
nand U3156 (N_3156,N_1433,N_642);
and U3157 (N_3157,N_549,N_2365);
nand U3158 (N_3158,N_1414,N_1975);
nor U3159 (N_3159,N_163,N_527);
and U3160 (N_3160,N_1697,N_1642);
or U3161 (N_3161,N_776,N_2076);
nor U3162 (N_3162,N_1490,N_726);
or U3163 (N_3163,N_1865,N_26);
nor U3164 (N_3164,N_401,N_2364);
nor U3165 (N_3165,N_1481,N_43);
nor U3166 (N_3166,N_142,N_753);
and U3167 (N_3167,N_999,N_1846);
or U3168 (N_3168,N_1035,N_2294);
and U3169 (N_3169,N_1951,N_1140);
nand U3170 (N_3170,N_692,N_871);
or U3171 (N_3171,N_570,N_1509);
nand U3172 (N_3172,N_766,N_423);
nor U3173 (N_3173,N_1266,N_1243);
and U3174 (N_3174,N_2115,N_1905);
nand U3175 (N_3175,N_386,N_639);
xnor U3176 (N_3176,N_2103,N_2348);
and U3177 (N_3177,N_1701,N_2159);
xor U3178 (N_3178,N_1430,N_1124);
or U3179 (N_3179,N_1721,N_1730);
xor U3180 (N_3180,N_1110,N_1473);
and U3181 (N_3181,N_846,N_517);
nor U3182 (N_3182,N_1018,N_834);
nand U3183 (N_3183,N_2066,N_1242);
nor U3184 (N_3184,N_2492,N_1602);
nor U3185 (N_3185,N_289,N_728);
nor U3186 (N_3186,N_1377,N_2169);
nand U3187 (N_3187,N_851,N_1788);
or U3188 (N_3188,N_2017,N_1735);
nor U3189 (N_3189,N_2418,N_347);
and U3190 (N_3190,N_1799,N_85);
nor U3191 (N_3191,N_709,N_59);
and U3192 (N_3192,N_1121,N_402);
and U3193 (N_3193,N_1028,N_2009);
nand U3194 (N_3194,N_260,N_755);
or U3195 (N_3195,N_69,N_619);
nor U3196 (N_3196,N_633,N_490);
and U3197 (N_3197,N_1294,N_2256);
nand U3198 (N_3198,N_56,N_844);
and U3199 (N_3199,N_2371,N_1040);
nand U3200 (N_3200,N_2321,N_139);
xor U3201 (N_3201,N_594,N_798);
or U3202 (N_3202,N_1482,N_417);
and U3203 (N_3203,N_180,N_2483);
or U3204 (N_3204,N_720,N_1958);
nor U3205 (N_3205,N_1676,N_733);
nor U3206 (N_3206,N_130,N_1834);
and U3207 (N_3207,N_494,N_1466);
nand U3208 (N_3208,N_483,N_2139);
or U3209 (N_3209,N_1628,N_1322);
nand U3210 (N_3210,N_1650,N_66);
nor U3211 (N_3211,N_1288,N_1632);
nand U3212 (N_3212,N_1500,N_2011);
xnor U3213 (N_3213,N_1034,N_1805);
nand U3214 (N_3214,N_320,N_407);
and U3215 (N_3215,N_2270,N_1195);
or U3216 (N_3216,N_2308,N_1703);
or U3217 (N_3217,N_1536,N_2064);
xor U3218 (N_3218,N_1912,N_1186);
and U3219 (N_3219,N_501,N_1911);
or U3220 (N_3220,N_1373,N_113);
nand U3221 (N_3221,N_2003,N_1292);
xor U3222 (N_3222,N_1707,N_2036);
nand U3223 (N_3223,N_393,N_217);
and U3224 (N_3224,N_370,N_1038);
and U3225 (N_3225,N_1393,N_2421);
nand U3226 (N_3226,N_2474,N_973);
xor U3227 (N_3227,N_1684,N_1097);
and U3228 (N_3228,N_892,N_1365);
or U3229 (N_3229,N_1666,N_1950);
and U3230 (N_3230,N_1268,N_1158);
nand U3231 (N_3231,N_1142,N_1783);
nor U3232 (N_3232,N_833,N_1177);
nor U3233 (N_3233,N_2397,N_1781);
and U3234 (N_3234,N_889,N_2180);
or U3235 (N_3235,N_2242,N_2479);
or U3236 (N_3236,N_1614,N_2493);
nand U3237 (N_3237,N_2168,N_1791);
nand U3238 (N_3238,N_2432,N_2227);
nand U3239 (N_3239,N_1946,N_1250);
or U3240 (N_3240,N_2248,N_581);
nor U3241 (N_3241,N_1774,N_1814);
nand U3242 (N_3242,N_1530,N_1659);
and U3243 (N_3243,N_436,N_2465);
and U3244 (N_3244,N_1257,N_1460);
and U3245 (N_3245,N_662,N_106);
nand U3246 (N_3246,N_9,N_521);
and U3247 (N_3247,N_2384,N_2132);
or U3248 (N_3248,N_1058,N_976);
or U3249 (N_3249,N_2296,N_388);
nand U3250 (N_3250,N_806,N_1839);
or U3251 (N_3251,N_724,N_2341);
nor U3252 (N_3252,N_469,N_64);
or U3253 (N_3253,N_206,N_742);
nand U3254 (N_3254,N_836,N_281);
and U3255 (N_3255,N_2181,N_1852);
nor U3256 (N_3256,N_1005,N_1077);
and U3257 (N_3257,N_2404,N_1437);
xor U3258 (N_3258,N_673,N_1255);
xnor U3259 (N_3259,N_2297,N_1417);
or U3260 (N_3260,N_2496,N_1868);
xnor U3261 (N_3261,N_2067,N_1625);
or U3262 (N_3262,N_1143,N_1087);
and U3263 (N_3263,N_12,N_1445);
and U3264 (N_3264,N_8,N_1344);
nor U3265 (N_3265,N_1366,N_1724);
and U3266 (N_3266,N_360,N_628);
xnor U3267 (N_3267,N_1339,N_2422);
nand U3268 (N_3268,N_546,N_1323);
nor U3269 (N_3269,N_2317,N_1451);
nand U3270 (N_3270,N_1403,N_2054);
or U3271 (N_3271,N_488,N_2006);
nand U3272 (N_3272,N_1495,N_884);
nand U3273 (N_3273,N_343,N_1899);
and U3274 (N_3274,N_943,N_731);
xor U3275 (N_3275,N_2494,N_696);
or U3276 (N_3276,N_2488,N_710);
nand U3277 (N_3277,N_1297,N_1939);
xnor U3278 (N_3278,N_1178,N_1843);
xnor U3279 (N_3279,N_1168,N_1785);
or U3280 (N_3280,N_2343,N_1390);
and U3281 (N_3281,N_1400,N_2392);
or U3282 (N_3282,N_1126,N_2455);
and U3283 (N_3283,N_568,N_2268);
or U3284 (N_3284,N_1869,N_237);
nor U3285 (N_3285,N_2260,N_705);
or U3286 (N_3286,N_1745,N_1815);
nor U3287 (N_3287,N_302,N_2391);
nor U3288 (N_3288,N_1291,N_2330);
nor U3289 (N_3289,N_1827,N_2289);
nor U3290 (N_3290,N_1644,N_513);
nor U3291 (N_3291,N_968,N_765);
nor U3292 (N_3292,N_2110,N_318);
or U3293 (N_3293,N_2039,N_2104);
and U3294 (N_3294,N_449,N_2349);
nor U3295 (N_3295,N_336,N_1020);
nor U3296 (N_3296,N_675,N_861);
and U3297 (N_3297,N_814,N_1256);
xnor U3298 (N_3298,N_2347,N_1216);
and U3299 (N_3299,N_1402,N_24);
xnor U3300 (N_3300,N_329,N_261);
nor U3301 (N_3301,N_531,N_379);
nand U3302 (N_3302,N_1906,N_2151);
or U3303 (N_3303,N_845,N_1164);
xnor U3304 (N_3304,N_389,N_159);
nor U3305 (N_3305,N_1429,N_785);
and U3306 (N_3306,N_1469,N_1638);
or U3307 (N_3307,N_435,N_2065);
and U3308 (N_3308,N_1263,N_22);
nor U3309 (N_3309,N_342,N_676);
nand U3310 (N_3310,N_134,N_1514);
or U3311 (N_3311,N_1853,N_1733);
nor U3312 (N_3312,N_171,N_345);
or U3313 (N_3313,N_344,N_1570);
or U3314 (N_3314,N_1172,N_936);
nand U3315 (N_3315,N_458,N_1563);
nand U3316 (N_3316,N_1588,N_2429);
or U3317 (N_3317,N_2063,N_110);
nor U3318 (N_3318,N_272,N_1306);
nor U3319 (N_3319,N_1687,N_1501);
or U3320 (N_3320,N_1547,N_512);
xor U3321 (N_3321,N_1850,N_1611);
and U3322 (N_3322,N_932,N_2025);
xor U3323 (N_3323,N_805,N_1947);
nand U3324 (N_3324,N_1134,N_773);
nor U3325 (N_3325,N_1675,N_2099);
nor U3326 (N_3326,N_1061,N_1078);
and U3327 (N_3327,N_1714,N_1873);
and U3328 (N_3328,N_768,N_2212);
nor U3329 (N_3329,N_1032,N_1369);
or U3330 (N_3330,N_1264,N_80);
or U3331 (N_3331,N_2271,N_1826);
nand U3332 (N_3332,N_1953,N_701);
or U3333 (N_3333,N_310,N_1516);
nor U3334 (N_3334,N_16,N_885);
and U3335 (N_3335,N_1732,N_756);
or U3336 (N_3336,N_1187,N_1534);
or U3337 (N_3337,N_2426,N_2291);
nor U3338 (N_3338,N_879,N_608);
nand U3339 (N_3339,N_1162,N_2490);
nand U3340 (N_3340,N_195,N_2261);
xnor U3341 (N_3341,N_544,N_505);
nor U3342 (N_3342,N_1508,N_2167);
and U3343 (N_3343,N_1978,N_194);
xnor U3344 (N_3344,N_848,N_2471);
and U3345 (N_3345,N_202,N_2443);
nand U3346 (N_3346,N_1204,N_463);
and U3347 (N_3347,N_659,N_2195);
nand U3348 (N_3348,N_1952,N_1318);
nand U3349 (N_3349,N_299,N_2015);
or U3350 (N_3350,N_1252,N_2214);
nor U3351 (N_3351,N_2028,N_498);
and U3352 (N_3352,N_523,N_707);
nor U3353 (N_3353,N_1535,N_1304);
or U3354 (N_3354,N_2106,N_1248);
nor U3355 (N_3355,N_190,N_683);
nand U3356 (N_3356,N_518,N_992);
nor U3357 (N_3357,N_1130,N_907);
nand U3358 (N_3358,N_67,N_492);
or U3359 (N_3359,N_605,N_1064);
nand U3360 (N_3360,N_1165,N_616);
nor U3361 (N_3361,N_1303,N_1878);
nor U3362 (N_3362,N_1985,N_783);
and U3363 (N_3363,N_35,N_690);
or U3364 (N_3364,N_225,N_1768);
nor U3365 (N_3365,N_201,N_262);
and U3366 (N_3366,N_196,N_1047);
nand U3367 (N_3367,N_603,N_1133);
nand U3368 (N_3368,N_2240,N_532);
nand U3369 (N_3369,N_296,N_1990);
and U3370 (N_3370,N_137,N_44);
nand U3371 (N_3371,N_1104,N_1079);
and U3372 (N_3372,N_2453,N_2026);
xnor U3373 (N_3373,N_598,N_1180);
and U3374 (N_3374,N_2081,N_966);
and U3375 (N_3375,N_689,N_780);
xnor U3376 (N_3376,N_591,N_390);
nor U3377 (N_3377,N_1421,N_368);
nor U3378 (N_3378,N_1289,N_2142);
or U3379 (N_3379,N_1022,N_503);
nand U3380 (N_3380,N_1900,N_782);
nor U3381 (N_3381,N_485,N_1039);
xor U3382 (N_3382,N_2462,N_933);
and U3383 (N_3383,N_1897,N_2315);
nand U3384 (N_3384,N_470,N_1275);
xnor U3385 (N_3385,N_2223,N_151);
nand U3386 (N_3386,N_1898,N_2447);
or U3387 (N_3387,N_827,N_694);
nand U3388 (N_3388,N_353,N_1859);
or U3389 (N_3389,N_1974,N_663);
and U3390 (N_3390,N_74,N_1411);
nand U3391 (N_3391,N_475,N_1353);
xor U3392 (N_3392,N_2033,N_1706);
nand U3393 (N_3393,N_1664,N_2201);
nand U3394 (N_3394,N_1904,N_930);
or U3395 (N_3395,N_2107,N_637);
or U3396 (N_3396,N_2100,N_1357);
nand U3397 (N_3397,N_47,N_1170);
nand U3398 (N_3398,N_479,N_1924);
nor U3399 (N_3399,N_1605,N_2457);
and U3400 (N_3400,N_428,N_2247);
nand U3401 (N_3401,N_1282,N_769);
and U3402 (N_3402,N_1136,N_250);
nand U3403 (N_3403,N_635,N_2148);
xor U3404 (N_3404,N_1211,N_1832);
nand U3405 (N_3405,N_1540,N_816);
nand U3406 (N_3406,N_63,N_444);
nor U3407 (N_3407,N_989,N_2184);
or U3408 (N_3408,N_1670,N_1337);
or U3409 (N_3409,N_2353,N_2281);
nand U3410 (N_3410,N_489,N_623);
xor U3411 (N_3411,N_397,N_184);
or U3412 (N_3412,N_38,N_1485);
nand U3413 (N_3413,N_652,N_405);
nand U3414 (N_3414,N_682,N_1656);
nand U3415 (N_3415,N_102,N_1092);
and U3416 (N_3416,N_1689,N_974);
nand U3417 (N_3417,N_265,N_107);
nor U3418 (N_3418,N_2359,N_2238);
xnor U3419 (N_3419,N_762,N_2182);
and U3420 (N_3420,N_1049,N_1931);
nor U3421 (N_3421,N_1063,N_668);
nor U3422 (N_3422,N_2109,N_2440);
xor U3423 (N_3423,N_303,N_259);
nor U3424 (N_3424,N_148,N_338);
xnor U3425 (N_3425,N_826,N_294);
and U3426 (N_3426,N_415,N_563);
nor U3427 (N_3427,N_290,N_1389);
nand U3428 (N_3428,N_11,N_865);
and U3429 (N_3429,N_172,N_1067);
and U3430 (N_3430,N_1123,N_1330);
nor U3431 (N_3431,N_2008,N_54);
or U3432 (N_3432,N_547,N_1699);
xor U3433 (N_3433,N_2410,N_1181);
and U3434 (N_3434,N_32,N_597);
nor U3435 (N_3435,N_1736,N_459);
or U3436 (N_3436,N_993,N_2283);
or U3437 (N_3437,N_583,N_108);
xnor U3438 (N_3438,N_346,N_1174);
and U3439 (N_3439,N_98,N_141);
nor U3440 (N_3440,N_147,N_702);
and U3441 (N_3441,N_1137,N_2010);
and U3442 (N_3442,N_1660,N_1669);
nand U3443 (N_3443,N_2029,N_37);
or U3444 (N_3444,N_2424,N_1333);
nand U3445 (N_3445,N_1809,N_2403);
nor U3446 (N_3446,N_2174,N_1996);
xor U3447 (N_3447,N_1394,N_1315);
and U3448 (N_3448,N_49,N_153);
or U3449 (N_3449,N_1746,N_4);
or U3450 (N_3450,N_713,N_1543);
or U3451 (N_3451,N_670,N_1138);
nand U3452 (N_3452,N_2020,N_2377);
xnor U3453 (N_3453,N_1796,N_1607);
and U3454 (N_3454,N_1057,N_1620);
xnor U3455 (N_3455,N_2361,N_1860);
nand U3456 (N_3456,N_1205,N_712);
nand U3457 (N_3457,N_1581,N_685);
and U3458 (N_3458,N_1474,N_1583);
nand U3459 (N_3459,N_1235,N_1663);
xnor U3460 (N_3460,N_204,N_2111);
and U3461 (N_3461,N_797,N_117);
nand U3462 (N_3462,N_657,N_971);
xor U3463 (N_3463,N_57,N_1105);
nor U3464 (N_3464,N_761,N_442);
nor U3465 (N_3465,N_2072,N_2134);
or U3466 (N_3466,N_1016,N_651);
nor U3467 (N_3467,N_866,N_1185);
and U3468 (N_3468,N_257,N_2272);
nand U3469 (N_3469,N_924,N_1094);
nor U3470 (N_3470,N_42,N_468);
xnor U3471 (N_3471,N_2303,N_1861);
nor U3472 (N_3472,N_1523,N_1464);
nor U3473 (N_3473,N_1800,N_1704);
and U3474 (N_3474,N_484,N_868);
nor U3475 (N_3475,N_622,N_373);
xor U3476 (N_3476,N_1476,N_2387);
and U3477 (N_3477,N_2122,N_2123);
and U3478 (N_3478,N_300,N_1992);
nand U3479 (N_3479,N_1107,N_1761);
nand U3480 (N_3480,N_2221,N_734);
xor U3481 (N_3481,N_883,N_516);
nor U3482 (N_3482,N_276,N_1129);
or U3483 (N_3483,N_2278,N_1560);
or U3484 (N_3484,N_1036,N_1144);
nand U3485 (N_3485,N_1100,N_964);
nor U3486 (N_3486,N_2414,N_1218);
and U3487 (N_3487,N_1770,N_1506);
and U3488 (N_3488,N_39,N_1465);
or U3489 (N_3489,N_1648,N_429);
nand U3490 (N_3490,N_1810,N_1794);
or U3491 (N_3491,N_1452,N_648);
xor U3492 (N_3492,N_1512,N_2030);
or U3493 (N_3493,N_2075,N_881);
xor U3494 (N_3494,N_244,N_1629);
and U3495 (N_3495,N_1253,N_584);
and U3496 (N_3496,N_794,N_813);
and U3497 (N_3497,N_2334,N_1139);
and U3498 (N_3498,N_2276,N_1773);
and U3499 (N_3499,N_1520,N_1532);
nand U3500 (N_3500,N_537,N_1615);
xor U3501 (N_3501,N_422,N_2022);
nand U3502 (N_3502,N_502,N_772);
and U3503 (N_3503,N_740,N_913);
or U3504 (N_3504,N_736,N_698);
nor U3505 (N_3505,N_2027,N_779);
or U3506 (N_3506,N_1088,N_197);
or U3507 (N_3507,N_1857,N_431);
and U3508 (N_3508,N_1332,N_253);
and U3509 (N_3509,N_126,N_1541);
and U3510 (N_3510,N_333,N_1497);
nor U3511 (N_3511,N_1491,N_1002);
nand U3512 (N_3512,N_2370,N_621);
and U3513 (N_3513,N_1589,N_233);
nor U3514 (N_3514,N_1215,N_354);
nor U3515 (N_3515,N_83,N_495);
or U3516 (N_3516,N_2079,N_1521);
nor U3517 (N_3517,N_1108,N_819);
nor U3518 (N_3518,N_903,N_1551);
or U3519 (N_3519,N_146,N_1986);
nand U3520 (N_3520,N_2206,N_1397);
nand U3521 (N_3521,N_1713,N_81);
and U3522 (N_3522,N_164,N_1739);
nor U3523 (N_3523,N_5,N_975);
or U3524 (N_3524,N_2068,N_815);
and U3525 (N_3525,N_1012,N_119);
or U3526 (N_3526,N_2306,N_2386);
or U3527 (N_3527,N_743,N_447);
nand U3528 (N_3528,N_630,N_1420);
nand U3529 (N_3529,N_392,N_1858);
nand U3530 (N_3530,N_1529,N_15);
nand U3531 (N_3531,N_669,N_298);
nor U3532 (N_3532,N_2452,N_1716);
or U3533 (N_3533,N_1617,N_1639);
or U3534 (N_3534,N_672,N_1837);
nand U3535 (N_3535,N_7,N_1118);
and U3536 (N_3536,N_1499,N_1549);
or U3537 (N_3537,N_2360,N_378);
xor U3538 (N_3538,N_2136,N_1043);
and U3539 (N_3539,N_1000,N_2434);
and U3540 (N_3540,N_2298,N_2277);
and U3541 (N_3541,N_615,N_2331);
and U3542 (N_3542,N_1624,N_1447);
nand U3543 (N_3543,N_601,N_247);
nor U3544 (N_3544,N_687,N_1434);
nand U3545 (N_3545,N_1979,N_121);
xnor U3546 (N_3546,N_2048,N_1808);
nor U3547 (N_3547,N_524,N_279);
xor U3548 (N_3548,N_1538,N_116);
and U3549 (N_3549,N_777,N_641);
xnor U3550 (N_3550,N_1576,N_288);
and U3551 (N_3551,N_2233,N_2205);
nor U3552 (N_3552,N_1479,N_340);
and U3553 (N_3553,N_291,N_823);
and U3554 (N_3554,N_2021,N_1362);
nor U3555 (N_3555,N_2173,N_2178);
nor U3556 (N_3556,N_2484,N_721);
nor U3557 (N_3557,N_2445,N_1962);
xnor U3558 (N_3558,N_228,N_437);
or U3559 (N_3559,N_954,N_1921);
xor U3560 (N_3560,N_451,N_1103);
or U3561 (N_3561,N_1608,N_278);
and U3562 (N_3562,N_1345,N_60);
and U3563 (N_3563,N_1001,N_1080);
nand U3564 (N_3564,N_95,N_876);
or U3565 (N_3565,N_2078,N_645);
xor U3566 (N_3566,N_2352,N_1959);
and U3567 (N_3567,N_174,N_277);
nor U3568 (N_3568,N_1091,N_1896);
and U3569 (N_3569,N_1385,N_292);
nor U3570 (N_3570,N_1686,N_1010);
xor U3571 (N_3571,N_923,N_1309);
or U3572 (N_3572,N_2345,N_445);
and U3573 (N_3573,N_997,N_220);
nor U3574 (N_3574,N_1492,N_2226);
nand U3575 (N_3575,N_2293,N_732);
nor U3576 (N_3576,N_454,N_526);
nor U3577 (N_3577,N_910,N_609);
and U3578 (N_3578,N_849,N_1927);
xnor U3579 (N_3579,N_1349,N_2325);
nor U3580 (N_3580,N_1633,N_2170);
nor U3581 (N_3581,N_366,N_825);
and U3582 (N_3582,N_1970,N_214);
nand U3583 (N_3583,N_811,N_500);
and U3584 (N_3584,N_1919,N_1153);
nor U3585 (N_3585,N_1743,N_571);
and U3586 (N_3586,N_1957,N_719);
or U3587 (N_3587,N_461,N_1206);
and U3588 (N_3588,N_2473,N_1406);
nand U3589 (N_3589,N_287,N_50);
nand U3590 (N_3590,N_2002,N_1449);
nand U3591 (N_3591,N_157,N_438);
and U3592 (N_3592,N_2097,N_1388);
nand U3593 (N_3593,N_19,N_2085);
nor U3594 (N_3594,N_341,N_385);
or U3595 (N_3595,N_2269,N_862);
nor U3596 (N_3596,N_1798,N_2162);
or U3597 (N_3597,N_2301,N_781);
and U3598 (N_3598,N_1234,N_280);
nand U3599 (N_3599,N_1046,N_439);
or U3600 (N_3600,N_2086,N_656);
nand U3601 (N_3601,N_2249,N_564);
nor U3602 (N_3602,N_1555,N_1674);
and U3603 (N_3603,N_775,N_1943);
xnor U3604 (N_3604,N_2070,N_1227);
and U3605 (N_3605,N_1587,N_1510);
and U3606 (N_3606,N_314,N_2062);
nand U3607 (N_3607,N_499,N_771);
and U3608 (N_3608,N_2018,N_2398);
and U3609 (N_3609,N_170,N_856);
and U3610 (N_3610,N_634,N_1886);
and U3611 (N_3611,N_1719,N_1740);
nand U3612 (N_3612,N_455,N_1609);
and U3613 (N_3613,N_2197,N_1678);
xor U3614 (N_3614,N_480,N_337);
nand U3615 (N_3615,N_588,N_2243);
nand U3616 (N_3616,N_926,N_693);
or U3617 (N_3617,N_1829,N_880);
and U3618 (N_3618,N_751,N_349);
nor U3619 (N_3619,N_977,N_129);
or U3620 (N_3620,N_2402,N_138);
and U3621 (N_3621,N_1157,N_2366);
nor U3622 (N_3622,N_179,N_758);
or U3623 (N_3623,N_841,N_2231);
nand U3624 (N_3624,N_2204,N_2092);
or U3625 (N_3625,N_161,N_2263);
and U3626 (N_3626,N_1573,N_1281);
nor U3627 (N_3627,N_511,N_285);
or U3628 (N_3628,N_1175,N_1192);
or U3629 (N_3629,N_156,N_1749);
and U3630 (N_3630,N_2019,N_2363);
nand U3631 (N_3631,N_767,N_1963);
or U3632 (N_3632,N_1111,N_1895);
nand U3633 (N_3633,N_398,N_606);
xnor U3634 (N_3634,N_1410,N_266);
nor U3635 (N_3635,N_358,N_2285);
and U3636 (N_3636,N_1223,N_2290);
nand U3637 (N_3637,N_1544,N_481);
or U3638 (N_3638,N_644,N_491);
nor U3639 (N_3639,N_981,N_1526);
or U3640 (N_3640,N_375,N_1381);
nand U3641 (N_3641,N_36,N_557);
or U3642 (N_3642,N_1937,N_2000);
nand U3643 (N_3643,N_820,N_1435);
or U3644 (N_3644,N_1847,N_2381);
or U3645 (N_3645,N_1209,N_589);
or U3646 (N_3646,N_1752,N_2130);
xor U3647 (N_3647,N_655,N_2090);
or U3648 (N_3648,N_114,N_1621);
nor U3649 (N_3649,N_241,N_1329);
xor U3650 (N_3650,N_1564,N_1191);
nor U3651 (N_3651,N_745,N_1127);
nand U3652 (N_3652,N_1048,N_496);
nor U3653 (N_3653,N_1848,N_2166);
and U3654 (N_3654,N_409,N_1051);
nor U3655 (N_3655,N_1461,N_1901);
nor U3656 (N_3656,N_760,N_1283);
nand U3657 (N_3657,N_1545,N_955);
nand U3658 (N_3658,N_1657,N_509);
nor U3659 (N_3659,N_1194,N_2497);
and U3660 (N_3660,N_160,N_2143);
nand U3661 (N_3661,N_1361,N_2305);
nor U3662 (N_3662,N_269,N_2172);
nand U3663 (N_3663,N_293,N_1665);
nand U3664 (N_3664,N_1976,N_1441);
or U3665 (N_3665,N_625,N_53);
nand U3666 (N_3666,N_1171,N_1238);
nand U3667 (N_3667,N_1750,N_198);
or U3668 (N_3668,N_448,N_18);
nand U3669 (N_3669,N_1760,N_486);
or U3670 (N_3670,N_1751,N_1169);
or U3671 (N_3671,N_235,N_122);
nor U3672 (N_3672,N_2313,N_1325);
nand U3673 (N_3673,N_1824,N_1462);
or U3674 (N_3674,N_1352,N_908);
xor U3675 (N_3675,N_1513,N_2416);
nand U3676 (N_3676,N_951,N_835);
nand U3677 (N_3677,N_230,N_801);
or U3678 (N_3678,N_2383,N_790);
or U3679 (N_3679,N_186,N_1471);
nand U3680 (N_3680,N_554,N_2186);
nand U3681 (N_3681,N_452,N_578);
nand U3682 (N_3682,N_893,N_545);
or U3683 (N_3683,N_1754,N_103);
or U3684 (N_3684,N_1806,N_2224);
or U3685 (N_3685,N_1062,N_328);
nor U3686 (N_3686,N_1183,N_207);
xor U3687 (N_3687,N_1934,N_1358);
and U3688 (N_3688,N_77,N_1915);
or U3689 (N_3689,N_1415,N_0);
xor U3690 (N_3690,N_1844,N_2061);
and U3691 (N_3691,N_1616,N_1935);
and U3692 (N_3692,N_1054,N_443);
nand U3693 (N_3693,N_793,N_2394);
and U3694 (N_3694,N_403,N_432);
nand U3695 (N_3695,N_1472,N_149);
xor U3696 (N_3696,N_1662,N_985);
or U3697 (N_3697,N_1095,N_561);
nor U3698 (N_3698,N_1910,N_2423);
nor U3699 (N_3699,N_2150,N_2149);
and U3700 (N_3700,N_1249,N_812);
or U3701 (N_3701,N_764,N_949);
or U3702 (N_3702,N_2327,N_359);
nand U3703 (N_3703,N_212,N_1093);
or U3704 (N_3704,N_2388,N_730);
nand U3705 (N_3705,N_2058,N_1418);
nand U3706 (N_3706,N_1710,N_1916);
or U3707 (N_3707,N_650,N_1190);
nand U3708 (N_3708,N_1866,N_787);
or U3709 (N_3709,N_2218,N_1300);
nand U3710 (N_3710,N_520,N_30);
nor U3711 (N_3711,N_1920,N_1109);
nand U3712 (N_3712,N_1208,N_377);
and U3713 (N_3713,N_748,N_1273);
nand U3714 (N_3714,N_553,N_1504);
nor U3715 (N_3715,N_1584,N_2158);
nand U3716 (N_3716,N_2335,N_984);
or U3717 (N_3717,N_1888,N_796);
nand U3718 (N_3718,N_1623,N_2089);
xor U3719 (N_3719,N_1070,N_1667);
xor U3720 (N_3720,N_282,N_1559);
nor U3721 (N_3721,N_2486,N_859);
nor U3722 (N_3722,N_78,N_1651);
nand U3723 (N_3723,N_1463,N_440);
xnor U3724 (N_3724,N_73,N_2259);
nor U3725 (N_3725,N_1889,N_263);
nor U3726 (N_3726,N_1324,N_1198);
and U3727 (N_3727,N_1683,N_569);
nand U3728 (N_3728,N_1725,N_2286);
or U3729 (N_3729,N_1871,N_667);
nor U3730 (N_3730,N_90,N_1784);
and U3731 (N_3731,N_144,N_595);
xor U3732 (N_3732,N_1856,N_1453);
and U3733 (N_3733,N_1870,N_931);
xor U3734 (N_3734,N_1556,N_2244);
nand U3735 (N_3735,N_1159,N_408);
and U3736 (N_3736,N_1580,N_2050);
nor U3737 (N_3737,N_875,N_362);
nand U3738 (N_3738,N_2145,N_1830);
or U3739 (N_3739,N_1596,N_1348);
and U3740 (N_3740,N_1731,N_1030);
xnor U3741 (N_3741,N_2385,N_70);
or U3742 (N_3742,N_1146,N_1863);
nand U3743 (N_3743,N_1239,N_1438);
or U3744 (N_3744,N_565,N_2323);
or U3745 (N_3745,N_248,N_132);
or U3746 (N_3746,N_807,N_538);
nor U3747 (N_3747,N_2056,N_638);
or U3748 (N_3748,N_886,N_1575);
nand U3749 (N_3749,N_472,N_525);
nor U3750 (N_3750,N_308,N_1038);
nor U3751 (N_3751,N_306,N_509);
xor U3752 (N_3752,N_632,N_1250);
nor U3753 (N_3753,N_2327,N_200);
and U3754 (N_3754,N_2381,N_1313);
or U3755 (N_3755,N_2128,N_694);
nor U3756 (N_3756,N_1617,N_439);
nand U3757 (N_3757,N_703,N_2180);
nor U3758 (N_3758,N_1545,N_643);
or U3759 (N_3759,N_1678,N_2439);
or U3760 (N_3760,N_2129,N_612);
nor U3761 (N_3761,N_621,N_2141);
nor U3762 (N_3762,N_2139,N_2356);
xnor U3763 (N_3763,N_1169,N_1042);
xor U3764 (N_3764,N_1823,N_946);
nor U3765 (N_3765,N_31,N_776);
nand U3766 (N_3766,N_1507,N_3);
and U3767 (N_3767,N_788,N_1600);
nor U3768 (N_3768,N_2075,N_1098);
or U3769 (N_3769,N_1747,N_1555);
and U3770 (N_3770,N_1585,N_446);
nand U3771 (N_3771,N_666,N_2283);
or U3772 (N_3772,N_1979,N_1070);
and U3773 (N_3773,N_925,N_2064);
or U3774 (N_3774,N_618,N_732);
nor U3775 (N_3775,N_2331,N_1361);
nor U3776 (N_3776,N_2126,N_477);
nand U3777 (N_3777,N_1444,N_2067);
nor U3778 (N_3778,N_699,N_393);
and U3779 (N_3779,N_205,N_1899);
nand U3780 (N_3780,N_1350,N_1039);
or U3781 (N_3781,N_1499,N_1190);
and U3782 (N_3782,N_1591,N_297);
nor U3783 (N_3783,N_1500,N_216);
nand U3784 (N_3784,N_1382,N_8);
nor U3785 (N_3785,N_875,N_51);
and U3786 (N_3786,N_1337,N_649);
nand U3787 (N_3787,N_1274,N_2269);
or U3788 (N_3788,N_55,N_1025);
or U3789 (N_3789,N_1763,N_2497);
nand U3790 (N_3790,N_1019,N_1222);
or U3791 (N_3791,N_2040,N_646);
nor U3792 (N_3792,N_275,N_1637);
or U3793 (N_3793,N_338,N_2080);
nor U3794 (N_3794,N_911,N_506);
nand U3795 (N_3795,N_2133,N_2011);
or U3796 (N_3796,N_241,N_2077);
nor U3797 (N_3797,N_878,N_227);
and U3798 (N_3798,N_407,N_787);
and U3799 (N_3799,N_117,N_596);
and U3800 (N_3800,N_322,N_2311);
nor U3801 (N_3801,N_93,N_70);
and U3802 (N_3802,N_2390,N_1351);
nor U3803 (N_3803,N_18,N_1103);
xnor U3804 (N_3804,N_2376,N_129);
nand U3805 (N_3805,N_135,N_1286);
or U3806 (N_3806,N_200,N_268);
nor U3807 (N_3807,N_553,N_705);
xor U3808 (N_3808,N_2103,N_1982);
nor U3809 (N_3809,N_1255,N_1700);
nor U3810 (N_3810,N_1497,N_313);
and U3811 (N_3811,N_1729,N_326);
and U3812 (N_3812,N_2454,N_521);
nand U3813 (N_3813,N_2434,N_181);
nor U3814 (N_3814,N_1480,N_2037);
or U3815 (N_3815,N_2056,N_1337);
xnor U3816 (N_3816,N_372,N_709);
nor U3817 (N_3817,N_1063,N_2097);
and U3818 (N_3818,N_2021,N_1030);
nand U3819 (N_3819,N_958,N_1925);
nor U3820 (N_3820,N_2491,N_1345);
or U3821 (N_3821,N_1588,N_965);
xor U3822 (N_3822,N_882,N_233);
nor U3823 (N_3823,N_122,N_311);
nor U3824 (N_3824,N_1818,N_236);
nor U3825 (N_3825,N_782,N_1794);
nand U3826 (N_3826,N_178,N_744);
nor U3827 (N_3827,N_877,N_939);
nor U3828 (N_3828,N_1840,N_579);
nand U3829 (N_3829,N_1296,N_605);
nand U3830 (N_3830,N_318,N_2262);
and U3831 (N_3831,N_1545,N_470);
and U3832 (N_3832,N_529,N_304);
and U3833 (N_3833,N_1756,N_1231);
or U3834 (N_3834,N_1221,N_1249);
nand U3835 (N_3835,N_87,N_938);
nor U3836 (N_3836,N_1755,N_1868);
and U3837 (N_3837,N_1511,N_1477);
and U3838 (N_3838,N_2301,N_1784);
or U3839 (N_3839,N_763,N_45);
and U3840 (N_3840,N_1823,N_2134);
and U3841 (N_3841,N_1717,N_2322);
xor U3842 (N_3842,N_1368,N_1261);
nand U3843 (N_3843,N_840,N_2409);
nand U3844 (N_3844,N_34,N_523);
or U3845 (N_3845,N_58,N_371);
or U3846 (N_3846,N_776,N_1566);
nand U3847 (N_3847,N_2332,N_1169);
nand U3848 (N_3848,N_1957,N_77);
nand U3849 (N_3849,N_975,N_774);
nand U3850 (N_3850,N_334,N_1048);
or U3851 (N_3851,N_1684,N_98);
or U3852 (N_3852,N_985,N_2423);
and U3853 (N_3853,N_1176,N_1463);
and U3854 (N_3854,N_218,N_1741);
nor U3855 (N_3855,N_2469,N_1847);
or U3856 (N_3856,N_1520,N_266);
or U3857 (N_3857,N_684,N_542);
xnor U3858 (N_3858,N_1040,N_2245);
nand U3859 (N_3859,N_2063,N_1344);
or U3860 (N_3860,N_215,N_2468);
nand U3861 (N_3861,N_1838,N_1724);
and U3862 (N_3862,N_108,N_449);
xnor U3863 (N_3863,N_2276,N_1222);
nand U3864 (N_3864,N_834,N_2224);
or U3865 (N_3865,N_593,N_2303);
nand U3866 (N_3866,N_1310,N_294);
or U3867 (N_3867,N_1494,N_1391);
or U3868 (N_3868,N_1173,N_2206);
nand U3869 (N_3869,N_1366,N_40);
and U3870 (N_3870,N_669,N_26);
and U3871 (N_3871,N_2333,N_260);
nor U3872 (N_3872,N_377,N_1247);
or U3873 (N_3873,N_2045,N_854);
and U3874 (N_3874,N_797,N_2301);
and U3875 (N_3875,N_687,N_2426);
nand U3876 (N_3876,N_56,N_1736);
nand U3877 (N_3877,N_2372,N_1142);
nand U3878 (N_3878,N_385,N_687);
nand U3879 (N_3879,N_697,N_265);
or U3880 (N_3880,N_2465,N_966);
nand U3881 (N_3881,N_926,N_545);
nand U3882 (N_3882,N_566,N_125);
nor U3883 (N_3883,N_2330,N_618);
and U3884 (N_3884,N_980,N_272);
nor U3885 (N_3885,N_1158,N_882);
xnor U3886 (N_3886,N_675,N_1190);
xnor U3887 (N_3887,N_698,N_1638);
and U3888 (N_3888,N_943,N_176);
and U3889 (N_3889,N_1855,N_114);
nand U3890 (N_3890,N_1772,N_950);
or U3891 (N_3891,N_2409,N_951);
and U3892 (N_3892,N_2308,N_427);
nor U3893 (N_3893,N_2343,N_1986);
xor U3894 (N_3894,N_1351,N_1370);
nand U3895 (N_3895,N_2176,N_2167);
or U3896 (N_3896,N_426,N_109);
or U3897 (N_3897,N_336,N_2105);
nor U3898 (N_3898,N_1561,N_392);
nand U3899 (N_3899,N_20,N_2147);
nand U3900 (N_3900,N_40,N_1483);
and U3901 (N_3901,N_1429,N_1295);
nand U3902 (N_3902,N_2352,N_1150);
nor U3903 (N_3903,N_1953,N_1584);
nand U3904 (N_3904,N_1310,N_1278);
and U3905 (N_3905,N_154,N_594);
xor U3906 (N_3906,N_581,N_2047);
or U3907 (N_3907,N_2349,N_574);
or U3908 (N_3908,N_2060,N_344);
xor U3909 (N_3909,N_2275,N_1623);
nor U3910 (N_3910,N_1840,N_1680);
or U3911 (N_3911,N_185,N_1801);
nand U3912 (N_3912,N_1557,N_876);
or U3913 (N_3913,N_1695,N_1399);
nand U3914 (N_3914,N_247,N_490);
nand U3915 (N_3915,N_1843,N_589);
or U3916 (N_3916,N_1792,N_416);
nor U3917 (N_3917,N_958,N_740);
nor U3918 (N_3918,N_2436,N_833);
and U3919 (N_3919,N_99,N_626);
or U3920 (N_3920,N_564,N_1687);
nor U3921 (N_3921,N_408,N_1807);
or U3922 (N_3922,N_2450,N_455);
and U3923 (N_3923,N_1109,N_243);
nor U3924 (N_3924,N_1230,N_1557);
or U3925 (N_3925,N_777,N_2114);
and U3926 (N_3926,N_554,N_1746);
and U3927 (N_3927,N_2019,N_1969);
xnor U3928 (N_3928,N_1204,N_394);
nor U3929 (N_3929,N_1448,N_1939);
and U3930 (N_3930,N_1594,N_124);
or U3931 (N_3931,N_1661,N_1723);
nand U3932 (N_3932,N_1504,N_2173);
and U3933 (N_3933,N_2366,N_1775);
and U3934 (N_3934,N_1243,N_489);
nor U3935 (N_3935,N_2230,N_392);
nand U3936 (N_3936,N_2138,N_1027);
and U3937 (N_3937,N_119,N_1382);
nor U3938 (N_3938,N_1398,N_2308);
and U3939 (N_3939,N_2450,N_766);
nand U3940 (N_3940,N_1855,N_387);
or U3941 (N_3941,N_1789,N_2423);
nor U3942 (N_3942,N_2126,N_930);
or U3943 (N_3943,N_73,N_1731);
or U3944 (N_3944,N_524,N_363);
nand U3945 (N_3945,N_905,N_234);
nor U3946 (N_3946,N_1004,N_2474);
and U3947 (N_3947,N_983,N_622);
xor U3948 (N_3948,N_1706,N_2475);
or U3949 (N_3949,N_1183,N_832);
nand U3950 (N_3950,N_442,N_675);
nand U3951 (N_3951,N_639,N_2033);
xor U3952 (N_3952,N_142,N_699);
nand U3953 (N_3953,N_1893,N_1990);
or U3954 (N_3954,N_1872,N_753);
nand U3955 (N_3955,N_1487,N_1752);
nor U3956 (N_3956,N_829,N_2243);
and U3957 (N_3957,N_64,N_2442);
nand U3958 (N_3958,N_551,N_855);
and U3959 (N_3959,N_1909,N_1459);
xnor U3960 (N_3960,N_797,N_1443);
and U3961 (N_3961,N_1021,N_1856);
and U3962 (N_3962,N_31,N_2371);
and U3963 (N_3963,N_1460,N_1284);
or U3964 (N_3964,N_2408,N_1550);
or U3965 (N_3965,N_2130,N_301);
or U3966 (N_3966,N_1343,N_1801);
nor U3967 (N_3967,N_1734,N_1970);
or U3968 (N_3968,N_1021,N_1855);
nand U3969 (N_3969,N_539,N_1485);
and U3970 (N_3970,N_594,N_1415);
nand U3971 (N_3971,N_859,N_901);
nand U3972 (N_3972,N_2040,N_715);
nor U3973 (N_3973,N_1712,N_2294);
or U3974 (N_3974,N_2112,N_1529);
nor U3975 (N_3975,N_1758,N_896);
nor U3976 (N_3976,N_490,N_854);
xor U3977 (N_3977,N_1496,N_610);
or U3978 (N_3978,N_494,N_125);
nand U3979 (N_3979,N_1367,N_1986);
or U3980 (N_3980,N_270,N_27);
and U3981 (N_3981,N_352,N_2268);
or U3982 (N_3982,N_911,N_1878);
nor U3983 (N_3983,N_1458,N_418);
nor U3984 (N_3984,N_352,N_2434);
nand U3985 (N_3985,N_2386,N_2475);
nand U3986 (N_3986,N_603,N_2385);
xor U3987 (N_3987,N_2021,N_2120);
nand U3988 (N_3988,N_1258,N_46);
nor U3989 (N_3989,N_2019,N_968);
xnor U3990 (N_3990,N_650,N_343);
nor U3991 (N_3991,N_1220,N_1837);
nand U3992 (N_3992,N_2004,N_1392);
xor U3993 (N_3993,N_1165,N_1667);
nor U3994 (N_3994,N_214,N_6);
and U3995 (N_3995,N_1813,N_47);
nand U3996 (N_3996,N_954,N_1625);
or U3997 (N_3997,N_1709,N_385);
and U3998 (N_3998,N_103,N_1521);
and U3999 (N_3999,N_1182,N_1124);
nor U4000 (N_4000,N_1402,N_2194);
nor U4001 (N_4001,N_1594,N_2256);
nor U4002 (N_4002,N_2485,N_912);
xnor U4003 (N_4003,N_672,N_1434);
and U4004 (N_4004,N_1666,N_1624);
and U4005 (N_4005,N_420,N_676);
or U4006 (N_4006,N_128,N_1526);
nand U4007 (N_4007,N_1710,N_1237);
and U4008 (N_4008,N_1557,N_1572);
or U4009 (N_4009,N_707,N_335);
and U4010 (N_4010,N_755,N_1703);
nor U4011 (N_4011,N_2019,N_2340);
nand U4012 (N_4012,N_1160,N_2314);
nor U4013 (N_4013,N_310,N_1662);
nand U4014 (N_4014,N_347,N_2290);
nand U4015 (N_4015,N_1012,N_1960);
nand U4016 (N_4016,N_1324,N_1537);
or U4017 (N_4017,N_1800,N_94);
or U4018 (N_4018,N_1252,N_61);
nand U4019 (N_4019,N_1009,N_1267);
or U4020 (N_4020,N_2373,N_1315);
nand U4021 (N_4021,N_66,N_2441);
nor U4022 (N_4022,N_1865,N_2256);
nand U4023 (N_4023,N_2247,N_1211);
nor U4024 (N_4024,N_2414,N_29);
or U4025 (N_4025,N_1872,N_1987);
or U4026 (N_4026,N_927,N_677);
xnor U4027 (N_4027,N_2429,N_914);
and U4028 (N_4028,N_546,N_987);
xnor U4029 (N_4029,N_2312,N_1765);
nor U4030 (N_4030,N_2317,N_128);
xor U4031 (N_4031,N_114,N_361);
and U4032 (N_4032,N_240,N_2268);
nor U4033 (N_4033,N_1285,N_2496);
and U4034 (N_4034,N_79,N_1301);
and U4035 (N_4035,N_1485,N_154);
nand U4036 (N_4036,N_569,N_2435);
and U4037 (N_4037,N_814,N_2350);
and U4038 (N_4038,N_1853,N_1466);
nand U4039 (N_4039,N_1426,N_522);
and U4040 (N_4040,N_2183,N_2070);
and U4041 (N_4041,N_2320,N_1263);
nor U4042 (N_4042,N_1384,N_1704);
xor U4043 (N_4043,N_1388,N_1457);
xnor U4044 (N_4044,N_2294,N_954);
nand U4045 (N_4045,N_1150,N_1249);
nand U4046 (N_4046,N_1405,N_2216);
and U4047 (N_4047,N_1841,N_2218);
nand U4048 (N_4048,N_2115,N_1166);
and U4049 (N_4049,N_561,N_1001);
and U4050 (N_4050,N_392,N_2044);
or U4051 (N_4051,N_1442,N_1538);
or U4052 (N_4052,N_2245,N_551);
nor U4053 (N_4053,N_346,N_577);
and U4054 (N_4054,N_2471,N_2241);
and U4055 (N_4055,N_543,N_2172);
or U4056 (N_4056,N_640,N_1293);
nor U4057 (N_4057,N_1878,N_769);
or U4058 (N_4058,N_1824,N_2136);
nand U4059 (N_4059,N_180,N_1589);
nor U4060 (N_4060,N_2041,N_459);
nor U4061 (N_4061,N_78,N_1570);
or U4062 (N_4062,N_2318,N_1043);
or U4063 (N_4063,N_644,N_1119);
nor U4064 (N_4064,N_670,N_960);
xor U4065 (N_4065,N_1565,N_1493);
nor U4066 (N_4066,N_1976,N_1421);
xnor U4067 (N_4067,N_1887,N_2234);
nor U4068 (N_4068,N_995,N_1698);
or U4069 (N_4069,N_601,N_156);
or U4070 (N_4070,N_633,N_1265);
and U4071 (N_4071,N_941,N_971);
or U4072 (N_4072,N_96,N_1030);
and U4073 (N_4073,N_2311,N_130);
nand U4074 (N_4074,N_494,N_1443);
and U4075 (N_4075,N_1889,N_1985);
xor U4076 (N_4076,N_1186,N_2178);
nor U4077 (N_4077,N_704,N_2394);
or U4078 (N_4078,N_603,N_1101);
and U4079 (N_4079,N_2068,N_1523);
nor U4080 (N_4080,N_1991,N_585);
or U4081 (N_4081,N_396,N_2074);
nand U4082 (N_4082,N_2300,N_929);
or U4083 (N_4083,N_1236,N_1588);
nand U4084 (N_4084,N_2210,N_399);
xnor U4085 (N_4085,N_1216,N_108);
nand U4086 (N_4086,N_458,N_198);
nor U4087 (N_4087,N_266,N_1982);
and U4088 (N_4088,N_551,N_615);
and U4089 (N_4089,N_39,N_668);
nand U4090 (N_4090,N_1739,N_228);
nand U4091 (N_4091,N_1814,N_1012);
xor U4092 (N_4092,N_2,N_2083);
nand U4093 (N_4093,N_418,N_1510);
nor U4094 (N_4094,N_1951,N_2008);
nor U4095 (N_4095,N_1836,N_598);
nor U4096 (N_4096,N_1929,N_1397);
nor U4097 (N_4097,N_2216,N_300);
xor U4098 (N_4098,N_170,N_2483);
and U4099 (N_4099,N_1172,N_1676);
and U4100 (N_4100,N_1385,N_2134);
or U4101 (N_4101,N_126,N_1960);
nand U4102 (N_4102,N_1349,N_2370);
and U4103 (N_4103,N_1415,N_1144);
or U4104 (N_4104,N_285,N_724);
nor U4105 (N_4105,N_939,N_425);
xor U4106 (N_4106,N_2042,N_2494);
nand U4107 (N_4107,N_749,N_1902);
or U4108 (N_4108,N_1142,N_1531);
nor U4109 (N_4109,N_1030,N_1294);
or U4110 (N_4110,N_1602,N_2313);
xnor U4111 (N_4111,N_447,N_599);
or U4112 (N_4112,N_1964,N_1250);
and U4113 (N_4113,N_426,N_243);
xor U4114 (N_4114,N_269,N_270);
nand U4115 (N_4115,N_955,N_230);
or U4116 (N_4116,N_1584,N_679);
and U4117 (N_4117,N_1672,N_1471);
or U4118 (N_4118,N_437,N_2236);
or U4119 (N_4119,N_1067,N_1454);
or U4120 (N_4120,N_2174,N_1071);
and U4121 (N_4121,N_2493,N_1095);
and U4122 (N_4122,N_1615,N_2015);
nand U4123 (N_4123,N_2328,N_919);
nand U4124 (N_4124,N_1762,N_1892);
nor U4125 (N_4125,N_2270,N_962);
nand U4126 (N_4126,N_552,N_2116);
and U4127 (N_4127,N_1567,N_1835);
nor U4128 (N_4128,N_527,N_1503);
nand U4129 (N_4129,N_2145,N_1560);
nor U4130 (N_4130,N_2425,N_1479);
nand U4131 (N_4131,N_2335,N_1622);
and U4132 (N_4132,N_1593,N_1844);
and U4133 (N_4133,N_2105,N_2089);
xor U4134 (N_4134,N_1830,N_1687);
nor U4135 (N_4135,N_2121,N_1817);
or U4136 (N_4136,N_2103,N_1921);
nand U4137 (N_4137,N_622,N_2385);
nor U4138 (N_4138,N_1771,N_184);
and U4139 (N_4139,N_2455,N_923);
and U4140 (N_4140,N_2002,N_2377);
nor U4141 (N_4141,N_144,N_1897);
and U4142 (N_4142,N_606,N_2000);
nand U4143 (N_4143,N_562,N_1213);
or U4144 (N_4144,N_324,N_1528);
and U4145 (N_4145,N_1134,N_2458);
and U4146 (N_4146,N_1746,N_1152);
nand U4147 (N_4147,N_2341,N_2242);
xnor U4148 (N_4148,N_1569,N_1439);
nor U4149 (N_4149,N_1029,N_2134);
nor U4150 (N_4150,N_1365,N_2316);
nand U4151 (N_4151,N_1357,N_448);
nor U4152 (N_4152,N_320,N_1834);
or U4153 (N_4153,N_1394,N_2264);
nor U4154 (N_4154,N_2450,N_414);
and U4155 (N_4155,N_828,N_570);
nand U4156 (N_4156,N_1386,N_858);
or U4157 (N_4157,N_308,N_80);
nor U4158 (N_4158,N_2189,N_573);
nand U4159 (N_4159,N_1395,N_2080);
nand U4160 (N_4160,N_250,N_2452);
or U4161 (N_4161,N_835,N_1358);
nor U4162 (N_4162,N_278,N_894);
nand U4163 (N_4163,N_1053,N_60);
nor U4164 (N_4164,N_1604,N_1571);
or U4165 (N_4165,N_69,N_2051);
nand U4166 (N_4166,N_1905,N_762);
and U4167 (N_4167,N_1583,N_1611);
and U4168 (N_4168,N_393,N_833);
or U4169 (N_4169,N_1006,N_216);
or U4170 (N_4170,N_185,N_1692);
nand U4171 (N_4171,N_1477,N_399);
nand U4172 (N_4172,N_826,N_1918);
nor U4173 (N_4173,N_169,N_180);
xor U4174 (N_4174,N_2497,N_935);
or U4175 (N_4175,N_1485,N_391);
nand U4176 (N_4176,N_2289,N_1999);
nand U4177 (N_4177,N_231,N_330);
and U4178 (N_4178,N_1241,N_846);
and U4179 (N_4179,N_1919,N_1989);
or U4180 (N_4180,N_672,N_1233);
and U4181 (N_4181,N_865,N_267);
nand U4182 (N_4182,N_424,N_209);
and U4183 (N_4183,N_296,N_839);
and U4184 (N_4184,N_1538,N_1385);
or U4185 (N_4185,N_2207,N_1807);
nor U4186 (N_4186,N_351,N_1975);
nand U4187 (N_4187,N_2457,N_2077);
nor U4188 (N_4188,N_2241,N_2179);
or U4189 (N_4189,N_291,N_1108);
nor U4190 (N_4190,N_2297,N_1670);
or U4191 (N_4191,N_2443,N_1204);
nor U4192 (N_4192,N_1767,N_771);
nand U4193 (N_4193,N_251,N_1007);
xnor U4194 (N_4194,N_875,N_2241);
nand U4195 (N_4195,N_1124,N_756);
nand U4196 (N_4196,N_1159,N_400);
or U4197 (N_4197,N_246,N_1599);
xor U4198 (N_4198,N_1626,N_1894);
xor U4199 (N_4199,N_1548,N_261);
xnor U4200 (N_4200,N_930,N_870);
or U4201 (N_4201,N_665,N_1700);
xor U4202 (N_4202,N_905,N_1122);
or U4203 (N_4203,N_2046,N_738);
or U4204 (N_4204,N_988,N_1530);
nand U4205 (N_4205,N_65,N_1184);
or U4206 (N_4206,N_1292,N_999);
or U4207 (N_4207,N_1806,N_2357);
nand U4208 (N_4208,N_543,N_132);
or U4209 (N_4209,N_597,N_166);
nand U4210 (N_4210,N_1250,N_1044);
and U4211 (N_4211,N_254,N_1879);
nand U4212 (N_4212,N_745,N_2189);
xor U4213 (N_4213,N_305,N_1446);
nand U4214 (N_4214,N_2180,N_1382);
and U4215 (N_4215,N_863,N_1257);
nor U4216 (N_4216,N_2334,N_624);
xor U4217 (N_4217,N_391,N_2327);
nand U4218 (N_4218,N_235,N_1942);
and U4219 (N_4219,N_1361,N_930);
nand U4220 (N_4220,N_14,N_233);
and U4221 (N_4221,N_2297,N_744);
nand U4222 (N_4222,N_1119,N_85);
nand U4223 (N_4223,N_560,N_2189);
or U4224 (N_4224,N_2232,N_2496);
nand U4225 (N_4225,N_2418,N_1716);
and U4226 (N_4226,N_59,N_1207);
and U4227 (N_4227,N_1600,N_1337);
nor U4228 (N_4228,N_1647,N_1337);
nand U4229 (N_4229,N_1936,N_1791);
or U4230 (N_4230,N_1495,N_130);
and U4231 (N_4231,N_2153,N_652);
nor U4232 (N_4232,N_710,N_1218);
or U4233 (N_4233,N_754,N_672);
or U4234 (N_4234,N_1029,N_223);
and U4235 (N_4235,N_927,N_564);
and U4236 (N_4236,N_708,N_790);
nand U4237 (N_4237,N_1500,N_1488);
nand U4238 (N_4238,N_2493,N_2020);
nand U4239 (N_4239,N_1383,N_970);
and U4240 (N_4240,N_1251,N_1467);
xor U4241 (N_4241,N_2434,N_2450);
or U4242 (N_4242,N_1845,N_795);
and U4243 (N_4243,N_299,N_2177);
nor U4244 (N_4244,N_2075,N_1755);
nand U4245 (N_4245,N_183,N_2287);
xor U4246 (N_4246,N_554,N_586);
nor U4247 (N_4247,N_442,N_723);
nand U4248 (N_4248,N_2337,N_1093);
nand U4249 (N_4249,N_1086,N_2096);
nand U4250 (N_4250,N_809,N_2486);
nand U4251 (N_4251,N_634,N_67);
or U4252 (N_4252,N_275,N_1663);
and U4253 (N_4253,N_1008,N_1619);
nand U4254 (N_4254,N_2420,N_1427);
and U4255 (N_4255,N_1835,N_173);
or U4256 (N_4256,N_230,N_305);
nand U4257 (N_4257,N_2244,N_1720);
nand U4258 (N_4258,N_2407,N_1278);
nor U4259 (N_4259,N_1582,N_2085);
nor U4260 (N_4260,N_2361,N_644);
and U4261 (N_4261,N_976,N_983);
or U4262 (N_4262,N_28,N_1127);
nand U4263 (N_4263,N_539,N_1127);
nand U4264 (N_4264,N_605,N_2460);
nor U4265 (N_4265,N_2483,N_517);
nor U4266 (N_4266,N_329,N_639);
or U4267 (N_4267,N_693,N_876);
xnor U4268 (N_4268,N_2266,N_1900);
nand U4269 (N_4269,N_1127,N_542);
nand U4270 (N_4270,N_1299,N_1745);
or U4271 (N_4271,N_763,N_1405);
or U4272 (N_4272,N_726,N_2382);
nor U4273 (N_4273,N_2187,N_48);
xor U4274 (N_4274,N_252,N_1898);
nor U4275 (N_4275,N_1365,N_1137);
and U4276 (N_4276,N_1492,N_2389);
nand U4277 (N_4277,N_610,N_1234);
nand U4278 (N_4278,N_610,N_496);
or U4279 (N_4279,N_1561,N_926);
nor U4280 (N_4280,N_1087,N_1021);
or U4281 (N_4281,N_849,N_584);
or U4282 (N_4282,N_1429,N_189);
nand U4283 (N_4283,N_48,N_826);
and U4284 (N_4284,N_820,N_2384);
nand U4285 (N_4285,N_843,N_679);
and U4286 (N_4286,N_1293,N_2232);
or U4287 (N_4287,N_759,N_1193);
or U4288 (N_4288,N_2229,N_2077);
or U4289 (N_4289,N_2291,N_891);
nor U4290 (N_4290,N_1222,N_1195);
xor U4291 (N_4291,N_1090,N_894);
nor U4292 (N_4292,N_305,N_195);
or U4293 (N_4293,N_1924,N_2402);
or U4294 (N_4294,N_700,N_922);
and U4295 (N_4295,N_2489,N_2096);
and U4296 (N_4296,N_1353,N_2177);
and U4297 (N_4297,N_1391,N_2417);
or U4298 (N_4298,N_1625,N_678);
nand U4299 (N_4299,N_2497,N_2045);
and U4300 (N_4300,N_428,N_212);
or U4301 (N_4301,N_2049,N_1569);
and U4302 (N_4302,N_1797,N_1732);
and U4303 (N_4303,N_789,N_1774);
nand U4304 (N_4304,N_1991,N_244);
or U4305 (N_4305,N_2210,N_2031);
nor U4306 (N_4306,N_1918,N_2110);
and U4307 (N_4307,N_355,N_146);
or U4308 (N_4308,N_43,N_441);
xnor U4309 (N_4309,N_1462,N_656);
or U4310 (N_4310,N_1467,N_907);
or U4311 (N_4311,N_103,N_316);
or U4312 (N_4312,N_369,N_2453);
and U4313 (N_4313,N_845,N_2298);
nor U4314 (N_4314,N_776,N_761);
and U4315 (N_4315,N_1005,N_2339);
nor U4316 (N_4316,N_1218,N_154);
nand U4317 (N_4317,N_1375,N_947);
or U4318 (N_4318,N_977,N_2003);
nand U4319 (N_4319,N_1460,N_620);
nand U4320 (N_4320,N_1540,N_1879);
or U4321 (N_4321,N_1805,N_2206);
or U4322 (N_4322,N_1134,N_715);
nor U4323 (N_4323,N_741,N_762);
nand U4324 (N_4324,N_2488,N_2060);
or U4325 (N_4325,N_1071,N_1821);
nand U4326 (N_4326,N_2491,N_2352);
nand U4327 (N_4327,N_1197,N_1650);
and U4328 (N_4328,N_2487,N_1244);
nor U4329 (N_4329,N_1365,N_669);
and U4330 (N_4330,N_371,N_369);
nand U4331 (N_4331,N_1425,N_291);
nor U4332 (N_4332,N_1746,N_1349);
nand U4333 (N_4333,N_1912,N_714);
nor U4334 (N_4334,N_95,N_2251);
nor U4335 (N_4335,N_591,N_2027);
and U4336 (N_4336,N_2256,N_810);
and U4337 (N_4337,N_822,N_170);
nand U4338 (N_4338,N_1560,N_2298);
or U4339 (N_4339,N_2437,N_1704);
nand U4340 (N_4340,N_1094,N_765);
nand U4341 (N_4341,N_1195,N_1784);
and U4342 (N_4342,N_1078,N_1577);
nor U4343 (N_4343,N_1784,N_393);
and U4344 (N_4344,N_1097,N_344);
and U4345 (N_4345,N_966,N_2495);
nor U4346 (N_4346,N_1680,N_1910);
nand U4347 (N_4347,N_538,N_2349);
or U4348 (N_4348,N_2436,N_1654);
nand U4349 (N_4349,N_2445,N_1226);
or U4350 (N_4350,N_1691,N_983);
nor U4351 (N_4351,N_1054,N_682);
and U4352 (N_4352,N_60,N_473);
and U4353 (N_4353,N_2175,N_345);
nor U4354 (N_4354,N_2186,N_975);
nor U4355 (N_4355,N_117,N_472);
or U4356 (N_4356,N_1639,N_2489);
or U4357 (N_4357,N_1416,N_358);
and U4358 (N_4358,N_775,N_487);
or U4359 (N_4359,N_2241,N_2225);
and U4360 (N_4360,N_1114,N_660);
nand U4361 (N_4361,N_703,N_2188);
nand U4362 (N_4362,N_869,N_1964);
and U4363 (N_4363,N_2091,N_1981);
and U4364 (N_4364,N_1522,N_176);
nor U4365 (N_4365,N_1332,N_2499);
nand U4366 (N_4366,N_1938,N_1918);
nand U4367 (N_4367,N_2478,N_1879);
nor U4368 (N_4368,N_1933,N_1185);
xor U4369 (N_4369,N_120,N_1313);
nor U4370 (N_4370,N_1865,N_519);
xor U4371 (N_4371,N_801,N_2160);
nand U4372 (N_4372,N_938,N_991);
or U4373 (N_4373,N_2401,N_750);
nand U4374 (N_4374,N_89,N_1523);
nor U4375 (N_4375,N_1394,N_800);
nand U4376 (N_4376,N_643,N_1484);
nand U4377 (N_4377,N_1394,N_2016);
or U4378 (N_4378,N_341,N_848);
or U4379 (N_4379,N_1476,N_328);
or U4380 (N_4380,N_1687,N_848);
nand U4381 (N_4381,N_2221,N_994);
and U4382 (N_4382,N_1991,N_837);
xnor U4383 (N_4383,N_2349,N_2200);
nand U4384 (N_4384,N_444,N_2346);
nand U4385 (N_4385,N_1573,N_2293);
or U4386 (N_4386,N_303,N_2076);
or U4387 (N_4387,N_518,N_2130);
and U4388 (N_4388,N_1363,N_509);
nor U4389 (N_4389,N_1065,N_53);
nor U4390 (N_4390,N_1282,N_294);
nand U4391 (N_4391,N_868,N_321);
or U4392 (N_4392,N_1700,N_360);
or U4393 (N_4393,N_874,N_422);
or U4394 (N_4394,N_2486,N_377);
and U4395 (N_4395,N_1921,N_2467);
or U4396 (N_4396,N_2104,N_197);
nor U4397 (N_4397,N_1499,N_2374);
nor U4398 (N_4398,N_1566,N_2231);
nand U4399 (N_4399,N_904,N_2131);
nand U4400 (N_4400,N_1229,N_1734);
and U4401 (N_4401,N_1335,N_791);
nor U4402 (N_4402,N_632,N_1408);
xnor U4403 (N_4403,N_182,N_297);
nand U4404 (N_4404,N_259,N_1630);
and U4405 (N_4405,N_706,N_451);
and U4406 (N_4406,N_1478,N_482);
or U4407 (N_4407,N_279,N_370);
and U4408 (N_4408,N_1257,N_107);
or U4409 (N_4409,N_526,N_1306);
nand U4410 (N_4410,N_2049,N_1682);
and U4411 (N_4411,N_2039,N_425);
and U4412 (N_4412,N_2011,N_696);
xor U4413 (N_4413,N_1801,N_910);
nand U4414 (N_4414,N_1994,N_911);
xnor U4415 (N_4415,N_2286,N_2022);
nor U4416 (N_4416,N_702,N_553);
or U4417 (N_4417,N_2329,N_2403);
nor U4418 (N_4418,N_2075,N_846);
nand U4419 (N_4419,N_973,N_2113);
xnor U4420 (N_4420,N_2016,N_1682);
xnor U4421 (N_4421,N_120,N_914);
nor U4422 (N_4422,N_444,N_651);
nor U4423 (N_4423,N_2196,N_1612);
nor U4424 (N_4424,N_1338,N_1896);
nor U4425 (N_4425,N_969,N_1099);
nand U4426 (N_4426,N_2446,N_1169);
and U4427 (N_4427,N_743,N_1522);
and U4428 (N_4428,N_1618,N_2219);
and U4429 (N_4429,N_1646,N_966);
and U4430 (N_4430,N_200,N_884);
or U4431 (N_4431,N_1518,N_922);
and U4432 (N_4432,N_2323,N_537);
xor U4433 (N_4433,N_1936,N_483);
nand U4434 (N_4434,N_1456,N_1368);
nor U4435 (N_4435,N_1773,N_2025);
xor U4436 (N_4436,N_556,N_485);
nor U4437 (N_4437,N_1354,N_2229);
or U4438 (N_4438,N_959,N_2320);
xnor U4439 (N_4439,N_1877,N_1571);
and U4440 (N_4440,N_2235,N_1648);
and U4441 (N_4441,N_464,N_891);
nand U4442 (N_4442,N_880,N_1558);
nand U4443 (N_4443,N_1471,N_1356);
nand U4444 (N_4444,N_419,N_1815);
or U4445 (N_4445,N_534,N_1866);
nand U4446 (N_4446,N_46,N_1370);
nand U4447 (N_4447,N_2141,N_1828);
or U4448 (N_4448,N_1657,N_836);
xnor U4449 (N_4449,N_215,N_2395);
nor U4450 (N_4450,N_1990,N_2367);
nand U4451 (N_4451,N_645,N_973);
xnor U4452 (N_4452,N_2129,N_1929);
and U4453 (N_4453,N_543,N_85);
and U4454 (N_4454,N_769,N_1239);
and U4455 (N_4455,N_1024,N_382);
nor U4456 (N_4456,N_1698,N_1815);
nand U4457 (N_4457,N_1186,N_1431);
or U4458 (N_4458,N_2162,N_209);
or U4459 (N_4459,N_1807,N_673);
nand U4460 (N_4460,N_1026,N_880);
nand U4461 (N_4461,N_338,N_1752);
and U4462 (N_4462,N_2386,N_1855);
or U4463 (N_4463,N_1911,N_1889);
nand U4464 (N_4464,N_94,N_890);
and U4465 (N_4465,N_2481,N_507);
nor U4466 (N_4466,N_788,N_1203);
or U4467 (N_4467,N_2346,N_2103);
or U4468 (N_4468,N_940,N_1);
nor U4469 (N_4469,N_925,N_1158);
or U4470 (N_4470,N_1175,N_664);
nor U4471 (N_4471,N_1638,N_1588);
and U4472 (N_4472,N_325,N_878);
nand U4473 (N_4473,N_870,N_2207);
nand U4474 (N_4474,N_656,N_1455);
xnor U4475 (N_4475,N_478,N_2114);
nand U4476 (N_4476,N_119,N_844);
and U4477 (N_4477,N_1055,N_2275);
and U4478 (N_4478,N_339,N_2186);
xnor U4479 (N_4479,N_2092,N_684);
or U4480 (N_4480,N_1095,N_2323);
nand U4481 (N_4481,N_1058,N_1163);
nand U4482 (N_4482,N_1024,N_68);
or U4483 (N_4483,N_1663,N_1714);
xnor U4484 (N_4484,N_1203,N_1363);
or U4485 (N_4485,N_2070,N_146);
xnor U4486 (N_4486,N_130,N_441);
xnor U4487 (N_4487,N_1539,N_669);
nand U4488 (N_4488,N_102,N_1208);
nand U4489 (N_4489,N_1445,N_1170);
and U4490 (N_4490,N_641,N_1180);
nand U4491 (N_4491,N_2482,N_203);
or U4492 (N_4492,N_309,N_247);
xnor U4493 (N_4493,N_2204,N_448);
or U4494 (N_4494,N_1930,N_1081);
xnor U4495 (N_4495,N_621,N_1238);
or U4496 (N_4496,N_1140,N_855);
or U4497 (N_4497,N_2197,N_1184);
xor U4498 (N_4498,N_1548,N_979);
xor U4499 (N_4499,N_2397,N_953);
nor U4500 (N_4500,N_714,N_10);
nand U4501 (N_4501,N_207,N_1105);
nand U4502 (N_4502,N_1157,N_1098);
nand U4503 (N_4503,N_1995,N_349);
nand U4504 (N_4504,N_2278,N_395);
nand U4505 (N_4505,N_1301,N_32);
and U4506 (N_4506,N_1902,N_2356);
nor U4507 (N_4507,N_1940,N_432);
or U4508 (N_4508,N_257,N_2308);
or U4509 (N_4509,N_178,N_1255);
and U4510 (N_4510,N_2133,N_8);
nand U4511 (N_4511,N_424,N_2133);
and U4512 (N_4512,N_317,N_2388);
and U4513 (N_4513,N_1591,N_1626);
nand U4514 (N_4514,N_161,N_2451);
nor U4515 (N_4515,N_1205,N_737);
nand U4516 (N_4516,N_873,N_894);
and U4517 (N_4517,N_1660,N_1891);
nand U4518 (N_4518,N_571,N_2338);
nand U4519 (N_4519,N_2158,N_2035);
and U4520 (N_4520,N_781,N_2462);
nor U4521 (N_4521,N_1088,N_415);
nor U4522 (N_4522,N_1940,N_1027);
nor U4523 (N_4523,N_1481,N_425);
and U4524 (N_4524,N_377,N_366);
nor U4525 (N_4525,N_275,N_1736);
xor U4526 (N_4526,N_509,N_471);
xor U4527 (N_4527,N_720,N_1090);
nor U4528 (N_4528,N_213,N_873);
nand U4529 (N_4529,N_971,N_1815);
xor U4530 (N_4530,N_1542,N_1099);
or U4531 (N_4531,N_1580,N_1196);
and U4532 (N_4532,N_2062,N_494);
xnor U4533 (N_4533,N_1971,N_279);
and U4534 (N_4534,N_359,N_1318);
nor U4535 (N_4535,N_1868,N_786);
or U4536 (N_4536,N_712,N_1511);
nand U4537 (N_4537,N_2034,N_49);
nor U4538 (N_4538,N_1710,N_2152);
nor U4539 (N_4539,N_683,N_1690);
or U4540 (N_4540,N_1590,N_415);
or U4541 (N_4541,N_154,N_754);
and U4542 (N_4542,N_1358,N_1218);
nor U4543 (N_4543,N_1678,N_2272);
xnor U4544 (N_4544,N_1280,N_345);
nor U4545 (N_4545,N_2351,N_2037);
nand U4546 (N_4546,N_2295,N_1236);
nand U4547 (N_4547,N_1566,N_63);
nand U4548 (N_4548,N_857,N_2205);
xor U4549 (N_4549,N_1158,N_1216);
nor U4550 (N_4550,N_242,N_2322);
and U4551 (N_4551,N_1030,N_1100);
nand U4552 (N_4552,N_325,N_738);
nor U4553 (N_4553,N_214,N_1259);
nor U4554 (N_4554,N_2453,N_74);
xnor U4555 (N_4555,N_281,N_1538);
nand U4556 (N_4556,N_139,N_1681);
and U4557 (N_4557,N_1434,N_1600);
and U4558 (N_4558,N_1020,N_1721);
nor U4559 (N_4559,N_1030,N_1834);
nor U4560 (N_4560,N_1877,N_1915);
nor U4561 (N_4561,N_2493,N_1784);
nand U4562 (N_4562,N_1364,N_2114);
and U4563 (N_4563,N_942,N_1360);
and U4564 (N_4564,N_404,N_2122);
nand U4565 (N_4565,N_1708,N_21);
or U4566 (N_4566,N_1150,N_657);
nor U4567 (N_4567,N_1008,N_888);
nor U4568 (N_4568,N_379,N_1002);
xnor U4569 (N_4569,N_1756,N_1477);
xor U4570 (N_4570,N_1132,N_134);
nand U4571 (N_4571,N_2327,N_1580);
or U4572 (N_4572,N_811,N_1379);
and U4573 (N_4573,N_1857,N_2146);
or U4574 (N_4574,N_1248,N_2020);
nor U4575 (N_4575,N_1791,N_900);
nand U4576 (N_4576,N_973,N_451);
nor U4577 (N_4577,N_135,N_2284);
nand U4578 (N_4578,N_1247,N_1747);
or U4579 (N_4579,N_933,N_2152);
and U4580 (N_4580,N_2308,N_753);
nor U4581 (N_4581,N_1049,N_1876);
xnor U4582 (N_4582,N_1200,N_53);
nor U4583 (N_4583,N_390,N_1758);
xor U4584 (N_4584,N_2058,N_2404);
and U4585 (N_4585,N_2269,N_1934);
nor U4586 (N_4586,N_1104,N_1597);
and U4587 (N_4587,N_1218,N_2387);
nand U4588 (N_4588,N_1213,N_289);
or U4589 (N_4589,N_873,N_356);
and U4590 (N_4590,N_1632,N_1625);
and U4591 (N_4591,N_1596,N_37);
nand U4592 (N_4592,N_1180,N_1414);
nor U4593 (N_4593,N_1637,N_2231);
xnor U4594 (N_4594,N_813,N_328);
nor U4595 (N_4595,N_1709,N_180);
nand U4596 (N_4596,N_1226,N_331);
or U4597 (N_4597,N_1178,N_1322);
or U4598 (N_4598,N_2123,N_1202);
nor U4599 (N_4599,N_2026,N_1301);
and U4600 (N_4600,N_105,N_1014);
nand U4601 (N_4601,N_1212,N_739);
nor U4602 (N_4602,N_1863,N_1156);
and U4603 (N_4603,N_290,N_1776);
nor U4604 (N_4604,N_1117,N_410);
xor U4605 (N_4605,N_1787,N_1280);
nand U4606 (N_4606,N_1242,N_1221);
nand U4607 (N_4607,N_1531,N_913);
or U4608 (N_4608,N_1788,N_781);
or U4609 (N_4609,N_973,N_1704);
nand U4610 (N_4610,N_2380,N_1470);
and U4611 (N_4611,N_1580,N_1019);
and U4612 (N_4612,N_2493,N_1651);
or U4613 (N_4613,N_1177,N_321);
nand U4614 (N_4614,N_1999,N_806);
or U4615 (N_4615,N_691,N_1663);
or U4616 (N_4616,N_2255,N_1271);
nor U4617 (N_4617,N_404,N_1343);
nand U4618 (N_4618,N_2094,N_1118);
nor U4619 (N_4619,N_2273,N_1384);
nand U4620 (N_4620,N_1757,N_2462);
or U4621 (N_4621,N_653,N_1905);
and U4622 (N_4622,N_1784,N_986);
nor U4623 (N_4623,N_1426,N_1009);
or U4624 (N_4624,N_785,N_303);
and U4625 (N_4625,N_2432,N_1251);
nand U4626 (N_4626,N_987,N_772);
or U4627 (N_4627,N_137,N_1804);
nor U4628 (N_4628,N_552,N_696);
nor U4629 (N_4629,N_933,N_2331);
xor U4630 (N_4630,N_472,N_1219);
nand U4631 (N_4631,N_703,N_2273);
nor U4632 (N_4632,N_693,N_1831);
or U4633 (N_4633,N_394,N_1316);
and U4634 (N_4634,N_1142,N_1683);
nand U4635 (N_4635,N_1272,N_2183);
nor U4636 (N_4636,N_1078,N_811);
and U4637 (N_4637,N_1013,N_268);
and U4638 (N_4638,N_35,N_1429);
or U4639 (N_4639,N_2178,N_44);
nand U4640 (N_4640,N_1044,N_828);
and U4641 (N_4641,N_64,N_2276);
or U4642 (N_4642,N_1251,N_824);
and U4643 (N_4643,N_2037,N_1403);
and U4644 (N_4644,N_2185,N_43);
or U4645 (N_4645,N_221,N_1884);
nand U4646 (N_4646,N_1429,N_1957);
nand U4647 (N_4647,N_347,N_2235);
nor U4648 (N_4648,N_2427,N_1816);
or U4649 (N_4649,N_1010,N_1415);
nand U4650 (N_4650,N_667,N_1368);
or U4651 (N_4651,N_2224,N_240);
nand U4652 (N_4652,N_2284,N_1107);
nor U4653 (N_4653,N_2422,N_411);
and U4654 (N_4654,N_2259,N_258);
or U4655 (N_4655,N_407,N_708);
or U4656 (N_4656,N_488,N_1882);
and U4657 (N_4657,N_879,N_1114);
and U4658 (N_4658,N_1352,N_1112);
or U4659 (N_4659,N_2344,N_2121);
nor U4660 (N_4660,N_1447,N_2030);
nand U4661 (N_4661,N_503,N_1064);
and U4662 (N_4662,N_2144,N_726);
nor U4663 (N_4663,N_1738,N_1768);
nor U4664 (N_4664,N_1787,N_1119);
nand U4665 (N_4665,N_2280,N_2489);
and U4666 (N_4666,N_2065,N_1410);
or U4667 (N_4667,N_231,N_59);
and U4668 (N_4668,N_598,N_488);
and U4669 (N_4669,N_2065,N_2304);
xor U4670 (N_4670,N_191,N_2217);
nor U4671 (N_4671,N_2205,N_632);
and U4672 (N_4672,N_819,N_1526);
nand U4673 (N_4673,N_1612,N_1082);
or U4674 (N_4674,N_1845,N_735);
nand U4675 (N_4675,N_985,N_1283);
or U4676 (N_4676,N_892,N_2171);
and U4677 (N_4677,N_641,N_322);
and U4678 (N_4678,N_1633,N_982);
nand U4679 (N_4679,N_1980,N_585);
nand U4680 (N_4680,N_2266,N_99);
nand U4681 (N_4681,N_327,N_837);
and U4682 (N_4682,N_837,N_2379);
nand U4683 (N_4683,N_968,N_2362);
or U4684 (N_4684,N_1483,N_1160);
nand U4685 (N_4685,N_2328,N_241);
and U4686 (N_4686,N_1554,N_752);
nand U4687 (N_4687,N_1971,N_2231);
or U4688 (N_4688,N_957,N_832);
nand U4689 (N_4689,N_523,N_106);
nor U4690 (N_4690,N_153,N_420);
or U4691 (N_4691,N_2064,N_250);
nand U4692 (N_4692,N_983,N_1010);
xnor U4693 (N_4693,N_1134,N_565);
and U4694 (N_4694,N_301,N_2038);
nand U4695 (N_4695,N_332,N_560);
nand U4696 (N_4696,N_2439,N_781);
nand U4697 (N_4697,N_1249,N_149);
nor U4698 (N_4698,N_1801,N_1056);
nor U4699 (N_4699,N_2499,N_303);
nand U4700 (N_4700,N_1290,N_1240);
nand U4701 (N_4701,N_1508,N_965);
and U4702 (N_4702,N_976,N_1615);
or U4703 (N_4703,N_1341,N_879);
nor U4704 (N_4704,N_1503,N_381);
and U4705 (N_4705,N_1864,N_650);
nor U4706 (N_4706,N_776,N_1236);
nor U4707 (N_4707,N_1134,N_2486);
and U4708 (N_4708,N_2462,N_1436);
or U4709 (N_4709,N_1822,N_2398);
or U4710 (N_4710,N_1004,N_1036);
nand U4711 (N_4711,N_2354,N_1774);
and U4712 (N_4712,N_1675,N_788);
and U4713 (N_4713,N_1559,N_635);
and U4714 (N_4714,N_308,N_715);
nor U4715 (N_4715,N_1721,N_1557);
xnor U4716 (N_4716,N_279,N_1246);
and U4717 (N_4717,N_1420,N_2058);
xor U4718 (N_4718,N_1798,N_818);
or U4719 (N_4719,N_366,N_634);
and U4720 (N_4720,N_2200,N_1919);
or U4721 (N_4721,N_2009,N_909);
and U4722 (N_4722,N_612,N_2481);
nor U4723 (N_4723,N_1414,N_1283);
nor U4724 (N_4724,N_2415,N_503);
and U4725 (N_4725,N_2278,N_927);
or U4726 (N_4726,N_1069,N_2495);
nand U4727 (N_4727,N_1293,N_2383);
and U4728 (N_4728,N_410,N_1984);
or U4729 (N_4729,N_1704,N_36);
nor U4730 (N_4730,N_342,N_2203);
and U4731 (N_4731,N_1277,N_803);
xor U4732 (N_4732,N_2185,N_1030);
nand U4733 (N_4733,N_981,N_1427);
and U4734 (N_4734,N_904,N_452);
or U4735 (N_4735,N_1520,N_276);
or U4736 (N_4736,N_476,N_1328);
nor U4737 (N_4737,N_1287,N_2273);
nor U4738 (N_4738,N_780,N_971);
and U4739 (N_4739,N_1433,N_1859);
nor U4740 (N_4740,N_817,N_2123);
and U4741 (N_4741,N_2221,N_2262);
nand U4742 (N_4742,N_25,N_593);
or U4743 (N_4743,N_479,N_419);
nand U4744 (N_4744,N_1349,N_625);
and U4745 (N_4745,N_2182,N_2428);
and U4746 (N_4746,N_1284,N_2234);
or U4747 (N_4747,N_588,N_1508);
and U4748 (N_4748,N_1313,N_1013);
xor U4749 (N_4749,N_1393,N_963);
or U4750 (N_4750,N_1796,N_228);
and U4751 (N_4751,N_2068,N_427);
nand U4752 (N_4752,N_2345,N_1919);
and U4753 (N_4753,N_62,N_1475);
nand U4754 (N_4754,N_2219,N_847);
nor U4755 (N_4755,N_2192,N_2225);
nor U4756 (N_4756,N_1773,N_1897);
and U4757 (N_4757,N_2049,N_506);
nor U4758 (N_4758,N_2495,N_1123);
nand U4759 (N_4759,N_2369,N_1014);
nand U4760 (N_4760,N_1981,N_1498);
nand U4761 (N_4761,N_1367,N_1533);
nor U4762 (N_4762,N_193,N_1134);
nor U4763 (N_4763,N_283,N_1852);
or U4764 (N_4764,N_69,N_1500);
and U4765 (N_4765,N_633,N_2335);
nand U4766 (N_4766,N_857,N_1215);
nor U4767 (N_4767,N_1288,N_1144);
or U4768 (N_4768,N_2154,N_930);
or U4769 (N_4769,N_2179,N_58);
nand U4770 (N_4770,N_1841,N_1296);
nor U4771 (N_4771,N_1259,N_2156);
nor U4772 (N_4772,N_719,N_1233);
and U4773 (N_4773,N_1347,N_496);
or U4774 (N_4774,N_556,N_587);
or U4775 (N_4775,N_1892,N_1765);
xnor U4776 (N_4776,N_738,N_753);
nor U4777 (N_4777,N_2430,N_539);
or U4778 (N_4778,N_80,N_790);
nand U4779 (N_4779,N_1060,N_261);
nor U4780 (N_4780,N_1559,N_1538);
or U4781 (N_4781,N_1945,N_1232);
nand U4782 (N_4782,N_1232,N_112);
and U4783 (N_4783,N_1508,N_1296);
and U4784 (N_4784,N_1229,N_1574);
nand U4785 (N_4785,N_864,N_852);
xnor U4786 (N_4786,N_1979,N_549);
or U4787 (N_4787,N_889,N_2353);
and U4788 (N_4788,N_2338,N_1796);
and U4789 (N_4789,N_1901,N_2112);
nor U4790 (N_4790,N_997,N_1716);
and U4791 (N_4791,N_1697,N_437);
nor U4792 (N_4792,N_1429,N_687);
nor U4793 (N_4793,N_1985,N_1879);
nand U4794 (N_4794,N_680,N_936);
nand U4795 (N_4795,N_1691,N_275);
and U4796 (N_4796,N_1023,N_1007);
or U4797 (N_4797,N_1523,N_1851);
or U4798 (N_4798,N_1785,N_260);
and U4799 (N_4799,N_295,N_214);
or U4800 (N_4800,N_1742,N_1867);
nor U4801 (N_4801,N_1075,N_1811);
nand U4802 (N_4802,N_1903,N_1995);
nor U4803 (N_4803,N_201,N_1458);
or U4804 (N_4804,N_241,N_362);
and U4805 (N_4805,N_1330,N_1005);
nand U4806 (N_4806,N_1280,N_154);
and U4807 (N_4807,N_1823,N_1311);
nor U4808 (N_4808,N_818,N_1186);
and U4809 (N_4809,N_2069,N_888);
or U4810 (N_4810,N_1894,N_2355);
or U4811 (N_4811,N_2246,N_497);
xor U4812 (N_4812,N_1841,N_2309);
nand U4813 (N_4813,N_924,N_2129);
and U4814 (N_4814,N_1612,N_334);
or U4815 (N_4815,N_139,N_1500);
nor U4816 (N_4816,N_1998,N_2430);
or U4817 (N_4817,N_547,N_1773);
or U4818 (N_4818,N_32,N_1089);
or U4819 (N_4819,N_39,N_1055);
or U4820 (N_4820,N_2095,N_1539);
nand U4821 (N_4821,N_2041,N_1144);
and U4822 (N_4822,N_2317,N_781);
and U4823 (N_4823,N_1378,N_106);
or U4824 (N_4824,N_897,N_739);
and U4825 (N_4825,N_339,N_465);
nand U4826 (N_4826,N_863,N_1018);
xnor U4827 (N_4827,N_1153,N_60);
and U4828 (N_4828,N_426,N_1175);
and U4829 (N_4829,N_760,N_1383);
or U4830 (N_4830,N_1845,N_1689);
nor U4831 (N_4831,N_965,N_2273);
nand U4832 (N_4832,N_28,N_2378);
xor U4833 (N_4833,N_2268,N_1211);
and U4834 (N_4834,N_52,N_803);
nand U4835 (N_4835,N_2446,N_1419);
nand U4836 (N_4836,N_1507,N_1184);
xor U4837 (N_4837,N_1452,N_418);
nor U4838 (N_4838,N_314,N_2201);
nor U4839 (N_4839,N_495,N_1300);
and U4840 (N_4840,N_1167,N_559);
nand U4841 (N_4841,N_1574,N_1549);
and U4842 (N_4842,N_252,N_2201);
nor U4843 (N_4843,N_123,N_1506);
and U4844 (N_4844,N_1591,N_2470);
xnor U4845 (N_4845,N_1520,N_1206);
nand U4846 (N_4846,N_1776,N_1976);
and U4847 (N_4847,N_2052,N_584);
nor U4848 (N_4848,N_1883,N_2076);
nand U4849 (N_4849,N_1158,N_1876);
nand U4850 (N_4850,N_937,N_417);
or U4851 (N_4851,N_543,N_1560);
or U4852 (N_4852,N_1770,N_2198);
and U4853 (N_4853,N_739,N_2083);
nor U4854 (N_4854,N_677,N_1988);
nand U4855 (N_4855,N_1430,N_1617);
or U4856 (N_4856,N_1112,N_570);
or U4857 (N_4857,N_1437,N_1982);
nor U4858 (N_4858,N_699,N_260);
and U4859 (N_4859,N_1830,N_2061);
and U4860 (N_4860,N_2000,N_2075);
or U4861 (N_4861,N_1616,N_588);
and U4862 (N_4862,N_1106,N_2204);
or U4863 (N_4863,N_2460,N_1169);
nor U4864 (N_4864,N_559,N_2443);
or U4865 (N_4865,N_1311,N_838);
and U4866 (N_4866,N_1923,N_2242);
xor U4867 (N_4867,N_11,N_855);
nor U4868 (N_4868,N_611,N_765);
or U4869 (N_4869,N_2161,N_761);
nand U4870 (N_4870,N_2050,N_1653);
nand U4871 (N_4871,N_401,N_528);
nand U4872 (N_4872,N_1584,N_456);
nand U4873 (N_4873,N_2214,N_374);
nor U4874 (N_4874,N_2038,N_766);
xor U4875 (N_4875,N_1080,N_2243);
xor U4876 (N_4876,N_977,N_1129);
xor U4877 (N_4877,N_487,N_1333);
or U4878 (N_4878,N_2209,N_2001);
and U4879 (N_4879,N_372,N_1871);
nor U4880 (N_4880,N_2285,N_2229);
or U4881 (N_4881,N_1531,N_437);
nor U4882 (N_4882,N_1993,N_362);
xnor U4883 (N_4883,N_1378,N_1107);
nand U4884 (N_4884,N_13,N_1022);
nor U4885 (N_4885,N_993,N_2035);
nor U4886 (N_4886,N_2218,N_1399);
and U4887 (N_4887,N_2322,N_1008);
nand U4888 (N_4888,N_936,N_1079);
or U4889 (N_4889,N_1924,N_752);
nand U4890 (N_4890,N_1747,N_2059);
nand U4891 (N_4891,N_1988,N_1725);
nor U4892 (N_4892,N_161,N_1367);
nor U4893 (N_4893,N_1537,N_42);
xor U4894 (N_4894,N_614,N_517);
and U4895 (N_4895,N_419,N_537);
or U4896 (N_4896,N_536,N_1315);
and U4897 (N_4897,N_2021,N_751);
nand U4898 (N_4898,N_1314,N_1157);
nor U4899 (N_4899,N_171,N_557);
nor U4900 (N_4900,N_1581,N_558);
nor U4901 (N_4901,N_1345,N_1400);
and U4902 (N_4902,N_1821,N_2077);
nor U4903 (N_4903,N_2134,N_55);
nand U4904 (N_4904,N_1126,N_2177);
and U4905 (N_4905,N_557,N_552);
nor U4906 (N_4906,N_1421,N_1892);
nand U4907 (N_4907,N_2255,N_2288);
nand U4908 (N_4908,N_1398,N_1944);
nand U4909 (N_4909,N_558,N_303);
and U4910 (N_4910,N_1977,N_873);
and U4911 (N_4911,N_2395,N_86);
or U4912 (N_4912,N_372,N_589);
nand U4913 (N_4913,N_1868,N_469);
xor U4914 (N_4914,N_444,N_1274);
xor U4915 (N_4915,N_923,N_1211);
or U4916 (N_4916,N_568,N_115);
nand U4917 (N_4917,N_335,N_60);
nor U4918 (N_4918,N_727,N_1942);
xnor U4919 (N_4919,N_900,N_441);
nand U4920 (N_4920,N_218,N_1506);
and U4921 (N_4921,N_2447,N_94);
and U4922 (N_4922,N_1850,N_314);
nand U4923 (N_4923,N_704,N_830);
xnor U4924 (N_4924,N_2320,N_2045);
nand U4925 (N_4925,N_470,N_1696);
or U4926 (N_4926,N_703,N_2162);
nor U4927 (N_4927,N_2136,N_2454);
or U4928 (N_4928,N_2068,N_2300);
nor U4929 (N_4929,N_180,N_855);
nand U4930 (N_4930,N_923,N_815);
nor U4931 (N_4931,N_1536,N_1693);
nor U4932 (N_4932,N_122,N_86);
nor U4933 (N_4933,N_1412,N_2194);
and U4934 (N_4934,N_646,N_1113);
or U4935 (N_4935,N_1829,N_1855);
or U4936 (N_4936,N_1628,N_221);
and U4937 (N_4937,N_1611,N_1404);
xor U4938 (N_4938,N_556,N_1675);
and U4939 (N_4939,N_1612,N_317);
and U4940 (N_4940,N_239,N_1774);
nand U4941 (N_4941,N_1805,N_1302);
nor U4942 (N_4942,N_1858,N_40);
or U4943 (N_4943,N_674,N_753);
nand U4944 (N_4944,N_611,N_2478);
xnor U4945 (N_4945,N_2458,N_1530);
and U4946 (N_4946,N_1894,N_147);
xor U4947 (N_4947,N_1170,N_2294);
nor U4948 (N_4948,N_1063,N_515);
nand U4949 (N_4949,N_1458,N_2420);
or U4950 (N_4950,N_1019,N_2076);
nor U4951 (N_4951,N_502,N_977);
nand U4952 (N_4952,N_1308,N_904);
nor U4953 (N_4953,N_66,N_2402);
or U4954 (N_4954,N_1036,N_1719);
and U4955 (N_4955,N_2169,N_937);
xnor U4956 (N_4956,N_17,N_1031);
nand U4957 (N_4957,N_1762,N_2280);
nand U4958 (N_4958,N_101,N_974);
nor U4959 (N_4959,N_1826,N_1497);
or U4960 (N_4960,N_821,N_2432);
or U4961 (N_4961,N_961,N_1358);
nor U4962 (N_4962,N_2047,N_1904);
or U4963 (N_4963,N_1025,N_1974);
nor U4964 (N_4964,N_386,N_1127);
nand U4965 (N_4965,N_949,N_1176);
or U4966 (N_4966,N_1157,N_293);
xor U4967 (N_4967,N_1292,N_1397);
and U4968 (N_4968,N_2371,N_846);
and U4969 (N_4969,N_988,N_1049);
and U4970 (N_4970,N_1049,N_603);
nand U4971 (N_4971,N_1133,N_1197);
xor U4972 (N_4972,N_1291,N_659);
nor U4973 (N_4973,N_1464,N_1199);
nand U4974 (N_4974,N_1695,N_2233);
nand U4975 (N_4975,N_1978,N_799);
and U4976 (N_4976,N_1647,N_2);
nor U4977 (N_4977,N_1968,N_943);
and U4978 (N_4978,N_94,N_1058);
nor U4979 (N_4979,N_1088,N_119);
xor U4980 (N_4980,N_527,N_1406);
or U4981 (N_4981,N_642,N_1180);
and U4982 (N_4982,N_2379,N_816);
xnor U4983 (N_4983,N_2262,N_348);
nor U4984 (N_4984,N_821,N_1946);
or U4985 (N_4985,N_544,N_89);
and U4986 (N_4986,N_2257,N_1699);
nand U4987 (N_4987,N_243,N_1250);
nor U4988 (N_4988,N_2013,N_1029);
or U4989 (N_4989,N_1020,N_1357);
or U4990 (N_4990,N_2089,N_2437);
or U4991 (N_4991,N_642,N_1352);
nor U4992 (N_4992,N_671,N_173);
nand U4993 (N_4993,N_605,N_1374);
nor U4994 (N_4994,N_170,N_1475);
or U4995 (N_4995,N_935,N_504);
nand U4996 (N_4996,N_847,N_2402);
nand U4997 (N_4997,N_2092,N_804);
xor U4998 (N_4998,N_2387,N_2490);
nor U4999 (N_4999,N_2375,N_2349);
nand U5000 (N_5000,N_2928,N_4532);
nor U5001 (N_5001,N_3459,N_3863);
and U5002 (N_5002,N_2854,N_4877);
nand U5003 (N_5003,N_4831,N_3775);
or U5004 (N_5004,N_4788,N_2639);
and U5005 (N_5005,N_4291,N_4215);
and U5006 (N_5006,N_3925,N_4141);
nand U5007 (N_5007,N_3632,N_3498);
xnor U5008 (N_5008,N_4167,N_3848);
or U5009 (N_5009,N_2815,N_2843);
or U5010 (N_5010,N_3698,N_4004);
nor U5011 (N_5011,N_2959,N_3267);
and U5012 (N_5012,N_2985,N_4903);
nor U5013 (N_5013,N_4949,N_4499);
nor U5014 (N_5014,N_4667,N_4270);
xnor U5015 (N_5015,N_4992,N_3549);
nor U5016 (N_5016,N_4401,N_4128);
nand U5017 (N_5017,N_3416,N_4720);
nand U5018 (N_5018,N_4165,N_4147);
nor U5019 (N_5019,N_4380,N_3676);
and U5020 (N_5020,N_4595,N_2666);
or U5021 (N_5021,N_3835,N_4111);
and U5022 (N_5022,N_4103,N_2915);
and U5023 (N_5023,N_2587,N_4072);
xnor U5024 (N_5024,N_2632,N_3983);
and U5025 (N_5025,N_2966,N_4222);
or U5026 (N_5026,N_4299,N_3051);
nor U5027 (N_5027,N_3011,N_4334);
or U5028 (N_5028,N_4540,N_3304);
nand U5029 (N_5029,N_4233,N_2547);
nor U5030 (N_5030,N_3747,N_4606);
or U5031 (N_5031,N_4089,N_3430);
nand U5032 (N_5032,N_4551,N_4657);
nand U5033 (N_5033,N_3212,N_4898);
and U5034 (N_5034,N_4488,N_3478);
nor U5035 (N_5035,N_3619,N_3724);
or U5036 (N_5036,N_2624,N_3474);
or U5037 (N_5037,N_2820,N_4535);
and U5038 (N_5038,N_3907,N_4712);
xnor U5039 (N_5039,N_3223,N_3448);
nor U5040 (N_5040,N_3940,N_2531);
xor U5041 (N_5041,N_3268,N_3510);
and U5042 (N_5042,N_3797,N_3854);
nand U5043 (N_5043,N_2855,N_2528);
and U5044 (N_5044,N_4655,N_4224);
nor U5045 (N_5045,N_2500,N_3326);
or U5046 (N_5046,N_2705,N_4560);
xnor U5047 (N_5047,N_2916,N_3528);
nand U5048 (N_5048,N_4910,N_3605);
nor U5049 (N_5049,N_4973,N_3948);
and U5050 (N_5050,N_2782,N_3229);
nor U5051 (N_5051,N_3045,N_2672);
or U5052 (N_5052,N_2912,N_3104);
xnor U5053 (N_5053,N_4410,N_4879);
and U5054 (N_5054,N_2670,N_3793);
nand U5055 (N_5055,N_2751,N_4544);
or U5056 (N_5056,N_3471,N_4867);
and U5057 (N_5057,N_4428,N_3396);
nand U5058 (N_5058,N_2623,N_3830);
nand U5059 (N_5059,N_4340,N_2834);
nand U5060 (N_5060,N_3672,N_4028);
nor U5061 (N_5061,N_2935,N_4901);
nand U5062 (N_5062,N_2700,N_3577);
or U5063 (N_5063,N_4304,N_2680);
nor U5064 (N_5064,N_2960,N_4302);
or U5065 (N_5065,N_3062,N_2553);
nand U5066 (N_5066,N_3462,N_3303);
or U5067 (N_5067,N_3222,N_3359);
or U5068 (N_5068,N_4939,N_3870);
nor U5069 (N_5069,N_2536,N_3939);
and U5070 (N_5070,N_4908,N_3754);
xor U5071 (N_5071,N_3923,N_3700);
nand U5072 (N_5072,N_3386,N_4433);
and U5073 (N_5073,N_3401,N_4126);
or U5074 (N_5074,N_4173,N_4647);
nor U5075 (N_5075,N_3002,N_3817);
nor U5076 (N_5076,N_4207,N_3084);
nor U5077 (N_5077,N_4639,N_2932);
xnor U5078 (N_5078,N_3112,N_4883);
or U5079 (N_5079,N_3217,N_3391);
and U5080 (N_5080,N_3365,N_4842);
nand U5081 (N_5081,N_4256,N_2699);
nor U5082 (N_5082,N_4691,N_4050);
nor U5083 (N_5083,N_3890,N_3746);
or U5084 (N_5084,N_3145,N_4443);
and U5085 (N_5085,N_2584,N_4286);
nor U5086 (N_5086,N_3137,N_4849);
or U5087 (N_5087,N_3331,N_3647);
or U5088 (N_5088,N_4725,N_4799);
or U5089 (N_5089,N_4959,N_4646);
nor U5090 (N_5090,N_4427,N_2723);
nand U5091 (N_5091,N_4569,N_3920);
and U5092 (N_5092,N_2669,N_4988);
nor U5093 (N_5093,N_3468,N_4912);
or U5094 (N_5094,N_4191,N_3434);
or U5095 (N_5095,N_3150,N_3418);
and U5096 (N_5096,N_4047,N_3133);
nor U5097 (N_5097,N_2571,N_3688);
or U5098 (N_5098,N_2636,N_4658);
or U5099 (N_5099,N_4529,N_2775);
nor U5100 (N_5100,N_2873,N_3839);
or U5101 (N_5101,N_3562,N_4746);
nand U5102 (N_5102,N_2545,N_3307);
and U5103 (N_5103,N_3057,N_4176);
or U5104 (N_5104,N_3806,N_3796);
nand U5105 (N_5105,N_3203,N_4208);
or U5106 (N_5106,N_4313,N_3291);
or U5107 (N_5107,N_2602,N_2538);
xnor U5108 (N_5108,N_3350,N_3515);
nor U5109 (N_5109,N_2607,N_4916);
nand U5110 (N_5110,N_3997,N_4837);
and U5111 (N_5111,N_3009,N_4836);
or U5112 (N_5112,N_3371,N_4461);
and U5113 (N_5113,N_2823,N_4755);
nand U5114 (N_5114,N_4818,N_3302);
nor U5115 (N_5115,N_3597,N_3574);
nor U5116 (N_5116,N_4926,N_2936);
and U5117 (N_5117,N_4151,N_3687);
and U5118 (N_5118,N_2885,N_2920);
xnor U5119 (N_5119,N_3306,N_4169);
nor U5120 (N_5120,N_3706,N_2662);
nor U5121 (N_5121,N_3224,N_4938);
or U5122 (N_5122,N_4360,N_3380);
and U5123 (N_5123,N_2786,N_3157);
xor U5124 (N_5124,N_3208,N_3893);
or U5125 (N_5125,N_3546,N_4106);
or U5126 (N_5126,N_2987,N_3548);
nor U5127 (N_5127,N_4697,N_3825);
and U5128 (N_5128,N_4174,N_4932);
or U5129 (N_5129,N_3666,N_4756);
nor U5130 (N_5130,N_4163,N_2948);
nor U5131 (N_5131,N_3385,N_3991);
nor U5132 (N_5132,N_3532,N_3878);
xnor U5133 (N_5133,N_2791,N_3637);
or U5134 (N_5134,N_3657,N_3384);
nand U5135 (N_5135,N_2645,N_3663);
and U5136 (N_5136,N_4227,N_3375);
nand U5137 (N_5137,N_2809,N_3937);
nand U5138 (N_5138,N_3942,N_2509);
nor U5139 (N_5139,N_4265,N_3076);
or U5140 (N_5140,N_4006,N_3193);
nand U5141 (N_5141,N_3495,N_4485);
and U5142 (N_5142,N_4087,N_3093);
or U5143 (N_5143,N_2781,N_3862);
nand U5144 (N_5144,N_2917,N_4424);
and U5145 (N_5145,N_4052,N_2958);
and U5146 (N_5146,N_2996,N_4924);
or U5147 (N_5147,N_3541,N_3564);
nor U5148 (N_5148,N_2761,N_2657);
and U5149 (N_5149,N_2530,N_4328);
and U5150 (N_5150,N_3711,N_3974);
nor U5151 (N_5151,N_2621,N_4094);
or U5152 (N_5152,N_3768,N_4796);
xor U5153 (N_5153,N_4001,N_2594);
nor U5154 (N_5154,N_2727,N_3503);
and U5155 (N_5155,N_2846,N_4195);
xnor U5156 (N_5156,N_2828,N_2541);
and U5157 (N_5157,N_2519,N_3833);
and U5158 (N_5158,N_4280,N_3636);
and U5159 (N_5159,N_3322,N_2909);
and U5160 (N_5160,N_3725,N_4586);
nand U5161 (N_5161,N_3432,N_4377);
or U5162 (N_5162,N_4777,N_3653);
xor U5163 (N_5163,N_3239,N_3684);
and U5164 (N_5164,N_3346,N_4391);
nand U5165 (N_5165,N_2676,N_4507);
and U5166 (N_5166,N_3595,N_2930);
nor U5167 (N_5167,N_3318,N_2655);
nor U5168 (N_5168,N_2914,N_2868);
nand U5169 (N_5169,N_3282,N_4858);
or U5170 (N_5170,N_3140,N_4269);
nor U5171 (N_5171,N_3590,N_3691);
nor U5172 (N_5172,N_4948,N_4951);
nand U5173 (N_5173,N_4766,N_4578);
xnor U5174 (N_5174,N_2738,N_3828);
nand U5175 (N_5175,N_3583,N_4735);
nor U5176 (N_5176,N_4374,N_3263);
or U5177 (N_5177,N_3857,N_3316);
or U5178 (N_5178,N_3629,N_4049);
and U5179 (N_5179,N_4656,N_2535);
nor U5180 (N_5180,N_4929,N_3994);
nand U5181 (N_5181,N_3230,N_3352);
nor U5182 (N_5182,N_2808,N_4022);
or U5183 (N_5183,N_2858,N_3205);
and U5184 (N_5184,N_4841,N_3177);
or U5185 (N_5185,N_4142,N_4534);
nor U5186 (N_5186,N_3146,N_2899);
and U5187 (N_5187,N_4415,N_4283);
or U5188 (N_5188,N_4029,N_3330);
xor U5189 (N_5189,N_3425,N_4585);
and U5190 (N_5190,N_2897,N_3873);
and U5191 (N_5191,N_4454,N_3399);
and U5192 (N_5192,N_3269,N_3074);
nor U5193 (N_5193,N_4827,N_3897);
nand U5194 (N_5194,N_4359,N_4431);
and U5195 (N_5195,N_4825,N_2522);
nand U5196 (N_5196,N_4348,N_4565);
nor U5197 (N_5197,N_2927,N_2992);
nand U5198 (N_5198,N_3850,N_3447);
or U5199 (N_5199,N_4486,N_3918);
and U5200 (N_5200,N_3098,N_2778);
nor U5201 (N_5201,N_4341,N_3034);
xnor U5202 (N_5202,N_3877,N_2622);
or U5203 (N_5203,N_2586,N_4465);
and U5204 (N_5204,N_4407,N_4617);
xnor U5205 (N_5205,N_2882,N_3790);
nand U5206 (N_5206,N_3395,N_2863);
nand U5207 (N_5207,N_4146,N_2982);
xor U5208 (N_5208,N_4297,N_4076);
xnor U5209 (N_5209,N_4091,N_2848);
and U5210 (N_5210,N_4744,N_3433);
nor U5211 (N_5211,N_3978,N_2902);
or U5212 (N_5212,N_2633,N_4798);
xor U5213 (N_5213,N_4213,N_4322);
nor U5214 (N_5214,N_2582,N_4596);
nand U5215 (N_5215,N_3644,N_3127);
or U5216 (N_5216,N_4139,N_4017);
nor U5217 (N_5217,N_3452,N_4400);
or U5218 (N_5218,N_3281,N_3547);
or U5219 (N_5219,N_3031,N_2593);
nor U5220 (N_5220,N_3606,N_4761);
nor U5221 (N_5221,N_4411,N_3161);
nand U5222 (N_5222,N_2729,N_3604);
and U5223 (N_5223,N_3845,N_2887);
nor U5224 (N_5224,N_3534,N_4150);
nor U5225 (N_5225,N_4320,N_4514);
nor U5226 (N_5226,N_4140,N_4218);
and U5227 (N_5227,N_3162,N_4610);
nand U5228 (N_5228,N_3591,N_2745);
and U5229 (N_5229,N_3444,N_3665);
and U5230 (N_5230,N_3277,N_3780);
nor U5231 (N_5231,N_3934,N_3245);
nor U5232 (N_5232,N_4983,N_4418);
nor U5233 (N_5233,N_3301,N_2773);
or U5234 (N_5234,N_4221,N_3569);
nor U5235 (N_5235,N_3238,N_3184);
and U5236 (N_5236,N_2544,N_3550);
nand U5237 (N_5237,N_2891,N_4007);
and U5238 (N_5238,N_2907,N_3694);
nor U5239 (N_5239,N_3731,N_4453);
and U5240 (N_5240,N_2683,N_4971);
and U5241 (N_5241,N_4084,N_4456);
or U5242 (N_5242,N_3270,N_2862);
or U5243 (N_5243,N_4928,N_3013);
or U5244 (N_5244,N_2661,N_4292);
or U5245 (N_5245,N_4326,N_3124);
or U5246 (N_5246,N_3435,N_3214);
nor U5247 (N_5247,N_3415,N_2949);
nand U5248 (N_5248,N_3895,N_3007);
and U5249 (N_5249,N_4458,N_3875);
nand U5250 (N_5250,N_3610,N_2563);
or U5251 (N_5251,N_4479,N_3297);
nand U5252 (N_5252,N_3414,N_2830);
and U5253 (N_5253,N_4708,N_3586);
nand U5254 (N_5254,N_3659,N_4351);
nand U5255 (N_5255,N_4580,N_3986);
nor U5256 (N_5256,N_3758,N_4274);
nor U5257 (N_5257,N_3608,N_3885);
and U5258 (N_5258,N_4957,N_3446);
nor U5259 (N_5259,N_4409,N_2641);
nor U5260 (N_5260,N_4918,N_2697);
and U5261 (N_5261,N_2921,N_4847);
or U5262 (N_5262,N_2849,N_2554);
nor U5263 (N_5263,N_4308,N_3976);
nand U5264 (N_5264,N_4327,N_4900);
and U5265 (N_5265,N_4564,N_4063);
or U5266 (N_5266,N_3048,N_3334);
nor U5267 (N_5267,N_4556,N_4890);
and U5268 (N_5268,N_3087,N_4369);
nand U5269 (N_5269,N_2507,N_2938);
and U5270 (N_5270,N_3437,N_2965);
or U5271 (N_5271,N_3037,N_3333);
nor U5272 (N_5272,N_4763,N_4554);
nand U5273 (N_5273,N_4388,N_4448);
and U5274 (N_5274,N_3693,N_3502);
or U5275 (N_5275,N_4743,N_3517);
or U5276 (N_5276,N_2910,N_3998);
nand U5277 (N_5277,N_4714,N_3669);
nor U5278 (N_5278,N_3180,N_3374);
nand U5279 (N_5279,N_4316,N_3860);
and U5280 (N_5280,N_2577,N_3894);
or U5281 (N_5281,N_2517,N_4857);
and U5282 (N_5282,N_3678,N_2784);
nand U5283 (N_5283,N_4417,N_3494);
and U5284 (N_5284,N_3965,N_4108);
and U5285 (N_5285,N_3054,N_3261);
and U5286 (N_5286,N_4966,N_3858);
nand U5287 (N_5287,N_3508,N_3442);
xor U5288 (N_5288,N_4430,N_2579);
xnor U5289 (N_5289,N_4099,N_2613);
nor U5290 (N_5290,N_4160,N_3292);
nor U5291 (N_5291,N_2501,N_2726);
nand U5292 (N_5292,N_4120,N_3079);
nand U5293 (N_5293,N_3525,N_3905);
and U5294 (N_5294,N_3373,N_2911);
nand U5295 (N_5295,N_2998,N_3671);
xor U5296 (N_5296,N_3592,N_2664);
nand U5297 (N_5297,N_4234,N_2894);
nor U5298 (N_5298,N_3393,N_2516);
nand U5299 (N_5299,N_3046,N_4709);
nand U5300 (N_5300,N_2728,N_4528);
and U5301 (N_5301,N_4517,N_2635);
nor U5302 (N_5302,N_3710,N_4981);
or U5303 (N_5303,N_3707,N_4078);
nor U5304 (N_5304,N_2779,N_4648);
or U5305 (N_5305,N_2603,N_3232);
or U5306 (N_5306,N_4522,N_4079);
and U5307 (N_5307,N_2599,N_4492);
nand U5308 (N_5308,N_4781,N_4085);
nand U5309 (N_5309,N_4166,N_3556);
nor U5310 (N_5310,N_4581,N_3368);
or U5311 (N_5311,N_3465,N_3101);
or U5312 (N_5312,N_3323,N_4622);
nand U5313 (N_5313,N_2798,N_2673);
or U5314 (N_5314,N_3518,N_4650);
and U5315 (N_5315,N_2590,N_3010);
and U5316 (N_5316,N_4591,N_4247);
and U5317 (N_5317,N_3419,N_3363);
or U5318 (N_5318,N_4695,N_4379);
and U5319 (N_5319,N_4116,N_3204);
nand U5320 (N_5320,N_4525,N_2580);
and U5321 (N_5321,N_2533,N_3540);
or U5322 (N_5322,N_4678,N_2962);
nand U5323 (N_5323,N_4549,N_4624);
and U5324 (N_5324,N_3417,N_2792);
nor U5325 (N_5325,N_4404,N_4716);
and U5326 (N_5326,N_4651,N_2569);
nor U5327 (N_5327,N_4513,N_4490);
xnor U5328 (N_5328,N_3717,N_3943);
nor U5329 (N_5329,N_3799,N_2968);
or U5330 (N_5330,N_3182,N_3008);
and U5331 (N_5331,N_4074,N_4721);
and U5332 (N_5332,N_3387,N_3543);
nand U5333 (N_5333,N_4035,N_3612);
and U5334 (N_5334,N_4906,N_3950);
and U5335 (N_5335,N_4179,N_4303);
nor U5336 (N_5336,N_4582,N_4909);
nand U5337 (N_5337,N_4186,N_3383);
nand U5338 (N_5338,N_2844,N_4866);
or U5339 (N_5339,N_2716,N_3134);
nor U5340 (N_5340,N_4253,N_3968);
nand U5341 (N_5341,N_2570,N_2768);
and U5342 (N_5342,N_2839,N_2955);
nand U5343 (N_5343,N_2600,N_4843);
or U5344 (N_5344,N_4987,N_2731);
nor U5345 (N_5345,N_3912,N_2588);
xor U5346 (N_5346,N_2617,N_4563);
xor U5347 (N_5347,N_2831,N_3774);
nand U5348 (N_5348,N_4432,N_3888);
nor U5349 (N_5349,N_4717,N_4032);
and U5350 (N_5350,N_4794,N_3170);
and U5351 (N_5351,N_2589,N_4362);
nor U5352 (N_5352,N_4955,N_4715);
or U5353 (N_5353,N_4088,N_3720);
nand U5354 (N_5354,N_2511,N_2742);
nor U5355 (N_5355,N_2997,N_3367);
or U5356 (N_5356,N_4538,N_2757);
or U5357 (N_5357,N_4686,N_2689);
or U5358 (N_5358,N_3926,N_3164);
nand U5359 (N_5359,N_3670,N_3552);
nor U5360 (N_5360,N_2988,N_2648);
and U5361 (N_5361,N_3741,N_3349);
and U5362 (N_5362,N_4602,N_2893);
or U5363 (N_5363,N_4305,N_2944);
xnor U5364 (N_5364,N_2693,N_4945);
nor U5365 (N_5365,N_4185,N_4661);
xor U5366 (N_5366,N_4839,N_3397);
nor U5367 (N_5367,N_2644,N_3344);
or U5368 (N_5368,N_3342,N_3189);
or U5369 (N_5369,N_3313,N_4476);
and U5370 (N_5370,N_4967,N_4641);
nand U5371 (N_5371,N_2707,N_3129);
and U5372 (N_5372,N_3100,N_2896);
nor U5373 (N_5373,N_3102,N_4092);
nor U5374 (N_5374,N_3259,N_4800);
or U5375 (N_5375,N_3685,N_4119);
nor U5376 (N_5376,N_4887,N_3190);
and U5377 (N_5377,N_3436,N_4765);
nor U5378 (N_5378,N_4259,N_3357);
nor U5379 (N_5379,N_3856,N_4629);
nand U5380 (N_5380,N_2979,N_3456);
nand U5381 (N_5381,N_4779,N_3132);
nand U5382 (N_5382,N_2609,N_4384);
and U5383 (N_5383,N_3406,N_3516);
nand U5384 (N_5384,N_4287,N_4509);
xor U5385 (N_5385,N_4683,N_4677);
and U5386 (N_5386,N_3389,N_4814);
nand U5387 (N_5387,N_4376,N_3967);
and U5388 (N_5388,N_3836,N_4117);
nand U5389 (N_5389,N_2913,N_4919);
or U5390 (N_5390,N_4357,N_3571);
and U5391 (N_5391,N_4364,N_3623);
nor U5392 (N_5392,N_3335,N_2677);
xnor U5393 (N_5393,N_4749,N_4389);
nand U5394 (N_5394,N_4552,N_4700);
nand U5395 (N_5395,N_3585,N_4129);
nand U5396 (N_5396,N_4336,N_2724);
nor U5397 (N_5397,N_3280,N_3135);
or U5398 (N_5398,N_2537,N_3689);
and U5399 (N_5399,N_3734,N_2640);
and U5400 (N_5400,N_3743,N_3382);
and U5401 (N_5401,N_3814,N_4450);
nand U5402 (N_5402,N_4868,N_2604);
nand U5403 (N_5403,N_4940,N_2895);
and U5404 (N_5404,N_3634,N_3773);
or U5405 (N_5405,N_3891,N_3580);
and U5406 (N_5406,N_2725,N_3058);
nand U5407 (N_5407,N_4862,N_4962);
nor U5408 (N_5408,N_3394,N_3366);
nand U5409 (N_5409,N_4876,N_4603);
and U5410 (N_5410,N_3911,N_2805);
nor U5411 (N_5411,N_4817,N_2523);
or U5412 (N_5412,N_3822,N_4026);
nand U5413 (N_5413,N_4811,N_3962);
nand U5414 (N_5414,N_4553,N_2933);
nand U5415 (N_5415,N_3354,N_4000);
nand U5416 (N_5416,N_4201,N_3255);
or U5417 (N_5417,N_2512,N_3169);
and U5418 (N_5418,N_3274,N_4408);
nor U5419 (N_5419,N_2951,N_3730);
or U5420 (N_5420,N_4220,N_4644);
and U5421 (N_5421,N_3513,N_4792);
xor U5422 (N_5422,N_4015,N_3370);
xnor U5423 (N_5423,N_4036,N_4860);
xnor U5424 (N_5424,N_4071,N_4758);
or U5425 (N_5425,N_4355,N_2627);
xor U5426 (N_5426,N_2663,N_2736);
or U5427 (N_5427,N_2859,N_3713);
nor U5428 (N_5428,N_2969,N_4943);
and U5429 (N_5429,N_2984,N_3109);
nand U5430 (N_5430,N_4865,N_4732);
and U5431 (N_5431,N_2616,N_4034);
or U5432 (N_5432,N_2900,N_3151);
or U5433 (N_5433,N_3412,N_4107);
and U5434 (N_5434,N_4009,N_4081);
nor U5435 (N_5435,N_4031,N_2954);
nand U5436 (N_5436,N_3812,N_2789);
and U5437 (N_5437,N_3613,N_3941);
or U5438 (N_5438,N_4976,N_4361);
and U5439 (N_5439,N_3464,N_3853);
and U5440 (N_5440,N_3044,N_3838);
nand U5441 (N_5441,N_3001,N_2654);
or U5442 (N_5442,N_2852,N_3343);
nand U5443 (N_5443,N_3661,N_4537);
or U5444 (N_5444,N_3183,N_3256);
or U5445 (N_5445,N_3826,N_3999);
and U5446 (N_5446,N_4601,N_4444);
nor U5447 (N_5447,N_4402,N_4130);
nand U5448 (N_5448,N_4193,N_4187);
nand U5449 (N_5449,N_4392,N_4874);
nand U5450 (N_5450,N_3902,N_4965);
and U5451 (N_5451,N_4054,N_4278);
nor U5452 (N_5452,N_4820,N_3656);
and U5453 (N_5453,N_3479,N_4737);
and U5454 (N_5454,N_3903,N_3047);
and U5455 (N_5455,N_3450,N_4852);
nor U5456 (N_5456,N_3246,N_3866);
or U5457 (N_5457,N_3461,N_3332);
nand U5458 (N_5458,N_4373,N_2630);
and U5459 (N_5459,N_3588,N_2973);
nand U5460 (N_5460,N_3431,N_3218);
and U5461 (N_5461,N_2514,N_2521);
nor U5462 (N_5462,N_3770,N_3003);
nand U5463 (N_5463,N_2860,N_4197);
nand U5464 (N_5464,N_3085,N_3199);
nand U5465 (N_5465,N_4589,N_2722);
or U5466 (N_5466,N_3023,N_4634);
or U5467 (N_5467,N_3545,N_2776);
nand U5468 (N_5468,N_3179,N_3823);
and U5469 (N_5469,N_3682,N_3409);
and U5470 (N_5470,N_4730,N_3113);
xor U5471 (N_5471,N_4263,N_2518);
nor U5472 (N_5472,N_4978,N_2733);
nor U5473 (N_5473,N_4970,N_3496);
and U5474 (N_5474,N_3195,N_2539);
nand U5475 (N_5475,N_4685,N_3692);
nor U5476 (N_5476,N_4338,N_2505);
and U5477 (N_5477,N_3544,N_3989);
nor U5478 (N_5478,N_2606,N_3015);
nand U5479 (N_5479,N_4861,N_4989);
nand U5480 (N_5480,N_3872,N_2562);
and U5481 (N_5481,N_3090,N_3136);
nor U5482 (N_5482,N_3611,N_4824);
and U5483 (N_5483,N_3067,N_3091);
or U5484 (N_5484,N_4101,N_4309);
or U5485 (N_5485,N_4859,N_3201);
or U5486 (N_5486,N_3961,N_3755);
and U5487 (N_5487,N_2918,N_3559);
and U5488 (N_5488,N_4387,N_3649);
nor U5489 (N_5489,N_4152,N_3573);
nand U5490 (N_5490,N_3081,N_4536);
and U5491 (N_5491,N_3587,N_4086);
or U5492 (N_5492,N_4975,N_4383);
nor U5493 (N_5493,N_2871,N_4854);
xor U5494 (N_5494,N_4102,N_3070);
or U5495 (N_5495,N_4358,N_3904);
or U5496 (N_5496,N_2818,N_2597);
and U5497 (N_5497,N_2740,N_4317);
and U5498 (N_5498,N_4626,N_4663);
or U5499 (N_5499,N_3012,N_3443);
and U5500 (N_5500,N_3336,N_2770);
nand U5501 (N_5501,N_4182,N_3798);
nand U5502 (N_5502,N_3648,N_4024);
and U5503 (N_5503,N_4719,N_3811);
and U5504 (N_5504,N_3491,N_2714);
or U5505 (N_5505,N_2625,N_3314);
nand U5506 (N_5506,N_3558,N_4627);
nor U5507 (N_5507,N_4572,N_3116);
xor U5508 (N_5508,N_4493,N_4982);
and U5509 (N_5509,N_2764,N_4673);
or U5510 (N_5510,N_4134,N_4046);
and U5511 (N_5511,N_4980,N_3679);
and U5512 (N_5512,N_4944,N_3438);
xor U5513 (N_5513,N_2550,N_3964);
xor U5514 (N_5514,N_3153,N_3566);
nand U5515 (N_5515,N_3757,N_4840);
or U5516 (N_5516,N_4368,N_4127);
nand U5517 (N_5517,N_2703,N_4964);
nor U5518 (N_5518,N_4751,N_4013);
or U5519 (N_5519,N_4920,N_4324);
nand U5520 (N_5520,N_4576,N_3876);
and U5521 (N_5521,N_4631,N_3772);
nand U5522 (N_5522,N_2975,N_4494);
and U5523 (N_5523,N_3563,N_4020);
and U5524 (N_5524,N_4830,N_3298);
nor U5525 (N_5525,N_3539,N_3681);
nand U5526 (N_5526,N_3732,N_3871);
nor U5527 (N_5527,N_3703,N_3581);
nor U5528 (N_5528,N_3381,N_3537);
and U5529 (N_5529,N_3938,N_2706);
nand U5530 (N_5530,N_4219,N_3123);
or U5531 (N_5531,N_3560,N_4922);
nor U5532 (N_5532,N_3695,N_4264);
and U5533 (N_5533,N_3924,N_2989);
nand U5534 (N_5534,N_3348,N_3922);
and U5535 (N_5535,N_2919,N_3192);
and U5536 (N_5536,N_3160,N_3990);
xnor U5537 (N_5537,N_3686,N_2986);
xnor U5538 (N_5538,N_4914,N_2585);
or U5539 (N_5539,N_4950,N_4497);
nor U5540 (N_5540,N_4642,N_3523);
or U5541 (N_5541,N_2581,N_2892);
nand U5542 (N_5542,N_2796,N_4053);
nor U5543 (N_5543,N_4199,N_3816);
nand U5544 (N_5544,N_3240,N_3021);
nor U5545 (N_5545,N_3844,N_4474);
nor U5546 (N_5546,N_3638,N_4726);
nand U5547 (N_5547,N_4002,N_4272);
and U5548 (N_5548,N_4649,N_3120);
nor U5549 (N_5549,N_3376,N_2564);
nand U5550 (N_5550,N_4475,N_4246);
or U5551 (N_5551,N_2845,N_4446);
nor U5552 (N_5552,N_3673,N_2686);
and U5553 (N_5553,N_2679,N_3841);
or U5554 (N_5554,N_4613,N_2734);
or U5555 (N_5555,N_2832,N_3933);
or U5556 (N_5556,N_4692,N_2901);
or U5557 (N_5557,N_4209,N_2869);
or U5558 (N_5558,N_4452,N_3078);
nor U5559 (N_5559,N_4917,N_3325);
or U5560 (N_5560,N_4516,N_3675);
nand U5561 (N_5561,N_2972,N_3759);
nand U5562 (N_5562,N_3421,N_3721);
nand U5563 (N_5563,N_4772,N_4097);
and U5564 (N_5564,N_4397,N_3782);
or U5565 (N_5565,N_4872,N_2513);
nor U5566 (N_5566,N_4289,N_3908);
and U5567 (N_5567,N_4654,N_4051);
xor U5568 (N_5568,N_3155,N_3206);
xor U5569 (N_5569,N_4027,N_2884);
nand U5570 (N_5570,N_3981,N_4321);
nor U5571 (N_5571,N_4385,N_4255);
or U5572 (N_5572,N_3809,N_3944);
and U5573 (N_5573,N_4774,N_3946);
nor U5574 (N_5574,N_4813,N_3535);
and U5575 (N_5575,N_3705,N_4921);
xor U5576 (N_5576,N_3122,N_3141);
nor U5577 (N_5577,N_4175,N_4330);
nand U5578 (N_5578,N_2886,N_4243);
and U5579 (N_5579,N_4997,N_4342);
or U5580 (N_5580,N_4615,N_2799);
or U5581 (N_5581,N_3016,N_4257);
nor U5582 (N_5582,N_3236,N_4323);
or U5583 (N_5583,N_3749,N_2598);
xor U5584 (N_5584,N_4510,N_4386);
and U5585 (N_5585,N_3227,N_4471);
or U5586 (N_5586,N_3052,N_4760);
nand U5587 (N_5587,N_3913,N_2929);
nand U5588 (N_5588,N_4062,N_2850);
nor U5589 (N_5589,N_3662,N_3859);
and U5590 (N_5590,N_3026,N_3379);
nand U5591 (N_5591,N_4607,N_4998);
and U5592 (N_5592,N_4467,N_3677);
nor U5593 (N_5593,N_3095,N_4815);
nand U5594 (N_5594,N_3618,N_3014);
nor U5595 (N_5595,N_3231,N_3089);
nand U5596 (N_5596,N_3060,N_4833);
nor U5597 (N_5597,N_3874,N_4896);
nor U5598 (N_5598,N_4232,N_4153);
or U5599 (N_5599,N_2974,N_3582);
nand U5600 (N_5600,N_3165,N_3704);
nor U5601 (N_5601,N_3355,N_4069);
and U5602 (N_5602,N_3804,N_3651);
and U5603 (N_5603,N_4435,N_3388);
nand U5604 (N_5604,N_3378,N_3119);
nand U5605 (N_5605,N_4786,N_3561);
nor U5606 (N_5606,N_4251,N_3072);
nor U5607 (N_5607,N_4873,N_4481);
xnor U5608 (N_5608,N_4170,N_3761);
xor U5609 (N_5609,N_4694,N_3305);
nand U5610 (N_5610,N_3094,N_3664);
and U5611 (N_5611,N_2692,N_4498);
or U5612 (N_5612,N_4584,N_4125);
xnor U5613 (N_5613,N_3785,N_3882);
xor U5614 (N_5614,N_3680,N_4331);
xor U5615 (N_5615,N_4194,N_4082);
nand U5616 (N_5616,N_4363,N_3805);
nand U5617 (N_5617,N_3993,N_3551);
nor U5618 (N_5618,N_4542,N_2735);
xnor U5619 (N_5619,N_3635,N_4241);
nor U5620 (N_5620,N_4339,N_3117);
xor U5621 (N_5621,N_4931,N_4795);
nand U5622 (N_5622,N_4003,N_4702);
or U5623 (N_5623,N_4671,N_3283);
nand U5624 (N_5624,N_2806,N_4592);
nor U5625 (N_5625,N_4895,N_3910);
and U5626 (N_5626,N_4994,N_3064);
and U5627 (N_5627,N_4070,N_4618);
or U5628 (N_5628,N_4472,N_3082);
and U5629 (N_5629,N_4740,N_3105);
or U5630 (N_5630,N_4770,N_4038);
nand U5631 (N_5631,N_3616,N_2906);
nand U5632 (N_5632,N_2819,N_3959);
nor U5633 (N_5633,N_3284,N_2671);
nand U5634 (N_5634,N_3837,N_3483);
and U5635 (N_5635,N_3898,N_2880);
nand U5636 (N_5636,N_4113,N_3320);
nand U5637 (N_5637,N_2650,N_3142);
or U5638 (N_5638,N_2957,N_3536);
nor U5639 (N_5639,N_3329,N_3807);
or U5640 (N_5640,N_3851,N_2565);
or U5641 (N_5641,N_4736,N_3765);
and U5642 (N_5642,N_3041,N_2552);
nor U5643 (N_5643,N_3622,N_2626);
or U5644 (N_5644,N_3130,N_3786);
nand U5645 (N_5645,N_4010,N_3131);
and U5646 (N_5646,N_4875,N_4343);
and U5647 (N_5647,N_4954,N_4148);
nand U5648 (N_5648,N_2701,N_2720);
nand U5649 (N_5649,N_4645,N_4356);
or U5650 (N_5650,N_4205,N_3156);
nand U5651 (N_5651,N_2822,N_2634);
and U5652 (N_5652,N_2780,N_2923);
xor U5653 (N_5653,N_3554,N_4281);
or U5654 (N_5654,N_4670,N_3602);
nand U5655 (N_5655,N_3795,N_3066);
or U5656 (N_5656,N_3645,N_4809);
nor U5657 (N_5657,N_2810,N_3803);
nor U5658 (N_5658,N_4635,N_2687);
and U5659 (N_5659,N_3029,N_3295);
nand U5660 (N_5660,N_4583,N_4750);
or U5661 (N_5661,N_4189,N_2527);
or U5662 (N_5662,N_4619,N_2756);
nand U5663 (N_5663,N_2875,N_2737);
xor U5664 (N_5664,N_4217,N_3784);
nor U5665 (N_5665,N_3215,N_3032);
or U5666 (N_5666,N_3341,N_4681);
and U5667 (N_5667,N_3568,N_3049);
nand U5668 (N_5668,N_4521,N_4952);
xor U5669 (N_5669,N_3800,N_3699);
or U5670 (N_5670,N_4604,N_4935);
xor U5671 (N_5671,N_2904,N_3764);
nor U5672 (N_5672,N_3402,N_3766);
or U5673 (N_5673,N_4061,N_2754);
and U5674 (N_5674,N_2956,N_4258);
nand U5675 (N_5675,N_4561,N_4999);
and U5676 (N_5676,N_3778,N_4159);
nand U5677 (N_5677,N_4718,N_4045);
nor U5678 (N_5678,N_4225,N_3080);
nor U5679 (N_5679,N_2947,N_4930);
or U5680 (N_5680,N_3235,N_4346);
xnor U5681 (N_5681,N_3043,N_4693);
nand U5682 (N_5682,N_4526,N_4137);
nor U5683 (N_5683,N_4350,N_3921);
nor U5684 (N_5684,N_3339,N_3207);
nand U5685 (N_5685,N_4459,N_3887);
or U5686 (N_5686,N_3919,N_4823);
and U5687 (N_5687,N_3209,N_3696);
and U5688 (N_5688,N_3470,N_2861);
and U5689 (N_5689,N_2867,N_4724);
nor U5690 (N_5690,N_2739,N_2642);
xnor U5691 (N_5691,N_3056,N_2926);
nand U5692 (N_5692,N_3392,N_3621);
and U5693 (N_5693,N_4850,N_3226);
and U5694 (N_5694,N_3099,N_4608);
nor U5695 (N_5695,N_4899,N_3951);
or U5696 (N_5696,N_4625,N_4881);
or U5697 (N_5697,N_4855,N_3260);
and U5698 (N_5698,N_2836,N_2842);
or U5699 (N_5699,N_2837,N_3752);
or U5700 (N_5700,N_4372,N_2567);
and U5701 (N_5701,N_3356,N_2548);
and U5702 (N_5702,N_4060,N_2816);
nand U5703 (N_5703,N_4687,N_3017);
or U5704 (N_5704,N_4742,N_4664);
and U5705 (N_5705,N_3760,N_4202);
nand U5706 (N_5706,N_2643,N_4226);
and U5707 (N_5707,N_2952,N_3973);
nand U5708 (N_5708,N_3053,N_4913);
or U5709 (N_5709,N_4806,N_3716);
or U5710 (N_5710,N_3247,N_4200);
nor U5711 (N_5711,N_2744,N_2990);
nor U5712 (N_5712,N_2838,N_3531);
nand U5713 (N_5713,N_4597,N_2995);
nor U5714 (N_5714,N_3506,N_3257);
nor U5715 (N_5715,N_4907,N_2638);
nor U5716 (N_5716,N_2963,N_2557);
or U5717 (N_5717,N_3627,N_2696);
nor U5718 (N_5718,N_4672,N_3762);
or U5719 (N_5719,N_3718,N_4969);
nor U5720 (N_5720,N_4731,N_4288);
nand U5721 (N_5721,N_4115,N_3626);
or U5722 (N_5722,N_4960,N_4300);
nand U5723 (N_5723,N_2759,N_4378);
and U5724 (N_5724,N_4095,N_3463);
nand U5725 (N_5725,N_3216,N_4039);
nand U5726 (N_5726,N_2583,N_4508);
and U5727 (N_5727,N_4043,N_3186);
nor U5728 (N_5728,N_2631,N_2898);
xnor U5729 (N_5729,N_4329,N_4429);
or U5730 (N_5730,N_3063,N_4745);
nor U5731 (N_5731,N_4279,N_4426);
or U5732 (N_5732,N_4238,N_3960);
or U5733 (N_5733,N_2717,N_3143);
nand U5734 (N_5734,N_4599,N_3427);
or U5735 (N_5735,N_3864,N_3055);
and U5736 (N_5736,N_4273,N_3712);
or U5737 (N_5737,N_4064,N_2835);
and U5738 (N_5738,N_3598,N_3906);
or U5739 (N_5739,N_4668,N_4974);
or U5740 (N_5740,N_4768,N_4523);
nor U5741 (N_5741,N_3865,N_4729);
nand U5742 (N_5742,N_2608,N_3213);
or U5743 (N_5743,N_3927,N_2812);
and U5744 (N_5744,N_3030,N_4856);
nand U5745 (N_5745,N_3490,N_4812);
nor U5746 (N_5746,N_4904,N_3737);
or U5747 (N_5747,N_4416,N_3738);
or U5748 (N_5748,N_2762,N_2821);
and U5749 (N_5749,N_3789,N_4478);
or U5750 (N_5750,N_3792,N_3018);
nor U5751 (N_5751,N_2755,N_3947);
nand U5752 (N_5752,N_2847,N_4611);
nor U5753 (N_5753,N_3299,N_3196);
and U5754 (N_5754,N_4019,N_2610);
and U5755 (N_5755,N_4680,N_4503);
and U5756 (N_5756,N_3620,N_4676);
nor U5757 (N_5757,N_3500,N_3522);
and U5758 (N_5758,N_2749,N_4254);
or U5759 (N_5759,N_4371,N_3273);
nor U5760 (N_5760,N_4703,N_3791);
and U5761 (N_5761,N_2758,N_2983);
and U5762 (N_5762,N_4885,N_3362);
or U5763 (N_5763,N_3181,N_2596);
nor U5764 (N_5764,N_3842,N_3279);
nand U5765 (N_5765,N_2851,N_3428);
or U5766 (N_5766,N_2685,N_4782);
nand U5767 (N_5767,N_4933,N_4953);
xnor U5768 (N_5768,N_3200,N_4889);
and U5769 (N_5769,N_2708,N_4395);
nor U5770 (N_5770,N_2618,N_4381);
or U5771 (N_5771,N_4437,N_2811);
and U5772 (N_5772,N_4778,N_2879);
nand U5773 (N_5773,N_3660,N_2652);
nor U5774 (N_5774,N_3744,N_4394);
xnor U5775 (N_5775,N_3953,N_3641);
and U5776 (N_5776,N_2743,N_3966);
or U5777 (N_5777,N_3173,N_4245);
nor U5778 (N_5778,N_4979,N_2876);
nand U5779 (N_5779,N_3351,N_4925);
xnor U5780 (N_5780,N_3915,N_3751);
and U5781 (N_5781,N_3211,N_4710);
nor U5782 (N_5782,N_4136,N_3977);
nor U5783 (N_5783,N_3077,N_2559);
nand U5784 (N_5784,N_4577,N_4041);
nand U5785 (N_5785,N_4306,N_4666);
nand U5786 (N_5786,N_2790,N_2510);
or U5787 (N_5787,N_2827,N_3278);
nand U5788 (N_5788,N_3275,N_4573);
or U5789 (N_5789,N_3956,N_3840);
nor U5790 (N_5790,N_4689,N_4168);
xnor U5791 (N_5791,N_3601,N_3530);
or U5792 (N_5792,N_4539,N_2715);
or U5793 (N_5793,N_4696,N_4271);
and U5794 (N_5794,N_4065,N_3630);
or U5795 (N_5795,N_3969,N_3972);
or U5796 (N_5796,N_3493,N_3068);
nand U5797 (N_5797,N_3039,N_3107);
nor U5798 (N_5798,N_4762,N_4669);
nand U5799 (N_5799,N_4704,N_3489);
xnor U5800 (N_5800,N_3958,N_4008);
or U5801 (N_5801,N_3521,N_4886);
xor U5802 (N_5802,N_4545,N_3439);
xor U5803 (N_5803,N_4728,N_4805);
or U5804 (N_5804,N_3249,N_3702);
nand U5805 (N_5805,N_4110,N_4942);
nor U5806 (N_5806,N_3369,N_4558);
or U5807 (N_5807,N_4441,N_3481);
nor U5808 (N_5808,N_2615,N_2710);
or U5809 (N_5809,N_3579,N_2748);
nor U5810 (N_5810,N_3572,N_2787);
and U5811 (N_5811,N_2719,N_4752);
nand U5812 (N_5812,N_4986,N_4638);
and U5813 (N_5813,N_4463,N_3250);
nor U5814 (N_5814,N_3198,N_3631);
or U5815 (N_5815,N_4505,N_2684);
xor U5816 (N_5816,N_4616,N_4759);
or U5817 (N_5817,N_3158,N_4804);
xor U5818 (N_5818,N_4797,N_3917);
xnor U5819 (N_5819,N_3609,N_3884);
or U5820 (N_5820,N_3219,N_3168);
and U5821 (N_5821,N_3174,N_3935);
nor U5822 (N_5822,N_4261,N_2829);
nand U5823 (N_5823,N_4044,N_3570);
nand U5824 (N_5824,N_3484,N_4164);
xnor U5825 (N_5825,N_3000,N_4311);
nand U5826 (N_5826,N_2591,N_4482);
nand U5827 (N_5827,N_3690,N_3340);
nor U5828 (N_5828,N_3783,N_3555);
xnor U5829 (N_5829,N_4500,N_3308);
and U5830 (N_5830,N_2942,N_3879);
xor U5831 (N_5831,N_4636,N_4405);
nand U5832 (N_5832,N_3197,N_4502);
xor U5833 (N_5833,N_4293,N_3529);
or U5834 (N_5834,N_3287,N_4210);
nand U5835 (N_5835,N_3519,N_4802);
nor U5836 (N_5836,N_4963,N_2788);
nor U5837 (N_5837,N_3413,N_2682);
xor U5838 (N_5838,N_4068,N_2765);
or U5839 (N_5839,N_3040,N_4005);
nand U5840 (N_5840,N_3042,N_4442);
nand U5841 (N_5841,N_2813,N_3567);
nand U5842 (N_5842,N_4114,N_3781);
nor U5843 (N_5843,N_4023,N_4016);
nor U5844 (N_5844,N_4819,N_2905);
xor U5845 (N_5845,N_4021,N_3138);
xor U5846 (N_5846,N_4177,N_4295);
and U5847 (N_5847,N_4977,N_4307);
nor U5848 (N_5848,N_4310,N_4425);
nor U5849 (N_5849,N_3652,N_3286);
or U5850 (N_5850,N_3264,N_3317);
or U5851 (N_5851,N_3639,N_4785);
and U5852 (N_5852,N_4653,N_3715);
and U5853 (N_5853,N_2611,N_3477);
or U5854 (N_5854,N_4353,N_2614);
or U5855 (N_5855,N_2857,N_4296);
and U5856 (N_5856,N_4354,N_4623);
and U5857 (N_5857,N_3745,N_2945);
nand U5858 (N_5858,N_4480,N_4230);
or U5859 (N_5859,N_2556,N_3108);
or U5860 (N_5860,N_4421,N_2675);
nor U5861 (N_5861,N_2712,N_2878);
xor U5862 (N_5862,N_3258,N_2702);
or U5863 (N_5863,N_4491,N_3658);
and U5864 (N_5864,N_4688,N_4707);
nor U5865 (N_5865,N_2970,N_3982);
and U5866 (N_5866,N_4555,N_2730);
or U5867 (N_5867,N_4570,N_3501);
and U5868 (N_5868,N_2777,N_4132);
or U5869 (N_5869,N_4882,N_4211);
xor U5870 (N_5870,N_4018,N_3083);
xnor U5871 (N_5871,N_4698,N_3149);
xnor U5872 (N_5872,N_4319,N_4801);
nand U5873 (N_5873,N_3936,N_4192);
or U5874 (N_5874,N_4934,N_4469);
nand U5875 (N_5875,N_4398,N_3426);
or U5876 (N_5876,N_3111,N_3361);
or U5877 (N_5877,N_2619,N_3288);
or U5878 (N_5878,N_4880,N_4844);
and U5879 (N_5879,N_3847,N_3148);
or U5880 (N_5880,N_2760,N_2772);
nand U5881 (N_5881,N_4853,N_3460);
or U5882 (N_5882,N_3372,N_3033);
nor U5883 (N_5883,N_4937,N_4640);
xor U5884 (N_5884,N_4665,N_4727);
nand U5885 (N_5885,N_2656,N_4941);
nor U5886 (N_5886,N_3449,N_3843);
and U5887 (N_5887,N_3869,N_4370);
and U5888 (N_5888,N_4574,N_2766);
xnor U5889 (N_5889,N_4093,N_2961);
nor U5890 (N_5890,N_4748,N_3319);
nand U5891 (N_5891,N_3808,N_4033);
xor U5892 (N_5892,N_3952,N_3603);
and U5893 (N_5893,N_4739,N_4285);
and U5894 (N_5894,N_4546,N_4375);
nor U5895 (N_5895,N_4878,N_2870);
or U5896 (N_5896,N_3834,N_2825);
nand U5897 (N_5897,N_2980,N_2658);
and U5898 (N_5898,N_2877,N_4990);
xor U5899 (N_5899,N_3701,N_4109);
or U5900 (N_5900,N_4675,N_4594);
nor U5901 (N_5901,N_4808,N_4519);
xnor U5902 (N_5902,N_3593,N_4793);
or U5903 (N_5903,N_4112,N_2529);
nand U5904 (N_5904,N_3565,N_4470);
or U5905 (N_5905,N_3251,N_4484);
and U5906 (N_5906,N_4449,N_3440);
or U5907 (N_5907,N_4846,N_3578);
xor U5908 (N_5908,N_4511,N_2978);
nand U5909 (N_5909,N_3262,N_2709);
xnor U5910 (N_5910,N_4204,N_4367);
nand U5911 (N_5911,N_2865,N_4284);
and U5912 (N_5912,N_3533,N_4301);
nor U5913 (N_5913,N_2620,N_4851);
and U5914 (N_5914,N_3668,N_4838);
nor U5915 (N_5915,N_4058,N_4131);
nor U5916 (N_5916,N_2595,N_4298);
or U5917 (N_5917,N_4684,N_2695);
nor U5918 (N_5918,N_2991,N_2568);
nand U5919 (N_5919,N_3756,N_4845);
or U5920 (N_5920,N_4333,N_4056);
xor U5921 (N_5921,N_4335,N_3553);
and U5922 (N_5922,N_2946,N_3787);
and U5923 (N_5923,N_3172,N_4180);
xnor U5924 (N_5924,N_2628,N_4420);
nor U5925 (N_5925,N_3771,N_2763);
nor U5926 (N_5926,N_4701,N_3422);
nand U5927 (N_5927,N_3005,N_2774);
nor U5928 (N_5928,N_3405,N_4240);
nor U5929 (N_5929,N_2841,N_4011);
and U5930 (N_5930,N_3683,N_4787);
or U5931 (N_5931,N_3234,N_4422);
nand U5932 (N_5932,N_4014,N_4181);
or U5933 (N_5933,N_3714,N_2888);
or U5934 (N_5934,N_3071,N_4104);
and U5935 (N_5935,N_3103,N_3110);
nor U5936 (N_5936,N_3832,N_3526);
xor U5937 (N_5937,N_2649,N_4863);
and U5938 (N_5938,N_4557,N_3979);
or U5939 (N_5939,N_3557,N_4439);
xnor U5940 (N_5940,N_3328,N_2601);
xnor U5941 (N_5941,N_3019,N_4419);
nor U5942 (N_5942,N_4460,N_4834);
xor U5943 (N_5943,N_4956,N_4524);
nand U5944 (N_5944,N_3290,N_4312);
nor U5945 (N_5945,N_4096,N_4620);
nor U5946 (N_5946,N_3996,N_3499);
xnor U5947 (N_5947,N_3411,N_3324);
nor U5948 (N_5948,N_3121,N_3294);
or U5949 (N_5949,N_4741,N_3624);
nand U5950 (N_5950,N_2558,N_4059);
nand U5951 (N_5951,N_3867,N_2573);
and U5952 (N_5952,N_4864,N_4807);
and U5953 (N_5953,N_3880,N_3599);
nand U5954 (N_5954,N_2612,N_2665);
or U5955 (N_5955,N_4135,N_3404);
and U5956 (N_5956,N_4789,N_4568);
nand U5957 (N_5957,N_3025,N_4156);
xor U5958 (N_5958,N_2605,N_3453);
and U5959 (N_5959,N_2794,N_4037);
and U5960 (N_5960,N_4771,N_3821);
nor U5961 (N_5961,N_4947,N_3930);
and U5962 (N_5962,N_3159,N_4144);
and U5963 (N_5963,N_4891,N_3727);
or U5964 (N_5964,N_2817,N_4440);
and U5965 (N_5965,N_3364,N_2647);
and U5966 (N_5966,N_4936,N_3617);
nor U5967 (N_5967,N_3144,N_4231);
xor U5968 (N_5968,N_2856,N_3241);
xor U5969 (N_5969,N_3128,N_4527);
or U5970 (N_5970,N_3244,N_4393);
xor U5971 (N_5971,N_3514,N_3788);
nor U5972 (N_5972,N_4946,N_3312);
or U5973 (N_5973,N_3646,N_4722);
and U5974 (N_5974,N_3271,N_4662);
nand U5975 (N_5975,N_2653,N_4884);
nand U5976 (N_5976,N_3050,N_4178);
or U5977 (N_5977,N_3779,N_2532);
or U5978 (N_5978,N_2964,N_3748);
or U5979 (N_5979,N_3027,N_3655);
nor U5980 (N_5980,N_3210,N_4124);
nand U5981 (N_5981,N_4275,N_4042);
and U5982 (N_5982,N_4848,N_3360);
and U5983 (N_5983,N_4643,N_2840);
nand U5984 (N_5984,N_4083,N_2824);
nor U5985 (N_5985,N_3445,N_2881);
or U5986 (N_5986,N_3600,N_3482);
or U5987 (N_5987,N_2807,N_3886);
nor U5988 (N_5988,N_4911,N_3576);
or U5989 (N_5989,N_3820,N_3118);
nand U5990 (N_5990,N_3980,N_4294);
and U5991 (N_5991,N_3221,N_4984);
xnor U5992 (N_5992,N_3220,N_4652);
or U5993 (N_5993,N_3667,N_4457);
and U5994 (N_5994,N_4249,N_3088);
nor U5995 (N_5995,N_4466,N_4587);
nand U5996 (N_5996,N_3248,N_3505);
or U5997 (N_5997,N_3633,N_2660);
and U5998 (N_5998,N_3242,N_3992);
and U5999 (N_5999,N_3733,N_4832);
nand U6000 (N_6000,N_2993,N_4464);
nand U6001 (N_6001,N_3086,N_2704);
or U6002 (N_6002,N_4870,N_3125);
and U6003 (N_6003,N_4162,N_3469);
xor U6004 (N_6004,N_4030,N_3115);
nand U6005 (N_6005,N_2753,N_2711);
nand U6006 (N_6006,N_3178,N_3916);
and U6007 (N_6007,N_4206,N_3455);
or U6008 (N_6008,N_4268,N_3831);
nand U6009 (N_6009,N_3347,N_4905);
or U6010 (N_6010,N_3065,N_4682);
nor U6011 (N_6011,N_3024,N_4090);
or U6012 (N_6012,N_4138,N_4747);
xor U6013 (N_6013,N_2937,N_3984);
xor U6014 (N_6014,N_3408,N_3321);
nor U6015 (N_6015,N_3300,N_2646);
or U6016 (N_6016,N_3643,N_3767);
and U6017 (N_6017,N_4775,N_3945);
and U6018 (N_6018,N_4548,N_3152);
nor U6019 (N_6019,N_3819,N_3995);
or U6020 (N_6020,N_2629,N_3650);
or U6021 (N_6021,N_3410,N_4477);
or U6022 (N_6022,N_4012,N_4533);
xnor U6023 (N_6023,N_4040,N_2939);
and U6024 (N_6024,N_2718,N_3486);
nor U6025 (N_6025,N_4614,N_3509);
nor U6026 (N_6026,N_4892,N_2637);
or U6027 (N_6027,N_2540,N_4366);
nor U6028 (N_6028,N_3596,N_4547);
xnor U6029 (N_6029,N_3849,N_4157);
or U6030 (N_6030,N_3276,N_3802);
nor U6031 (N_6031,N_2574,N_4436);
nor U6032 (N_6032,N_4562,N_3114);
nand U6033 (N_6033,N_3187,N_4705);
or U6034 (N_6034,N_3188,N_3139);
and U6035 (N_6035,N_4633,N_4315);
or U6036 (N_6036,N_2803,N_3931);
or U6037 (N_6037,N_3338,N_2943);
or U6038 (N_6038,N_4972,N_2883);
xor U6039 (N_6039,N_3697,N_3473);
nor U6040 (N_6040,N_3932,N_4995);
or U6041 (N_6041,N_4145,N_3488);
and U6042 (N_6042,N_3006,N_4897);
xor U6043 (N_6043,N_3777,N_4566);
or U6044 (N_6044,N_3311,N_3801);
and U6045 (N_6045,N_3337,N_4567);
nand U6046 (N_6046,N_3584,N_2783);
and U6047 (N_6047,N_4347,N_3310);
or U6048 (N_6048,N_4414,N_4133);
or U6049 (N_6049,N_4822,N_4184);
nor U6050 (N_6050,N_2542,N_3429);
nor U6051 (N_6051,N_3846,N_3073);
nor U6052 (N_6052,N_3769,N_4630);
nand U6053 (N_6053,N_2651,N_4100);
and U6054 (N_6054,N_3092,N_4345);
and U6055 (N_6055,N_4501,N_2572);
or U6056 (N_6056,N_3472,N_2678);
nor U6057 (N_6057,N_4600,N_2866);
or U6058 (N_6058,N_3289,N_2506);
nand U6059 (N_6059,N_4262,N_4183);
and U6060 (N_6060,N_4816,N_2922);
and U6061 (N_6061,N_2890,N_4968);
or U6062 (N_6062,N_4985,N_4434);
nor U6063 (N_6063,N_2667,N_4337);
xnor U6064 (N_6064,N_2578,N_4413);
or U6065 (N_6065,N_3753,N_3899);
and U6066 (N_6066,N_2795,N_4266);
nor U6067 (N_6067,N_4344,N_3527);
and U6068 (N_6068,N_4780,N_3729);
xnor U6069 (N_6069,N_4504,N_3928);
nand U6070 (N_6070,N_3424,N_4790);
and U6071 (N_6071,N_3512,N_4674);
nor U6072 (N_6072,N_4066,N_4571);
nand U6073 (N_6073,N_3815,N_3520);
and U6074 (N_6074,N_4406,N_3454);
and U6075 (N_6075,N_4776,N_4198);
and U6076 (N_6076,N_2575,N_4541);
and U6077 (N_6077,N_2931,N_4810);
xnor U6078 (N_6078,N_4250,N_4252);
xor U6079 (N_6079,N_4550,N_3327);
and U6080 (N_6080,N_3167,N_2801);
nor U6081 (N_6081,N_4290,N_2502);
nand U6082 (N_6082,N_3607,N_4228);
nor U6083 (N_6083,N_4239,N_4057);
or U6084 (N_6084,N_3476,N_4991);
nor U6085 (N_6085,N_3719,N_4888);
and U6086 (N_6086,N_4483,N_2934);
xor U6087 (N_6087,N_2688,N_3987);
and U6088 (N_6088,N_4518,N_3466);
or U6089 (N_6089,N_4869,N_3735);
or U6090 (N_6090,N_2732,N_3901);
or U6091 (N_6091,N_4260,N_3345);
or U6092 (N_6092,N_2555,N_4143);
xor U6093 (N_6093,N_2503,N_4077);
or U6094 (N_6094,N_3233,N_4236);
and U6095 (N_6095,N_4396,N_4512);
nor U6096 (N_6096,N_3708,N_4783);
nor U6097 (N_6097,N_3243,N_2560);
nand U6098 (N_6098,N_3309,N_3059);
nor U6099 (N_6099,N_4075,N_3485);
nand U6100 (N_6100,N_4267,N_4915);
nand U6101 (N_6101,N_2691,N_3035);
nor U6102 (N_6102,N_4893,N_3069);
or U6103 (N_6103,N_3524,N_4699);
and U6104 (N_6104,N_4067,N_4612);
nand U6105 (N_6105,N_3154,N_3254);
nand U6106 (N_6106,N_4495,N_4118);
and U6107 (N_6107,N_3475,N_3949);
nand U6108 (N_6108,N_3407,N_3829);
nand U6109 (N_6109,N_3742,N_4706);
or U6110 (N_6110,N_4277,N_4190);
or U6111 (N_6111,N_3315,N_2967);
and U6112 (N_6112,N_2826,N_4025);
nand U6113 (N_6113,N_3202,N_2549);
nor U6114 (N_6114,N_4828,N_4216);
nor U6115 (N_6115,N_4172,N_3589);
xnor U6116 (N_6116,N_4713,N_4506);
or U6117 (N_6117,N_2767,N_3296);
and U6118 (N_6118,N_4123,N_3575);
and U6119 (N_6119,N_2690,N_3542);
or U6120 (N_6120,N_3909,N_4628);
and U6121 (N_6121,N_4171,N_4826);
nand U6122 (N_6122,N_4462,N_2694);
or U6123 (N_6123,N_3147,N_4690);
nand U6124 (N_6124,N_3827,N_3963);
or U6125 (N_6125,N_3722,N_4349);
and U6126 (N_6126,N_3813,N_4605);
or U6127 (N_6127,N_4996,N_3900);
nor U6128 (N_6128,N_4154,N_4754);
nand U6129 (N_6129,N_4902,N_4496);
nor U6130 (N_6130,N_3881,N_2674);
or U6131 (N_6131,N_4829,N_3358);
and U6132 (N_6132,N_3810,N_4711);
xor U6133 (N_6133,N_4149,N_4188);
nor U6134 (N_6134,N_3740,N_3614);
and U6135 (N_6135,N_3403,N_2721);
or U6136 (N_6136,N_4632,N_3293);
nand U6137 (N_6137,N_4203,N_3487);
xor U6138 (N_6138,N_4821,N_4487);
or U6139 (N_6139,N_2546,N_2520);
nand U6140 (N_6140,N_3390,N_3739);
and U6141 (N_6141,N_3868,N_2526);
and U6142 (N_6142,N_4121,N_2769);
nor U6143 (N_6143,N_4105,N_4927);
nor U6144 (N_6144,N_2908,N_4242);
and U6145 (N_6145,N_3726,N_3272);
nor U6146 (N_6146,N_4579,N_3723);
xor U6147 (N_6147,N_3985,N_2681);
nand U6148 (N_6148,N_4598,N_3861);
nor U6149 (N_6149,N_2750,N_4455);
xnor U6150 (N_6150,N_4158,N_4588);
or U6151 (N_6151,N_4382,N_3457);
nor U6152 (N_6152,N_3794,N_4403);
nor U6153 (N_6153,N_4679,N_4520);
or U6154 (N_6154,N_3728,N_4229);
xnor U6155 (N_6155,N_2981,N_3628);
and U6156 (N_6156,N_3654,N_4080);
or U6157 (N_6157,N_3028,N_3266);
and U6158 (N_6158,N_4399,N_2994);
and U6159 (N_6159,N_3126,N_4048);
or U6160 (N_6160,N_2925,N_3776);
nor U6161 (N_6161,N_4314,N_4445);
nand U6162 (N_6162,N_3818,N_3175);
nand U6163 (N_6163,N_2713,N_4055);
nand U6164 (N_6164,N_3253,N_4530);
xnor U6165 (N_6165,N_4764,N_3423);
and U6166 (N_6166,N_4757,N_4423);
nand U6167 (N_6167,N_4412,N_3892);
nand U6168 (N_6168,N_3004,N_3955);
nand U6169 (N_6169,N_3020,N_2940);
nor U6170 (N_6170,N_3750,N_3615);
and U6171 (N_6171,N_4769,N_3763);
and U6172 (N_6172,N_4489,N_2747);
nor U6173 (N_6173,N_3852,N_4773);
xnor U6174 (N_6174,N_3480,N_3163);
and U6175 (N_6175,N_4733,N_3883);
xor U6176 (N_6176,N_2504,N_2746);
and U6177 (N_6177,N_4575,N_3975);
nand U6178 (N_6178,N_4803,N_3458);
nor U6179 (N_6179,N_3022,N_4352);
and U6180 (N_6180,N_2752,N_3855);
nand U6181 (N_6181,N_3674,N_2953);
and U6182 (N_6182,N_4609,N_4438);
and U6183 (N_6183,N_2524,N_2924);
and U6184 (N_6184,N_3971,N_3492);
nand U6185 (N_6185,N_3507,N_4590);
nand U6186 (N_6186,N_4894,N_3988);
nor U6187 (N_6187,N_3441,N_2534);
or U6188 (N_6188,N_3497,N_2592);
or U6189 (N_6189,N_3377,N_3957);
nor U6190 (N_6190,N_2800,N_3451);
and U6191 (N_6191,N_2543,N_4559);
and U6192 (N_6192,N_4468,N_4767);
nor U6193 (N_6193,N_2864,N_4637);
nand U6194 (N_6194,N_3824,N_3504);
or U6195 (N_6195,N_4593,N_4660);
and U6196 (N_6196,N_4325,N_2950);
nor U6197 (N_6197,N_4734,N_2793);
nand U6198 (N_6198,N_2853,N_3265);
and U6199 (N_6199,N_3889,N_4122);
and U6200 (N_6200,N_4196,N_3061);
xnor U6201 (N_6201,N_4161,N_3185);
and U6202 (N_6202,N_3106,N_2566);
nor U6203 (N_6203,N_2508,N_4738);
or U6204 (N_6204,N_4723,N_2797);
and U6205 (N_6205,N_2576,N_3166);
and U6206 (N_6206,N_3594,N_4248);
xnor U6207 (N_6207,N_3252,N_3625);
or U6208 (N_6208,N_4923,N_4871);
nor U6209 (N_6209,N_2668,N_2741);
and U6210 (N_6210,N_3538,N_4961);
xnor U6211 (N_6211,N_2814,N_4621);
or U6212 (N_6212,N_2941,N_2999);
nor U6213 (N_6213,N_3237,N_4451);
nand U6214 (N_6214,N_3736,N_3467);
nor U6215 (N_6215,N_3075,N_2889);
and U6216 (N_6216,N_4318,N_2833);
nand U6217 (N_6217,N_4365,N_3176);
and U6218 (N_6218,N_2659,N_4543);
and U6219 (N_6219,N_2525,N_3285);
nand U6220 (N_6220,N_2785,N_3896);
nor U6221 (N_6221,N_3096,N_4958);
and U6222 (N_6222,N_4223,N_4784);
and U6223 (N_6223,N_4276,N_3398);
nand U6224 (N_6224,N_4155,N_3353);
nand U6225 (N_6225,N_3914,N_3038);
nand U6226 (N_6226,N_4214,N_2874);
and U6227 (N_6227,N_3511,N_4332);
xnor U6228 (N_6228,N_2515,N_3642);
xnor U6229 (N_6229,N_4993,N_4212);
and U6230 (N_6230,N_3036,N_2804);
nor U6231 (N_6231,N_2872,N_2903);
nand U6232 (N_6232,N_3954,N_3420);
nor U6233 (N_6233,N_4098,N_3970);
xnor U6234 (N_6234,N_3400,N_4515);
or U6235 (N_6235,N_4073,N_4282);
nor U6236 (N_6236,N_4447,N_2971);
nor U6237 (N_6237,N_4235,N_4473);
nand U6238 (N_6238,N_2802,N_4659);
or U6239 (N_6239,N_4237,N_2551);
or U6240 (N_6240,N_4244,N_3640);
nand U6241 (N_6241,N_3194,N_3709);
nor U6242 (N_6242,N_2977,N_4753);
or U6243 (N_6243,N_2976,N_3225);
or U6244 (N_6244,N_3929,N_3228);
and U6245 (N_6245,N_4791,N_4835);
nand U6246 (N_6246,N_3171,N_4531);
or U6247 (N_6247,N_2698,N_3191);
nor U6248 (N_6248,N_4390,N_2561);
xnor U6249 (N_6249,N_3097,N_2771);
nor U6250 (N_6250,N_3710,N_4193);
nor U6251 (N_6251,N_2834,N_4900);
nand U6252 (N_6252,N_4541,N_3698);
nand U6253 (N_6253,N_4596,N_3839);
and U6254 (N_6254,N_4521,N_3881);
xnor U6255 (N_6255,N_4273,N_3968);
or U6256 (N_6256,N_4975,N_2668);
and U6257 (N_6257,N_3264,N_4703);
and U6258 (N_6258,N_2998,N_2736);
and U6259 (N_6259,N_4261,N_4918);
xor U6260 (N_6260,N_4289,N_3521);
nand U6261 (N_6261,N_3180,N_4651);
xor U6262 (N_6262,N_4666,N_2942);
nand U6263 (N_6263,N_4885,N_2970);
nand U6264 (N_6264,N_3216,N_4050);
or U6265 (N_6265,N_3673,N_3840);
nor U6266 (N_6266,N_4456,N_3460);
or U6267 (N_6267,N_2904,N_4804);
or U6268 (N_6268,N_2710,N_4985);
xnor U6269 (N_6269,N_4537,N_4637);
and U6270 (N_6270,N_4941,N_3868);
nand U6271 (N_6271,N_2903,N_4584);
or U6272 (N_6272,N_2947,N_4589);
nor U6273 (N_6273,N_4299,N_4564);
nand U6274 (N_6274,N_4925,N_4429);
nand U6275 (N_6275,N_4404,N_2654);
xor U6276 (N_6276,N_3958,N_4588);
and U6277 (N_6277,N_2914,N_4452);
nand U6278 (N_6278,N_3381,N_3600);
or U6279 (N_6279,N_3524,N_4850);
xnor U6280 (N_6280,N_4828,N_4996);
and U6281 (N_6281,N_2986,N_3643);
xnor U6282 (N_6282,N_3662,N_3119);
nor U6283 (N_6283,N_3494,N_4233);
and U6284 (N_6284,N_3163,N_4618);
and U6285 (N_6285,N_3131,N_2617);
nor U6286 (N_6286,N_3951,N_3783);
nand U6287 (N_6287,N_3894,N_4486);
nor U6288 (N_6288,N_3991,N_3338);
and U6289 (N_6289,N_3062,N_3291);
or U6290 (N_6290,N_4663,N_4538);
or U6291 (N_6291,N_3681,N_3669);
nor U6292 (N_6292,N_2900,N_2857);
xor U6293 (N_6293,N_3875,N_4857);
or U6294 (N_6294,N_2634,N_4536);
and U6295 (N_6295,N_4452,N_2597);
and U6296 (N_6296,N_4214,N_2528);
nor U6297 (N_6297,N_3567,N_4846);
nand U6298 (N_6298,N_2856,N_3134);
xor U6299 (N_6299,N_4058,N_4172);
and U6300 (N_6300,N_4245,N_3109);
nand U6301 (N_6301,N_4285,N_4031);
or U6302 (N_6302,N_2623,N_2503);
or U6303 (N_6303,N_3286,N_3624);
nand U6304 (N_6304,N_3843,N_4211);
and U6305 (N_6305,N_4466,N_2503);
and U6306 (N_6306,N_3778,N_3602);
nor U6307 (N_6307,N_3630,N_3593);
nor U6308 (N_6308,N_4095,N_2958);
nor U6309 (N_6309,N_4915,N_3357);
nor U6310 (N_6310,N_4125,N_3221);
nand U6311 (N_6311,N_4946,N_4963);
nand U6312 (N_6312,N_2665,N_3608);
nor U6313 (N_6313,N_4625,N_4603);
nor U6314 (N_6314,N_3486,N_2581);
nand U6315 (N_6315,N_3433,N_4478);
and U6316 (N_6316,N_4798,N_3039);
nand U6317 (N_6317,N_4250,N_3889);
nand U6318 (N_6318,N_4684,N_3674);
or U6319 (N_6319,N_4992,N_3049);
nand U6320 (N_6320,N_2526,N_3419);
nor U6321 (N_6321,N_2745,N_2958);
or U6322 (N_6322,N_3137,N_2516);
nor U6323 (N_6323,N_3736,N_3023);
nand U6324 (N_6324,N_4911,N_3472);
or U6325 (N_6325,N_4995,N_3189);
nand U6326 (N_6326,N_4544,N_3008);
nand U6327 (N_6327,N_4322,N_3930);
nand U6328 (N_6328,N_4424,N_3317);
and U6329 (N_6329,N_4097,N_4575);
nand U6330 (N_6330,N_4427,N_3005);
and U6331 (N_6331,N_4808,N_4440);
and U6332 (N_6332,N_4384,N_4578);
and U6333 (N_6333,N_4562,N_3622);
and U6334 (N_6334,N_2574,N_2892);
and U6335 (N_6335,N_3111,N_3285);
or U6336 (N_6336,N_4338,N_4534);
nor U6337 (N_6337,N_3484,N_3632);
nand U6338 (N_6338,N_4412,N_4863);
nand U6339 (N_6339,N_4853,N_3232);
and U6340 (N_6340,N_3912,N_3467);
and U6341 (N_6341,N_3016,N_2553);
or U6342 (N_6342,N_4126,N_3677);
or U6343 (N_6343,N_3546,N_2906);
nand U6344 (N_6344,N_3213,N_3800);
nor U6345 (N_6345,N_3414,N_3371);
or U6346 (N_6346,N_3657,N_3728);
nor U6347 (N_6347,N_4928,N_4835);
xnor U6348 (N_6348,N_3735,N_3497);
nor U6349 (N_6349,N_3976,N_3300);
nor U6350 (N_6350,N_4504,N_4406);
and U6351 (N_6351,N_2638,N_4362);
nand U6352 (N_6352,N_3187,N_4751);
xor U6353 (N_6353,N_4156,N_4030);
or U6354 (N_6354,N_4987,N_4715);
and U6355 (N_6355,N_4495,N_3113);
or U6356 (N_6356,N_3422,N_4708);
or U6357 (N_6357,N_3425,N_3550);
or U6358 (N_6358,N_3897,N_3831);
or U6359 (N_6359,N_4679,N_4856);
and U6360 (N_6360,N_4767,N_3612);
nor U6361 (N_6361,N_4069,N_3366);
and U6362 (N_6362,N_2769,N_4461);
nor U6363 (N_6363,N_4767,N_4512);
nand U6364 (N_6364,N_2914,N_2702);
or U6365 (N_6365,N_3939,N_3134);
and U6366 (N_6366,N_4854,N_3592);
or U6367 (N_6367,N_2732,N_3850);
and U6368 (N_6368,N_3051,N_4025);
nor U6369 (N_6369,N_3295,N_2613);
and U6370 (N_6370,N_3071,N_4789);
nand U6371 (N_6371,N_4975,N_3132);
or U6372 (N_6372,N_3784,N_3430);
or U6373 (N_6373,N_2535,N_3057);
or U6374 (N_6374,N_3503,N_4581);
nand U6375 (N_6375,N_4613,N_3679);
and U6376 (N_6376,N_4866,N_3710);
xor U6377 (N_6377,N_3847,N_2998);
and U6378 (N_6378,N_4983,N_3736);
and U6379 (N_6379,N_4000,N_2912);
or U6380 (N_6380,N_3109,N_3114);
nand U6381 (N_6381,N_2635,N_3351);
or U6382 (N_6382,N_4037,N_4562);
nand U6383 (N_6383,N_4913,N_3454);
and U6384 (N_6384,N_2654,N_3525);
nand U6385 (N_6385,N_4857,N_4946);
xor U6386 (N_6386,N_4738,N_3788);
and U6387 (N_6387,N_3585,N_4838);
xnor U6388 (N_6388,N_3735,N_2948);
nor U6389 (N_6389,N_3250,N_3394);
nor U6390 (N_6390,N_2978,N_2582);
nand U6391 (N_6391,N_3054,N_4463);
or U6392 (N_6392,N_3121,N_3536);
or U6393 (N_6393,N_4083,N_4700);
and U6394 (N_6394,N_4911,N_3533);
nand U6395 (N_6395,N_3864,N_4269);
nand U6396 (N_6396,N_3392,N_4097);
nand U6397 (N_6397,N_4952,N_3277);
or U6398 (N_6398,N_2826,N_2909);
xnor U6399 (N_6399,N_3308,N_3916);
nor U6400 (N_6400,N_4343,N_3361);
nor U6401 (N_6401,N_3540,N_3878);
nor U6402 (N_6402,N_3447,N_4172);
or U6403 (N_6403,N_3570,N_3366);
xor U6404 (N_6404,N_3718,N_4986);
or U6405 (N_6405,N_4392,N_3459);
nand U6406 (N_6406,N_2677,N_3801);
nand U6407 (N_6407,N_3926,N_3334);
nand U6408 (N_6408,N_3639,N_4566);
and U6409 (N_6409,N_3806,N_4378);
nor U6410 (N_6410,N_3266,N_3655);
and U6411 (N_6411,N_4591,N_4530);
or U6412 (N_6412,N_4111,N_4097);
nand U6413 (N_6413,N_3786,N_3708);
nand U6414 (N_6414,N_3763,N_3947);
nand U6415 (N_6415,N_3973,N_4688);
nor U6416 (N_6416,N_3442,N_4902);
nand U6417 (N_6417,N_4249,N_4679);
nand U6418 (N_6418,N_4287,N_4787);
and U6419 (N_6419,N_3330,N_3755);
nand U6420 (N_6420,N_3130,N_3231);
nand U6421 (N_6421,N_3013,N_4169);
and U6422 (N_6422,N_3529,N_3487);
nor U6423 (N_6423,N_3455,N_4077);
nand U6424 (N_6424,N_3197,N_4729);
nand U6425 (N_6425,N_4451,N_2960);
or U6426 (N_6426,N_3877,N_3008);
or U6427 (N_6427,N_3773,N_4923);
or U6428 (N_6428,N_4705,N_2827);
and U6429 (N_6429,N_4970,N_3862);
or U6430 (N_6430,N_2604,N_2510);
xor U6431 (N_6431,N_2691,N_4206);
or U6432 (N_6432,N_3245,N_3709);
or U6433 (N_6433,N_3217,N_4300);
nor U6434 (N_6434,N_3280,N_4510);
or U6435 (N_6435,N_4449,N_4086);
nand U6436 (N_6436,N_4311,N_3127);
or U6437 (N_6437,N_4365,N_4400);
nand U6438 (N_6438,N_2649,N_3126);
or U6439 (N_6439,N_4942,N_3932);
and U6440 (N_6440,N_2562,N_4813);
or U6441 (N_6441,N_3140,N_3525);
nor U6442 (N_6442,N_3850,N_4049);
nand U6443 (N_6443,N_4254,N_4580);
and U6444 (N_6444,N_4473,N_4676);
and U6445 (N_6445,N_2940,N_3071);
and U6446 (N_6446,N_2869,N_3780);
or U6447 (N_6447,N_3592,N_3924);
nand U6448 (N_6448,N_3002,N_3644);
or U6449 (N_6449,N_3055,N_4807);
or U6450 (N_6450,N_2537,N_3493);
xnor U6451 (N_6451,N_3200,N_3367);
or U6452 (N_6452,N_2951,N_3280);
or U6453 (N_6453,N_4265,N_4216);
or U6454 (N_6454,N_4004,N_3112);
and U6455 (N_6455,N_3647,N_3853);
or U6456 (N_6456,N_4992,N_3015);
and U6457 (N_6457,N_3719,N_4449);
nand U6458 (N_6458,N_4608,N_2978);
or U6459 (N_6459,N_4499,N_3118);
nor U6460 (N_6460,N_4384,N_4184);
or U6461 (N_6461,N_3540,N_2662);
nor U6462 (N_6462,N_2929,N_3580);
or U6463 (N_6463,N_4019,N_3317);
nor U6464 (N_6464,N_3837,N_4733);
nand U6465 (N_6465,N_3996,N_4054);
nor U6466 (N_6466,N_4917,N_4534);
nand U6467 (N_6467,N_4139,N_2750);
and U6468 (N_6468,N_4176,N_3875);
nor U6469 (N_6469,N_4304,N_3976);
nor U6470 (N_6470,N_2900,N_3909);
and U6471 (N_6471,N_3755,N_4870);
nand U6472 (N_6472,N_3626,N_4655);
or U6473 (N_6473,N_4081,N_3687);
nand U6474 (N_6474,N_2913,N_4095);
xnor U6475 (N_6475,N_4605,N_3609);
nor U6476 (N_6476,N_2561,N_3441);
nor U6477 (N_6477,N_4483,N_2534);
nor U6478 (N_6478,N_3613,N_2997);
nand U6479 (N_6479,N_4866,N_2723);
or U6480 (N_6480,N_2623,N_3486);
nand U6481 (N_6481,N_2513,N_4300);
nand U6482 (N_6482,N_3041,N_3591);
nor U6483 (N_6483,N_3608,N_2686);
or U6484 (N_6484,N_4555,N_3431);
nor U6485 (N_6485,N_2991,N_4867);
xor U6486 (N_6486,N_3271,N_2816);
or U6487 (N_6487,N_4675,N_2675);
or U6488 (N_6488,N_2788,N_4733);
and U6489 (N_6489,N_4533,N_2509);
nor U6490 (N_6490,N_3087,N_3972);
nand U6491 (N_6491,N_3383,N_4669);
and U6492 (N_6492,N_4814,N_3642);
nor U6493 (N_6493,N_3239,N_3667);
or U6494 (N_6494,N_4563,N_3759);
and U6495 (N_6495,N_4467,N_4636);
or U6496 (N_6496,N_4334,N_4273);
xor U6497 (N_6497,N_2732,N_4860);
nor U6498 (N_6498,N_3580,N_4170);
or U6499 (N_6499,N_3892,N_3001);
nand U6500 (N_6500,N_4206,N_2670);
xor U6501 (N_6501,N_4329,N_4837);
and U6502 (N_6502,N_4331,N_3208);
nor U6503 (N_6503,N_2791,N_2702);
or U6504 (N_6504,N_2978,N_4659);
and U6505 (N_6505,N_2629,N_4282);
or U6506 (N_6506,N_4323,N_4179);
or U6507 (N_6507,N_4492,N_2709);
xor U6508 (N_6508,N_4850,N_4088);
nand U6509 (N_6509,N_3615,N_4324);
xnor U6510 (N_6510,N_4864,N_3308);
or U6511 (N_6511,N_2673,N_3002);
and U6512 (N_6512,N_3604,N_2764);
nand U6513 (N_6513,N_3576,N_2827);
nor U6514 (N_6514,N_3274,N_3821);
nor U6515 (N_6515,N_4836,N_4860);
nor U6516 (N_6516,N_4196,N_3965);
nor U6517 (N_6517,N_4003,N_2726);
nor U6518 (N_6518,N_4661,N_4751);
or U6519 (N_6519,N_3302,N_4921);
nand U6520 (N_6520,N_3388,N_4928);
nor U6521 (N_6521,N_4155,N_4158);
or U6522 (N_6522,N_3491,N_3151);
nor U6523 (N_6523,N_4295,N_2889);
and U6524 (N_6524,N_4289,N_4501);
nor U6525 (N_6525,N_3628,N_4071);
nand U6526 (N_6526,N_4383,N_3141);
or U6527 (N_6527,N_4334,N_4634);
or U6528 (N_6528,N_3162,N_3249);
and U6529 (N_6529,N_2863,N_3511);
or U6530 (N_6530,N_4864,N_3391);
or U6531 (N_6531,N_4886,N_4100);
and U6532 (N_6532,N_2581,N_2722);
or U6533 (N_6533,N_3779,N_3771);
nand U6534 (N_6534,N_3797,N_4100);
and U6535 (N_6535,N_3711,N_3338);
nand U6536 (N_6536,N_2922,N_3264);
nand U6537 (N_6537,N_4348,N_3566);
and U6538 (N_6538,N_3721,N_2852);
or U6539 (N_6539,N_3733,N_4585);
nor U6540 (N_6540,N_2652,N_3104);
or U6541 (N_6541,N_4109,N_4674);
nand U6542 (N_6542,N_4557,N_3942);
or U6543 (N_6543,N_3706,N_4528);
or U6544 (N_6544,N_4352,N_3654);
and U6545 (N_6545,N_3224,N_4271);
nor U6546 (N_6546,N_4891,N_2511);
nand U6547 (N_6547,N_3253,N_4580);
and U6548 (N_6548,N_2693,N_4967);
nand U6549 (N_6549,N_3068,N_3308);
and U6550 (N_6550,N_3889,N_4709);
or U6551 (N_6551,N_4784,N_4582);
and U6552 (N_6552,N_4829,N_2919);
or U6553 (N_6553,N_3944,N_4816);
or U6554 (N_6554,N_3520,N_4960);
nand U6555 (N_6555,N_4762,N_4938);
or U6556 (N_6556,N_3937,N_3085);
or U6557 (N_6557,N_3014,N_2684);
or U6558 (N_6558,N_3495,N_4953);
nand U6559 (N_6559,N_3145,N_2958);
nand U6560 (N_6560,N_4454,N_3330);
nand U6561 (N_6561,N_2975,N_3594);
and U6562 (N_6562,N_2924,N_4691);
xor U6563 (N_6563,N_3900,N_2772);
and U6564 (N_6564,N_2759,N_3817);
xor U6565 (N_6565,N_4668,N_3016);
xor U6566 (N_6566,N_3816,N_3605);
nor U6567 (N_6567,N_4282,N_3500);
or U6568 (N_6568,N_3820,N_2683);
or U6569 (N_6569,N_3482,N_3740);
nand U6570 (N_6570,N_4038,N_4234);
or U6571 (N_6571,N_2763,N_3323);
nand U6572 (N_6572,N_4911,N_2705);
and U6573 (N_6573,N_3628,N_3644);
and U6574 (N_6574,N_4841,N_3756);
nand U6575 (N_6575,N_4183,N_4347);
and U6576 (N_6576,N_3649,N_3953);
nand U6577 (N_6577,N_3172,N_3896);
and U6578 (N_6578,N_4253,N_3062);
and U6579 (N_6579,N_3149,N_3733);
and U6580 (N_6580,N_4255,N_3875);
nor U6581 (N_6581,N_4146,N_2889);
xor U6582 (N_6582,N_4094,N_4061);
nor U6583 (N_6583,N_4907,N_3189);
nor U6584 (N_6584,N_2691,N_3093);
nor U6585 (N_6585,N_3186,N_2842);
xnor U6586 (N_6586,N_3264,N_3529);
nand U6587 (N_6587,N_4029,N_3631);
nand U6588 (N_6588,N_3636,N_2629);
or U6589 (N_6589,N_2906,N_3050);
or U6590 (N_6590,N_4365,N_4410);
or U6591 (N_6591,N_4683,N_4407);
and U6592 (N_6592,N_4026,N_3932);
and U6593 (N_6593,N_4233,N_3556);
or U6594 (N_6594,N_4086,N_4673);
and U6595 (N_6595,N_4861,N_4432);
or U6596 (N_6596,N_3772,N_4693);
and U6597 (N_6597,N_2586,N_3422);
and U6598 (N_6598,N_2912,N_2650);
and U6599 (N_6599,N_4601,N_4156);
or U6600 (N_6600,N_4982,N_4616);
and U6601 (N_6601,N_2552,N_2683);
nor U6602 (N_6602,N_3365,N_3936);
or U6603 (N_6603,N_4029,N_2791);
or U6604 (N_6604,N_3092,N_4483);
nor U6605 (N_6605,N_2924,N_4777);
nor U6606 (N_6606,N_3025,N_4012);
or U6607 (N_6607,N_3737,N_4897);
nor U6608 (N_6608,N_3190,N_3859);
and U6609 (N_6609,N_3928,N_4037);
or U6610 (N_6610,N_2655,N_2743);
nor U6611 (N_6611,N_3341,N_3646);
and U6612 (N_6612,N_3031,N_3853);
nand U6613 (N_6613,N_2645,N_4970);
and U6614 (N_6614,N_3387,N_2727);
or U6615 (N_6615,N_3044,N_4578);
nor U6616 (N_6616,N_3334,N_4591);
nand U6617 (N_6617,N_3332,N_4962);
or U6618 (N_6618,N_3475,N_4653);
or U6619 (N_6619,N_4726,N_4176);
and U6620 (N_6620,N_2531,N_4237);
xor U6621 (N_6621,N_3223,N_3522);
nor U6622 (N_6622,N_4770,N_4794);
and U6623 (N_6623,N_4000,N_3599);
nor U6624 (N_6624,N_4022,N_2630);
nor U6625 (N_6625,N_3621,N_2911);
nor U6626 (N_6626,N_4078,N_3701);
or U6627 (N_6627,N_3749,N_4355);
or U6628 (N_6628,N_4421,N_3513);
xnor U6629 (N_6629,N_3775,N_3047);
nand U6630 (N_6630,N_2825,N_4729);
or U6631 (N_6631,N_4554,N_2674);
nand U6632 (N_6632,N_4242,N_4401);
or U6633 (N_6633,N_3221,N_4297);
nand U6634 (N_6634,N_3928,N_4525);
or U6635 (N_6635,N_2963,N_4546);
nand U6636 (N_6636,N_2673,N_3653);
or U6637 (N_6637,N_3065,N_2905);
and U6638 (N_6638,N_4076,N_4151);
xnor U6639 (N_6639,N_4795,N_3036);
nor U6640 (N_6640,N_2932,N_3857);
or U6641 (N_6641,N_3899,N_3126);
or U6642 (N_6642,N_3657,N_4282);
nand U6643 (N_6643,N_3767,N_3120);
nand U6644 (N_6644,N_4122,N_4007);
or U6645 (N_6645,N_4527,N_3836);
and U6646 (N_6646,N_3582,N_2736);
and U6647 (N_6647,N_3518,N_3439);
nand U6648 (N_6648,N_3389,N_3649);
nor U6649 (N_6649,N_4715,N_2910);
nor U6650 (N_6650,N_3706,N_3058);
nand U6651 (N_6651,N_3665,N_2592);
nand U6652 (N_6652,N_3653,N_3662);
or U6653 (N_6653,N_2966,N_4294);
or U6654 (N_6654,N_4649,N_4999);
xnor U6655 (N_6655,N_3074,N_3064);
nand U6656 (N_6656,N_2725,N_2695);
nand U6657 (N_6657,N_4484,N_3443);
and U6658 (N_6658,N_4526,N_2661);
and U6659 (N_6659,N_4946,N_4395);
xor U6660 (N_6660,N_4477,N_3145);
xor U6661 (N_6661,N_3974,N_2815);
or U6662 (N_6662,N_3849,N_3901);
nor U6663 (N_6663,N_4557,N_4130);
nor U6664 (N_6664,N_3685,N_3740);
and U6665 (N_6665,N_3098,N_4546);
or U6666 (N_6666,N_4960,N_4764);
or U6667 (N_6667,N_4983,N_3244);
nor U6668 (N_6668,N_3553,N_4556);
or U6669 (N_6669,N_3319,N_3992);
nor U6670 (N_6670,N_4996,N_4980);
nor U6671 (N_6671,N_4040,N_4986);
nor U6672 (N_6672,N_3631,N_3752);
nor U6673 (N_6673,N_4849,N_3741);
nand U6674 (N_6674,N_4414,N_4082);
nand U6675 (N_6675,N_4805,N_3952);
xnor U6676 (N_6676,N_3055,N_3531);
nand U6677 (N_6677,N_2808,N_2931);
and U6678 (N_6678,N_3963,N_4482);
nand U6679 (N_6679,N_4185,N_4422);
nor U6680 (N_6680,N_4734,N_4064);
and U6681 (N_6681,N_3357,N_4073);
nand U6682 (N_6682,N_4831,N_3778);
xor U6683 (N_6683,N_2691,N_4823);
nand U6684 (N_6684,N_4200,N_2917);
and U6685 (N_6685,N_2822,N_3228);
and U6686 (N_6686,N_4180,N_3339);
xnor U6687 (N_6687,N_2646,N_4112);
nor U6688 (N_6688,N_3588,N_3595);
nor U6689 (N_6689,N_3666,N_2739);
nor U6690 (N_6690,N_4221,N_4453);
nor U6691 (N_6691,N_4940,N_3540);
xnor U6692 (N_6692,N_4057,N_3044);
or U6693 (N_6693,N_3095,N_4616);
or U6694 (N_6694,N_4854,N_4243);
nand U6695 (N_6695,N_3174,N_2989);
nor U6696 (N_6696,N_4464,N_4972);
xor U6697 (N_6697,N_4797,N_4398);
nor U6698 (N_6698,N_3394,N_4202);
nor U6699 (N_6699,N_4892,N_2944);
and U6700 (N_6700,N_3492,N_4463);
nor U6701 (N_6701,N_3417,N_2714);
nor U6702 (N_6702,N_3633,N_4145);
nor U6703 (N_6703,N_2812,N_3967);
nor U6704 (N_6704,N_2742,N_2983);
nor U6705 (N_6705,N_2852,N_2832);
and U6706 (N_6706,N_4876,N_4769);
or U6707 (N_6707,N_4985,N_4943);
and U6708 (N_6708,N_3677,N_2946);
or U6709 (N_6709,N_3558,N_3302);
or U6710 (N_6710,N_3229,N_4466);
nand U6711 (N_6711,N_2643,N_3805);
and U6712 (N_6712,N_4106,N_3893);
xor U6713 (N_6713,N_3086,N_3775);
nor U6714 (N_6714,N_3277,N_4186);
nand U6715 (N_6715,N_3855,N_2735);
or U6716 (N_6716,N_4910,N_3227);
nor U6717 (N_6717,N_2976,N_4507);
nand U6718 (N_6718,N_4788,N_4631);
and U6719 (N_6719,N_3502,N_3248);
or U6720 (N_6720,N_3458,N_3118);
or U6721 (N_6721,N_3764,N_3426);
or U6722 (N_6722,N_3148,N_4093);
xor U6723 (N_6723,N_4655,N_4342);
and U6724 (N_6724,N_3356,N_4117);
nor U6725 (N_6725,N_4156,N_4299);
nor U6726 (N_6726,N_3040,N_4792);
nand U6727 (N_6727,N_3924,N_4036);
and U6728 (N_6728,N_4554,N_3937);
nor U6729 (N_6729,N_4775,N_3705);
and U6730 (N_6730,N_3320,N_4073);
nand U6731 (N_6731,N_4875,N_2777);
and U6732 (N_6732,N_4029,N_4657);
nand U6733 (N_6733,N_4277,N_4442);
or U6734 (N_6734,N_3532,N_4348);
and U6735 (N_6735,N_3517,N_2621);
and U6736 (N_6736,N_4978,N_4762);
nor U6737 (N_6737,N_3735,N_4975);
or U6738 (N_6738,N_3697,N_2540);
and U6739 (N_6739,N_2594,N_2679);
nor U6740 (N_6740,N_3599,N_4386);
nor U6741 (N_6741,N_2829,N_3406);
or U6742 (N_6742,N_2694,N_4125);
nor U6743 (N_6743,N_3556,N_3392);
or U6744 (N_6744,N_3014,N_2512);
nor U6745 (N_6745,N_2689,N_3003);
or U6746 (N_6746,N_4048,N_4284);
nor U6747 (N_6747,N_4770,N_4457);
or U6748 (N_6748,N_4486,N_3548);
and U6749 (N_6749,N_3083,N_3740);
nor U6750 (N_6750,N_3265,N_4253);
and U6751 (N_6751,N_4059,N_3324);
nand U6752 (N_6752,N_4430,N_3389);
nor U6753 (N_6753,N_3760,N_3346);
nand U6754 (N_6754,N_3965,N_3984);
and U6755 (N_6755,N_3424,N_4963);
or U6756 (N_6756,N_4950,N_4777);
nor U6757 (N_6757,N_4087,N_3939);
nor U6758 (N_6758,N_3512,N_3837);
or U6759 (N_6759,N_3509,N_2719);
or U6760 (N_6760,N_4449,N_3356);
nor U6761 (N_6761,N_4709,N_3708);
or U6762 (N_6762,N_2677,N_3922);
nor U6763 (N_6763,N_4075,N_3567);
nand U6764 (N_6764,N_2886,N_2785);
or U6765 (N_6765,N_3540,N_4510);
or U6766 (N_6766,N_2805,N_3119);
nor U6767 (N_6767,N_4559,N_2590);
nor U6768 (N_6768,N_4480,N_4855);
xor U6769 (N_6769,N_3754,N_4250);
or U6770 (N_6770,N_3055,N_2914);
nand U6771 (N_6771,N_2967,N_3188);
xor U6772 (N_6772,N_4887,N_4752);
xor U6773 (N_6773,N_3414,N_4118);
nor U6774 (N_6774,N_4857,N_4745);
xor U6775 (N_6775,N_3969,N_3686);
or U6776 (N_6776,N_3873,N_3418);
nor U6777 (N_6777,N_2899,N_2797);
nand U6778 (N_6778,N_3236,N_2548);
nor U6779 (N_6779,N_4216,N_4176);
or U6780 (N_6780,N_3400,N_4958);
and U6781 (N_6781,N_2524,N_4243);
nand U6782 (N_6782,N_4003,N_3300);
nand U6783 (N_6783,N_2963,N_4610);
nor U6784 (N_6784,N_3610,N_3647);
and U6785 (N_6785,N_3685,N_3052);
nor U6786 (N_6786,N_4489,N_4592);
or U6787 (N_6787,N_3824,N_4729);
xnor U6788 (N_6788,N_4465,N_3331);
nor U6789 (N_6789,N_4518,N_3422);
nand U6790 (N_6790,N_4524,N_3993);
xor U6791 (N_6791,N_3305,N_4568);
nor U6792 (N_6792,N_3948,N_2665);
xor U6793 (N_6793,N_3438,N_2975);
and U6794 (N_6794,N_2716,N_4133);
or U6795 (N_6795,N_4444,N_4710);
and U6796 (N_6796,N_4843,N_3230);
or U6797 (N_6797,N_3785,N_2878);
nor U6798 (N_6798,N_3427,N_3272);
or U6799 (N_6799,N_4240,N_4187);
nand U6800 (N_6800,N_4126,N_3330);
nand U6801 (N_6801,N_4434,N_3228);
and U6802 (N_6802,N_3856,N_4349);
and U6803 (N_6803,N_4029,N_4584);
nand U6804 (N_6804,N_4626,N_3824);
nor U6805 (N_6805,N_4827,N_4523);
nand U6806 (N_6806,N_4404,N_4344);
nor U6807 (N_6807,N_2840,N_3590);
or U6808 (N_6808,N_3665,N_4635);
and U6809 (N_6809,N_4077,N_3473);
and U6810 (N_6810,N_4878,N_4967);
and U6811 (N_6811,N_2740,N_3743);
nor U6812 (N_6812,N_2678,N_3636);
nor U6813 (N_6813,N_2610,N_3570);
nor U6814 (N_6814,N_4129,N_4295);
and U6815 (N_6815,N_3950,N_3215);
nand U6816 (N_6816,N_2769,N_4901);
nor U6817 (N_6817,N_4329,N_4797);
nand U6818 (N_6818,N_2895,N_2592);
or U6819 (N_6819,N_2907,N_4055);
nor U6820 (N_6820,N_4785,N_3983);
or U6821 (N_6821,N_3629,N_3772);
or U6822 (N_6822,N_2704,N_2560);
nand U6823 (N_6823,N_2587,N_2596);
and U6824 (N_6824,N_2801,N_3212);
nand U6825 (N_6825,N_2546,N_3640);
or U6826 (N_6826,N_4897,N_3302);
or U6827 (N_6827,N_3113,N_3805);
or U6828 (N_6828,N_3010,N_3273);
and U6829 (N_6829,N_4179,N_3430);
xor U6830 (N_6830,N_2858,N_4075);
xnor U6831 (N_6831,N_2668,N_4962);
and U6832 (N_6832,N_3445,N_4527);
nor U6833 (N_6833,N_4797,N_4640);
and U6834 (N_6834,N_3248,N_3571);
nor U6835 (N_6835,N_2504,N_3716);
and U6836 (N_6836,N_4865,N_4581);
or U6837 (N_6837,N_4273,N_2778);
nor U6838 (N_6838,N_4574,N_3825);
and U6839 (N_6839,N_3509,N_4658);
nand U6840 (N_6840,N_2864,N_4803);
xor U6841 (N_6841,N_3598,N_3612);
nand U6842 (N_6842,N_4480,N_3310);
xnor U6843 (N_6843,N_3136,N_3494);
nand U6844 (N_6844,N_3656,N_4273);
nand U6845 (N_6845,N_2952,N_3186);
or U6846 (N_6846,N_3007,N_3158);
nor U6847 (N_6847,N_4381,N_4968);
nor U6848 (N_6848,N_3386,N_2964);
and U6849 (N_6849,N_4355,N_3731);
or U6850 (N_6850,N_3145,N_2956);
nand U6851 (N_6851,N_4920,N_4802);
or U6852 (N_6852,N_3330,N_3021);
or U6853 (N_6853,N_4442,N_3413);
or U6854 (N_6854,N_3119,N_3402);
nor U6855 (N_6855,N_4984,N_2532);
and U6856 (N_6856,N_4531,N_2656);
nor U6857 (N_6857,N_3568,N_3797);
and U6858 (N_6858,N_4984,N_3595);
and U6859 (N_6859,N_3046,N_4652);
and U6860 (N_6860,N_3585,N_4954);
nand U6861 (N_6861,N_4873,N_4674);
xor U6862 (N_6862,N_2514,N_3383);
nor U6863 (N_6863,N_4552,N_3244);
or U6864 (N_6864,N_4297,N_3379);
xnor U6865 (N_6865,N_4946,N_4109);
nand U6866 (N_6866,N_2968,N_2579);
and U6867 (N_6867,N_3591,N_4349);
or U6868 (N_6868,N_4077,N_3651);
or U6869 (N_6869,N_3763,N_3008);
nand U6870 (N_6870,N_2521,N_3293);
nand U6871 (N_6871,N_4661,N_3578);
and U6872 (N_6872,N_4817,N_4338);
nand U6873 (N_6873,N_2956,N_4699);
nor U6874 (N_6874,N_4517,N_3954);
and U6875 (N_6875,N_3682,N_2901);
nor U6876 (N_6876,N_2918,N_3529);
and U6877 (N_6877,N_3732,N_2838);
or U6878 (N_6878,N_2615,N_4123);
nor U6879 (N_6879,N_3087,N_3015);
and U6880 (N_6880,N_2894,N_4173);
or U6881 (N_6881,N_3082,N_4384);
nor U6882 (N_6882,N_3195,N_3419);
or U6883 (N_6883,N_4850,N_4818);
or U6884 (N_6884,N_3112,N_4261);
xnor U6885 (N_6885,N_3642,N_2647);
or U6886 (N_6886,N_2781,N_2538);
nor U6887 (N_6887,N_2989,N_2700);
and U6888 (N_6888,N_4199,N_2699);
or U6889 (N_6889,N_2798,N_3673);
nand U6890 (N_6890,N_3080,N_3609);
nand U6891 (N_6891,N_3837,N_4119);
nand U6892 (N_6892,N_3171,N_4076);
nor U6893 (N_6893,N_3247,N_4213);
and U6894 (N_6894,N_3380,N_3429);
nor U6895 (N_6895,N_2669,N_4328);
and U6896 (N_6896,N_4546,N_4634);
nor U6897 (N_6897,N_3401,N_3412);
nor U6898 (N_6898,N_2582,N_4610);
xnor U6899 (N_6899,N_3713,N_2962);
or U6900 (N_6900,N_3014,N_3123);
and U6901 (N_6901,N_4184,N_3071);
nor U6902 (N_6902,N_4368,N_3060);
nor U6903 (N_6903,N_3332,N_2776);
or U6904 (N_6904,N_4799,N_3171);
xor U6905 (N_6905,N_3990,N_4404);
nor U6906 (N_6906,N_3563,N_4265);
nor U6907 (N_6907,N_4202,N_3912);
or U6908 (N_6908,N_4771,N_4308);
nor U6909 (N_6909,N_3993,N_4935);
or U6910 (N_6910,N_4674,N_3798);
xnor U6911 (N_6911,N_4743,N_4202);
and U6912 (N_6912,N_3045,N_2751);
nand U6913 (N_6913,N_2578,N_4544);
xor U6914 (N_6914,N_3876,N_2843);
nand U6915 (N_6915,N_3352,N_3126);
and U6916 (N_6916,N_3997,N_2948);
nor U6917 (N_6917,N_4339,N_3618);
xnor U6918 (N_6918,N_2653,N_4289);
or U6919 (N_6919,N_4927,N_2519);
nor U6920 (N_6920,N_3447,N_3690);
nand U6921 (N_6921,N_4417,N_3959);
nor U6922 (N_6922,N_4740,N_4669);
nor U6923 (N_6923,N_2985,N_4124);
nand U6924 (N_6924,N_4971,N_2681);
and U6925 (N_6925,N_2975,N_3669);
nor U6926 (N_6926,N_4938,N_4223);
nand U6927 (N_6927,N_4765,N_2782);
nand U6928 (N_6928,N_2789,N_3158);
nor U6929 (N_6929,N_3195,N_4137);
nand U6930 (N_6930,N_3968,N_4585);
or U6931 (N_6931,N_4983,N_2875);
nor U6932 (N_6932,N_3497,N_3412);
nand U6933 (N_6933,N_4354,N_2982);
or U6934 (N_6934,N_2811,N_4921);
nor U6935 (N_6935,N_2717,N_4234);
nand U6936 (N_6936,N_3814,N_3455);
and U6937 (N_6937,N_3874,N_4759);
and U6938 (N_6938,N_4847,N_4650);
and U6939 (N_6939,N_3375,N_3661);
and U6940 (N_6940,N_3320,N_3273);
and U6941 (N_6941,N_4016,N_4462);
nor U6942 (N_6942,N_4172,N_4229);
nor U6943 (N_6943,N_4904,N_4687);
nand U6944 (N_6944,N_3631,N_4372);
and U6945 (N_6945,N_3734,N_4258);
nand U6946 (N_6946,N_2673,N_3298);
and U6947 (N_6947,N_4760,N_3694);
nor U6948 (N_6948,N_3350,N_3207);
nor U6949 (N_6949,N_4766,N_3469);
or U6950 (N_6950,N_4079,N_2874);
nand U6951 (N_6951,N_4436,N_4277);
and U6952 (N_6952,N_3229,N_3190);
nand U6953 (N_6953,N_4188,N_4537);
nand U6954 (N_6954,N_4064,N_3808);
or U6955 (N_6955,N_4783,N_3911);
or U6956 (N_6956,N_2966,N_3435);
nand U6957 (N_6957,N_4570,N_2683);
nor U6958 (N_6958,N_4413,N_3240);
nand U6959 (N_6959,N_3404,N_4880);
nand U6960 (N_6960,N_3351,N_4721);
and U6961 (N_6961,N_4226,N_3957);
nor U6962 (N_6962,N_2783,N_4099);
nand U6963 (N_6963,N_4554,N_2527);
nand U6964 (N_6964,N_3207,N_4866);
nor U6965 (N_6965,N_3679,N_2918);
nand U6966 (N_6966,N_2807,N_4178);
and U6967 (N_6967,N_3267,N_4251);
xor U6968 (N_6968,N_3800,N_3694);
or U6969 (N_6969,N_4773,N_3537);
or U6970 (N_6970,N_3542,N_3786);
nor U6971 (N_6971,N_2500,N_3371);
nand U6972 (N_6972,N_3439,N_4241);
nor U6973 (N_6973,N_3986,N_4808);
nor U6974 (N_6974,N_3015,N_4040);
and U6975 (N_6975,N_3858,N_3357);
nand U6976 (N_6976,N_2596,N_3015);
nand U6977 (N_6977,N_4155,N_4513);
and U6978 (N_6978,N_2663,N_4351);
and U6979 (N_6979,N_3982,N_3214);
nor U6980 (N_6980,N_3169,N_4313);
or U6981 (N_6981,N_3314,N_3174);
and U6982 (N_6982,N_4821,N_2763);
xor U6983 (N_6983,N_3286,N_4691);
or U6984 (N_6984,N_2694,N_3423);
nand U6985 (N_6985,N_3355,N_4225);
nand U6986 (N_6986,N_4331,N_4917);
or U6987 (N_6987,N_3498,N_2519);
nand U6988 (N_6988,N_4964,N_4631);
and U6989 (N_6989,N_3511,N_4799);
nand U6990 (N_6990,N_3384,N_3235);
xnor U6991 (N_6991,N_4167,N_4424);
nand U6992 (N_6992,N_3095,N_4902);
nand U6993 (N_6993,N_3056,N_4274);
nor U6994 (N_6994,N_3252,N_4679);
or U6995 (N_6995,N_2744,N_3163);
nand U6996 (N_6996,N_3297,N_3643);
nand U6997 (N_6997,N_3750,N_3828);
and U6998 (N_6998,N_3086,N_3340);
or U6999 (N_6999,N_3425,N_4966);
nor U7000 (N_7000,N_4825,N_2928);
and U7001 (N_7001,N_3348,N_2538);
nor U7002 (N_7002,N_4530,N_4866);
or U7003 (N_7003,N_3889,N_3251);
and U7004 (N_7004,N_3164,N_4749);
and U7005 (N_7005,N_4749,N_4198);
and U7006 (N_7006,N_4998,N_3416);
and U7007 (N_7007,N_4067,N_3977);
nand U7008 (N_7008,N_4697,N_4776);
and U7009 (N_7009,N_3977,N_4220);
nand U7010 (N_7010,N_4534,N_4067);
xor U7011 (N_7011,N_4472,N_4759);
or U7012 (N_7012,N_4755,N_4654);
nor U7013 (N_7013,N_3337,N_4631);
xor U7014 (N_7014,N_2739,N_4822);
or U7015 (N_7015,N_4161,N_4155);
nand U7016 (N_7016,N_4404,N_4489);
and U7017 (N_7017,N_3454,N_4345);
nor U7018 (N_7018,N_4306,N_2571);
nand U7019 (N_7019,N_3166,N_2668);
nor U7020 (N_7020,N_4901,N_2919);
nor U7021 (N_7021,N_4721,N_4205);
nand U7022 (N_7022,N_4693,N_3511);
and U7023 (N_7023,N_4028,N_3776);
nand U7024 (N_7024,N_3021,N_3207);
xor U7025 (N_7025,N_3462,N_2506);
or U7026 (N_7026,N_4450,N_4877);
or U7027 (N_7027,N_3564,N_2651);
nand U7028 (N_7028,N_2516,N_2821);
nor U7029 (N_7029,N_4991,N_3692);
or U7030 (N_7030,N_2624,N_3057);
or U7031 (N_7031,N_4197,N_3855);
or U7032 (N_7032,N_4485,N_4542);
nand U7033 (N_7033,N_2776,N_3999);
xor U7034 (N_7034,N_4040,N_2501);
and U7035 (N_7035,N_4307,N_3878);
xnor U7036 (N_7036,N_4169,N_2602);
nand U7037 (N_7037,N_3238,N_2521);
nor U7038 (N_7038,N_4973,N_3832);
or U7039 (N_7039,N_4628,N_2656);
or U7040 (N_7040,N_3740,N_3549);
or U7041 (N_7041,N_3266,N_4711);
nand U7042 (N_7042,N_2935,N_4372);
and U7043 (N_7043,N_3778,N_3686);
nand U7044 (N_7044,N_3729,N_3089);
and U7045 (N_7045,N_4139,N_4625);
or U7046 (N_7046,N_3481,N_4490);
xnor U7047 (N_7047,N_2894,N_3604);
nor U7048 (N_7048,N_2691,N_4433);
and U7049 (N_7049,N_3535,N_3761);
or U7050 (N_7050,N_4589,N_4634);
or U7051 (N_7051,N_2874,N_3037);
nand U7052 (N_7052,N_3913,N_4477);
and U7053 (N_7053,N_4365,N_4526);
or U7054 (N_7054,N_4706,N_4985);
xnor U7055 (N_7055,N_2786,N_4088);
xnor U7056 (N_7056,N_4688,N_4594);
or U7057 (N_7057,N_4119,N_2536);
nor U7058 (N_7058,N_4215,N_3184);
nor U7059 (N_7059,N_4168,N_3936);
and U7060 (N_7060,N_2546,N_3100);
and U7061 (N_7061,N_4735,N_3824);
or U7062 (N_7062,N_4456,N_3731);
nand U7063 (N_7063,N_3109,N_3366);
nor U7064 (N_7064,N_4038,N_2559);
and U7065 (N_7065,N_3488,N_3106);
nor U7066 (N_7066,N_3236,N_4400);
or U7067 (N_7067,N_3481,N_4710);
or U7068 (N_7068,N_3603,N_4215);
nor U7069 (N_7069,N_4609,N_2958);
nand U7070 (N_7070,N_2662,N_3614);
nor U7071 (N_7071,N_2927,N_3110);
and U7072 (N_7072,N_4847,N_3904);
xor U7073 (N_7073,N_4784,N_2961);
or U7074 (N_7074,N_2565,N_2654);
nand U7075 (N_7075,N_3912,N_4558);
or U7076 (N_7076,N_4861,N_2575);
nand U7077 (N_7077,N_3890,N_3866);
nor U7078 (N_7078,N_4761,N_2705);
nor U7079 (N_7079,N_2960,N_4365);
nor U7080 (N_7080,N_2890,N_3666);
or U7081 (N_7081,N_2762,N_3467);
nand U7082 (N_7082,N_4416,N_3173);
nor U7083 (N_7083,N_3122,N_4238);
or U7084 (N_7084,N_3736,N_2517);
nand U7085 (N_7085,N_4504,N_2709);
nand U7086 (N_7086,N_3573,N_4134);
nor U7087 (N_7087,N_2512,N_4025);
nor U7088 (N_7088,N_4942,N_3674);
or U7089 (N_7089,N_2866,N_4075);
nor U7090 (N_7090,N_3976,N_4361);
nor U7091 (N_7091,N_2654,N_2857);
and U7092 (N_7092,N_4287,N_3405);
and U7093 (N_7093,N_3409,N_3152);
nor U7094 (N_7094,N_4849,N_3228);
nand U7095 (N_7095,N_4649,N_3457);
xor U7096 (N_7096,N_4500,N_2613);
nor U7097 (N_7097,N_3808,N_2550);
or U7098 (N_7098,N_4101,N_3308);
xor U7099 (N_7099,N_4010,N_4881);
nor U7100 (N_7100,N_3744,N_4430);
and U7101 (N_7101,N_4778,N_3103);
or U7102 (N_7102,N_3655,N_4214);
or U7103 (N_7103,N_4448,N_3465);
and U7104 (N_7104,N_2891,N_4178);
and U7105 (N_7105,N_4823,N_2618);
or U7106 (N_7106,N_3071,N_4970);
and U7107 (N_7107,N_3070,N_4881);
or U7108 (N_7108,N_4279,N_2803);
and U7109 (N_7109,N_4830,N_4062);
nor U7110 (N_7110,N_2559,N_2939);
and U7111 (N_7111,N_2764,N_3757);
nand U7112 (N_7112,N_4880,N_4539);
nand U7113 (N_7113,N_4877,N_2926);
nand U7114 (N_7114,N_3136,N_2902);
nand U7115 (N_7115,N_2622,N_4249);
or U7116 (N_7116,N_4148,N_2982);
nand U7117 (N_7117,N_3259,N_3290);
and U7118 (N_7118,N_2556,N_4762);
and U7119 (N_7119,N_3654,N_2587);
or U7120 (N_7120,N_4097,N_4465);
nand U7121 (N_7121,N_3156,N_3533);
nor U7122 (N_7122,N_4699,N_3502);
nand U7123 (N_7123,N_4549,N_4693);
and U7124 (N_7124,N_4797,N_4838);
nand U7125 (N_7125,N_3306,N_4894);
nor U7126 (N_7126,N_3226,N_3709);
nor U7127 (N_7127,N_4752,N_2674);
nor U7128 (N_7128,N_3293,N_4010);
nand U7129 (N_7129,N_3963,N_3727);
nand U7130 (N_7130,N_4518,N_2949);
nor U7131 (N_7131,N_3778,N_4146);
or U7132 (N_7132,N_4462,N_3770);
xor U7133 (N_7133,N_3327,N_2868);
nor U7134 (N_7134,N_4355,N_4619);
xor U7135 (N_7135,N_3129,N_3173);
nor U7136 (N_7136,N_3063,N_2750);
nor U7137 (N_7137,N_4082,N_2569);
nand U7138 (N_7138,N_4153,N_4335);
or U7139 (N_7139,N_3063,N_4306);
or U7140 (N_7140,N_3390,N_4790);
nor U7141 (N_7141,N_4315,N_3419);
nand U7142 (N_7142,N_2776,N_4171);
nor U7143 (N_7143,N_3487,N_4550);
nor U7144 (N_7144,N_3593,N_3612);
nand U7145 (N_7145,N_3559,N_4966);
nand U7146 (N_7146,N_4275,N_3375);
nor U7147 (N_7147,N_3799,N_4519);
and U7148 (N_7148,N_3215,N_3977);
and U7149 (N_7149,N_3772,N_4907);
nor U7150 (N_7150,N_4895,N_4747);
or U7151 (N_7151,N_4940,N_4129);
and U7152 (N_7152,N_4331,N_4342);
nand U7153 (N_7153,N_4311,N_3110);
and U7154 (N_7154,N_4587,N_3866);
and U7155 (N_7155,N_2977,N_4610);
nor U7156 (N_7156,N_4812,N_2583);
nand U7157 (N_7157,N_3251,N_2804);
nor U7158 (N_7158,N_3714,N_3851);
and U7159 (N_7159,N_4668,N_3281);
and U7160 (N_7160,N_3766,N_2920);
nor U7161 (N_7161,N_3683,N_2580);
and U7162 (N_7162,N_3901,N_4169);
and U7163 (N_7163,N_3297,N_2655);
nor U7164 (N_7164,N_4477,N_2734);
nor U7165 (N_7165,N_3158,N_4143);
xor U7166 (N_7166,N_3596,N_3170);
or U7167 (N_7167,N_3033,N_3343);
nor U7168 (N_7168,N_4642,N_4761);
and U7169 (N_7169,N_4707,N_4278);
xor U7170 (N_7170,N_4731,N_2889);
and U7171 (N_7171,N_3341,N_2878);
nand U7172 (N_7172,N_2639,N_4141);
and U7173 (N_7173,N_4976,N_3559);
xnor U7174 (N_7174,N_4363,N_3979);
nand U7175 (N_7175,N_2783,N_4473);
nand U7176 (N_7176,N_2882,N_4954);
nand U7177 (N_7177,N_2970,N_2640);
and U7178 (N_7178,N_4679,N_3141);
xor U7179 (N_7179,N_4291,N_3576);
nor U7180 (N_7180,N_2617,N_3217);
nand U7181 (N_7181,N_2811,N_3661);
nand U7182 (N_7182,N_4686,N_4264);
nor U7183 (N_7183,N_4986,N_3321);
or U7184 (N_7184,N_3681,N_2850);
and U7185 (N_7185,N_2949,N_4035);
and U7186 (N_7186,N_4525,N_3209);
nor U7187 (N_7187,N_3083,N_2528);
or U7188 (N_7188,N_4037,N_3274);
nor U7189 (N_7189,N_3483,N_4201);
nand U7190 (N_7190,N_3960,N_2763);
nor U7191 (N_7191,N_4557,N_3042);
nand U7192 (N_7192,N_4162,N_4636);
and U7193 (N_7193,N_3299,N_3501);
nand U7194 (N_7194,N_2558,N_4043);
nor U7195 (N_7195,N_3506,N_4379);
or U7196 (N_7196,N_4611,N_2775);
or U7197 (N_7197,N_4931,N_3536);
nor U7198 (N_7198,N_3990,N_4144);
xor U7199 (N_7199,N_2606,N_4582);
nor U7200 (N_7200,N_3308,N_2748);
nand U7201 (N_7201,N_3947,N_3515);
or U7202 (N_7202,N_3776,N_3485);
nor U7203 (N_7203,N_3253,N_4600);
nand U7204 (N_7204,N_4989,N_2718);
xor U7205 (N_7205,N_3425,N_4424);
nand U7206 (N_7206,N_3330,N_3237);
nand U7207 (N_7207,N_3438,N_4986);
or U7208 (N_7208,N_4954,N_4421);
or U7209 (N_7209,N_3711,N_3118);
nor U7210 (N_7210,N_4537,N_2735);
xor U7211 (N_7211,N_3472,N_3718);
nor U7212 (N_7212,N_2630,N_3941);
nor U7213 (N_7213,N_3667,N_2963);
xor U7214 (N_7214,N_2598,N_4762);
and U7215 (N_7215,N_4553,N_4860);
xnor U7216 (N_7216,N_2547,N_3904);
or U7217 (N_7217,N_4327,N_4947);
and U7218 (N_7218,N_3881,N_3294);
and U7219 (N_7219,N_3250,N_4237);
nand U7220 (N_7220,N_2843,N_2655);
or U7221 (N_7221,N_3717,N_4222);
nand U7222 (N_7222,N_3486,N_2865);
and U7223 (N_7223,N_2756,N_3029);
or U7224 (N_7224,N_4253,N_3234);
nor U7225 (N_7225,N_3873,N_3905);
xnor U7226 (N_7226,N_4140,N_3094);
nor U7227 (N_7227,N_3245,N_2618);
and U7228 (N_7228,N_4458,N_3477);
xnor U7229 (N_7229,N_4515,N_3911);
nor U7230 (N_7230,N_2920,N_4881);
or U7231 (N_7231,N_4227,N_4592);
nand U7232 (N_7232,N_3190,N_3182);
nand U7233 (N_7233,N_3072,N_3678);
nand U7234 (N_7234,N_3352,N_3146);
nor U7235 (N_7235,N_3743,N_2600);
nand U7236 (N_7236,N_2512,N_4095);
nor U7237 (N_7237,N_2855,N_3682);
and U7238 (N_7238,N_3020,N_4281);
xnor U7239 (N_7239,N_2643,N_2600);
nand U7240 (N_7240,N_4564,N_4271);
or U7241 (N_7241,N_2843,N_4572);
xor U7242 (N_7242,N_3909,N_2734);
xnor U7243 (N_7243,N_2577,N_2598);
nor U7244 (N_7244,N_3566,N_4970);
nand U7245 (N_7245,N_4047,N_3281);
xnor U7246 (N_7246,N_4160,N_4913);
nor U7247 (N_7247,N_3990,N_3633);
or U7248 (N_7248,N_3911,N_2765);
and U7249 (N_7249,N_2697,N_3186);
or U7250 (N_7250,N_2663,N_2837);
nand U7251 (N_7251,N_4173,N_3682);
or U7252 (N_7252,N_4587,N_4309);
or U7253 (N_7253,N_4700,N_4868);
nand U7254 (N_7254,N_3404,N_4057);
xor U7255 (N_7255,N_4390,N_2822);
or U7256 (N_7256,N_4536,N_3019);
nor U7257 (N_7257,N_3673,N_4316);
or U7258 (N_7258,N_3614,N_4839);
and U7259 (N_7259,N_3444,N_2524);
nand U7260 (N_7260,N_2516,N_2936);
and U7261 (N_7261,N_4467,N_3457);
nor U7262 (N_7262,N_4675,N_4111);
nand U7263 (N_7263,N_3531,N_2797);
and U7264 (N_7264,N_4486,N_3008);
or U7265 (N_7265,N_4369,N_3647);
or U7266 (N_7266,N_4814,N_3671);
nor U7267 (N_7267,N_3885,N_2546);
nand U7268 (N_7268,N_3171,N_3997);
nor U7269 (N_7269,N_4775,N_4484);
nand U7270 (N_7270,N_2916,N_4931);
nor U7271 (N_7271,N_4806,N_2847);
nor U7272 (N_7272,N_3348,N_4224);
or U7273 (N_7273,N_3007,N_3828);
or U7274 (N_7274,N_4889,N_4270);
xor U7275 (N_7275,N_4876,N_4376);
or U7276 (N_7276,N_2929,N_4694);
nand U7277 (N_7277,N_4351,N_3359);
nand U7278 (N_7278,N_3257,N_3249);
and U7279 (N_7279,N_3684,N_3176);
nand U7280 (N_7280,N_4602,N_3367);
or U7281 (N_7281,N_4875,N_4825);
or U7282 (N_7282,N_2639,N_4362);
nor U7283 (N_7283,N_3152,N_3039);
or U7284 (N_7284,N_2528,N_2917);
or U7285 (N_7285,N_4807,N_3057);
nand U7286 (N_7286,N_4466,N_4170);
nand U7287 (N_7287,N_4751,N_2590);
and U7288 (N_7288,N_4423,N_3939);
xnor U7289 (N_7289,N_3922,N_2802);
and U7290 (N_7290,N_4219,N_3935);
or U7291 (N_7291,N_4606,N_3586);
or U7292 (N_7292,N_4748,N_3747);
xnor U7293 (N_7293,N_3195,N_2926);
nor U7294 (N_7294,N_2730,N_4348);
xor U7295 (N_7295,N_3535,N_4173);
or U7296 (N_7296,N_3838,N_3334);
or U7297 (N_7297,N_4424,N_2968);
nor U7298 (N_7298,N_3603,N_2668);
nor U7299 (N_7299,N_4984,N_4105);
nor U7300 (N_7300,N_4051,N_3423);
and U7301 (N_7301,N_4662,N_2507);
nand U7302 (N_7302,N_4462,N_4704);
and U7303 (N_7303,N_4190,N_4279);
nand U7304 (N_7304,N_3612,N_3232);
nand U7305 (N_7305,N_2695,N_3012);
and U7306 (N_7306,N_2896,N_3178);
and U7307 (N_7307,N_3083,N_3999);
xor U7308 (N_7308,N_4069,N_3635);
nand U7309 (N_7309,N_4634,N_2722);
nand U7310 (N_7310,N_3030,N_4365);
or U7311 (N_7311,N_4022,N_3979);
nand U7312 (N_7312,N_3777,N_4980);
nand U7313 (N_7313,N_2875,N_3499);
or U7314 (N_7314,N_4734,N_2533);
xor U7315 (N_7315,N_3648,N_2531);
or U7316 (N_7316,N_2663,N_3681);
xnor U7317 (N_7317,N_2628,N_2611);
nor U7318 (N_7318,N_2541,N_4118);
and U7319 (N_7319,N_2684,N_3352);
xnor U7320 (N_7320,N_4059,N_4523);
and U7321 (N_7321,N_4518,N_3116);
nor U7322 (N_7322,N_3809,N_4221);
nand U7323 (N_7323,N_4313,N_4602);
or U7324 (N_7324,N_2568,N_4375);
nand U7325 (N_7325,N_4117,N_2617);
nor U7326 (N_7326,N_2907,N_4009);
xor U7327 (N_7327,N_3737,N_3535);
nor U7328 (N_7328,N_3177,N_2542);
or U7329 (N_7329,N_3109,N_4488);
and U7330 (N_7330,N_3359,N_4945);
or U7331 (N_7331,N_3449,N_2737);
or U7332 (N_7332,N_4713,N_3180);
and U7333 (N_7333,N_4977,N_2696);
nor U7334 (N_7334,N_4797,N_3018);
nand U7335 (N_7335,N_3851,N_3807);
and U7336 (N_7336,N_3142,N_4330);
nand U7337 (N_7337,N_4033,N_2539);
nor U7338 (N_7338,N_2839,N_4696);
and U7339 (N_7339,N_3078,N_3778);
and U7340 (N_7340,N_2647,N_4742);
nor U7341 (N_7341,N_2922,N_4511);
or U7342 (N_7342,N_3927,N_4969);
nand U7343 (N_7343,N_4726,N_4800);
or U7344 (N_7344,N_3222,N_4030);
nor U7345 (N_7345,N_3528,N_4960);
nand U7346 (N_7346,N_2733,N_2516);
nand U7347 (N_7347,N_3961,N_4436);
or U7348 (N_7348,N_4497,N_4557);
and U7349 (N_7349,N_4822,N_2924);
nor U7350 (N_7350,N_4190,N_4939);
or U7351 (N_7351,N_4445,N_2749);
xor U7352 (N_7352,N_4844,N_3822);
nand U7353 (N_7353,N_3229,N_2652);
and U7354 (N_7354,N_2794,N_3436);
or U7355 (N_7355,N_3659,N_2539);
and U7356 (N_7356,N_4613,N_3855);
nor U7357 (N_7357,N_4136,N_2986);
or U7358 (N_7358,N_4041,N_3243);
xor U7359 (N_7359,N_4508,N_4408);
or U7360 (N_7360,N_4383,N_4328);
nand U7361 (N_7361,N_3825,N_2743);
xnor U7362 (N_7362,N_3866,N_4459);
nor U7363 (N_7363,N_2731,N_3872);
nand U7364 (N_7364,N_2830,N_2678);
nand U7365 (N_7365,N_4308,N_2817);
nor U7366 (N_7366,N_4307,N_2824);
nand U7367 (N_7367,N_2787,N_3445);
xnor U7368 (N_7368,N_3296,N_2590);
nand U7369 (N_7369,N_3501,N_4929);
xor U7370 (N_7370,N_4636,N_2742);
and U7371 (N_7371,N_4101,N_3956);
nand U7372 (N_7372,N_3354,N_2791);
or U7373 (N_7373,N_4440,N_4768);
nor U7374 (N_7374,N_3816,N_3350);
and U7375 (N_7375,N_4120,N_3987);
or U7376 (N_7376,N_3875,N_3669);
and U7377 (N_7377,N_3838,N_2617);
and U7378 (N_7378,N_4774,N_3423);
nor U7379 (N_7379,N_3367,N_3435);
and U7380 (N_7380,N_2755,N_3812);
and U7381 (N_7381,N_3095,N_2559);
and U7382 (N_7382,N_4063,N_3631);
nand U7383 (N_7383,N_3683,N_2778);
nor U7384 (N_7384,N_3626,N_4001);
and U7385 (N_7385,N_4322,N_4840);
and U7386 (N_7386,N_3906,N_4924);
and U7387 (N_7387,N_4814,N_4426);
or U7388 (N_7388,N_4822,N_4397);
nand U7389 (N_7389,N_3435,N_4929);
or U7390 (N_7390,N_2657,N_3415);
nor U7391 (N_7391,N_2723,N_4625);
or U7392 (N_7392,N_2828,N_2862);
or U7393 (N_7393,N_2583,N_3357);
or U7394 (N_7394,N_4070,N_4592);
or U7395 (N_7395,N_2924,N_4169);
nor U7396 (N_7396,N_2789,N_2686);
nand U7397 (N_7397,N_3864,N_3197);
or U7398 (N_7398,N_4724,N_2778);
nand U7399 (N_7399,N_4924,N_3233);
and U7400 (N_7400,N_3472,N_4103);
nand U7401 (N_7401,N_4901,N_3986);
or U7402 (N_7402,N_4061,N_3915);
and U7403 (N_7403,N_2588,N_4515);
xor U7404 (N_7404,N_4067,N_3000);
nand U7405 (N_7405,N_3936,N_3057);
and U7406 (N_7406,N_4046,N_4379);
or U7407 (N_7407,N_3659,N_3370);
nand U7408 (N_7408,N_3955,N_4295);
and U7409 (N_7409,N_4011,N_4532);
and U7410 (N_7410,N_2595,N_2891);
and U7411 (N_7411,N_4773,N_4396);
nor U7412 (N_7412,N_3030,N_3173);
nor U7413 (N_7413,N_3448,N_4765);
nand U7414 (N_7414,N_3399,N_3722);
and U7415 (N_7415,N_3324,N_3517);
nand U7416 (N_7416,N_2646,N_4950);
xnor U7417 (N_7417,N_4553,N_3917);
nand U7418 (N_7418,N_3839,N_4862);
nand U7419 (N_7419,N_2757,N_3564);
or U7420 (N_7420,N_3801,N_3911);
nand U7421 (N_7421,N_3419,N_2925);
or U7422 (N_7422,N_2862,N_4598);
xor U7423 (N_7423,N_4492,N_3460);
xor U7424 (N_7424,N_4099,N_4628);
or U7425 (N_7425,N_2684,N_4694);
and U7426 (N_7426,N_3267,N_3120);
xnor U7427 (N_7427,N_4243,N_4437);
and U7428 (N_7428,N_4341,N_3935);
and U7429 (N_7429,N_4042,N_3407);
nor U7430 (N_7430,N_4960,N_4975);
or U7431 (N_7431,N_3052,N_4116);
nand U7432 (N_7432,N_4751,N_3625);
or U7433 (N_7433,N_3374,N_4457);
nor U7434 (N_7434,N_4210,N_4720);
nand U7435 (N_7435,N_4323,N_4533);
nor U7436 (N_7436,N_3734,N_4121);
or U7437 (N_7437,N_4483,N_2660);
or U7438 (N_7438,N_4524,N_4128);
or U7439 (N_7439,N_2705,N_3691);
and U7440 (N_7440,N_2697,N_3760);
or U7441 (N_7441,N_3605,N_3273);
or U7442 (N_7442,N_3185,N_4774);
nand U7443 (N_7443,N_3349,N_4011);
or U7444 (N_7444,N_4808,N_2596);
and U7445 (N_7445,N_3755,N_2744);
nand U7446 (N_7446,N_4486,N_3692);
nand U7447 (N_7447,N_3900,N_3035);
or U7448 (N_7448,N_4106,N_2518);
and U7449 (N_7449,N_4780,N_4076);
and U7450 (N_7450,N_4039,N_2822);
nor U7451 (N_7451,N_4731,N_2547);
or U7452 (N_7452,N_4050,N_3213);
xnor U7453 (N_7453,N_2969,N_4268);
and U7454 (N_7454,N_4903,N_3568);
xnor U7455 (N_7455,N_4939,N_4123);
nand U7456 (N_7456,N_4094,N_3668);
or U7457 (N_7457,N_2782,N_3449);
or U7458 (N_7458,N_2598,N_4645);
nor U7459 (N_7459,N_4215,N_2925);
and U7460 (N_7460,N_4182,N_3648);
nor U7461 (N_7461,N_4417,N_3381);
or U7462 (N_7462,N_3063,N_3164);
and U7463 (N_7463,N_4332,N_3181);
or U7464 (N_7464,N_3573,N_4421);
and U7465 (N_7465,N_4050,N_4985);
or U7466 (N_7466,N_2787,N_4715);
and U7467 (N_7467,N_4752,N_3184);
xnor U7468 (N_7468,N_4386,N_4801);
and U7469 (N_7469,N_3159,N_3797);
or U7470 (N_7470,N_3459,N_2768);
or U7471 (N_7471,N_3599,N_2897);
or U7472 (N_7472,N_4897,N_4535);
and U7473 (N_7473,N_2538,N_2733);
nor U7474 (N_7474,N_3367,N_3399);
or U7475 (N_7475,N_4366,N_4891);
or U7476 (N_7476,N_3816,N_2743);
nand U7477 (N_7477,N_2705,N_4638);
xor U7478 (N_7478,N_3443,N_2654);
nor U7479 (N_7479,N_2697,N_3248);
nor U7480 (N_7480,N_2686,N_2854);
nor U7481 (N_7481,N_4418,N_4137);
nand U7482 (N_7482,N_4049,N_4039);
and U7483 (N_7483,N_2654,N_4705);
nand U7484 (N_7484,N_3597,N_4362);
nand U7485 (N_7485,N_2896,N_4566);
nand U7486 (N_7486,N_3840,N_4421);
and U7487 (N_7487,N_2787,N_4440);
nand U7488 (N_7488,N_4935,N_3361);
xnor U7489 (N_7489,N_2700,N_2832);
and U7490 (N_7490,N_2743,N_3100);
and U7491 (N_7491,N_4589,N_4806);
or U7492 (N_7492,N_4609,N_2957);
nor U7493 (N_7493,N_2653,N_3956);
nand U7494 (N_7494,N_4069,N_3961);
nand U7495 (N_7495,N_4097,N_2678);
nand U7496 (N_7496,N_4654,N_4307);
and U7497 (N_7497,N_2560,N_4600);
or U7498 (N_7498,N_2984,N_2535);
and U7499 (N_7499,N_4551,N_3030);
or U7500 (N_7500,N_5603,N_6029);
nor U7501 (N_7501,N_5035,N_6636);
nand U7502 (N_7502,N_5357,N_6725);
nor U7503 (N_7503,N_5042,N_5749);
or U7504 (N_7504,N_6253,N_5914);
or U7505 (N_7505,N_5919,N_6432);
and U7506 (N_7506,N_6291,N_7149);
nand U7507 (N_7507,N_6495,N_7152);
nand U7508 (N_7508,N_6184,N_6148);
and U7509 (N_7509,N_7093,N_7478);
and U7510 (N_7510,N_6706,N_6252);
nor U7511 (N_7511,N_5554,N_5187);
nand U7512 (N_7512,N_5727,N_5798);
nor U7513 (N_7513,N_5828,N_7063);
or U7514 (N_7514,N_6943,N_5496);
nand U7515 (N_7515,N_6180,N_7313);
nand U7516 (N_7516,N_5250,N_7499);
xor U7517 (N_7517,N_7332,N_5204);
nand U7518 (N_7518,N_5097,N_6624);
nor U7519 (N_7519,N_5656,N_6189);
or U7520 (N_7520,N_7166,N_6031);
or U7521 (N_7521,N_5982,N_5634);
nand U7522 (N_7522,N_7398,N_5655);
nor U7523 (N_7523,N_6425,N_6016);
nand U7524 (N_7524,N_7148,N_5251);
and U7525 (N_7525,N_6006,N_7133);
or U7526 (N_7526,N_7316,N_6849);
and U7527 (N_7527,N_7037,N_7338);
or U7528 (N_7528,N_6910,N_5908);
or U7529 (N_7529,N_7319,N_6550);
nor U7530 (N_7530,N_7119,N_7223);
nand U7531 (N_7531,N_5861,N_5882);
or U7532 (N_7532,N_6328,N_6799);
xor U7533 (N_7533,N_6632,N_5299);
or U7534 (N_7534,N_5811,N_6535);
and U7535 (N_7535,N_6571,N_5645);
nand U7536 (N_7536,N_6999,N_5781);
nand U7537 (N_7537,N_6801,N_5207);
or U7538 (N_7538,N_6674,N_5384);
nand U7539 (N_7539,N_6585,N_7365);
xnor U7540 (N_7540,N_5394,N_6883);
nor U7541 (N_7541,N_5827,N_6879);
nand U7542 (N_7542,N_7050,N_5853);
and U7543 (N_7543,N_6622,N_5627);
nor U7544 (N_7544,N_5743,N_5557);
nand U7545 (N_7545,N_5849,N_5677);
or U7546 (N_7546,N_5801,N_5964);
and U7547 (N_7547,N_6247,N_7009);
and U7548 (N_7548,N_6409,N_6465);
nand U7549 (N_7549,N_5142,N_5401);
and U7550 (N_7550,N_6234,N_7187);
and U7551 (N_7551,N_6556,N_7217);
or U7552 (N_7552,N_7011,N_7195);
nand U7553 (N_7553,N_6742,N_6317);
nor U7554 (N_7554,N_5717,N_5129);
and U7555 (N_7555,N_5376,N_5210);
nor U7556 (N_7556,N_7078,N_6603);
and U7557 (N_7557,N_6287,N_5336);
nand U7558 (N_7558,N_6797,N_6990);
and U7559 (N_7559,N_7402,N_5577);
xor U7560 (N_7560,N_5074,N_6439);
and U7561 (N_7561,N_6908,N_5807);
nand U7562 (N_7562,N_5124,N_6975);
xor U7563 (N_7563,N_6577,N_6601);
and U7564 (N_7564,N_7378,N_5578);
or U7565 (N_7565,N_5597,N_7437);
or U7566 (N_7566,N_7482,N_6055);
nor U7567 (N_7567,N_6431,N_5423);
or U7568 (N_7568,N_5747,N_5093);
nor U7569 (N_7569,N_6336,N_7264);
nor U7570 (N_7570,N_6623,N_6634);
or U7571 (N_7571,N_6829,N_6812);
and U7572 (N_7572,N_6940,N_5509);
and U7573 (N_7573,N_6030,N_6335);
nor U7574 (N_7574,N_6824,N_5347);
nor U7575 (N_7575,N_6613,N_6131);
or U7576 (N_7576,N_6348,N_7470);
nor U7577 (N_7577,N_5813,N_7479);
nor U7578 (N_7578,N_6479,N_5967);
and U7579 (N_7579,N_5199,N_5342);
nand U7580 (N_7580,N_6384,N_5815);
and U7581 (N_7581,N_6862,N_5864);
nor U7582 (N_7582,N_5147,N_7222);
and U7583 (N_7583,N_5069,N_6010);
xnor U7584 (N_7584,N_5959,N_6281);
or U7585 (N_7585,N_5773,N_6542);
and U7586 (N_7586,N_5934,N_6041);
xor U7587 (N_7587,N_6160,N_5793);
and U7588 (N_7588,N_7436,N_7370);
nor U7589 (N_7589,N_6490,N_6821);
or U7590 (N_7590,N_5200,N_5909);
and U7591 (N_7591,N_7333,N_5545);
or U7592 (N_7592,N_5650,N_5448);
or U7593 (N_7593,N_5633,N_7045);
xor U7594 (N_7594,N_6618,N_5497);
and U7595 (N_7595,N_6688,N_5283);
and U7596 (N_7596,N_6283,N_5365);
or U7597 (N_7597,N_5456,N_6173);
and U7598 (N_7598,N_5211,N_6497);
and U7599 (N_7599,N_6049,N_5024);
nor U7600 (N_7600,N_7024,N_5975);
and U7601 (N_7601,N_5198,N_5281);
and U7602 (N_7602,N_7134,N_5382);
and U7603 (N_7603,N_5078,N_6878);
and U7604 (N_7604,N_6593,N_6259);
nor U7605 (N_7605,N_7385,N_5977);
and U7606 (N_7606,N_5572,N_6566);
and U7607 (N_7607,N_6840,N_6111);
and U7608 (N_7608,N_5182,N_7128);
or U7609 (N_7609,N_5623,N_6786);
nand U7610 (N_7610,N_5540,N_6671);
or U7611 (N_7611,N_5895,N_5957);
xnor U7612 (N_7612,N_6779,N_7043);
nor U7613 (N_7613,N_6715,N_6099);
and U7614 (N_7614,N_7487,N_5296);
and U7615 (N_7615,N_6166,N_6196);
xnor U7616 (N_7616,N_5291,N_7038);
or U7617 (N_7617,N_6732,N_5167);
and U7618 (N_7618,N_5820,N_6702);
nor U7619 (N_7619,N_6302,N_7412);
or U7620 (N_7620,N_5151,N_6536);
nor U7621 (N_7621,N_5569,N_6858);
and U7622 (N_7622,N_5407,N_5141);
and U7623 (N_7623,N_5720,N_7295);
and U7624 (N_7624,N_6953,N_6164);
or U7625 (N_7625,N_5831,N_6848);
nor U7626 (N_7626,N_5966,N_6907);
nor U7627 (N_7627,N_6061,N_5945);
xor U7628 (N_7628,N_6905,N_6126);
nand U7629 (N_7629,N_5832,N_5073);
and U7630 (N_7630,N_5707,N_6755);
nand U7631 (N_7631,N_7022,N_5206);
or U7632 (N_7632,N_6417,N_5128);
and U7633 (N_7633,N_5759,N_5348);
and U7634 (N_7634,N_7254,N_6219);
nor U7635 (N_7635,N_5123,N_5009);
or U7636 (N_7636,N_6323,N_5659);
or U7637 (N_7637,N_6985,N_6653);
nand U7638 (N_7638,N_7293,N_6441);
nand U7639 (N_7639,N_6820,N_6557);
and U7640 (N_7640,N_5981,N_7253);
nor U7641 (N_7641,N_7342,N_6021);
nor U7642 (N_7642,N_5556,N_6095);
nor U7643 (N_7643,N_6500,N_6675);
or U7644 (N_7644,N_6997,N_7323);
nand U7645 (N_7645,N_6218,N_5955);
nand U7646 (N_7646,N_5121,N_6340);
nand U7647 (N_7647,N_5535,N_5332);
and U7648 (N_7648,N_7389,N_6946);
xnor U7649 (N_7649,N_5399,N_5692);
or U7650 (N_7650,N_5753,N_6169);
or U7651 (N_7651,N_7344,N_7335);
and U7652 (N_7652,N_7360,N_7079);
or U7653 (N_7653,N_5002,N_5404);
nor U7654 (N_7654,N_5192,N_6244);
nor U7655 (N_7655,N_5610,N_7170);
nand U7656 (N_7656,N_5534,N_6109);
nor U7657 (N_7657,N_6044,N_6359);
or U7658 (N_7658,N_6414,N_7320);
nor U7659 (N_7659,N_5051,N_5704);
and U7660 (N_7660,N_6691,N_7440);
nand U7661 (N_7661,N_6746,N_5880);
xor U7662 (N_7662,N_5438,N_6949);
nand U7663 (N_7663,N_5086,N_5290);
or U7664 (N_7664,N_5263,N_6969);
or U7665 (N_7665,N_6912,N_6208);
nor U7666 (N_7666,N_5653,N_6651);
or U7667 (N_7667,N_6738,N_5059);
and U7668 (N_7668,N_5089,N_5470);
nor U7669 (N_7669,N_5661,N_7445);
nand U7670 (N_7670,N_6512,N_6137);
or U7671 (N_7671,N_6664,N_6757);
nand U7672 (N_7672,N_6804,N_7294);
and U7673 (N_7673,N_5777,N_5865);
or U7674 (N_7674,N_5169,N_6619);
and U7675 (N_7675,N_6637,N_6163);
nand U7676 (N_7676,N_7248,N_6343);
nor U7677 (N_7677,N_5635,N_5092);
xnor U7678 (N_7678,N_5261,N_5023);
nor U7679 (N_7679,N_5758,N_5709);
and U7680 (N_7680,N_5277,N_5622);
and U7681 (N_7681,N_7107,N_5493);
and U7682 (N_7682,N_6312,N_6805);
and U7683 (N_7683,N_7240,N_5235);
nand U7684 (N_7684,N_6920,N_6264);
or U7685 (N_7685,N_6324,N_5276);
and U7686 (N_7686,N_5657,N_5640);
and U7687 (N_7687,N_5842,N_7064);
or U7688 (N_7688,N_7000,N_5953);
or U7689 (N_7689,N_6641,N_7065);
nand U7690 (N_7690,N_6238,N_7194);
nor U7691 (N_7691,N_6059,N_5008);
or U7692 (N_7692,N_7260,N_6043);
or U7693 (N_7693,N_5370,N_5462);
nand U7694 (N_7694,N_6373,N_6760);
or U7695 (N_7695,N_7180,N_5071);
nor U7696 (N_7696,N_6337,N_7444);
and U7697 (N_7697,N_5005,N_5028);
or U7698 (N_7698,N_6209,N_6051);
nand U7699 (N_7699,N_6352,N_6934);
or U7700 (N_7700,N_5512,N_5333);
nor U7701 (N_7701,N_5120,N_5927);
nand U7702 (N_7702,N_7363,N_5396);
nand U7703 (N_7703,N_5651,N_5736);
xnor U7704 (N_7704,N_6257,N_5504);
or U7705 (N_7705,N_6683,N_5702);
and U7706 (N_7706,N_7467,N_7446);
nand U7707 (N_7707,N_6827,N_6358);
nand U7708 (N_7708,N_6187,N_5343);
nand U7709 (N_7709,N_6696,N_6771);
or U7710 (N_7710,N_5383,N_6522);
and U7711 (N_7711,N_7307,N_7279);
nor U7712 (N_7712,N_5878,N_6455);
or U7713 (N_7713,N_6230,N_6501);
or U7714 (N_7714,N_5574,N_5271);
nor U7715 (N_7715,N_6235,N_6311);
nand U7716 (N_7716,N_5220,N_7273);
or U7717 (N_7717,N_6579,N_5551);
or U7718 (N_7718,N_7483,N_5698);
or U7719 (N_7719,N_5979,N_5676);
or U7720 (N_7720,N_7372,N_7272);
nand U7721 (N_7721,N_6182,N_7076);
nor U7722 (N_7722,N_7181,N_7464);
nor U7723 (N_7723,N_5483,N_5963);
nor U7724 (N_7724,N_5242,N_5756);
or U7725 (N_7725,N_5113,N_5033);
and U7726 (N_7726,N_5014,N_5986);
and U7727 (N_7727,N_6492,N_5782);
and U7728 (N_7728,N_6316,N_6011);
or U7729 (N_7729,N_6661,N_6047);
and U7730 (N_7730,N_7104,N_6523);
nor U7731 (N_7731,N_5745,N_5178);
nor U7732 (N_7732,N_7186,N_5951);
xnor U7733 (N_7733,N_5549,N_6525);
or U7734 (N_7734,N_5416,N_7017);
nor U7735 (N_7735,N_7085,N_6306);
nor U7736 (N_7736,N_7089,N_5428);
nor U7737 (N_7737,N_6548,N_6551);
nand U7738 (N_7738,N_6958,N_6205);
xor U7739 (N_7739,N_7314,N_6847);
and U7740 (N_7740,N_6159,N_6236);
and U7741 (N_7741,N_7377,N_6584);
or U7742 (N_7742,N_5246,N_7121);
nand U7743 (N_7743,N_6604,N_5232);
nand U7744 (N_7744,N_5592,N_7315);
nand U7745 (N_7745,N_6091,N_6605);
nand U7746 (N_7746,N_7031,N_5391);
nor U7747 (N_7747,N_6450,N_6977);
and U7748 (N_7748,N_7101,N_6890);
nor U7749 (N_7749,N_5713,N_5993);
xnor U7750 (N_7750,N_5328,N_6646);
or U7751 (N_7751,N_7484,N_5511);
nand U7752 (N_7752,N_6001,N_5475);
nor U7753 (N_7753,N_6916,N_5648);
nor U7754 (N_7754,N_5526,N_6456);
nand U7755 (N_7755,N_5525,N_5668);
nor U7756 (N_7756,N_6592,N_6193);
and U7757 (N_7757,N_5409,N_5352);
nor U7758 (N_7758,N_7206,N_6243);
and U7759 (N_7759,N_5432,N_7127);
and U7760 (N_7760,N_6489,N_5044);
xnor U7761 (N_7761,N_5329,N_5612);
nand U7762 (N_7762,N_5364,N_7238);
nor U7763 (N_7763,N_7371,N_6246);
or U7764 (N_7764,N_7156,N_6083);
nand U7765 (N_7765,N_5886,N_5703);
and U7766 (N_7766,N_5297,N_5938);
and U7767 (N_7767,N_5224,N_6058);
nor U7768 (N_7768,N_5020,N_5268);
nand U7769 (N_7769,N_5941,N_5601);
and U7770 (N_7770,N_5355,N_7459);
nand U7771 (N_7771,N_6116,N_5195);
and U7772 (N_7772,N_5602,N_5029);
and U7773 (N_7773,N_7305,N_7441);
nand U7774 (N_7774,N_5390,N_5079);
or U7775 (N_7775,N_6428,N_6533);
or U7776 (N_7776,N_6144,N_5331);
or U7777 (N_7777,N_5260,N_5395);
nor U7778 (N_7778,N_6947,N_7171);
and U7779 (N_7779,N_6297,N_6069);
and U7780 (N_7780,N_5724,N_5875);
and U7781 (N_7781,N_5122,N_5065);
nor U7782 (N_7782,N_7154,N_7334);
xnor U7783 (N_7783,N_5311,N_5792);
nand U7784 (N_7784,N_5553,N_5313);
xnor U7785 (N_7785,N_6104,N_6354);
or U7786 (N_7786,N_5607,N_5543);
nand U7787 (N_7787,N_6591,N_7391);
xor U7788 (N_7788,N_7241,N_5775);
or U7789 (N_7789,N_5523,N_7346);
or U7790 (N_7790,N_6078,N_5733);
and U7791 (N_7791,N_5244,N_5082);
or U7792 (N_7792,N_6033,N_6514);
or U7793 (N_7793,N_5295,N_5294);
nor U7794 (N_7794,N_5011,N_6830);
and U7795 (N_7795,N_6416,N_6463);
and U7796 (N_7796,N_5208,N_6057);
or U7797 (N_7797,N_5137,N_5628);
nor U7798 (N_7798,N_7161,N_5776);
or U7799 (N_7799,N_5334,N_7480);
nand U7800 (N_7800,N_7350,N_5769);
nor U7801 (N_7801,N_6188,N_7364);
and U7802 (N_7802,N_6457,N_5802);
xnor U7803 (N_7803,N_6063,N_6945);
and U7804 (N_7804,N_7120,N_6087);
or U7805 (N_7805,N_6539,N_7027);
or U7806 (N_7806,N_5726,N_6617);
and U7807 (N_7807,N_5117,N_6315);
nand U7808 (N_7808,N_5529,N_7086);
nor U7809 (N_7809,N_6784,N_5317);
or U7810 (N_7810,N_7392,N_6405);
xor U7811 (N_7811,N_5859,N_7066);
nor U7812 (N_7812,N_6660,N_6367);
or U7813 (N_7813,N_7137,N_7353);
nor U7814 (N_7814,N_5790,N_5146);
and U7815 (N_7815,N_6050,N_5976);
xor U7816 (N_7816,N_7454,N_5680);
nand U7817 (N_7817,N_6192,N_6039);
and U7818 (N_7818,N_6644,N_5422);
or U7819 (N_7819,N_6381,N_5728);
nand U7820 (N_7820,N_5643,N_6752);
or U7821 (N_7821,N_6909,N_5319);
nand U7822 (N_7822,N_6608,N_6722);
or U7823 (N_7823,N_5550,N_5960);
or U7824 (N_7824,N_5503,N_6005);
or U7825 (N_7825,N_6240,N_7111);
xor U7826 (N_7826,N_5135,N_6761);
and U7827 (N_7827,N_5388,N_7039);
or U7828 (N_7828,N_6298,N_5971);
nand U7829 (N_7829,N_6368,N_7369);
and U7830 (N_7830,N_6831,N_6615);
nand U7831 (N_7831,N_5338,N_6206);
nand U7832 (N_7832,N_7103,N_6914);
and U7833 (N_7833,N_6794,N_5708);
and U7834 (N_7834,N_7481,N_6017);
or U7835 (N_7835,N_7362,N_6642);
or U7836 (N_7836,N_6587,N_5025);
and U7837 (N_7837,N_7290,N_6911);
nor U7838 (N_7838,N_5420,N_6446);
nor U7839 (N_7839,N_6334,N_5439);
xnor U7840 (N_7840,N_5454,N_6952);
or U7841 (N_7841,N_7176,N_7390);
and U7842 (N_7842,N_6633,N_6165);
nand U7843 (N_7843,N_7282,N_6447);
and U7844 (N_7844,N_6694,N_6279);
or U7845 (N_7845,N_6103,N_6494);
and U7846 (N_7846,N_5588,N_7008);
xor U7847 (N_7847,N_6775,N_6627);
nand U7848 (N_7848,N_6024,N_6509);
xor U7849 (N_7849,N_5258,N_6009);
or U7850 (N_7850,N_6388,N_7136);
nand U7851 (N_7851,N_6881,N_7105);
and U7852 (N_7852,N_6598,N_5316);
and U7853 (N_7853,N_7173,N_5230);
and U7854 (N_7854,N_6762,N_5403);
or U7855 (N_7855,N_6275,N_7297);
and U7856 (N_7856,N_7144,N_6296);
nand U7857 (N_7857,N_6255,N_6004);
and U7858 (N_7858,N_7150,N_6519);
xor U7859 (N_7859,N_5822,N_5145);
nand U7860 (N_7860,N_7488,N_6781);
nor U7861 (N_7861,N_6555,N_5887);
and U7862 (N_7862,N_7041,N_6527);
nand U7863 (N_7863,N_7244,N_6473);
or U7864 (N_7864,N_6245,N_7496);
nand U7865 (N_7865,N_6716,N_5126);
nand U7866 (N_7866,N_6709,N_5176);
xnor U7867 (N_7867,N_5685,N_5808);
nor U7868 (N_7868,N_6353,N_6318);
nor U7869 (N_7869,N_6986,N_7061);
xor U7870 (N_7870,N_5508,N_7108);
xor U7871 (N_7871,N_7213,N_6976);
or U7872 (N_7872,N_5444,N_5196);
and U7873 (N_7873,N_5797,N_5599);
or U7874 (N_7874,N_5898,N_6552);
and U7875 (N_7875,N_7081,N_6394);
nor U7876 (N_7876,N_5153,N_6402);
nor U7877 (N_7877,N_6919,N_5314);
nand U7878 (N_7878,N_7006,N_5936);
or U7879 (N_7879,N_5445,N_7084);
or U7880 (N_7880,N_6819,N_6356);
nand U7881 (N_7881,N_6964,N_5191);
or U7882 (N_7882,N_7139,N_5515);
nand U7883 (N_7883,N_7439,N_5636);
nand U7884 (N_7884,N_5273,N_6915);
nand U7885 (N_7885,N_6177,N_6037);
nor U7886 (N_7886,N_5320,N_6770);
and U7887 (N_7887,N_7374,N_5922);
or U7888 (N_7888,N_5046,N_5965);
nor U7889 (N_7889,N_5852,N_6731);
and U7890 (N_7890,N_7280,N_5048);
nand U7891 (N_7891,N_6150,N_5030);
or U7892 (N_7892,N_6422,N_7249);
or U7893 (N_7893,N_5487,N_6669);
or U7894 (N_7894,N_5323,N_5860);
nand U7895 (N_7895,N_6857,N_7200);
and U7896 (N_7896,N_7277,N_5751);
xor U7897 (N_7897,N_6565,N_6475);
and U7898 (N_7898,N_6429,N_6493);
and U7899 (N_7899,N_6504,N_6136);
and U7900 (N_7900,N_6032,N_6682);
or U7901 (N_7901,N_7020,N_6773);
xnor U7902 (N_7902,N_6948,N_6939);
and U7903 (N_7903,N_5996,N_6151);
or U7904 (N_7904,N_7347,N_5559);
or U7905 (N_7905,N_5590,N_6719);
nor U7906 (N_7906,N_5162,N_5893);
and U7907 (N_7907,N_5339,N_5871);
nand U7908 (N_7908,N_6506,N_6075);
nand U7909 (N_7909,N_5414,N_6226);
nand U7910 (N_7910,N_5841,N_6376);
nand U7911 (N_7911,N_6530,N_7267);
nor U7912 (N_7912,N_6942,N_7339);
and U7913 (N_7913,N_6684,N_5737);
nand U7914 (N_7914,N_6053,N_7151);
or U7915 (N_7915,N_5215,N_6657);
nand U7916 (N_7916,N_5609,N_5595);
nor U7917 (N_7917,N_6411,N_5638);
xor U7918 (N_7918,N_5858,N_5083);
or U7919 (N_7919,N_6341,N_7400);
or U7920 (N_7920,N_5202,N_6290);
nor U7921 (N_7921,N_5900,N_6461);
or U7922 (N_7922,N_7055,N_5763);
nor U7923 (N_7923,N_6221,N_5476);
or U7924 (N_7924,N_6581,N_5731);
nand U7925 (N_7925,N_5754,N_5541);
nand U7926 (N_7926,N_6503,N_7417);
nand U7927 (N_7927,N_6711,N_5181);
nor U7928 (N_7928,N_6896,N_7474);
nor U7929 (N_7929,N_6129,N_6120);
and U7930 (N_7930,N_5940,N_5946);
or U7931 (N_7931,N_7189,N_5041);
nand U7932 (N_7932,N_6629,N_5868);
and U7933 (N_7933,N_7211,N_5318);
xnor U7934 (N_7934,N_5378,N_5359);
or U7935 (N_7935,N_5873,N_5999);
nand U7936 (N_7936,N_6442,N_6270);
or U7937 (N_7937,N_5434,N_6887);
and U7938 (N_7938,N_5696,N_5765);
and U7939 (N_7939,N_5649,N_6028);
and U7940 (N_7940,N_5995,N_7491);
nor U7941 (N_7941,N_5621,N_7415);
or U7942 (N_7942,N_5571,N_6899);
nand U7943 (N_7943,N_5386,N_7199);
nand U7944 (N_7944,N_5016,N_5506);
and U7945 (N_7945,N_6654,N_7147);
nor U7946 (N_7946,N_5062,N_5642);
nor U7947 (N_7947,N_5278,N_6080);
nand U7948 (N_7948,N_6124,N_6586);
nand U7949 (N_7949,N_6190,N_7367);
and U7950 (N_7950,N_6237,N_5288);
and U7951 (N_7951,N_5134,N_7435);
and U7952 (N_7952,N_6232,N_6987);
nor U7953 (N_7953,N_5102,N_6751);
or U7954 (N_7954,N_5920,N_5788);
nand U7955 (N_7955,N_5767,N_7092);
nor U7956 (N_7956,N_6876,N_7427);
and U7957 (N_7957,N_5690,N_6718);
nor U7958 (N_7958,N_5618,N_5824);
nor U7959 (N_7959,N_6267,N_7208);
nor U7960 (N_7960,N_5315,N_6485);
nor U7961 (N_7961,N_6139,N_7406);
nand U7962 (N_7962,N_6970,N_5091);
or U7963 (N_7963,N_6285,N_6607);
nor U7964 (N_7964,N_6650,N_6885);
xnor U7965 (N_7965,N_5589,N_6640);
or U7966 (N_7966,N_7115,N_7138);
and U7967 (N_7967,N_6766,N_6596);
xor U7968 (N_7968,N_5087,N_6470);
nor U7969 (N_7969,N_5784,N_6998);
xnor U7970 (N_7970,N_6228,N_5249);
nand U7971 (N_7971,N_6480,N_6498);
nor U7972 (N_7972,N_7431,N_6092);
or U7973 (N_7973,N_7197,N_5983);
nor U7974 (N_7974,N_7410,N_6564);
or U7975 (N_7975,N_5679,N_5287);
and U7976 (N_7976,N_6902,N_5490);
nor U7977 (N_7977,N_7308,N_6540);
nand U7978 (N_7978,N_6765,N_7351);
and U7979 (N_7979,N_6085,N_7049);
xnor U7980 (N_7980,N_6145,N_7287);
nor U7981 (N_7981,N_5639,N_6927);
or U7982 (N_7982,N_6396,N_6710);
or U7983 (N_7983,N_6906,N_6965);
nand U7984 (N_7984,N_6677,N_6346);
nand U7985 (N_7985,N_6146,N_6496);
nor U7986 (N_7986,N_5568,N_5712);
nand U7987 (N_7987,N_7384,N_5233);
nand U7988 (N_7988,N_6630,N_5531);
or U7989 (N_7989,N_5750,N_5884);
or U7990 (N_7990,N_5505,N_6865);
xor U7991 (N_7991,N_6476,N_6515);
nand U7992 (N_7992,N_6127,N_7257);
and U7993 (N_7993,N_6904,N_6866);
nand U7994 (N_7994,N_6748,N_6410);
xnor U7995 (N_7995,N_5174,N_6265);
or U7996 (N_7996,N_7330,N_5410);
or U7997 (N_7997,N_5039,N_7358);
xor U7998 (N_7998,N_5757,N_7227);
nand U7999 (N_7999,N_7232,N_6981);
nand U8000 (N_8000,N_5746,N_7207);
nor U8001 (N_8001,N_6486,N_5632);
nor U8002 (N_8002,N_5143,N_7091);
nand U8003 (N_8003,N_5562,N_7096);
xnor U8004 (N_8004,N_7341,N_7221);
nand U8005 (N_8005,N_7060,N_5771);
and U8006 (N_8006,N_5442,N_7386);
or U8007 (N_8007,N_5166,N_5050);
nand U8008 (N_8008,N_5671,N_5103);
nor U8009 (N_8009,N_6806,N_6599);
nand U8010 (N_8010,N_5214,N_7422);
nand U8011 (N_8011,N_5904,N_5265);
nand U8012 (N_8012,N_7449,N_6991);
nand U8013 (N_8013,N_5748,N_6851);
nor U8014 (N_8014,N_7265,N_6303);
nand U8015 (N_8015,N_6074,N_6957);
nand U8016 (N_8016,N_7419,N_7250);
nor U8017 (N_8017,N_5611,N_5243);
nor U8018 (N_8018,N_5544,N_6777);
xnor U8019 (N_8019,N_5575,N_7465);
nand U8020 (N_8020,N_7463,N_7396);
nand U8021 (N_8021,N_5459,N_5040);
or U8022 (N_8022,N_7196,N_6167);
nor U8023 (N_8023,N_5561,N_5385);
or U8024 (N_8024,N_6213,N_7345);
nor U8025 (N_8025,N_5138,N_7070);
and U8026 (N_8026,N_5026,N_5430);
nor U8027 (N_8027,N_5652,N_6926);
and U8028 (N_8028,N_6435,N_5108);
and U8029 (N_8029,N_6117,N_6382);
or U8030 (N_8030,N_6156,N_5453);
xnor U8031 (N_8031,N_5673,N_7302);
nand U8032 (N_8032,N_7340,N_6778);
nand U8033 (N_8033,N_7274,N_5901);
xor U8034 (N_8034,N_5840,N_7193);
and U8035 (N_8035,N_6045,N_6951);
nor U8036 (N_8036,N_6096,N_5095);
nand U8037 (N_8037,N_6231,N_5156);
nor U8038 (N_8038,N_7116,N_6407);
xnor U8039 (N_8039,N_6520,N_6048);
nor U8040 (N_8040,N_6220,N_6241);
nor U8041 (N_8041,N_6813,N_5667);
or U8042 (N_8042,N_5105,N_5337);
and U8043 (N_8043,N_6448,N_6606);
and U8044 (N_8044,N_6764,N_6121);
and U8045 (N_8045,N_7432,N_5604);
xor U8046 (N_8046,N_6133,N_6466);
nand U8047 (N_8047,N_6672,N_6505);
nor U8048 (N_8048,N_7420,N_6638);
and U8049 (N_8049,N_6153,N_5915);
and U8050 (N_8050,N_6294,N_5471);
nand U8051 (N_8051,N_5565,N_5043);
nor U8052 (N_8052,N_6843,N_6673);
or U8053 (N_8053,N_6125,N_5458);
xor U8054 (N_8054,N_7472,N_6304);
and U8055 (N_8055,N_6389,N_5560);
nand U8056 (N_8056,N_5310,N_5038);
nand U8057 (N_8057,N_7243,N_6850);
or U8058 (N_8058,N_7209,N_6750);
and U8059 (N_8059,N_7141,N_6293);
or U8060 (N_8060,N_5817,N_6454);
and U8061 (N_8061,N_6793,N_6477);
nand U8062 (N_8062,N_6143,N_5440);
nand U8063 (N_8063,N_6481,N_6787);
nor U8064 (N_8064,N_7284,N_6903);
nand U8065 (N_8065,N_6329,N_5854);
nand U8066 (N_8066,N_6880,N_6714);
and U8067 (N_8067,N_6007,N_5697);
or U8068 (N_8068,N_6783,N_5158);
and U8069 (N_8069,N_6079,N_6225);
and U8070 (N_8070,N_7322,N_5241);
nand U8071 (N_8071,N_5354,N_6274);
nand U8072 (N_8072,N_7130,N_7382);
and U8073 (N_8073,N_6838,N_5755);
or U8074 (N_8074,N_6983,N_7292);
nand U8075 (N_8075,N_5335,N_5032);
and U8076 (N_8076,N_6543,N_5835);
or U8077 (N_8077,N_5566,N_5057);
and U8078 (N_8078,N_5721,N_6443);
and U8079 (N_8079,N_5441,N_6361);
nand U8080 (N_8080,N_5876,N_6737);
nand U8081 (N_8081,N_6576,N_7035);
or U8082 (N_8082,N_7067,N_5286);
and U8083 (N_8083,N_6772,N_6802);
nand U8084 (N_8084,N_6689,N_5184);
nand U8085 (N_8085,N_6172,N_6898);
or U8086 (N_8086,N_6583,N_5163);
nand U8087 (N_8087,N_5877,N_7443);
and U8088 (N_8088,N_6464,N_7004);
xor U8089 (N_8089,N_5061,N_7106);
or U8090 (N_8090,N_6362,N_5903);
nand U8091 (N_8091,N_5699,N_6413);
nand U8092 (N_8092,N_7160,N_6073);
or U8093 (N_8093,N_7082,N_6269);
nand U8094 (N_8094,N_6614,N_7113);
xnor U8095 (N_8095,N_6484,N_5764);
nand U8096 (N_8096,N_7220,N_7143);
nor U8097 (N_8097,N_5109,N_6963);
nand U8098 (N_8098,N_5942,N_6286);
xnor U8099 (N_8099,N_5034,N_5171);
and U8100 (N_8100,N_5485,N_5906);
and U8101 (N_8101,N_5932,N_5950);
nand U8102 (N_8102,N_6474,N_6836);
and U8103 (N_8103,N_5015,N_6272);
nor U8104 (N_8104,N_5888,N_5587);
or U8105 (N_8105,N_5170,N_5716);
nor U8106 (N_8106,N_6989,N_6929);
nor U8107 (N_8107,N_7188,N_7460);
or U8108 (N_8108,N_7185,N_5845);
nor U8109 (N_8109,N_5264,N_5608);
nor U8110 (N_8110,N_5252,N_7118);
and U8111 (N_8111,N_5010,N_6399);
or U8112 (N_8112,N_6186,N_5688);
nand U8113 (N_8113,N_6008,N_7015);
and U8114 (N_8114,N_5447,N_7018);
or U8115 (N_8115,N_7033,N_6098);
nand U8116 (N_8116,N_7495,N_6152);
nand U8117 (N_8117,N_7395,N_6891);
nand U8118 (N_8118,N_6808,N_5267);
nand U8119 (N_8119,N_7424,N_5047);
and U8120 (N_8120,N_6444,N_5658);
and U8121 (N_8121,N_7318,N_5361);
nand U8122 (N_8122,N_7457,N_5558);
or U8123 (N_8123,N_7215,N_6863);
nor U8124 (N_8124,N_6483,N_6322);
nand U8125 (N_8125,N_7214,N_6421);
or U8126 (N_8126,N_6157,N_6502);
and U8127 (N_8127,N_6810,N_6181);
nor U8128 (N_8128,N_5896,N_7205);
or U8129 (N_8129,N_7485,N_5855);
nand U8130 (N_8130,N_5725,N_7190);
nand U8131 (N_8131,N_5691,N_5466);
or U8132 (N_8132,N_7468,N_7283);
or U8133 (N_8133,N_7140,N_5341);
nand U8134 (N_8134,N_5076,N_7256);
or U8135 (N_8135,N_7126,N_6321);
nor U8136 (N_8136,N_6698,N_6871);
or U8137 (N_8137,N_5848,N_5257);
nor U8138 (N_8138,N_5522,N_5114);
nor U8139 (N_8139,N_7281,N_5136);
or U8140 (N_8140,N_7239,N_5785);
nor U8141 (N_8141,N_5766,N_5507);
or U8142 (N_8142,N_5274,N_5400);
xor U8143 (N_8143,N_6768,N_6134);
nand U8144 (N_8144,N_6666,N_5806);
nor U8145 (N_8145,N_7321,N_5881);
nor U8146 (N_8146,N_6625,N_6511);
nand U8147 (N_8147,N_6162,N_5734);
nor U8148 (N_8148,N_6488,N_5446);
nor U8149 (N_8149,N_5973,N_7356);
nor U8150 (N_8150,N_7047,N_5826);
or U8151 (N_8151,N_5066,N_5307);
nand U8152 (N_8152,N_5968,N_5226);
nand U8153 (N_8153,N_5096,N_5894);
and U8154 (N_8154,N_7229,N_6776);
or U8155 (N_8155,N_5972,N_6835);
nand U8156 (N_8156,N_6852,N_5054);
nor U8157 (N_8157,N_5270,N_7179);
nand U8158 (N_8158,N_6420,N_6419);
and U8159 (N_8159,N_5256,N_6655);
nor U8160 (N_8160,N_5660,N_7021);
nor U8161 (N_8161,N_7252,N_7354);
nand U8162 (N_8162,N_5664,N_5001);
or U8163 (N_8163,N_6357,N_6580);
nand U8164 (N_8164,N_5863,N_6194);
or U8165 (N_8165,N_5431,N_7379);
nand U8166 (N_8166,N_6728,N_5177);
xor U8167 (N_8167,N_5457,N_5923);
and U8168 (N_8168,N_6355,N_5952);
and U8169 (N_8169,N_7309,N_5408);
nor U8170 (N_8170,N_5866,N_6211);
nand U8171 (N_8171,N_7010,N_5521);
nor U8172 (N_8172,N_5846,N_7486);
nand U8173 (N_8173,N_5730,N_7278);
xor U8174 (N_8174,N_5131,N_6788);
nor U8175 (N_8175,N_5990,N_5678);
nand U8176 (N_8176,N_6678,N_5197);
or U8177 (N_8177,N_6708,N_5988);
nand U8178 (N_8178,N_6263,N_5829);
or U8179 (N_8179,N_7097,N_5060);
nand U8180 (N_8180,N_5693,N_6130);
xnor U8181 (N_8181,N_6081,N_6401);
nand U8182 (N_8182,N_6954,N_6663);
and U8183 (N_8183,N_6872,N_5536);
nand U8184 (N_8184,N_7473,N_5682);
and U8185 (N_8185,N_7132,N_6217);
and U8186 (N_8186,N_6936,N_6168);
or U8187 (N_8187,N_6686,N_6140);
nor U8188 (N_8188,N_5579,N_6561);
nand U8189 (N_8189,N_6308,N_7030);
nor U8190 (N_8190,N_7304,N_5212);
nor U8191 (N_8191,N_7411,N_5080);
or U8192 (N_8192,N_6300,N_5222);
nand U8193 (N_8193,N_6962,N_5930);
nand U8194 (N_8194,N_6224,N_6562);
and U8195 (N_8195,N_6482,N_5489);
or U8196 (N_8196,N_7327,N_7425);
or U8197 (N_8197,N_5292,N_6563);
nand U8198 (N_8198,N_6097,N_5794);
and U8199 (N_8199,N_7122,N_6700);
or U8200 (N_8200,N_5426,N_6392);
and U8201 (N_8201,N_7230,N_7336);
nand U8202 (N_8202,N_7456,N_6380);
nand U8203 (N_8203,N_7178,N_5107);
and U8204 (N_8204,N_5814,N_5351);
and U8205 (N_8205,N_5237,N_7489);
or U8206 (N_8206,N_5686,N_5427);
nand U8207 (N_8207,N_6273,N_5072);
or U8208 (N_8208,N_5449,N_6889);
or U8209 (N_8209,N_5053,N_5998);
nor U8210 (N_8210,N_7032,N_6631);
or U8211 (N_8211,N_7476,N_6400);
and U8212 (N_8212,N_6982,N_6278);
nor U8213 (N_8213,N_6467,N_6518);
nand U8214 (N_8214,N_6873,N_7475);
xnor U8215 (N_8215,N_5718,N_5464);
or U8216 (N_8216,N_5644,N_6753);
nor U8217 (N_8217,N_5654,N_5027);
and U8218 (N_8218,N_5219,N_6724);
or U8219 (N_8219,N_6877,N_5897);
and U8220 (N_8220,N_7450,N_6106);
and U8221 (N_8221,N_7216,N_5672);
and U8222 (N_8222,N_5662,N_5168);
nand U8223 (N_8223,N_5312,N_5018);
nand U8224 (N_8224,N_5481,N_6035);
xor U8225 (N_8225,N_7163,N_7157);
nor U8226 (N_8226,N_7234,N_5081);
nor U8227 (N_8227,N_5706,N_6438);
nor U8228 (N_8228,N_5947,N_5463);
and U8229 (N_8229,N_6289,N_5929);
or U8230 (N_8230,N_6854,N_5978);
nand U8231 (N_8231,N_5115,N_7416);
nand U8232 (N_8232,N_5874,N_5474);
and U8233 (N_8233,N_5804,N_5101);
and U8234 (N_8234,N_5477,N_6460);
nand U8235 (N_8235,N_6171,N_5254);
xnor U8236 (N_8236,N_5741,N_5436);
nand U8237 (N_8237,N_5537,N_5381);
and U8238 (N_8238,N_6178,N_6993);
nand U8239 (N_8239,N_7080,N_7044);
or U8240 (N_8240,N_6309,N_6101);
nor U8241 (N_8241,N_6391,N_6925);
nor U8242 (N_8242,N_5624,N_7331);
xor U8243 (N_8243,N_5799,N_5593);
and U8244 (N_8244,N_6423,N_5567);
or U8245 (N_8245,N_5402,N_6090);
or U8246 (N_8246,N_5637,N_7426);
and U8247 (N_8247,N_6730,N_6612);
nand U8248 (N_8248,N_7025,N_7383);
nand U8249 (N_8249,N_6726,N_5774);
nor U8250 (N_8250,N_5787,N_6928);
and U8251 (N_8251,N_5349,N_7068);
and U8252 (N_8252,N_6602,N_6349);
nor U8253 (N_8253,N_5161,N_5705);
xor U8254 (N_8254,N_5580,N_5293);
and U8255 (N_8255,N_5847,N_7202);
and U8256 (N_8256,N_5284,N_7310);
nor U8257 (N_8257,N_6248,N_5253);
xnor U8258 (N_8258,N_6478,N_6076);
xor U8259 (N_8259,N_6108,N_5594);
nor U8260 (N_8260,N_6817,N_7268);
and U8261 (N_8261,N_7159,N_5094);
nor U8262 (N_8262,N_5450,N_6841);
nor U8263 (N_8263,N_6690,N_6344);
nand U8264 (N_8264,N_6200,N_6754);
or U8265 (N_8265,N_5694,N_6521);
and U8266 (N_8266,N_5600,N_5012);
xor U8267 (N_8267,N_7042,N_5417);
and U8268 (N_8268,N_5068,N_7014);
nand U8269 (N_8269,N_6800,N_5205);
nand U8270 (N_8270,N_6900,N_6935);
nand U8271 (N_8271,N_5324,N_6002);
and U8272 (N_8272,N_5280,N_6310);
nand U8273 (N_8273,N_6138,N_6692);
and U8274 (N_8274,N_6364,N_6679);
nor U8275 (N_8275,N_6427,N_5377);
or U8276 (N_8276,N_6094,N_7404);
and U8277 (N_8277,N_6922,N_6544);
nand U8278 (N_8278,N_7433,N_6616);
and U8279 (N_8279,N_5918,N_6471);
and U8280 (N_8280,N_6763,N_7237);
and U8281 (N_8281,N_7145,N_6780);
nor U8282 (N_8282,N_6901,N_5714);
nand U8283 (N_8283,N_6393,N_7114);
or U8284 (N_8284,N_6767,N_6207);
nor U8285 (N_8285,N_5467,N_5954);
and U8286 (N_8286,N_5225,N_7359);
nand U8287 (N_8287,N_6216,N_6743);
nand U8288 (N_8288,N_5533,N_5548);
or U8289 (N_8289,N_5985,N_5371);
and U8290 (N_8290,N_5492,N_6842);
nand U8291 (N_8291,N_5889,N_5465);
nand U8292 (N_8292,N_6553,N_6326);
xnor U8293 (N_8293,N_7451,N_6398);
or U8294 (N_8294,N_6036,N_7407);
or U8295 (N_8295,N_5674,N_5149);
and U8296 (N_8296,N_6620,N_7183);
and U8297 (N_8297,N_6662,N_6268);
and U8298 (N_8298,N_7071,N_5372);
and U8299 (N_8299,N_5902,N_7129);
nor U8300 (N_8300,N_5563,N_7447);
nor U8301 (N_8301,N_6796,N_5221);
nor U8302 (N_8302,N_7158,N_6967);
nand U8303 (N_8303,N_5380,N_6575);
nor U8304 (N_8304,N_6534,N_6212);
nor U8305 (N_8305,N_5524,N_5913);
nor U8306 (N_8306,N_7286,N_5369);
nand U8307 (N_8307,N_7349,N_5494);
or U8308 (N_8308,N_6437,N_6175);
nand U8309 (N_8309,N_5017,N_5304);
or U8310 (N_8310,N_6332,N_6918);
nor U8311 (N_8311,N_6258,N_7036);
or U8312 (N_8312,N_7124,N_6424);
or U8313 (N_8313,N_6508,N_5879);
nor U8314 (N_8314,N_5098,N_7403);
xor U8315 (N_8315,N_6020,N_6345);
nand U8316 (N_8316,N_6086,N_6023);
and U8317 (N_8317,N_7090,N_7430);
and U8318 (N_8318,N_5616,N_5321);
and U8319 (N_8319,N_5004,N_6837);
and U8320 (N_8320,N_6699,N_6060);
and U8321 (N_8321,N_6517,N_5987);
and U8322 (N_8322,N_6210,N_6284);
nand U8323 (N_8323,N_6734,N_5173);
nand U8324 (N_8324,N_5683,N_5830);
or U8325 (N_8325,N_6288,N_6703);
nor U8326 (N_8326,N_6531,N_7083);
nor U8327 (N_8327,N_5980,N_7285);
xor U8328 (N_8328,N_7329,N_6342);
and U8329 (N_8329,N_6893,N_6973);
and U8330 (N_8330,N_6590,N_5160);
or U8331 (N_8331,N_5596,N_5742);
xnor U8332 (N_8332,N_5796,N_7026);
and U8333 (N_8333,N_6792,N_5738);
nand U8334 (N_8334,N_6695,N_5255);
nand U8335 (N_8335,N_6064,N_5266);
or U8336 (N_8336,N_6833,N_6227);
and U8337 (N_8337,N_7259,N_5127);
nand U8338 (N_8338,N_6874,N_5598);
or U8339 (N_8339,N_5112,N_7380);
xnor U8340 (N_8340,N_5193,N_5305);
nand U8341 (N_8341,N_6147,N_6803);
nor U8342 (N_8342,N_7153,N_6014);
nor U8343 (N_8343,N_6370,N_5373);
nand U8344 (N_8344,N_7458,N_6701);
xor U8345 (N_8345,N_6070,N_5867);
and U8346 (N_8346,N_6301,N_5387);
nand U8347 (N_8347,N_6717,N_5739);
nor U8348 (N_8348,N_6524,N_7052);
and U8349 (N_8349,N_5921,N_5928);
and U8350 (N_8350,N_5301,N_6541);
nor U8351 (N_8351,N_5605,N_7172);
nand U8352 (N_8352,N_7434,N_6077);
nor U8353 (N_8353,N_5375,N_7023);
nand U8354 (N_8354,N_6680,N_5539);
or U8355 (N_8355,N_5231,N_5300);
nor U8356 (N_8356,N_6249,N_6733);
and U8357 (N_8357,N_6179,N_5912);
nand U8358 (N_8358,N_5768,N_6972);
and U8359 (N_8359,N_6434,N_6676);
or U8360 (N_8360,N_7224,N_5869);
nand U8361 (N_8361,N_6740,N_5397);
and U8362 (N_8362,N_6685,N_5106);
or U8363 (N_8363,N_6327,N_7123);
nand U8364 (N_8364,N_7165,N_6875);
nand U8365 (N_8365,N_6649,N_6113);
and U8366 (N_8366,N_6383,N_5910);
xnor U8367 (N_8367,N_5989,N_7393);
nand U8368 (N_8368,N_6128,N_6068);
nand U8369 (N_8369,N_5948,N_6363);
and U8370 (N_8370,N_6377,N_7058);
or U8371 (N_8371,N_5130,N_5582);
and U8372 (N_8372,N_5547,N_5891);
nor U8373 (N_8373,N_6229,N_7219);
or U8374 (N_8374,N_6114,N_7262);
or U8375 (N_8375,N_7461,N_5905);
nor U8376 (N_8376,N_5723,N_5856);
nor U8377 (N_8377,N_6966,N_5500);
nor U8378 (N_8378,N_6491,N_6736);
and U8379 (N_8379,N_5021,N_7448);
nand U8380 (N_8380,N_5478,N_5007);
nor U8381 (N_8381,N_5234,N_6529);
and U8382 (N_8382,N_6729,N_5665);
nor U8383 (N_8383,N_5045,N_5970);
nor U8384 (N_8384,N_5180,N_7087);
nand U8385 (N_8385,N_5625,N_5272);
xor U8386 (N_8386,N_7002,N_5837);
nor U8387 (N_8387,N_7112,N_7210);
or U8388 (N_8388,N_6727,N_5259);
and U8389 (N_8389,N_5302,N_6735);
nand U8390 (N_8390,N_5488,N_6320);
or U8391 (N_8391,N_6994,N_7201);
or U8392 (N_8392,N_6313,N_5778);
nand U8393 (N_8393,N_6594,N_7174);
or U8394 (N_8394,N_5552,N_6436);
xnor U8395 (N_8395,N_6578,N_5345);
or U8396 (N_8396,N_5172,N_7296);
and U8397 (N_8397,N_5519,N_6012);
xnor U8398 (N_8398,N_5099,N_5502);
nor U8399 (N_8399,N_5189,N_5116);
or U8400 (N_8400,N_6924,N_5433);
and U8401 (N_8401,N_6499,N_5368);
nor U8402 (N_8402,N_6971,N_5479);
nor U8403 (N_8403,N_7303,N_5825);
nor U8404 (N_8404,N_6822,N_5363);
nand U8405 (N_8405,N_5984,N_6921);
nor U8406 (N_8406,N_5125,N_6658);
and U8407 (N_8407,N_7413,N_5614);
or U8408 (N_8408,N_7494,N_6239);
nand U8409 (N_8409,N_5424,N_7266);
and U8410 (N_8410,N_7034,N_7007);
and U8411 (N_8411,N_6628,N_6198);
and U8412 (N_8412,N_6119,N_6704);
nand U8413 (N_8413,N_5937,N_5836);
or U8414 (N_8414,N_6795,N_6547);
nand U8415 (N_8415,N_5056,N_7326);
nand U8416 (N_8416,N_5326,N_6870);
and U8417 (N_8417,N_6042,N_5870);
nand U8418 (N_8418,N_6387,N_6360);
and U8419 (N_8419,N_5289,N_7438);
or U8420 (N_8420,N_5501,N_6798);
or U8421 (N_8421,N_5538,N_5821);
nand U8422 (N_8422,N_5935,N_6894);
nand U8423 (N_8423,N_6532,N_6826);
and U8424 (N_8424,N_7233,N_6365);
nand U8425 (N_8425,N_7387,N_6065);
nor U8426 (N_8426,N_6818,N_5356);
nand U8427 (N_8427,N_5236,N_5843);
nor U8428 (N_8428,N_5527,N_7046);
or U8429 (N_8429,N_7263,N_6462);
or U8430 (N_8430,N_6330,N_7301);
nand U8431 (N_8431,N_6056,N_7477);
or U8432 (N_8432,N_5070,N_6811);
or U8433 (N_8433,N_6067,N_5358);
nor U8434 (N_8434,N_7236,N_5228);
and U8435 (N_8435,N_7312,N_7493);
nand U8436 (N_8436,N_5405,N_5367);
nand U8437 (N_8437,N_5063,N_5415);
and U8438 (N_8438,N_5911,N_5647);
and U8439 (N_8439,N_5631,N_7054);
nand U8440 (N_8440,N_5322,N_5013);
or U8441 (N_8441,N_6888,N_6088);
or U8442 (N_8442,N_6687,N_5418);
and U8443 (N_8443,N_6950,N_6018);
nand U8444 (N_8444,N_5992,N_5425);
nand U8445 (N_8445,N_5997,N_6626);
nor U8446 (N_8446,N_6271,N_6155);
xor U8447 (N_8447,N_5949,N_6331);
nand U8448 (N_8448,N_6262,N_6510);
nand U8449 (N_8449,N_5795,N_6333);
nand U8450 (N_8450,N_5974,N_6516);
nand U8451 (N_8451,N_6445,N_7469);
and U8452 (N_8452,N_6745,N_5818);
nand U8453 (N_8453,N_6807,N_6572);
nor U8454 (N_8454,N_6559,N_7271);
nand U8455 (N_8455,N_5803,N_5513);
nand U8456 (N_8456,N_6897,N_6537);
and U8457 (N_8457,N_7317,N_7247);
and U8458 (N_8458,N_6412,N_5067);
nor U8459 (N_8459,N_5393,N_6276);
nor U8460 (N_8460,N_5058,N_6647);
xor U8461 (N_8461,N_7357,N_5719);
and U8462 (N_8462,N_5772,N_6756);
and U8463 (N_8463,N_5800,N_7228);
nand U8464 (N_8464,N_6197,N_5711);
nand U8465 (N_8465,N_7098,N_6720);
nor U8466 (N_8466,N_5217,N_7013);
nand U8467 (N_8467,N_6084,N_5100);
nand U8468 (N_8468,N_6453,N_6656);
xor U8469 (N_8469,N_6351,N_5780);
and U8470 (N_8470,N_6513,N_6440);
nor U8471 (N_8471,N_5770,N_7376);
nor U8472 (N_8472,N_6853,N_5584);
or U8473 (N_8473,N_6823,N_6869);
and U8474 (N_8474,N_7348,N_5591);
nor U8475 (N_8475,N_5689,N_6621);
nand U8476 (N_8476,N_5546,N_6741);
and U8477 (N_8477,N_7325,N_5555);
nand U8478 (N_8478,N_5366,N_5353);
nor U8479 (N_8479,N_5629,N_7408);
and U8480 (N_8480,N_7255,N_5885);
nand U8481 (N_8481,N_6390,N_6941);
nor U8482 (N_8482,N_5482,N_5729);
nor U8483 (N_8483,N_5480,N_6378);
nor U8484 (N_8484,N_5245,N_6595);
nand U8485 (N_8485,N_6828,N_6379);
and U8486 (N_8486,N_5360,N_6215);
nor U8487 (N_8487,N_5419,N_7299);
and U8488 (N_8488,N_5443,N_7077);
nor U8489 (N_8489,N_5762,N_5451);
nand U8490 (N_8490,N_6149,N_5944);
or U8491 (N_8491,N_7168,N_6809);
xnor U8492 (N_8492,N_5209,N_6789);
nor U8493 (N_8493,N_7110,N_6214);
or U8494 (N_8494,N_7352,N_6707);
and U8495 (N_8495,N_6895,N_6082);
nand U8496 (N_8496,N_6046,N_5460);
nor U8497 (N_8497,N_7048,N_6667);
and U8498 (N_8498,N_5406,N_5486);
and U8499 (N_8499,N_7289,N_5003);
or U8500 (N_8500,N_5308,N_5899);
or U8501 (N_8501,N_5710,N_6135);
nor U8502 (N_8502,N_7095,N_5530);
or U8503 (N_8503,N_6859,N_7062);
xor U8504 (N_8504,N_6176,N_5084);
and U8505 (N_8505,N_5943,N_6917);
nand U8506 (N_8506,N_7019,N_5484);
xor U8507 (N_8507,N_7270,N_7074);
and U8508 (N_8508,N_6526,N_5851);
or U8509 (N_8509,N_6093,N_7231);
nand U8510 (N_8510,N_6174,N_5695);
and U8511 (N_8511,N_6668,N_6299);
nor U8512 (N_8512,N_5350,N_5247);
nand U8513 (N_8513,N_5389,N_6546);
nand U8514 (N_8514,N_5344,N_6856);
and U8515 (N_8515,N_7428,N_6892);
and U8516 (N_8516,N_6978,N_7375);
or U8517 (N_8517,N_6122,N_6223);
xnor U8518 (N_8518,N_6832,N_5285);
nor U8519 (N_8519,N_7429,N_6825);
xnor U8520 (N_8520,N_5190,N_6314);
or U8521 (N_8521,N_5783,N_5991);
and U8522 (N_8522,N_5646,N_5133);
or U8523 (N_8523,N_6325,N_6956);
xnor U8524 (N_8524,N_5227,N_6112);
or U8525 (N_8525,N_5049,N_5429);
nor U8526 (N_8526,N_5340,N_6816);
nand U8527 (N_8527,N_6415,N_6886);
and U8528 (N_8528,N_6705,N_6589);
and U8529 (N_8529,N_5392,N_5619);
xor U8530 (N_8530,N_7072,N_5085);
nand U8531 (N_8531,N_6062,N_5185);
and U8532 (N_8532,N_5779,N_5617);
or U8533 (N_8533,N_5186,N_6102);
and U8534 (N_8534,N_7421,N_6123);
or U8535 (N_8535,N_5684,N_7040);
nand U8536 (N_8536,N_6974,N_7275);
or U8537 (N_8537,N_6665,N_6403);
or U8538 (N_8538,N_5528,N_6000);
and U8539 (N_8539,N_7169,N_5179);
nand U8540 (N_8540,N_5468,N_6697);
xor U8541 (N_8541,N_6459,N_5298);
nand U8542 (N_8542,N_5006,N_5132);
or U8543 (N_8543,N_6659,N_6026);
nand U8544 (N_8544,N_6774,N_5398);
nand U8545 (N_8545,N_6242,N_6712);
or U8546 (N_8546,N_6574,N_5346);
xnor U8547 (N_8547,N_6744,N_6961);
and U8548 (N_8548,N_7056,N_5715);
or U8549 (N_8549,N_5201,N_6884);
nand U8550 (N_8550,N_7490,N_5229);
nor U8551 (N_8551,N_5670,N_5961);
and U8552 (N_8552,N_5675,N_5140);
nand U8553 (N_8553,N_5000,N_5740);
nor U8554 (N_8554,N_7051,N_7191);
xnor U8555 (N_8555,N_5844,N_7261);
and U8556 (N_8556,N_7235,N_5437);
or U8557 (N_8557,N_7497,N_5435);
or U8558 (N_8558,N_5088,N_6996);
nor U8559 (N_8559,N_5064,N_6713);
or U8560 (N_8560,N_7498,N_6758);
xnor U8561 (N_8561,N_5994,N_6645);
nand U8562 (N_8562,N_6968,N_6937);
and U8563 (N_8563,N_5154,N_7399);
nand U8564 (N_8564,N_7401,N_7251);
nand U8565 (N_8565,N_5520,N_6054);
nor U8566 (N_8566,N_6022,N_5838);
nor U8567 (N_8567,N_6643,N_6089);
and U8568 (N_8568,N_6860,N_5262);
or U8569 (N_8569,N_7311,N_5761);
nand U8570 (N_8570,N_5279,N_5119);
nor U8571 (N_8571,N_6375,N_7337);
and U8572 (N_8572,N_6027,N_6385);
nor U8573 (N_8573,N_6118,N_7102);
or U8574 (N_8574,N_6115,N_6834);
xor U8575 (N_8575,N_6339,N_5223);
nand U8576 (N_8576,N_7167,N_6487);
nor U8577 (N_8577,N_6203,N_5542);
nand U8578 (N_8578,N_6013,N_5732);
nand U8579 (N_8579,N_7146,N_6988);
or U8580 (N_8580,N_5857,N_5532);
nor U8581 (N_8581,N_6307,N_5564);
nand U8582 (N_8582,N_5789,N_6468);
nor U8583 (N_8583,N_7269,N_5570);
and U8584 (N_8584,N_7099,N_5819);
nand U8585 (N_8585,N_7028,N_7455);
xnor U8586 (N_8586,N_7069,N_6204);
nor U8587 (N_8587,N_5630,N_5883);
nand U8588 (N_8588,N_6992,N_6959);
and U8589 (N_8589,N_5152,N_5917);
nor U8590 (N_8590,N_7075,N_6979);
or U8591 (N_8591,N_6195,N_5282);
or U8592 (N_8592,N_5238,N_5306);
or U8593 (N_8593,N_6280,N_5275);
nand U8594 (N_8594,N_5461,N_6110);
nor U8595 (N_8595,N_7100,N_6072);
nand U8596 (N_8596,N_5681,N_7276);
and U8597 (N_8597,N_7324,N_6635);
nand U8598 (N_8598,N_5722,N_6256);
or U8599 (N_8599,N_6569,N_6791);
or U8600 (N_8600,N_6845,N_6199);
or U8601 (N_8601,N_5812,N_5956);
nor U8602 (N_8602,N_5239,N_6251);
xor U8603 (N_8603,N_6844,N_5890);
nand U8604 (N_8604,N_6639,N_5744);
nor U8605 (N_8605,N_6185,N_6611);
nand U8606 (N_8606,N_5218,N_5330);
xnor U8607 (N_8607,N_5150,N_6406);
or U8608 (N_8608,N_6749,N_6350);
nand U8609 (N_8609,N_7016,N_5452);
nor U8610 (N_8610,N_6132,N_7361);
and U8611 (N_8611,N_5491,N_5805);
xor U8612 (N_8612,N_5752,N_6923);
nand U8613 (N_8613,N_6449,N_6739);
and U8614 (N_8614,N_6944,N_6292);
and U8615 (N_8615,N_7462,N_7005);
xnor U8616 (N_8616,N_7218,N_7300);
nand U8617 (N_8617,N_6610,N_6282);
nand U8618 (N_8618,N_6769,N_6408);
nand U8619 (N_8619,N_7203,N_6538);
nor U8620 (N_8620,N_6932,N_5248);
xnor U8621 (N_8621,N_6052,N_5666);
and U8622 (N_8622,N_5183,N_5669);
or U8623 (N_8623,N_5892,N_6960);
and U8624 (N_8624,N_6570,N_7094);
nand U8625 (N_8625,N_6105,N_5413);
or U8626 (N_8626,N_6670,N_6588);
or U8627 (N_8627,N_5175,N_6864);
and U8628 (N_8628,N_5019,N_5157);
or U8629 (N_8629,N_5816,N_5309);
and U8630 (N_8630,N_5498,N_7226);
nand U8631 (N_8631,N_5926,N_7204);
xor U8632 (N_8632,N_5194,N_5586);
or U8633 (N_8633,N_7466,N_6451);
nand U8634 (N_8634,N_5075,N_7471);
or U8635 (N_8635,N_7291,N_7184);
nor U8636 (N_8636,N_6980,N_5118);
or U8637 (N_8637,N_7057,N_6558);
nor U8638 (N_8638,N_5495,N_5925);
nor U8639 (N_8639,N_5469,N_6938);
or U8640 (N_8640,N_7328,N_5620);
xor U8641 (N_8641,N_7492,N_5613);
and U8642 (N_8642,N_7177,N_5421);
nor U8643 (N_8643,N_7088,N_6161);
and U8644 (N_8644,N_5510,N_6142);
and U8645 (N_8645,N_5472,N_5090);
nor U8646 (N_8646,N_5823,N_6573);
and U8647 (N_8647,N_5022,N_6855);
nand U8648 (N_8648,N_5810,N_7109);
nor U8649 (N_8649,N_5916,N_6652);
nand U8650 (N_8650,N_5833,N_7012);
nor U8651 (N_8651,N_6426,N_7164);
nand U8652 (N_8652,N_6430,N_6846);
and U8653 (N_8653,N_6759,N_6790);
nand U8654 (N_8654,N_5924,N_6040);
nor U8655 (N_8655,N_5809,N_5412);
xnor U8656 (N_8656,N_6681,N_6261);
and U8657 (N_8657,N_7198,N_6418);
and U8658 (N_8658,N_6071,N_6395);
nand U8659 (N_8659,N_5939,N_5907);
and U8660 (N_8660,N_6597,N_6868);
nor U8661 (N_8661,N_6233,N_7288);
or U8662 (N_8662,N_6183,N_6984);
or U8663 (N_8663,N_6721,N_5188);
xor U8664 (N_8664,N_5110,N_6545);
and U8665 (N_8665,N_5327,N_5641);
or U8666 (N_8666,N_6038,N_7373);
nand U8667 (N_8667,N_5144,N_7155);
or U8668 (N_8668,N_6723,N_6995);
and U8669 (N_8669,N_7182,N_6782);
nor U8670 (N_8670,N_5036,N_5052);
xor U8671 (N_8671,N_6154,N_5687);
nor U8672 (N_8672,N_6191,N_7059);
or U8673 (N_8673,N_5933,N_5159);
and U8674 (N_8674,N_6609,N_7117);
or U8675 (N_8675,N_6366,N_6913);
nand U8676 (N_8676,N_5862,N_6347);
and U8677 (N_8677,N_5735,N_6250);
xor U8678 (N_8678,N_5269,N_6338);
and U8679 (N_8679,N_7125,N_5213);
nor U8680 (N_8680,N_5663,N_5077);
or U8681 (N_8681,N_7355,N_5031);
nor U8682 (N_8682,N_5615,N_6469);
nor U8683 (N_8683,N_7306,N_6019);
nand U8684 (N_8684,N_7175,N_6600);
and U8685 (N_8685,N_6277,N_5581);
nand U8686 (N_8686,N_6568,N_6305);
nand U8687 (N_8687,N_7142,N_6861);
nand U8688 (N_8688,N_6371,N_7135);
or U8689 (N_8689,N_5969,N_5139);
nor U8690 (N_8690,N_7073,N_6882);
and U8691 (N_8691,N_6025,N_5362);
nand U8692 (N_8692,N_6404,N_5240);
or U8693 (N_8693,N_5962,N_7242);
or U8694 (N_8694,N_6158,N_6567);
nor U8695 (N_8695,N_6201,N_6066);
nor U8696 (N_8696,N_5931,N_6170);
and U8697 (N_8697,N_6582,N_7053);
nand U8698 (N_8698,N_7131,N_5411);
or U8699 (N_8699,N_6319,N_5791);
and U8700 (N_8700,N_5583,N_6867);
or U8701 (N_8701,N_7343,N_7409);
nor U8702 (N_8702,N_5055,N_5325);
and U8703 (N_8703,N_7192,N_5760);
nor U8704 (N_8704,N_6458,N_5379);
or U8705 (N_8705,N_7368,N_7418);
nor U8706 (N_8706,N_6003,N_6785);
nor U8707 (N_8707,N_6372,N_7442);
or U8708 (N_8708,N_5701,N_5958);
nor U8709 (N_8709,N_5516,N_7452);
or U8710 (N_8710,N_6141,N_5104);
and U8711 (N_8711,N_6528,N_6554);
and U8712 (N_8712,N_6260,N_6266);
nor U8713 (N_8713,N_5203,N_5700);
or U8714 (N_8714,N_5517,N_6955);
and U8715 (N_8715,N_6472,N_5514);
and U8716 (N_8716,N_6814,N_6747);
or U8717 (N_8717,N_7246,N_5164);
or U8718 (N_8718,N_5037,N_6560);
nor U8719 (N_8719,N_5850,N_5165);
nand U8720 (N_8720,N_6100,N_7029);
nor U8721 (N_8721,N_6386,N_6549);
or U8722 (N_8722,N_7212,N_6933);
nor U8723 (N_8723,N_5455,N_7414);
nand U8724 (N_8724,N_6648,N_7388);
xor U8725 (N_8725,N_6015,N_5786);
or U8726 (N_8726,N_6254,N_5148);
or U8727 (N_8727,N_5303,N_7298);
and U8728 (N_8728,N_7394,N_5473);
and U8729 (N_8729,N_7245,N_6202);
or U8730 (N_8730,N_6839,N_6222);
xor U8731 (N_8731,N_6034,N_7405);
nor U8732 (N_8732,N_6295,N_7453);
and U8733 (N_8733,N_7001,N_6433);
or U8734 (N_8734,N_6397,N_6930);
or U8735 (N_8735,N_6107,N_6369);
xnor U8736 (N_8736,N_7423,N_7397);
and U8737 (N_8737,N_7162,N_7003);
or U8738 (N_8738,N_5626,N_5374);
nand U8739 (N_8739,N_6931,N_5518);
nand U8740 (N_8740,N_7381,N_6507);
nor U8741 (N_8741,N_5606,N_5155);
nor U8742 (N_8742,N_7225,N_5111);
xnor U8743 (N_8743,N_6815,N_7258);
nand U8744 (N_8744,N_5872,N_5585);
nand U8745 (N_8745,N_5839,N_5834);
nand U8746 (N_8746,N_7366,N_5576);
or U8747 (N_8747,N_5573,N_5499);
nor U8748 (N_8748,N_6452,N_6374);
nor U8749 (N_8749,N_6693,N_5216);
and U8750 (N_8750,N_6461,N_5661);
and U8751 (N_8751,N_5833,N_5761);
nor U8752 (N_8752,N_5567,N_6481);
nor U8753 (N_8753,N_6135,N_5234);
or U8754 (N_8754,N_6165,N_5064);
nand U8755 (N_8755,N_5102,N_6817);
xor U8756 (N_8756,N_5440,N_5315);
or U8757 (N_8757,N_5646,N_5299);
or U8758 (N_8758,N_5264,N_5976);
or U8759 (N_8759,N_5087,N_6909);
nand U8760 (N_8760,N_5076,N_5884);
nor U8761 (N_8761,N_5845,N_5797);
and U8762 (N_8762,N_7240,N_5486);
nand U8763 (N_8763,N_6766,N_6188);
nor U8764 (N_8764,N_6239,N_6956);
nand U8765 (N_8765,N_5284,N_7006);
nand U8766 (N_8766,N_5382,N_5568);
nor U8767 (N_8767,N_5893,N_5921);
xnor U8768 (N_8768,N_6341,N_5150);
or U8769 (N_8769,N_5220,N_6571);
nand U8770 (N_8770,N_7080,N_5223);
or U8771 (N_8771,N_7359,N_5341);
and U8772 (N_8772,N_6520,N_6536);
or U8773 (N_8773,N_6763,N_7346);
or U8774 (N_8774,N_6891,N_5010);
nand U8775 (N_8775,N_5171,N_6183);
nor U8776 (N_8776,N_6059,N_6612);
and U8777 (N_8777,N_5840,N_5777);
and U8778 (N_8778,N_5238,N_5360);
and U8779 (N_8779,N_6300,N_5867);
xnor U8780 (N_8780,N_6316,N_5862);
nor U8781 (N_8781,N_7198,N_5254);
nand U8782 (N_8782,N_6864,N_5590);
nor U8783 (N_8783,N_6676,N_5202);
nor U8784 (N_8784,N_7310,N_6198);
nor U8785 (N_8785,N_6615,N_5986);
or U8786 (N_8786,N_7461,N_5445);
or U8787 (N_8787,N_6463,N_5218);
and U8788 (N_8788,N_6784,N_5197);
xor U8789 (N_8789,N_6917,N_5549);
xnor U8790 (N_8790,N_6466,N_6314);
and U8791 (N_8791,N_5217,N_6752);
nand U8792 (N_8792,N_6245,N_6719);
xor U8793 (N_8793,N_5351,N_5555);
xnor U8794 (N_8794,N_5615,N_6399);
or U8795 (N_8795,N_5035,N_7053);
nor U8796 (N_8796,N_5038,N_6693);
nor U8797 (N_8797,N_7258,N_5642);
nand U8798 (N_8798,N_6009,N_7384);
nand U8799 (N_8799,N_6363,N_6021);
nand U8800 (N_8800,N_5789,N_6453);
nor U8801 (N_8801,N_5644,N_6864);
nor U8802 (N_8802,N_6345,N_6931);
nand U8803 (N_8803,N_6442,N_7383);
nand U8804 (N_8804,N_6396,N_6718);
and U8805 (N_8805,N_5809,N_5892);
nand U8806 (N_8806,N_5065,N_7032);
or U8807 (N_8807,N_6080,N_5073);
nand U8808 (N_8808,N_6170,N_6928);
nor U8809 (N_8809,N_7033,N_5214);
nand U8810 (N_8810,N_5209,N_6873);
nor U8811 (N_8811,N_5501,N_5813);
nand U8812 (N_8812,N_5916,N_6353);
or U8813 (N_8813,N_6247,N_6008);
and U8814 (N_8814,N_5599,N_5948);
nand U8815 (N_8815,N_7165,N_5397);
nand U8816 (N_8816,N_6640,N_5411);
or U8817 (N_8817,N_5741,N_6915);
or U8818 (N_8818,N_6654,N_6832);
or U8819 (N_8819,N_5380,N_5292);
nor U8820 (N_8820,N_7206,N_6927);
or U8821 (N_8821,N_6111,N_5517);
nand U8822 (N_8822,N_6466,N_5343);
nand U8823 (N_8823,N_5011,N_6413);
nand U8824 (N_8824,N_5704,N_5982);
nand U8825 (N_8825,N_7487,N_7184);
and U8826 (N_8826,N_6912,N_7409);
xor U8827 (N_8827,N_5283,N_5150);
nand U8828 (N_8828,N_6773,N_5387);
nand U8829 (N_8829,N_5404,N_5378);
nor U8830 (N_8830,N_6647,N_5845);
nand U8831 (N_8831,N_5688,N_7343);
xnor U8832 (N_8832,N_5886,N_6121);
or U8833 (N_8833,N_5430,N_5792);
xnor U8834 (N_8834,N_6476,N_6027);
and U8835 (N_8835,N_5470,N_6726);
nor U8836 (N_8836,N_5257,N_5104);
or U8837 (N_8837,N_7067,N_6129);
nor U8838 (N_8838,N_7394,N_7395);
xnor U8839 (N_8839,N_5186,N_6862);
nor U8840 (N_8840,N_6970,N_7115);
xor U8841 (N_8841,N_5326,N_7085);
nor U8842 (N_8842,N_7037,N_5425);
or U8843 (N_8843,N_6492,N_6069);
or U8844 (N_8844,N_5430,N_7273);
nand U8845 (N_8845,N_5851,N_5492);
and U8846 (N_8846,N_5565,N_7357);
and U8847 (N_8847,N_6913,N_5152);
nand U8848 (N_8848,N_6604,N_7096);
and U8849 (N_8849,N_6190,N_6936);
xor U8850 (N_8850,N_6723,N_5555);
and U8851 (N_8851,N_6492,N_6515);
and U8852 (N_8852,N_7359,N_5355);
or U8853 (N_8853,N_5657,N_7137);
nand U8854 (N_8854,N_5344,N_6080);
or U8855 (N_8855,N_6927,N_5948);
or U8856 (N_8856,N_5127,N_5067);
and U8857 (N_8857,N_7334,N_6784);
and U8858 (N_8858,N_5513,N_6497);
nor U8859 (N_8859,N_5385,N_5420);
nor U8860 (N_8860,N_7161,N_7013);
xnor U8861 (N_8861,N_7207,N_5077);
or U8862 (N_8862,N_6336,N_7106);
or U8863 (N_8863,N_6945,N_7094);
or U8864 (N_8864,N_7164,N_5870);
nor U8865 (N_8865,N_6773,N_5526);
nor U8866 (N_8866,N_5453,N_6169);
xnor U8867 (N_8867,N_6290,N_7269);
and U8868 (N_8868,N_7154,N_6880);
nand U8869 (N_8869,N_5859,N_7027);
nand U8870 (N_8870,N_6513,N_6059);
nand U8871 (N_8871,N_5509,N_5618);
or U8872 (N_8872,N_5721,N_5618);
or U8873 (N_8873,N_5477,N_6892);
nand U8874 (N_8874,N_6977,N_7040);
nor U8875 (N_8875,N_5550,N_7494);
nor U8876 (N_8876,N_7144,N_5399);
or U8877 (N_8877,N_6427,N_5279);
or U8878 (N_8878,N_6661,N_5546);
nand U8879 (N_8879,N_6794,N_6966);
and U8880 (N_8880,N_5412,N_6237);
or U8881 (N_8881,N_6882,N_6738);
or U8882 (N_8882,N_5822,N_5805);
or U8883 (N_8883,N_5500,N_7100);
nand U8884 (N_8884,N_6601,N_5649);
nand U8885 (N_8885,N_5798,N_5838);
or U8886 (N_8886,N_6841,N_5316);
or U8887 (N_8887,N_5293,N_5125);
nor U8888 (N_8888,N_6622,N_6156);
and U8889 (N_8889,N_5599,N_6285);
xor U8890 (N_8890,N_7116,N_6304);
nor U8891 (N_8891,N_5689,N_7425);
or U8892 (N_8892,N_6521,N_7240);
and U8893 (N_8893,N_6475,N_5381);
xnor U8894 (N_8894,N_7170,N_5438);
or U8895 (N_8895,N_5069,N_7361);
and U8896 (N_8896,N_7330,N_7198);
or U8897 (N_8897,N_5480,N_7312);
and U8898 (N_8898,N_6277,N_7071);
xnor U8899 (N_8899,N_5775,N_5140);
nor U8900 (N_8900,N_5769,N_6218);
nor U8901 (N_8901,N_6096,N_6536);
and U8902 (N_8902,N_5336,N_7407);
or U8903 (N_8903,N_7178,N_5571);
or U8904 (N_8904,N_5800,N_7189);
and U8905 (N_8905,N_6547,N_6314);
or U8906 (N_8906,N_6090,N_7094);
or U8907 (N_8907,N_5082,N_6402);
xnor U8908 (N_8908,N_5858,N_5969);
nand U8909 (N_8909,N_5462,N_6050);
or U8910 (N_8910,N_6159,N_6948);
nor U8911 (N_8911,N_6497,N_7211);
and U8912 (N_8912,N_6143,N_7076);
and U8913 (N_8913,N_6076,N_5216);
nand U8914 (N_8914,N_5889,N_5739);
nor U8915 (N_8915,N_6508,N_6480);
and U8916 (N_8916,N_5121,N_5716);
or U8917 (N_8917,N_5153,N_6090);
nand U8918 (N_8918,N_6481,N_6468);
and U8919 (N_8919,N_6041,N_5781);
and U8920 (N_8920,N_5079,N_5738);
and U8921 (N_8921,N_5184,N_5435);
or U8922 (N_8922,N_5046,N_6335);
nor U8923 (N_8923,N_6496,N_6968);
or U8924 (N_8924,N_6172,N_5704);
and U8925 (N_8925,N_5494,N_6273);
and U8926 (N_8926,N_6721,N_5659);
or U8927 (N_8927,N_5047,N_7356);
and U8928 (N_8928,N_6600,N_6913);
or U8929 (N_8929,N_5942,N_6804);
nand U8930 (N_8930,N_7240,N_6466);
and U8931 (N_8931,N_5956,N_5275);
or U8932 (N_8932,N_7093,N_5531);
nor U8933 (N_8933,N_5650,N_5293);
and U8934 (N_8934,N_5085,N_6043);
or U8935 (N_8935,N_5311,N_6744);
nand U8936 (N_8936,N_6584,N_6566);
and U8937 (N_8937,N_7284,N_6212);
xor U8938 (N_8938,N_6465,N_5163);
nand U8939 (N_8939,N_6602,N_6391);
or U8940 (N_8940,N_6598,N_6439);
nand U8941 (N_8941,N_6674,N_6029);
and U8942 (N_8942,N_6267,N_5681);
nor U8943 (N_8943,N_7152,N_5987);
nor U8944 (N_8944,N_6020,N_6835);
nor U8945 (N_8945,N_5866,N_6151);
and U8946 (N_8946,N_6628,N_5792);
nand U8947 (N_8947,N_5450,N_5160);
and U8948 (N_8948,N_6912,N_6414);
nor U8949 (N_8949,N_5334,N_7415);
or U8950 (N_8950,N_5513,N_7334);
nor U8951 (N_8951,N_7049,N_5840);
or U8952 (N_8952,N_5577,N_5505);
or U8953 (N_8953,N_7465,N_7253);
or U8954 (N_8954,N_6462,N_6293);
nand U8955 (N_8955,N_6767,N_6721);
or U8956 (N_8956,N_5018,N_6392);
nand U8957 (N_8957,N_6493,N_5821);
or U8958 (N_8958,N_6881,N_6959);
and U8959 (N_8959,N_6473,N_5372);
nor U8960 (N_8960,N_7156,N_6898);
and U8961 (N_8961,N_6256,N_5871);
or U8962 (N_8962,N_5695,N_5759);
nor U8963 (N_8963,N_6179,N_6050);
and U8964 (N_8964,N_5341,N_7351);
or U8965 (N_8965,N_7206,N_6802);
nand U8966 (N_8966,N_5791,N_6256);
and U8967 (N_8967,N_5691,N_5017);
and U8968 (N_8968,N_5027,N_5348);
and U8969 (N_8969,N_7201,N_5892);
and U8970 (N_8970,N_6989,N_6833);
or U8971 (N_8971,N_7231,N_5950);
nor U8972 (N_8972,N_7241,N_5241);
or U8973 (N_8973,N_7174,N_6677);
nand U8974 (N_8974,N_6696,N_6297);
nand U8975 (N_8975,N_5431,N_6778);
or U8976 (N_8976,N_5889,N_6316);
nand U8977 (N_8977,N_7073,N_7272);
xnor U8978 (N_8978,N_6924,N_6947);
nor U8979 (N_8979,N_6975,N_5818);
nand U8980 (N_8980,N_5367,N_7235);
nor U8981 (N_8981,N_6496,N_5304);
xor U8982 (N_8982,N_5514,N_5058);
and U8983 (N_8983,N_6454,N_7192);
and U8984 (N_8984,N_6621,N_5729);
or U8985 (N_8985,N_6202,N_5543);
nor U8986 (N_8986,N_7191,N_6758);
nand U8987 (N_8987,N_5758,N_6775);
and U8988 (N_8988,N_5782,N_6008);
nand U8989 (N_8989,N_6711,N_5215);
nand U8990 (N_8990,N_5525,N_6853);
nand U8991 (N_8991,N_5694,N_7407);
nand U8992 (N_8992,N_6194,N_6129);
or U8993 (N_8993,N_5484,N_7205);
xnor U8994 (N_8994,N_7244,N_7083);
or U8995 (N_8995,N_6663,N_6356);
nor U8996 (N_8996,N_7017,N_6779);
nor U8997 (N_8997,N_5770,N_6270);
and U8998 (N_8998,N_6300,N_6442);
nand U8999 (N_8999,N_6321,N_5993);
and U9000 (N_9000,N_7252,N_6397);
nor U9001 (N_9001,N_5333,N_5987);
nand U9002 (N_9002,N_6579,N_5270);
nand U9003 (N_9003,N_6566,N_6911);
nor U9004 (N_9004,N_6225,N_5985);
or U9005 (N_9005,N_5376,N_5546);
or U9006 (N_9006,N_6133,N_6339);
nand U9007 (N_9007,N_7291,N_6428);
nor U9008 (N_9008,N_6235,N_7110);
nand U9009 (N_9009,N_5571,N_6102);
and U9010 (N_9010,N_6711,N_7269);
or U9011 (N_9011,N_7414,N_5955);
nand U9012 (N_9012,N_6776,N_5032);
and U9013 (N_9013,N_6268,N_6197);
nand U9014 (N_9014,N_6633,N_5028);
nand U9015 (N_9015,N_7483,N_5797);
and U9016 (N_9016,N_7359,N_6559);
nor U9017 (N_9017,N_6553,N_6323);
nor U9018 (N_9018,N_6712,N_6599);
or U9019 (N_9019,N_5196,N_5439);
nor U9020 (N_9020,N_7161,N_6873);
or U9021 (N_9021,N_6377,N_7089);
or U9022 (N_9022,N_7059,N_5454);
nor U9023 (N_9023,N_6468,N_5903);
xnor U9024 (N_9024,N_5609,N_6617);
and U9025 (N_9025,N_7362,N_6906);
and U9026 (N_9026,N_5077,N_6669);
nand U9027 (N_9027,N_6716,N_5601);
or U9028 (N_9028,N_7094,N_6888);
nand U9029 (N_9029,N_5016,N_5015);
xor U9030 (N_9030,N_5346,N_6868);
nor U9031 (N_9031,N_7284,N_5824);
nand U9032 (N_9032,N_6279,N_6102);
nand U9033 (N_9033,N_6507,N_5238);
and U9034 (N_9034,N_6375,N_6838);
xor U9035 (N_9035,N_5522,N_6897);
xor U9036 (N_9036,N_7240,N_5375);
and U9037 (N_9037,N_5380,N_5242);
nor U9038 (N_9038,N_6271,N_6611);
nor U9039 (N_9039,N_7485,N_6171);
nor U9040 (N_9040,N_7166,N_7117);
nor U9041 (N_9041,N_6923,N_6687);
or U9042 (N_9042,N_5475,N_6570);
and U9043 (N_9043,N_5308,N_5866);
and U9044 (N_9044,N_6151,N_6105);
nand U9045 (N_9045,N_5618,N_5946);
or U9046 (N_9046,N_5350,N_5082);
xor U9047 (N_9047,N_6162,N_5118);
nand U9048 (N_9048,N_5744,N_6346);
nand U9049 (N_9049,N_5268,N_5720);
nor U9050 (N_9050,N_6206,N_6131);
and U9051 (N_9051,N_6612,N_7280);
nand U9052 (N_9052,N_7452,N_5938);
and U9053 (N_9053,N_6490,N_5123);
nor U9054 (N_9054,N_5220,N_6410);
and U9055 (N_9055,N_6827,N_6047);
or U9056 (N_9056,N_5749,N_7351);
or U9057 (N_9057,N_7151,N_7115);
or U9058 (N_9058,N_5681,N_6559);
and U9059 (N_9059,N_5993,N_5285);
and U9060 (N_9060,N_6316,N_5610);
nand U9061 (N_9061,N_7130,N_5925);
and U9062 (N_9062,N_5529,N_6998);
nor U9063 (N_9063,N_6196,N_7024);
or U9064 (N_9064,N_5738,N_6045);
and U9065 (N_9065,N_6468,N_5319);
and U9066 (N_9066,N_6808,N_6629);
xnor U9067 (N_9067,N_6011,N_7127);
nor U9068 (N_9068,N_5856,N_6740);
nor U9069 (N_9069,N_5298,N_5655);
and U9070 (N_9070,N_6395,N_5174);
nor U9071 (N_9071,N_6623,N_5524);
nand U9072 (N_9072,N_6272,N_6860);
nor U9073 (N_9073,N_6575,N_5494);
nand U9074 (N_9074,N_6900,N_6068);
and U9075 (N_9075,N_7329,N_6727);
or U9076 (N_9076,N_5685,N_6343);
nor U9077 (N_9077,N_6374,N_6029);
nand U9078 (N_9078,N_7497,N_6599);
nand U9079 (N_9079,N_5554,N_5208);
and U9080 (N_9080,N_7328,N_5201);
and U9081 (N_9081,N_5902,N_7013);
or U9082 (N_9082,N_7271,N_7337);
nor U9083 (N_9083,N_6458,N_6485);
and U9084 (N_9084,N_5483,N_7312);
and U9085 (N_9085,N_6016,N_6053);
and U9086 (N_9086,N_6989,N_6585);
nand U9087 (N_9087,N_5560,N_5232);
and U9088 (N_9088,N_6480,N_5413);
nand U9089 (N_9089,N_5007,N_6080);
nor U9090 (N_9090,N_5590,N_6878);
and U9091 (N_9091,N_7318,N_6566);
or U9092 (N_9092,N_6815,N_7297);
and U9093 (N_9093,N_6170,N_5613);
xor U9094 (N_9094,N_6330,N_5523);
nand U9095 (N_9095,N_5714,N_5163);
and U9096 (N_9096,N_5229,N_5771);
nand U9097 (N_9097,N_5207,N_6889);
xor U9098 (N_9098,N_7235,N_5676);
nor U9099 (N_9099,N_6048,N_5135);
nor U9100 (N_9100,N_6142,N_6464);
xor U9101 (N_9101,N_6845,N_5988);
or U9102 (N_9102,N_5564,N_5651);
nand U9103 (N_9103,N_7095,N_5641);
nand U9104 (N_9104,N_5063,N_5011);
nand U9105 (N_9105,N_5616,N_6670);
and U9106 (N_9106,N_5743,N_6812);
or U9107 (N_9107,N_5820,N_6991);
and U9108 (N_9108,N_7017,N_6602);
nor U9109 (N_9109,N_5299,N_7424);
or U9110 (N_9110,N_6401,N_6354);
nand U9111 (N_9111,N_7288,N_5586);
xnor U9112 (N_9112,N_7379,N_5335);
nor U9113 (N_9113,N_5464,N_6235);
nand U9114 (N_9114,N_5349,N_6116);
xnor U9115 (N_9115,N_5688,N_7479);
nand U9116 (N_9116,N_5426,N_5172);
or U9117 (N_9117,N_7126,N_5409);
and U9118 (N_9118,N_6356,N_6785);
or U9119 (N_9119,N_6166,N_5779);
and U9120 (N_9120,N_6478,N_5565);
nor U9121 (N_9121,N_6349,N_5565);
nor U9122 (N_9122,N_7029,N_5822);
xor U9123 (N_9123,N_5836,N_5199);
and U9124 (N_9124,N_7403,N_6022);
nor U9125 (N_9125,N_5954,N_5403);
nand U9126 (N_9126,N_5535,N_5980);
nor U9127 (N_9127,N_6043,N_6201);
xor U9128 (N_9128,N_6652,N_7304);
xor U9129 (N_9129,N_5427,N_7115);
and U9130 (N_9130,N_7346,N_6760);
nand U9131 (N_9131,N_6458,N_6379);
nor U9132 (N_9132,N_5524,N_5886);
or U9133 (N_9133,N_5256,N_5952);
nand U9134 (N_9134,N_7262,N_6566);
xnor U9135 (N_9135,N_6384,N_6929);
nand U9136 (N_9136,N_6915,N_6787);
nand U9137 (N_9137,N_5351,N_6288);
or U9138 (N_9138,N_5479,N_5279);
or U9139 (N_9139,N_7250,N_6302);
nor U9140 (N_9140,N_7188,N_5115);
and U9141 (N_9141,N_6879,N_7071);
and U9142 (N_9142,N_7353,N_6033);
nand U9143 (N_9143,N_5212,N_6187);
and U9144 (N_9144,N_5468,N_5632);
nand U9145 (N_9145,N_5587,N_5925);
nor U9146 (N_9146,N_7198,N_6517);
nand U9147 (N_9147,N_7376,N_5603);
and U9148 (N_9148,N_7136,N_6849);
and U9149 (N_9149,N_5747,N_6928);
and U9150 (N_9150,N_5011,N_6515);
xor U9151 (N_9151,N_6903,N_6264);
nand U9152 (N_9152,N_5351,N_7172);
and U9153 (N_9153,N_6764,N_7305);
nand U9154 (N_9154,N_5989,N_5638);
or U9155 (N_9155,N_6174,N_7110);
and U9156 (N_9156,N_6974,N_7207);
nor U9157 (N_9157,N_6266,N_6965);
nand U9158 (N_9158,N_7131,N_6200);
nand U9159 (N_9159,N_6922,N_5926);
or U9160 (N_9160,N_5205,N_5636);
nor U9161 (N_9161,N_5623,N_7381);
nor U9162 (N_9162,N_6893,N_5074);
and U9163 (N_9163,N_5708,N_5766);
and U9164 (N_9164,N_7291,N_6382);
nand U9165 (N_9165,N_6328,N_7319);
or U9166 (N_9166,N_7459,N_7469);
nand U9167 (N_9167,N_6615,N_5332);
nand U9168 (N_9168,N_7215,N_7355);
or U9169 (N_9169,N_6121,N_5124);
and U9170 (N_9170,N_7386,N_7319);
and U9171 (N_9171,N_5032,N_5008);
and U9172 (N_9172,N_5881,N_6076);
and U9173 (N_9173,N_6394,N_6073);
nand U9174 (N_9174,N_5416,N_5666);
and U9175 (N_9175,N_5540,N_5861);
nor U9176 (N_9176,N_6009,N_6033);
and U9177 (N_9177,N_6677,N_5522);
nand U9178 (N_9178,N_6817,N_6870);
nand U9179 (N_9179,N_5598,N_6208);
and U9180 (N_9180,N_5103,N_5322);
and U9181 (N_9181,N_5168,N_6787);
nand U9182 (N_9182,N_5457,N_6543);
nor U9183 (N_9183,N_5918,N_6296);
or U9184 (N_9184,N_5643,N_7228);
xor U9185 (N_9185,N_5101,N_7090);
nand U9186 (N_9186,N_7046,N_6580);
and U9187 (N_9187,N_7235,N_6195);
and U9188 (N_9188,N_5192,N_6863);
and U9189 (N_9189,N_6357,N_7250);
nor U9190 (N_9190,N_6956,N_6169);
and U9191 (N_9191,N_6404,N_6186);
or U9192 (N_9192,N_6295,N_6410);
nand U9193 (N_9193,N_7461,N_6352);
or U9194 (N_9194,N_5613,N_7401);
or U9195 (N_9195,N_6700,N_7486);
nor U9196 (N_9196,N_6402,N_6127);
xnor U9197 (N_9197,N_5506,N_5101);
or U9198 (N_9198,N_6398,N_5157);
nor U9199 (N_9199,N_6902,N_7130);
or U9200 (N_9200,N_6056,N_5515);
nand U9201 (N_9201,N_6811,N_7364);
nand U9202 (N_9202,N_7023,N_6039);
nor U9203 (N_9203,N_5568,N_7333);
and U9204 (N_9204,N_5271,N_6395);
and U9205 (N_9205,N_6199,N_7308);
nand U9206 (N_9206,N_5385,N_7208);
or U9207 (N_9207,N_6707,N_5364);
xnor U9208 (N_9208,N_6140,N_7104);
or U9209 (N_9209,N_6866,N_7186);
nor U9210 (N_9210,N_6906,N_6385);
or U9211 (N_9211,N_6103,N_6269);
nor U9212 (N_9212,N_5593,N_6271);
nor U9213 (N_9213,N_6658,N_6668);
and U9214 (N_9214,N_5521,N_7268);
nand U9215 (N_9215,N_5307,N_5938);
xnor U9216 (N_9216,N_6339,N_5567);
or U9217 (N_9217,N_6430,N_6929);
nor U9218 (N_9218,N_6219,N_6994);
nor U9219 (N_9219,N_7132,N_7144);
and U9220 (N_9220,N_6606,N_6895);
or U9221 (N_9221,N_7310,N_5762);
or U9222 (N_9222,N_6921,N_6724);
nor U9223 (N_9223,N_6651,N_6349);
nand U9224 (N_9224,N_6618,N_5079);
nand U9225 (N_9225,N_7399,N_6169);
or U9226 (N_9226,N_5337,N_5311);
nor U9227 (N_9227,N_6669,N_7437);
or U9228 (N_9228,N_7463,N_5139);
or U9229 (N_9229,N_5344,N_5439);
and U9230 (N_9230,N_5427,N_5991);
and U9231 (N_9231,N_6849,N_5871);
and U9232 (N_9232,N_5556,N_7115);
nand U9233 (N_9233,N_6568,N_6015);
or U9234 (N_9234,N_5184,N_5561);
nor U9235 (N_9235,N_5682,N_5511);
or U9236 (N_9236,N_7496,N_6621);
nand U9237 (N_9237,N_5168,N_6468);
xnor U9238 (N_9238,N_6358,N_6801);
or U9239 (N_9239,N_7122,N_5614);
nand U9240 (N_9240,N_6211,N_5480);
or U9241 (N_9241,N_6979,N_5831);
xor U9242 (N_9242,N_5157,N_6635);
nor U9243 (N_9243,N_6913,N_7056);
and U9244 (N_9244,N_6745,N_7146);
or U9245 (N_9245,N_5736,N_5602);
nand U9246 (N_9246,N_5217,N_5476);
and U9247 (N_9247,N_6219,N_6040);
nor U9248 (N_9248,N_5014,N_7134);
or U9249 (N_9249,N_6255,N_7293);
nand U9250 (N_9250,N_6158,N_6396);
nand U9251 (N_9251,N_5247,N_6582);
nand U9252 (N_9252,N_6175,N_6732);
xor U9253 (N_9253,N_5775,N_5362);
nor U9254 (N_9254,N_5989,N_5441);
and U9255 (N_9255,N_6924,N_5435);
nor U9256 (N_9256,N_6466,N_5793);
nand U9257 (N_9257,N_6733,N_5554);
nor U9258 (N_9258,N_5988,N_6168);
or U9259 (N_9259,N_6689,N_6044);
and U9260 (N_9260,N_6360,N_6146);
nand U9261 (N_9261,N_5108,N_7037);
nor U9262 (N_9262,N_6816,N_5945);
nor U9263 (N_9263,N_6967,N_6922);
and U9264 (N_9264,N_7113,N_5840);
or U9265 (N_9265,N_5332,N_7146);
nor U9266 (N_9266,N_6623,N_6770);
and U9267 (N_9267,N_7230,N_6434);
or U9268 (N_9268,N_6588,N_5290);
nor U9269 (N_9269,N_5004,N_5424);
or U9270 (N_9270,N_5420,N_6604);
and U9271 (N_9271,N_6253,N_6927);
nand U9272 (N_9272,N_7451,N_5038);
and U9273 (N_9273,N_5582,N_5430);
nand U9274 (N_9274,N_6021,N_6720);
nor U9275 (N_9275,N_5496,N_5882);
nor U9276 (N_9276,N_6654,N_5696);
nor U9277 (N_9277,N_5054,N_5956);
and U9278 (N_9278,N_7065,N_6468);
nand U9279 (N_9279,N_5692,N_5024);
nor U9280 (N_9280,N_5643,N_6921);
nand U9281 (N_9281,N_6329,N_5352);
and U9282 (N_9282,N_6780,N_6358);
or U9283 (N_9283,N_6430,N_6253);
nor U9284 (N_9284,N_5104,N_6497);
nor U9285 (N_9285,N_6022,N_5157);
nor U9286 (N_9286,N_5421,N_5132);
nand U9287 (N_9287,N_6313,N_5690);
and U9288 (N_9288,N_6646,N_7474);
or U9289 (N_9289,N_6049,N_5513);
nand U9290 (N_9290,N_5628,N_5133);
or U9291 (N_9291,N_5420,N_6728);
or U9292 (N_9292,N_7304,N_5923);
nor U9293 (N_9293,N_5014,N_5013);
nor U9294 (N_9294,N_6132,N_7294);
nor U9295 (N_9295,N_6209,N_7364);
nand U9296 (N_9296,N_6781,N_5861);
nor U9297 (N_9297,N_5158,N_5747);
or U9298 (N_9298,N_5563,N_7072);
nor U9299 (N_9299,N_7319,N_5959);
or U9300 (N_9300,N_5999,N_5442);
and U9301 (N_9301,N_5514,N_6760);
and U9302 (N_9302,N_6253,N_7285);
nand U9303 (N_9303,N_5006,N_6128);
nor U9304 (N_9304,N_6429,N_5253);
xor U9305 (N_9305,N_5223,N_5221);
and U9306 (N_9306,N_5467,N_5514);
or U9307 (N_9307,N_7006,N_5934);
nor U9308 (N_9308,N_6352,N_5694);
nand U9309 (N_9309,N_7028,N_5455);
and U9310 (N_9310,N_6372,N_7310);
nor U9311 (N_9311,N_5320,N_5685);
nand U9312 (N_9312,N_5268,N_5966);
nor U9313 (N_9313,N_6130,N_6978);
nand U9314 (N_9314,N_5970,N_7071);
xnor U9315 (N_9315,N_7038,N_7478);
nand U9316 (N_9316,N_5745,N_5869);
nand U9317 (N_9317,N_6782,N_6849);
nor U9318 (N_9318,N_5821,N_6030);
nor U9319 (N_9319,N_7038,N_5013);
and U9320 (N_9320,N_6987,N_5863);
nand U9321 (N_9321,N_6008,N_7272);
or U9322 (N_9322,N_5651,N_7362);
nor U9323 (N_9323,N_6593,N_5647);
nand U9324 (N_9324,N_5897,N_7285);
nor U9325 (N_9325,N_6855,N_7302);
nor U9326 (N_9326,N_5895,N_7070);
and U9327 (N_9327,N_7029,N_5424);
nor U9328 (N_9328,N_6237,N_5602);
nor U9329 (N_9329,N_6379,N_6052);
and U9330 (N_9330,N_6907,N_5474);
and U9331 (N_9331,N_5051,N_5229);
xor U9332 (N_9332,N_5486,N_7390);
xor U9333 (N_9333,N_6807,N_7365);
nand U9334 (N_9334,N_5809,N_6892);
nand U9335 (N_9335,N_5721,N_5567);
nand U9336 (N_9336,N_7354,N_5408);
nand U9337 (N_9337,N_5765,N_6039);
or U9338 (N_9338,N_7136,N_6457);
xnor U9339 (N_9339,N_6102,N_7164);
nand U9340 (N_9340,N_6450,N_5810);
nor U9341 (N_9341,N_6103,N_6682);
or U9342 (N_9342,N_5514,N_6410);
nand U9343 (N_9343,N_6382,N_5538);
nor U9344 (N_9344,N_7059,N_5691);
or U9345 (N_9345,N_5967,N_5219);
nand U9346 (N_9346,N_6558,N_7235);
and U9347 (N_9347,N_6370,N_5338);
nor U9348 (N_9348,N_6397,N_5038);
nor U9349 (N_9349,N_5324,N_5452);
nand U9350 (N_9350,N_6541,N_6351);
nand U9351 (N_9351,N_6485,N_6158);
xnor U9352 (N_9352,N_5195,N_5792);
nand U9353 (N_9353,N_6458,N_7168);
nand U9354 (N_9354,N_6103,N_5962);
nand U9355 (N_9355,N_6786,N_5365);
or U9356 (N_9356,N_5540,N_5845);
nor U9357 (N_9357,N_5872,N_6707);
and U9358 (N_9358,N_5563,N_5068);
or U9359 (N_9359,N_6061,N_5020);
or U9360 (N_9360,N_5950,N_6830);
nand U9361 (N_9361,N_6602,N_5461);
nor U9362 (N_9362,N_5126,N_7382);
nand U9363 (N_9363,N_7074,N_5425);
or U9364 (N_9364,N_5147,N_6497);
nand U9365 (N_9365,N_5067,N_6551);
xnor U9366 (N_9366,N_5594,N_7212);
nand U9367 (N_9367,N_6462,N_6152);
or U9368 (N_9368,N_5150,N_5816);
nor U9369 (N_9369,N_5887,N_5540);
nor U9370 (N_9370,N_6295,N_7217);
and U9371 (N_9371,N_5926,N_5789);
or U9372 (N_9372,N_7482,N_5758);
nand U9373 (N_9373,N_6479,N_6022);
nand U9374 (N_9374,N_6927,N_6490);
nor U9375 (N_9375,N_6490,N_5962);
nand U9376 (N_9376,N_5865,N_7308);
nor U9377 (N_9377,N_6358,N_7203);
nor U9378 (N_9378,N_7450,N_5178);
and U9379 (N_9379,N_5213,N_7013);
and U9380 (N_9380,N_5402,N_7016);
nor U9381 (N_9381,N_5662,N_6439);
xnor U9382 (N_9382,N_5750,N_5062);
and U9383 (N_9383,N_5602,N_5335);
and U9384 (N_9384,N_6926,N_5765);
and U9385 (N_9385,N_6158,N_7335);
and U9386 (N_9386,N_6662,N_6584);
nor U9387 (N_9387,N_5535,N_6779);
nand U9388 (N_9388,N_5920,N_7486);
nand U9389 (N_9389,N_6831,N_5173);
nand U9390 (N_9390,N_6718,N_6282);
or U9391 (N_9391,N_5942,N_7193);
nand U9392 (N_9392,N_5230,N_5673);
xor U9393 (N_9393,N_5665,N_5017);
nor U9394 (N_9394,N_5052,N_6319);
nand U9395 (N_9395,N_5735,N_6775);
nor U9396 (N_9396,N_7132,N_5310);
nand U9397 (N_9397,N_6968,N_7128);
nor U9398 (N_9398,N_6470,N_5565);
and U9399 (N_9399,N_6039,N_6541);
or U9400 (N_9400,N_7240,N_6866);
xnor U9401 (N_9401,N_6146,N_5329);
xor U9402 (N_9402,N_5087,N_6976);
nand U9403 (N_9403,N_7045,N_5818);
and U9404 (N_9404,N_6772,N_5672);
or U9405 (N_9405,N_7223,N_5925);
nand U9406 (N_9406,N_7284,N_5087);
xor U9407 (N_9407,N_5254,N_6009);
and U9408 (N_9408,N_7276,N_7119);
xnor U9409 (N_9409,N_7298,N_6778);
or U9410 (N_9410,N_5749,N_6927);
nand U9411 (N_9411,N_7186,N_5929);
nor U9412 (N_9412,N_6465,N_6076);
and U9413 (N_9413,N_6843,N_5706);
and U9414 (N_9414,N_5024,N_6871);
or U9415 (N_9415,N_7182,N_7381);
nor U9416 (N_9416,N_7098,N_7258);
nand U9417 (N_9417,N_5157,N_5587);
nand U9418 (N_9418,N_6261,N_7478);
nor U9419 (N_9419,N_6773,N_5051);
and U9420 (N_9420,N_7243,N_5329);
and U9421 (N_9421,N_5453,N_5634);
nor U9422 (N_9422,N_5593,N_6780);
nand U9423 (N_9423,N_5393,N_5404);
xnor U9424 (N_9424,N_6532,N_7186);
or U9425 (N_9425,N_6472,N_5845);
nand U9426 (N_9426,N_7266,N_5171);
nand U9427 (N_9427,N_6019,N_7029);
nor U9428 (N_9428,N_5069,N_5530);
nor U9429 (N_9429,N_6306,N_5289);
nand U9430 (N_9430,N_5245,N_6901);
or U9431 (N_9431,N_5901,N_5312);
nor U9432 (N_9432,N_5995,N_5052);
nor U9433 (N_9433,N_7310,N_6513);
nand U9434 (N_9434,N_5851,N_5607);
and U9435 (N_9435,N_6838,N_7000);
and U9436 (N_9436,N_7292,N_5791);
nand U9437 (N_9437,N_5486,N_6051);
or U9438 (N_9438,N_5455,N_6793);
and U9439 (N_9439,N_6584,N_5518);
or U9440 (N_9440,N_7272,N_5800);
or U9441 (N_9441,N_7267,N_5129);
nor U9442 (N_9442,N_6528,N_6007);
xor U9443 (N_9443,N_6464,N_5508);
or U9444 (N_9444,N_5801,N_6779);
nand U9445 (N_9445,N_5285,N_6600);
or U9446 (N_9446,N_5782,N_5764);
nor U9447 (N_9447,N_5220,N_6471);
or U9448 (N_9448,N_5749,N_7036);
xor U9449 (N_9449,N_5041,N_7385);
or U9450 (N_9450,N_7496,N_5742);
nor U9451 (N_9451,N_6158,N_6418);
nor U9452 (N_9452,N_6593,N_6404);
and U9453 (N_9453,N_5911,N_5657);
nand U9454 (N_9454,N_6854,N_6053);
or U9455 (N_9455,N_6860,N_5181);
nand U9456 (N_9456,N_5590,N_6737);
or U9457 (N_9457,N_5413,N_5602);
and U9458 (N_9458,N_5930,N_6367);
nor U9459 (N_9459,N_6628,N_5484);
nor U9460 (N_9460,N_6496,N_5305);
nor U9461 (N_9461,N_7079,N_6893);
and U9462 (N_9462,N_7462,N_6001);
or U9463 (N_9463,N_5748,N_5713);
nand U9464 (N_9464,N_5497,N_5768);
or U9465 (N_9465,N_7052,N_6218);
nand U9466 (N_9466,N_6420,N_6325);
nor U9467 (N_9467,N_5945,N_5462);
nor U9468 (N_9468,N_6154,N_7331);
nor U9469 (N_9469,N_5168,N_6095);
and U9470 (N_9470,N_5303,N_5544);
and U9471 (N_9471,N_6881,N_5805);
nand U9472 (N_9472,N_5217,N_6007);
nor U9473 (N_9473,N_5006,N_6843);
nor U9474 (N_9474,N_7423,N_6048);
and U9475 (N_9475,N_6909,N_5507);
nand U9476 (N_9476,N_5336,N_5513);
nor U9477 (N_9477,N_6033,N_5814);
xnor U9478 (N_9478,N_6091,N_6427);
and U9479 (N_9479,N_6344,N_7054);
and U9480 (N_9480,N_5599,N_7227);
nor U9481 (N_9481,N_5409,N_6365);
nor U9482 (N_9482,N_7261,N_6793);
nand U9483 (N_9483,N_5966,N_5089);
nor U9484 (N_9484,N_6153,N_7042);
nand U9485 (N_9485,N_5182,N_5808);
nor U9486 (N_9486,N_7300,N_7020);
or U9487 (N_9487,N_5303,N_6287);
and U9488 (N_9488,N_7182,N_7110);
nand U9489 (N_9489,N_6518,N_6121);
and U9490 (N_9490,N_7249,N_5725);
or U9491 (N_9491,N_6015,N_6259);
nand U9492 (N_9492,N_7240,N_5820);
and U9493 (N_9493,N_5388,N_6024);
and U9494 (N_9494,N_5977,N_5384);
xor U9495 (N_9495,N_5539,N_6322);
or U9496 (N_9496,N_6124,N_7097);
and U9497 (N_9497,N_5920,N_6126);
and U9498 (N_9498,N_6544,N_6064);
nor U9499 (N_9499,N_6867,N_5895);
nor U9500 (N_9500,N_7024,N_7374);
xnor U9501 (N_9501,N_7331,N_5082);
nor U9502 (N_9502,N_5764,N_5583);
nand U9503 (N_9503,N_5411,N_6020);
and U9504 (N_9504,N_5346,N_5615);
or U9505 (N_9505,N_6329,N_5265);
or U9506 (N_9506,N_5883,N_7347);
or U9507 (N_9507,N_5232,N_5845);
and U9508 (N_9508,N_5402,N_5267);
and U9509 (N_9509,N_7132,N_5047);
nand U9510 (N_9510,N_7248,N_6363);
and U9511 (N_9511,N_5124,N_6797);
nand U9512 (N_9512,N_7056,N_5413);
and U9513 (N_9513,N_5294,N_7341);
nand U9514 (N_9514,N_5269,N_7458);
nor U9515 (N_9515,N_6966,N_6530);
and U9516 (N_9516,N_6849,N_5874);
and U9517 (N_9517,N_5467,N_5003);
nand U9518 (N_9518,N_5749,N_7157);
xnor U9519 (N_9519,N_5487,N_5741);
xor U9520 (N_9520,N_7043,N_7297);
nor U9521 (N_9521,N_7011,N_5484);
nand U9522 (N_9522,N_5629,N_7171);
or U9523 (N_9523,N_5059,N_6265);
nor U9524 (N_9524,N_7098,N_7122);
nand U9525 (N_9525,N_5050,N_5106);
and U9526 (N_9526,N_5098,N_5030);
nand U9527 (N_9527,N_6211,N_7498);
nand U9528 (N_9528,N_5830,N_5989);
or U9529 (N_9529,N_7123,N_5416);
nand U9530 (N_9530,N_6673,N_6063);
nor U9531 (N_9531,N_5553,N_6184);
or U9532 (N_9532,N_7459,N_6092);
or U9533 (N_9533,N_6864,N_6660);
nor U9534 (N_9534,N_5338,N_5948);
xor U9535 (N_9535,N_6526,N_5375);
or U9536 (N_9536,N_7289,N_5522);
or U9537 (N_9537,N_5265,N_7179);
nand U9538 (N_9538,N_5337,N_5966);
or U9539 (N_9539,N_6727,N_5495);
and U9540 (N_9540,N_5468,N_6146);
or U9541 (N_9541,N_6613,N_5824);
and U9542 (N_9542,N_5482,N_5240);
or U9543 (N_9543,N_7384,N_5286);
and U9544 (N_9544,N_5923,N_6185);
nor U9545 (N_9545,N_6292,N_5760);
xor U9546 (N_9546,N_7224,N_6234);
nand U9547 (N_9547,N_7056,N_6632);
and U9548 (N_9548,N_7365,N_5792);
nor U9549 (N_9549,N_6004,N_6290);
nor U9550 (N_9550,N_7244,N_5500);
and U9551 (N_9551,N_5304,N_5814);
nand U9552 (N_9552,N_6144,N_5869);
or U9553 (N_9553,N_5383,N_5586);
nor U9554 (N_9554,N_5809,N_7499);
and U9555 (N_9555,N_6466,N_7320);
or U9556 (N_9556,N_5802,N_6653);
nand U9557 (N_9557,N_5209,N_7381);
or U9558 (N_9558,N_6482,N_6171);
and U9559 (N_9559,N_5586,N_6806);
nand U9560 (N_9560,N_5169,N_6808);
nor U9561 (N_9561,N_6248,N_6614);
nand U9562 (N_9562,N_5935,N_6254);
or U9563 (N_9563,N_6578,N_5867);
xnor U9564 (N_9564,N_7041,N_5368);
or U9565 (N_9565,N_6601,N_5882);
nand U9566 (N_9566,N_6675,N_6877);
or U9567 (N_9567,N_5124,N_7403);
nor U9568 (N_9568,N_5752,N_5231);
nor U9569 (N_9569,N_5481,N_7335);
and U9570 (N_9570,N_7109,N_7093);
nor U9571 (N_9571,N_6078,N_6126);
nor U9572 (N_9572,N_5569,N_5080);
nor U9573 (N_9573,N_6415,N_7337);
xnor U9574 (N_9574,N_6769,N_5331);
and U9575 (N_9575,N_7187,N_6912);
nand U9576 (N_9576,N_5880,N_7435);
and U9577 (N_9577,N_5221,N_5647);
nand U9578 (N_9578,N_7347,N_6310);
or U9579 (N_9579,N_6428,N_7120);
nand U9580 (N_9580,N_6409,N_5195);
nand U9581 (N_9581,N_5880,N_7421);
xnor U9582 (N_9582,N_5875,N_7395);
nor U9583 (N_9583,N_7357,N_5109);
or U9584 (N_9584,N_6021,N_5755);
nand U9585 (N_9585,N_6079,N_6148);
nor U9586 (N_9586,N_6082,N_5312);
nor U9587 (N_9587,N_5481,N_6612);
and U9588 (N_9588,N_5498,N_5802);
nor U9589 (N_9589,N_5439,N_7257);
nor U9590 (N_9590,N_5104,N_5182);
nor U9591 (N_9591,N_6218,N_5875);
or U9592 (N_9592,N_5919,N_6023);
nand U9593 (N_9593,N_5196,N_7464);
nor U9594 (N_9594,N_5755,N_6086);
xor U9595 (N_9595,N_6910,N_6502);
or U9596 (N_9596,N_6190,N_5176);
nand U9597 (N_9597,N_6982,N_5169);
xnor U9598 (N_9598,N_5271,N_5245);
and U9599 (N_9599,N_6659,N_6364);
xor U9600 (N_9600,N_7203,N_7322);
or U9601 (N_9601,N_6335,N_6481);
nand U9602 (N_9602,N_5785,N_6475);
nor U9603 (N_9603,N_6804,N_7123);
nand U9604 (N_9604,N_6440,N_5917);
and U9605 (N_9605,N_6187,N_7056);
and U9606 (N_9606,N_6710,N_7030);
and U9607 (N_9607,N_6567,N_6298);
nor U9608 (N_9608,N_5661,N_5233);
nor U9609 (N_9609,N_5283,N_6451);
and U9610 (N_9610,N_6094,N_6110);
and U9611 (N_9611,N_5932,N_5364);
nor U9612 (N_9612,N_7137,N_6824);
or U9613 (N_9613,N_6414,N_5899);
nand U9614 (N_9614,N_6382,N_5742);
nor U9615 (N_9615,N_7007,N_6934);
nand U9616 (N_9616,N_5645,N_5655);
and U9617 (N_9617,N_5106,N_6900);
nand U9618 (N_9618,N_5264,N_6012);
and U9619 (N_9619,N_5822,N_7398);
nand U9620 (N_9620,N_5567,N_6966);
xor U9621 (N_9621,N_5923,N_6853);
nor U9622 (N_9622,N_7361,N_7305);
nand U9623 (N_9623,N_5123,N_5073);
nor U9624 (N_9624,N_5977,N_5255);
nor U9625 (N_9625,N_6817,N_6643);
and U9626 (N_9626,N_5115,N_6156);
nor U9627 (N_9627,N_6988,N_7127);
nor U9628 (N_9628,N_7286,N_5138);
nand U9629 (N_9629,N_5949,N_5281);
nand U9630 (N_9630,N_5754,N_6832);
or U9631 (N_9631,N_6992,N_6087);
nor U9632 (N_9632,N_6862,N_6354);
nand U9633 (N_9633,N_5026,N_5732);
or U9634 (N_9634,N_6488,N_6190);
nand U9635 (N_9635,N_6711,N_5941);
nand U9636 (N_9636,N_7428,N_6357);
nor U9637 (N_9637,N_6797,N_7280);
nand U9638 (N_9638,N_5127,N_6308);
or U9639 (N_9639,N_6065,N_7030);
xor U9640 (N_9640,N_6949,N_5558);
or U9641 (N_9641,N_6708,N_6576);
nand U9642 (N_9642,N_6350,N_5085);
and U9643 (N_9643,N_5044,N_7129);
and U9644 (N_9644,N_6240,N_5317);
or U9645 (N_9645,N_6558,N_5843);
nand U9646 (N_9646,N_6132,N_5359);
xor U9647 (N_9647,N_7042,N_5123);
nand U9648 (N_9648,N_5568,N_6472);
nand U9649 (N_9649,N_6677,N_7474);
and U9650 (N_9650,N_5268,N_6969);
nand U9651 (N_9651,N_6467,N_7345);
nor U9652 (N_9652,N_5398,N_6452);
nor U9653 (N_9653,N_5873,N_5826);
or U9654 (N_9654,N_6684,N_6192);
or U9655 (N_9655,N_7452,N_5387);
nand U9656 (N_9656,N_5939,N_6794);
nor U9657 (N_9657,N_5773,N_7430);
or U9658 (N_9658,N_6468,N_7210);
or U9659 (N_9659,N_5970,N_5684);
nand U9660 (N_9660,N_6443,N_6594);
nand U9661 (N_9661,N_7488,N_7206);
or U9662 (N_9662,N_6922,N_5067);
or U9663 (N_9663,N_5632,N_5595);
or U9664 (N_9664,N_7299,N_7361);
nand U9665 (N_9665,N_6548,N_5498);
nand U9666 (N_9666,N_7366,N_5122);
or U9667 (N_9667,N_5328,N_6721);
nor U9668 (N_9668,N_7323,N_6105);
or U9669 (N_9669,N_5304,N_5006);
or U9670 (N_9670,N_5221,N_6823);
nor U9671 (N_9671,N_7229,N_5738);
nor U9672 (N_9672,N_6494,N_5300);
xor U9673 (N_9673,N_6268,N_5003);
nor U9674 (N_9674,N_5996,N_5479);
or U9675 (N_9675,N_5009,N_5426);
and U9676 (N_9676,N_5381,N_5363);
or U9677 (N_9677,N_5252,N_6257);
nor U9678 (N_9678,N_6122,N_5080);
xor U9679 (N_9679,N_5090,N_5408);
xor U9680 (N_9680,N_5894,N_6527);
nand U9681 (N_9681,N_5401,N_6532);
or U9682 (N_9682,N_6216,N_5582);
nand U9683 (N_9683,N_6797,N_6227);
nand U9684 (N_9684,N_6184,N_5768);
xnor U9685 (N_9685,N_5692,N_6708);
and U9686 (N_9686,N_6908,N_6888);
nor U9687 (N_9687,N_5338,N_6047);
or U9688 (N_9688,N_7157,N_5143);
and U9689 (N_9689,N_5105,N_6214);
nand U9690 (N_9690,N_6537,N_5621);
and U9691 (N_9691,N_5030,N_5581);
or U9692 (N_9692,N_6647,N_7474);
and U9693 (N_9693,N_6241,N_7073);
nor U9694 (N_9694,N_6936,N_6517);
nor U9695 (N_9695,N_6526,N_6614);
and U9696 (N_9696,N_6346,N_7239);
or U9697 (N_9697,N_7470,N_5008);
nor U9698 (N_9698,N_5730,N_5477);
or U9699 (N_9699,N_5075,N_5482);
or U9700 (N_9700,N_7220,N_5698);
and U9701 (N_9701,N_7014,N_5269);
or U9702 (N_9702,N_6852,N_6397);
nand U9703 (N_9703,N_7127,N_5369);
or U9704 (N_9704,N_5445,N_5804);
nand U9705 (N_9705,N_5089,N_7374);
and U9706 (N_9706,N_5468,N_5018);
nor U9707 (N_9707,N_6925,N_6001);
or U9708 (N_9708,N_7020,N_5221);
xor U9709 (N_9709,N_6008,N_6394);
nand U9710 (N_9710,N_7314,N_6171);
nor U9711 (N_9711,N_5794,N_5290);
nand U9712 (N_9712,N_6399,N_6406);
nor U9713 (N_9713,N_5118,N_7079);
nor U9714 (N_9714,N_7295,N_7199);
or U9715 (N_9715,N_6636,N_7364);
nand U9716 (N_9716,N_5631,N_5362);
nor U9717 (N_9717,N_5040,N_6564);
and U9718 (N_9718,N_6033,N_6534);
nand U9719 (N_9719,N_7067,N_5261);
xor U9720 (N_9720,N_7397,N_6421);
nor U9721 (N_9721,N_6946,N_6491);
xnor U9722 (N_9722,N_6492,N_7221);
nand U9723 (N_9723,N_6219,N_6241);
nor U9724 (N_9724,N_5047,N_5004);
nor U9725 (N_9725,N_6382,N_5935);
xnor U9726 (N_9726,N_7479,N_7160);
nor U9727 (N_9727,N_6676,N_6829);
or U9728 (N_9728,N_5576,N_6068);
or U9729 (N_9729,N_5344,N_6069);
or U9730 (N_9730,N_6338,N_5131);
nor U9731 (N_9731,N_5207,N_6414);
nor U9732 (N_9732,N_6954,N_5069);
xnor U9733 (N_9733,N_6006,N_5002);
nor U9734 (N_9734,N_5632,N_5204);
nor U9735 (N_9735,N_6594,N_6431);
xor U9736 (N_9736,N_5851,N_7189);
and U9737 (N_9737,N_7002,N_6421);
and U9738 (N_9738,N_6626,N_5373);
or U9739 (N_9739,N_5697,N_6870);
or U9740 (N_9740,N_5817,N_6225);
or U9741 (N_9741,N_6841,N_6106);
or U9742 (N_9742,N_7406,N_5007);
xnor U9743 (N_9743,N_6963,N_7022);
nor U9744 (N_9744,N_7450,N_7271);
nor U9745 (N_9745,N_5069,N_6038);
or U9746 (N_9746,N_5192,N_5249);
nand U9747 (N_9747,N_7159,N_6086);
or U9748 (N_9748,N_6676,N_6011);
or U9749 (N_9749,N_6258,N_7034);
and U9750 (N_9750,N_7178,N_5377);
and U9751 (N_9751,N_6021,N_5138);
and U9752 (N_9752,N_5344,N_6698);
nor U9753 (N_9753,N_7066,N_7249);
or U9754 (N_9754,N_6649,N_6759);
xnor U9755 (N_9755,N_7064,N_6792);
nand U9756 (N_9756,N_5530,N_5395);
nor U9757 (N_9757,N_7243,N_5899);
nor U9758 (N_9758,N_6363,N_7167);
or U9759 (N_9759,N_6359,N_5590);
nor U9760 (N_9760,N_6055,N_6297);
or U9761 (N_9761,N_5889,N_5265);
nor U9762 (N_9762,N_7002,N_7005);
or U9763 (N_9763,N_6431,N_6297);
nor U9764 (N_9764,N_5209,N_5316);
xnor U9765 (N_9765,N_6541,N_5227);
and U9766 (N_9766,N_5995,N_6243);
or U9767 (N_9767,N_5538,N_5957);
nand U9768 (N_9768,N_6407,N_6690);
nor U9769 (N_9769,N_7086,N_6557);
nand U9770 (N_9770,N_6287,N_7285);
nand U9771 (N_9771,N_5267,N_7296);
or U9772 (N_9772,N_7115,N_6046);
or U9773 (N_9773,N_7268,N_5243);
or U9774 (N_9774,N_5771,N_7039);
and U9775 (N_9775,N_5359,N_6857);
and U9776 (N_9776,N_5189,N_5761);
and U9777 (N_9777,N_6342,N_5403);
or U9778 (N_9778,N_6057,N_5493);
or U9779 (N_9779,N_6771,N_6605);
nand U9780 (N_9780,N_6623,N_6479);
or U9781 (N_9781,N_5889,N_5769);
and U9782 (N_9782,N_6407,N_6879);
nor U9783 (N_9783,N_5860,N_5446);
or U9784 (N_9784,N_5762,N_7395);
nor U9785 (N_9785,N_5039,N_6499);
xnor U9786 (N_9786,N_6787,N_5826);
or U9787 (N_9787,N_6665,N_5838);
and U9788 (N_9788,N_7275,N_6210);
nand U9789 (N_9789,N_6373,N_5424);
nand U9790 (N_9790,N_6203,N_6423);
nand U9791 (N_9791,N_6734,N_6390);
xor U9792 (N_9792,N_6024,N_6473);
and U9793 (N_9793,N_6491,N_6394);
and U9794 (N_9794,N_5252,N_5340);
and U9795 (N_9795,N_6271,N_5679);
nand U9796 (N_9796,N_5300,N_5377);
nand U9797 (N_9797,N_5472,N_6559);
nor U9798 (N_9798,N_6181,N_5024);
nand U9799 (N_9799,N_5104,N_5486);
nor U9800 (N_9800,N_5087,N_5985);
and U9801 (N_9801,N_7357,N_7259);
xnor U9802 (N_9802,N_6851,N_7270);
nand U9803 (N_9803,N_5015,N_6524);
nand U9804 (N_9804,N_6977,N_6295);
xor U9805 (N_9805,N_7048,N_6425);
or U9806 (N_9806,N_6545,N_5310);
nor U9807 (N_9807,N_5960,N_7047);
nor U9808 (N_9808,N_5130,N_5677);
and U9809 (N_9809,N_7352,N_6241);
or U9810 (N_9810,N_6852,N_5215);
and U9811 (N_9811,N_6766,N_7347);
xnor U9812 (N_9812,N_6308,N_6226);
or U9813 (N_9813,N_7261,N_7011);
nand U9814 (N_9814,N_5971,N_5669);
and U9815 (N_9815,N_5890,N_6922);
or U9816 (N_9816,N_6992,N_5686);
nand U9817 (N_9817,N_7269,N_5211);
and U9818 (N_9818,N_5872,N_7119);
or U9819 (N_9819,N_6127,N_5942);
and U9820 (N_9820,N_7085,N_6377);
or U9821 (N_9821,N_7172,N_5540);
nand U9822 (N_9822,N_5907,N_6765);
or U9823 (N_9823,N_5378,N_5108);
or U9824 (N_9824,N_6780,N_5778);
nand U9825 (N_9825,N_5266,N_5420);
nor U9826 (N_9826,N_5628,N_5428);
nor U9827 (N_9827,N_6465,N_5152);
nand U9828 (N_9828,N_6042,N_5942);
and U9829 (N_9829,N_5892,N_5276);
nand U9830 (N_9830,N_5358,N_7328);
or U9831 (N_9831,N_6631,N_6871);
and U9832 (N_9832,N_5846,N_7082);
nor U9833 (N_9833,N_6088,N_6963);
nor U9834 (N_9834,N_5548,N_5240);
nand U9835 (N_9835,N_6878,N_7272);
nor U9836 (N_9836,N_5796,N_5522);
or U9837 (N_9837,N_7239,N_5030);
and U9838 (N_9838,N_5191,N_5104);
or U9839 (N_9839,N_6043,N_5970);
nor U9840 (N_9840,N_7414,N_6910);
or U9841 (N_9841,N_6390,N_6725);
nor U9842 (N_9842,N_6313,N_5932);
or U9843 (N_9843,N_7156,N_7295);
nor U9844 (N_9844,N_7005,N_6726);
or U9845 (N_9845,N_5217,N_5091);
xor U9846 (N_9846,N_5558,N_6693);
nor U9847 (N_9847,N_7481,N_7200);
or U9848 (N_9848,N_5193,N_5609);
and U9849 (N_9849,N_6022,N_6013);
nand U9850 (N_9850,N_6742,N_6599);
and U9851 (N_9851,N_7372,N_6095);
or U9852 (N_9852,N_6809,N_6967);
and U9853 (N_9853,N_5144,N_5781);
xor U9854 (N_9854,N_5169,N_6523);
or U9855 (N_9855,N_5277,N_5322);
nor U9856 (N_9856,N_7041,N_5804);
or U9857 (N_9857,N_7296,N_6831);
nor U9858 (N_9858,N_5634,N_7178);
xnor U9859 (N_9859,N_6381,N_5195);
xnor U9860 (N_9860,N_6470,N_6857);
nand U9861 (N_9861,N_6999,N_6606);
nor U9862 (N_9862,N_6125,N_6956);
or U9863 (N_9863,N_6780,N_5134);
nand U9864 (N_9864,N_6634,N_6374);
nor U9865 (N_9865,N_6462,N_5238);
or U9866 (N_9866,N_7088,N_6513);
nand U9867 (N_9867,N_6001,N_6905);
nor U9868 (N_9868,N_5286,N_5298);
and U9869 (N_9869,N_5753,N_5372);
or U9870 (N_9870,N_6011,N_5238);
nor U9871 (N_9871,N_7335,N_6672);
nand U9872 (N_9872,N_7009,N_6859);
nand U9873 (N_9873,N_6239,N_5454);
xor U9874 (N_9874,N_6085,N_6443);
nor U9875 (N_9875,N_5248,N_5191);
or U9876 (N_9876,N_6297,N_6565);
or U9877 (N_9877,N_7285,N_7474);
or U9878 (N_9878,N_6779,N_5127);
or U9879 (N_9879,N_6265,N_5297);
or U9880 (N_9880,N_5719,N_6295);
nand U9881 (N_9881,N_6098,N_6613);
or U9882 (N_9882,N_7459,N_7305);
and U9883 (N_9883,N_6472,N_6811);
or U9884 (N_9884,N_5850,N_7171);
nor U9885 (N_9885,N_6482,N_6676);
nand U9886 (N_9886,N_5028,N_7299);
xnor U9887 (N_9887,N_5950,N_6182);
xnor U9888 (N_9888,N_5255,N_5206);
xnor U9889 (N_9889,N_5683,N_5298);
or U9890 (N_9890,N_7360,N_5933);
and U9891 (N_9891,N_5072,N_6613);
and U9892 (N_9892,N_6168,N_6961);
or U9893 (N_9893,N_6713,N_6759);
or U9894 (N_9894,N_6260,N_6974);
nor U9895 (N_9895,N_6044,N_7430);
nor U9896 (N_9896,N_5822,N_7441);
nor U9897 (N_9897,N_6468,N_5369);
nand U9898 (N_9898,N_6238,N_5458);
nand U9899 (N_9899,N_6091,N_7170);
xnor U9900 (N_9900,N_6728,N_5698);
nor U9901 (N_9901,N_5407,N_6668);
and U9902 (N_9902,N_7233,N_6348);
nand U9903 (N_9903,N_7022,N_5471);
and U9904 (N_9904,N_6400,N_5279);
nor U9905 (N_9905,N_6122,N_5005);
nor U9906 (N_9906,N_5702,N_6064);
nor U9907 (N_9907,N_6868,N_7346);
nor U9908 (N_9908,N_6526,N_6840);
xor U9909 (N_9909,N_6100,N_6033);
nand U9910 (N_9910,N_6602,N_7204);
and U9911 (N_9911,N_5958,N_6720);
nand U9912 (N_9912,N_6803,N_5579);
xor U9913 (N_9913,N_6955,N_7460);
xnor U9914 (N_9914,N_5332,N_7259);
nor U9915 (N_9915,N_5738,N_5057);
or U9916 (N_9916,N_6198,N_5805);
nor U9917 (N_9917,N_6319,N_7325);
nor U9918 (N_9918,N_6844,N_6192);
and U9919 (N_9919,N_6650,N_6601);
or U9920 (N_9920,N_5615,N_6835);
nor U9921 (N_9921,N_7172,N_6119);
and U9922 (N_9922,N_5560,N_7433);
and U9923 (N_9923,N_5314,N_5816);
nand U9924 (N_9924,N_7272,N_5377);
nand U9925 (N_9925,N_6095,N_5519);
or U9926 (N_9926,N_7411,N_6103);
nand U9927 (N_9927,N_6858,N_5538);
and U9928 (N_9928,N_6308,N_5386);
nor U9929 (N_9929,N_7274,N_6911);
nor U9930 (N_9930,N_5579,N_5002);
and U9931 (N_9931,N_6337,N_5050);
or U9932 (N_9932,N_6709,N_5073);
nand U9933 (N_9933,N_7497,N_5967);
nor U9934 (N_9934,N_7128,N_6185);
or U9935 (N_9935,N_5243,N_7347);
nor U9936 (N_9936,N_6481,N_5705);
or U9937 (N_9937,N_7108,N_7057);
or U9938 (N_9938,N_5110,N_7207);
and U9939 (N_9939,N_5111,N_6907);
nand U9940 (N_9940,N_6362,N_6648);
and U9941 (N_9941,N_6051,N_7172);
and U9942 (N_9942,N_6100,N_5097);
xnor U9943 (N_9943,N_6971,N_6589);
nand U9944 (N_9944,N_6678,N_5809);
nand U9945 (N_9945,N_6178,N_5843);
nor U9946 (N_9946,N_7003,N_5168);
xnor U9947 (N_9947,N_6708,N_7249);
and U9948 (N_9948,N_5802,N_5927);
or U9949 (N_9949,N_6441,N_5851);
xnor U9950 (N_9950,N_5236,N_5787);
nor U9951 (N_9951,N_6174,N_6573);
nand U9952 (N_9952,N_6744,N_5076);
nand U9953 (N_9953,N_6461,N_5381);
nand U9954 (N_9954,N_5035,N_5393);
nand U9955 (N_9955,N_5608,N_6414);
and U9956 (N_9956,N_5389,N_5998);
xor U9957 (N_9957,N_6457,N_6647);
and U9958 (N_9958,N_7199,N_6780);
nand U9959 (N_9959,N_5042,N_7250);
or U9960 (N_9960,N_5885,N_7319);
nand U9961 (N_9961,N_6936,N_6336);
and U9962 (N_9962,N_6959,N_7498);
or U9963 (N_9963,N_6423,N_5542);
or U9964 (N_9964,N_6215,N_6595);
xor U9965 (N_9965,N_5194,N_6840);
xnor U9966 (N_9966,N_6293,N_5020);
nand U9967 (N_9967,N_7365,N_6478);
nand U9968 (N_9968,N_6467,N_6510);
xor U9969 (N_9969,N_6198,N_6082);
nor U9970 (N_9970,N_6369,N_6662);
and U9971 (N_9971,N_6498,N_7221);
or U9972 (N_9972,N_5459,N_5994);
nor U9973 (N_9973,N_5826,N_5378);
nor U9974 (N_9974,N_5938,N_6966);
nand U9975 (N_9975,N_5380,N_5067);
nand U9976 (N_9976,N_5235,N_7128);
and U9977 (N_9977,N_7027,N_6415);
and U9978 (N_9978,N_6489,N_6959);
nand U9979 (N_9979,N_7356,N_5880);
nor U9980 (N_9980,N_6024,N_5667);
and U9981 (N_9981,N_5366,N_7493);
or U9982 (N_9982,N_6852,N_6382);
or U9983 (N_9983,N_6896,N_7059);
and U9984 (N_9984,N_6643,N_7219);
nand U9985 (N_9985,N_7252,N_5890);
and U9986 (N_9986,N_5761,N_6612);
xnor U9987 (N_9987,N_6611,N_7363);
or U9988 (N_9988,N_6390,N_5654);
or U9989 (N_9989,N_5777,N_5098);
nand U9990 (N_9990,N_5835,N_5280);
nand U9991 (N_9991,N_6103,N_7270);
and U9992 (N_9992,N_5749,N_7207);
or U9993 (N_9993,N_6219,N_5552);
nor U9994 (N_9994,N_6501,N_7194);
nand U9995 (N_9995,N_6048,N_6142);
nand U9996 (N_9996,N_7238,N_5927);
and U9997 (N_9997,N_5823,N_5699);
and U9998 (N_9998,N_5815,N_5550);
xnor U9999 (N_9999,N_6715,N_7261);
or UO_0 (O_0,N_8702,N_8445);
nor UO_1 (O_1,N_8262,N_8648);
or UO_2 (O_2,N_9033,N_9237);
xnor UO_3 (O_3,N_9175,N_8683);
nor UO_4 (O_4,N_8208,N_8097);
and UO_5 (O_5,N_9099,N_9433);
nand UO_6 (O_6,N_7717,N_7760);
nor UO_7 (O_7,N_9494,N_8092);
or UO_8 (O_8,N_8940,N_8539);
nand UO_9 (O_9,N_7854,N_7707);
nor UO_10 (O_10,N_7708,N_8623);
nor UO_11 (O_11,N_9809,N_7981);
xor UO_12 (O_12,N_7975,N_9343);
nand UO_13 (O_13,N_9934,N_7518);
and UO_14 (O_14,N_7862,N_7933);
nand UO_15 (O_15,N_9739,N_8575);
and UO_16 (O_16,N_7609,N_9651);
nor UO_17 (O_17,N_8266,N_9171);
nor UO_18 (O_18,N_9473,N_7555);
nor UO_19 (O_19,N_8602,N_7857);
or UO_20 (O_20,N_8244,N_8870);
and UO_21 (O_21,N_7739,N_9224);
nand UO_22 (O_22,N_8863,N_8204);
and UO_23 (O_23,N_9789,N_8419);
and UO_24 (O_24,N_9654,N_7901);
nand UO_25 (O_25,N_8641,N_9527);
and UO_26 (O_26,N_8311,N_9490);
nand UO_27 (O_27,N_8316,N_8912);
xor UO_28 (O_28,N_9474,N_8778);
and UO_29 (O_29,N_8213,N_9991);
or UO_30 (O_30,N_8987,N_9188);
or UO_31 (O_31,N_9357,N_9440);
and UO_32 (O_32,N_7568,N_9984);
nand UO_33 (O_33,N_8808,N_8815);
nor UO_34 (O_34,N_8110,N_9954);
and UO_35 (O_35,N_9782,N_9959);
and UO_36 (O_36,N_9716,N_8788);
or UO_37 (O_37,N_8588,N_9987);
nor UO_38 (O_38,N_9656,N_8856);
and UO_39 (O_39,N_9747,N_7956);
nand UO_40 (O_40,N_9381,N_9865);
nor UO_41 (O_41,N_8177,N_7722);
nand UO_42 (O_42,N_9724,N_8955);
nand UO_43 (O_43,N_9314,N_8621);
nor UO_44 (O_44,N_9287,N_9606);
nand UO_45 (O_45,N_7972,N_8592);
nand UO_46 (O_46,N_9818,N_9136);
or UO_47 (O_47,N_7848,N_8625);
nand UO_48 (O_48,N_9070,N_7619);
nor UO_49 (O_49,N_9297,N_8735);
and UO_50 (O_50,N_9678,N_9332);
or UO_51 (O_51,N_7825,N_7606);
and UO_52 (O_52,N_8030,N_7940);
and UO_53 (O_53,N_9373,N_8489);
and UO_54 (O_54,N_7799,N_9115);
nand UO_55 (O_55,N_7873,N_8949);
nor UO_56 (O_56,N_8239,N_7993);
nand UO_57 (O_57,N_8139,N_7761);
or UO_58 (O_58,N_8281,N_9014);
or UO_59 (O_59,N_9770,N_9869);
nand UO_60 (O_60,N_9650,N_8170);
or UO_61 (O_61,N_7770,N_8394);
nand UO_62 (O_62,N_9484,N_9498);
nor UO_63 (O_63,N_8728,N_7645);
or UO_64 (O_64,N_8104,N_7696);
xnor UO_65 (O_65,N_7856,N_8328);
nand UO_66 (O_66,N_8103,N_9477);
xnor UO_67 (O_67,N_7627,N_8527);
or UO_68 (O_68,N_7811,N_9466);
nand UO_69 (O_69,N_7970,N_7698);
or UO_70 (O_70,N_9333,N_7727);
or UO_71 (O_71,N_8136,N_9290);
or UO_72 (O_72,N_7711,N_7959);
nor UO_73 (O_73,N_7505,N_9783);
nand UO_74 (O_74,N_8721,N_8712);
nor UO_75 (O_75,N_9249,N_8167);
and UO_76 (O_76,N_8355,N_9049);
or UO_77 (O_77,N_8832,N_8306);
nand UO_78 (O_78,N_9980,N_9199);
and UO_79 (O_79,N_8288,N_8834);
nand UO_80 (O_80,N_9826,N_8564);
nor UO_81 (O_81,N_7923,N_9812);
xor UO_82 (O_82,N_7520,N_7971);
nand UO_83 (O_83,N_8759,N_7570);
nand UO_84 (O_84,N_8901,N_8669);
nor UO_85 (O_85,N_8523,N_9503);
and UO_86 (O_86,N_8447,N_9036);
nand UO_87 (O_87,N_7566,N_8862);
nand UO_88 (O_88,N_8697,N_8854);
nand UO_89 (O_89,N_8145,N_9540);
or UO_90 (O_90,N_8607,N_9534);
xnor UO_91 (O_91,N_8764,N_8522);
and UO_92 (O_92,N_8687,N_8091);
nand UO_93 (O_93,N_7903,N_9203);
or UO_94 (O_94,N_9345,N_8981);
nor UO_95 (O_95,N_8922,N_9380);
or UO_96 (O_96,N_9997,N_8658);
nor UO_97 (O_97,N_9080,N_8884);
nand UO_98 (O_98,N_8510,N_9879);
and UO_99 (O_99,N_9130,N_9748);
or UO_100 (O_100,N_9031,N_9384);
nand UO_101 (O_101,N_9492,N_9754);
nor UO_102 (O_102,N_8500,N_7652);
xor UO_103 (O_103,N_9504,N_9050);
nand UO_104 (O_104,N_7503,N_8017);
or UO_105 (O_105,N_9006,N_8406);
nand UO_106 (O_106,N_9127,N_9730);
and UO_107 (O_107,N_8939,N_8127);
nor UO_108 (O_108,N_7614,N_9548);
nor UO_109 (O_109,N_9363,N_8879);
nand UO_110 (O_110,N_8422,N_9082);
nor UO_111 (O_111,N_9276,N_8554);
nor UO_112 (O_112,N_8849,N_9221);
nor UO_113 (O_113,N_8726,N_9429);
and UO_114 (O_114,N_7967,N_9841);
nand UO_115 (O_115,N_8556,N_9568);
nor UO_116 (O_116,N_8787,N_9698);
nand UO_117 (O_117,N_8671,N_7908);
xor UO_118 (O_118,N_9536,N_8518);
nand UO_119 (O_119,N_8694,N_8289);
or UO_120 (O_120,N_8062,N_8709);
and UO_121 (O_121,N_7507,N_9254);
xor UO_122 (O_122,N_8317,N_8951);
and UO_123 (O_123,N_9419,N_8781);
and UO_124 (O_124,N_9881,N_8644);
and UO_125 (O_125,N_7751,N_9761);
or UO_126 (O_126,N_7607,N_8148);
nor UO_127 (O_127,N_9884,N_9220);
nand UO_128 (O_128,N_8878,N_7852);
nand UO_129 (O_129,N_8670,N_9391);
nor UO_130 (O_130,N_9686,N_8072);
and UO_131 (O_131,N_9637,N_9864);
and UO_132 (O_132,N_7596,N_8366);
nor UO_133 (O_133,N_9444,N_8075);
nor UO_134 (O_134,N_9787,N_7641);
or UO_135 (O_135,N_9110,N_8255);
or UO_136 (O_136,N_9704,N_8034);
and UO_137 (O_137,N_8055,N_9766);
or UO_138 (O_138,N_7579,N_9862);
or UO_139 (O_139,N_9305,N_7618);
or UO_140 (O_140,N_9705,N_8358);
nor UO_141 (O_141,N_7747,N_9772);
and UO_142 (O_142,N_8600,N_8268);
or UO_143 (O_143,N_9346,N_9848);
or UO_144 (O_144,N_7748,N_8341);
nand UO_145 (O_145,N_8713,N_8277);
nor UO_146 (O_146,N_7658,N_9159);
and UO_147 (O_147,N_9587,N_8198);
or UO_148 (O_148,N_9134,N_8546);
nand UO_149 (O_149,N_9608,N_7752);
nor UO_150 (O_150,N_9905,N_7807);
or UO_151 (O_151,N_8356,N_9633);
nand UO_152 (O_152,N_8555,N_9908);
nand UO_153 (O_153,N_8482,N_9668);
or UO_154 (O_154,N_8704,N_7872);
or UO_155 (O_155,N_8013,N_9952);
or UO_156 (O_156,N_7945,N_8583);
or UO_157 (O_157,N_7947,N_9740);
xor UO_158 (O_158,N_8639,N_9547);
and UO_159 (O_159,N_9328,N_7954);
and UO_160 (O_160,N_8819,N_8467);
nor UO_161 (O_161,N_9154,N_9522);
or UO_162 (O_162,N_7858,N_9893);
nand UO_163 (O_163,N_9349,N_9227);
and UO_164 (O_164,N_8488,N_7720);
and UO_165 (O_165,N_7528,N_9008);
or UO_166 (O_166,N_7815,N_8001);
xor UO_167 (O_167,N_8312,N_8654);
nand UO_168 (O_168,N_7828,N_9009);
nand UO_169 (O_169,N_8258,N_9330);
nor UO_170 (O_170,N_9193,N_9933);
nor UO_171 (O_171,N_9844,N_9128);
xor UO_172 (O_172,N_9538,N_7690);
or UO_173 (O_173,N_9040,N_8932);
nor UO_174 (O_174,N_8885,N_9774);
nand UO_175 (O_175,N_9410,N_9415);
nor UO_176 (O_176,N_9635,N_8586);
or UO_177 (O_177,N_8401,N_7500);
nand UO_178 (O_178,N_8615,N_9423);
and UO_179 (O_179,N_7949,N_9574);
nor UO_180 (O_180,N_8182,N_9518);
nor UO_181 (O_181,N_8507,N_8746);
nand UO_182 (O_182,N_9260,N_9197);
xor UO_183 (O_183,N_8763,N_9471);
nor UO_184 (O_184,N_7691,N_9375);
and UO_185 (O_185,N_8750,N_9849);
and UO_186 (O_186,N_9830,N_9513);
and UO_187 (O_187,N_9383,N_8631);
and UO_188 (O_188,N_8047,N_9463);
and UO_189 (O_189,N_9960,N_9268);
nor UO_190 (O_190,N_8984,N_8881);
and UO_191 (O_191,N_9813,N_7796);
or UO_192 (O_192,N_7938,N_8428);
and UO_193 (O_193,N_9597,N_9112);
nand UO_194 (O_194,N_8042,N_9507);
nand UO_195 (O_195,N_8462,N_8083);
and UO_196 (O_196,N_9392,N_9092);
nor UO_197 (O_197,N_7794,N_8534);
nand UO_198 (O_198,N_9921,N_7578);
nand UO_199 (O_199,N_8407,N_8649);
nand UO_200 (O_200,N_9222,N_8526);
nand UO_201 (O_201,N_8577,N_8221);
nor UO_202 (O_202,N_8905,N_7869);
nand UO_203 (O_203,N_8098,N_8494);
nor UO_204 (O_204,N_9455,N_8132);
nand UO_205 (O_205,N_7800,N_8188);
or UO_206 (O_206,N_8099,N_9184);
nand UO_207 (O_207,N_9946,N_9255);
nand UO_208 (O_208,N_8918,N_8847);
nand UO_209 (O_209,N_9262,N_8578);
nor UO_210 (O_210,N_8044,N_7847);
nor UO_211 (O_211,N_8659,N_9537);
nand UO_212 (O_212,N_7642,N_8838);
xnor UO_213 (O_213,N_9676,N_8995);
and UO_214 (O_214,N_9454,N_9364);
nand UO_215 (O_215,N_9016,N_8842);
and UO_216 (O_216,N_9386,N_8199);
nand UO_217 (O_217,N_8519,N_9405);
xnor UO_218 (O_218,N_7654,N_8882);
nand UO_219 (O_219,N_7764,N_7544);
and UO_220 (O_220,N_9706,N_9662);
nand UO_221 (O_221,N_8053,N_7661);
nand UO_222 (O_222,N_9183,N_9252);
or UO_223 (O_223,N_8181,N_7976);
or UO_224 (O_224,N_7501,N_7721);
and UO_225 (O_225,N_7826,N_7502);
nor UO_226 (O_226,N_8865,N_8516);
or UO_227 (O_227,N_9143,N_7870);
and UO_228 (O_228,N_7835,N_8929);
or UO_229 (O_229,N_9118,N_7737);
nor UO_230 (O_230,N_8023,N_8008);
or UO_231 (O_231,N_8056,N_8684);
and UO_232 (O_232,N_8175,N_9552);
nand UO_233 (O_233,N_7767,N_8895);
nor UO_234 (O_234,N_8531,N_8194);
xnor UO_235 (O_235,N_9393,N_7887);
and UO_236 (O_236,N_9069,N_9779);
and UO_237 (O_237,N_8021,N_9989);
nor UO_238 (O_238,N_9907,N_9251);
nor UO_239 (O_239,N_9596,N_7886);
nand UO_240 (O_240,N_9480,N_9304);
nor UO_241 (O_241,N_8423,N_8817);
or UO_242 (O_242,N_8988,N_7631);
or UO_243 (O_243,N_9874,N_9969);
nor UO_244 (O_244,N_9432,N_7875);
and UO_245 (O_245,N_8968,N_7689);
or UO_246 (O_246,N_9925,N_9915);
nand UO_247 (O_247,N_9068,N_8907);
nor UO_248 (O_248,N_7673,N_8063);
xnor UO_249 (O_249,N_7936,N_9448);
nand UO_250 (O_250,N_9121,N_9324);
and UO_251 (O_251,N_9794,N_9059);
or UO_252 (O_252,N_9291,N_7939);
or UO_253 (O_253,N_9028,N_8459);
or UO_254 (O_254,N_8685,N_9022);
xor UO_255 (O_255,N_7790,N_9801);
or UO_256 (O_256,N_7723,N_8923);
and UO_257 (O_257,N_9603,N_7669);
or UO_258 (O_258,N_7622,N_9722);
and UO_259 (O_259,N_8769,N_8541);
and UO_260 (O_260,N_8424,N_9030);
nand UO_261 (O_261,N_7628,N_9963);
or UO_262 (O_262,N_9938,N_9837);
nand UO_263 (O_263,N_8814,N_8786);
or UO_264 (O_264,N_7738,N_9181);
and UO_265 (O_265,N_9799,N_8229);
nor UO_266 (O_266,N_9365,N_7977);
and UO_267 (O_267,N_8903,N_7917);
or UO_268 (O_268,N_7843,N_9586);
nand UO_269 (O_269,N_8942,N_7814);
nand UO_270 (O_270,N_7771,N_8889);
nand UO_271 (O_271,N_7575,N_8810);
nand UO_272 (O_272,N_8481,N_8632);
nor UO_273 (O_273,N_7793,N_7749);
nand UO_274 (O_274,N_9388,N_9340);
nor UO_275 (O_275,N_8688,N_7924);
and UO_276 (O_276,N_7657,N_8603);
or UO_277 (O_277,N_8926,N_9264);
nor UO_278 (O_278,N_7550,N_8580);
or UO_279 (O_279,N_7552,N_9161);
xor UO_280 (O_280,N_8813,N_9495);
nor UO_281 (O_281,N_9447,N_8686);
and UO_282 (O_282,N_7930,N_9728);
nand UO_283 (O_283,N_9247,N_8758);
xor UO_284 (O_284,N_8200,N_8384);
or UO_285 (O_285,N_8404,N_7633);
and UO_286 (O_286,N_9579,N_7832);
nor UO_287 (O_287,N_9097,N_9942);
nor UO_288 (O_288,N_7978,N_9168);
nand UO_289 (O_289,N_7590,N_7980);
and UO_290 (O_290,N_9267,N_9093);
nor UO_291 (O_291,N_9751,N_8653);
nand UO_292 (O_292,N_7663,N_7659);
or UO_293 (O_293,N_7526,N_9904);
and UO_294 (O_294,N_9400,N_8322);
xnor UO_295 (O_295,N_8176,N_8413);
and UO_296 (O_296,N_7944,N_8570);
or UO_297 (O_297,N_7876,N_9711);
and UO_298 (O_298,N_8663,N_8318);
nor UO_299 (O_299,N_9967,N_7778);
or UO_300 (O_300,N_7741,N_9506);
nand UO_301 (O_301,N_9853,N_9821);
nor UO_302 (O_302,N_8853,N_9024);
nand UO_303 (O_303,N_8624,N_8894);
nand UO_304 (O_304,N_8528,N_8720);
nor UO_305 (O_305,N_8264,N_9376);
and UO_306 (O_306,N_8361,N_9733);
and UO_307 (O_307,N_7610,N_9981);
nand UO_308 (O_308,N_9002,N_9833);
nand UO_309 (O_309,N_9216,N_8031);
or UO_310 (O_310,N_9233,N_9019);
nor UO_311 (O_311,N_7605,N_8752);
nor UO_312 (O_312,N_9824,N_8770);
or UO_313 (O_313,N_9529,N_9056);
nor UO_314 (O_314,N_8393,N_9558);
nand UO_315 (O_315,N_9496,N_9029);
and UO_316 (O_316,N_9459,N_7644);
nor UO_317 (O_317,N_7880,N_9993);
nand UO_318 (O_318,N_9348,N_7603);
or UO_319 (O_319,N_9556,N_9158);
xor UO_320 (O_320,N_9857,N_8714);
nand UO_321 (O_321,N_9478,N_8248);
xnor UO_322 (O_322,N_8509,N_9005);
nand UO_323 (O_323,N_8193,N_8730);
and UO_324 (O_324,N_7553,N_8003);
or UO_325 (O_325,N_7671,N_8723);
nand UO_326 (O_326,N_7624,N_7791);
and UO_327 (O_327,N_7905,N_7823);
nand UO_328 (O_328,N_8339,N_7795);
xnor UO_329 (O_329,N_9890,N_7929);
or UO_330 (O_330,N_9658,N_8666);
xnor UO_331 (O_331,N_8771,N_8395);
or UO_332 (O_332,N_9525,N_8891);
or UO_333 (O_333,N_8503,N_8087);
nor UO_334 (O_334,N_8906,N_9106);
nor UO_335 (O_335,N_9929,N_8065);
or UO_336 (O_336,N_8795,N_9013);
nand UO_337 (O_337,N_9044,N_9791);
nand UO_338 (O_338,N_8498,N_8337);
or UO_339 (O_339,N_9684,N_8405);
and UO_340 (O_340,N_9817,N_8024);
nor UO_341 (O_341,N_8657,N_9932);
nor UO_342 (O_342,N_7849,N_9067);
or UO_343 (O_343,N_8005,N_9045);
nor UO_344 (O_344,N_8126,N_9156);
or UO_345 (O_345,N_9631,N_9424);
and UO_346 (O_346,N_9920,N_9725);
nor UO_347 (O_347,N_9749,N_9404);
or UO_348 (O_348,N_8451,N_7899);
nor UO_349 (O_349,N_8477,N_9572);
nor UO_350 (O_350,N_8524,N_9177);
or UO_351 (O_351,N_9955,N_9999);
nand UO_352 (O_352,N_9066,N_8610);
or UO_353 (O_353,N_9577,N_9394);
nand UO_354 (O_354,N_9780,N_7968);
or UO_355 (O_355,N_7884,N_9261);
and UO_356 (O_356,N_8599,N_9750);
and UO_357 (O_357,N_8803,N_7672);
or UO_358 (O_358,N_9887,N_8944);
and UO_359 (O_359,N_8448,N_9311);
and UO_360 (O_360,N_8682,N_9342);
xor UO_361 (O_361,N_8216,N_7931);
xor UO_362 (O_362,N_9661,N_9659);
or UO_363 (O_363,N_7602,N_9951);
xnor UO_364 (O_364,N_8235,N_8616);
nor UO_365 (O_365,N_9061,N_8105);
or UO_366 (O_366,N_8614,N_8517);
nand UO_367 (O_367,N_7516,N_9299);
or UO_368 (O_368,N_9253,N_7920);
and UO_369 (O_369,N_7514,N_9695);
and UO_370 (O_370,N_9325,N_8233);
nor UO_371 (O_371,N_8253,N_8574);
and UO_372 (O_372,N_8418,N_7692);
nand UO_373 (O_373,N_8532,N_7517);
or UO_374 (O_374,N_9563,N_7705);
nand UO_375 (O_375,N_9528,N_7639);
nand UO_376 (O_376,N_8784,N_8943);
or UO_377 (O_377,N_8945,N_9509);
or UO_378 (O_378,N_9703,N_9569);
and UO_379 (O_379,N_8598,N_7632);
and UO_380 (O_380,N_9591,N_8079);
nand UO_381 (O_381,N_9859,N_8417);
nand UO_382 (O_382,N_7871,N_9457);
nand UO_383 (O_383,N_8157,N_8368);
nor UO_384 (O_384,N_7889,N_9673);
nor UO_385 (O_385,N_8511,N_8159);
xor UO_386 (O_386,N_7616,N_8756);
nor UO_387 (O_387,N_8890,N_8293);
or UO_388 (O_388,N_8470,N_7678);
nand UO_389 (O_389,N_9018,N_9578);
nor UO_390 (O_390,N_7593,N_9524);
and UO_391 (O_391,N_8634,N_8766);
and UO_392 (O_392,N_8195,N_7772);
and UO_393 (O_393,N_9209,N_9323);
or UO_394 (O_394,N_9017,N_8504);
xnor UO_395 (O_395,N_7704,N_8680);
or UO_396 (O_396,N_9442,N_7860);
xnor UO_397 (O_397,N_9570,N_7964);
nor UO_398 (O_398,N_9902,N_9788);
and UO_399 (O_399,N_9822,N_9037);
nand UO_400 (O_400,N_7574,N_8256);
nand UO_401 (O_401,N_7942,N_8656);
xor UO_402 (O_402,N_9882,N_7675);
or UO_403 (O_403,N_8388,N_9814);
and UO_404 (O_404,N_8980,N_7617);
and UO_405 (O_405,N_8963,N_9776);
nor UO_406 (O_406,N_8877,N_9420);
or UO_407 (O_407,N_8237,N_8976);
and UO_408 (O_408,N_8520,N_7532);
nor UO_409 (O_409,N_8718,N_9257);
and UO_410 (O_410,N_9897,N_8054);
or UO_411 (O_411,N_7996,N_9521);
and UO_412 (O_412,N_9163,N_9378);
nor UO_413 (O_413,N_7781,N_9609);
nand UO_414 (O_414,N_7867,N_8158);
nand UO_415 (O_415,N_8036,N_9727);
or UO_416 (O_416,N_9852,N_7987);
nor UO_417 (O_417,N_9590,N_8557);
or UO_418 (O_418,N_9743,N_9277);
nor UO_419 (O_419,N_9189,N_7635);
and UO_420 (O_420,N_9437,N_7997);
nand UO_421 (O_421,N_9773,N_8346);
xor UO_422 (O_422,N_9060,N_8131);
and UO_423 (O_423,N_9894,N_8782);
nor UO_424 (O_424,N_7538,N_8699);
and UO_425 (O_425,N_9811,N_8094);
nand UO_426 (O_426,N_7878,N_8828);
and UO_427 (O_427,N_7543,N_7948);
nand UO_428 (O_428,N_9258,N_9622);
nor UO_429 (O_429,N_8156,N_9407);
or UO_430 (O_430,N_9962,N_8660);
nor UO_431 (O_431,N_9145,N_8722);
nor UO_432 (O_432,N_9871,N_9395);
or UO_433 (O_433,N_7776,N_8172);
or UO_434 (O_434,N_8403,N_9338);
nor UO_435 (O_435,N_9628,N_9341);
xor UO_436 (O_436,N_8387,N_8364);
and UO_437 (O_437,N_8749,N_9157);
nand UO_438 (O_438,N_9301,N_8662);
or UO_439 (O_439,N_7726,N_8455);
and UO_440 (O_440,N_9767,N_8076);
nand UO_441 (O_441,N_9958,N_8111);
or UO_442 (O_442,N_8296,N_9977);
nand UO_443 (O_443,N_7925,N_8617);
nor UO_444 (O_444,N_8472,N_9804);
nand UO_445 (O_445,N_9079,N_7833);
nand UO_446 (O_446,N_7511,N_9639);
or UO_447 (O_447,N_8941,N_9458);
nor UO_448 (O_448,N_9055,N_9983);
and UO_449 (O_449,N_8875,N_7918);
nand UO_450 (O_450,N_7589,N_9807);
and UO_451 (O_451,N_8961,N_9169);
nand UO_452 (O_452,N_8390,N_9827);
and UO_453 (O_453,N_8252,N_7665);
or UO_454 (O_454,N_8218,N_9217);
or UO_455 (O_455,N_9976,N_9845);
or UO_456 (O_456,N_8806,N_9550);
and UO_457 (O_457,N_7829,N_8342);
and UO_458 (O_458,N_8802,N_9062);
nand UO_459 (O_459,N_8568,N_9083);
nand UO_460 (O_460,N_7851,N_9273);
xor UO_461 (O_461,N_8140,N_7824);
and UO_462 (O_462,N_9487,N_9803);
nand UO_463 (O_463,N_7649,N_8184);
xnor UO_464 (O_464,N_8552,N_8433);
nand UO_465 (O_465,N_9359,N_8947);
nor UO_466 (O_466,N_8740,N_7608);
nand UO_467 (O_467,N_8826,N_7934);
nand UO_468 (O_468,N_8597,N_9948);
and UO_469 (O_469,N_8590,N_8137);
xnor UO_470 (O_470,N_7706,N_8874);
nand UO_471 (O_471,N_9876,N_8261);
or UO_472 (O_472,N_9909,N_7580);
and UO_473 (O_473,N_7900,N_9191);
and UO_474 (O_474,N_9599,N_7683);
and UO_475 (O_475,N_8737,N_9034);
nand UO_476 (O_476,N_8000,N_8774);
and UO_477 (O_477,N_9007,N_9182);
and UO_478 (O_478,N_9207,N_9286);
nor UO_479 (O_479,N_9781,N_9011);
nand UO_480 (O_480,N_8135,N_7557);
xnor UO_481 (O_481,N_7662,N_9741);
and UO_482 (O_482,N_9327,N_7809);
nand UO_483 (O_483,N_7830,N_7955);
nor UO_484 (O_484,N_9850,N_9982);
or UO_485 (O_485,N_9120,N_7914);
xor UO_486 (O_486,N_8606,N_7636);
or UO_487 (O_487,N_9051,N_9797);
and UO_488 (O_488,N_8291,N_8985);
nand UO_489 (O_489,N_8924,N_9488);
nand UO_490 (O_490,N_8593,N_8402);
or UO_491 (O_491,N_9610,N_9123);
nand UO_492 (O_492,N_7594,N_8335);
nor UO_493 (O_493,N_8192,N_8561);
or UO_494 (O_494,N_8080,N_8128);
xor UO_495 (O_495,N_7513,N_8247);
nor UO_496 (O_496,N_8934,N_9298);
or UO_497 (O_497,N_8348,N_9551);
nand UO_498 (O_498,N_8226,N_7730);
nor UO_499 (O_499,N_9076,N_9071);
nor UO_500 (O_500,N_7740,N_9961);
xor UO_501 (O_501,N_9995,N_7834);
nor UO_502 (O_502,N_9469,N_7890);
or UO_503 (O_503,N_9228,N_8102);
or UO_504 (O_504,N_9472,N_7600);
nor UO_505 (O_505,N_9300,N_8319);
or UO_506 (O_506,N_8975,N_9126);
and UO_507 (O_507,N_8619,N_8755);
xor UO_508 (O_508,N_7784,N_7983);
xor UO_509 (O_509,N_9218,N_8888);
nor UO_510 (O_510,N_8274,N_9358);
xnor UO_511 (O_511,N_8392,N_8868);
and UO_512 (O_512,N_9053,N_9165);
or UO_513 (O_513,N_8761,N_8692);
nand UO_514 (O_514,N_9720,N_8363);
nand UO_515 (O_515,N_9052,N_8640);
nor UO_516 (O_516,N_9414,N_9390);
and UO_517 (O_517,N_8169,N_7775);
xnor UO_518 (O_518,N_7537,N_7932);
nor UO_519 (O_519,N_8480,N_7601);
and UO_520 (O_520,N_7732,N_8867);
or UO_521 (O_521,N_8130,N_9039);
or UO_522 (O_522,N_7536,N_9174);
nand UO_523 (O_523,N_8041,N_9428);
or UO_524 (O_524,N_7935,N_7891);
or UO_525 (O_525,N_9401,N_8837);
nand UO_526 (O_526,N_9530,N_9246);
and UO_527 (O_527,N_8948,N_7587);
nor UO_528 (O_528,N_9514,N_9671);
nand UO_529 (O_529,N_8367,N_8138);
nor UO_530 (O_530,N_9422,N_7746);
nand UO_531 (O_531,N_8977,N_7789);
nor UO_532 (O_532,N_9917,N_8129);
and UO_533 (O_533,N_7743,N_9119);
nand UO_534 (O_534,N_9344,N_9895);
nor UO_535 (O_535,N_8043,N_7842);
nor UO_536 (O_536,N_8821,N_8440);
xnor UO_537 (O_537,N_8805,N_8275);
or UO_538 (O_538,N_8214,N_9867);
and UO_539 (O_539,N_8371,N_9225);
nor UO_540 (O_540,N_7973,N_8112);
xnor UO_541 (O_541,N_7991,N_8466);
nand UO_542 (O_542,N_7837,N_9992);
or UO_543 (O_543,N_8930,N_9035);
nand UO_544 (O_544,N_7810,N_8038);
nand UO_545 (O_545,N_8349,N_9234);
and UO_546 (O_546,N_8971,N_7845);
and UO_547 (O_547,N_7571,N_9861);
and UO_548 (O_548,N_9545,N_8303);
nand UO_549 (O_549,N_7629,N_8914);
or UO_550 (O_550,N_8049,N_7564);
nor UO_551 (O_551,N_9742,N_8628);
nor UO_552 (O_552,N_9935,N_9308);
or UO_553 (O_553,N_8301,N_9138);
nor UO_554 (O_554,N_8777,N_7734);
or UO_555 (O_555,N_7687,N_8521);
and UO_556 (O_556,N_9445,N_7960);
nor UO_557 (O_557,N_9707,N_8010);
or UO_558 (O_558,N_8376,N_8321);
and UO_559 (O_559,N_8979,N_9713);
xnor UO_560 (O_560,N_8972,N_7615);
nand UO_561 (O_561,N_9192,N_8196);
or UO_562 (O_562,N_7926,N_9208);
and UO_563 (O_563,N_8265,N_9107);
and UO_564 (O_564,N_8990,N_8909);
nand UO_565 (O_565,N_9315,N_8589);
nand UO_566 (O_566,N_7569,N_9900);
and UO_567 (O_567,N_7699,N_9892);
nor UO_568 (O_568,N_9584,N_8025);
nor UO_569 (O_569,N_8068,N_8202);
xnor UO_570 (O_570,N_7893,N_8695);
xnor UO_571 (O_571,N_8633,N_8858);
or UO_572 (O_572,N_9499,N_9316);
xnor UO_573 (O_573,N_7680,N_8465);
and UO_574 (O_574,N_9940,N_7694);
or UO_575 (O_575,N_8676,N_8851);
and UO_576 (O_576,N_8855,N_7577);
nand UO_577 (O_577,N_8974,N_7735);
and UO_578 (O_578,N_7591,N_7961);
and UO_579 (O_579,N_9883,N_7962);
xor UO_580 (O_580,N_8779,N_8463);
xnor UO_581 (O_581,N_7679,N_7879);
or UO_582 (O_582,N_9708,N_9690);
nor UO_583 (O_583,N_8673,N_8067);
nor UO_584 (O_584,N_8471,N_9602);
nor UO_585 (O_585,N_9140,N_9238);
or UO_586 (O_586,N_8453,N_8026);
and UO_587 (O_587,N_9846,N_9403);
or UO_588 (O_588,N_9116,N_9945);
nor UO_589 (O_589,N_9283,N_9446);
nor UO_590 (O_590,N_8964,N_8240);
or UO_591 (O_591,N_9914,N_8378);
or UO_592 (O_592,N_9571,N_7674);
or UO_593 (O_593,N_7895,N_8443);
xnor UO_594 (O_594,N_8391,N_9726);
or UO_595 (O_595,N_9379,N_8731);
nor UO_596 (O_596,N_8753,N_8379);
or UO_597 (O_597,N_9353,N_7630);
and UO_598 (O_598,N_8305,N_9643);
nor UO_599 (O_599,N_8514,N_8090);
nand UO_600 (O_600,N_9027,N_9347);
nor UO_601 (O_601,N_7539,N_8242);
xnor UO_602 (O_602,N_7855,N_8572);
nor UO_603 (O_603,N_9753,N_8377);
or UO_604 (O_604,N_7643,N_9137);
or UO_605 (O_605,N_8738,N_8927);
and UO_606 (O_606,N_8872,N_8681);
xnor UO_607 (O_607,N_9760,N_9411);
nor UO_608 (O_608,N_9564,N_9927);
nand UO_609 (O_609,N_9326,N_7541);
nor UO_610 (O_610,N_9715,N_7729);
or UO_611 (O_611,N_9737,N_7716);
and UO_612 (O_612,N_8499,N_8234);
and UO_613 (O_613,N_7813,N_8732);
or UO_614 (O_614,N_8217,N_9680);
and UO_615 (O_615,N_8210,N_9710);
or UO_616 (O_616,N_9368,N_9944);
xor UO_617 (O_617,N_9834,N_8449);
and UO_618 (O_618,N_8835,N_9292);
or UO_619 (O_619,N_9250,N_8427);
nor UO_620 (O_620,N_9354,N_7703);
xor UO_621 (O_621,N_7892,N_8037);
nor UO_622 (O_622,N_8164,N_8432);
and UO_623 (O_623,N_7974,N_7554);
or UO_624 (O_624,N_7763,N_9103);
nor UO_625 (O_625,N_9464,N_9350);
nor UO_626 (O_626,N_9205,N_9618);
or UO_627 (O_627,N_8152,N_7902);
nor UO_628 (O_628,N_9306,N_7988);
nor UO_629 (O_629,N_9612,N_9336);
or UO_630 (O_630,N_8706,N_9000);
and UO_631 (O_631,N_8304,N_9734);
and UO_632 (O_632,N_7909,N_8816);
nor UO_633 (O_633,N_9270,N_7838);
and UO_634 (O_634,N_7766,N_7786);
or UO_635 (O_635,N_7995,N_9607);
nand UO_636 (O_636,N_8409,N_8560);
or UO_637 (O_637,N_7982,N_7572);
xor UO_638 (O_638,N_7588,N_8966);
and UO_639 (O_639,N_8101,N_7780);
nor UO_640 (O_640,N_8679,N_7684);
nand UO_641 (O_641,N_7812,N_8078);
nor UO_642 (O_642,N_9588,N_8074);
nand UO_643 (O_643,N_9280,N_8959);
nand UO_644 (O_644,N_8230,N_8513);
nand UO_645 (O_645,N_8767,N_7525);
and UO_646 (O_646,N_7668,N_8928);
xnor UO_647 (O_647,N_8626,N_8315);
nand UO_648 (O_648,N_8620,N_8359);
or UO_649 (O_649,N_9426,N_8772);
or UO_650 (O_650,N_7648,N_9239);
and UO_651 (O_651,N_8844,N_8565);
and UO_652 (O_652,N_8790,N_8609);
nor UO_653 (O_653,N_9786,N_8124);
nand UO_654 (O_654,N_9784,N_7530);
nand UO_655 (O_655,N_8897,N_8484);
and UO_656 (O_656,N_8636,N_9167);
and UO_657 (O_657,N_9461,N_8045);
nor UO_658 (O_658,N_8209,N_8412);
nand UO_659 (O_659,N_8246,N_9451);
nand UO_660 (O_660,N_8107,N_9465);
and UO_661 (O_661,N_8850,N_7759);
xnor UO_662 (O_662,N_8292,N_8260);
or UO_663 (O_663,N_9047,N_9632);
nor UO_664 (O_664,N_7782,N_8512);
nor UO_665 (O_665,N_7820,N_8071);
nor UO_666 (O_666,N_8436,N_9575);
xnor UO_667 (O_667,N_7604,N_7731);
or UO_668 (O_668,N_9712,N_9793);
and UO_669 (O_669,N_8562,N_9810);
and UO_670 (O_670,N_9757,N_9924);
nor UO_671 (O_671,N_9585,N_9835);
nand UO_672 (O_672,N_9660,N_8314);
nand UO_673 (O_673,N_8206,N_9289);
nor UO_674 (O_674,N_9582,N_9906);
and UO_675 (O_675,N_8326,N_9815);
xor UO_676 (O_676,N_8796,N_8027);
nor UO_677 (O_677,N_9693,N_7545);
and UO_678 (O_678,N_7640,N_9259);
xnor UO_679 (O_679,N_8201,N_7979);
or UO_680 (O_680,N_9533,N_7802);
nor UO_681 (O_681,N_9402,N_9337);
nand UO_682 (O_682,N_9949,N_9832);
nor UO_683 (O_683,N_8707,N_8121);
nor UO_684 (O_684,N_7798,N_8300);
or UO_685 (O_685,N_9162,N_7821);
nor UO_686 (O_686,N_8456,N_9889);
or UO_687 (O_687,N_8151,N_9968);
nor UO_688 (O_688,N_8798,N_9738);
and UO_689 (O_689,N_9666,N_8495);
nand UO_690 (O_690,N_9593,N_9369);
xnor UO_691 (O_691,N_8100,N_7957);
and UO_692 (O_692,N_7509,N_8587);
nor UO_693 (O_693,N_9542,N_9729);
and UO_694 (O_694,N_8250,N_9421);
nand UO_695 (O_695,N_7753,N_7836);
and UO_696 (O_696,N_9064,N_9888);
nand UO_697 (O_697,N_8675,N_8887);
and UO_698 (O_698,N_9219,N_8742);
nand UO_699 (O_699,N_8958,N_8150);
and UO_700 (O_700,N_9274,N_7831);
or UO_701 (O_701,N_9108,N_7714);
xnor UO_702 (O_702,N_9088,N_8998);
nand UO_703 (O_703,N_8165,N_8343);
nor UO_704 (O_704,N_9164,N_9670);
xor UO_705 (O_705,N_9755,N_7817);
and UO_706 (O_706,N_9947,N_9166);
xor UO_707 (O_707,N_9172,N_7805);
xor UO_708 (O_708,N_8953,N_9615);
nor UO_709 (O_709,N_7853,N_9335);
or UO_710 (O_710,N_8046,N_8160);
or UO_711 (O_711,N_9800,N_8604);
nor UO_712 (O_712,N_9310,N_8302);
nand UO_713 (O_713,N_9416,N_8693);
nor UO_714 (O_714,N_9178,N_8340);
and UO_715 (O_715,N_7666,N_8334);
xor UO_716 (O_716,N_8332,N_8398);
nand UO_717 (O_717,N_8015,N_9377);
nand UO_718 (O_718,N_7904,N_7695);
nor UO_719 (O_719,N_9759,N_8096);
xor UO_720 (O_720,N_9544,N_7651);
and UO_721 (O_721,N_8655,N_8385);
or UO_722 (O_722,N_8088,N_9689);
nand UO_723 (O_723,N_9723,N_9078);
and UO_724 (O_724,N_8845,N_8051);
and UO_725 (O_725,N_9627,N_7912);
and UO_726 (O_726,N_8629,N_8185);
xnor UO_727 (O_727,N_9176,N_9081);
and UO_728 (O_728,N_9312,N_7797);
and UO_729 (O_729,N_9674,N_9839);
xor UO_730 (O_730,N_7758,N_9644);
or UO_731 (O_731,N_8820,N_8745);
nor UO_732 (O_732,N_8748,N_8757);
or UO_733 (O_733,N_8989,N_7611);
nor UO_734 (O_734,N_8163,N_9777);
xor UO_735 (O_735,N_8608,N_8672);
nor UO_736 (O_736,N_9990,N_8501);
nand UO_737 (O_737,N_8215,N_7951);
nand UO_738 (O_738,N_9409,N_7534);
and UO_739 (O_739,N_8119,N_9441);
or UO_740 (O_740,N_8818,N_9387);
or UO_741 (O_741,N_7969,N_8081);
and UO_742 (O_742,N_7542,N_9279);
and UO_743 (O_743,N_9285,N_8050);
or UO_744 (O_744,N_8014,N_8117);
or UO_745 (O_745,N_7623,N_9714);
or UO_746 (O_746,N_9758,N_7736);
xor UO_747 (O_747,N_8259,N_9516);
or UO_748 (O_748,N_8701,N_8543);
nand UO_749 (O_749,N_7989,N_9870);
xnor UO_750 (O_750,N_9655,N_8093);
nor UO_751 (O_751,N_8271,N_9687);
and UO_752 (O_752,N_9601,N_8061);
or UO_753 (O_753,N_7559,N_7634);
or UO_754 (O_754,N_8381,N_9589);
xor UO_755 (O_755,N_9493,N_9719);
nand UO_756 (O_756,N_8284,N_9604);
nor UO_757 (O_757,N_8290,N_9792);
and UO_758 (O_758,N_7913,N_9057);
xor UO_759 (O_759,N_7676,N_9139);
and UO_760 (O_760,N_8238,N_9105);
nor UO_761 (O_761,N_9026,N_8573);
or UO_762 (O_762,N_7803,N_8040);
and UO_763 (O_763,N_8896,N_9836);
or UO_764 (O_764,N_9567,N_7874);
nor UO_765 (O_765,N_7916,N_8611);
xnor UO_766 (O_766,N_7688,N_8651);
nand UO_767 (O_767,N_9796,N_8386);
xor UO_768 (O_768,N_9696,N_9190);
or UO_769 (O_769,N_9646,N_8983);
nand UO_770 (O_770,N_9688,N_9752);
nor UO_771 (O_771,N_8383,N_8162);
nand UO_772 (O_772,N_8991,N_8286);
nor UO_773 (O_773,N_8674,N_7515);
and UO_774 (O_774,N_9854,N_9701);
nand UO_775 (O_775,N_9847,N_8496);
nor UO_776 (O_776,N_9543,N_8298);
nor UO_777 (O_777,N_9417,N_9647);
or UO_778 (O_778,N_9931,N_8917);
or UO_779 (O_779,N_8475,N_9595);
xnor UO_780 (O_780,N_9860,N_9032);
nor UO_781 (O_781,N_8362,N_8039);
xnor UO_782 (O_782,N_7808,N_8347);
nor UO_783 (O_783,N_8113,N_9975);
xnor UO_784 (O_784,N_9681,N_7864);
and UO_785 (O_785,N_9928,N_8374);
and UO_786 (O_786,N_9204,N_8141);
nand UO_787 (O_787,N_9101,N_8434);
xor UO_788 (O_788,N_8751,N_7990);
and UO_789 (O_789,N_9973,N_7562);
nor UO_790 (O_790,N_8344,N_8994);
and UO_791 (O_791,N_7898,N_7647);
or UO_792 (O_792,N_8822,N_9468);
nand UO_793 (O_793,N_8925,N_9100);
and UO_794 (O_794,N_9397,N_8146);
nor UO_795 (O_795,N_9916,N_9598);
nor UO_796 (O_796,N_8785,N_9012);
nor UO_797 (O_797,N_8920,N_8908);
or UO_798 (O_798,N_9820,N_9746);
and UO_799 (O_799,N_8936,N_7818);
nor UO_800 (O_800,N_9560,N_8211);
or UO_801 (O_801,N_9745,N_7965);
or UO_802 (O_802,N_7655,N_8812);
nand UO_803 (O_803,N_8114,N_9559);
and UO_804 (O_804,N_8904,N_7745);
nor UO_805 (O_805,N_8754,N_8535);
or UO_806 (O_806,N_9483,N_8569);
and UO_807 (O_807,N_9913,N_7840);
nor UO_808 (O_808,N_9275,N_9736);
or UO_809 (O_809,N_9109,N_9266);
nand UO_810 (O_810,N_9427,N_8506);
xnor UO_811 (O_811,N_9307,N_9978);
nand UO_812 (O_812,N_8622,N_9941);
nand UO_813 (O_813,N_8308,N_9485);
xnor UO_814 (O_814,N_9823,N_8396);
nand UO_815 (O_815,N_7839,N_8186);
nor UO_816 (O_816,N_7911,N_8950);
or UO_817 (O_817,N_7785,N_8397);
nor UO_818 (O_818,N_7952,N_9592);
nor UO_819 (O_819,N_9664,N_9269);
or UO_820 (O_820,N_8696,N_7523);
nand UO_821 (O_821,N_7685,N_8747);
and UO_822 (O_822,N_8883,N_7994);
xor UO_823 (O_823,N_9322,N_7561);
and UO_824 (O_824,N_8760,N_9382);
nor UO_825 (O_825,N_7919,N_7844);
and UO_826 (O_826,N_8647,N_7558);
or UO_827 (O_827,N_9095,N_9180);
and UO_828 (O_828,N_8365,N_9972);
nor UO_829 (O_829,N_8893,N_7941);
nand UO_830 (O_830,N_8848,N_8646);
nand UO_831 (O_831,N_8508,N_9851);
nand UO_832 (O_832,N_9594,N_9362);
nand UO_833 (O_833,N_8938,N_9329);
and UO_834 (O_834,N_8783,N_9094);
or UO_835 (O_835,N_8576,N_8276);
nand UO_836 (O_836,N_9085,N_8665);
nor UO_837 (O_837,N_9434,N_9360);
nor UO_838 (O_838,N_7921,N_8705);
and UO_839 (O_839,N_9798,N_8143);
and UO_840 (O_840,N_9245,N_9957);
or UO_841 (O_841,N_7762,N_8762);
nor UO_842 (O_842,N_8408,N_7681);
or UO_843 (O_843,N_7992,N_8497);
nor UO_844 (O_844,N_9196,N_7725);
and UO_845 (O_845,N_8115,N_9918);
nor UO_846 (O_846,N_9272,N_9546);
and UO_847 (O_847,N_7620,N_9389);
nor UO_848 (O_848,N_8916,N_8581);
nand UO_849 (O_849,N_7894,N_9717);
or UO_850 (O_850,N_9086,N_7637);
and UO_851 (O_851,N_8739,N_7686);
nand UO_852 (O_852,N_9135,N_7906);
or UO_853 (O_853,N_9321,N_8551);
and UO_854 (O_854,N_8605,N_8549);
or UO_855 (O_855,N_8155,N_9131);
nand UO_856 (O_856,N_8085,N_8537);
and UO_857 (O_857,N_8108,N_9374);
xnor UO_858 (O_858,N_8515,N_9084);
nand UO_859 (O_859,N_7863,N_7804);
nor UO_860 (O_860,N_7827,N_7922);
or UO_861 (O_861,N_9576,N_8254);
or UO_862 (O_862,N_8563,N_9371);
or UO_863 (O_863,N_8553,N_9430);
or UO_864 (O_864,N_8529,N_8464);
and UO_865 (O_865,N_9912,N_9295);
nand UO_866 (O_866,N_9361,N_8149);
nor UO_867 (O_867,N_7533,N_9149);
and UO_868 (O_868,N_8861,N_9985);
and UO_869 (O_869,N_9505,N_8876);
nand UO_870 (O_870,N_9663,N_7709);
nand UO_871 (O_871,N_9790,N_9486);
nand UO_872 (O_872,N_9731,N_8650);
and UO_873 (O_873,N_9816,N_8070);
or UO_874 (O_874,N_9555,N_9413);
or UO_875 (O_875,N_7757,N_7664);
nand UO_876 (O_876,N_8807,N_8095);
nand UO_877 (O_877,N_9966,N_8134);
or UO_878 (O_878,N_8585,N_7660);
nand UO_879 (O_879,N_8236,N_8373);
or UO_880 (O_880,N_8913,N_9089);
nand UO_881 (O_881,N_7595,N_8118);
or UO_882 (O_882,N_8122,N_8429);
nor UO_883 (O_883,N_8069,N_9526);
nand UO_884 (O_884,N_9230,N_9425);
nor UO_885 (O_885,N_8273,N_7719);
and UO_886 (O_886,N_9113,N_7882);
xnor UO_887 (O_887,N_7859,N_9150);
or UO_888 (O_888,N_7563,N_7963);
nand UO_889 (O_889,N_8992,N_8241);
xor UO_890 (O_890,N_8353,N_8638);
and UO_891 (O_891,N_7801,N_8154);
or UO_892 (O_892,N_8147,N_7522);
nand UO_893 (O_893,N_9683,N_9937);
or UO_894 (O_894,N_8642,N_7656);
and UO_895 (O_895,N_8973,N_8245);
nand UO_896 (O_896,N_8171,N_9950);
or UO_897 (O_897,N_9303,N_8006);
and UO_898 (O_898,N_8540,N_9111);
and UO_899 (O_899,N_9206,N_9004);
xnor UO_900 (O_900,N_9911,N_8915);
or UO_901 (O_901,N_7583,N_8431);
or UO_902 (O_902,N_7861,N_8937);
nor UO_903 (O_903,N_9763,N_9124);
and UO_904 (O_904,N_8450,N_9640);
or UO_905 (O_905,N_9769,N_8873);
or UO_906 (O_906,N_9141,N_9974);
or UO_907 (O_907,N_8579,N_9732);
and UO_908 (O_908,N_9244,N_8612);
nor UO_909 (O_909,N_8280,N_9764);
nor UO_910 (O_910,N_7504,N_9919);
nand UO_911 (O_911,N_9697,N_8430);
nor UO_912 (O_912,N_7713,N_7865);
and UO_913 (O_913,N_9896,N_9580);
and UO_914 (O_914,N_7682,N_9021);
and UO_915 (O_915,N_8360,N_8892);
and UO_916 (O_916,N_9573,N_9186);
nor UO_917 (O_917,N_9986,N_9248);
and UO_918 (O_918,N_9500,N_9549);
and UO_919 (O_919,N_9623,N_8223);
nand UO_920 (O_920,N_7527,N_9367);
and UO_921 (O_921,N_8232,N_8710);
xnor UO_922 (O_922,N_8698,N_9491);
nor UO_923 (O_923,N_9979,N_7512);
nand UO_924 (O_924,N_9682,N_9939);
nor UO_925 (O_925,N_8792,N_7710);
and UO_926 (O_926,N_8824,N_9838);
and UO_927 (O_927,N_8717,N_9077);
and UO_928 (O_928,N_7946,N_7765);
nor UO_929 (O_929,N_8270,N_9399);
and UO_930 (O_930,N_9709,N_8109);
and UO_931 (O_931,N_8996,N_9475);
and UO_932 (O_932,N_9271,N_9117);
and UO_933 (O_933,N_8057,N_7881);
nor UO_934 (O_934,N_9616,N_9649);
nor UO_935 (O_935,N_9515,N_9331);
xor UO_936 (O_936,N_9553,N_8708);
or UO_937 (O_937,N_8691,N_9293);
xor UO_938 (O_938,N_9317,N_7850);
and UO_939 (O_939,N_8898,N_9319);
and UO_940 (O_940,N_7531,N_9241);
xor UO_941 (O_941,N_9613,N_7819);
or UO_942 (O_942,N_8969,N_8811);
or UO_943 (O_943,N_8677,N_8458);
or UO_944 (O_944,N_8993,N_8116);
or UO_945 (O_945,N_9185,N_8833);
and UO_946 (O_946,N_9449,N_8630);
nor UO_947 (O_947,N_8839,N_9318);
nor UO_948 (O_948,N_8283,N_9243);
nor UO_949 (O_949,N_9229,N_9825);
and UO_950 (O_950,N_8416,N_8860);
nor UO_951 (O_951,N_9170,N_9936);
and UO_952 (O_952,N_9795,N_8438);
nand UO_953 (O_953,N_8227,N_9700);
or UO_954 (O_954,N_9872,N_9211);
nor UO_955 (O_955,N_8734,N_9510);
and UO_956 (O_956,N_8664,N_8970);
xnor UO_957 (O_957,N_8009,N_7519);
nor UO_958 (O_958,N_8287,N_8307);
and UO_959 (O_959,N_8372,N_9583);
and UO_960 (O_960,N_9048,N_7927);
nand UO_961 (O_961,N_8375,N_8846);
nor UO_962 (O_962,N_9768,N_8727);
and UO_963 (O_963,N_9840,N_9235);
nor UO_964 (O_964,N_9875,N_7788);
nor UO_965 (O_965,N_8794,N_8954);
or UO_966 (O_966,N_9450,N_8857);
and UO_967 (O_967,N_9672,N_7928);
nor UO_968 (O_968,N_9611,N_8775);
nor UO_969 (O_969,N_8168,N_7667);
and UO_970 (O_970,N_8133,N_9431);
and UO_971 (O_971,N_9645,N_9880);
or UO_972 (O_972,N_9866,N_8982);
nor UO_973 (O_973,N_9899,N_9242);
and UO_974 (O_974,N_7597,N_8700);
nor UO_975 (O_975,N_7560,N_8871);
nor UO_976 (O_976,N_9160,N_8823);
and UO_977 (O_977,N_7592,N_9621);
nand UO_978 (O_978,N_7877,N_9231);
xnor UO_979 (O_979,N_8773,N_7769);
xor UO_980 (O_980,N_8173,N_8596);
and UO_981 (O_981,N_7868,N_8505);
nor UO_982 (O_982,N_9479,N_8558);
and UO_983 (O_983,N_9501,N_9539);
nand UO_984 (O_984,N_7567,N_9619);
and UO_985 (O_985,N_7576,N_8946);
nand UO_986 (O_986,N_9842,N_8197);
and UO_987 (O_987,N_8479,N_8435);
and UO_988 (O_988,N_9212,N_9561);
xor UO_989 (O_989,N_9642,N_8880);
or UO_990 (O_990,N_9885,N_9481);
or UO_991 (O_991,N_7625,N_9614);
or UO_992 (O_992,N_9508,N_9073);
and UO_993 (O_993,N_9001,N_9236);
and UO_994 (O_994,N_7582,N_8962);
and UO_995 (O_995,N_8836,N_7565);
and UO_996 (O_996,N_8768,N_9476);
or UO_997 (O_997,N_8548,N_8594);
nand UO_998 (O_998,N_9132,N_9309);
nor UO_999 (O_999,N_8668,N_8719);
nand UO_1000 (O_1000,N_8645,N_9278);
nor UO_1001 (O_1001,N_8190,N_9808);
nor UO_1002 (O_1002,N_8900,N_8336);
and UO_1003 (O_1003,N_7985,N_8120);
nor UO_1004 (O_1004,N_8059,N_7547);
nor UO_1005 (O_1005,N_9657,N_9923);
or UO_1006 (O_1006,N_9147,N_9438);
or UO_1007 (O_1007,N_9858,N_9873);
or UO_1008 (O_1008,N_9042,N_8956);
xor UO_1009 (O_1009,N_9855,N_8582);
nor UO_1010 (O_1010,N_7822,N_8469);
or UO_1011 (O_1011,N_7584,N_8799);
nor UO_1012 (O_1012,N_9805,N_9517);
and UO_1013 (O_1013,N_8689,N_9213);
and UO_1014 (O_1014,N_7506,N_8144);
nand UO_1015 (O_1015,N_9829,N_9406);
nand UO_1016 (O_1016,N_9629,N_7715);
nand UO_1017 (O_1017,N_9641,N_8461);
or UO_1018 (O_1018,N_7556,N_9063);
or UO_1019 (O_1019,N_8457,N_9396);
xor UO_1020 (O_1020,N_9038,N_8724);
xnor UO_1021 (O_1021,N_8191,N_7650);
and UO_1022 (O_1022,N_8487,N_9497);
or UO_1023 (O_1023,N_7806,N_9133);
nand UO_1024 (O_1024,N_9891,N_8460);
and UO_1025 (O_1025,N_8736,N_8330);
and UO_1026 (O_1026,N_9226,N_8825);
and UO_1027 (O_1027,N_8525,N_7907);
nand UO_1028 (O_1028,N_7999,N_8106);
or UO_1029 (O_1029,N_8219,N_9718);
and UO_1030 (O_1030,N_7792,N_8831);
or UO_1031 (O_1031,N_8643,N_9087);
nand UO_1032 (O_1032,N_9096,N_8345);
xor UO_1033 (O_1033,N_8382,N_9532);
and UO_1034 (O_1034,N_8545,N_9104);
and UO_1035 (O_1035,N_8711,N_8829);
nand UO_1036 (O_1036,N_9439,N_8399);
nor UO_1037 (O_1037,N_8299,N_9557);
nand UO_1038 (O_1038,N_9232,N_8425);
nor UO_1039 (O_1039,N_9511,N_7718);
nand UO_1040 (O_1040,N_7700,N_8542);
xnor UO_1041 (O_1041,N_8550,N_9562);
nor UO_1042 (O_1042,N_7612,N_9806);
nand UO_1043 (O_1043,N_9624,N_9625);
and UO_1044 (O_1044,N_7998,N_9863);
or UO_1045 (O_1045,N_8295,N_9023);
nand UO_1046 (O_1046,N_8491,N_9074);
xor UO_1047 (O_1047,N_9856,N_9922);
xor UO_1048 (O_1048,N_7742,N_9901);
xor UO_1049 (O_1049,N_9965,N_8886);
nand UO_1050 (O_1050,N_8703,N_9356);
and UO_1051 (O_1051,N_9194,N_9281);
xnor UO_1052 (O_1052,N_9744,N_7599);
nand UO_1053 (O_1053,N_9355,N_9994);
nor UO_1054 (O_1054,N_8179,N_8743);
nor UO_1055 (O_1055,N_7728,N_9370);
nor UO_1056 (O_1056,N_9398,N_7841);
and UO_1057 (O_1057,N_8733,N_9201);
and UO_1058 (O_1058,N_8744,N_9366);
nand UO_1059 (O_1059,N_9412,N_9626);
nor UO_1060 (O_1060,N_8411,N_9620);
and UO_1061 (O_1061,N_9090,N_9956);
nand UO_1062 (O_1062,N_8082,N_8483);
xor UO_1063 (O_1063,N_8910,N_8827);
or UO_1064 (O_1064,N_7846,N_8297);
nand UO_1065 (O_1065,N_8011,N_9187);
nor UO_1066 (O_1066,N_9630,N_8022);
nand UO_1067 (O_1067,N_8442,N_8485);
nor UO_1068 (O_1068,N_9677,N_8899);
nand UO_1069 (O_1069,N_8935,N_8502);
and UO_1070 (O_1070,N_9685,N_9482);
nand UO_1071 (O_1071,N_9531,N_9775);
nor UO_1072 (O_1072,N_8064,N_9877);
or UO_1073 (O_1073,N_8267,N_9223);
or UO_1074 (O_1074,N_7783,N_9122);
or UO_1075 (O_1075,N_8729,N_8220);
and UO_1076 (O_1076,N_9003,N_8715);
and UO_1077 (O_1077,N_9153,N_9263);
or UO_1078 (O_1078,N_7888,N_7958);
xor UO_1079 (O_1079,N_8243,N_8441);
or UO_1080 (O_1080,N_8869,N_7750);
and UO_1081 (O_1081,N_8591,N_8566);
and UO_1082 (O_1082,N_8690,N_8780);
or UO_1083 (O_1083,N_9694,N_9638);
and UO_1084 (O_1084,N_9210,N_7984);
nand UO_1085 (O_1085,N_9653,N_8957);
nor UO_1086 (O_1086,N_9819,N_8426);
nand UO_1087 (O_1087,N_8801,N_9179);
and UO_1088 (O_1088,N_9566,N_9886);
nor UO_1089 (O_1089,N_8437,N_8357);
or UO_1090 (O_1090,N_8544,N_9195);
or UO_1091 (O_1091,N_7754,N_8476);
nand UO_1092 (O_1092,N_9320,N_8571);
or UO_1093 (O_1093,N_8020,N_8161);
or UO_1094 (O_1094,N_7586,N_8327);
or UO_1095 (O_1095,N_9408,N_7702);
or UO_1096 (O_1096,N_9930,N_9648);
or UO_1097 (O_1097,N_9372,N_9778);
nand UO_1098 (O_1098,N_8601,N_8350);
nor UO_1099 (O_1099,N_8741,N_9910);
nor UO_1100 (O_1100,N_8613,N_9903);
or UO_1101 (O_1101,N_8547,N_8089);
and UO_1102 (O_1102,N_9702,N_8212);
nand UO_1103 (O_1103,N_8016,N_8492);
xor UO_1104 (O_1104,N_8986,N_9691);
xor UO_1105 (O_1105,N_9288,N_9173);
and UO_1106 (O_1106,N_9058,N_8414);
nor UO_1107 (O_1107,N_8249,N_8066);
nand UO_1108 (O_1108,N_8840,N_8325);
nor UO_1109 (O_1109,N_8635,N_7551);
xor UO_1110 (O_1110,N_7573,N_8052);
and UO_1111 (O_1111,N_8187,N_8029);
or UO_1112 (O_1112,N_8380,N_9456);
nor UO_1113 (O_1113,N_9843,N_7546);
and UO_1114 (O_1114,N_7787,N_7521);
and UO_1115 (O_1115,N_9098,N_9334);
nor UO_1116 (O_1116,N_7953,N_7883);
nor UO_1117 (O_1117,N_9385,N_7744);
nor UO_1118 (O_1118,N_9785,N_8048);
nand UO_1119 (O_1119,N_8627,N_8530);
and UO_1120 (O_1120,N_7724,N_9953);
and UO_1121 (O_1121,N_8032,N_8257);
nor UO_1122 (O_1122,N_8921,N_8142);
xnor UO_1123 (O_1123,N_8595,N_9669);
nand UO_1124 (O_1124,N_8474,N_9214);
or UO_1125 (O_1125,N_9652,N_7585);
nand UO_1126 (O_1126,N_9462,N_9452);
nor UO_1127 (O_1127,N_8859,N_7621);
nor UO_1128 (O_1128,N_8310,N_7937);
nor UO_1129 (O_1129,N_9215,N_9054);
nor UO_1130 (O_1130,N_7774,N_9102);
nand UO_1131 (O_1131,N_8978,N_9502);
nor UO_1132 (O_1132,N_8278,N_9148);
or UO_1133 (O_1133,N_7896,N_8852);
nor UO_1134 (O_1134,N_8389,N_9765);
and UO_1135 (O_1135,N_7670,N_7677);
xor UO_1136 (O_1136,N_8415,N_8282);
or UO_1137 (O_1137,N_9520,N_8444);
nor UO_1138 (O_1138,N_9470,N_9151);
and UO_1139 (O_1139,N_7755,N_9600);
and UO_1140 (O_1140,N_8263,N_7773);
nor UO_1141 (O_1141,N_8331,N_9735);
nor UO_1142 (O_1142,N_8060,N_9971);
nand UO_1143 (O_1143,N_8661,N_9240);
nor UO_1144 (O_1144,N_8251,N_9046);
and UO_1145 (O_1145,N_7915,N_7910);
or UO_1146 (O_1146,N_9265,N_7535);
nor UO_1147 (O_1147,N_8125,N_8864);
nand UO_1148 (O_1148,N_9155,N_8843);
nor UO_1149 (O_1149,N_7693,N_8486);
nand UO_1150 (O_1150,N_8329,N_9302);
nand UO_1151 (O_1151,N_8473,N_8866);
and UO_1152 (O_1152,N_8012,N_8279);
or UO_1153 (O_1153,N_7966,N_9152);
nand UO_1154 (O_1154,N_8205,N_9535);
or UO_1155 (O_1155,N_8536,N_9943);
xor UO_1156 (O_1156,N_9996,N_8019);
nor UO_1157 (O_1157,N_9256,N_9771);
or UO_1158 (O_1158,N_9988,N_9634);
nand UO_1159 (O_1159,N_8716,N_9868);
and UO_1160 (O_1160,N_9313,N_9198);
nand UO_1161 (O_1161,N_8269,N_8999);
or UO_1162 (O_1162,N_9142,N_8567);
nor UO_1163 (O_1163,N_8007,N_9025);
or UO_1164 (O_1164,N_8207,N_8231);
and UO_1165 (O_1165,N_7697,N_9565);
or UO_1166 (O_1166,N_7779,N_8033);
or UO_1167 (O_1167,N_7885,N_8454);
xor UO_1168 (O_1168,N_7701,N_9010);
and UO_1169 (O_1169,N_8902,N_8478);
nor UO_1170 (O_1170,N_7986,N_8439);
nor UO_1171 (O_1171,N_9581,N_9202);
or UO_1172 (O_1172,N_9041,N_8320);
nand UO_1173 (O_1173,N_8952,N_8997);
nor UO_1174 (O_1174,N_9435,N_7653);
nand UO_1175 (O_1175,N_9898,N_9489);
nand UO_1176 (O_1176,N_8791,N_9519);
and UO_1177 (O_1177,N_8180,N_8351);
xor UO_1178 (O_1178,N_9667,N_7549);
and UO_1179 (O_1179,N_8446,N_8166);
nand UO_1180 (O_1180,N_8793,N_8203);
or UO_1181 (O_1181,N_9284,N_9453);
nand UO_1182 (O_1182,N_8789,N_9756);
or UO_1183 (O_1183,N_7548,N_9970);
xor UO_1184 (O_1184,N_7866,N_8058);
and UO_1185 (O_1185,N_7943,N_8667);
and UO_1186 (O_1186,N_9699,N_8294);
or UO_1187 (O_1187,N_8123,N_9964);
nand UO_1188 (O_1188,N_8468,N_8028);
nand UO_1189 (O_1189,N_8018,N_9460);
xnor UO_1190 (O_1190,N_8841,N_9665);
and UO_1191 (O_1191,N_9339,N_9072);
and UO_1192 (O_1192,N_9541,N_8678);
and UO_1193 (O_1193,N_9721,N_8369);
nand UO_1194 (O_1194,N_8285,N_8309);
nand UO_1195 (O_1195,N_7626,N_8222);
nor UO_1196 (O_1196,N_8919,N_8338);
or UO_1197 (O_1197,N_8776,N_9467);
or UO_1198 (O_1198,N_7816,N_8178);
nor UO_1199 (O_1199,N_9762,N_8086);
nand UO_1200 (O_1200,N_8224,N_9554);
nor UO_1201 (O_1201,N_8637,N_9352);
nand UO_1202 (O_1202,N_8323,N_9926);
nor UO_1203 (O_1203,N_8765,N_8911);
and UO_1204 (O_1204,N_7540,N_8073);
nor UO_1205 (O_1205,N_8830,N_7777);
and UO_1206 (O_1206,N_8533,N_8002);
and UO_1207 (O_1207,N_7613,N_8490);
and UO_1208 (O_1208,N_7598,N_9043);
or UO_1209 (O_1209,N_9114,N_9091);
nor UO_1210 (O_1210,N_8370,N_8559);
nand UO_1211 (O_1211,N_8652,N_9831);
and UO_1212 (O_1212,N_8352,N_9523);
and UO_1213 (O_1213,N_8960,N_9802);
and UO_1214 (O_1214,N_8931,N_7733);
or UO_1215 (O_1215,N_7950,N_7524);
or UO_1216 (O_1216,N_7581,N_9200);
nand UO_1217 (O_1217,N_8035,N_8272);
xnor UO_1218 (O_1218,N_7510,N_9125);
nor UO_1219 (O_1219,N_8183,N_8809);
nor UO_1220 (O_1220,N_8452,N_9144);
nor UO_1221 (O_1221,N_9828,N_7646);
nand UO_1222 (O_1222,N_9679,N_9065);
nand UO_1223 (O_1223,N_8084,N_9146);
xnor UO_1224 (O_1224,N_9129,N_8800);
or UO_1225 (O_1225,N_9282,N_9617);
nor UO_1226 (O_1226,N_8313,N_8725);
and UO_1227 (O_1227,N_9998,N_8189);
and UO_1228 (O_1228,N_7529,N_7638);
xnor UO_1229 (O_1229,N_9294,N_8420);
xnor UO_1230 (O_1230,N_7897,N_8324);
nor UO_1231 (O_1231,N_9075,N_8077);
and UO_1232 (O_1232,N_9636,N_9296);
and UO_1233 (O_1233,N_7768,N_8804);
nand UO_1234 (O_1234,N_9443,N_8967);
nor UO_1235 (O_1235,N_9605,N_8333);
and UO_1236 (O_1236,N_9436,N_8421);
and UO_1237 (O_1237,N_8153,N_7508);
xor UO_1238 (O_1238,N_8618,N_9692);
and UO_1239 (O_1239,N_8174,N_8584);
and UO_1240 (O_1240,N_8410,N_9675);
or UO_1241 (O_1241,N_8228,N_9015);
nor UO_1242 (O_1242,N_8538,N_8493);
nor UO_1243 (O_1243,N_7756,N_8225);
nor UO_1244 (O_1244,N_8004,N_8797);
or UO_1245 (O_1245,N_8400,N_9351);
nor UO_1246 (O_1246,N_9512,N_8933);
and UO_1247 (O_1247,N_7712,N_8354);
and UO_1248 (O_1248,N_9878,N_8965);
or UO_1249 (O_1249,N_9020,N_9418);
or UO_1250 (O_1250,N_8027,N_9006);
nand UO_1251 (O_1251,N_8782,N_7841);
nor UO_1252 (O_1252,N_9536,N_9479);
or UO_1253 (O_1253,N_7927,N_8056);
nand UO_1254 (O_1254,N_8885,N_8510);
nand UO_1255 (O_1255,N_9881,N_9243);
and UO_1256 (O_1256,N_7627,N_8312);
or UO_1257 (O_1257,N_9610,N_9478);
or UO_1258 (O_1258,N_9219,N_8368);
xor UO_1259 (O_1259,N_7987,N_8762);
or UO_1260 (O_1260,N_8798,N_7848);
nor UO_1261 (O_1261,N_9841,N_9828);
and UO_1262 (O_1262,N_9744,N_8841);
xor UO_1263 (O_1263,N_9660,N_8516);
nor UO_1264 (O_1264,N_8342,N_8611);
nor UO_1265 (O_1265,N_8066,N_7849);
nand UO_1266 (O_1266,N_8390,N_8555);
or UO_1267 (O_1267,N_9125,N_9145);
xor UO_1268 (O_1268,N_9127,N_7625);
xor UO_1269 (O_1269,N_9473,N_9526);
nand UO_1270 (O_1270,N_8927,N_9375);
nor UO_1271 (O_1271,N_9145,N_8304);
nor UO_1272 (O_1272,N_9578,N_9380);
nand UO_1273 (O_1273,N_9920,N_8466);
nor UO_1274 (O_1274,N_7663,N_8810);
nand UO_1275 (O_1275,N_9850,N_8616);
nand UO_1276 (O_1276,N_7537,N_9696);
nand UO_1277 (O_1277,N_9764,N_9479);
and UO_1278 (O_1278,N_9669,N_8387);
and UO_1279 (O_1279,N_7815,N_8334);
or UO_1280 (O_1280,N_7546,N_9816);
or UO_1281 (O_1281,N_8774,N_9434);
and UO_1282 (O_1282,N_9325,N_8557);
nand UO_1283 (O_1283,N_9735,N_8134);
or UO_1284 (O_1284,N_8244,N_9051);
or UO_1285 (O_1285,N_9860,N_9729);
or UO_1286 (O_1286,N_7624,N_9799);
or UO_1287 (O_1287,N_9953,N_8988);
nand UO_1288 (O_1288,N_8585,N_9662);
nand UO_1289 (O_1289,N_9061,N_7803);
nand UO_1290 (O_1290,N_9998,N_7691);
nand UO_1291 (O_1291,N_8552,N_8146);
or UO_1292 (O_1292,N_8701,N_8315);
nand UO_1293 (O_1293,N_8570,N_9924);
nand UO_1294 (O_1294,N_8535,N_9209);
or UO_1295 (O_1295,N_8787,N_7913);
nand UO_1296 (O_1296,N_8979,N_9232);
or UO_1297 (O_1297,N_9784,N_8100);
and UO_1298 (O_1298,N_8122,N_9300);
and UO_1299 (O_1299,N_9519,N_8877);
and UO_1300 (O_1300,N_8776,N_9972);
or UO_1301 (O_1301,N_9266,N_9535);
nand UO_1302 (O_1302,N_9850,N_8796);
and UO_1303 (O_1303,N_9859,N_9280);
nor UO_1304 (O_1304,N_9784,N_7729);
nand UO_1305 (O_1305,N_8209,N_8409);
or UO_1306 (O_1306,N_9848,N_7698);
or UO_1307 (O_1307,N_8850,N_9137);
or UO_1308 (O_1308,N_9960,N_9589);
and UO_1309 (O_1309,N_9171,N_9475);
nor UO_1310 (O_1310,N_9777,N_9956);
or UO_1311 (O_1311,N_8957,N_8850);
and UO_1312 (O_1312,N_8950,N_7559);
nand UO_1313 (O_1313,N_8132,N_9080);
or UO_1314 (O_1314,N_9206,N_7865);
or UO_1315 (O_1315,N_9647,N_7788);
and UO_1316 (O_1316,N_7959,N_9222);
nand UO_1317 (O_1317,N_7766,N_8179);
and UO_1318 (O_1318,N_9459,N_8825);
nand UO_1319 (O_1319,N_9159,N_8291);
nand UO_1320 (O_1320,N_8837,N_8623);
nor UO_1321 (O_1321,N_8920,N_7883);
nor UO_1322 (O_1322,N_8858,N_8282);
nor UO_1323 (O_1323,N_7865,N_9138);
and UO_1324 (O_1324,N_9901,N_8367);
and UO_1325 (O_1325,N_8475,N_9159);
and UO_1326 (O_1326,N_9465,N_8102);
or UO_1327 (O_1327,N_8570,N_8064);
or UO_1328 (O_1328,N_7843,N_8272);
nor UO_1329 (O_1329,N_9110,N_9642);
and UO_1330 (O_1330,N_7786,N_9012);
nand UO_1331 (O_1331,N_8441,N_9389);
or UO_1332 (O_1332,N_9158,N_9942);
and UO_1333 (O_1333,N_9994,N_9572);
nor UO_1334 (O_1334,N_8722,N_8768);
and UO_1335 (O_1335,N_8044,N_8757);
and UO_1336 (O_1336,N_8851,N_8117);
and UO_1337 (O_1337,N_8523,N_9637);
or UO_1338 (O_1338,N_8601,N_8421);
nor UO_1339 (O_1339,N_9930,N_9505);
or UO_1340 (O_1340,N_8766,N_8175);
nand UO_1341 (O_1341,N_7602,N_9167);
nor UO_1342 (O_1342,N_7800,N_8650);
or UO_1343 (O_1343,N_7899,N_9579);
nand UO_1344 (O_1344,N_8819,N_8627);
and UO_1345 (O_1345,N_7809,N_8578);
nor UO_1346 (O_1346,N_8734,N_7822);
or UO_1347 (O_1347,N_9745,N_8744);
nor UO_1348 (O_1348,N_9780,N_8131);
nand UO_1349 (O_1349,N_8526,N_7958);
and UO_1350 (O_1350,N_7795,N_7906);
nor UO_1351 (O_1351,N_8564,N_7530);
or UO_1352 (O_1352,N_7927,N_9189);
nor UO_1353 (O_1353,N_8889,N_9925);
or UO_1354 (O_1354,N_9810,N_8017);
nor UO_1355 (O_1355,N_8882,N_9405);
and UO_1356 (O_1356,N_8617,N_9458);
and UO_1357 (O_1357,N_8081,N_7718);
nor UO_1358 (O_1358,N_9311,N_9392);
or UO_1359 (O_1359,N_8793,N_8639);
and UO_1360 (O_1360,N_9643,N_7631);
xnor UO_1361 (O_1361,N_9852,N_8838);
nand UO_1362 (O_1362,N_8405,N_9384);
and UO_1363 (O_1363,N_9037,N_9523);
nor UO_1364 (O_1364,N_9714,N_9390);
nor UO_1365 (O_1365,N_9354,N_9360);
nor UO_1366 (O_1366,N_8207,N_8894);
nor UO_1367 (O_1367,N_9416,N_8380);
or UO_1368 (O_1368,N_7969,N_9411);
and UO_1369 (O_1369,N_8148,N_9356);
xor UO_1370 (O_1370,N_8604,N_7512);
nand UO_1371 (O_1371,N_8224,N_8250);
or UO_1372 (O_1372,N_8796,N_8749);
nand UO_1373 (O_1373,N_8964,N_8766);
and UO_1374 (O_1374,N_8887,N_9318);
or UO_1375 (O_1375,N_7673,N_8508);
or UO_1376 (O_1376,N_7629,N_9125);
or UO_1377 (O_1377,N_9550,N_9700);
and UO_1378 (O_1378,N_8745,N_8252);
or UO_1379 (O_1379,N_8642,N_7753);
nor UO_1380 (O_1380,N_9721,N_8477);
nand UO_1381 (O_1381,N_8842,N_9227);
nor UO_1382 (O_1382,N_7951,N_9934);
and UO_1383 (O_1383,N_9155,N_8749);
xnor UO_1384 (O_1384,N_8467,N_8890);
nand UO_1385 (O_1385,N_9277,N_9241);
and UO_1386 (O_1386,N_9036,N_8522);
and UO_1387 (O_1387,N_9282,N_8041);
or UO_1388 (O_1388,N_8931,N_7866);
xnor UO_1389 (O_1389,N_8750,N_8159);
and UO_1390 (O_1390,N_8580,N_8100);
nand UO_1391 (O_1391,N_9065,N_8361);
or UO_1392 (O_1392,N_7654,N_9288);
nand UO_1393 (O_1393,N_7704,N_9748);
and UO_1394 (O_1394,N_7804,N_8530);
nand UO_1395 (O_1395,N_8063,N_9502);
or UO_1396 (O_1396,N_8274,N_8883);
or UO_1397 (O_1397,N_8694,N_9308);
and UO_1398 (O_1398,N_9027,N_9863);
nand UO_1399 (O_1399,N_9716,N_7588);
or UO_1400 (O_1400,N_7554,N_8464);
nor UO_1401 (O_1401,N_9171,N_9491);
nand UO_1402 (O_1402,N_8215,N_8989);
nor UO_1403 (O_1403,N_8104,N_9841);
nor UO_1404 (O_1404,N_9227,N_7696);
nand UO_1405 (O_1405,N_9306,N_9358);
or UO_1406 (O_1406,N_8359,N_9965);
and UO_1407 (O_1407,N_8884,N_8909);
or UO_1408 (O_1408,N_7797,N_7867);
and UO_1409 (O_1409,N_7679,N_9288);
and UO_1410 (O_1410,N_9390,N_7872);
or UO_1411 (O_1411,N_8083,N_9162);
or UO_1412 (O_1412,N_8759,N_8813);
or UO_1413 (O_1413,N_8470,N_7696);
nor UO_1414 (O_1414,N_9927,N_7762);
or UO_1415 (O_1415,N_8896,N_9951);
or UO_1416 (O_1416,N_8523,N_8927);
nand UO_1417 (O_1417,N_9890,N_7653);
xor UO_1418 (O_1418,N_7573,N_8012);
nor UO_1419 (O_1419,N_7972,N_9937);
and UO_1420 (O_1420,N_7948,N_9555);
and UO_1421 (O_1421,N_9064,N_8200);
nor UO_1422 (O_1422,N_8199,N_7817);
or UO_1423 (O_1423,N_8783,N_8582);
or UO_1424 (O_1424,N_8589,N_8163);
xnor UO_1425 (O_1425,N_9117,N_7856);
xor UO_1426 (O_1426,N_7975,N_8463);
nor UO_1427 (O_1427,N_7596,N_8911);
and UO_1428 (O_1428,N_9820,N_9524);
nor UO_1429 (O_1429,N_8689,N_7942);
nand UO_1430 (O_1430,N_7594,N_8676);
and UO_1431 (O_1431,N_9458,N_8337);
nand UO_1432 (O_1432,N_9598,N_8849);
or UO_1433 (O_1433,N_9895,N_8183);
nand UO_1434 (O_1434,N_8607,N_9321);
or UO_1435 (O_1435,N_8079,N_8491);
nor UO_1436 (O_1436,N_9311,N_9445);
or UO_1437 (O_1437,N_8857,N_9213);
nor UO_1438 (O_1438,N_9523,N_8131);
or UO_1439 (O_1439,N_8840,N_7556);
nor UO_1440 (O_1440,N_8053,N_9746);
nor UO_1441 (O_1441,N_9768,N_9501);
or UO_1442 (O_1442,N_9001,N_9451);
or UO_1443 (O_1443,N_7576,N_9670);
and UO_1444 (O_1444,N_9729,N_9740);
and UO_1445 (O_1445,N_8946,N_9350);
nand UO_1446 (O_1446,N_9858,N_9017);
and UO_1447 (O_1447,N_9877,N_8116);
xnor UO_1448 (O_1448,N_7511,N_7657);
nand UO_1449 (O_1449,N_8128,N_8878);
nor UO_1450 (O_1450,N_7968,N_8442);
nor UO_1451 (O_1451,N_8396,N_8932);
nor UO_1452 (O_1452,N_8925,N_9220);
and UO_1453 (O_1453,N_9836,N_7752);
xor UO_1454 (O_1454,N_9644,N_9022);
nand UO_1455 (O_1455,N_9238,N_8732);
nand UO_1456 (O_1456,N_8218,N_8462);
xnor UO_1457 (O_1457,N_8209,N_7871);
and UO_1458 (O_1458,N_9600,N_8676);
and UO_1459 (O_1459,N_7663,N_8678);
and UO_1460 (O_1460,N_9553,N_7982);
nand UO_1461 (O_1461,N_7752,N_7700);
nand UO_1462 (O_1462,N_8750,N_9510);
or UO_1463 (O_1463,N_8999,N_8237);
xnor UO_1464 (O_1464,N_7895,N_9288);
nand UO_1465 (O_1465,N_9978,N_8329);
nor UO_1466 (O_1466,N_8822,N_9115);
and UO_1467 (O_1467,N_8519,N_9329);
xor UO_1468 (O_1468,N_9047,N_9682);
nand UO_1469 (O_1469,N_8094,N_7898);
nor UO_1470 (O_1470,N_8841,N_8872);
xor UO_1471 (O_1471,N_9211,N_9808);
nand UO_1472 (O_1472,N_9820,N_9895);
or UO_1473 (O_1473,N_9302,N_8361);
nand UO_1474 (O_1474,N_9694,N_8287);
or UO_1475 (O_1475,N_7614,N_8203);
and UO_1476 (O_1476,N_9006,N_9131);
xnor UO_1477 (O_1477,N_9898,N_8344);
and UO_1478 (O_1478,N_8751,N_8893);
and UO_1479 (O_1479,N_9917,N_9124);
nor UO_1480 (O_1480,N_8362,N_9473);
xor UO_1481 (O_1481,N_9248,N_9935);
nand UO_1482 (O_1482,N_8255,N_7525);
and UO_1483 (O_1483,N_7867,N_8869);
nand UO_1484 (O_1484,N_9839,N_9740);
and UO_1485 (O_1485,N_8820,N_7732);
nand UO_1486 (O_1486,N_8707,N_9641);
and UO_1487 (O_1487,N_8310,N_8959);
or UO_1488 (O_1488,N_8056,N_7800);
nor UO_1489 (O_1489,N_8265,N_8986);
or UO_1490 (O_1490,N_9410,N_8091);
nand UO_1491 (O_1491,N_8680,N_8829);
nor UO_1492 (O_1492,N_9890,N_8441);
nand UO_1493 (O_1493,N_9281,N_9365);
or UO_1494 (O_1494,N_7583,N_8334);
or UO_1495 (O_1495,N_8874,N_9461);
nor UO_1496 (O_1496,N_8738,N_8250);
or UO_1497 (O_1497,N_8654,N_7793);
xor UO_1498 (O_1498,N_9913,N_7649);
nor UO_1499 (O_1499,N_8246,N_7674);
endmodule