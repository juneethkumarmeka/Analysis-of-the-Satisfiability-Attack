module basic_1000_10000_1500_5_levels_2xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_995,In_952);
or U1 (N_1,In_314,In_512);
or U2 (N_2,In_644,In_351);
and U3 (N_3,In_554,In_780);
and U4 (N_4,In_155,In_65);
nor U5 (N_5,In_169,In_982);
or U6 (N_6,In_781,In_165);
and U7 (N_7,In_366,In_503);
or U8 (N_8,In_413,In_343);
nand U9 (N_9,In_590,In_215);
or U10 (N_10,In_531,In_726);
nand U11 (N_11,In_346,In_153);
or U12 (N_12,In_546,In_792);
and U13 (N_13,In_632,In_885);
or U14 (N_14,In_800,In_776);
and U15 (N_15,In_206,In_504);
or U16 (N_16,In_331,In_812);
and U17 (N_17,In_87,In_52);
nor U18 (N_18,In_595,In_485);
or U19 (N_19,In_691,In_316);
or U20 (N_20,In_362,In_476);
nand U21 (N_21,In_954,In_439);
and U22 (N_22,In_647,In_152);
nand U23 (N_23,In_741,In_565);
or U24 (N_24,In_139,In_886);
xor U25 (N_25,In_245,In_402);
nand U26 (N_26,In_602,In_703);
xnor U27 (N_27,In_455,In_729);
and U28 (N_28,In_748,In_149);
nor U29 (N_29,In_851,In_274);
nor U30 (N_30,In_850,In_18);
nand U31 (N_31,In_306,In_289);
and U32 (N_32,In_57,In_174);
or U33 (N_33,In_650,In_712);
or U34 (N_34,In_103,In_100);
and U35 (N_35,In_624,In_154);
nor U36 (N_36,In_129,In_612);
nor U37 (N_37,In_763,In_633);
or U38 (N_38,In_478,In_387);
or U39 (N_39,In_965,In_251);
or U40 (N_40,In_482,In_81);
nand U41 (N_41,In_583,In_10);
and U42 (N_42,In_842,In_575);
nand U43 (N_43,In_496,In_921);
or U44 (N_44,In_643,In_560);
or U45 (N_45,In_588,In_769);
and U46 (N_46,In_446,In_819);
or U47 (N_47,In_460,In_194);
nand U48 (N_48,In_16,In_871);
and U49 (N_49,In_19,In_852);
and U50 (N_50,In_755,In_766);
nor U51 (N_51,In_41,In_203);
nand U52 (N_52,In_121,In_158);
nor U53 (N_53,In_22,In_487);
nor U54 (N_54,In_700,In_209);
nor U55 (N_55,In_530,In_931);
or U56 (N_56,In_281,In_96);
and U57 (N_57,In_617,In_344);
nand U58 (N_58,In_679,In_704);
or U59 (N_59,In_266,In_735);
nor U60 (N_60,In_687,In_436);
nand U61 (N_61,In_297,In_7);
or U62 (N_62,In_867,In_923);
nor U63 (N_63,In_414,In_90);
nand U64 (N_64,In_142,In_649);
and U65 (N_65,In_743,In_205);
nand U66 (N_66,In_53,In_359);
nand U67 (N_67,In_872,In_779);
and U68 (N_68,In_311,In_645);
and U69 (N_69,In_86,In_72);
nand U70 (N_70,In_901,In_141);
nor U71 (N_71,In_299,In_592);
nor U72 (N_72,In_146,In_345);
or U73 (N_73,In_138,In_528);
and U74 (N_74,In_929,In_773);
nand U75 (N_75,In_191,In_60);
or U76 (N_76,In_278,In_888);
nor U77 (N_77,In_811,In_290);
and U78 (N_78,In_899,In_127);
and U79 (N_79,In_616,In_124);
and U80 (N_80,In_390,In_581);
and U81 (N_81,In_144,In_211);
or U82 (N_82,In_606,In_688);
or U83 (N_83,In_986,In_109);
or U84 (N_84,In_935,In_39);
nand U85 (N_85,In_913,In_628);
nor U86 (N_86,In_705,In_309);
and U87 (N_87,In_574,In_557);
nand U88 (N_88,In_454,In_707);
nand U89 (N_89,In_128,In_475);
and U90 (N_90,In_586,In_608);
or U91 (N_91,In_302,In_938);
and U92 (N_92,In_429,In_552);
or U93 (N_93,In_962,In_568);
nand U94 (N_94,In_925,In_898);
nor U95 (N_95,In_843,In_930);
or U96 (N_96,In_917,In_132);
nor U97 (N_97,In_862,In_909);
or U98 (N_98,In_48,In_515);
nor U99 (N_99,In_201,In_682);
nor U100 (N_100,In_280,In_622);
nand U101 (N_101,In_942,In_808);
nand U102 (N_102,In_58,In_210);
nand U103 (N_103,In_196,In_880);
or U104 (N_104,In_564,In_105);
nor U105 (N_105,In_63,In_364);
and U106 (N_106,In_431,In_330);
xnor U107 (N_107,In_67,In_613);
nor U108 (N_108,In_791,In_988);
nand U109 (N_109,In_559,In_859);
or U110 (N_110,In_118,In_591);
or U111 (N_111,In_549,In_320);
or U112 (N_112,In_534,In_269);
nand U113 (N_113,In_114,In_864);
nor U114 (N_114,In_927,In_156);
or U115 (N_115,In_777,In_524);
or U116 (N_116,In_458,In_976);
nor U117 (N_117,In_884,In_656);
or U118 (N_118,In_248,In_569);
and U119 (N_119,In_835,In_971);
and U120 (N_120,In_652,In_604);
and U121 (N_121,In_268,In_657);
nor U122 (N_122,In_409,In_64);
or U123 (N_123,In_974,In_2);
and U124 (N_124,In_500,In_912);
nand U125 (N_125,In_881,In_379);
or U126 (N_126,In_464,In_618);
nand U127 (N_127,In_33,In_133);
or U128 (N_128,In_902,In_603);
nor U129 (N_129,In_360,In_893);
nand U130 (N_130,In_733,In_438);
nand U131 (N_131,In_312,In_221);
nor U132 (N_132,In_709,In_456);
or U133 (N_133,In_826,In_523);
nand U134 (N_134,In_265,In_228);
or U135 (N_135,In_80,In_508);
nor U136 (N_136,In_329,In_375);
or U137 (N_137,In_999,In_273);
nor U138 (N_138,In_240,In_372);
nand U139 (N_139,In_101,In_598);
and U140 (N_140,In_467,In_510);
and U141 (N_141,In_45,In_382);
or U142 (N_142,In_261,In_572);
or U143 (N_143,In_753,In_148);
and U144 (N_144,In_36,In_627);
nor U145 (N_145,In_257,In_846);
and U146 (N_146,In_6,In_896);
nand U147 (N_147,In_630,In_635);
and U148 (N_148,In_411,In_989);
nand U149 (N_149,In_365,In_834);
nand U150 (N_150,In_352,In_388);
or U151 (N_151,In_170,In_21);
and U152 (N_152,In_180,In_15);
and U153 (N_153,In_31,In_746);
nand U154 (N_154,In_533,In_50);
or U155 (N_155,In_936,In_181);
nor U156 (N_156,In_997,In_399);
nand U157 (N_157,In_803,In_767);
nor U158 (N_158,In_651,In_298);
and U159 (N_159,In_789,In_354);
nand U160 (N_160,In_810,In_192);
nand U161 (N_161,In_561,In_163);
nor U162 (N_162,In_878,In_293);
nand U163 (N_163,In_304,In_88);
nand U164 (N_164,In_111,In_120);
and U165 (N_165,In_959,In_906);
and U166 (N_166,In_793,In_224);
or U167 (N_167,In_469,In_232);
or U168 (N_168,In_914,In_162);
and U169 (N_169,In_507,In_951);
nor U170 (N_170,In_126,In_684);
nor U171 (N_171,In_958,In_573);
nor U172 (N_172,In_903,In_911);
and U173 (N_173,In_778,In_77);
nand U174 (N_174,In_668,In_840);
and U175 (N_175,In_380,In_782);
nand U176 (N_176,In_695,In_44);
and U177 (N_177,In_42,In_193);
nor U178 (N_178,In_747,In_806);
or U179 (N_179,In_59,In_607);
nor U180 (N_180,In_356,In_757);
nand U181 (N_181,In_736,In_368);
and U182 (N_182,In_593,In_374);
and U183 (N_183,In_673,In_236);
nor U184 (N_184,In_887,In_870);
or U185 (N_185,In_879,In_285);
and U186 (N_186,In_519,In_889);
nand U187 (N_187,In_212,In_488);
nor U188 (N_188,In_981,In_646);
nand U189 (N_189,In_355,In_30);
nand U190 (N_190,In_397,In_279);
and U191 (N_191,In_823,In_648);
and U192 (N_192,In_764,In_979);
nor U193 (N_193,In_226,In_238);
and U194 (N_194,In_953,In_214);
or U195 (N_195,In_417,In_816);
or U196 (N_196,In_875,In_449);
nand U197 (N_197,In_966,In_112);
and U198 (N_198,In_532,In_548);
nand U199 (N_199,In_396,In_415);
xnor U200 (N_200,In_809,In_805);
nand U201 (N_201,In_94,In_398);
or U202 (N_202,In_246,In_945);
nand U203 (N_203,In_336,In_734);
and U204 (N_204,In_738,In_333);
nor U205 (N_205,In_264,In_494);
and U206 (N_206,In_916,In_13);
nor U207 (N_207,In_724,In_623);
nand U208 (N_208,In_424,In_972);
nor U209 (N_209,In_699,In_970);
nor U210 (N_210,In_451,In_854);
xnor U211 (N_211,In_327,In_85);
and U212 (N_212,In_183,In_667);
nor U213 (N_213,In_401,In_949);
nand U214 (N_214,In_75,In_754);
and U215 (N_215,In_964,In_577);
and U216 (N_216,In_296,In_908);
nand U217 (N_217,In_73,In_242);
or U218 (N_218,In_253,In_479);
or U219 (N_219,In_828,In_615);
and U220 (N_220,In_115,In_877);
nor U221 (N_221,In_459,In_317);
nor U222 (N_222,In_340,In_218);
nor U223 (N_223,In_117,In_465);
and U224 (N_224,In_489,In_940);
or U225 (N_225,In_220,In_318);
or U226 (N_226,In_334,In_861);
xor U227 (N_227,In_762,In_0);
and U228 (N_228,In_693,In_701);
nand U229 (N_229,In_186,In_230);
and U230 (N_230,In_787,In_710);
nand U231 (N_231,In_654,In_660);
and U232 (N_232,In_737,In_659);
nand U233 (N_233,In_594,In_468);
or U234 (N_234,In_1,In_928);
and U235 (N_235,In_43,In_625);
nor U236 (N_236,In_509,In_807);
and U237 (N_237,In_957,In_676);
nor U238 (N_238,In_639,In_335);
and U239 (N_239,In_70,In_948);
and U240 (N_240,In_377,In_664);
or U241 (N_241,In_815,In_786);
nor U242 (N_242,In_794,In_521);
or U243 (N_243,In_994,In_444);
nand U244 (N_244,In_943,In_255);
and U245 (N_245,In_430,In_984);
nor U246 (N_246,In_99,In_410);
and U247 (N_247,In_185,In_801);
nor U248 (N_248,In_730,In_308);
nor U249 (N_249,In_599,In_977);
and U250 (N_250,In_140,In_821);
nand U251 (N_251,In_744,In_865);
and U252 (N_252,In_631,In_461);
nand U253 (N_253,In_547,In_428);
nor U254 (N_254,In_349,In_225);
or U255 (N_255,In_605,In_731);
and U256 (N_256,In_262,In_25);
nand U257 (N_257,In_391,In_27);
xor U258 (N_258,In_434,In_670);
nand U259 (N_259,In_157,In_207);
nand U260 (N_260,In_969,In_291);
nand U261 (N_261,In_924,In_204);
nand U262 (N_262,In_529,In_235);
nand U263 (N_263,In_34,In_381);
or U264 (N_264,In_250,In_24);
and U265 (N_265,In_714,In_991);
or U266 (N_266,In_395,In_389);
nor U267 (N_267,In_915,In_130);
and U268 (N_268,In_371,In_23);
or U269 (N_269,In_818,In_239);
nand U270 (N_270,In_946,In_102);
xor U271 (N_271,In_171,In_498);
and U272 (N_272,In_740,In_227);
and U273 (N_273,In_824,In_759);
nor U274 (N_274,In_677,In_956);
xnor U275 (N_275,In_722,In_200);
or U276 (N_276,In_907,In_166);
or U277 (N_277,In_696,In_527);
nand U278 (N_278,In_983,In_283);
and U279 (N_279,In_442,In_955);
nor U280 (N_280,In_135,In_987);
and U281 (N_281,In_28,In_985);
nor U282 (N_282,In_990,In_678);
nor U283 (N_283,In_520,In_725);
nand U284 (N_284,In_890,In_937);
and U285 (N_285,In_29,In_868);
nor U286 (N_286,In_944,In_502);
nand U287 (N_287,In_178,In_347);
xor U288 (N_288,In_544,In_324);
nor U289 (N_289,In_416,In_752);
nor U290 (N_290,In_536,In_258);
or U291 (N_291,In_638,In_721);
or U292 (N_292,In_55,In_11);
nand U293 (N_293,In_910,In_838);
and U294 (N_294,In_136,In_892);
nand U295 (N_295,In_483,In_975);
nand U296 (N_296,In_551,In_217);
nand U297 (N_297,In_939,In_686);
nor U298 (N_298,In_137,In_405);
nand U299 (N_299,In_400,In_849);
and U300 (N_300,In_611,In_471);
xor U301 (N_301,In_159,In_481);
nor U302 (N_302,In_751,In_827);
or U303 (N_303,In_62,In_681);
nor U304 (N_304,In_576,In_69);
or U305 (N_305,In_784,In_474);
nor U306 (N_306,In_869,In_276);
nand U307 (N_307,In_855,In_727);
nor U308 (N_308,In_950,In_272);
or U309 (N_309,In_435,In_768);
nand U310 (N_310,In_873,In_104);
nand U311 (N_311,In_589,In_83);
or U312 (N_312,In_516,In_300);
or U313 (N_313,In_295,In_814);
or U314 (N_314,In_216,In_145);
nor U315 (N_315,In_56,In_848);
and U316 (N_316,In_685,In_219);
and U317 (N_317,In_383,In_199);
and U318 (N_318,In_4,In_369);
and U319 (N_319,In_963,In_263);
nand U320 (N_320,In_202,In_406);
nand U321 (N_321,In_378,In_17);
nor U322 (N_322,In_143,In_629);
nor U323 (N_323,In_46,In_897);
nand U324 (N_324,In_506,In_614);
xnor U325 (N_325,In_175,In_698);
or U326 (N_326,In_817,In_342);
nor U327 (N_327,In_790,In_282);
or U328 (N_328,In_47,In_92);
nand U329 (N_329,In_79,In_732);
and U330 (N_330,In_425,In_426);
nor U331 (N_331,In_339,In_980);
and U332 (N_332,In_462,In_131);
nor U333 (N_333,In_244,In_905);
and U334 (N_334,In_486,In_961);
nand U335 (N_335,In_788,In_495);
nor U336 (N_336,In_452,In_770);
nand U337 (N_337,In_665,In_717);
nand U338 (N_338,In_641,In_470);
and U339 (N_339,In_233,In_177);
nor U340 (N_340,In_992,In_771);
nand U341 (N_341,In_582,In_5);
and U342 (N_342,In_445,In_553);
nor U343 (N_343,In_195,In_484);
or U344 (N_344,In_107,In_433);
or U345 (N_345,In_728,In_960);
nor U346 (N_346,In_243,In_539);
nor U347 (N_347,In_198,In_497);
nand U348 (N_348,In_421,In_491);
nor U349 (N_349,In_453,In_837);
xnor U350 (N_350,In_514,In_825);
and U351 (N_351,In_662,In_671);
or U352 (N_352,In_190,In_920);
nor U353 (N_353,In_739,In_348);
and U354 (N_354,In_719,In_550);
nor U355 (N_355,In_796,In_95);
xor U356 (N_356,In_847,In_213);
nand U357 (N_357,In_353,In_579);
or U358 (N_358,In_254,In_61);
or U359 (N_359,In_222,In_723);
or U360 (N_360,In_761,In_658);
or U361 (N_361,In_493,In_844);
nand U362 (N_362,In_229,In_501);
and U363 (N_363,In_918,In_363);
and U364 (N_364,In_967,In_772);
or U365 (N_365,In_116,In_669);
and U366 (N_366,In_742,In_537);
and U367 (N_367,In_125,In_160);
nand U368 (N_368,In_247,In_610);
and U369 (N_369,In_328,In_596);
nor U370 (N_370,In_288,In_386);
nand U371 (N_371,In_692,In_443);
or U372 (N_372,In_179,In_545);
and U373 (N_373,In_423,In_968);
or U374 (N_374,In_231,In_799);
and U375 (N_375,In_267,In_926);
nand U376 (N_376,In_525,In_934);
xnor U377 (N_377,In_511,In_35);
nand U378 (N_378,In_820,In_40);
and U379 (N_379,In_370,In_8);
and U380 (N_380,In_20,In_853);
nand U381 (N_381,In_490,In_275);
or U382 (N_382,In_492,In_978);
and U383 (N_383,In_601,In_188);
or U384 (N_384,In_91,In_715);
nand U385 (N_385,In_284,In_919);
nand U386 (N_386,In_566,In_341);
or U387 (N_387,In_313,In_271);
nor U388 (N_388,In_385,In_797);
nor U389 (N_389,In_798,In_173);
and U390 (N_390,In_350,In_82);
and U391 (N_391,In_774,In_882);
nand U392 (N_392,In_325,In_876);
nor U393 (N_393,In_836,In_640);
or U394 (N_394,In_113,In_642);
and U395 (N_395,In_277,In_357);
and U396 (N_396,In_249,In_89);
nand U397 (N_397,In_147,In_287);
and U398 (N_398,In_542,In_326);
or U399 (N_399,In_26,In_332);
or U400 (N_400,In_110,In_321);
and U401 (N_401,In_78,In_857);
nor U402 (N_402,In_440,In_480);
and U403 (N_403,In_252,In_338);
and U404 (N_404,In_432,In_562);
or U405 (N_405,In_637,In_653);
nand U406 (N_406,In_718,In_563);
nor U407 (N_407,In_535,In_322);
nand U408 (N_408,In_393,In_663);
or U409 (N_409,In_765,In_310);
or U410 (N_410,In_555,In_674);
or U411 (N_411,In_567,In_418);
nand U412 (N_412,In_839,In_74);
or U413 (N_413,In_473,In_151);
or U414 (N_414,In_833,In_499);
nand U415 (N_415,In_466,In_37);
xor U416 (N_416,In_237,In_150);
and U417 (N_417,In_197,In_900);
and U418 (N_418,In_384,In_973);
nand U419 (N_419,In_14,In_775);
and U420 (N_420,In_472,In_795);
nand U421 (N_421,In_32,In_634);
nor U422 (N_422,In_98,In_9);
nand U423 (N_423,In_51,In_675);
or U424 (N_424,In_578,In_690);
or U425 (N_425,In_571,In_441);
nor U426 (N_426,In_760,In_403);
and U427 (N_427,In_505,In_609);
and U428 (N_428,In_168,In_305);
nand U429 (N_429,In_758,In_860);
or U430 (N_430,In_477,In_404);
nor U431 (N_431,In_672,In_680);
nor U432 (N_432,In_711,In_785);
or U433 (N_433,In_376,In_38);
nand U434 (N_434,In_412,In_182);
nand U435 (N_435,In_941,In_526);
nor U436 (N_436,In_694,In_319);
nor U437 (N_437,In_303,In_292);
nor U438 (N_438,In_241,In_161);
nand U439 (N_439,In_831,In_891);
or U440 (N_440,In_3,In_518);
and U441 (N_441,In_301,In_904);
nand U442 (N_442,In_373,In_702);
and U443 (N_443,In_394,In_450);
nor U444 (N_444,In_619,In_866);
nand U445 (N_445,In_858,In_68);
and U446 (N_446,In_187,In_337);
or U447 (N_447,In_749,In_716);
nor U448 (N_448,In_66,In_448);
and U449 (N_449,In_367,In_260);
nand U450 (N_450,In_845,In_189);
nand U451 (N_451,In_713,In_184);
nand U452 (N_452,In_256,In_932);
or U453 (N_453,In_106,In_286);
xor U454 (N_454,In_108,In_708);
and U455 (N_455,In_558,In_122);
nor U456 (N_456,In_856,In_407);
or U457 (N_457,In_993,In_541);
xor U458 (N_458,In_683,In_830);
nand U459 (N_459,In_208,In_874);
nor U460 (N_460,In_538,In_176);
nor U461 (N_461,In_392,In_783);
and U462 (N_462,In_12,In_587);
or U463 (N_463,In_756,In_802);
xnor U464 (N_464,In_996,In_585);
xnor U465 (N_465,In_822,In_636);
or U466 (N_466,In_49,In_307);
and U467 (N_467,In_71,In_750);
nor U468 (N_468,In_164,In_570);
xor U469 (N_469,In_97,In_223);
or U470 (N_470,In_358,In_361);
nor U471 (N_471,In_895,In_259);
nand U472 (N_472,In_580,In_998);
or U473 (N_473,In_894,In_804);
xnor U474 (N_474,In_947,In_463);
and U475 (N_475,In_119,In_522);
nand U476 (N_476,In_841,In_123);
xnor U477 (N_477,In_620,In_621);
or U478 (N_478,In_167,In_666);
nand U479 (N_479,In_883,In_447);
nand U480 (N_480,In_720,In_427);
nand U481 (N_481,In_513,In_234);
xnor U482 (N_482,In_832,In_745);
nand U483 (N_483,In_134,In_93);
and U484 (N_484,In_270,In_597);
nand U485 (N_485,In_543,In_54);
or U486 (N_486,In_422,In_315);
and U487 (N_487,In_689,In_706);
nor U488 (N_488,In_294,In_323);
nor U489 (N_489,In_517,In_933);
nor U490 (N_490,In_437,In_829);
and U491 (N_491,In_600,In_813);
nor U492 (N_492,In_556,In_655);
xnor U493 (N_493,In_457,In_922);
and U494 (N_494,In_420,In_863);
nor U495 (N_495,In_76,In_661);
nand U496 (N_496,In_626,In_172);
and U497 (N_497,In_419,In_84);
and U498 (N_498,In_408,In_697);
or U499 (N_499,In_584,In_540);
xnor U500 (N_500,In_318,In_817);
nor U501 (N_501,In_963,In_200);
and U502 (N_502,In_137,In_877);
nand U503 (N_503,In_70,In_62);
nand U504 (N_504,In_285,In_860);
nand U505 (N_505,In_802,In_715);
nor U506 (N_506,In_568,In_257);
or U507 (N_507,In_978,In_471);
nand U508 (N_508,In_504,In_163);
and U509 (N_509,In_532,In_436);
nor U510 (N_510,In_574,In_318);
nor U511 (N_511,In_983,In_273);
nand U512 (N_512,In_618,In_445);
nor U513 (N_513,In_268,In_495);
or U514 (N_514,In_732,In_713);
or U515 (N_515,In_638,In_596);
and U516 (N_516,In_351,In_763);
and U517 (N_517,In_391,In_965);
nand U518 (N_518,In_175,In_926);
and U519 (N_519,In_114,In_91);
nor U520 (N_520,In_262,In_412);
nand U521 (N_521,In_544,In_428);
or U522 (N_522,In_259,In_592);
nand U523 (N_523,In_309,In_580);
or U524 (N_524,In_182,In_108);
and U525 (N_525,In_196,In_304);
nor U526 (N_526,In_355,In_285);
nand U527 (N_527,In_923,In_496);
or U528 (N_528,In_175,In_598);
nor U529 (N_529,In_963,In_326);
and U530 (N_530,In_44,In_368);
nor U531 (N_531,In_197,In_675);
nor U532 (N_532,In_974,In_149);
nand U533 (N_533,In_697,In_282);
nand U534 (N_534,In_70,In_99);
and U535 (N_535,In_508,In_598);
nor U536 (N_536,In_828,In_883);
nor U537 (N_537,In_111,In_880);
or U538 (N_538,In_364,In_767);
or U539 (N_539,In_355,In_259);
and U540 (N_540,In_120,In_794);
nor U541 (N_541,In_855,In_914);
or U542 (N_542,In_826,In_743);
nor U543 (N_543,In_7,In_138);
nand U544 (N_544,In_295,In_61);
nand U545 (N_545,In_127,In_693);
or U546 (N_546,In_151,In_518);
or U547 (N_547,In_669,In_149);
or U548 (N_548,In_682,In_834);
nand U549 (N_549,In_830,In_465);
nand U550 (N_550,In_997,In_436);
or U551 (N_551,In_890,In_515);
nor U552 (N_552,In_799,In_241);
nand U553 (N_553,In_930,In_774);
nand U554 (N_554,In_336,In_154);
nand U555 (N_555,In_888,In_244);
nor U556 (N_556,In_548,In_714);
nor U557 (N_557,In_813,In_798);
or U558 (N_558,In_482,In_394);
and U559 (N_559,In_781,In_345);
and U560 (N_560,In_84,In_680);
and U561 (N_561,In_140,In_559);
and U562 (N_562,In_83,In_494);
or U563 (N_563,In_601,In_900);
nand U564 (N_564,In_91,In_954);
and U565 (N_565,In_224,In_261);
and U566 (N_566,In_859,In_122);
or U567 (N_567,In_189,In_401);
nor U568 (N_568,In_917,In_75);
or U569 (N_569,In_654,In_239);
nand U570 (N_570,In_893,In_602);
nor U571 (N_571,In_872,In_878);
xnor U572 (N_572,In_202,In_312);
and U573 (N_573,In_430,In_402);
or U574 (N_574,In_709,In_312);
and U575 (N_575,In_856,In_699);
nor U576 (N_576,In_826,In_309);
nand U577 (N_577,In_124,In_732);
nor U578 (N_578,In_249,In_730);
nand U579 (N_579,In_895,In_757);
nor U580 (N_580,In_833,In_339);
and U581 (N_581,In_591,In_607);
nor U582 (N_582,In_749,In_901);
and U583 (N_583,In_950,In_852);
nor U584 (N_584,In_43,In_244);
nand U585 (N_585,In_414,In_563);
and U586 (N_586,In_104,In_599);
or U587 (N_587,In_608,In_227);
or U588 (N_588,In_553,In_959);
and U589 (N_589,In_283,In_847);
or U590 (N_590,In_757,In_369);
nor U591 (N_591,In_875,In_806);
nor U592 (N_592,In_461,In_974);
or U593 (N_593,In_182,In_173);
nand U594 (N_594,In_95,In_543);
nand U595 (N_595,In_494,In_173);
nand U596 (N_596,In_874,In_902);
or U597 (N_597,In_745,In_378);
nor U598 (N_598,In_804,In_257);
nand U599 (N_599,In_695,In_652);
nor U600 (N_600,In_62,In_235);
or U601 (N_601,In_394,In_337);
and U602 (N_602,In_366,In_239);
nand U603 (N_603,In_112,In_30);
and U604 (N_604,In_714,In_604);
or U605 (N_605,In_352,In_751);
and U606 (N_606,In_431,In_392);
and U607 (N_607,In_510,In_551);
or U608 (N_608,In_457,In_880);
and U609 (N_609,In_933,In_792);
and U610 (N_610,In_455,In_26);
or U611 (N_611,In_140,In_772);
and U612 (N_612,In_262,In_792);
or U613 (N_613,In_163,In_434);
nor U614 (N_614,In_952,In_546);
nor U615 (N_615,In_377,In_395);
nor U616 (N_616,In_92,In_42);
xnor U617 (N_617,In_433,In_19);
nand U618 (N_618,In_528,In_598);
nor U619 (N_619,In_296,In_126);
nor U620 (N_620,In_624,In_871);
nand U621 (N_621,In_454,In_703);
nand U622 (N_622,In_341,In_455);
or U623 (N_623,In_570,In_413);
and U624 (N_624,In_441,In_754);
nand U625 (N_625,In_987,In_823);
or U626 (N_626,In_115,In_865);
nor U627 (N_627,In_930,In_278);
nand U628 (N_628,In_893,In_190);
nand U629 (N_629,In_699,In_688);
nand U630 (N_630,In_441,In_445);
nor U631 (N_631,In_102,In_247);
and U632 (N_632,In_256,In_308);
or U633 (N_633,In_636,In_7);
nand U634 (N_634,In_808,In_997);
and U635 (N_635,In_604,In_159);
nor U636 (N_636,In_716,In_203);
nand U637 (N_637,In_990,In_822);
nand U638 (N_638,In_727,In_460);
xnor U639 (N_639,In_572,In_485);
and U640 (N_640,In_219,In_843);
nor U641 (N_641,In_212,In_948);
nor U642 (N_642,In_436,In_847);
nand U643 (N_643,In_713,In_61);
xnor U644 (N_644,In_854,In_827);
or U645 (N_645,In_458,In_456);
and U646 (N_646,In_590,In_905);
and U647 (N_647,In_486,In_350);
nand U648 (N_648,In_443,In_837);
nand U649 (N_649,In_235,In_415);
nor U650 (N_650,In_349,In_642);
or U651 (N_651,In_608,In_627);
nor U652 (N_652,In_737,In_832);
or U653 (N_653,In_894,In_72);
and U654 (N_654,In_718,In_311);
or U655 (N_655,In_439,In_678);
xnor U656 (N_656,In_201,In_551);
and U657 (N_657,In_467,In_523);
or U658 (N_658,In_476,In_136);
or U659 (N_659,In_862,In_234);
and U660 (N_660,In_427,In_713);
or U661 (N_661,In_392,In_308);
and U662 (N_662,In_642,In_105);
nor U663 (N_663,In_801,In_889);
xnor U664 (N_664,In_406,In_83);
nor U665 (N_665,In_397,In_92);
and U666 (N_666,In_451,In_69);
and U667 (N_667,In_680,In_400);
nand U668 (N_668,In_193,In_447);
nor U669 (N_669,In_913,In_709);
and U670 (N_670,In_701,In_715);
nand U671 (N_671,In_149,In_960);
or U672 (N_672,In_348,In_265);
or U673 (N_673,In_908,In_76);
xor U674 (N_674,In_635,In_920);
nor U675 (N_675,In_786,In_446);
or U676 (N_676,In_206,In_44);
nand U677 (N_677,In_559,In_545);
nor U678 (N_678,In_476,In_359);
and U679 (N_679,In_60,In_808);
nor U680 (N_680,In_13,In_585);
nor U681 (N_681,In_187,In_727);
and U682 (N_682,In_117,In_162);
nor U683 (N_683,In_115,In_836);
nand U684 (N_684,In_122,In_744);
nor U685 (N_685,In_625,In_644);
xnor U686 (N_686,In_498,In_250);
nor U687 (N_687,In_446,In_579);
nand U688 (N_688,In_421,In_341);
nor U689 (N_689,In_401,In_641);
nor U690 (N_690,In_113,In_920);
or U691 (N_691,In_622,In_629);
or U692 (N_692,In_343,In_777);
and U693 (N_693,In_141,In_466);
nand U694 (N_694,In_158,In_693);
or U695 (N_695,In_459,In_867);
nand U696 (N_696,In_581,In_498);
and U697 (N_697,In_284,In_465);
nor U698 (N_698,In_706,In_604);
nor U699 (N_699,In_449,In_638);
and U700 (N_700,In_695,In_99);
nand U701 (N_701,In_46,In_610);
nor U702 (N_702,In_198,In_503);
nor U703 (N_703,In_16,In_820);
nand U704 (N_704,In_464,In_505);
nand U705 (N_705,In_562,In_873);
and U706 (N_706,In_756,In_482);
or U707 (N_707,In_352,In_814);
and U708 (N_708,In_802,In_895);
nand U709 (N_709,In_89,In_849);
nand U710 (N_710,In_915,In_163);
and U711 (N_711,In_5,In_382);
nand U712 (N_712,In_980,In_847);
and U713 (N_713,In_498,In_169);
or U714 (N_714,In_839,In_345);
nor U715 (N_715,In_765,In_645);
nor U716 (N_716,In_394,In_449);
and U717 (N_717,In_68,In_115);
xor U718 (N_718,In_86,In_20);
and U719 (N_719,In_20,In_621);
or U720 (N_720,In_762,In_67);
nor U721 (N_721,In_366,In_865);
nand U722 (N_722,In_132,In_911);
nand U723 (N_723,In_417,In_782);
or U724 (N_724,In_533,In_459);
or U725 (N_725,In_154,In_47);
or U726 (N_726,In_935,In_144);
or U727 (N_727,In_121,In_772);
nand U728 (N_728,In_391,In_768);
nor U729 (N_729,In_835,In_207);
and U730 (N_730,In_879,In_682);
nor U731 (N_731,In_668,In_451);
nand U732 (N_732,In_764,In_601);
nor U733 (N_733,In_567,In_252);
or U734 (N_734,In_305,In_608);
and U735 (N_735,In_990,In_160);
and U736 (N_736,In_75,In_805);
or U737 (N_737,In_566,In_217);
and U738 (N_738,In_555,In_309);
or U739 (N_739,In_107,In_68);
nor U740 (N_740,In_791,In_765);
nor U741 (N_741,In_605,In_592);
and U742 (N_742,In_33,In_616);
nor U743 (N_743,In_706,In_894);
and U744 (N_744,In_275,In_421);
nor U745 (N_745,In_446,In_992);
and U746 (N_746,In_46,In_231);
nand U747 (N_747,In_17,In_521);
and U748 (N_748,In_229,In_607);
nand U749 (N_749,In_912,In_255);
nor U750 (N_750,In_162,In_756);
nor U751 (N_751,In_939,In_280);
or U752 (N_752,In_929,In_805);
nor U753 (N_753,In_163,In_785);
nand U754 (N_754,In_462,In_163);
or U755 (N_755,In_629,In_495);
nor U756 (N_756,In_145,In_128);
xnor U757 (N_757,In_536,In_8);
or U758 (N_758,In_744,In_582);
or U759 (N_759,In_117,In_407);
or U760 (N_760,In_326,In_649);
and U761 (N_761,In_537,In_367);
and U762 (N_762,In_212,In_684);
nand U763 (N_763,In_840,In_741);
nand U764 (N_764,In_223,In_773);
xor U765 (N_765,In_769,In_347);
nand U766 (N_766,In_280,In_122);
and U767 (N_767,In_819,In_260);
nor U768 (N_768,In_889,In_86);
nand U769 (N_769,In_813,In_632);
and U770 (N_770,In_62,In_638);
nor U771 (N_771,In_841,In_365);
or U772 (N_772,In_733,In_381);
nor U773 (N_773,In_0,In_832);
and U774 (N_774,In_992,In_191);
or U775 (N_775,In_991,In_925);
and U776 (N_776,In_298,In_765);
nor U777 (N_777,In_8,In_943);
nor U778 (N_778,In_433,In_207);
nor U779 (N_779,In_925,In_943);
nor U780 (N_780,In_942,In_95);
or U781 (N_781,In_666,In_19);
nand U782 (N_782,In_517,In_156);
nor U783 (N_783,In_472,In_830);
and U784 (N_784,In_564,In_171);
and U785 (N_785,In_56,In_186);
or U786 (N_786,In_490,In_798);
nand U787 (N_787,In_14,In_337);
or U788 (N_788,In_83,In_250);
xnor U789 (N_789,In_336,In_265);
and U790 (N_790,In_863,In_462);
and U791 (N_791,In_859,In_886);
or U792 (N_792,In_634,In_436);
xnor U793 (N_793,In_648,In_239);
and U794 (N_794,In_36,In_618);
and U795 (N_795,In_22,In_92);
nand U796 (N_796,In_683,In_862);
and U797 (N_797,In_714,In_92);
nand U798 (N_798,In_770,In_932);
nor U799 (N_799,In_414,In_63);
or U800 (N_800,In_916,In_700);
nor U801 (N_801,In_784,In_59);
and U802 (N_802,In_1,In_980);
nand U803 (N_803,In_609,In_754);
nand U804 (N_804,In_737,In_446);
nand U805 (N_805,In_45,In_692);
or U806 (N_806,In_724,In_640);
or U807 (N_807,In_580,In_11);
nand U808 (N_808,In_457,In_586);
or U809 (N_809,In_24,In_447);
nand U810 (N_810,In_842,In_250);
and U811 (N_811,In_696,In_410);
nand U812 (N_812,In_635,In_231);
and U813 (N_813,In_516,In_207);
and U814 (N_814,In_682,In_572);
and U815 (N_815,In_510,In_292);
nand U816 (N_816,In_88,In_489);
nor U817 (N_817,In_404,In_328);
nor U818 (N_818,In_816,In_46);
nand U819 (N_819,In_976,In_402);
nand U820 (N_820,In_276,In_449);
nor U821 (N_821,In_483,In_33);
nor U822 (N_822,In_356,In_675);
nand U823 (N_823,In_678,In_659);
nor U824 (N_824,In_877,In_682);
nand U825 (N_825,In_201,In_104);
nor U826 (N_826,In_307,In_542);
or U827 (N_827,In_515,In_223);
nor U828 (N_828,In_690,In_987);
and U829 (N_829,In_950,In_264);
or U830 (N_830,In_492,In_21);
nor U831 (N_831,In_22,In_999);
nand U832 (N_832,In_675,In_288);
or U833 (N_833,In_755,In_953);
or U834 (N_834,In_929,In_42);
nand U835 (N_835,In_172,In_671);
nand U836 (N_836,In_391,In_668);
nor U837 (N_837,In_419,In_768);
nor U838 (N_838,In_612,In_252);
or U839 (N_839,In_64,In_528);
nand U840 (N_840,In_45,In_326);
or U841 (N_841,In_51,In_135);
nor U842 (N_842,In_370,In_850);
nand U843 (N_843,In_923,In_491);
xnor U844 (N_844,In_275,In_373);
or U845 (N_845,In_201,In_68);
and U846 (N_846,In_443,In_610);
nand U847 (N_847,In_854,In_229);
and U848 (N_848,In_192,In_586);
and U849 (N_849,In_794,In_309);
nor U850 (N_850,In_710,In_815);
nand U851 (N_851,In_506,In_836);
and U852 (N_852,In_900,In_151);
or U853 (N_853,In_475,In_691);
nor U854 (N_854,In_179,In_363);
or U855 (N_855,In_762,In_243);
or U856 (N_856,In_634,In_150);
and U857 (N_857,In_181,In_714);
nand U858 (N_858,In_397,In_468);
nor U859 (N_859,In_389,In_251);
nand U860 (N_860,In_339,In_409);
nand U861 (N_861,In_761,In_934);
or U862 (N_862,In_257,In_328);
nand U863 (N_863,In_917,In_679);
and U864 (N_864,In_586,In_973);
or U865 (N_865,In_157,In_698);
and U866 (N_866,In_303,In_92);
or U867 (N_867,In_811,In_489);
and U868 (N_868,In_1,In_905);
nand U869 (N_869,In_514,In_802);
and U870 (N_870,In_769,In_372);
nand U871 (N_871,In_867,In_555);
nor U872 (N_872,In_319,In_948);
nor U873 (N_873,In_239,In_681);
nor U874 (N_874,In_22,In_533);
or U875 (N_875,In_471,In_712);
nand U876 (N_876,In_956,In_839);
and U877 (N_877,In_753,In_58);
nand U878 (N_878,In_513,In_546);
nor U879 (N_879,In_204,In_512);
or U880 (N_880,In_76,In_196);
or U881 (N_881,In_370,In_85);
nand U882 (N_882,In_23,In_937);
nand U883 (N_883,In_148,In_873);
nor U884 (N_884,In_483,In_75);
nor U885 (N_885,In_189,In_783);
nand U886 (N_886,In_661,In_107);
and U887 (N_887,In_254,In_65);
nor U888 (N_888,In_88,In_75);
and U889 (N_889,In_17,In_703);
and U890 (N_890,In_318,In_315);
nor U891 (N_891,In_75,In_944);
nor U892 (N_892,In_435,In_329);
and U893 (N_893,In_208,In_638);
and U894 (N_894,In_179,In_610);
nor U895 (N_895,In_757,In_692);
and U896 (N_896,In_384,In_829);
and U897 (N_897,In_526,In_29);
and U898 (N_898,In_620,In_407);
and U899 (N_899,In_436,In_321);
nand U900 (N_900,In_889,In_44);
nand U901 (N_901,In_825,In_684);
xor U902 (N_902,In_305,In_686);
nand U903 (N_903,In_50,In_345);
or U904 (N_904,In_532,In_557);
and U905 (N_905,In_547,In_759);
nand U906 (N_906,In_754,In_171);
or U907 (N_907,In_241,In_400);
and U908 (N_908,In_938,In_677);
and U909 (N_909,In_943,In_340);
nor U910 (N_910,In_379,In_529);
and U911 (N_911,In_32,In_107);
nand U912 (N_912,In_84,In_800);
nor U913 (N_913,In_405,In_35);
or U914 (N_914,In_500,In_804);
and U915 (N_915,In_286,In_909);
and U916 (N_916,In_469,In_754);
xor U917 (N_917,In_217,In_671);
and U918 (N_918,In_276,In_673);
nand U919 (N_919,In_869,In_92);
nor U920 (N_920,In_211,In_691);
nand U921 (N_921,In_955,In_819);
nand U922 (N_922,In_8,In_721);
and U923 (N_923,In_899,In_131);
nor U924 (N_924,In_200,In_202);
nor U925 (N_925,In_26,In_754);
nor U926 (N_926,In_440,In_197);
nor U927 (N_927,In_481,In_582);
and U928 (N_928,In_24,In_633);
and U929 (N_929,In_251,In_987);
nor U930 (N_930,In_252,In_883);
nor U931 (N_931,In_451,In_715);
and U932 (N_932,In_31,In_823);
or U933 (N_933,In_539,In_969);
and U934 (N_934,In_175,In_479);
and U935 (N_935,In_256,In_4);
nand U936 (N_936,In_96,In_622);
or U937 (N_937,In_681,In_405);
and U938 (N_938,In_552,In_689);
nor U939 (N_939,In_800,In_916);
nor U940 (N_940,In_662,In_376);
nor U941 (N_941,In_206,In_243);
nand U942 (N_942,In_35,In_426);
nand U943 (N_943,In_723,In_886);
nor U944 (N_944,In_969,In_309);
nand U945 (N_945,In_931,In_145);
and U946 (N_946,In_172,In_442);
nand U947 (N_947,In_923,In_156);
nor U948 (N_948,In_305,In_563);
nor U949 (N_949,In_125,In_984);
and U950 (N_950,In_753,In_512);
nor U951 (N_951,In_347,In_581);
or U952 (N_952,In_804,In_70);
nand U953 (N_953,In_606,In_938);
nand U954 (N_954,In_443,In_675);
nor U955 (N_955,In_515,In_380);
nor U956 (N_956,In_838,In_598);
or U957 (N_957,In_878,In_1);
nand U958 (N_958,In_556,In_829);
and U959 (N_959,In_788,In_797);
xor U960 (N_960,In_62,In_705);
and U961 (N_961,In_134,In_863);
nor U962 (N_962,In_800,In_992);
nand U963 (N_963,In_475,In_123);
nor U964 (N_964,In_521,In_559);
and U965 (N_965,In_888,In_520);
or U966 (N_966,In_806,In_13);
or U967 (N_967,In_11,In_722);
or U968 (N_968,In_934,In_943);
nand U969 (N_969,In_328,In_510);
nor U970 (N_970,In_114,In_361);
or U971 (N_971,In_924,In_835);
or U972 (N_972,In_659,In_492);
nand U973 (N_973,In_67,In_686);
or U974 (N_974,In_679,In_393);
or U975 (N_975,In_67,In_713);
or U976 (N_976,In_401,In_405);
xnor U977 (N_977,In_163,In_37);
and U978 (N_978,In_823,In_107);
and U979 (N_979,In_250,In_692);
or U980 (N_980,In_147,In_247);
and U981 (N_981,In_198,In_846);
nand U982 (N_982,In_177,In_657);
nor U983 (N_983,In_617,In_281);
and U984 (N_984,In_184,In_709);
or U985 (N_985,In_28,In_728);
and U986 (N_986,In_954,In_70);
nand U987 (N_987,In_413,In_323);
nor U988 (N_988,In_370,In_959);
nand U989 (N_989,In_737,In_356);
or U990 (N_990,In_53,In_852);
nor U991 (N_991,In_725,In_762);
nand U992 (N_992,In_166,In_609);
nand U993 (N_993,In_662,In_624);
or U994 (N_994,In_527,In_345);
or U995 (N_995,In_328,In_656);
or U996 (N_996,In_145,In_232);
xor U997 (N_997,In_629,In_488);
or U998 (N_998,In_733,In_330);
nor U999 (N_999,In_33,In_145);
nand U1000 (N_1000,In_537,In_532);
or U1001 (N_1001,In_326,In_944);
nor U1002 (N_1002,In_815,In_485);
and U1003 (N_1003,In_13,In_166);
and U1004 (N_1004,In_835,In_520);
or U1005 (N_1005,In_141,In_893);
or U1006 (N_1006,In_270,In_770);
nor U1007 (N_1007,In_926,In_941);
nand U1008 (N_1008,In_395,In_851);
xnor U1009 (N_1009,In_364,In_122);
nor U1010 (N_1010,In_892,In_864);
nor U1011 (N_1011,In_584,In_500);
and U1012 (N_1012,In_159,In_810);
and U1013 (N_1013,In_284,In_427);
nor U1014 (N_1014,In_396,In_52);
nand U1015 (N_1015,In_911,In_929);
nand U1016 (N_1016,In_299,In_103);
and U1017 (N_1017,In_74,In_726);
nor U1018 (N_1018,In_963,In_792);
and U1019 (N_1019,In_4,In_2);
nor U1020 (N_1020,In_525,In_517);
nand U1021 (N_1021,In_911,In_457);
and U1022 (N_1022,In_634,In_895);
or U1023 (N_1023,In_464,In_203);
nor U1024 (N_1024,In_582,In_305);
nand U1025 (N_1025,In_451,In_154);
or U1026 (N_1026,In_914,In_700);
or U1027 (N_1027,In_683,In_69);
nor U1028 (N_1028,In_664,In_825);
and U1029 (N_1029,In_759,In_433);
nand U1030 (N_1030,In_848,In_90);
nor U1031 (N_1031,In_978,In_385);
nor U1032 (N_1032,In_482,In_326);
nand U1033 (N_1033,In_436,In_153);
nand U1034 (N_1034,In_100,In_154);
and U1035 (N_1035,In_121,In_846);
and U1036 (N_1036,In_302,In_564);
or U1037 (N_1037,In_868,In_86);
or U1038 (N_1038,In_538,In_518);
xnor U1039 (N_1039,In_522,In_248);
nand U1040 (N_1040,In_715,In_302);
or U1041 (N_1041,In_301,In_292);
and U1042 (N_1042,In_592,In_890);
xor U1043 (N_1043,In_909,In_234);
nor U1044 (N_1044,In_895,In_362);
and U1045 (N_1045,In_789,In_157);
and U1046 (N_1046,In_475,In_479);
nand U1047 (N_1047,In_293,In_605);
or U1048 (N_1048,In_372,In_420);
or U1049 (N_1049,In_942,In_147);
nand U1050 (N_1050,In_526,In_586);
nor U1051 (N_1051,In_28,In_311);
nand U1052 (N_1052,In_719,In_389);
and U1053 (N_1053,In_152,In_702);
nor U1054 (N_1054,In_102,In_279);
xnor U1055 (N_1055,In_605,In_429);
nand U1056 (N_1056,In_798,In_500);
nand U1057 (N_1057,In_92,In_791);
or U1058 (N_1058,In_486,In_804);
or U1059 (N_1059,In_453,In_245);
and U1060 (N_1060,In_913,In_81);
nand U1061 (N_1061,In_327,In_241);
nand U1062 (N_1062,In_978,In_943);
or U1063 (N_1063,In_671,In_899);
nor U1064 (N_1064,In_724,In_184);
nor U1065 (N_1065,In_66,In_705);
nor U1066 (N_1066,In_171,In_713);
or U1067 (N_1067,In_531,In_202);
nand U1068 (N_1068,In_60,In_873);
or U1069 (N_1069,In_304,In_350);
nand U1070 (N_1070,In_556,In_863);
nor U1071 (N_1071,In_979,In_740);
nor U1072 (N_1072,In_634,In_545);
or U1073 (N_1073,In_230,In_529);
or U1074 (N_1074,In_562,In_138);
xnor U1075 (N_1075,In_537,In_807);
and U1076 (N_1076,In_479,In_815);
nand U1077 (N_1077,In_532,In_832);
nor U1078 (N_1078,In_882,In_221);
and U1079 (N_1079,In_190,In_480);
or U1080 (N_1080,In_698,In_721);
or U1081 (N_1081,In_445,In_337);
and U1082 (N_1082,In_113,In_964);
or U1083 (N_1083,In_533,In_649);
and U1084 (N_1084,In_791,In_38);
and U1085 (N_1085,In_830,In_422);
nor U1086 (N_1086,In_829,In_890);
or U1087 (N_1087,In_351,In_742);
nand U1088 (N_1088,In_825,In_734);
and U1089 (N_1089,In_397,In_420);
and U1090 (N_1090,In_676,In_827);
and U1091 (N_1091,In_119,In_515);
nor U1092 (N_1092,In_503,In_392);
or U1093 (N_1093,In_512,In_563);
or U1094 (N_1094,In_465,In_50);
or U1095 (N_1095,In_621,In_468);
and U1096 (N_1096,In_898,In_199);
or U1097 (N_1097,In_963,In_462);
and U1098 (N_1098,In_844,In_192);
or U1099 (N_1099,In_968,In_831);
nor U1100 (N_1100,In_251,In_254);
and U1101 (N_1101,In_424,In_273);
or U1102 (N_1102,In_84,In_794);
and U1103 (N_1103,In_546,In_135);
or U1104 (N_1104,In_466,In_650);
and U1105 (N_1105,In_233,In_142);
nand U1106 (N_1106,In_864,In_74);
nor U1107 (N_1107,In_431,In_489);
nand U1108 (N_1108,In_345,In_887);
or U1109 (N_1109,In_40,In_341);
nand U1110 (N_1110,In_896,In_262);
nand U1111 (N_1111,In_956,In_890);
and U1112 (N_1112,In_698,In_95);
or U1113 (N_1113,In_11,In_930);
and U1114 (N_1114,In_836,In_587);
nand U1115 (N_1115,In_69,In_982);
nor U1116 (N_1116,In_792,In_791);
and U1117 (N_1117,In_307,In_702);
nor U1118 (N_1118,In_302,In_495);
and U1119 (N_1119,In_129,In_564);
or U1120 (N_1120,In_201,In_202);
or U1121 (N_1121,In_341,In_974);
nor U1122 (N_1122,In_680,In_94);
or U1123 (N_1123,In_531,In_158);
nor U1124 (N_1124,In_995,In_198);
nand U1125 (N_1125,In_964,In_422);
nor U1126 (N_1126,In_448,In_45);
nor U1127 (N_1127,In_206,In_784);
nand U1128 (N_1128,In_677,In_319);
nor U1129 (N_1129,In_596,In_778);
and U1130 (N_1130,In_621,In_992);
nand U1131 (N_1131,In_482,In_959);
and U1132 (N_1132,In_119,In_576);
nand U1133 (N_1133,In_309,In_36);
or U1134 (N_1134,In_799,In_964);
or U1135 (N_1135,In_723,In_430);
nor U1136 (N_1136,In_850,In_92);
or U1137 (N_1137,In_215,In_200);
nand U1138 (N_1138,In_806,In_554);
nor U1139 (N_1139,In_409,In_488);
nand U1140 (N_1140,In_567,In_350);
and U1141 (N_1141,In_126,In_152);
nor U1142 (N_1142,In_891,In_116);
and U1143 (N_1143,In_106,In_873);
nor U1144 (N_1144,In_999,In_918);
nor U1145 (N_1145,In_946,In_281);
and U1146 (N_1146,In_474,In_334);
nand U1147 (N_1147,In_14,In_411);
nand U1148 (N_1148,In_821,In_966);
or U1149 (N_1149,In_616,In_513);
and U1150 (N_1150,In_445,In_827);
nand U1151 (N_1151,In_862,In_478);
nand U1152 (N_1152,In_155,In_599);
nand U1153 (N_1153,In_587,In_8);
and U1154 (N_1154,In_375,In_134);
nand U1155 (N_1155,In_960,In_956);
nor U1156 (N_1156,In_681,In_624);
and U1157 (N_1157,In_229,In_125);
nand U1158 (N_1158,In_373,In_767);
xor U1159 (N_1159,In_189,In_909);
nand U1160 (N_1160,In_452,In_1);
and U1161 (N_1161,In_415,In_513);
or U1162 (N_1162,In_69,In_142);
nor U1163 (N_1163,In_608,In_27);
nor U1164 (N_1164,In_253,In_682);
nor U1165 (N_1165,In_494,In_139);
nand U1166 (N_1166,In_797,In_191);
nand U1167 (N_1167,In_876,In_951);
or U1168 (N_1168,In_459,In_288);
and U1169 (N_1169,In_550,In_261);
nor U1170 (N_1170,In_560,In_207);
and U1171 (N_1171,In_520,In_161);
nor U1172 (N_1172,In_934,In_366);
and U1173 (N_1173,In_273,In_570);
nor U1174 (N_1174,In_123,In_144);
nor U1175 (N_1175,In_880,In_244);
xnor U1176 (N_1176,In_726,In_722);
or U1177 (N_1177,In_169,In_833);
nor U1178 (N_1178,In_635,In_930);
and U1179 (N_1179,In_590,In_709);
and U1180 (N_1180,In_430,In_695);
and U1181 (N_1181,In_294,In_192);
nor U1182 (N_1182,In_485,In_159);
or U1183 (N_1183,In_510,In_355);
and U1184 (N_1184,In_887,In_76);
nand U1185 (N_1185,In_33,In_971);
or U1186 (N_1186,In_281,In_791);
nor U1187 (N_1187,In_829,In_254);
nand U1188 (N_1188,In_379,In_97);
or U1189 (N_1189,In_580,In_50);
or U1190 (N_1190,In_417,In_647);
or U1191 (N_1191,In_850,In_33);
nor U1192 (N_1192,In_539,In_5);
xnor U1193 (N_1193,In_768,In_481);
nand U1194 (N_1194,In_535,In_18);
and U1195 (N_1195,In_322,In_682);
or U1196 (N_1196,In_631,In_370);
nor U1197 (N_1197,In_934,In_902);
and U1198 (N_1198,In_23,In_597);
xor U1199 (N_1199,In_318,In_234);
nand U1200 (N_1200,In_87,In_111);
nand U1201 (N_1201,In_153,In_301);
and U1202 (N_1202,In_677,In_273);
nand U1203 (N_1203,In_468,In_97);
nand U1204 (N_1204,In_419,In_828);
nor U1205 (N_1205,In_418,In_308);
or U1206 (N_1206,In_136,In_959);
or U1207 (N_1207,In_498,In_305);
and U1208 (N_1208,In_452,In_109);
nor U1209 (N_1209,In_398,In_430);
or U1210 (N_1210,In_646,In_74);
nand U1211 (N_1211,In_950,In_443);
or U1212 (N_1212,In_607,In_329);
nand U1213 (N_1213,In_793,In_369);
nor U1214 (N_1214,In_924,In_970);
or U1215 (N_1215,In_457,In_456);
or U1216 (N_1216,In_64,In_739);
nand U1217 (N_1217,In_867,In_9);
and U1218 (N_1218,In_370,In_1);
or U1219 (N_1219,In_965,In_990);
or U1220 (N_1220,In_671,In_351);
nor U1221 (N_1221,In_269,In_508);
or U1222 (N_1222,In_559,In_147);
nor U1223 (N_1223,In_142,In_309);
and U1224 (N_1224,In_224,In_316);
nand U1225 (N_1225,In_749,In_686);
nor U1226 (N_1226,In_943,In_1);
or U1227 (N_1227,In_250,In_503);
nand U1228 (N_1228,In_865,In_333);
or U1229 (N_1229,In_130,In_587);
or U1230 (N_1230,In_421,In_205);
and U1231 (N_1231,In_697,In_976);
and U1232 (N_1232,In_649,In_594);
nor U1233 (N_1233,In_891,In_820);
or U1234 (N_1234,In_582,In_48);
or U1235 (N_1235,In_99,In_106);
or U1236 (N_1236,In_537,In_255);
xor U1237 (N_1237,In_241,In_756);
or U1238 (N_1238,In_180,In_473);
nor U1239 (N_1239,In_521,In_594);
and U1240 (N_1240,In_458,In_656);
xor U1241 (N_1241,In_292,In_49);
or U1242 (N_1242,In_294,In_579);
nand U1243 (N_1243,In_355,In_815);
or U1244 (N_1244,In_850,In_369);
nor U1245 (N_1245,In_727,In_801);
or U1246 (N_1246,In_891,In_71);
nand U1247 (N_1247,In_635,In_147);
xnor U1248 (N_1248,In_56,In_475);
and U1249 (N_1249,In_528,In_127);
nand U1250 (N_1250,In_77,In_14);
nor U1251 (N_1251,In_281,In_704);
and U1252 (N_1252,In_592,In_604);
nor U1253 (N_1253,In_185,In_644);
and U1254 (N_1254,In_35,In_108);
nor U1255 (N_1255,In_317,In_848);
and U1256 (N_1256,In_939,In_937);
nand U1257 (N_1257,In_833,In_739);
and U1258 (N_1258,In_590,In_671);
nand U1259 (N_1259,In_723,In_25);
and U1260 (N_1260,In_613,In_225);
xnor U1261 (N_1261,In_758,In_50);
and U1262 (N_1262,In_75,In_926);
and U1263 (N_1263,In_343,In_140);
and U1264 (N_1264,In_324,In_673);
nand U1265 (N_1265,In_882,In_842);
nand U1266 (N_1266,In_121,In_292);
nand U1267 (N_1267,In_976,In_588);
or U1268 (N_1268,In_177,In_971);
nand U1269 (N_1269,In_596,In_39);
nand U1270 (N_1270,In_121,In_63);
nand U1271 (N_1271,In_533,In_290);
or U1272 (N_1272,In_21,In_679);
nand U1273 (N_1273,In_306,In_550);
nor U1274 (N_1274,In_956,In_629);
nor U1275 (N_1275,In_366,In_953);
and U1276 (N_1276,In_410,In_94);
nand U1277 (N_1277,In_785,In_792);
or U1278 (N_1278,In_351,In_855);
or U1279 (N_1279,In_641,In_809);
nor U1280 (N_1280,In_459,In_736);
and U1281 (N_1281,In_957,In_441);
nor U1282 (N_1282,In_417,In_74);
nor U1283 (N_1283,In_564,In_235);
and U1284 (N_1284,In_459,In_606);
nor U1285 (N_1285,In_868,In_555);
nand U1286 (N_1286,In_378,In_301);
and U1287 (N_1287,In_829,In_935);
or U1288 (N_1288,In_903,In_731);
nand U1289 (N_1289,In_231,In_702);
and U1290 (N_1290,In_161,In_503);
nor U1291 (N_1291,In_623,In_581);
and U1292 (N_1292,In_389,In_8);
and U1293 (N_1293,In_97,In_747);
nor U1294 (N_1294,In_386,In_264);
nor U1295 (N_1295,In_562,In_179);
nand U1296 (N_1296,In_557,In_934);
and U1297 (N_1297,In_762,In_327);
nand U1298 (N_1298,In_226,In_579);
nand U1299 (N_1299,In_414,In_281);
and U1300 (N_1300,In_287,In_293);
or U1301 (N_1301,In_505,In_858);
or U1302 (N_1302,In_236,In_204);
or U1303 (N_1303,In_425,In_594);
or U1304 (N_1304,In_59,In_158);
nor U1305 (N_1305,In_869,In_116);
nor U1306 (N_1306,In_475,In_421);
or U1307 (N_1307,In_270,In_233);
and U1308 (N_1308,In_274,In_684);
or U1309 (N_1309,In_460,In_170);
nor U1310 (N_1310,In_89,In_183);
and U1311 (N_1311,In_740,In_180);
nor U1312 (N_1312,In_14,In_444);
and U1313 (N_1313,In_971,In_331);
xnor U1314 (N_1314,In_252,In_641);
or U1315 (N_1315,In_598,In_422);
and U1316 (N_1316,In_227,In_752);
and U1317 (N_1317,In_186,In_898);
nor U1318 (N_1318,In_111,In_802);
and U1319 (N_1319,In_653,In_230);
and U1320 (N_1320,In_864,In_822);
nor U1321 (N_1321,In_73,In_809);
and U1322 (N_1322,In_632,In_552);
or U1323 (N_1323,In_317,In_415);
and U1324 (N_1324,In_644,In_689);
nand U1325 (N_1325,In_649,In_897);
and U1326 (N_1326,In_341,In_114);
and U1327 (N_1327,In_158,In_836);
nand U1328 (N_1328,In_118,In_200);
and U1329 (N_1329,In_545,In_814);
nand U1330 (N_1330,In_716,In_178);
and U1331 (N_1331,In_388,In_419);
or U1332 (N_1332,In_47,In_538);
and U1333 (N_1333,In_518,In_134);
nor U1334 (N_1334,In_342,In_229);
or U1335 (N_1335,In_328,In_72);
or U1336 (N_1336,In_91,In_975);
nor U1337 (N_1337,In_89,In_163);
nor U1338 (N_1338,In_538,In_252);
nand U1339 (N_1339,In_168,In_676);
and U1340 (N_1340,In_847,In_381);
nand U1341 (N_1341,In_772,In_392);
nand U1342 (N_1342,In_137,In_168);
and U1343 (N_1343,In_884,In_692);
xnor U1344 (N_1344,In_657,In_454);
nand U1345 (N_1345,In_160,In_263);
nor U1346 (N_1346,In_317,In_766);
or U1347 (N_1347,In_774,In_874);
nor U1348 (N_1348,In_887,In_958);
or U1349 (N_1349,In_310,In_449);
nor U1350 (N_1350,In_937,In_950);
or U1351 (N_1351,In_302,In_894);
nor U1352 (N_1352,In_702,In_926);
nor U1353 (N_1353,In_292,In_505);
nand U1354 (N_1354,In_740,In_724);
nand U1355 (N_1355,In_870,In_193);
nand U1356 (N_1356,In_1,In_683);
and U1357 (N_1357,In_848,In_405);
or U1358 (N_1358,In_997,In_867);
and U1359 (N_1359,In_454,In_957);
nor U1360 (N_1360,In_216,In_346);
nand U1361 (N_1361,In_451,In_561);
nor U1362 (N_1362,In_29,In_924);
nand U1363 (N_1363,In_490,In_363);
nand U1364 (N_1364,In_910,In_188);
and U1365 (N_1365,In_796,In_446);
or U1366 (N_1366,In_441,In_93);
or U1367 (N_1367,In_456,In_861);
and U1368 (N_1368,In_774,In_532);
or U1369 (N_1369,In_951,In_796);
nor U1370 (N_1370,In_196,In_981);
nor U1371 (N_1371,In_758,In_842);
or U1372 (N_1372,In_929,In_523);
and U1373 (N_1373,In_822,In_709);
and U1374 (N_1374,In_365,In_239);
xnor U1375 (N_1375,In_775,In_741);
nor U1376 (N_1376,In_926,In_123);
nor U1377 (N_1377,In_568,In_705);
or U1378 (N_1378,In_95,In_567);
and U1379 (N_1379,In_892,In_894);
and U1380 (N_1380,In_76,In_605);
and U1381 (N_1381,In_2,In_96);
nand U1382 (N_1382,In_213,In_746);
or U1383 (N_1383,In_973,In_773);
nand U1384 (N_1384,In_292,In_30);
and U1385 (N_1385,In_478,In_298);
nand U1386 (N_1386,In_461,In_96);
nor U1387 (N_1387,In_284,In_603);
or U1388 (N_1388,In_461,In_535);
nor U1389 (N_1389,In_966,In_888);
and U1390 (N_1390,In_925,In_658);
and U1391 (N_1391,In_791,In_274);
xnor U1392 (N_1392,In_96,In_91);
nand U1393 (N_1393,In_771,In_994);
nor U1394 (N_1394,In_105,In_75);
nand U1395 (N_1395,In_111,In_293);
nand U1396 (N_1396,In_470,In_968);
and U1397 (N_1397,In_578,In_327);
and U1398 (N_1398,In_75,In_583);
and U1399 (N_1399,In_204,In_601);
and U1400 (N_1400,In_365,In_49);
nand U1401 (N_1401,In_444,In_653);
xnor U1402 (N_1402,In_0,In_112);
and U1403 (N_1403,In_764,In_671);
and U1404 (N_1404,In_235,In_520);
nand U1405 (N_1405,In_997,In_637);
or U1406 (N_1406,In_262,In_592);
nand U1407 (N_1407,In_923,In_531);
or U1408 (N_1408,In_550,In_736);
nor U1409 (N_1409,In_956,In_324);
or U1410 (N_1410,In_797,In_669);
nand U1411 (N_1411,In_457,In_356);
and U1412 (N_1412,In_22,In_537);
nor U1413 (N_1413,In_830,In_667);
or U1414 (N_1414,In_453,In_807);
nand U1415 (N_1415,In_544,In_728);
nor U1416 (N_1416,In_924,In_115);
nand U1417 (N_1417,In_123,In_150);
nand U1418 (N_1418,In_770,In_978);
and U1419 (N_1419,In_647,In_886);
nand U1420 (N_1420,In_459,In_205);
and U1421 (N_1421,In_495,In_688);
nor U1422 (N_1422,In_531,In_777);
and U1423 (N_1423,In_326,In_411);
nand U1424 (N_1424,In_978,In_777);
or U1425 (N_1425,In_917,In_443);
or U1426 (N_1426,In_93,In_897);
nor U1427 (N_1427,In_238,In_680);
xor U1428 (N_1428,In_912,In_662);
nor U1429 (N_1429,In_822,In_226);
or U1430 (N_1430,In_118,In_764);
or U1431 (N_1431,In_340,In_833);
xor U1432 (N_1432,In_813,In_121);
and U1433 (N_1433,In_988,In_599);
nand U1434 (N_1434,In_467,In_343);
or U1435 (N_1435,In_187,In_768);
and U1436 (N_1436,In_179,In_810);
nor U1437 (N_1437,In_107,In_482);
nand U1438 (N_1438,In_260,In_796);
or U1439 (N_1439,In_214,In_663);
and U1440 (N_1440,In_485,In_996);
and U1441 (N_1441,In_319,In_137);
nor U1442 (N_1442,In_202,In_398);
nand U1443 (N_1443,In_355,In_575);
or U1444 (N_1444,In_172,In_446);
nand U1445 (N_1445,In_561,In_754);
nor U1446 (N_1446,In_661,In_144);
or U1447 (N_1447,In_754,In_786);
nand U1448 (N_1448,In_82,In_924);
and U1449 (N_1449,In_607,In_541);
nand U1450 (N_1450,In_805,In_263);
and U1451 (N_1451,In_639,In_894);
nand U1452 (N_1452,In_851,In_502);
nor U1453 (N_1453,In_879,In_613);
nand U1454 (N_1454,In_944,In_909);
nand U1455 (N_1455,In_701,In_232);
nor U1456 (N_1456,In_29,In_263);
and U1457 (N_1457,In_812,In_306);
nand U1458 (N_1458,In_530,In_357);
and U1459 (N_1459,In_644,In_959);
nor U1460 (N_1460,In_67,In_968);
or U1461 (N_1461,In_776,In_949);
nand U1462 (N_1462,In_149,In_783);
nor U1463 (N_1463,In_669,In_448);
nand U1464 (N_1464,In_198,In_183);
or U1465 (N_1465,In_490,In_18);
nor U1466 (N_1466,In_33,In_642);
or U1467 (N_1467,In_361,In_850);
nand U1468 (N_1468,In_875,In_400);
nor U1469 (N_1469,In_459,In_457);
nand U1470 (N_1470,In_483,In_575);
xnor U1471 (N_1471,In_888,In_449);
nor U1472 (N_1472,In_350,In_150);
nor U1473 (N_1473,In_353,In_89);
nor U1474 (N_1474,In_26,In_110);
nand U1475 (N_1475,In_248,In_673);
and U1476 (N_1476,In_411,In_436);
xnor U1477 (N_1477,In_957,In_945);
nand U1478 (N_1478,In_177,In_427);
nand U1479 (N_1479,In_85,In_962);
nand U1480 (N_1480,In_990,In_386);
nor U1481 (N_1481,In_786,In_761);
nor U1482 (N_1482,In_795,In_354);
nand U1483 (N_1483,In_327,In_55);
nor U1484 (N_1484,In_801,In_510);
or U1485 (N_1485,In_311,In_601);
nand U1486 (N_1486,In_812,In_827);
or U1487 (N_1487,In_926,In_399);
nand U1488 (N_1488,In_123,In_410);
nor U1489 (N_1489,In_262,In_37);
and U1490 (N_1490,In_690,In_719);
nand U1491 (N_1491,In_2,In_255);
nand U1492 (N_1492,In_908,In_349);
nor U1493 (N_1493,In_263,In_848);
nor U1494 (N_1494,In_580,In_685);
or U1495 (N_1495,In_682,In_100);
nor U1496 (N_1496,In_717,In_288);
nand U1497 (N_1497,In_998,In_44);
nand U1498 (N_1498,In_375,In_282);
nor U1499 (N_1499,In_111,In_291);
nand U1500 (N_1500,In_494,In_686);
nand U1501 (N_1501,In_312,In_83);
and U1502 (N_1502,In_950,In_845);
or U1503 (N_1503,In_44,In_757);
nand U1504 (N_1504,In_611,In_186);
and U1505 (N_1505,In_77,In_920);
nand U1506 (N_1506,In_144,In_365);
nor U1507 (N_1507,In_226,In_853);
nand U1508 (N_1508,In_429,In_617);
or U1509 (N_1509,In_878,In_753);
or U1510 (N_1510,In_403,In_926);
nand U1511 (N_1511,In_890,In_657);
nor U1512 (N_1512,In_601,In_93);
and U1513 (N_1513,In_1,In_43);
xor U1514 (N_1514,In_159,In_360);
and U1515 (N_1515,In_394,In_809);
nor U1516 (N_1516,In_73,In_357);
and U1517 (N_1517,In_180,In_80);
nor U1518 (N_1518,In_638,In_502);
or U1519 (N_1519,In_485,In_790);
xor U1520 (N_1520,In_237,In_502);
nand U1521 (N_1521,In_804,In_506);
and U1522 (N_1522,In_435,In_455);
nor U1523 (N_1523,In_101,In_729);
nor U1524 (N_1524,In_866,In_790);
nor U1525 (N_1525,In_414,In_628);
or U1526 (N_1526,In_505,In_146);
nor U1527 (N_1527,In_153,In_955);
nor U1528 (N_1528,In_582,In_58);
or U1529 (N_1529,In_274,In_60);
or U1530 (N_1530,In_316,In_839);
xor U1531 (N_1531,In_833,In_983);
or U1532 (N_1532,In_367,In_233);
or U1533 (N_1533,In_948,In_983);
nor U1534 (N_1534,In_875,In_574);
nand U1535 (N_1535,In_572,In_520);
and U1536 (N_1536,In_206,In_713);
nand U1537 (N_1537,In_555,In_676);
or U1538 (N_1538,In_971,In_746);
and U1539 (N_1539,In_192,In_316);
nand U1540 (N_1540,In_330,In_771);
and U1541 (N_1541,In_736,In_7);
nor U1542 (N_1542,In_448,In_627);
or U1543 (N_1543,In_922,In_224);
nand U1544 (N_1544,In_240,In_113);
or U1545 (N_1545,In_647,In_578);
or U1546 (N_1546,In_11,In_359);
or U1547 (N_1547,In_152,In_18);
nor U1548 (N_1548,In_528,In_806);
nor U1549 (N_1549,In_399,In_78);
nand U1550 (N_1550,In_422,In_140);
nor U1551 (N_1551,In_625,In_775);
or U1552 (N_1552,In_130,In_237);
nand U1553 (N_1553,In_770,In_118);
nor U1554 (N_1554,In_221,In_75);
nor U1555 (N_1555,In_544,In_700);
and U1556 (N_1556,In_501,In_85);
nand U1557 (N_1557,In_529,In_353);
and U1558 (N_1558,In_329,In_778);
nor U1559 (N_1559,In_454,In_367);
and U1560 (N_1560,In_510,In_157);
or U1561 (N_1561,In_610,In_595);
and U1562 (N_1562,In_63,In_802);
and U1563 (N_1563,In_514,In_715);
nor U1564 (N_1564,In_646,In_162);
and U1565 (N_1565,In_409,In_724);
nor U1566 (N_1566,In_580,In_348);
nor U1567 (N_1567,In_235,In_136);
and U1568 (N_1568,In_395,In_214);
and U1569 (N_1569,In_262,In_427);
or U1570 (N_1570,In_12,In_317);
nor U1571 (N_1571,In_662,In_53);
or U1572 (N_1572,In_417,In_721);
and U1573 (N_1573,In_52,In_910);
or U1574 (N_1574,In_612,In_535);
nand U1575 (N_1575,In_471,In_984);
nand U1576 (N_1576,In_950,In_598);
and U1577 (N_1577,In_41,In_471);
nand U1578 (N_1578,In_89,In_536);
nand U1579 (N_1579,In_173,In_811);
nand U1580 (N_1580,In_400,In_239);
nor U1581 (N_1581,In_21,In_408);
nor U1582 (N_1582,In_389,In_90);
xnor U1583 (N_1583,In_938,In_283);
or U1584 (N_1584,In_661,In_738);
and U1585 (N_1585,In_435,In_889);
and U1586 (N_1586,In_114,In_480);
or U1587 (N_1587,In_616,In_675);
nand U1588 (N_1588,In_529,In_561);
nor U1589 (N_1589,In_802,In_668);
or U1590 (N_1590,In_889,In_199);
and U1591 (N_1591,In_224,In_169);
and U1592 (N_1592,In_530,In_466);
or U1593 (N_1593,In_395,In_520);
and U1594 (N_1594,In_216,In_256);
nor U1595 (N_1595,In_382,In_567);
and U1596 (N_1596,In_298,In_732);
and U1597 (N_1597,In_116,In_614);
and U1598 (N_1598,In_389,In_42);
nor U1599 (N_1599,In_750,In_110);
nor U1600 (N_1600,In_249,In_888);
and U1601 (N_1601,In_986,In_918);
nor U1602 (N_1602,In_135,In_405);
and U1603 (N_1603,In_575,In_476);
nor U1604 (N_1604,In_768,In_396);
nor U1605 (N_1605,In_755,In_120);
or U1606 (N_1606,In_265,In_681);
nand U1607 (N_1607,In_300,In_470);
or U1608 (N_1608,In_696,In_320);
and U1609 (N_1609,In_342,In_850);
or U1610 (N_1610,In_533,In_514);
or U1611 (N_1611,In_988,In_288);
and U1612 (N_1612,In_216,In_161);
nand U1613 (N_1613,In_160,In_643);
nand U1614 (N_1614,In_0,In_686);
and U1615 (N_1615,In_124,In_159);
and U1616 (N_1616,In_894,In_838);
nor U1617 (N_1617,In_535,In_953);
nand U1618 (N_1618,In_227,In_945);
nor U1619 (N_1619,In_493,In_183);
and U1620 (N_1620,In_899,In_809);
nor U1621 (N_1621,In_66,In_472);
or U1622 (N_1622,In_166,In_359);
or U1623 (N_1623,In_177,In_307);
nand U1624 (N_1624,In_758,In_601);
or U1625 (N_1625,In_206,In_104);
and U1626 (N_1626,In_348,In_833);
or U1627 (N_1627,In_781,In_609);
xnor U1628 (N_1628,In_94,In_503);
nor U1629 (N_1629,In_247,In_869);
nand U1630 (N_1630,In_905,In_534);
nand U1631 (N_1631,In_909,In_192);
nand U1632 (N_1632,In_39,In_994);
or U1633 (N_1633,In_18,In_854);
or U1634 (N_1634,In_922,In_929);
nand U1635 (N_1635,In_766,In_70);
nor U1636 (N_1636,In_662,In_643);
nor U1637 (N_1637,In_589,In_22);
nand U1638 (N_1638,In_273,In_290);
nand U1639 (N_1639,In_627,In_385);
nor U1640 (N_1640,In_548,In_948);
nor U1641 (N_1641,In_962,In_143);
and U1642 (N_1642,In_388,In_411);
and U1643 (N_1643,In_441,In_406);
and U1644 (N_1644,In_56,In_556);
nand U1645 (N_1645,In_672,In_925);
and U1646 (N_1646,In_984,In_817);
or U1647 (N_1647,In_974,In_267);
or U1648 (N_1648,In_995,In_945);
nand U1649 (N_1649,In_85,In_592);
and U1650 (N_1650,In_863,In_886);
nand U1651 (N_1651,In_963,In_933);
or U1652 (N_1652,In_93,In_46);
nor U1653 (N_1653,In_188,In_913);
nor U1654 (N_1654,In_288,In_944);
nor U1655 (N_1655,In_819,In_608);
or U1656 (N_1656,In_15,In_736);
nor U1657 (N_1657,In_251,In_260);
or U1658 (N_1658,In_679,In_836);
or U1659 (N_1659,In_520,In_448);
or U1660 (N_1660,In_226,In_264);
or U1661 (N_1661,In_132,In_800);
or U1662 (N_1662,In_31,In_680);
nand U1663 (N_1663,In_685,In_222);
nor U1664 (N_1664,In_77,In_987);
nand U1665 (N_1665,In_354,In_449);
nor U1666 (N_1666,In_377,In_588);
and U1667 (N_1667,In_797,In_219);
and U1668 (N_1668,In_477,In_306);
or U1669 (N_1669,In_839,In_782);
and U1670 (N_1670,In_644,In_755);
and U1671 (N_1671,In_919,In_456);
nand U1672 (N_1672,In_747,In_599);
or U1673 (N_1673,In_416,In_485);
nand U1674 (N_1674,In_532,In_100);
nand U1675 (N_1675,In_425,In_209);
or U1676 (N_1676,In_179,In_206);
or U1677 (N_1677,In_452,In_724);
and U1678 (N_1678,In_153,In_408);
nor U1679 (N_1679,In_448,In_754);
or U1680 (N_1680,In_449,In_975);
and U1681 (N_1681,In_729,In_640);
nor U1682 (N_1682,In_858,In_565);
nand U1683 (N_1683,In_737,In_178);
nor U1684 (N_1684,In_374,In_3);
nand U1685 (N_1685,In_977,In_602);
or U1686 (N_1686,In_787,In_256);
xor U1687 (N_1687,In_115,In_867);
or U1688 (N_1688,In_636,In_683);
or U1689 (N_1689,In_334,In_991);
or U1690 (N_1690,In_30,In_780);
or U1691 (N_1691,In_52,In_143);
and U1692 (N_1692,In_852,In_938);
nor U1693 (N_1693,In_449,In_32);
and U1694 (N_1694,In_323,In_139);
nor U1695 (N_1695,In_114,In_107);
or U1696 (N_1696,In_822,In_608);
and U1697 (N_1697,In_690,In_425);
and U1698 (N_1698,In_227,In_526);
and U1699 (N_1699,In_133,In_489);
nor U1700 (N_1700,In_776,In_541);
nand U1701 (N_1701,In_169,In_999);
or U1702 (N_1702,In_433,In_558);
and U1703 (N_1703,In_329,In_400);
nor U1704 (N_1704,In_859,In_842);
nand U1705 (N_1705,In_40,In_885);
xnor U1706 (N_1706,In_30,In_56);
nand U1707 (N_1707,In_380,In_108);
and U1708 (N_1708,In_199,In_598);
and U1709 (N_1709,In_590,In_956);
or U1710 (N_1710,In_497,In_890);
and U1711 (N_1711,In_385,In_772);
or U1712 (N_1712,In_931,In_817);
nor U1713 (N_1713,In_652,In_395);
nor U1714 (N_1714,In_422,In_575);
nand U1715 (N_1715,In_618,In_682);
or U1716 (N_1716,In_967,In_902);
nand U1717 (N_1717,In_190,In_785);
or U1718 (N_1718,In_246,In_90);
nand U1719 (N_1719,In_742,In_370);
nand U1720 (N_1720,In_41,In_442);
nand U1721 (N_1721,In_28,In_544);
nor U1722 (N_1722,In_164,In_851);
nand U1723 (N_1723,In_663,In_384);
and U1724 (N_1724,In_833,In_22);
or U1725 (N_1725,In_57,In_106);
nor U1726 (N_1726,In_795,In_744);
or U1727 (N_1727,In_844,In_223);
or U1728 (N_1728,In_369,In_787);
or U1729 (N_1729,In_546,In_467);
and U1730 (N_1730,In_415,In_950);
nor U1731 (N_1731,In_617,In_764);
and U1732 (N_1732,In_624,In_397);
or U1733 (N_1733,In_500,In_935);
nand U1734 (N_1734,In_983,In_488);
nand U1735 (N_1735,In_284,In_827);
or U1736 (N_1736,In_629,In_244);
or U1737 (N_1737,In_807,In_570);
or U1738 (N_1738,In_2,In_580);
and U1739 (N_1739,In_769,In_962);
nand U1740 (N_1740,In_798,In_807);
and U1741 (N_1741,In_978,In_942);
nand U1742 (N_1742,In_462,In_181);
nor U1743 (N_1743,In_190,In_759);
nand U1744 (N_1744,In_72,In_347);
nand U1745 (N_1745,In_322,In_394);
nor U1746 (N_1746,In_949,In_67);
and U1747 (N_1747,In_798,In_137);
or U1748 (N_1748,In_440,In_986);
or U1749 (N_1749,In_730,In_891);
or U1750 (N_1750,In_346,In_554);
nand U1751 (N_1751,In_55,In_864);
nand U1752 (N_1752,In_561,In_297);
nand U1753 (N_1753,In_22,In_933);
nor U1754 (N_1754,In_221,In_131);
nor U1755 (N_1755,In_359,In_30);
or U1756 (N_1756,In_125,In_536);
and U1757 (N_1757,In_330,In_354);
nand U1758 (N_1758,In_995,In_978);
nor U1759 (N_1759,In_52,In_953);
and U1760 (N_1760,In_605,In_36);
nor U1761 (N_1761,In_940,In_730);
or U1762 (N_1762,In_69,In_377);
and U1763 (N_1763,In_585,In_419);
and U1764 (N_1764,In_212,In_517);
nor U1765 (N_1765,In_712,In_478);
xor U1766 (N_1766,In_858,In_889);
nor U1767 (N_1767,In_667,In_3);
or U1768 (N_1768,In_732,In_295);
nor U1769 (N_1769,In_878,In_911);
nor U1770 (N_1770,In_664,In_2);
nor U1771 (N_1771,In_190,In_725);
nor U1772 (N_1772,In_189,In_168);
nand U1773 (N_1773,In_467,In_885);
and U1774 (N_1774,In_211,In_312);
and U1775 (N_1775,In_931,In_900);
or U1776 (N_1776,In_159,In_572);
nor U1777 (N_1777,In_991,In_456);
nand U1778 (N_1778,In_666,In_356);
xnor U1779 (N_1779,In_675,In_900);
and U1780 (N_1780,In_385,In_277);
nand U1781 (N_1781,In_911,In_164);
or U1782 (N_1782,In_692,In_590);
and U1783 (N_1783,In_715,In_676);
or U1784 (N_1784,In_597,In_41);
nand U1785 (N_1785,In_411,In_36);
nand U1786 (N_1786,In_504,In_627);
and U1787 (N_1787,In_536,In_558);
nor U1788 (N_1788,In_660,In_193);
and U1789 (N_1789,In_116,In_576);
or U1790 (N_1790,In_756,In_674);
or U1791 (N_1791,In_160,In_487);
or U1792 (N_1792,In_793,In_428);
nand U1793 (N_1793,In_970,In_656);
and U1794 (N_1794,In_443,In_244);
and U1795 (N_1795,In_985,In_739);
or U1796 (N_1796,In_195,In_573);
and U1797 (N_1797,In_940,In_699);
xor U1798 (N_1798,In_971,In_72);
nand U1799 (N_1799,In_429,In_505);
and U1800 (N_1800,In_281,In_724);
or U1801 (N_1801,In_131,In_241);
nand U1802 (N_1802,In_364,In_232);
nor U1803 (N_1803,In_237,In_341);
and U1804 (N_1804,In_21,In_205);
and U1805 (N_1805,In_378,In_38);
nor U1806 (N_1806,In_726,In_374);
nor U1807 (N_1807,In_731,In_539);
nor U1808 (N_1808,In_100,In_131);
nor U1809 (N_1809,In_166,In_567);
and U1810 (N_1810,In_732,In_683);
nand U1811 (N_1811,In_480,In_359);
xnor U1812 (N_1812,In_853,In_168);
nand U1813 (N_1813,In_816,In_917);
and U1814 (N_1814,In_711,In_452);
nand U1815 (N_1815,In_265,In_437);
or U1816 (N_1816,In_988,In_575);
nand U1817 (N_1817,In_12,In_310);
and U1818 (N_1818,In_591,In_299);
nand U1819 (N_1819,In_644,In_55);
or U1820 (N_1820,In_910,In_189);
or U1821 (N_1821,In_16,In_831);
and U1822 (N_1822,In_543,In_129);
nand U1823 (N_1823,In_965,In_83);
nor U1824 (N_1824,In_968,In_111);
and U1825 (N_1825,In_947,In_327);
nor U1826 (N_1826,In_996,In_818);
or U1827 (N_1827,In_504,In_448);
nor U1828 (N_1828,In_337,In_855);
and U1829 (N_1829,In_113,In_860);
or U1830 (N_1830,In_64,In_456);
and U1831 (N_1831,In_52,In_261);
nor U1832 (N_1832,In_332,In_547);
nor U1833 (N_1833,In_978,In_228);
or U1834 (N_1834,In_129,In_317);
nor U1835 (N_1835,In_151,In_676);
xnor U1836 (N_1836,In_834,In_976);
or U1837 (N_1837,In_862,In_167);
xor U1838 (N_1838,In_753,In_557);
and U1839 (N_1839,In_718,In_929);
nor U1840 (N_1840,In_391,In_226);
nor U1841 (N_1841,In_532,In_282);
and U1842 (N_1842,In_392,In_912);
nor U1843 (N_1843,In_686,In_383);
nor U1844 (N_1844,In_769,In_548);
and U1845 (N_1845,In_203,In_76);
nor U1846 (N_1846,In_318,In_250);
and U1847 (N_1847,In_958,In_580);
nor U1848 (N_1848,In_537,In_102);
xnor U1849 (N_1849,In_318,In_712);
nand U1850 (N_1850,In_352,In_607);
nand U1851 (N_1851,In_7,In_855);
nand U1852 (N_1852,In_613,In_282);
or U1853 (N_1853,In_250,In_376);
nand U1854 (N_1854,In_630,In_911);
and U1855 (N_1855,In_448,In_235);
or U1856 (N_1856,In_957,In_886);
nand U1857 (N_1857,In_695,In_442);
or U1858 (N_1858,In_838,In_458);
nand U1859 (N_1859,In_177,In_997);
or U1860 (N_1860,In_8,In_435);
nand U1861 (N_1861,In_609,In_654);
or U1862 (N_1862,In_911,In_739);
nor U1863 (N_1863,In_261,In_930);
nor U1864 (N_1864,In_442,In_750);
or U1865 (N_1865,In_696,In_138);
and U1866 (N_1866,In_841,In_149);
nand U1867 (N_1867,In_804,In_887);
and U1868 (N_1868,In_410,In_672);
and U1869 (N_1869,In_481,In_774);
and U1870 (N_1870,In_407,In_806);
and U1871 (N_1871,In_269,In_348);
nor U1872 (N_1872,In_621,In_605);
nand U1873 (N_1873,In_189,In_558);
or U1874 (N_1874,In_952,In_59);
or U1875 (N_1875,In_986,In_795);
nand U1876 (N_1876,In_967,In_373);
or U1877 (N_1877,In_848,In_883);
nand U1878 (N_1878,In_38,In_807);
and U1879 (N_1879,In_236,In_844);
or U1880 (N_1880,In_300,In_592);
or U1881 (N_1881,In_196,In_796);
and U1882 (N_1882,In_444,In_837);
nand U1883 (N_1883,In_9,In_11);
or U1884 (N_1884,In_6,In_972);
nor U1885 (N_1885,In_561,In_797);
and U1886 (N_1886,In_68,In_204);
nor U1887 (N_1887,In_861,In_298);
and U1888 (N_1888,In_294,In_888);
nor U1889 (N_1889,In_411,In_13);
xor U1890 (N_1890,In_355,In_296);
nor U1891 (N_1891,In_272,In_419);
nand U1892 (N_1892,In_426,In_533);
or U1893 (N_1893,In_40,In_782);
nand U1894 (N_1894,In_198,In_717);
xor U1895 (N_1895,In_107,In_801);
nor U1896 (N_1896,In_101,In_825);
or U1897 (N_1897,In_510,In_613);
xnor U1898 (N_1898,In_49,In_551);
or U1899 (N_1899,In_635,In_887);
nand U1900 (N_1900,In_124,In_243);
nor U1901 (N_1901,In_835,In_353);
nand U1902 (N_1902,In_86,In_385);
nor U1903 (N_1903,In_603,In_287);
and U1904 (N_1904,In_801,In_482);
nor U1905 (N_1905,In_781,In_569);
nand U1906 (N_1906,In_862,In_406);
nand U1907 (N_1907,In_261,In_289);
and U1908 (N_1908,In_204,In_607);
and U1909 (N_1909,In_525,In_406);
and U1910 (N_1910,In_429,In_5);
nand U1911 (N_1911,In_544,In_349);
and U1912 (N_1912,In_804,In_96);
nor U1913 (N_1913,In_314,In_628);
nand U1914 (N_1914,In_639,In_462);
and U1915 (N_1915,In_932,In_246);
nand U1916 (N_1916,In_726,In_632);
nand U1917 (N_1917,In_273,In_110);
nand U1918 (N_1918,In_422,In_665);
or U1919 (N_1919,In_827,In_316);
nand U1920 (N_1920,In_329,In_841);
or U1921 (N_1921,In_205,In_563);
nand U1922 (N_1922,In_535,In_339);
nor U1923 (N_1923,In_815,In_478);
nor U1924 (N_1924,In_300,In_605);
or U1925 (N_1925,In_270,In_999);
nor U1926 (N_1926,In_749,In_352);
and U1927 (N_1927,In_649,In_452);
or U1928 (N_1928,In_511,In_985);
and U1929 (N_1929,In_528,In_596);
nand U1930 (N_1930,In_827,In_578);
xnor U1931 (N_1931,In_195,In_492);
and U1932 (N_1932,In_207,In_736);
and U1933 (N_1933,In_653,In_601);
nand U1934 (N_1934,In_700,In_234);
and U1935 (N_1935,In_964,In_723);
nor U1936 (N_1936,In_758,In_365);
nand U1937 (N_1937,In_973,In_353);
nor U1938 (N_1938,In_948,In_83);
nand U1939 (N_1939,In_20,In_296);
nand U1940 (N_1940,In_973,In_481);
nor U1941 (N_1941,In_552,In_288);
nor U1942 (N_1942,In_450,In_610);
or U1943 (N_1943,In_35,In_997);
nand U1944 (N_1944,In_503,In_889);
and U1945 (N_1945,In_985,In_109);
and U1946 (N_1946,In_809,In_646);
nor U1947 (N_1947,In_252,In_361);
or U1948 (N_1948,In_173,In_864);
nand U1949 (N_1949,In_998,In_750);
nor U1950 (N_1950,In_518,In_493);
nand U1951 (N_1951,In_521,In_28);
and U1952 (N_1952,In_242,In_199);
nand U1953 (N_1953,In_287,In_481);
nand U1954 (N_1954,In_625,In_685);
or U1955 (N_1955,In_333,In_444);
nand U1956 (N_1956,In_177,In_205);
nand U1957 (N_1957,In_598,In_602);
xnor U1958 (N_1958,In_285,In_600);
and U1959 (N_1959,In_733,In_209);
and U1960 (N_1960,In_545,In_922);
and U1961 (N_1961,In_285,In_815);
xnor U1962 (N_1962,In_791,In_420);
or U1963 (N_1963,In_991,In_734);
or U1964 (N_1964,In_565,In_826);
nor U1965 (N_1965,In_762,In_482);
nand U1966 (N_1966,In_280,In_634);
or U1967 (N_1967,In_687,In_742);
and U1968 (N_1968,In_330,In_695);
nand U1969 (N_1969,In_535,In_560);
nor U1970 (N_1970,In_64,In_941);
nand U1971 (N_1971,In_553,In_254);
nor U1972 (N_1972,In_876,In_659);
and U1973 (N_1973,In_129,In_433);
nor U1974 (N_1974,In_34,In_788);
or U1975 (N_1975,In_61,In_460);
and U1976 (N_1976,In_339,In_842);
nor U1977 (N_1977,In_479,In_691);
and U1978 (N_1978,In_584,In_51);
and U1979 (N_1979,In_788,In_505);
nor U1980 (N_1980,In_361,In_113);
or U1981 (N_1981,In_433,In_376);
and U1982 (N_1982,In_662,In_362);
and U1983 (N_1983,In_84,In_183);
xor U1984 (N_1984,In_764,In_358);
and U1985 (N_1985,In_391,In_880);
xnor U1986 (N_1986,In_965,In_53);
nor U1987 (N_1987,In_340,In_543);
nand U1988 (N_1988,In_212,In_692);
nor U1989 (N_1989,In_73,In_230);
nor U1990 (N_1990,In_740,In_818);
nor U1991 (N_1991,In_808,In_585);
or U1992 (N_1992,In_748,In_432);
or U1993 (N_1993,In_143,In_175);
nor U1994 (N_1994,In_894,In_472);
nand U1995 (N_1995,In_652,In_157);
nor U1996 (N_1996,In_158,In_780);
and U1997 (N_1997,In_976,In_865);
nand U1998 (N_1998,In_380,In_208);
and U1999 (N_1999,In_509,In_657);
or U2000 (N_2000,N_1253,N_1480);
or U2001 (N_2001,N_131,N_2);
and U2002 (N_2002,N_1319,N_505);
and U2003 (N_2003,N_1608,N_1040);
and U2004 (N_2004,N_1476,N_1672);
or U2005 (N_2005,N_1020,N_1396);
and U2006 (N_2006,N_1953,N_1428);
nand U2007 (N_2007,N_313,N_1970);
or U2008 (N_2008,N_1891,N_916);
nor U2009 (N_2009,N_253,N_632);
or U2010 (N_2010,N_67,N_172);
and U2011 (N_2011,N_878,N_1645);
nor U2012 (N_2012,N_1489,N_165);
and U2013 (N_2013,N_1644,N_19);
and U2014 (N_2014,N_1575,N_107);
or U2015 (N_2015,N_1071,N_514);
nor U2016 (N_2016,N_6,N_1643);
nor U2017 (N_2017,N_1900,N_877);
and U2018 (N_2018,N_963,N_1877);
and U2019 (N_2019,N_1101,N_1393);
nor U2020 (N_2020,N_1895,N_1652);
and U2021 (N_2021,N_731,N_1191);
and U2022 (N_2022,N_894,N_89);
or U2023 (N_2023,N_694,N_1036);
or U2024 (N_2024,N_1421,N_1367);
xnor U2025 (N_2025,N_570,N_1340);
or U2026 (N_2026,N_1297,N_511);
and U2027 (N_2027,N_1347,N_194);
nor U2028 (N_2028,N_1038,N_515);
nor U2029 (N_2029,N_1507,N_973);
nand U2030 (N_2030,N_1424,N_1129);
nand U2031 (N_2031,N_1680,N_723);
and U2032 (N_2032,N_1632,N_1143);
nand U2033 (N_2033,N_1812,N_1250);
and U2034 (N_2034,N_1899,N_798);
or U2035 (N_2035,N_1230,N_162);
and U2036 (N_2036,N_1994,N_1093);
nor U2037 (N_2037,N_222,N_292);
and U2038 (N_2038,N_1099,N_1752);
nand U2039 (N_2039,N_1098,N_0);
nor U2040 (N_2040,N_1602,N_249);
or U2041 (N_2041,N_1966,N_308);
nand U2042 (N_2042,N_1948,N_937);
or U2043 (N_2043,N_1998,N_1554);
nor U2044 (N_2044,N_1302,N_845);
nor U2045 (N_2045,N_1350,N_491);
nor U2046 (N_2046,N_522,N_1579);
nand U2047 (N_2047,N_1238,N_1282);
nor U2048 (N_2048,N_881,N_14);
or U2049 (N_2049,N_1638,N_527);
and U2050 (N_2050,N_1373,N_1597);
and U2051 (N_2051,N_1068,N_1648);
nor U2052 (N_2052,N_525,N_133);
or U2053 (N_2053,N_214,N_1235);
nor U2054 (N_2054,N_535,N_1357);
or U2055 (N_2055,N_1097,N_584);
or U2056 (N_2056,N_1770,N_608);
or U2057 (N_2057,N_1805,N_68);
nor U2058 (N_2058,N_1195,N_585);
nand U2059 (N_2059,N_1843,N_1668);
xor U2060 (N_2060,N_1288,N_628);
nand U2061 (N_2061,N_1066,N_352);
or U2062 (N_2062,N_1688,N_267);
or U2063 (N_2063,N_1317,N_1385);
and U2064 (N_2064,N_640,N_157);
xor U2065 (N_2065,N_235,N_960);
and U2066 (N_2066,N_71,N_1291);
nand U2067 (N_2067,N_8,N_1580);
nor U2068 (N_2068,N_775,N_695);
or U2069 (N_2069,N_1646,N_1723);
and U2070 (N_2070,N_1403,N_237);
nand U2071 (N_2071,N_247,N_243);
and U2072 (N_2072,N_650,N_1362);
or U2073 (N_2073,N_1369,N_793);
and U2074 (N_2074,N_1087,N_1278);
and U2075 (N_2075,N_61,N_73);
nand U2076 (N_2076,N_1592,N_431);
and U2077 (N_2077,N_552,N_1758);
nand U2078 (N_2078,N_251,N_1492);
or U2079 (N_2079,N_241,N_818);
or U2080 (N_2080,N_476,N_1659);
nor U2081 (N_2081,N_633,N_423);
nand U2082 (N_2082,N_875,N_1841);
nand U2083 (N_2083,N_899,N_1354);
nor U2084 (N_2084,N_1786,N_850);
or U2085 (N_2085,N_1784,N_849);
nand U2086 (N_2086,N_626,N_897);
nand U2087 (N_2087,N_123,N_1574);
or U2088 (N_2088,N_1446,N_1635);
nor U2089 (N_2089,N_1207,N_1154);
nor U2090 (N_2090,N_929,N_1828);
nor U2091 (N_2091,N_977,N_1193);
and U2092 (N_2092,N_78,N_983);
or U2093 (N_2093,N_579,N_817);
or U2094 (N_2094,N_443,N_786);
or U2095 (N_2095,N_1616,N_3);
and U2096 (N_2096,N_299,N_912);
or U2097 (N_2097,N_190,N_1307);
or U2098 (N_2098,N_1477,N_1522);
nand U2099 (N_2099,N_1830,N_1494);
nand U2100 (N_2100,N_1995,N_1621);
and U2101 (N_2101,N_662,N_872);
or U2102 (N_2102,N_1219,N_35);
nand U2103 (N_2103,N_160,N_90);
or U2104 (N_2104,N_368,N_781);
and U2105 (N_2105,N_905,N_199);
or U2106 (N_2106,N_23,N_571);
and U2107 (N_2107,N_398,N_36);
xnor U2108 (N_2108,N_480,N_1342);
or U2109 (N_2109,N_997,N_1807);
or U2110 (N_2110,N_1562,N_1206);
and U2111 (N_2111,N_1790,N_170);
nor U2112 (N_2112,N_291,N_1440);
nand U2113 (N_2113,N_1439,N_772);
or U2114 (N_2114,N_210,N_27);
nor U2115 (N_2115,N_196,N_10);
and U2116 (N_2116,N_16,N_1400);
nand U2117 (N_2117,N_147,N_389);
or U2118 (N_2118,N_599,N_919);
or U2119 (N_2119,N_754,N_1556);
and U2120 (N_2120,N_490,N_699);
or U2121 (N_2121,N_751,N_322);
nor U2122 (N_2122,N_787,N_114);
nor U2123 (N_2123,N_1280,N_1115);
nor U2124 (N_2124,N_1388,N_1510);
nand U2125 (N_2125,N_171,N_1054);
nand U2126 (N_2126,N_670,N_1955);
and U2127 (N_2127,N_17,N_1922);
or U2128 (N_2128,N_207,N_1775);
and U2129 (N_2129,N_1442,N_1447);
nor U2130 (N_2130,N_1868,N_1410);
nand U2131 (N_2131,N_1986,N_1697);
nor U2132 (N_2132,N_1460,N_212);
nor U2133 (N_2133,N_601,N_1058);
or U2134 (N_2134,N_166,N_1589);
and U2135 (N_2135,N_489,N_1566);
nor U2136 (N_2136,N_1525,N_1503);
or U2137 (N_2137,N_1512,N_1055);
nor U2138 (N_2138,N_1051,N_1352);
and U2139 (N_2139,N_1853,N_433);
nand U2140 (N_2140,N_1013,N_808);
or U2141 (N_2141,N_942,N_922);
or U2142 (N_2142,N_607,N_419);
nor U2143 (N_2143,N_979,N_783);
nor U2144 (N_2144,N_1618,N_1015);
nand U2145 (N_2145,N_1835,N_874);
and U2146 (N_2146,N_804,N_1227);
nor U2147 (N_2147,N_302,N_1331);
or U2148 (N_2148,N_1289,N_1582);
and U2149 (N_2149,N_1002,N_1785);
or U2150 (N_2150,N_1878,N_20);
and U2151 (N_2151,N_1263,N_803);
and U2152 (N_2152,N_913,N_624);
nand U2153 (N_2153,N_315,N_1631);
nand U2154 (N_2154,N_1852,N_962);
or U2155 (N_2155,N_732,N_26);
or U2156 (N_2156,N_375,N_1451);
nor U2157 (N_2157,N_1208,N_83);
or U2158 (N_2158,N_448,N_1558);
or U2159 (N_2159,N_466,N_57);
and U2160 (N_2160,N_1022,N_283);
or U2161 (N_2161,N_1728,N_1174);
nor U2162 (N_2162,N_1605,N_1990);
and U2163 (N_2163,N_1281,N_583);
and U2164 (N_2164,N_988,N_1718);
or U2165 (N_2165,N_430,N_1759);
nor U2166 (N_2166,N_1074,N_1706);
and U2167 (N_2167,N_667,N_102);
nor U2168 (N_2168,N_896,N_1760);
nor U2169 (N_2169,N_178,N_1103);
or U2170 (N_2170,N_1563,N_45);
and U2171 (N_2171,N_138,N_314);
or U2172 (N_2172,N_1792,N_829);
xor U2173 (N_2173,N_100,N_209);
or U2174 (N_2174,N_1418,N_1704);
or U2175 (N_2175,N_1046,N_106);
or U2176 (N_2176,N_873,N_1001);
and U2177 (N_2177,N_717,N_592);
or U2178 (N_2178,N_226,N_1356);
xnor U2179 (N_2179,N_658,N_1908);
nand U2180 (N_2180,N_1992,N_1665);
and U2181 (N_2181,N_507,N_42);
nand U2182 (N_2182,N_1315,N_1274);
or U2183 (N_2183,N_892,N_441);
and U2184 (N_2184,N_611,N_1229);
nor U2185 (N_2185,N_1177,N_1468);
nand U2186 (N_2186,N_1633,N_1676);
or U2187 (N_2187,N_1650,N_317);
nor U2188 (N_2188,N_1909,N_697);
nor U2189 (N_2189,N_1742,N_816);
and U2190 (N_2190,N_1889,N_1801);
nor U2191 (N_2191,N_153,N_1765);
and U2192 (N_2192,N_1532,N_482);
nor U2193 (N_2193,N_562,N_631);
and U2194 (N_2194,N_11,N_1032);
nand U2195 (N_2195,N_1249,N_1606);
or U2196 (N_2196,N_812,N_884);
and U2197 (N_2197,N_1610,N_21);
and U2198 (N_2198,N_1200,N_1931);
nor U2199 (N_2199,N_290,N_734);
or U2200 (N_2200,N_1176,N_1333);
and U2201 (N_2201,N_1422,N_1234);
or U2202 (N_2202,N_1581,N_682);
xnor U2203 (N_2203,N_1194,N_1452);
nor U2204 (N_2204,N_1779,N_1989);
and U2205 (N_2205,N_1951,N_1226);
nor U2206 (N_2206,N_519,N_428);
nand U2207 (N_2207,N_1484,N_424);
and U2208 (N_2208,N_1096,N_546);
and U2209 (N_2209,N_1247,N_805);
nand U2210 (N_2210,N_856,N_116);
nor U2211 (N_2211,N_834,N_1660);
and U2212 (N_2212,N_774,N_835);
or U2213 (N_2213,N_1392,N_1542);
nor U2214 (N_2214,N_1839,N_342);
nand U2215 (N_2215,N_596,N_966);
and U2216 (N_2216,N_228,N_312);
or U2217 (N_2217,N_1000,N_737);
nand U2218 (N_2218,N_729,N_1771);
nor U2219 (N_2219,N_1475,N_412);
and U2220 (N_2220,N_1689,N_330);
or U2221 (N_2221,N_971,N_1316);
nand U2222 (N_2222,N_76,N_288);
or U2223 (N_2223,N_521,N_1182);
nand U2224 (N_2224,N_47,N_410);
nand U2225 (N_2225,N_1034,N_82);
or U2226 (N_2226,N_60,N_1886);
nor U2227 (N_2227,N_589,N_1667);
or U2228 (N_2228,N_1823,N_1945);
and U2229 (N_2229,N_768,N_1736);
or U2230 (N_2230,N_861,N_726);
nor U2231 (N_2231,N_255,N_1138);
nand U2232 (N_2232,N_533,N_568);
nand U2233 (N_2233,N_1466,N_1520);
nand U2234 (N_2234,N_436,N_1598);
nand U2235 (N_2235,N_495,N_1493);
and U2236 (N_2236,N_846,N_524);
nor U2237 (N_2237,N_456,N_1919);
or U2238 (N_2238,N_1106,N_1056);
and U2239 (N_2239,N_746,N_1117);
and U2240 (N_2240,N_1590,N_1464);
or U2241 (N_2241,N_1600,N_1438);
and U2242 (N_2242,N_24,N_1186);
or U2243 (N_2243,N_1938,N_1150);
or U2244 (N_2244,N_397,N_517);
or U2245 (N_2245,N_512,N_1259);
nor U2246 (N_2246,N_625,N_407);
nand U2247 (N_2247,N_1377,N_941);
or U2248 (N_2248,N_219,N_725);
nor U2249 (N_2249,N_1012,N_1072);
or U2250 (N_2250,N_1415,N_854);
or U2251 (N_2251,N_779,N_526);
and U2252 (N_2252,N_1470,N_1500);
and U2253 (N_2253,N_1491,N_842);
and U2254 (N_2254,N_262,N_472);
and U2255 (N_2255,N_461,N_270);
nand U2256 (N_2256,N_827,N_677);
or U2257 (N_2257,N_1890,N_1047);
and U2258 (N_2258,N_1968,N_558);
and U2259 (N_2259,N_1809,N_548);
nor U2260 (N_2260,N_1538,N_1233);
nor U2261 (N_2261,N_387,N_654);
nor U2262 (N_2262,N_471,N_1813);
or U2263 (N_2263,N_711,N_1634);
and U2264 (N_2264,N_1465,N_1329);
or U2265 (N_2265,N_738,N_1677);
or U2266 (N_2266,N_1498,N_1271);
nand U2267 (N_2267,N_1764,N_523);
nand U2268 (N_2268,N_260,N_981);
and U2269 (N_2269,N_1528,N_1975);
or U2270 (N_2270,N_380,N_156);
and U2271 (N_2271,N_72,N_151);
or U2272 (N_2272,N_70,N_1654);
nor U2273 (N_2273,N_684,N_477);
or U2274 (N_2274,N_1957,N_1016);
xnor U2275 (N_2275,N_1243,N_1947);
and U2276 (N_2276,N_366,N_188);
nand U2277 (N_2277,N_840,N_126);
and U2278 (N_2278,N_229,N_1425);
nand U2279 (N_2279,N_295,N_1173);
nor U2280 (N_2280,N_1467,N_815);
nor U2281 (N_2281,N_1078,N_192);
and U2282 (N_2282,N_1946,N_1856);
or U2283 (N_2283,N_1640,N_1299);
and U2284 (N_2284,N_1144,N_259);
or U2285 (N_2285,N_688,N_25);
or U2286 (N_2286,N_1880,N_529);
nand U2287 (N_2287,N_1690,N_344);
and U2288 (N_2288,N_135,N_227);
xor U2289 (N_2289,N_197,N_555);
and U2290 (N_2290,N_22,N_1146);
and U2291 (N_2291,N_382,N_52);
and U2292 (N_2292,N_492,N_1405);
and U2293 (N_2293,N_554,N_1323);
nor U2294 (N_2294,N_1549,N_1006);
nor U2295 (N_2295,N_65,N_353);
or U2296 (N_2296,N_1678,N_1321);
nor U2297 (N_2297,N_739,N_683);
and U2298 (N_2298,N_1359,N_1241);
or U2299 (N_2299,N_414,N_591);
or U2300 (N_2300,N_455,N_791);
and U2301 (N_2301,N_1171,N_544);
and U2302 (N_2302,N_895,N_797);
and U2303 (N_2303,N_108,N_1504);
or U2304 (N_2304,N_478,N_1430);
nor U2305 (N_2305,N_112,N_1049);
nor U2306 (N_2306,N_356,N_1565);
and U2307 (N_2307,N_1435,N_618);
or U2308 (N_2308,N_394,N_689);
nand U2309 (N_2309,N_1787,N_365);
or U2310 (N_2310,N_824,N_164);
and U2311 (N_2311,N_128,N_1381);
nor U2312 (N_2312,N_1903,N_1747);
or U2313 (N_2313,N_144,N_615);
or U2314 (N_2314,N_225,N_1887);
and U2315 (N_2315,N_1983,N_174);
nand U2316 (N_2316,N_263,N_934);
nor U2317 (N_2317,N_801,N_1658);
nand U2318 (N_2318,N_1050,N_360);
nor U2319 (N_2319,N_348,N_325);
nand U2320 (N_2320,N_459,N_254);
nand U2321 (N_2321,N_902,N_1985);
or U2322 (N_2322,N_1408,N_733);
and U2323 (N_2323,N_1883,N_125);
nor U2324 (N_2324,N_1698,N_1626);
and U2325 (N_2325,N_621,N_778);
or U2326 (N_2326,N_409,N_1857);
and U2327 (N_2327,N_1337,N_557);
and U2328 (N_2328,N_675,N_553);
or U2329 (N_2329,N_1105,N_1413);
nor U2330 (N_2330,N_1863,N_1472);
nor U2331 (N_2331,N_866,N_1722);
nor U2332 (N_2332,N_1014,N_1960);
nor U2333 (N_2333,N_784,N_1596);
nand U2334 (N_2334,N_1937,N_66);
or U2335 (N_2335,N_1712,N_720);
and U2336 (N_2336,N_705,N_576);
and U2337 (N_2337,N_1979,N_279);
or U2338 (N_2338,N_904,N_917);
or U2339 (N_2339,N_885,N_1346);
nand U2340 (N_2340,N_1025,N_1628);
or U2341 (N_2341,N_1152,N_1204);
or U2342 (N_2342,N_1670,N_285);
nor U2343 (N_2343,N_1007,N_1637);
xnor U2344 (N_2344,N_1534,N_943);
and U2345 (N_2345,N_272,N_105);
and U2346 (N_2346,N_1694,N_1192);
and U2347 (N_2347,N_362,N_1964);
and U2348 (N_2348,N_69,N_924);
nand U2349 (N_2349,N_1763,N_1292);
and U2350 (N_2350,N_1509,N_1332);
nor U2351 (N_2351,N_763,N_501);
nand U2352 (N_2352,N_434,N_142);
nor U2353 (N_2353,N_539,N_1344);
nand U2354 (N_2354,N_1486,N_1820);
nor U2355 (N_2355,N_1188,N_680);
xnor U2356 (N_2356,N_284,N_503);
and U2357 (N_2357,N_146,N_953);
nor U2358 (N_2358,N_1501,N_1523);
and U2359 (N_2359,N_1157,N_173);
and U2360 (N_2360,N_1481,N_1057);
or U2361 (N_2361,N_976,N_331);
or U2362 (N_2362,N_1816,N_499);
nor U2363 (N_2363,N_109,N_1613);
or U2364 (N_2364,N_990,N_96);
and U2365 (N_2365,N_416,N_657);
or U2366 (N_2366,N_1578,N_1490);
nand U2367 (N_2367,N_1312,N_678);
nand U2368 (N_2368,N_1821,N_1896);
nand U2369 (N_2369,N_1619,N_1730);
xnor U2370 (N_2370,N_612,N_1443);
or U2371 (N_2371,N_1448,N_1358);
nor U2372 (N_2372,N_437,N_93);
or U2373 (N_2373,N_1603,N_371);
nor U2374 (N_2374,N_1180,N_1541);
or U2375 (N_2375,N_1686,N_1855);
nand U2376 (N_2376,N_646,N_337);
nor U2377 (N_2377,N_771,N_1151);
nor U2378 (N_2378,N_1485,N_882);
nand U2379 (N_2379,N_656,N_673);
nand U2380 (N_2380,N_1065,N_1379);
or U2381 (N_2381,N_915,N_1551);
nor U2382 (N_2382,N_1286,N_316);
or U2383 (N_2383,N_1750,N_1089);
nor U2384 (N_2384,N_821,N_859);
nand U2385 (N_2385,N_1705,N_460);
and U2386 (N_2386,N_415,N_374);
or U2387 (N_2387,N_613,N_1727);
or U2388 (N_2388,N_1876,N_1735);
nor U2389 (N_2389,N_1866,N_782);
nand U2390 (N_2390,N_1162,N_996);
nor U2391 (N_2391,N_1588,N_1818);
nand U2392 (N_2392,N_378,N_1649);
or U2393 (N_2393,N_1720,N_1745);
nor U2394 (N_2394,N_610,N_789);
and U2395 (N_2395,N_1757,N_1796);
and U2396 (N_2396,N_1725,N_645);
and U2397 (N_2397,N_175,N_1819);
and U2398 (N_2398,N_1328,N_651);
or U2399 (N_2399,N_1904,N_1683);
or U2400 (N_2400,N_1374,N_1595);
nor U2401 (N_2401,N_335,N_810);
or U2402 (N_2402,N_439,N_1617);
nand U2403 (N_2403,N_248,N_1700);
or U2404 (N_2404,N_1348,N_298);
and U2405 (N_2405,N_1406,N_975);
nor U2406 (N_2406,N_1806,N_1726);
or U2407 (N_2407,N_989,N_593);
nor U2408 (N_2408,N_29,N_1755);
or U2409 (N_2409,N_1426,N_869);
and U2410 (N_2410,N_246,N_1095);
nand U2411 (N_2411,N_629,N_238);
or U2412 (N_2412,N_536,N_1875);
or U2413 (N_2413,N_1228,N_1441);
or U2414 (N_2414,N_838,N_163);
nor U2415 (N_2415,N_1614,N_940);
nand U2416 (N_2416,N_587,N_391);
or U2417 (N_2417,N_1060,N_422);
nor U2418 (N_2418,N_1155,N_1540);
nand U2419 (N_2419,N_99,N_1343);
and U2420 (N_2420,N_427,N_1547);
and U2421 (N_2421,N_1607,N_122);
nand U2422 (N_2422,N_1939,N_1112);
or U2423 (N_2423,N_271,N_278);
xor U2424 (N_2424,N_1090,N_34);
nor U2425 (N_2425,N_676,N_413);
nor U2426 (N_2426,N_659,N_1145);
nand U2427 (N_2427,N_1397,N_1133);
nand U2428 (N_2428,N_1811,N_1766);
and U2429 (N_2429,N_321,N_75);
nor U2430 (N_2430,N_1300,N_479);
or U2431 (N_2431,N_935,N_1197);
nor U2432 (N_2432,N_860,N_1178);
or U2433 (N_2433,N_1461,N_1181);
nor U2434 (N_2434,N_336,N_1902);
nor U2435 (N_2435,N_541,N_1559);
and U2436 (N_2436,N_319,N_454);
and U2437 (N_2437,N_294,N_1364);
or U2438 (N_2438,N_145,N_1334);
or U2439 (N_2439,N_998,N_1815);
or U2440 (N_2440,N_987,N_528);
nand U2441 (N_2441,N_531,N_1248);
or U2442 (N_2442,N_1682,N_1685);
and U2443 (N_2443,N_1761,N_1018);
nand U2444 (N_2444,N_381,N_1266);
nand U2445 (N_2445,N_1167,N_547);
nor U2446 (N_2446,N_1240,N_634);
or U2447 (N_2447,N_762,N_1187);
nor U2448 (N_2448,N_446,N_1061);
nand U2449 (N_2449,N_749,N_847);
nor U2450 (N_2450,N_111,N_9);
and U2451 (N_2451,N_1283,N_757);
and U2452 (N_2452,N_1965,N_1417);
xnor U2453 (N_2453,N_1526,N_1833);
and U2454 (N_2454,N_1185,N_1516);
and U2455 (N_2455,N_1859,N_1918);
and U2456 (N_2456,N_203,N_1211);
or U2457 (N_2457,N_1402,N_870);
or U2458 (N_2458,N_1548,N_1892);
nor U2459 (N_2459,N_1630,N_666);
and U2460 (N_2460,N_1108,N_469);
xor U2461 (N_2461,N_1808,N_1232);
nand U2462 (N_2462,N_181,N_642);
or U2463 (N_2463,N_1829,N_597);
nor U2464 (N_2464,N_1862,N_1166);
or U2465 (N_2465,N_806,N_1279);
nor U2466 (N_2466,N_691,N_58);
nor U2467 (N_2467,N_1380,N_1684);
nor U2468 (N_2468,N_1390,N_328);
nor U2469 (N_2469,N_1997,N_402);
nor U2470 (N_2470,N_1719,N_619);
nor U2471 (N_2471,N_700,N_844);
nand U2472 (N_2472,N_1827,N_236);
xnor U2473 (N_2473,N_211,N_964);
nor U2474 (N_2474,N_216,N_550);
and U2475 (N_2475,N_758,N_97);
nand U2476 (N_2476,N_1778,N_372);
nor U2477 (N_2477,N_119,N_1782);
nor U2478 (N_2478,N_1314,N_442);
nor U2479 (N_2479,N_282,N_1462);
nor U2480 (N_2480,N_1483,N_710);
nand U2481 (N_2481,N_1010,N_813);
and U2482 (N_2482,N_1132,N_1793);
nand U2483 (N_2483,N_1431,N_1734);
nand U2484 (N_2484,N_573,N_405);
or U2485 (N_2485,N_217,N_1748);
or U2486 (N_2486,N_117,N_668);
nand U2487 (N_2487,N_928,N_1218);
or U2488 (N_2488,N_1391,N_655);
nor U2489 (N_2489,N_986,N_1252);
nor U2490 (N_2490,N_1715,N_1309);
or U2491 (N_2491,N_1732,N_1119);
xnor U2492 (N_2492,N_1433,N_1024);
or U2493 (N_2493,N_653,N_1508);
or U2494 (N_2494,N_1,N_1881);
and U2495 (N_2495,N_49,N_1324);
nand U2496 (N_2496,N_377,N_1361);
or U2497 (N_2497,N_129,N_127);
nor U2498 (N_2498,N_1749,N_1661);
and U2499 (N_2499,N_1262,N_1463);
and U2500 (N_2500,N_168,N_1335);
nand U2501 (N_2501,N_1221,N_1159);
and U2502 (N_2502,N_1781,N_1800);
and U2503 (N_2503,N_616,N_623);
or U2504 (N_2504,N_1041,N_1962);
nor U2505 (N_2505,N_18,N_351);
nand U2506 (N_2506,N_909,N_1127);
and U2507 (N_2507,N_1026,N_324);
and U2508 (N_2508,N_234,N_276);
and U2509 (N_2509,N_418,N_1754);
and U2510 (N_2510,N_1555,N_1858);
and U2511 (N_2511,N_149,N_1854);
nand U2512 (N_2512,N_1237,N_88);
and U2513 (N_2513,N_1679,N_86);
and U2514 (N_2514,N_300,N_1774);
nor U2515 (N_2515,N_767,N_636);
nand U2516 (N_2516,N_551,N_582);
nand U2517 (N_2517,N_1669,N_560);
nand U2518 (N_2518,N_1936,N_903);
and U2519 (N_2519,N_396,N_1242);
nor U2520 (N_2520,N_1707,N_1977);
nor U2521 (N_2521,N_564,N_1455);
and U2522 (N_2522,N_841,N_1687);
or U2523 (N_2523,N_139,N_1326);
nor U2524 (N_2524,N_1220,N_927);
or U2525 (N_2525,N_1416,N_265);
and U2526 (N_2526,N_1436,N_1214);
or U2527 (N_2527,N_500,N_376);
nor U2528 (N_2528,N_532,N_1043);
nor U2529 (N_2529,N_855,N_1142);
nor U2530 (N_2530,N_741,N_239);
nor U2531 (N_2531,N_1120,N_85);
nand U2532 (N_2532,N_1524,N_823);
or U2533 (N_2533,N_303,N_886);
or U2534 (N_2534,N_575,N_1378);
and U2535 (N_2535,N_310,N_622);
or U2536 (N_2536,N_1851,N_1088);
nand U2537 (N_2537,N_1053,N_1272);
or U2538 (N_2538,N_132,N_712);
nand U2539 (N_2539,N_770,N_648);
or U2540 (N_2540,N_1737,N_258);
and U2541 (N_2541,N_1620,N_969);
nor U2542 (N_2542,N_1570,N_1623);
and U2543 (N_2543,N_1743,N_1277);
nand U2544 (N_2544,N_1269,N_745);
and U2545 (N_2545,N_421,N_386);
nor U2546 (N_2546,N_1663,N_232);
nor U2547 (N_2547,N_617,N_1161);
nor U2548 (N_2548,N_1276,N_1407);
xnor U2549 (N_2549,N_1137,N_465);
nor U2550 (N_2550,N_1083,N_177);
nand U2551 (N_2551,N_184,N_425);
or U2552 (N_2552,N_1432,N_84);
and U2553 (N_2553,N_727,N_242);
or U2554 (N_2554,N_708,N_951);
and U2555 (N_2555,N_1336,N_268);
nand U2556 (N_2556,N_932,N_1973);
nand U2557 (N_2557,N_1030,N_218);
or U2558 (N_2558,N_1365,N_408);
nor U2559 (N_2559,N_939,N_641);
and U2560 (N_2560,N_233,N_200);
and U2561 (N_2561,N_488,N_464);
and U2562 (N_2562,N_257,N_1478);
nor U2563 (N_2563,N_1147,N_1664);
and U2564 (N_2564,N_1310,N_487);
nor U2565 (N_2565,N_13,N_1371);
or U2566 (N_2566,N_1543,N_766);
nor U2567 (N_2567,N_724,N_581);
nand U2568 (N_2568,N_1789,N_1585);
nand U2569 (N_2569,N_980,N_1768);
nand U2570 (N_2570,N_1411,N_534);
or U2571 (N_2571,N_457,N_1136);
and U2572 (N_2572,N_639,N_1810);
nor U2573 (N_2573,N_1934,N_1203);
or U2574 (N_2574,N_256,N_1783);
nand U2575 (N_2575,N_1028,N_605);
nor U2576 (N_2576,N_1959,N_1874);
nor U2577 (N_2577,N_1170,N_1586);
and U2578 (N_2578,N_152,N_671);
or U2579 (N_2579,N_1224,N_598);
nor U2580 (N_2580,N_1515,N_1533);
nand U2581 (N_2581,N_721,N_1039);
nor U2582 (N_2582,N_1926,N_179);
or U2583 (N_2583,N_31,N_914);
nor U2584 (N_2584,N_1553,N_1693);
nand U2585 (N_2585,N_865,N_494);
or U2586 (N_2586,N_1831,N_1376);
nor U2587 (N_2587,N_728,N_1967);
and U2588 (N_2588,N_1134,N_1791);
and U2589 (N_2589,N_1943,N_118);
and U2590 (N_2590,N_1434,N_740);
nor U2591 (N_2591,N_41,N_1941);
and U2592 (N_2592,N_837,N_1445);
or U2593 (N_2593,N_307,N_37);
nand U2594 (N_2594,N_287,N_1940);
nand U2595 (N_2595,N_1651,N_1917);
nor U2596 (N_2596,N_193,N_756);
nand U2597 (N_2597,N_1008,N_44);
or U2598 (N_2598,N_1202,N_467);
or U2599 (N_2599,N_1383,N_540);
and U2600 (N_2600,N_1773,N_1882);
and U2601 (N_2601,N_1313,N_333);
and U2602 (N_2602,N_1780,N_98);
nor U2603 (N_2603,N_182,N_1389);
and U2604 (N_2604,N_1885,N_1996);
and U2605 (N_2605,N_692,N_811);
and U2606 (N_2606,N_901,N_753);
nand U2607 (N_2607,N_269,N_1703);
and U2608 (N_2608,N_1799,N_1519);
nand U2609 (N_2609,N_752,N_120);
nor U2610 (N_2610,N_716,N_1496);
nor U2611 (N_2611,N_484,N_347);
and U2612 (N_2612,N_385,N_1497);
or U2613 (N_2613,N_1444,N_580);
nand U2614 (N_2614,N_1537,N_1454);
nor U2615 (N_2615,N_350,N_1573);
and U2616 (N_2616,N_395,N_1308);
and U2617 (N_2617,N_1295,N_652);
and U2618 (N_2618,N_137,N_1842);
and U2619 (N_2619,N_1724,N_1419);
nand U2620 (N_2620,N_411,N_792);
and U2621 (N_2621,N_958,N_62);
nand U2622 (N_2622,N_1615,N_556);
or U2623 (N_2623,N_910,N_920);
nand U2624 (N_2624,N_747,N_1871);
nor U2625 (N_2625,N_1169,N_1429);
and U2626 (N_2626,N_440,N_999);
nand U2627 (N_2627,N_1495,N_669);
or U2628 (N_2628,N_1135,N_150);
nand U2629 (N_2629,N_1505,N_930);
nand U2630 (N_2630,N_158,N_445);
xor U2631 (N_2631,N_1729,N_1674);
and U2632 (N_2632,N_1035,N_1942);
nand U2633 (N_2633,N_851,N_794);
nand U2634 (N_2634,N_1382,N_1033);
nor U2635 (N_2635,N_449,N_588);
or U2636 (N_2636,N_161,N_1777);
nor U2637 (N_2637,N_124,N_392);
nor U2638 (N_2638,N_1125,N_1924);
or U2639 (N_2639,N_765,N_340);
nand U2640 (N_2640,N_1363,N_1834);
nor U2641 (N_2641,N_1550,N_1070);
or U2642 (N_2642,N_698,N_64);
nor U2643 (N_2643,N_826,N_1535);
nor U2644 (N_2644,N_799,N_868);
nor U2645 (N_2645,N_318,N_140);
and U2646 (N_2646,N_984,N_1270);
nand U2647 (N_2647,N_609,N_1052);
nand U2648 (N_2648,N_1629,N_252);
nand U2649 (N_2649,N_1306,N_1318);
and U2650 (N_2650,N_802,N_363);
or U2651 (N_2651,N_945,N_289);
nand U2652 (N_2652,N_858,N_1675);
nor U2653 (N_2653,N_742,N_1102);
nor U2654 (N_2654,N_871,N_577);
or U2655 (N_2655,N_1122,N_722);
nor U2656 (N_2656,N_1844,N_79);
nor U2657 (N_2657,N_1861,N_447);
nand U2658 (N_2658,N_1884,N_898);
nand U2659 (N_2659,N_1702,N_1701);
and U2660 (N_2660,N_220,N_1952);
and U2661 (N_2661,N_1225,N_1158);
and U2662 (N_2662,N_1287,N_687);
nand U2663 (N_2663,N_406,N_561);
and U2664 (N_2664,N_369,N_907);
nand U2665 (N_2665,N_148,N_1275);
nand U2666 (N_2666,N_508,N_1804);
and U2667 (N_2667,N_936,N_1265);
or U2668 (N_2668,N_349,N_187);
xnor U2669 (N_2669,N_959,N_1149);
and U2670 (N_2670,N_1925,N_565);
or U2671 (N_2671,N_1172,N_1912);
nand U2672 (N_2672,N_92,N_563);
nor U2673 (N_2673,N_1268,N_1398);
and U2674 (N_2674,N_438,N_690);
xnor U2675 (N_2675,N_879,N_1647);
nand U2676 (N_2676,N_355,N_703);
and U2677 (N_2677,N_404,N_832);
and U2678 (N_2678,N_1209,N_230);
and U2679 (N_2679,N_1076,N_167);
and U2680 (N_2680,N_311,N_603);
nand U2681 (N_2681,N_224,N_911);
and U2682 (N_2682,N_1929,N_543);
and U2683 (N_2683,N_1351,N_730);
nand U2684 (N_2684,N_1244,N_320);
nor U2685 (N_2685,N_574,N_326);
or U2686 (N_2686,N_1864,N_1260);
nand U2687 (N_2687,N_848,N_1625);
nand U2688 (N_2688,N_1982,N_1353);
nor U2689 (N_2689,N_1544,N_51);
nor U2690 (N_2690,N_1639,N_426);
nor U2691 (N_2691,N_836,N_1017);
nor U2692 (N_2692,N_309,N_250);
nor U2693 (N_2693,N_101,N_944);
nand U2694 (N_2694,N_993,N_1213);
xor U2695 (N_2695,N_1594,N_567);
or U2696 (N_2696,N_1205,N_136);
nor U2697 (N_2697,N_839,N_1949);
nor U2698 (N_2698,N_1978,N_862);
or U2699 (N_2699,N_91,N_1914);
nor U2700 (N_2700,N_566,N_1254);
and U2701 (N_2701,N_297,N_1999);
or U2702 (N_2702,N_470,N_1518);
or U2703 (N_2703,N_1298,N_1984);
and U2704 (N_2704,N_889,N_890);
nor U2705 (N_2705,N_195,N_1338);
nand U2706 (N_2706,N_1264,N_830);
nor U2707 (N_2707,N_1251,N_735);
and U2708 (N_2708,N_1837,N_154);
nor U2709 (N_2709,N_1906,N_760);
nor U2710 (N_2710,N_1037,N_1141);
nand U2711 (N_2711,N_1459,N_38);
xor U2712 (N_2712,N_1082,N_1655);
nor U2713 (N_2713,N_1976,N_274);
and U2714 (N_2714,N_1894,N_1009);
nand U2715 (N_2715,N_1604,N_1427);
nor U2716 (N_2716,N_367,N_1094);
nor U2717 (N_2717,N_1708,N_1746);
nand U2718 (N_2718,N_908,N_1245);
nor U2719 (N_2719,N_569,N_947);
nand U2720 (N_2720,N_828,N_1304);
and U2721 (N_2721,N_1681,N_1536);
nand U2722 (N_2722,N_509,N_1846);
or U2723 (N_2723,N_134,N_176);
nand U2724 (N_2724,N_502,N_1609);
or U2725 (N_2725,N_1153,N_1930);
and U2726 (N_2726,N_198,N_359);
or U2727 (N_2727,N_1560,N_809);
nor U2728 (N_2728,N_948,N_1591);
and U2729 (N_2729,N_1897,N_1273);
nor U2730 (N_2730,N_950,N_1988);
and U2731 (N_2731,N_1710,N_1156);
or U2732 (N_2732,N_788,N_1870);
or U2733 (N_2733,N_1116,N_952);
nor U2734 (N_2734,N_900,N_518);
and U2735 (N_2735,N_681,N_595);
nand U2736 (N_2736,N_1222,N_1160);
nor U2737 (N_2737,N_1471,N_1969);
nor U2738 (N_2738,N_663,N_305);
nand U2739 (N_2739,N_143,N_48);
and U2740 (N_2740,N_1404,N_974);
nor U2741 (N_2741,N_665,N_893);
or U2742 (N_2742,N_1772,N_281);
nor U2743 (N_2743,N_1092,N_1869);
nand U2744 (N_2744,N_1974,N_1502);
nor U2745 (N_2745,N_1063,N_1104);
nor U2746 (N_2746,N_452,N_946);
nand U2747 (N_2747,N_707,N_1109);
or U2748 (N_2748,N_1368,N_755);
nor U2749 (N_2749,N_1873,N_520);
nor U2750 (N_2750,N_1571,N_1482);
and U2751 (N_2751,N_1414,N_1458);
nand U2752 (N_2752,N_1322,N_776);
or U2753 (N_2753,N_306,N_1355);
nor U2754 (N_2754,N_991,N_1569);
or U2755 (N_2755,N_510,N_590);
nor U2756 (N_2756,N_661,N_343);
and U2757 (N_2757,N_12,N_1601);
nand U2758 (N_2758,N_244,N_1473);
or U2759 (N_2759,N_1184,N_965);
nor U2760 (N_2760,N_1662,N_1062);
nor U2761 (N_2761,N_586,N_1691);
and U2762 (N_2762,N_1148,N_1583);
and U2763 (N_2763,N_280,N_777);
and U2764 (N_2764,N_822,N_77);
and U2765 (N_2765,N_1673,N_1696);
nand U2766 (N_2766,N_1163,N_435);
nor U2767 (N_2767,N_1913,N_1488);
nand U2768 (N_2768,N_1450,N_1042);
nor U2769 (N_2769,N_1370,N_463);
and U2770 (N_2770,N_949,N_1479);
or U2771 (N_2771,N_864,N_1666);
and U2772 (N_2772,N_453,N_1420);
and U2773 (N_2773,N_1739,N_223);
and U2774 (N_2774,N_1091,N_1695);
and U2775 (N_2775,N_55,N_1064);
nand U2776 (N_2776,N_332,N_714);
nand U2777 (N_2777,N_831,N_1107);
nor U2778 (N_2778,N_483,N_1972);
nand U2779 (N_2779,N_679,N_1423);
or U2780 (N_2780,N_1121,N_713);
or U2781 (N_2781,N_780,N_293);
or U2782 (N_2782,N_759,N_180);
or U2783 (N_2783,N_1325,N_458);
or U2784 (N_2784,N_393,N_1216);
nand U2785 (N_2785,N_1059,N_1636);
nor U2786 (N_2786,N_1721,N_1223);
nand U2787 (N_2787,N_43,N_1100);
and U2788 (N_2788,N_709,N_1794);
nand U2789 (N_2789,N_1713,N_1751);
nor U2790 (N_2790,N_1958,N_1907);
or U2791 (N_2791,N_883,N_1256);
nand U2792 (N_2792,N_1517,N_354);
nand U2793 (N_2793,N_5,N_1756);
and U2794 (N_2794,N_1552,N_530);
nor U2795 (N_2795,N_820,N_800);
nand U2796 (N_2796,N_1175,N_334);
nor U2797 (N_2797,N_1067,N_1653);
nor U2798 (N_2798,N_4,N_130);
nand U2799 (N_2799,N_696,N_327);
nand U2800 (N_2800,N_204,N_277);
or U2801 (N_2801,N_1075,N_1021);
nand U2802 (N_2802,N_1627,N_660);
or U2803 (N_2803,N_1375,N_538);
nand U2804 (N_2804,N_1802,N_1529);
nor U2805 (N_2805,N_1212,N_888);
and U2806 (N_2806,N_388,N_115);
nor U2807 (N_2807,N_403,N_1044);
and U2808 (N_2808,N_80,N_1246);
nor U2809 (N_2809,N_1915,N_1085);
nor U2810 (N_2810,N_1671,N_451);
nand U2811 (N_2811,N_1031,N_702);
nand U2812 (N_2812,N_1165,N_1898);
nand U2813 (N_2813,N_1850,N_1305);
nand U2814 (N_2814,N_1910,N_1769);
and U2815 (N_2815,N_649,N_1164);
nand U2816 (N_2816,N_400,N_1168);
nor U2817 (N_2817,N_468,N_245);
xnor U2818 (N_2818,N_81,N_627);
nand U2819 (N_2819,N_159,N_1527);
nor U2820 (N_2820,N_304,N_1029);
and U2821 (N_2821,N_240,N_206);
nor U2822 (N_2822,N_506,N_1327);
or U2823 (N_2823,N_87,N_549);
nand U2824 (N_2824,N_1003,N_95);
nor U2825 (N_2825,N_429,N_1303);
nand U2826 (N_2826,N_925,N_1879);
nor U2827 (N_2827,N_1469,N_1201);
nor U2828 (N_2828,N_1048,N_1954);
nand U2829 (N_2829,N_462,N_1183);
or U2830 (N_2830,N_215,N_59);
or U2831 (N_2831,N_1126,N_863);
or U2832 (N_2832,N_1296,N_498);
or U2833 (N_2833,N_1980,N_1546);
or U2834 (N_2834,N_1257,N_485);
nand U2835 (N_2835,N_1401,N_1506);
or U2836 (N_2836,N_399,N_1612);
nor U2837 (N_2837,N_972,N_1901);
and U2838 (N_2838,N_54,N_825);
and U2839 (N_2839,N_1215,N_513);
nand U2840 (N_2840,N_1210,N_1840);
or U2841 (N_2841,N_1179,N_1795);
nand U2842 (N_2842,N_715,N_814);
nor U2843 (N_2843,N_205,N_1836);
nand U2844 (N_2844,N_1611,N_718);
nor U2845 (N_2845,N_906,N_1294);
or U2846 (N_2846,N_1692,N_202);
and U2847 (N_2847,N_1113,N_56);
or U2848 (N_2848,N_1825,N_1258);
and U2849 (N_2849,N_1339,N_1568);
and U2850 (N_2850,N_103,N_1019);
and U2851 (N_2851,N_647,N_339);
and U2852 (N_2852,N_1577,N_630);
or U2853 (N_2853,N_1762,N_364);
and U2854 (N_2854,N_1255,N_1409);
or U2855 (N_2855,N_1341,N_921);
and U2856 (N_2856,N_795,N_39);
nand U2857 (N_2857,N_338,N_1261);
nor U2858 (N_2858,N_28,N_104);
or U2859 (N_2859,N_744,N_1776);
and U2860 (N_2860,N_1349,N_957);
and U2861 (N_2861,N_420,N_1530);
nand U2862 (N_2862,N_231,N_1872);
and U2863 (N_2863,N_473,N_1932);
nand U2864 (N_2864,N_1921,N_383);
and U2865 (N_2865,N_1387,N_516);
and U2866 (N_2866,N_1584,N_1656);
nand U2867 (N_2867,N_475,N_273);
nand U2868 (N_2868,N_1539,N_1084);
or U2869 (N_2869,N_1847,N_769);
nand U2870 (N_2870,N_1832,N_1236);
nor U2871 (N_2871,N_1731,N_559);
or U2872 (N_2872,N_417,N_486);
and U2873 (N_2873,N_1824,N_432);
nand U2874 (N_2874,N_1360,N_113);
nor U2875 (N_2875,N_926,N_15);
nor U2876 (N_2876,N_481,N_931);
and U2877 (N_2877,N_1198,N_1456);
and U2878 (N_2878,N_1118,N_1077);
or U2879 (N_2879,N_978,N_1699);
nor U2880 (N_2880,N_1865,N_785);
nor U2881 (N_2881,N_1767,N_50);
nand U2882 (N_2882,N_545,N_1927);
and U2883 (N_2883,N_1867,N_1888);
nand U2884 (N_2884,N_1961,N_1130);
or U2885 (N_2885,N_1826,N_1004);
xnor U2886 (N_2886,N_701,N_1950);
or U2887 (N_2887,N_706,N_1576);
nor U2888 (N_2888,N_497,N_578);
nor U2889 (N_2889,N_275,N_614);
nand U2890 (N_2890,N_1711,N_833);
nand U2891 (N_2891,N_736,N_346);
and U2892 (N_2892,N_266,N_1709);
or U2893 (N_2893,N_1641,N_1301);
nor U2894 (N_2894,N_933,N_357);
nor U2895 (N_2895,N_644,N_110);
nand U2896 (N_2896,N_1928,N_384);
and U2897 (N_2897,N_853,N_1657);
and U2898 (N_2898,N_341,N_1412);
nand U2899 (N_2899,N_1027,N_1110);
and U2900 (N_2900,N_761,N_693);
nor U2901 (N_2901,N_183,N_956);
nor U2902 (N_2902,N_602,N_1798);
and U2903 (N_2903,N_1714,N_1293);
nand U2904 (N_2904,N_1190,N_155);
nor U2905 (N_2905,N_1557,N_1860);
nor U2906 (N_2906,N_968,N_1567);
and U2907 (N_2907,N_686,N_1624);
and U2908 (N_2908,N_1386,N_719);
or U2909 (N_2909,N_1599,N_221);
nor U2910 (N_2910,N_189,N_1893);
nand U2911 (N_2911,N_674,N_857);
or U2912 (N_2912,N_1564,N_672);
nand U2913 (N_2913,N_1399,N_1838);
or U2914 (N_2914,N_1944,N_992);
nand U2915 (N_2915,N_1267,N_1956);
and U2916 (N_2916,N_743,N_1717);
or U2917 (N_2917,N_843,N_1740);
nand U2918 (N_2918,N_1487,N_594);
nand U2919 (N_2919,N_1073,N_1079);
and U2920 (N_2920,N_201,N_1788);
and U2921 (N_2921,N_1081,N_955);
or U2922 (N_2922,N_358,N_1935);
nor U2923 (N_2923,N_572,N_1231);
and U2924 (N_2924,N_773,N_1848);
and U2925 (N_2925,N_970,N_796);
and U2926 (N_2926,N_191,N_1437);
nor U2927 (N_2927,N_1733,N_637);
and U2928 (N_2928,N_32,N_1394);
nor U2929 (N_2929,N_329,N_1449);
and U2930 (N_2930,N_121,N_764);
nor U2931 (N_2931,N_643,N_891);
nor U2932 (N_2932,N_1905,N_186);
or U2933 (N_2933,N_169,N_918);
or U2934 (N_2934,N_1993,N_1124);
or U2935 (N_2935,N_1330,N_704);
and U2936 (N_2936,N_750,N_664);
and U2937 (N_2937,N_1991,N_1531);
nand U2938 (N_2938,N_1545,N_390);
nor U2939 (N_2939,N_1797,N_1511);
nand U2940 (N_2940,N_53,N_923);
nor U2941 (N_2941,N_1217,N_1803);
nand U2942 (N_2942,N_379,N_185);
or U2943 (N_2943,N_1916,N_1716);
and U2944 (N_2944,N_444,N_1642);
nor U2945 (N_2945,N_213,N_345);
nand U2946 (N_2946,N_1366,N_1285);
and U2947 (N_2947,N_208,N_967);
nor U2948 (N_2948,N_600,N_1817);
or U2949 (N_2949,N_1981,N_496);
or U2950 (N_2950,N_1933,N_1572);
nor U2951 (N_2951,N_286,N_638);
nand U2952 (N_2952,N_1457,N_63);
and U2953 (N_2953,N_1239,N_1139);
nor U2954 (N_2954,N_635,N_1845);
nor U2955 (N_2955,N_1011,N_1384);
and U2956 (N_2956,N_1587,N_1499);
and U2957 (N_2957,N_94,N_748);
and U2958 (N_2958,N_1453,N_1123);
xor U2959 (N_2959,N_887,N_301);
or U2960 (N_2960,N_1738,N_1069);
nor U2961 (N_2961,N_852,N_373);
or U2962 (N_2962,N_7,N_1045);
or U2963 (N_2963,N_370,N_1963);
or U2964 (N_2964,N_1744,N_1199);
nor U2965 (N_2965,N_790,N_994);
nor U2966 (N_2966,N_1196,N_264);
or U2967 (N_2967,N_606,N_985);
nand U2968 (N_2968,N_1005,N_1513);
or U2969 (N_2969,N_1395,N_537);
or U2970 (N_2970,N_1284,N_46);
nor U2971 (N_2971,N_542,N_604);
and U2972 (N_2972,N_74,N_1114);
nor U2973 (N_2973,N_1080,N_1514);
and U2974 (N_2974,N_867,N_807);
nor U2975 (N_2975,N_961,N_493);
nand U2976 (N_2976,N_401,N_1971);
nor U2977 (N_2977,N_361,N_474);
and U2978 (N_2978,N_1345,N_1128);
nand U2979 (N_2979,N_1140,N_504);
nor U2980 (N_2980,N_1923,N_450);
and U2981 (N_2981,N_819,N_982);
nand U2982 (N_2982,N_1920,N_938);
or U2983 (N_2983,N_1290,N_880);
or U2984 (N_2984,N_954,N_1987);
nor U2985 (N_2985,N_1474,N_40);
nor U2986 (N_2986,N_1622,N_1741);
and U2987 (N_2987,N_1131,N_1320);
or U2988 (N_2988,N_1911,N_620);
nand U2989 (N_2989,N_876,N_1814);
and U2990 (N_2990,N_33,N_995);
nand U2991 (N_2991,N_30,N_1822);
and U2992 (N_2992,N_1086,N_296);
and U2993 (N_2993,N_1372,N_1593);
or U2994 (N_2994,N_1111,N_1561);
nand U2995 (N_2995,N_1189,N_685);
and U2996 (N_2996,N_1311,N_323);
nor U2997 (N_2997,N_261,N_1023);
or U2998 (N_2998,N_141,N_1753);
and U2999 (N_2999,N_1521,N_1849);
and U3000 (N_3000,N_1655,N_334);
nor U3001 (N_3001,N_201,N_786);
or U3002 (N_3002,N_875,N_1100);
nor U3003 (N_3003,N_1184,N_514);
nand U3004 (N_3004,N_618,N_541);
and U3005 (N_3005,N_1219,N_446);
nor U3006 (N_3006,N_1892,N_136);
nor U3007 (N_3007,N_191,N_1276);
or U3008 (N_3008,N_454,N_1894);
and U3009 (N_3009,N_1471,N_1499);
or U3010 (N_3010,N_618,N_1084);
nor U3011 (N_3011,N_1337,N_1209);
or U3012 (N_3012,N_756,N_405);
or U3013 (N_3013,N_743,N_705);
nor U3014 (N_3014,N_1343,N_1597);
nor U3015 (N_3015,N_1696,N_1184);
and U3016 (N_3016,N_144,N_1790);
and U3017 (N_3017,N_1692,N_871);
or U3018 (N_3018,N_1519,N_1886);
nor U3019 (N_3019,N_1065,N_1019);
nand U3020 (N_3020,N_1694,N_1534);
nand U3021 (N_3021,N_1502,N_153);
nand U3022 (N_3022,N_411,N_1341);
nand U3023 (N_3023,N_1228,N_898);
or U3024 (N_3024,N_736,N_392);
nor U3025 (N_3025,N_1805,N_1973);
nor U3026 (N_3026,N_1744,N_1225);
and U3027 (N_3027,N_946,N_625);
nand U3028 (N_3028,N_827,N_858);
nor U3029 (N_3029,N_1766,N_1373);
or U3030 (N_3030,N_16,N_1731);
nand U3031 (N_3031,N_1942,N_524);
or U3032 (N_3032,N_100,N_1234);
nand U3033 (N_3033,N_188,N_1041);
nor U3034 (N_3034,N_614,N_746);
nand U3035 (N_3035,N_1395,N_305);
or U3036 (N_3036,N_1848,N_442);
nand U3037 (N_3037,N_729,N_799);
or U3038 (N_3038,N_757,N_1570);
nor U3039 (N_3039,N_1529,N_1967);
nor U3040 (N_3040,N_754,N_770);
or U3041 (N_3041,N_560,N_214);
nand U3042 (N_3042,N_593,N_712);
and U3043 (N_3043,N_167,N_58);
and U3044 (N_3044,N_1151,N_1648);
nand U3045 (N_3045,N_1991,N_843);
nand U3046 (N_3046,N_521,N_1157);
and U3047 (N_3047,N_1703,N_51);
nand U3048 (N_3048,N_266,N_639);
or U3049 (N_3049,N_515,N_1384);
nor U3050 (N_3050,N_281,N_1292);
xor U3051 (N_3051,N_1391,N_491);
nor U3052 (N_3052,N_1569,N_1122);
and U3053 (N_3053,N_145,N_1651);
nor U3054 (N_3054,N_1056,N_686);
or U3055 (N_3055,N_967,N_1083);
nand U3056 (N_3056,N_836,N_1477);
and U3057 (N_3057,N_94,N_1984);
and U3058 (N_3058,N_619,N_1880);
or U3059 (N_3059,N_1367,N_1495);
and U3060 (N_3060,N_1605,N_375);
nand U3061 (N_3061,N_46,N_1149);
nand U3062 (N_3062,N_384,N_1694);
nor U3063 (N_3063,N_1185,N_1767);
nand U3064 (N_3064,N_1802,N_917);
nand U3065 (N_3065,N_1836,N_1944);
nor U3066 (N_3066,N_1779,N_590);
or U3067 (N_3067,N_94,N_29);
nand U3068 (N_3068,N_1586,N_1784);
or U3069 (N_3069,N_984,N_1854);
nor U3070 (N_3070,N_1015,N_1329);
nand U3071 (N_3071,N_1295,N_176);
and U3072 (N_3072,N_1066,N_139);
or U3073 (N_3073,N_1671,N_761);
nor U3074 (N_3074,N_742,N_1320);
and U3075 (N_3075,N_218,N_163);
or U3076 (N_3076,N_1462,N_1681);
or U3077 (N_3077,N_460,N_75);
or U3078 (N_3078,N_216,N_1328);
or U3079 (N_3079,N_724,N_1646);
and U3080 (N_3080,N_121,N_1521);
and U3081 (N_3081,N_1777,N_960);
and U3082 (N_3082,N_898,N_1204);
and U3083 (N_3083,N_1755,N_1131);
nor U3084 (N_3084,N_243,N_1121);
nor U3085 (N_3085,N_1604,N_1311);
xnor U3086 (N_3086,N_1620,N_418);
xnor U3087 (N_3087,N_1919,N_823);
and U3088 (N_3088,N_80,N_1780);
nor U3089 (N_3089,N_302,N_166);
or U3090 (N_3090,N_1424,N_1302);
and U3091 (N_3091,N_1721,N_637);
nand U3092 (N_3092,N_1,N_1966);
nand U3093 (N_3093,N_1466,N_81);
or U3094 (N_3094,N_719,N_1228);
or U3095 (N_3095,N_1631,N_1615);
and U3096 (N_3096,N_903,N_86);
or U3097 (N_3097,N_1716,N_1090);
and U3098 (N_3098,N_1779,N_45);
or U3099 (N_3099,N_1369,N_1649);
and U3100 (N_3100,N_314,N_355);
nor U3101 (N_3101,N_738,N_940);
nand U3102 (N_3102,N_1491,N_1022);
or U3103 (N_3103,N_1127,N_661);
or U3104 (N_3104,N_1384,N_407);
and U3105 (N_3105,N_1197,N_907);
nand U3106 (N_3106,N_121,N_728);
or U3107 (N_3107,N_1033,N_174);
nor U3108 (N_3108,N_345,N_1725);
nor U3109 (N_3109,N_400,N_1189);
nor U3110 (N_3110,N_1157,N_658);
and U3111 (N_3111,N_449,N_994);
or U3112 (N_3112,N_1130,N_1032);
nor U3113 (N_3113,N_3,N_641);
and U3114 (N_3114,N_1364,N_1550);
nor U3115 (N_3115,N_640,N_1485);
xor U3116 (N_3116,N_34,N_1699);
or U3117 (N_3117,N_798,N_870);
nand U3118 (N_3118,N_1480,N_1042);
nand U3119 (N_3119,N_358,N_267);
nor U3120 (N_3120,N_949,N_1276);
nor U3121 (N_3121,N_1100,N_1430);
nand U3122 (N_3122,N_1733,N_1226);
or U3123 (N_3123,N_499,N_177);
or U3124 (N_3124,N_56,N_1717);
nor U3125 (N_3125,N_412,N_1477);
and U3126 (N_3126,N_1356,N_876);
nand U3127 (N_3127,N_1803,N_132);
nor U3128 (N_3128,N_1529,N_1304);
or U3129 (N_3129,N_830,N_1789);
nor U3130 (N_3130,N_1592,N_1008);
or U3131 (N_3131,N_862,N_1163);
and U3132 (N_3132,N_1010,N_1114);
nand U3133 (N_3133,N_266,N_1669);
nand U3134 (N_3134,N_1244,N_229);
nand U3135 (N_3135,N_682,N_396);
or U3136 (N_3136,N_356,N_70);
and U3137 (N_3137,N_589,N_760);
or U3138 (N_3138,N_1132,N_1803);
nor U3139 (N_3139,N_1439,N_1680);
and U3140 (N_3140,N_1944,N_365);
nand U3141 (N_3141,N_1479,N_899);
nand U3142 (N_3142,N_1347,N_1512);
nand U3143 (N_3143,N_820,N_1220);
nand U3144 (N_3144,N_205,N_225);
and U3145 (N_3145,N_465,N_577);
nor U3146 (N_3146,N_1043,N_1202);
nand U3147 (N_3147,N_1008,N_260);
or U3148 (N_3148,N_813,N_1952);
or U3149 (N_3149,N_1143,N_638);
or U3150 (N_3150,N_1571,N_1707);
and U3151 (N_3151,N_1466,N_762);
nor U3152 (N_3152,N_1779,N_1189);
nand U3153 (N_3153,N_1960,N_861);
or U3154 (N_3154,N_1002,N_63);
or U3155 (N_3155,N_1180,N_1308);
and U3156 (N_3156,N_1703,N_324);
and U3157 (N_3157,N_692,N_890);
and U3158 (N_3158,N_542,N_1792);
or U3159 (N_3159,N_246,N_929);
and U3160 (N_3160,N_454,N_1904);
nor U3161 (N_3161,N_1153,N_1963);
or U3162 (N_3162,N_618,N_751);
and U3163 (N_3163,N_1710,N_1561);
nor U3164 (N_3164,N_1889,N_1925);
nor U3165 (N_3165,N_1511,N_1436);
or U3166 (N_3166,N_1495,N_610);
or U3167 (N_3167,N_906,N_1313);
and U3168 (N_3168,N_809,N_1971);
or U3169 (N_3169,N_466,N_1834);
nor U3170 (N_3170,N_1986,N_767);
and U3171 (N_3171,N_817,N_266);
or U3172 (N_3172,N_24,N_1545);
and U3173 (N_3173,N_511,N_1642);
nor U3174 (N_3174,N_1624,N_1665);
and U3175 (N_3175,N_602,N_1929);
nand U3176 (N_3176,N_1551,N_1856);
nand U3177 (N_3177,N_972,N_250);
nand U3178 (N_3178,N_310,N_53);
and U3179 (N_3179,N_935,N_558);
nand U3180 (N_3180,N_700,N_1512);
nor U3181 (N_3181,N_588,N_407);
nor U3182 (N_3182,N_774,N_1067);
nor U3183 (N_3183,N_732,N_1644);
or U3184 (N_3184,N_102,N_1783);
or U3185 (N_3185,N_1297,N_725);
xnor U3186 (N_3186,N_1100,N_1715);
or U3187 (N_3187,N_299,N_98);
nor U3188 (N_3188,N_1609,N_1379);
nor U3189 (N_3189,N_1210,N_23);
and U3190 (N_3190,N_985,N_776);
and U3191 (N_3191,N_20,N_784);
nor U3192 (N_3192,N_1625,N_1595);
nand U3193 (N_3193,N_1342,N_1798);
nand U3194 (N_3194,N_1573,N_1051);
nor U3195 (N_3195,N_378,N_1638);
nor U3196 (N_3196,N_60,N_367);
or U3197 (N_3197,N_551,N_826);
nand U3198 (N_3198,N_948,N_1218);
or U3199 (N_3199,N_1769,N_374);
or U3200 (N_3200,N_1512,N_1269);
nor U3201 (N_3201,N_1549,N_1639);
nand U3202 (N_3202,N_935,N_1659);
nand U3203 (N_3203,N_1277,N_1869);
nand U3204 (N_3204,N_749,N_1391);
xnor U3205 (N_3205,N_1103,N_1522);
nand U3206 (N_3206,N_812,N_1440);
or U3207 (N_3207,N_783,N_905);
xor U3208 (N_3208,N_513,N_1678);
nand U3209 (N_3209,N_303,N_16);
nor U3210 (N_3210,N_1445,N_1229);
or U3211 (N_3211,N_1332,N_1104);
nand U3212 (N_3212,N_312,N_1924);
xor U3213 (N_3213,N_921,N_885);
nor U3214 (N_3214,N_781,N_946);
or U3215 (N_3215,N_332,N_418);
or U3216 (N_3216,N_1359,N_234);
and U3217 (N_3217,N_1881,N_1534);
or U3218 (N_3218,N_1985,N_1475);
nor U3219 (N_3219,N_802,N_871);
nand U3220 (N_3220,N_501,N_1445);
nor U3221 (N_3221,N_652,N_1982);
or U3222 (N_3222,N_1970,N_1161);
nand U3223 (N_3223,N_1938,N_1987);
and U3224 (N_3224,N_374,N_1923);
nor U3225 (N_3225,N_537,N_760);
or U3226 (N_3226,N_676,N_1236);
nor U3227 (N_3227,N_628,N_1942);
and U3228 (N_3228,N_1787,N_472);
nand U3229 (N_3229,N_717,N_1074);
nand U3230 (N_3230,N_866,N_572);
or U3231 (N_3231,N_1514,N_818);
nor U3232 (N_3232,N_1496,N_1532);
and U3233 (N_3233,N_240,N_364);
nor U3234 (N_3234,N_737,N_608);
or U3235 (N_3235,N_937,N_1930);
nor U3236 (N_3236,N_934,N_861);
and U3237 (N_3237,N_40,N_1928);
and U3238 (N_3238,N_1339,N_297);
nand U3239 (N_3239,N_1446,N_267);
nand U3240 (N_3240,N_814,N_1540);
nor U3241 (N_3241,N_584,N_874);
and U3242 (N_3242,N_1673,N_275);
or U3243 (N_3243,N_295,N_1927);
nor U3244 (N_3244,N_1467,N_134);
and U3245 (N_3245,N_1859,N_144);
and U3246 (N_3246,N_1890,N_263);
nand U3247 (N_3247,N_1124,N_244);
or U3248 (N_3248,N_1702,N_1010);
or U3249 (N_3249,N_300,N_274);
nand U3250 (N_3250,N_207,N_1308);
nor U3251 (N_3251,N_1983,N_817);
nand U3252 (N_3252,N_939,N_404);
nor U3253 (N_3253,N_189,N_884);
nand U3254 (N_3254,N_808,N_1176);
or U3255 (N_3255,N_171,N_77);
nor U3256 (N_3256,N_627,N_759);
and U3257 (N_3257,N_1933,N_432);
nand U3258 (N_3258,N_1722,N_1658);
nor U3259 (N_3259,N_1648,N_121);
and U3260 (N_3260,N_1448,N_1518);
and U3261 (N_3261,N_1073,N_1397);
and U3262 (N_3262,N_59,N_502);
and U3263 (N_3263,N_1575,N_968);
xnor U3264 (N_3264,N_479,N_1791);
nand U3265 (N_3265,N_1971,N_1643);
nand U3266 (N_3266,N_1564,N_729);
nor U3267 (N_3267,N_1020,N_278);
nor U3268 (N_3268,N_404,N_1889);
or U3269 (N_3269,N_256,N_590);
or U3270 (N_3270,N_1728,N_1536);
or U3271 (N_3271,N_1347,N_894);
nor U3272 (N_3272,N_1984,N_1297);
nand U3273 (N_3273,N_817,N_531);
nand U3274 (N_3274,N_1367,N_925);
or U3275 (N_3275,N_969,N_1365);
nand U3276 (N_3276,N_1834,N_1332);
nand U3277 (N_3277,N_1492,N_66);
and U3278 (N_3278,N_553,N_1703);
and U3279 (N_3279,N_637,N_1214);
nand U3280 (N_3280,N_1922,N_260);
and U3281 (N_3281,N_1225,N_693);
nand U3282 (N_3282,N_106,N_1127);
or U3283 (N_3283,N_1327,N_615);
nand U3284 (N_3284,N_1331,N_1616);
and U3285 (N_3285,N_1177,N_153);
and U3286 (N_3286,N_301,N_92);
or U3287 (N_3287,N_959,N_523);
nand U3288 (N_3288,N_1507,N_388);
nor U3289 (N_3289,N_527,N_1858);
nand U3290 (N_3290,N_1968,N_1092);
and U3291 (N_3291,N_727,N_1869);
nor U3292 (N_3292,N_665,N_249);
or U3293 (N_3293,N_1653,N_1613);
and U3294 (N_3294,N_1413,N_730);
and U3295 (N_3295,N_193,N_435);
and U3296 (N_3296,N_484,N_962);
and U3297 (N_3297,N_325,N_1727);
or U3298 (N_3298,N_745,N_1221);
nor U3299 (N_3299,N_620,N_1947);
and U3300 (N_3300,N_859,N_1734);
nand U3301 (N_3301,N_1191,N_708);
or U3302 (N_3302,N_1948,N_1371);
and U3303 (N_3303,N_622,N_335);
nand U3304 (N_3304,N_88,N_159);
nand U3305 (N_3305,N_1411,N_1647);
or U3306 (N_3306,N_393,N_133);
and U3307 (N_3307,N_882,N_224);
nand U3308 (N_3308,N_1678,N_252);
and U3309 (N_3309,N_38,N_910);
nand U3310 (N_3310,N_717,N_1138);
and U3311 (N_3311,N_834,N_1783);
nor U3312 (N_3312,N_1888,N_1395);
and U3313 (N_3313,N_1041,N_399);
nand U3314 (N_3314,N_331,N_631);
nand U3315 (N_3315,N_1746,N_1214);
nor U3316 (N_3316,N_1462,N_501);
nor U3317 (N_3317,N_943,N_339);
nand U3318 (N_3318,N_163,N_547);
and U3319 (N_3319,N_1282,N_1969);
nor U3320 (N_3320,N_1067,N_1390);
or U3321 (N_3321,N_692,N_48);
nor U3322 (N_3322,N_1539,N_1649);
or U3323 (N_3323,N_197,N_515);
and U3324 (N_3324,N_549,N_981);
nor U3325 (N_3325,N_1478,N_221);
and U3326 (N_3326,N_788,N_222);
nor U3327 (N_3327,N_969,N_1254);
nand U3328 (N_3328,N_170,N_929);
or U3329 (N_3329,N_18,N_1666);
nand U3330 (N_3330,N_480,N_225);
nand U3331 (N_3331,N_580,N_466);
or U3332 (N_3332,N_1676,N_1203);
nand U3333 (N_3333,N_373,N_1494);
nor U3334 (N_3334,N_1815,N_862);
or U3335 (N_3335,N_734,N_181);
or U3336 (N_3336,N_637,N_742);
nor U3337 (N_3337,N_1429,N_1321);
nand U3338 (N_3338,N_1086,N_394);
nor U3339 (N_3339,N_1282,N_1994);
nand U3340 (N_3340,N_1186,N_292);
xnor U3341 (N_3341,N_1823,N_225);
and U3342 (N_3342,N_200,N_1023);
or U3343 (N_3343,N_1870,N_414);
nor U3344 (N_3344,N_341,N_808);
nand U3345 (N_3345,N_1448,N_168);
nor U3346 (N_3346,N_1134,N_715);
and U3347 (N_3347,N_644,N_1053);
nor U3348 (N_3348,N_146,N_785);
or U3349 (N_3349,N_1943,N_1897);
or U3350 (N_3350,N_1660,N_1913);
xor U3351 (N_3351,N_638,N_870);
and U3352 (N_3352,N_889,N_1416);
and U3353 (N_3353,N_1457,N_1250);
nand U3354 (N_3354,N_1149,N_677);
nand U3355 (N_3355,N_234,N_1814);
nand U3356 (N_3356,N_452,N_1358);
nor U3357 (N_3357,N_1673,N_658);
and U3358 (N_3358,N_1962,N_424);
or U3359 (N_3359,N_1957,N_516);
nor U3360 (N_3360,N_1122,N_1288);
or U3361 (N_3361,N_145,N_127);
and U3362 (N_3362,N_1798,N_1918);
nand U3363 (N_3363,N_1347,N_686);
and U3364 (N_3364,N_1148,N_1721);
and U3365 (N_3365,N_1640,N_279);
nor U3366 (N_3366,N_727,N_1836);
nor U3367 (N_3367,N_700,N_660);
or U3368 (N_3368,N_314,N_1522);
and U3369 (N_3369,N_1692,N_376);
nand U3370 (N_3370,N_1712,N_1066);
xnor U3371 (N_3371,N_324,N_158);
or U3372 (N_3372,N_447,N_458);
and U3373 (N_3373,N_1833,N_16);
and U3374 (N_3374,N_1530,N_373);
nand U3375 (N_3375,N_1835,N_67);
and U3376 (N_3376,N_750,N_1823);
nor U3377 (N_3377,N_907,N_549);
and U3378 (N_3378,N_664,N_600);
and U3379 (N_3379,N_23,N_463);
nand U3380 (N_3380,N_207,N_820);
or U3381 (N_3381,N_1342,N_302);
or U3382 (N_3382,N_1437,N_878);
and U3383 (N_3383,N_23,N_1293);
nor U3384 (N_3384,N_826,N_11);
nand U3385 (N_3385,N_1694,N_1550);
or U3386 (N_3386,N_1611,N_620);
or U3387 (N_3387,N_404,N_662);
nor U3388 (N_3388,N_1199,N_1534);
nor U3389 (N_3389,N_1208,N_1539);
or U3390 (N_3390,N_559,N_1791);
and U3391 (N_3391,N_785,N_1875);
or U3392 (N_3392,N_1764,N_983);
nor U3393 (N_3393,N_909,N_132);
and U3394 (N_3394,N_953,N_451);
nor U3395 (N_3395,N_1053,N_1265);
nand U3396 (N_3396,N_743,N_827);
nor U3397 (N_3397,N_238,N_1755);
nand U3398 (N_3398,N_635,N_1277);
nor U3399 (N_3399,N_1935,N_1689);
nor U3400 (N_3400,N_524,N_770);
nor U3401 (N_3401,N_1684,N_93);
nand U3402 (N_3402,N_84,N_583);
nor U3403 (N_3403,N_1424,N_700);
or U3404 (N_3404,N_261,N_1431);
nand U3405 (N_3405,N_1816,N_1638);
and U3406 (N_3406,N_1762,N_1098);
or U3407 (N_3407,N_167,N_53);
and U3408 (N_3408,N_1102,N_1950);
nor U3409 (N_3409,N_1211,N_1225);
and U3410 (N_3410,N_156,N_1213);
nor U3411 (N_3411,N_1315,N_398);
and U3412 (N_3412,N_335,N_1024);
or U3413 (N_3413,N_797,N_1737);
and U3414 (N_3414,N_249,N_1368);
nor U3415 (N_3415,N_1786,N_575);
nor U3416 (N_3416,N_922,N_1860);
nand U3417 (N_3417,N_1221,N_110);
xnor U3418 (N_3418,N_1637,N_782);
or U3419 (N_3419,N_1579,N_941);
nor U3420 (N_3420,N_1060,N_993);
or U3421 (N_3421,N_590,N_1019);
and U3422 (N_3422,N_375,N_426);
or U3423 (N_3423,N_651,N_680);
nor U3424 (N_3424,N_559,N_1079);
and U3425 (N_3425,N_1766,N_859);
nor U3426 (N_3426,N_1971,N_906);
and U3427 (N_3427,N_130,N_459);
nor U3428 (N_3428,N_957,N_193);
and U3429 (N_3429,N_1220,N_884);
nor U3430 (N_3430,N_333,N_1263);
and U3431 (N_3431,N_100,N_219);
nand U3432 (N_3432,N_114,N_1635);
nand U3433 (N_3433,N_352,N_1360);
or U3434 (N_3434,N_748,N_1571);
nor U3435 (N_3435,N_478,N_1786);
and U3436 (N_3436,N_1841,N_1685);
or U3437 (N_3437,N_1865,N_1765);
nand U3438 (N_3438,N_773,N_1457);
and U3439 (N_3439,N_520,N_1174);
nand U3440 (N_3440,N_1153,N_233);
or U3441 (N_3441,N_2,N_1318);
nand U3442 (N_3442,N_151,N_1822);
or U3443 (N_3443,N_1449,N_756);
nor U3444 (N_3444,N_1461,N_1232);
and U3445 (N_3445,N_865,N_1237);
xor U3446 (N_3446,N_1094,N_1766);
nor U3447 (N_3447,N_310,N_1911);
nor U3448 (N_3448,N_1395,N_489);
and U3449 (N_3449,N_1837,N_170);
nand U3450 (N_3450,N_1440,N_845);
and U3451 (N_3451,N_1420,N_1632);
or U3452 (N_3452,N_898,N_600);
nand U3453 (N_3453,N_536,N_272);
or U3454 (N_3454,N_1334,N_239);
and U3455 (N_3455,N_1707,N_1435);
or U3456 (N_3456,N_1855,N_411);
nor U3457 (N_3457,N_5,N_1669);
nor U3458 (N_3458,N_1441,N_1681);
and U3459 (N_3459,N_528,N_521);
or U3460 (N_3460,N_45,N_1085);
nand U3461 (N_3461,N_1368,N_1655);
nand U3462 (N_3462,N_1316,N_1098);
or U3463 (N_3463,N_1605,N_1630);
nor U3464 (N_3464,N_1550,N_1267);
or U3465 (N_3465,N_976,N_1537);
nor U3466 (N_3466,N_1816,N_1643);
nand U3467 (N_3467,N_327,N_1904);
and U3468 (N_3468,N_1501,N_802);
or U3469 (N_3469,N_1970,N_589);
nand U3470 (N_3470,N_1718,N_1146);
nor U3471 (N_3471,N_508,N_1271);
nor U3472 (N_3472,N_1855,N_1922);
nand U3473 (N_3473,N_867,N_987);
and U3474 (N_3474,N_310,N_1734);
nor U3475 (N_3475,N_101,N_1944);
nor U3476 (N_3476,N_231,N_375);
nand U3477 (N_3477,N_1363,N_91);
or U3478 (N_3478,N_1158,N_1105);
nor U3479 (N_3479,N_1920,N_1813);
nand U3480 (N_3480,N_20,N_555);
nand U3481 (N_3481,N_1616,N_906);
and U3482 (N_3482,N_1994,N_1763);
or U3483 (N_3483,N_333,N_1192);
or U3484 (N_3484,N_335,N_1658);
or U3485 (N_3485,N_597,N_838);
nor U3486 (N_3486,N_392,N_1607);
or U3487 (N_3487,N_1378,N_590);
nor U3488 (N_3488,N_97,N_513);
xor U3489 (N_3489,N_151,N_1324);
nand U3490 (N_3490,N_1475,N_185);
and U3491 (N_3491,N_1957,N_1677);
and U3492 (N_3492,N_1111,N_1532);
xor U3493 (N_3493,N_52,N_477);
nor U3494 (N_3494,N_710,N_1167);
nor U3495 (N_3495,N_1495,N_827);
and U3496 (N_3496,N_1736,N_67);
or U3497 (N_3497,N_948,N_1678);
and U3498 (N_3498,N_1794,N_513);
nor U3499 (N_3499,N_1568,N_1575);
nor U3500 (N_3500,N_1797,N_1992);
nand U3501 (N_3501,N_1140,N_1545);
and U3502 (N_3502,N_949,N_1037);
nand U3503 (N_3503,N_1143,N_1584);
nor U3504 (N_3504,N_784,N_778);
nor U3505 (N_3505,N_1857,N_873);
nor U3506 (N_3506,N_1058,N_463);
and U3507 (N_3507,N_125,N_739);
xor U3508 (N_3508,N_983,N_1094);
nor U3509 (N_3509,N_981,N_212);
nor U3510 (N_3510,N_1530,N_1787);
and U3511 (N_3511,N_1582,N_981);
nand U3512 (N_3512,N_1988,N_1518);
nor U3513 (N_3513,N_886,N_518);
nand U3514 (N_3514,N_688,N_817);
or U3515 (N_3515,N_463,N_114);
xnor U3516 (N_3516,N_879,N_1312);
and U3517 (N_3517,N_231,N_964);
nor U3518 (N_3518,N_1388,N_409);
nand U3519 (N_3519,N_335,N_1010);
nor U3520 (N_3520,N_1430,N_254);
or U3521 (N_3521,N_1911,N_1658);
or U3522 (N_3522,N_155,N_257);
or U3523 (N_3523,N_614,N_846);
and U3524 (N_3524,N_136,N_118);
or U3525 (N_3525,N_583,N_869);
nand U3526 (N_3526,N_1711,N_622);
and U3527 (N_3527,N_829,N_1878);
nor U3528 (N_3528,N_1387,N_1615);
nand U3529 (N_3529,N_1575,N_785);
or U3530 (N_3530,N_390,N_1405);
nand U3531 (N_3531,N_1952,N_1514);
and U3532 (N_3532,N_873,N_683);
nor U3533 (N_3533,N_1552,N_1844);
or U3534 (N_3534,N_1019,N_1173);
or U3535 (N_3535,N_1528,N_855);
xnor U3536 (N_3536,N_400,N_329);
xor U3537 (N_3537,N_794,N_429);
xor U3538 (N_3538,N_625,N_1051);
nand U3539 (N_3539,N_410,N_598);
nor U3540 (N_3540,N_621,N_1273);
or U3541 (N_3541,N_1932,N_1533);
nor U3542 (N_3542,N_1510,N_1367);
nor U3543 (N_3543,N_1214,N_512);
nor U3544 (N_3544,N_688,N_591);
or U3545 (N_3545,N_1840,N_1877);
and U3546 (N_3546,N_1801,N_359);
or U3547 (N_3547,N_1106,N_1029);
or U3548 (N_3548,N_1406,N_1286);
or U3549 (N_3549,N_617,N_1187);
or U3550 (N_3550,N_1777,N_1447);
and U3551 (N_3551,N_1813,N_907);
nand U3552 (N_3552,N_400,N_1105);
nand U3553 (N_3553,N_1225,N_1088);
nand U3554 (N_3554,N_717,N_1360);
and U3555 (N_3555,N_612,N_1683);
nand U3556 (N_3556,N_192,N_245);
nand U3557 (N_3557,N_1413,N_1320);
and U3558 (N_3558,N_212,N_790);
nand U3559 (N_3559,N_1475,N_574);
or U3560 (N_3560,N_207,N_1847);
or U3561 (N_3561,N_1899,N_566);
and U3562 (N_3562,N_1398,N_57);
nor U3563 (N_3563,N_21,N_1396);
nand U3564 (N_3564,N_1834,N_285);
or U3565 (N_3565,N_131,N_1543);
xnor U3566 (N_3566,N_1273,N_580);
xnor U3567 (N_3567,N_1199,N_736);
nor U3568 (N_3568,N_1405,N_724);
or U3569 (N_3569,N_1951,N_676);
or U3570 (N_3570,N_1020,N_190);
nor U3571 (N_3571,N_1190,N_1469);
nor U3572 (N_3572,N_1279,N_1255);
or U3573 (N_3573,N_1525,N_1162);
nor U3574 (N_3574,N_1024,N_408);
and U3575 (N_3575,N_1482,N_24);
or U3576 (N_3576,N_1111,N_873);
and U3577 (N_3577,N_100,N_1591);
nor U3578 (N_3578,N_920,N_1887);
nor U3579 (N_3579,N_1803,N_1579);
nor U3580 (N_3580,N_1598,N_40);
nand U3581 (N_3581,N_1611,N_1014);
and U3582 (N_3582,N_1439,N_678);
or U3583 (N_3583,N_1359,N_849);
nand U3584 (N_3584,N_1038,N_912);
xnor U3585 (N_3585,N_159,N_1484);
and U3586 (N_3586,N_1788,N_915);
or U3587 (N_3587,N_1318,N_70);
nor U3588 (N_3588,N_1768,N_282);
nor U3589 (N_3589,N_508,N_203);
nor U3590 (N_3590,N_892,N_788);
nand U3591 (N_3591,N_1287,N_1339);
nor U3592 (N_3592,N_1761,N_25);
nand U3593 (N_3593,N_980,N_1804);
or U3594 (N_3594,N_270,N_597);
or U3595 (N_3595,N_1171,N_770);
nand U3596 (N_3596,N_1311,N_545);
nand U3597 (N_3597,N_71,N_252);
nor U3598 (N_3598,N_1372,N_1819);
or U3599 (N_3599,N_552,N_1223);
or U3600 (N_3600,N_932,N_532);
and U3601 (N_3601,N_30,N_113);
or U3602 (N_3602,N_479,N_535);
nand U3603 (N_3603,N_1578,N_1939);
nor U3604 (N_3604,N_1297,N_531);
and U3605 (N_3605,N_702,N_933);
nand U3606 (N_3606,N_1113,N_712);
nor U3607 (N_3607,N_1498,N_1060);
or U3608 (N_3608,N_82,N_818);
and U3609 (N_3609,N_1818,N_828);
nor U3610 (N_3610,N_1978,N_214);
nor U3611 (N_3611,N_1903,N_1347);
nor U3612 (N_3612,N_1223,N_803);
and U3613 (N_3613,N_75,N_1784);
nand U3614 (N_3614,N_620,N_1575);
or U3615 (N_3615,N_1786,N_1026);
and U3616 (N_3616,N_1177,N_58);
or U3617 (N_3617,N_795,N_1997);
nand U3618 (N_3618,N_1858,N_949);
nor U3619 (N_3619,N_263,N_366);
and U3620 (N_3620,N_1222,N_1558);
and U3621 (N_3621,N_1485,N_50);
nor U3622 (N_3622,N_331,N_1326);
and U3623 (N_3623,N_1038,N_1116);
and U3624 (N_3624,N_386,N_988);
nand U3625 (N_3625,N_12,N_11);
or U3626 (N_3626,N_1647,N_218);
and U3627 (N_3627,N_1927,N_1206);
and U3628 (N_3628,N_1411,N_230);
or U3629 (N_3629,N_1174,N_197);
nand U3630 (N_3630,N_1818,N_1655);
and U3631 (N_3631,N_674,N_1175);
xor U3632 (N_3632,N_1196,N_1109);
and U3633 (N_3633,N_1358,N_1414);
and U3634 (N_3634,N_783,N_1473);
nand U3635 (N_3635,N_1706,N_442);
nand U3636 (N_3636,N_779,N_764);
or U3637 (N_3637,N_877,N_1236);
nand U3638 (N_3638,N_347,N_1909);
and U3639 (N_3639,N_1367,N_1587);
nor U3640 (N_3640,N_548,N_641);
nand U3641 (N_3641,N_82,N_986);
nand U3642 (N_3642,N_1161,N_1195);
nand U3643 (N_3643,N_1640,N_420);
or U3644 (N_3644,N_173,N_1780);
nor U3645 (N_3645,N_1950,N_1166);
nor U3646 (N_3646,N_858,N_610);
nand U3647 (N_3647,N_503,N_1421);
xor U3648 (N_3648,N_1683,N_497);
nand U3649 (N_3649,N_1848,N_1320);
or U3650 (N_3650,N_114,N_1877);
nor U3651 (N_3651,N_1044,N_1407);
nor U3652 (N_3652,N_949,N_389);
nor U3653 (N_3653,N_9,N_1793);
or U3654 (N_3654,N_1076,N_1962);
nand U3655 (N_3655,N_628,N_631);
nand U3656 (N_3656,N_854,N_1195);
nor U3657 (N_3657,N_1126,N_1307);
and U3658 (N_3658,N_1056,N_538);
nand U3659 (N_3659,N_1531,N_697);
or U3660 (N_3660,N_780,N_1376);
or U3661 (N_3661,N_1813,N_1387);
and U3662 (N_3662,N_1856,N_1479);
and U3663 (N_3663,N_1421,N_1246);
nor U3664 (N_3664,N_862,N_1530);
and U3665 (N_3665,N_1049,N_1150);
and U3666 (N_3666,N_1093,N_112);
nor U3667 (N_3667,N_1683,N_215);
nor U3668 (N_3668,N_722,N_1760);
xnor U3669 (N_3669,N_719,N_71);
or U3670 (N_3670,N_168,N_735);
or U3671 (N_3671,N_1296,N_1760);
nand U3672 (N_3672,N_1568,N_1861);
nor U3673 (N_3673,N_1059,N_983);
and U3674 (N_3674,N_1767,N_741);
or U3675 (N_3675,N_194,N_1413);
and U3676 (N_3676,N_773,N_1364);
nand U3677 (N_3677,N_1955,N_1222);
and U3678 (N_3678,N_610,N_1470);
nand U3679 (N_3679,N_655,N_220);
nor U3680 (N_3680,N_1536,N_782);
nand U3681 (N_3681,N_1650,N_744);
or U3682 (N_3682,N_810,N_749);
nand U3683 (N_3683,N_403,N_184);
and U3684 (N_3684,N_1324,N_1896);
nand U3685 (N_3685,N_1763,N_616);
and U3686 (N_3686,N_1870,N_1353);
and U3687 (N_3687,N_61,N_88);
nor U3688 (N_3688,N_365,N_1873);
and U3689 (N_3689,N_191,N_1236);
nand U3690 (N_3690,N_681,N_1296);
nor U3691 (N_3691,N_1982,N_1658);
and U3692 (N_3692,N_671,N_1299);
nor U3693 (N_3693,N_302,N_1798);
nand U3694 (N_3694,N_787,N_196);
or U3695 (N_3695,N_1278,N_1255);
and U3696 (N_3696,N_1319,N_812);
nor U3697 (N_3697,N_368,N_1134);
or U3698 (N_3698,N_1985,N_265);
and U3699 (N_3699,N_150,N_1644);
nand U3700 (N_3700,N_678,N_1729);
nor U3701 (N_3701,N_1848,N_3);
nor U3702 (N_3702,N_417,N_1475);
nand U3703 (N_3703,N_1228,N_1001);
and U3704 (N_3704,N_1762,N_1304);
or U3705 (N_3705,N_851,N_89);
and U3706 (N_3706,N_617,N_1682);
nor U3707 (N_3707,N_1658,N_1772);
and U3708 (N_3708,N_889,N_272);
nand U3709 (N_3709,N_161,N_1450);
and U3710 (N_3710,N_1178,N_1200);
nor U3711 (N_3711,N_1078,N_762);
nor U3712 (N_3712,N_1147,N_1771);
and U3713 (N_3713,N_833,N_89);
and U3714 (N_3714,N_1309,N_1585);
or U3715 (N_3715,N_14,N_1682);
nand U3716 (N_3716,N_1938,N_1245);
or U3717 (N_3717,N_1412,N_296);
nor U3718 (N_3718,N_798,N_10);
and U3719 (N_3719,N_639,N_1309);
or U3720 (N_3720,N_631,N_1620);
nand U3721 (N_3721,N_709,N_1761);
or U3722 (N_3722,N_247,N_1931);
and U3723 (N_3723,N_325,N_1979);
or U3724 (N_3724,N_227,N_1310);
nand U3725 (N_3725,N_461,N_1351);
nand U3726 (N_3726,N_694,N_1267);
nor U3727 (N_3727,N_1216,N_1167);
nand U3728 (N_3728,N_963,N_362);
or U3729 (N_3729,N_49,N_1842);
or U3730 (N_3730,N_371,N_993);
nor U3731 (N_3731,N_1090,N_825);
or U3732 (N_3732,N_1994,N_417);
and U3733 (N_3733,N_694,N_360);
and U3734 (N_3734,N_1156,N_451);
nand U3735 (N_3735,N_1503,N_271);
nor U3736 (N_3736,N_1171,N_634);
nand U3737 (N_3737,N_1550,N_1371);
and U3738 (N_3738,N_1376,N_953);
and U3739 (N_3739,N_52,N_1845);
or U3740 (N_3740,N_1370,N_633);
or U3741 (N_3741,N_1040,N_627);
and U3742 (N_3742,N_706,N_287);
or U3743 (N_3743,N_1510,N_222);
and U3744 (N_3744,N_1249,N_1663);
nand U3745 (N_3745,N_934,N_1869);
nand U3746 (N_3746,N_807,N_1351);
nand U3747 (N_3747,N_333,N_1953);
and U3748 (N_3748,N_1277,N_346);
nor U3749 (N_3749,N_251,N_204);
xnor U3750 (N_3750,N_741,N_1642);
nand U3751 (N_3751,N_717,N_1573);
or U3752 (N_3752,N_330,N_1323);
nand U3753 (N_3753,N_1534,N_67);
nand U3754 (N_3754,N_1132,N_1071);
nand U3755 (N_3755,N_1508,N_828);
and U3756 (N_3756,N_409,N_1150);
and U3757 (N_3757,N_3,N_491);
and U3758 (N_3758,N_993,N_1774);
or U3759 (N_3759,N_1243,N_890);
nor U3760 (N_3760,N_1416,N_1991);
xnor U3761 (N_3761,N_1444,N_673);
or U3762 (N_3762,N_1116,N_1950);
nor U3763 (N_3763,N_730,N_1777);
and U3764 (N_3764,N_741,N_1507);
nand U3765 (N_3765,N_399,N_309);
or U3766 (N_3766,N_1623,N_518);
or U3767 (N_3767,N_976,N_318);
and U3768 (N_3768,N_1615,N_826);
or U3769 (N_3769,N_1119,N_1187);
nor U3770 (N_3770,N_1174,N_675);
nor U3771 (N_3771,N_1028,N_1565);
and U3772 (N_3772,N_278,N_155);
or U3773 (N_3773,N_331,N_249);
nor U3774 (N_3774,N_1454,N_1322);
and U3775 (N_3775,N_267,N_977);
nor U3776 (N_3776,N_1290,N_771);
and U3777 (N_3777,N_1288,N_884);
and U3778 (N_3778,N_1211,N_982);
nor U3779 (N_3779,N_1652,N_301);
nand U3780 (N_3780,N_624,N_1847);
nor U3781 (N_3781,N_911,N_1452);
and U3782 (N_3782,N_1302,N_1784);
nor U3783 (N_3783,N_1092,N_707);
nand U3784 (N_3784,N_244,N_882);
and U3785 (N_3785,N_1533,N_4);
nor U3786 (N_3786,N_713,N_1600);
and U3787 (N_3787,N_1012,N_1526);
and U3788 (N_3788,N_954,N_1811);
nand U3789 (N_3789,N_1488,N_1861);
nand U3790 (N_3790,N_1915,N_816);
or U3791 (N_3791,N_1124,N_1025);
and U3792 (N_3792,N_301,N_1853);
and U3793 (N_3793,N_1384,N_1675);
and U3794 (N_3794,N_1942,N_410);
nor U3795 (N_3795,N_1371,N_445);
nor U3796 (N_3796,N_1216,N_7);
nand U3797 (N_3797,N_12,N_1696);
nor U3798 (N_3798,N_263,N_689);
nand U3799 (N_3799,N_1017,N_450);
xnor U3800 (N_3800,N_1661,N_1036);
nor U3801 (N_3801,N_914,N_908);
or U3802 (N_3802,N_1895,N_572);
nor U3803 (N_3803,N_413,N_1646);
or U3804 (N_3804,N_1031,N_280);
nand U3805 (N_3805,N_1395,N_970);
or U3806 (N_3806,N_237,N_1200);
nor U3807 (N_3807,N_856,N_1634);
or U3808 (N_3808,N_10,N_1570);
and U3809 (N_3809,N_1101,N_1952);
or U3810 (N_3810,N_1973,N_1411);
and U3811 (N_3811,N_1096,N_1134);
and U3812 (N_3812,N_608,N_174);
or U3813 (N_3813,N_1389,N_1477);
nor U3814 (N_3814,N_22,N_1606);
nor U3815 (N_3815,N_1088,N_150);
or U3816 (N_3816,N_945,N_353);
nor U3817 (N_3817,N_1015,N_1305);
or U3818 (N_3818,N_1892,N_1904);
and U3819 (N_3819,N_491,N_196);
or U3820 (N_3820,N_1922,N_423);
nor U3821 (N_3821,N_1766,N_1884);
nor U3822 (N_3822,N_1768,N_1842);
xnor U3823 (N_3823,N_1113,N_1967);
nor U3824 (N_3824,N_1289,N_1185);
nor U3825 (N_3825,N_811,N_1070);
nor U3826 (N_3826,N_1640,N_430);
and U3827 (N_3827,N_1307,N_1412);
nor U3828 (N_3828,N_1587,N_1774);
nor U3829 (N_3829,N_577,N_1951);
nand U3830 (N_3830,N_1114,N_575);
or U3831 (N_3831,N_27,N_1079);
nand U3832 (N_3832,N_689,N_794);
nor U3833 (N_3833,N_1146,N_259);
or U3834 (N_3834,N_549,N_1244);
or U3835 (N_3835,N_1536,N_171);
or U3836 (N_3836,N_12,N_697);
nor U3837 (N_3837,N_725,N_979);
or U3838 (N_3838,N_1610,N_1567);
and U3839 (N_3839,N_901,N_1924);
and U3840 (N_3840,N_1078,N_1696);
nand U3841 (N_3841,N_1347,N_780);
nand U3842 (N_3842,N_1092,N_1205);
and U3843 (N_3843,N_1852,N_1902);
nand U3844 (N_3844,N_802,N_912);
nand U3845 (N_3845,N_1428,N_1276);
nor U3846 (N_3846,N_925,N_1935);
nor U3847 (N_3847,N_742,N_1543);
nand U3848 (N_3848,N_166,N_1762);
or U3849 (N_3849,N_374,N_1379);
nand U3850 (N_3850,N_1020,N_625);
nand U3851 (N_3851,N_1409,N_1776);
and U3852 (N_3852,N_1032,N_241);
nand U3853 (N_3853,N_1983,N_1010);
and U3854 (N_3854,N_1711,N_1752);
or U3855 (N_3855,N_4,N_791);
nor U3856 (N_3856,N_1167,N_967);
and U3857 (N_3857,N_1544,N_378);
nand U3858 (N_3858,N_462,N_1150);
nand U3859 (N_3859,N_1160,N_910);
nand U3860 (N_3860,N_1057,N_404);
nand U3861 (N_3861,N_1815,N_168);
or U3862 (N_3862,N_1035,N_1973);
nor U3863 (N_3863,N_213,N_1157);
nand U3864 (N_3864,N_1046,N_1075);
nand U3865 (N_3865,N_1277,N_967);
nand U3866 (N_3866,N_1563,N_1591);
or U3867 (N_3867,N_1256,N_1951);
and U3868 (N_3868,N_263,N_830);
nor U3869 (N_3869,N_46,N_227);
nor U3870 (N_3870,N_711,N_1025);
and U3871 (N_3871,N_1696,N_416);
nand U3872 (N_3872,N_975,N_354);
or U3873 (N_3873,N_1610,N_1864);
nand U3874 (N_3874,N_1741,N_682);
or U3875 (N_3875,N_1708,N_1850);
nand U3876 (N_3876,N_1679,N_850);
and U3877 (N_3877,N_1742,N_702);
nor U3878 (N_3878,N_1588,N_1873);
nand U3879 (N_3879,N_1100,N_1405);
nand U3880 (N_3880,N_1987,N_344);
nor U3881 (N_3881,N_874,N_754);
nor U3882 (N_3882,N_1926,N_1513);
nor U3883 (N_3883,N_1871,N_377);
nor U3884 (N_3884,N_817,N_1730);
nor U3885 (N_3885,N_999,N_649);
xnor U3886 (N_3886,N_1745,N_1468);
nor U3887 (N_3887,N_1139,N_1316);
or U3888 (N_3888,N_398,N_658);
nor U3889 (N_3889,N_1560,N_1153);
or U3890 (N_3890,N_1089,N_559);
nor U3891 (N_3891,N_441,N_1298);
nor U3892 (N_3892,N_1735,N_473);
or U3893 (N_3893,N_470,N_1124);
nor U3894 (N_3894,N_740,N_30);
nor U3895 (N_3895,N_462,N_899);
and U3896 (N_3896,N_1678,N_863);
or U3897 (N_3897,N_1994,N_1413);
nand U3898 (N_3898,N_335,N_955);
nor U3899 (N_3899,N_666,N_784);
xnor U3900 (N_3900,N_1347,N_1511);
nor U3901 (N_3901,N_595,N_938);
nand U3902 (N_3902,N_422,N_1130);
xnor U3903 (N_3903,N_886,N_119);
nor U3904 (N_3904,N_666,N_1666);
nor U3905 (N_3905,N_407,N_1294);
or U3906 (N_3906,N_1280,N_1297);
and U3907 (N_3907,N_774,N_130);
nand U3908 (N_3908,N_1341,N_1758);
or U3909 (N_3909,N_1569,N_1349);
nor U3910 (N_3910,N_62,N_420);
nand U3911 (N_3911,N_1096,N_1408);
and U3912 (N_3912,N_1394,N_1571);
nor U3913 (N_3913,N_1503,N_1304);
nor U3914 (N_3914,N_225,N_565);
nand U3915 (N_3915,N_1488,N_1284);
nor U3916 (N_3916,N_76,N_1655);
or U3917 (N_3917,N_215,N_1507);
or U3918 (N_3918,N_859,N_36);
and U3919 (N_3919,N_818,N_496);
and U3920 (N_3920,N_1483,N_1140);
nor U3921 (N_3921,N_1050,N_609);
nand U3922 (N_3922,N_536,N_375);
xnor U3923 (N_3923,N_762,N_776);
and U3924 (N_3924,N_1228,N_94);
nor U3925 (N_3925,N_1025,N_3);
nand U3926 (N_3926,N_689,N_1315);
nand U3927 (N_3927,N_1780,N_1127);
and U3928 (N_3928,N_1028,N_1364);
nand U3929 (N_3929,N_1970,N_211);
nand U3930 (N_3930,N_1090,N_961);
or U3931 (N_3931,N_737,N_1951);
and U3932 (N_3932,N_1625,N_968);
nand U3933 (N_3933,N_104,N_1935);
nor U3934 (N_3934,N_438,N_1979);
nor U3935 (N_3935,N_646,N_1809);
nand U3936 (N_3936,N_316,N_672);
and U3937 (N_3937,N_618,N_1892);
or U3938 (N_3938,N_980,N_1413);
and U3939 (N_3939,N_602,N_1380);
nor U3940 (N_3940,N_1313,N_1595);
nand U3941 (N_3941,N_1276,N_1193);
and U3942 (N_3942,N_1332,N_113);
or U3943 (N_3943,N_961,N_1967);
and U3944 (N_3944,N_1403,N_1918);
or U3945 (N_3945,N_226,N_443);
nand U3946 (N_3946,N_1420,N_992);
nand U3947 (N_3947,N_1685,N_1484);
nor U3948 (N_3948,N_1373,N_1416);
or U3949 (N_3949,N_358,N_1321);
or U3950 (N_3950,N_1808,N_1244);
or U3951 (N_3951,N_1725,N_1808);
or U3952 (N_3952,N_1794,N_1962);
and U3953 (N_3953,N_22,N_395);
and U3954 (N_3954,N_10,N_732);
and U3955 (N_3955,N_979,N_1189);
nand U3956 (N_3956,N_225,N_1485);
and U3957 (N_3957,N_1789,N_1548);
nand U3958 (N_3958,N_254,N_1928);
nand U3959 (N_3959,N_914,N_728);
xnor U3960 (N_3960,N_1878,N_534);
nand U3961 (N_3961,N_329,N_167);
and U3962 (N_3962,N_1236,N_1470);
or U3963 (N_3963,N_211,N_1683);
and U3964 (N_3964,N_1033,N_233);
or U3965 (N_3965,N_1841,N_1775);
nand U3966 (N_3966,N_1188,N_1651);
and U3967 (N_3967,N_1369,N_1889);
or U3968 (N_3968,N_1762,N_572);
or U3969 (N_3969,N_1457,N_1128);
and U3970 (N_3970,N_575,N_12);
or U3971 (N_3971,N_595,N_993);
xor U3972 (N_3972,N_1219,N_1289);
or U3973 (N_3973,N_1884,N_45);
nand U3974 (N_3974,N_1510,N_1555);
nand U3975 (N_3975,N_433,N_931);
and U3976 (N_3976,N_1751,N_1680);
and U3977 (N_3977,N_820,N_518);
and U3978 (N_3978,N_1382,N_880);
nand U3979 (N_3979,N_1350,N_648);
nor U3980 (N_3980,N_1949,N_781);
or U3981 (N_3981,N_209,N_1516);
nor U3982 (N_3982,N_1193,N_1419);
and U3983 (N_3983,N_1705,N_561);
or U3984 (N_3984,N_834,N_688);
or U3985 (N_3985,N_1457,N_143);
xnor U3986 (N_3986,N_1852,N_878);
nand U3987 (N_3987,N_712,N_1678);
xnor U3988 (N_3988,N_872,N_927);
or U3989 (N_3989,N_1783,N_289);
nand U3990 (N_3990,N_442,N_433);
or U3991 (N_3991,N_229,N_2);
nor U3992 (N_3992,N_626,N_1044);
or U3993 (N_3993,N_34,N_588);
nand U3994 (N_3994,N_512,N_237);
nand U3995 (N_3995,N_1444,N_1763);
nand U3996 (N_3996,N_35,N_1981);
and U3997 (N_3997,N_1015,N_923);
or U3998 (N_3998,N_747,N_587);
and U3999 (N_3999,N_1745,N_625);
nand U4000 (N_4000,N_3632,N_2189);
or U4001 (N_4001,N_2404,N_2341);
or U4002 (N_4002,N_2610,N_2432);
and U4003 (N_4003,N_2310,N_2063);
nand U4004 (N_4004,N_2410,N_2913);
nor U4005 (N_4005,N_3672,N_2200);
and U4006 (N_4006,N_2338,N_2125);
nor U4007 (N_4007,N_3739,N_2226);
and U4008 (N_4008,N_2465,N_2412);
and U4009 (N_4009,N_3494,N_3357);
nand U4010 (N_4010,N_3190,N_2786);
or U4011 (N_4011,N_2113,N_3653);
nor U4012 (N_4012,N_2866,N_2037);
xor U4013 (N_4013,N_3413,N_2122);
and U4014 (N_4014,N_3451,N_2936);
or U4015 (N_4015,N_3279,N_2130);
or U4016 (N_4016,N_3216,N_2639);
or U4017 (N_4017,N_2058,N_3024);
nand U4018 (N_4018,N_3970,N_3060);
nor U4019 (N_4019,N_3404,N_3186);
nor U4020 (N_4020,N_2585,N_3601);
nor U4021 (N_4021,N_2179,N_3348);
or U4022 (N_4022,N_3550,N_3432);
or U4023 (N_4023,N_2419,N_3806);
nor U4024 (N_4024,N_3500,N_3296);
nor U4025 (N_4025,N_2114,N_3517);
nor U4026 (N_4026,N_3000,N_3016);
xor U4027 (N_4027,N_2761,N_3912);
nand U4028 (N_4028,N_2031,N_2408);
or U4029 (N_4029,N_3893,N_2323);
or U4030 (N_4030,N_2388,N_3396);
and U4031 (N_4031,N_2135,N_2060);
and U4032 (N_4032,N_3213,N_3159);
nor U4033 (N_4033,N_2477,N_2378);
and U4034 (N_4034,N_2915,N_3239);
or U4035 (N_4035,N_3709,N_2912);
nand U4036 (N_4036,N_2846,N_3525);
or U4037 (N_4037,N_3485,N_3052);
or U4038 (N_4038,N_3483,N_2269);
and U4039 (N_4039,N_2097,N_2690);
or U4040 (N_4040,N_3128,N_2844);
nand U4041 (N_4041,N_2084,N_3565);
nand U4042 (N_4042,N_2005,N_2677);
nor U4043 (N_4043,N_2997,N_2329);
or U4044 (N_4044,N_2923,N_2293);
nor U4045 (N_4045,N_3789,N_2029);
and U4046 (N_4046,N_2916,N_3229);
or U4047 (N_4047,N_3725,N_3753);
or U4048 (N_4048,N_3926,N_2445);
or U4049 (N_4049,N_3945,N_3959);
and U4050 (N_4050,N_3620,N_2056);
nor U4051 (N_4051,N_3956,N_3014);
or U4052 (N_4052,N_3009,N_2235);
and U4053 (N_4053,N_3965,N_2655);
and U4054 (N_4054,N_2612,N_2175);
nor U4055 (N_4055,N_3030,N_2316);
nand U4056 (N_4056,N_3683,N_3978);
nand U4057 (N_4057,N_2115,N_2149);
or U4058 (N_4058,N_3145,N_3054);
nand U4059 (N_4059,N_2103,N_3252);
nand U4060 (N_4060,N_3933,N_3176);
and U4061 (N_4061,N_3658,N_3953);
nor U4062 (N_4062,N_2586,N_2036);
and U4063 (N_4063,N_2145,N_2631);
nand U4064 (N_4064,N_2163,N_3749);
or U4065 (N_4065,N_2238,N_2570);
or U4066 (N_4066,N_2210,N_2271);
nand U4067 (N_4067,N_3822,N_2253);
nor U4068 (N_4068,N_3082,N_2955);
and U4069 (N_4069,N_3745,N_3392);
nor U4070 (N_4070,N_3985,N_3942);
and U4071 (N_4071,N_3811,N_2721);
or U4072 (N_4072,N_2061,N_2298);
nand U4073 (N_4073,N_3809,N_3701);
nor U4074 (N_4074,N_3760,N_3962);
nor U4075 (N_4075,N_2478,N_3692);
nor U4076 (N_4076,N_2795,N_3671);
or U4077 (N_4077,N_2972,N_2898);
nor U4078 (N_4078,N_3028,N_2220);
or U4079 (N_4079,N_2977,N_2140);
or U4080 (N_4080,N_2660,N_2359);
or U4081 (N_4081,N_3579,N_3208);
nand U4082 (N_4082,N_2257,N_3539);
and U4083 (N_4083,N_2862,N_2925);
nor U4084 (N_4084,N_3750,N_3036);
nor U4085 (N_4085,N_2101,N_2292);
or U4086 (N_4086,N_2067,N_2420);
nand U4087 (N_4087,N_2502,N_3061);
or U4088 (N_4088,N_2042,N_2134);
nor U4089 (N_4089,N_2129,N_2489);
xor U4090 (N_4090,N_3981,N_3311);
and U4091 (N_4091,N_3065,N_3260);
and U4092 (N_4092,N_2322,N_3347);
and U4093 (N_4093,N_3497,N_2849);
and U4094 (N_4094,N_2205,N_3441);
nand U4095 (N_4095,N_2604,N_2890);
and U4096 (N_4096,N_3118,N_2208);
nor U4097 (N_4097,N_3997,N_3918);
and U4098 (N_4098,N_2924,N_3874);
nor U4099 (N_4099,N_2334,N_2476);
or U4100 (N_4100,N_2073,N_2559);
nor U4101 (N_4101,N_3310,N_3569);
nor U4102 (N_4102,N_2427,N_3573);
or U4103 (N_4103,N_3540,N_3097);
or U4104 (N_4104,N_2059,N_3303);
nand U4105 (N_4105,N_3264,N_3585);
and U4106 (N_4106,N_3026,N_3940);
and U4107 (N_4107,N_2927,N_2630);
nand U4108 (N_4108,N_3453,N_3361);
nand U4109 (N_4109,N_2305,N_3547);
nor U4110 (N_4110,N_3111,N_2000);
and U4111 (N_4111,N_3998,N_2856);
nand U4112 (N_4112,N_3022,N_2254);
nor U4113 (N_4113,N_3382,N_3717);
and U4114 (N_4114,N_3304,N_2109);
or U4115 (N_4115,N_3526,N_2398);
or U4116 (N_4116,N_3056,N_3733);
and U4117 (N_4117,N_2289,N_2777);
and U4118 (N_4118,N_2947,N_2068);
nand U4119 (N_4119,N_3449,N_3673);
and U4120 (N_4120,N_2687,N_2242);
or U4121 (N_4121,N_3629,N_2221);
nor U4122 (N_4122,N_3858,N_3420);
and U4123 (N_4123,N_2191,N_2483);
nand U4124 (N_4124,N_2789,N_3813);
or U4125 (N_4125,N_3235,N_2845);
nand U4126 (N_4126,N_2193,N_3042);
nand U4127 (N_4127,N_2118,N_3136);
or U4128 (N_4128,N_2296,N_2550);
and U4129 (N_4129,N_3726,N_3409);
nor U4130 (N_4130,N_2547,N_2780);
nand U4131 (N_4131,N_2211,N_3805);
or U4132 (N_4132,N_2202,N_3468);
nand U4133 (N_4133,N_2750,N_2348);
nor U4134 (N_4134,N_3455,N_2536);
nor U4135 (N_4135,N_3198,N_3883);
nand U4136 (N_4136,N_3333,N_3882);
nor U4137 (N_4137,N_2116,N_3752);
and U4138 (N_4138,N_3920,N_2815);
nand U4139 (N_4139,N_3716,N_3895);
or U4140 (N_4140,N_2691,N_2929);
or U4141 (N_4141,N_2009,N_3532);
or U4142 (N_4142,N_3742,N_2356);
nand U4143 (N_4143,N_2365,N_2820);
and U4144 (N_4144,N_2993,N_2791);
and U4145 (N_4145,N_2194,N_3330);
nand U4146 (N_4146,N_2326,N_2635);
or U4147 (N_4147,N_3143,N_2453);
nand U4148 (N_4148,N_3634,N_2911);
nor U4149 (N_4149,N_2718,N_3043);
or U4150 (N_4150,N_2654,N_2506);
nand U4151 (N_4151,N_2987,N_2546);
or U4152 (N_4152,N_3217,N_3631);
nor U4153 (N_4153,N_2669,N_3243);
nand U4154 (N_4154,N_3439,N_3511);
nor U4155 (N_4155,N_3248,N_3234);
xnor U4156 (N_4156,N_2433,N_3106);
and U4157 (N_4157,N_2708,N_2075);
nand U4158 (N_4158,N_2263,N_3285);
nand U4159 (N_4159,N_2937,N_2394);
nor U4160 (N_4160,N_3318,N_2473);
nand U4161 (N_4161,N_3514,N_2794);
or U4162 (N_4162,N_2170,N_2539);
xnor U4163 (N_4163,N_2672,N_3275);
nand U4164 (N_4164,N_3801,N_2798);
nor U4165 (N_4165,N_3126,N_2367);
nor U4166 (N_4166,N_2426,N_2318);
and U4167 (N_4167,N_2537,N_2531);
nand U4168 (N_4168,N_2739,N_2282);
nand U4169 (N_4169,N_3331,N_3964);
or U4170 (N_4170,N_3067,N_2567);
or U4171 (N_4171,N_3712,N_3093);
nand U4172 (N_4172,N_3320,N_2406);
and U4173 (N_4173,N_3663,N_3084);
nor U4174 (N_4174,N_3381,N_3740);
nand U4175 (N_4175,N_2379,N_2555);
or U4176 (N_4176,N_2907,N_3486);
and U4177 (N_4177,N_2858,N_3635);
nand U4178 (N_4178,N_3161,N_3616);
and U4179 (N_4179,N_2275,N_2983);
nand U4180 (N_4180,N_2981,N_2201);
nand U4181 (N_4181,N_3821,N_2239);
nand U4182 (N_4182,N_3884,N_2371);
nand U4183 (N_4183,N_3649,N_2891);
nor U4184 (N_4184,N_3522,N_2773);
or U4185 (N_4185,N_3085,N_3559);
nor U4186 (N_4186,N_3328,N_3887);
xnor U4187 (N_4187,N_3183,N_3510);
nor U4188 (N_4188,N_2989,N_2261);
nor U4189 (N_4189,N_2222,N_3851);
nor U4190 (N_4190,N_2589,N_2720);
nor U4191 (N_4191,N_3790,N_3737);
or U4192 (N_4192,N_3447,N_2033);
nand U4193 (N_4193,N_3930,N_2574);
and U4194 (N_4194,N_2049,N_3076);
nor U4195 (N_4195,N_2328,N_2124);
or U4196 (N_4196,N_3627,N_3181);
or U4197 (N_4197,N_3309,N_3113);
nand U4198 (N_4198,N_3211,N_2992);
or U4199 (N_4199,N_2309,N_2681);
or U4200 (N_4200,N_3495,N_2990);
nand U4201 (N_4201,N_2542,N_2668);
nor U4202 (N_4202,N_3125,N_3202);
and U4203 (N_4203,N_3975,N_3520);
nor U4204 (N_4204,N_2047,N_2072);
nor U4205 (N_4205,N_3864,N_3957);
nor U4206 (N_4206,N_2692,N_3951);
nor U4207 (N_4207,N_2581,N_2760);
or U4208 (N_4208,N_3578,N_2299);
nor U4209 (N_4209,N_2642,N_3687);
nor U4210 (N_4210,N_3581,N_2885);
nor U4211 (N_4211,N_3702,N_2474);
nor U4212 (N_4212,N_3377,N_2504);
xor U4213 (N_4213,N_2045,N_2251);
and U4214 (N_4214,N_3542,N_3480);
and U4215 (N_4215,N_2472,N_3002);
or U4216 (N_4216,N_3277,N_3134);
nor U4217 (N_4217,N_3506,N_3850);
nor U4218 (N_4218,N_2311,N_3855);
and U4219 (N_4219,N_3120,N_2843);
and U4220 (N_4220,N_2648,N_3639);
and U4221 (N_4221,N_2920,N_3936);
or U4222 (N_4222,N_3242,N_2250);
or U4223 (N_4223,N_3463,N_3301);
and U4224 (N_4224,N_3624,N_3744);
and U4225 (N_4225,N_3466,N_3139);
nand U4226 (N_4226,N_3718,N_3488);
nand U4227 (N_4227,N_3808,N_2874);
or U4228 (N_4228,N_2022,N_3602);
nor U4229 (N_4229,N_2454,N_3358);
nor U4230 (N_4230,N_2225,N_3390);
and U4231 (N_4231,N_3681,N_3141);
nand U4232 (N_4232,N_3854,N_2169);
and U4233 (N_4233,N_3767,N_2150);
nand U4234 (N_4234,N_3349,N_2959);
and U4235 (N_4235,N_3195,N_3741);
nand U4236 (N_4236,N_3316,N_3429);
and U4237 (N_4237,N_3035,N_3329);
nor U4238 (N_4238,N_2808,N_2197);
xor U4239 (N_4239,N_2561,N_2636);
or U4240 (N_4240,N_2556,N_3656);
or U4241 (N_4241,N_3170,N_2355);
and U4242 (N_4242,N_3149,N_2580);
nor U4243 (N_4243,N_2434,N_3492);
and U4244 (N_4244,N_2627,N_3313);
and U4245 (N_4245,N_3612,N_3852);
and U4246 (N_4246,N_3778,N_2715);
nand U4247 (N_4247,N_3297,N_3866);
nor U4248 (N_4248,N_2023,N_3846);
or U4249 (N_4249,N_2390,N_3047);
nor U4250 (N_4250,N_3481,N_2244);
nor U4251 (N_4251,N_2594,N_3350);
or U4252 (N_4252,N_3008,N_2260);
or U4253 (N_4253,N_3816,N_3664);
and U4254 (N_4254,N_2688,N_2368);
and U4255 (N_4255,N_3682,N_3469);
nand U4256 (N_4256,N_3798,N_2183);
or U4257 (N_4257,N_2304,N_2219);
and U4258 (N_4258,N_2952,N_2479);
and U4259 (N_4259,N_2797,N_3595);
nor U4260 (N_4260,N_3580,N_2956);
or U4261 (N_4261,N_3119,N_3426);
nand U4262 (N_4262,N_2375,N_3324);
or U4263 (N_4263,N_3533,N_2682);
nor U4264 (N_4264,N_3570,N_2906);
nand U4265 (N_4265,N_2778,N_2693);
and U4266 (N_4266,N_2686,N_2230);
or U4267 (N_4267,N_2343,N_3241);
and U4268 (N_4268,N_2839,N_2618);
nand U4269 (N_4269,N_2889,N_3132);
nor U4270 (N_4270,N_2733,N_2768);
nand U4271 (N_4271,N_3236,N_2850);
and U4272 (N_4272,N_3223,N_3166);
or U4273 (N_4273,N_2548,N_2493);
nand U4274 (N_4274,N_3867,N_2520);
nor U4275 (N_4275,N_3189,N_2883);
nand U4276 (N_4276,N_3456,N_2784);
or U4277 (N_4277,N_2117,N_2827);
nor U4278 (N_4278,N_2016,N_3169);
xnor U4279 (N_4279,N_3342,N_2481);
nor U4280 (N_4280,N_2015,N_2098);
or U4281 (N_4281,N_3129,N_3465);
and U4282 (N_4282,N_3937,N_2389);
nor U4283 (N_4283,N_3605,N_3888);
or U4284 (N_4284,N_3491,N_2273);
or U4285 (N_4285,N_3844,N_2128);
and U4286 (N_4286,N_2841,N_2048);
nor U4287 (N_4287,N_2484,N_2980);
nor U4288 (N_4288,N_3954,N_2737);
or U4289 (N_4289,N_3856,N_3057);
or U4290 (N_4290,N_2111,N_3587);
or U4291 (N_4291,N_2800,N_3379);
nand U4292 (N_4292,N_3218,N_3552);
or U4293 (N_4293,N_2352,N_3910);
nor U4294 (N_4294,N_3448,N_3317);
nor U4295 (N_4295,N_3025,N_3558);
or U4296 (N_4296,N_2951,N_2694);
nor U4297 (N_4297,N_3151,N_2206);
nand U4298 (N_4298,N_3519,N_2008);
or U4299 (N_4299,N_3776,N_2457);
and U4300 (N_4300,N_2076,N_3295);
or U4301 (N_4301,N_3986,N_2280);
nand U4302 (N_4302,N_2517,N_2425);
and U4303 (N_4303,N_3068,N_3294);
nor U4304 (N_4304,N_3859,N_2510);
nand U4305 (N_4305,N_3323,N_3932);
or U4306 (N_4306,N_2180,N_2727);
nand U4307 (N_4307,N_2946,N_2450);
and U4308 (N_4308,N_3645,N_2775);
and U4309 (N_4309,N_3479,N_2902);
or U4310 (N_4310,N_2879,N_3660);
nor U4311 (N_4311,N_3140,N_3273);
and U4312 (N_4312,N_3630,N_3765);
and U4313 (N_4313,N_2615,N_3501);
nand U4314 (N_4314,N_3372,N_2069);
or U4315 (N_4315,N_2495,N_2057);
nor U4316 (N_4316,N_2557,N_2840);
nor U4317 (N_4317,N_3029,N_2161);
nand U4318 (N_4318,N_3411,N_2383);
or U4319 (N_4319,N_3362,N_3450);
and U4320 (N_4320,N_3751,N_2892);
and U4321 (N_4321,N_2712,N_2870);
or U4322 (N_4322,N_3768,N_2264);
and U4323 (N_4323,N_3898,N_3677);
nand U4324 (N_4324,N_3326,N_3446);
nor U4325 (N_4325,N_3144,N_2471);
nand U4326 (N_4326,N_3865,N_3384);
or U4327 (N_4327,N_2325,N_3387);
and U4328 (N_4328,N_2700,N_2975);
nor U4329 (N_4329,N_2358,N_3225);
nor U4330 (N_4330,N_2706,N_3493);
nor U4331 (N_4331,N_3464,N_2285);
and U4332 (N_4332,N_3689,N_2595);
or U4333 (N_4333,N_3648,N_2793);
nor U4334 (N_4334,N_2649,N_2698);
nor U4335 (N_4335,N_3902,N_3529);
nand U4336 (N_4336,N_3268,N_3032);
nand U4337 (N_4337,N_3412,N_2710);
and U4338 (N_4338,N_2307,N_2277);
nand U4339 (N_4339,N_2541,N_3165);
nand U4340 (N_4340,N_2602,N_2154);
nand U4341 (N_4341,N_3562,N_3598);
and U4342 (N_4342,N_3607,N_3394);
nand U4343 (N_4343,N_2848,N_2090);
and U4344 (N_4344,N_2174,N_2021);
or U4345 (N_4345,N_3452,N_3210);
nor U4346 (N_4346,N_3205,N_3794);
and U4347 (N_4347,N_3781,N_2428);
and U4348 (N_4348,N_3299,N_2132);
and U4349 (N_4349,N_2684,N_3315);
nand U4350 (N_4350,N_2665,N_2342);
or U4351 (N_4351,N_3738,N_2657);
and U4352 (N_4352,N_2185,N_3280);
and U4353 (N_4353,N_3188,N_3440);
and U4354 (N_4354,N_2153,N_2932);
and U4355 (N_4355,N_3247,N_3665);
or U4356 (N_4356,N_3334,N_3594);
or U4357 (N_4357,N_2351,N_2449);
nor U4358 (N_4358,N_3582,N_3960);
nor U4359 (N_4359,N_3990,N_2492);
or U4360 (N_4360,N_3459,N_3661);
or U4361 (N_4361,N_2463,N_3389);
and U4362 (N_4362,N_2417,N_3088);
nor U4363 (N_4363,N_3788,N_3471);
and U4364 (N_4364,N_3475,N_3355);
nand U4365 (N_4365,N_3840,N_2620);
nand U4366 (N_4366,N_3947,N_2447);
and U4367 (N_4367,N_2816,N_3916);
or U4368 (N_4368,N_3819,N_2772);
or U4369 (N_4369,N_3828,N_2507);
and U4370 (N_4370,N_2270,N_2978);
nor U4371 (N_4371,N_2386,N_2944);
or U4372 (N_4372,N_3040,N_3020);
nor U4373 (N_4373,N_2044,N_2213);
or U4374 (N_4374,N_2078,N_2357);
or U4375 (N_4375,N_3684,N_3713);
nor U4376 (N_4376,N_3319,N_2207);
or U4377 (N_4377,N_3626,N_2742);
or U4378 (N_4378,N_3160,N_2019);
and U4379 (N_4379,N_2231,N_3676);
or U4380 (N_4380,N_2579,N_2626);
and U4381 (N_4381,N_3064,N_3278);
nand U4382 (N_4382,N_3604,N_2976);
nand U4383 (N_4383,N_2014,N_3422);
nor U4384 (N_4384,N_3051,N_3445);
nand U4385 (N_4385,N_2486,N_3793);
nor U4386 (N_4386,N_2647,N_3290);
nand U4387 (N_4387,N_3695,N_3655);
nor U4388 (N_4388,N_3261,N_2158);
nor U4389 (N_4389,N_3747,N_3150);
nand U4390 (N_4390,N_3619,N_2624);
or U4391 (N_4391,N_3398,N_2893);
nor U4392 (N_4392,N_2832,N_3325);
or U4393 (N_4393,N_2746,N_3091);
nand U4394 (N_4394,N_2919,N_2948);
nand U4395 (N_4395,N_3039,N_2258);
and U4396 (N_4396,N_2817,N_2743);
nor U4397 (N_4397,N_3062,N_3368);
xnor U4398 (N_4398,N_3536,N_2731);
nor U4399 (N_4399,N_3842,N_2511);
nand U4400 (N_4400,N_3354,N_2198);
nand U4401 (N_4401,N_3286,N_2041);
and U4402 (N_4402,N_2184,N_2591);
nor U4403 (N_4403,N_2435,N_2966);
nor U4404 (N_4404,N_2818,N_3906);
and U4405 (N_4405,N_3836,N_2488);
nor U4406 (N_4406,N_2092,N_3576);
nor U4407 (N_4407,N_2835,N_2652);
nor U4408 (N_4408,N_2998,N_2335);
nand U4409 (N_4409,N_3516,N_3094);
nand U4410 (N_4410,N_3667,N_3697);
and U4411 (N_4411,N_3670,N_2645);
and U4412 (N_4412,N_2910,N_3180);
and U4413 (N_4413,N_2246,N_3857);
and U4414 (N_4414,N_3803,N_3001);
and U4415 (N_4415,N_3182,N_2600);
nor U4416 (N_4416,N_3504,N_3224);
nor U4417 (N_4417,N_3096,N_2704);
nor U4418 (N_4418,N_2991,N_3853);
or U4419 (N_4419,N_2745,N_3623);
nand U4420 (N_4420,N_2136,N_2529);
nand U4421 (N_4421,N_2763,N_2518);
nand U4422 (N_4422,N_2249,N_3652);
nand U4423 (N_4423,N_2317,N_3050);
nand U4424 (N_4424,N_3237,N_2823);
xor U4425 (N_4425,N_2160,N_3560);
or U4426 (N_4426,N_2364,N_3722);
and U4427 (N_4427,N_2689,N_2968);
nand U4428 (N_4428,N_3427,N_2327);
nand U4429 (N_4429,N_3924,N_2578);
or U4430 (N_4430,N_3685,N_2152);
nand U4431 (N_4431,N_3693,N_3704);
or U4432 (N_4432,N_2411,N_3457);
nor U4433 (N_4433,N_3383,N_3941);
nor U4434 (N_4434,N_2830,N_2462);
nand U4435 (N_4435,N_2377,N_3757);
nand U4436 (N_4436,N_2590,N_2888);
and U4437 (N_4437,N_2528,N_2851);
and U4438 (N_4438,N_3996,N_2515);
or U4439 (N_4439,N_3730,N_3003);
nand U4440 (N_4440,N_2679,N_3621);
nand U4441 (N_4441,N_3131,N_2468);
or U4442 (N_4442,N_3415,N_3152);
or U4443 (N_4443,N_2740,N_2942);
nand U4444 (N_4444,N_3779,N_3431);
or U4445 (N_4445,N_3834,N_2637);
and U4446 (N_4446,N_3706,N_2464);
nor U4447 (N_4447,N_3544,N_2928);
nor U4448 (N_4448,N_2809,N_2619);
nand U4449 (N_4449,N_3499,N_2878);
nor U4450 (N_4450,N_3838,N_3507);
nor U4451 (N_4451,N_2792,N_2563);
nand U4452 (N_4452,N_2051,N_3546);
and U4453 (N_4453,N_3458,N_3231);
xnor U4454 (N_4454,N_3974,N_3592);
nand U4455 (N_4455,N_3291,N_3123);
nor U4456 (N_4456,N_2683,N_3045);
or U4457 (N_4457,N_2131,N_2165);
xnor U4458 (N_4458,N_3462,N_3265);
and U4459 (N_4459,N_2667,N_2460);
nor U4460 (N_4460,N_2774,N_2926);
or U4461 (N_4461,N_2224,N_3336);
nand U4462 (N_4462,N_3403,N_3414);
or U4463 (N_4463,N_2141,N_3896);
and U4464 (N_4464,N_2573,N_2521);
or U4465 (N_4465,N_2921,N_3928);
nor U4466 (N_4466,N_2027,N_3146);
nor U4467 (N_4467,N_3553,N_3175);
or U4468 (N_4468,N_2705,N_2958);
nor U4469 (N_4469,N_3564,N_3395);
xor U4470 (N_4470,N_3015,N_3346);
or U4471 (N_4471,N_3332,N_2505);
nand U4472 (N_4472,N_3474,N_3171);
nor U4473 (N_4473,N_3890,N_3642);
nor U4474 (N_4474,N_2569,N_2281);
and U4475 (N_4475,N_3069,N_3758);
nand U4476 (N_4476,N_2759,N_3433);
nand U4477 (N_4477,N_2064,N_2480);
nand U4478 (N_4478,N_3708,N_3966);
nor U4479 (N_4479,N_2960,N_3797);
nor U4480 (N_4480,N_2728,N_2192);
or U4481 (N_4481,N_3786,N_3509);
and U4482 (N_4482,N_3774,N_3438);
xor U4483 (N_4483,N_3787,N_3643);
nand U4484 (N_4484,N_3696,N_2810);
nor U4485 (N_4485,N_3103,N_3977);
or U4486 (N_4486,N_2104,N_3258);
nand U4487 (N_4487,N_2905,N_2405);
and U4488 (N_4488,N_3982,N_3720);
or U4489 (N_4489,N_3269,N_3262);
nand U4490 (N_4490,N_3829,N_3168);
nor U4491 (N_4491,N_2622,N_2094);
or U4492 (N_4492,N_3352,N_3081);
or U4493 (N_4493,N_3058,N_3688);
or U4494 (N_4494,N_2181,N_2957);
nand U4495 (N_4495,N_3430,N_3341);
and U4496 (N_4496,N_2909,N_2709);
nor U4497 (N_4497,N_2599,N_2525);
and U4498 (N_4498,N_3548,N_2714);
nand U4499 (N_4499,N_2262,N_2685);
or U4500 (N_4500,N_2984,N_2629);
nand U4501 (N_4501,N_3215,N_2102);
and U4502 (N_4502,N_2918,N_3976);
nand U4503 (N_4503,N_2232,N_2996);
nand U4504 (N_4504,N_3791,N_3603);
or U4505 (N_4505,N_2606,N_2279);
nor U4506 (N_4506,N_2875,N_2287);
and U4507 (N_4507,N_2218,N_2291);
nand U4508 (N_4508,N_3675,N_3782);
nand U4509 (N_4509,N_3807,N_3613);
xnor U4510 (N_4510,N_3538,N_2703);
nand U4511 (N_4511,N_3527,N_2553);
xor U4512 (N_4512,N_3321,N_2801);
and U4513 (N_4513,N_2146,N_2565);
nand U4514 (N_4514,N_2509,N_2234);
nor U4515 (N_4515,N_3482,N_2829);
or U4516 (N_4516,N_2508,N_2302);
or U4517 (N_4517,N_3968,N_2988);
nor U4518 (N_4518,N_3221,N_2994);
or U4519 (N_4519,N_3899,N_3154);
nor U4520 (N_4520,N_3245,N_3005);
nor U4521 (N_4521,N_3199,N_3574);
xnor U4522 (N_4522,N_3046,N_2598);
or U4523 (N_4523,N_2717,N_2121);
nand U4524 (N_4524,N_3083,N_3338);
nand U4525 (N_4525,N_3992,N_3135);
or U4526 (N_4526,N_3041,N_3824);
nor U4527 (N_4527,N_3272,N_2857);
xor U4528 (N_4528,N_2954,N_3531);
or U4529 (N_4529,N_2695,N_2696);
nand U4530 (N_4530,N_2482,N_3847);
or U4531 (N_4531,N_3393,N_2392);
and U4532 (N_4532,N_2204,N_2333);
nor U4533 (N_4533,N_2112,N_3994);
and U4534 (N_4534,N_3121,N_3638);
and U4535 (N_4535,N_3873,N_2422);
nor U4536 (N_4536,N_3351,N_3679);
or U4537 (N_4537,N_2512,N_2741);
or U4538 (N_4538,N_2188,N_2038);
nor U4539 (N_4539,N_3929,N_2723);
or U4540 (N_4540,N_2965,N_3657);
nand U4541 (N_4541,N_2475,N_2713);
and U4542 (N_4542,N_3487,N_2625);
nor U4543 (N_4543,N_3875,N_2771);
nand U4544 (N_4544,N_3340,N_2455);
or U4545 (N_4545,N_2628,N_3314);
xor U4546 (N_4546,N_2834,N_2324);
nor U4547 (N_4547,N_3007,N_3470);
nand U4548 (N_4548,N_3376,N_3206);
and U4549 (N_4549,N_3818,N_3618);
and U4550 (N_4550,N_3878,N_3018);
nand U4551 (N_4551,N_2757,N_2634);
nor U4552 (N_4552,N_3955,N_3437);
and U4553 (N_4553,N_2303,N_2349);
nor U4554 (N_4554,N_3907,N_2173);
and U4555 (N_4555,N_2007,N_2143);
nand U4556 (N_4556,N_2755,N_2609);
nor U4557 (N_4557,N_2344,N_2466);
and U4558 (N_4558,N_3919,N_3724);
nor U4559 (N_4559,N_3399,N_2999);
and U4560 (N_4560,N_2514,N_2004);
nand U4561 (N_4561,N_3053,N_2155);
nand U4562 (N_4562,N_2982,N_2052);
nor U4563 (N_4563,N_2562,N_3153);
nor U4564 (N_4564,N_3909,N_2490);
or U4565 (N_4565,N_3792,N_3711);
and U4566 (N_4566,N_2608,N_3795);
nor U4567 (N_4567,N_3641,N_3777);
or U4568 (N_4568,N_3911,N_3212);
and U4569 (N_4569,N_3417,N_2551);
and U4570 (N_4570,N_2877,N_2002);
or U4571 (N_4571,N_3785,N_3108);
nand U4572 (N_4572,N_2596,N_3835);
or U4573 (N_4573,N_2332,N_3732);
and U4574 (N_4574,N_2656,N_3375);
nor U4575 (N_4575,N_2025,N_3203);
and U4576 (N_4576,N_2836,N_3654);
nor U4577 (N_4577,N_3367,N_2666);
and U4578 (N_4578,N_2886,N_2491);
and U4579 (N_4579,N_2217,N_3425);
and U4580 (N_4580,N_2283,N_2190);
and U4581 (N_4581,N_3993,N_2077);
nand U4582 (N_4582,N_3727,N_3100);
nor U4583 (N_4583,N_2837,N_3467);
nor U4584 (N_4584,N_3939,N_3019);
and U4585 (N_4585,N_2498,N_2538);
xnor U4586 (N_4586,N_3644,N_2516);
or U4587 (N_4587,N_2765,N_2833);
and U4588 (N_4588,N_3705,N_3922);
or U4589 (N_4589,N_2871,N_2148);
or U4590 (N_4590,N_2969,N_3596);
and U4591 (N_4591,N_2540,N_3796);
nand U4592 (N_4592,N_2577,N_2545);
or U4593 (N_4593,N_3263,N_3766);
and U4594 (N_4594,N_3079,N_2900);
nor U4595 (N_4595,N_2861,N_3622);
nor U4596 (N_4596,N_2215,N_3059);
and U4597 (N_4597,N_2452,N_3897);
or U4598 (N_4598,N_3098,N_3551);
nor U4599 (N_4599,N_3513,N_3736);
xor U4600 (N_4600,N_2223,N_3259);
nor U4601 (N_4601,N_3691,N_3386);
and U4602 (N_4602,N_3049,N_2825);
nor U4603 (N_4603,N_3698,N_2640);
nand U4604 (N_4604,N_3254,N_3253);
or U4605 (N_4605,N_3282,N_3870);
or U4606 (N_4606,N_2441,N_3549);
and U4607 (N_4607,N_3577,N_3952);
nor U4608 (N_4608,N_3980,N_3201);
nor U4609 (N_4609,N_2524,N_3680);
and U4610 (N_4610,N_2503,N_3012);
nor U4611 (N_4611,N_2985,N_2295);
nor U4612 (N_4612,N_2252,N_3138);
or U4613 (N_4613,N_2724,N_2526);
nand U4614 (N_4614,N_3860,N_2922);
nor U4615 (N_4615,N_3037,N_2272);
and U4616 (N_4616,N_2576,N_2401);
and U4617 (N_4617,N_3943,N_3204);
nor U4618 (N_4618,N_2337,N_2804);
or U4619 (N_4619,N_2028,N_3886);
and U4620 (N_4620,N_3961,N_2088);
nor U4621 (N_4621,N_2549,N_2350);
nand U4622 (N_4622,N_3308,N_2340);
or U4623 (N_4623,N_2632,N_2868);
nor U4624 (N_4624,N_2722,N_2587);
nand U4625 (N_4625,N_3583,N_3973);
nand U4626 (N_4626,N_3443,N_3999);
nor U4627 (N_4627,N_3921,N_2881);
nor U4628 (N_4628,N_2783,N_2354);
or U4629 (N_4629,N_2864,N_2268);
nand U4630 (N_4630,N_3289,N_2167);
nor U4631 (N_4631,N_2353,N_2500);
or U4632 (N_4632,N_3238,N_2729);
nor U4633 (N_4633,N_3668,N_2013);
and U4634 (N_4634,N_3274,N_2133);
nand U4635 (N_4635,N_3388,N_2440);
nand U4636 (N_4636,N_3107,N_2026);
and U4637 (N_4637,N_3073,N_2882);
nand U4638 (N_4638,N_3196,N_2237);
nor U4639 (N_4639,N_2738,N_2079);
and U4640 (N_4640,N_3178,N_3112);
or U4641 (N_4641,N_3116,N_2439);
nor U4642 (N_4642,N_3192,N_2872);
or U4643 (N_4643,N_2011,N_3363);
or U4644 (N_4644,N_3287,N_3322);
or U4645 (N_4645,N_3694,N_2865);
or U4646 (N_4646,N_2697,N_3841);
or U4647 (N_4647,N_3979,N_2020);
nand U4648 (N_4648,N_2611,N_3461);
xnor U4649 (N_4649,N_2424,N_3972);
or U4650 (N_4650,N_3087,N_3266);
xor U4651 (N_4651,N_2796,N_2790);
nor U4652 (N_4652,N_3748,N_3055);
nor U4653 (N_4653,N_3518,N_3590);
or U4654 (N_4654,N_3735,N_3650);
and U4655 (N_4655,N_2397,N_2527);
nor U4656 (N_4656,N_3117,N_2284);
and U4657 (N_4657,N_3880,N_2934);
nor U4658 (N_4658,N_3614,N_2497);
or U4659 (N_4659,N_3066,N_3292);
nor U4660 (N_4660,N_2407,N_2601);
or U4661 (N_4661,N_2286,N_3004);
or U4662 (N_4662,N_2276,N_3074);
nor U4663 (N_4663,N_2431,N_2838);
nor U4664 (N_4664,N_3721,N_2572);
nand U4665 (N_4665,N_3366,N_2854);
nor U4666 (N_4666,N_3370,N_3498);
nor U4667 (N_4667,N_2967,N_3207);
or U4668 (N_4668,N_3764,N_2962);
and U4669 (N_4669,N_3031,N_2662);
nand U4670 (N_4670,N_3715,N_3876);
nand U4671 (N_4671,N_3755,N_2605);
nand U4672 (N_4672,N_3163,N_3615);
nor U4673 (N_4673,N_3219,N_3267);
nand U4674 (N_4674,N_2055,N_3044);
or U4675 (N_4675,N_3246,N_3010);
and U4676 (N_4676,N_2336,N_2093);
and U4677 (N_4677,N_2806,N_3659);
nor U4678 (N_4678,N_3416,N_2418);
or U4679 (N_4679,N_3861,N_2046);
and U4680 (N_4680,N_2321,N_2314);
and U4681 (N_4681,N_2664,N_3174);
nand U4682 (N_4682,N_2151,N_3608);
and U4683 (N_4683,N_3339,N_3408);
nor U4684 (N_4684,N_2054,N_2267);
and U4685 (N_4685,N_2867,N_2730);
nand U4686 (N_4686,N_2396,N_3380);
nand U4687 (N_4687,N_3162,N_3651);
or U4688 (N_4688,N_2071,N_3256);
nor U4689 (N_4689,N_2597,N_2248);
and U4690 (N_4690,N_3194,N_3761);
nand U4691 (N_4691,N_2534,N_3783);
and U4692 (N_4692,N_2614,N_3554);
or U4693 (N_4693,N_3110,N_2748);
or U4694 (N_4694,N_3476,N_3048);
and U4695 (N_4695,N_3222,N_3023);
and U4696 (N_4696,N_2266,N_2039);
nand U4697 (N_4697,N_3164,N_2096);
or U4698 (N_4698,N_2895,N_2083);
and U4699 (N_4699,N_3837,N_2209);
and U4700 (N_4700,N_2904,N_3600);
and U4701 (N_4701,N_2873,N_2265);
and U4702 (N_4702,N_3923,N_2187);
and U4703 (N_4703,N_3034,N_2945);
and U4704 (N_4704,N_2747,N_2487);
or U4705 (N_4705,N_3989,N_2347);
and U4706 (N_4706,N_3775,N_3122);
or U4707 (N_4707,N_2675,N_2108);
nor U4708 (N_4708,N_2166,N_3815);
nor U4709 (N_4709,N_2752,N_2552);
nor U4710 (N_4710,N_3894,N_2139);
and U4711 (N_4711,N_2753,N_2241);
or U4712 (N_4712,N_2674,N_2395);
nand U4713 (N_4713,N_3934,N_3889);
nor U4714 (N_4714,N_2788,N_2331);
or U4715 (N_4715,N_2678,N_3903);
and U4716 (N_4716,N_3508,N_3863);
xor U4717 (N_4717,N_2256,N_3185);
nor U4718 (N_4718,N_2451,N_2399);
xor U4719 (N_4719,N_2429,N_3137);
or U4720 (N_4720,N_2081,N_3477);
nand U4721 (N_4721,N_3072,N_3812);
or U4722 (N_4722,N_3027,N_2233);
or U4723 (N_4723,N_2533,N_3541);
nor U4724 (N_4724,N_2961,N_3572);
and U4725 (N_4725,N_3869,N_3759);
or U4726 (N_4726,N_3307,N_2040);
and U4727 (N_4727,N_2070,N_2584);
or U4728 (N_4728,N_2702,N_2880);
and U4729 (N_4729,N_2442,N_3646);
nor U4730 (N_4730,N_3988,N_3364);
xor U4731 (N_4731,N_3610,N_3571);
or U4732 (N_4732,N_2621,N_2159);
nand U4733 (N_4733,N_3105,N_3157);
or U4734 (N_4734,N_3515,N_2887);
and U4735 (N_4735,N_2711,N_3770);
and U4736 (N_4736,N_3401,N_3021);
nor U4737 (N_4737,N_2313,N_3563);
nand U4738 (N_4738,N_2938,N_3523);
and U4739 (N_4739,N_3545,N_3156);
and U4740 (N_4740,N_2633,N_2855);
nand U4741 (N_4741,N_2393,N_2373);
and U4742 (N_4742,N_3512,N_2430);
or U4743 (N_4743,N_3700,N_3543);
and U4744 (N_4744,N_2171,N_3769);
nor U4745 (N_4745,N_3155,N_2443);
nor U4746 (N_4746,N_2811,N_3927);
or U4747 (N_4747,N_3647,N_3734);
nor U4748 (N_4748,N_3365,N_2091);
and U4749 (N_4749,N_3800,N_3086);
nor U4750 (N_4750,N_2082,N_2680);
and U4751 (N_4751,N_3662,N_2470);
and U4752 (N_4752,N_3802,N_2869);
and U4753 (N_4753,N_3359,N_2053);
nor U4754 (N_4754,N_3353,N_2749);
and U4755 (N_4755,N_3946,N_3033);
and U4756 (N_4756,N_3833,N_2725);
nor U4757 (N_4757,N_2519,N_3773);
or U4758 (N_4758,N_2372,N_2259);
nand U4759 (N_4759,N_2650,N_3421);
nor U4760 (N_4760,N_3830,N_2699);
and U4761 (N_4761,N_2085,N_3606);
nand U4762 (N_4762,N_2963,N_2380);
and U4763 (N_4763,N_3276,N_2199);
nor U4764 (N_4764,N_2884,N_2494);
and U4765 (N_4765,N_2701,N_3995);
or U4766 (N_4766,N_3901,N_2345);
nand U4767 (N_4767,N_2762,N_3674);
or U4768 (N_4768,N_3820,N_2764);
nand U4769 (N_4769,N_2779,N_2564);
nand U4770 (N_4770,N_2227,N_3699);
or U4771 (N_4771,N_3095,N_2339);
nand U4772 (N_4772,N_2935,N_2178);
or U4773 (N_4773,N_2095,N_3078);
nor U4774 (N_4774,N_3473,N_3496);
or U4775 (N_4775,N_2588,N_2535);
or U4776 (N_4776,N_3077,N_2214);
nor U4777 (N_4777,N_3935,N_3080);
and U4778 (N_4778,N_3187,N_3784);
or U4779 (N_4779,N_2374,N_2182);
or U4780 (N_4780,N_3915,N_3232);
nor U4781 (N_4781,N_2144,N_3013);
or U4782 (N_4782,N_3756,N_2831);
nor U4783 (N_4783,N_2024,N_2914);
and U4784 (N_4784,N_2459,N_3987);
or U4785 (N_4785,N_2361,N_2799);
nand U4786 (N_4786,N_3343,N_3371);
or U4787 (N_4787,N_3419,N_2583);
or U4788 (N_4788,N_3369,N_3435);
nand U4789 (N_4789,N_2080,N_3686);
nand U4790 (N_4790,N_3424,N_2416);
or U4791 (N_4791,N_3402,N_2876);
nand U4792 (N_4792,N_2950,N_2501);
or U4793 (N_4793,N_3305,N_3406);
and U4794 (N_4794,N_3312,N_2930);
nand U4795 (N_4795,N_2415,N_2658);
or U4796 (N_4796,N_2754,N_2050);
or U4797 (N_4797,N_3410,N_3609);
nand U4798 (N_4798,N_3561,N_2274);
and U4799 (N_4799,N_2575,N_3293);
nand U4800 (N_4800,N_3849,N_3391);
nand U4801 (N_4801,N_3589,N_3710);
or U4802 (N_4802,N_2939,N_2613);
nand U4803 (N_4803,N_3038,N_2370);
nor U4804 (N_4804,N_2312,N_2863);
nor U4805 (N_4805,N_3678,N_2123);
and U4806 (N_4806,N_3938,N_2641);
and U4807 (N_4807,N_2933,N_3892);
and U4808 (N_4808,N_2168,N_2805);
nand U4809 (N_4809,N_3167,N_2964);
nor U4810 (N_4810,N_3597,N_2953);
nand U4811 (N_4811,N_3385,N_2544);
or U4812 (N_4812,N_3436,N_3089);
nand U4813 (N_4813,N_3345,N_2812);
nand U4814 (N_4814,N_3772,N_2243);
nor U4815 (N_4815,N_3991,N_3640);
and U4816 (N_4816,N_2385,N_3799);
or U4817 (N_4817,N_2853,N_2530);
and U4818 (N_4818,N_3133,N_3227);
or U4819 (N_4819,N_2228,N_3593);
or U4820 (N_4820,N_2736,N_2106);
nand U4821 (N_4821,N_2897,N_2369);
or U4822 (N_4822,N_2766,N_3848);
nand U4823 (N_4823,N_3233,N_2767);
nand U4824 (N_4824,N_2814,N_3070);
nand U4825 (N_4825,N_2670,N_3397);
or U4826 (N_4826,N_2087,N_2802);
and U4827 (N_4827,N_2147,N_3763);
and U4828 (N_4828,N_2086,N_3804);
or U4829 (N_4829,N_3270,N_2707);
and U4830 (N_4830,N_2110,N_3306);
and U4831 (N_4831,N_3555,N_2826);
or U4832 (N_4832,N_3209,N_2360);
or U4833 (N_4833,N_2756,N_2229);
or U4834 (N_4834,N_2973,N_3104);
nor U4835 (N_4835,N_2162,N_2315);
or U4836 (N_4836,N_2732,N_3690);
nand U4837 (N_4837,N_3230,N_3537);
nand U4838 (N_4838,N_3114,N_3826);
and U4839 (N_4839,N_3831,N_2126);
and U4840 (N_4840,N_3092,N_3703);
and U4841 (N_4841,N_3130,N_3599);
nand U4842 (N_4842,N_2119,N_3428);
and U4843 (N_4843,N_3729,N_2446);
and U4844 (N_4844,N_2066,N_3011);
nand U4845 (N_4845,N_2785,N_3839);
and U4846 (N_4846,N_3200,N_2543);
nand U4847 (N_4847,N_2297,N_3148);
or U4848 (N_4848,N_3244,N_3407);
and U4849 (N_4849,N_3249,N_2821);
nor U4850 (N_4850,N_2363,N_3271);
nor U4851 (N_4851,N_3568,N_3173);
nor U4852 (N_4852,N_2301,N_3124);
nor U4853 (N_4853,N_3418,N_2593);
nor U4854 (N_4854,N_2986,N_2142);
and U4855 (N_4855,N_2366,N_3827);
nand U4856 (N_4856,N_3075,N_3197);
nor U4857 (N_4857,N_3099,N_3142);
and U4858 (N_4858,N_3490,N_2908);
and U4859 (N_4859,N_2676,N_3284);
and U4860 (N_4860,N_2172,N_3158);
or U4861 (N_4861,N_2896,N_3127);
xnor U4862 (N_4862,N_2673,N_2496);
nand U4863 (N_4863,N_3255,N_3505);
and U4864 (N_4864,N_2247,N_3877);
or U4865 (N_4865,N_2089,N_2164);
nand U4866 (N_4866,N_2807,N_3754);
and U4867 (N_4867,N_2288,N_3823);
or U4868 (N_4868,N_2558,N_2438);
nand U4869 (N_4869,N_3484,N_2646);
or U4870 (N_4870,N_3825,N_3963);
nand U4871 (N_4871,N_3908,N_3914);
or U4872 (N_4872,N_2157,N_2860);
nor U4873 (N_4873,N_3925,N_2899);
and U4874 (N_4874,N_3746,N_2402);
nor U4875 (N_4875,N_3969,N_2995);
or U4876 (N_4876,N_3400,N_2643);
and U4877 (N_4877,N_2444,N_3948);
nor U4878 (N_4878,N_3071,N_2300);
nor U4879 (N_4879,N_2403,N_3528);
or U4880 (N_4880,N_2062,N_2436);
or U4881 (N_4881,N_2105,N_2617);
nor U4882 (N_4882,N_3885,N_3240);
nand U4883 (N_4883,N_3868,N_2010);
nor U4884 (N_4884,N_3871,N_3472);
or U4885 (N_4885,N_3281,N_3967);
or U4886 (N_4886,N_2653,N_3251);
or U4887 (N_4887,N_2822,N_3879);
or U4888 (N_4888,N_2032,N_3327);
or U4889 (N_4889,N_3177,N_2177);
or U4890 (N_4890,N_2751,N_3714);
and U4891 (N_4891,N_3983,N_3147);
nor U4892 (N_4892,N_3405,N_2568);
or U4893 (N_4893,N_2847,N_2787);
nor U4894 (N_4894,N_3636,N_2917);
or U4895 (N_4895,N_2156,N_2560);
nand U4896 (N_4896,N_2824,N_2671);
nand U4897 (N_4897,N_2362,N_3115);
nand U4898 (N_4898,N_2744,N_2030);
nor U4899 (N_4899,N_3984,N_2726);
xor U4900 (N_4900,N_3958,N_3288);
nand U4901 (N_4901,N_2894,N_2974);
nor U4902 (N_4902,N_3556,N_3374);
nor U4903 (N_4903,N_2661,N_2074);
and U4904 (N_4904,N_2651,N_3454);
or U4905 (N_4905,N_2940,N_3628);
xor U4906 (N_4906,N_2381,N_2448);
nor U4907 (N_4907,N_3335,N_2456);
and U4908 (N_4908,N_2571,N_2901);
nor U4909 (N_4909,N_2245,N_2776);
nor U4910 (N_4910,N_2781,N_2663);
nor U4911 (N_4911,N_2499,N_2828);
or U4912 (N_4912,N_2319,N_3220);
and U4913 (N_4913,N_3949,N_2176);
or U4914 (N_4914,N_2099,N_2003);
or U4915 (N_4915,N_2290,N_2943);
nor U4916 (N_4916,N_2107,N_3373);
nor U4917 (N_4917,N_2813,N_3179);
nor U4918 (N_4918,N_3434,N_3524);
or U4919 (N_4919,N_2644,N_3378);
nand U4920 (N_4920,N_2409,N_2522);
and U4921 (N_4921,N_2400,N_3302);
nor U4922 (N_4922,N_3502,N_2803);
and U4923 (N_4923,N_2017,N_2018);
nor U4924 (N_4924,N_2532,N_2979);
nor U4925 (N_4925,N_2770,N_3566);
or U4926 (N_4926,N_2603,N_2255);
nand U4927 (N_4927,N_3172,N_3250);
and U4928 (N_4928,N_3283,N_3944);
nand U4929 (N_4929,N_2240,N_3728);
or U4930 (N_4930,N_2734,N_2320);
nand U4931 (N_4931,N_3534,N_2852);
nand U4932 (N_4932,N_2949,N_3586);
nand U4933 (N_4933,N_3611,N_3862);
nand U4934 (N_4934,N_2638,N_2012);
or U4935 (N_4935,N_3535,N_3109);
and U4936 (N_4936,N_2034,N_2196);
nand U4937 (N_4937,N_3478,N_3719);
and U4938 (N_4938,N_2278,N_3971);
or U4939 (N_4939,N_3063,N_2859);
nor U4940 (N_4940,N_3298,N_3575);
nor U4941 (N_4941,N_3584,N_3356);
nor U4942 (N_4942,N_3591,N_3503);
nor U4943 (N_4943,N_3214,N_3006);
or U4944 (N_4944,N_2616,N_2236);
nand U4945 (N_4945,N_2513,N_2623);
or U4946 (N_4946,N_2469,N_2294);
nand U4947 (N_4947,N_2127,N_3931);
or U4948 (N_4948,N_3567,N_2346);
nor U4949 (N_4949,N_2186,N_2384);
and U4950 (N_4950,N_3444,N_3625);
or U4951 (N_4951,N_3633,N_2137);
and U4952 (N_4952,N_3017,N_2523);
nor U4953 (N_4953,N_3904,N_2941);
and U4954 (N_4954,N_2461,N_3191);
nor U4955 (N_4955,N_2719,N_3588);
and U4956 (N_4956,N_2306,N_3780);
nand U4957 (N_4957,N_2413,N_3442);
nand U4958 (N_4958,N_2971,N_3843);
and U4959 (N_4959,N_3743,N_2203);
nand U4960 (N_4960,N_3360,N_3228);
nor U4961 (N_4961,N_2554,N_2437);
or U4962 (N_4962,N_2387,N_2782);
and U4963 (N_4963,N_2735,N_2592);
or U4964 (N_4964,N_3184,N_3226);
nand U4965 (N_4965,N_3845,N_3637);
and U4966 (N_4966,N_3090,N_2212);
nand U4967 (N_4967,N_2308,N_3460);
and U4968 (N_4968,N_2330,N_3530);
nand U4969 (N_4969,N_3950,N_3872);
and U4970 (N_4970,N_2467,N_2006);
and U4971 (N_4971,N_2216,N_3762);
nor U4972 (N_4972,N_2769,N_3707);
or U4973 (N_4973,N_2138,N_3257);
and U4974 (N_4974,N_3617,N_3723);
or U4975 (N_4975,N_2195,N_3337);
nor U4976 (N_4976,N_3905,N_3489);
nor U4977 (N_4977,N_2566,N_3832);
nor U4978 (N_4978,N_2485,N_2001);
nand U4979 (N_4979,N_2931,N_3101);
nor U4980 (N_4980,N_3521,N_2065);
nand U4981 (N_4981,N_3102,N_2970);
or U4982 (N_4982,N_3881,N_2414);
and U4983 (N_4983,N_3814,N_2421);
or U4984 (N_4984,N_3917,N_2043);
nand U4985 (N_4985,N_2716,N_3771);
nor U4986 (N_4986,N_3817,N_2035);
and U4987 (N_4987,N_3900,N_3810);
or U4988 (N_4988,N_2842,N_2819);
nor U4989 (N_4989,N_2607,N_2659);
or U4990 (N_4990,N_3669,N_2903);
or U4991 (N_4991,N_2458,N_2391);
or U4992 (N_4992,N_2758,N_3891);
nand U4993 (N_4993,N_2100,N_2120);
and U4994 (N_4994,N_3344,N_3300);
or U4995 (N_4995,N_2423,N_3423);
and U4996 (N_4996,N_3731,N_3193);
or U4997 (N_4997,N_2382,N_3666);
nand U4998 (N_4998,N_2582,N_3913);
nand U4999 (N_4999,N_3557,N_2376);
nand U5000 (N_5000,N_3206,N_3736);
nor U5001 (N_5001,N_3072,N_3329);
nor U5002 (N_5002,N_3457,N_2470);
or U5003 (N_5003,N_2463,N_2352);
or U5004 (N_5004,N_2839,N_2644);
nor U5005 (N_5005,N_3186,N_2642);
or U5006 (N_5006,N_2169,N_3592);
nand U5007 (N_5007,N_2338,N_3260);
nand U5008 (N_5008,N_2576,N_3170);
nor U5009 (N_5009,N_3028,N_2426);
and U5010 (N_5010,N_2683,N_2869);
and U5011 (N_5011,N_2732,N_3329);
or U5012 (N_5012,N_3889,N_2064);
nand U5013 (N_5013,N_3866,N_3846);
nand U5014 (N_5014,N_3125,N_3182);
and U5015 (N_5015,N_3470,N_3673);
nand U5016 (N_5016,N_2009,N_2444);
nor U5017 (N_5017,N_3482,N_3333);
nor U5018 (N_5018,N_3657,N_2589);
and U5019 (N_5019,N_2190,N_2967);
or U5020 (N_5020,N_3540,N_3848);
xor U5021 (N_5021,N_2484,N_2730);
nand U5022 (N_5022,N_2417,N_2756);
xnor U5023 (N_5023,N_3399,N_3048);
or U5024 (N_5024,N_3674,N_3751);
nor U5025 (N_5025,N_2148,N_2749);
and U5026 (N_5026,N_2989,N_3304);
nand U5027 (N_5027,N_3969,N_2569);
nand U5028 (N_5028,N_3313,N_2660);
or U5029 (N_5029,N_2060,N_2040);
and U5030 (N_5030,N_3817,N_2612);
or U5031 (N_5031,N_3995,N_3417);
and U5032 (N_5032,N_3540,N_2293);
nor U5033 (N_5033,N_3141,N_3521);
nor U5034 (N_5034,N_3022,N_2483);
nand U5035 (N_5035,N_3424,N_3287);
nor U5036 (N_5036,N_2697,N_3262);
nand U5037 (N_5037,N_2678,N_2136);
nor U5038 (N_5038,N_3588,N_3353);
or U5039 (N_5039,N_2248,N_3276);
nor U5040 (N_5040,N_3606,N_3268);
or U5041 (N_5041,N_3564,N_3205);
and U5042 (N_5042,N_3539,N_2124);
nor U5043 (N_5043,N_2943,N_3270);
and U5044 (N_5044,N_3175,N_2007);
and U5045 (N_5045,N_3829,N_2909);
or U5046 (N_5046,N_2073,N_3256);
and U5047 (N_5047,N_2308,N_3766);
and U5048 (N_5048,N_3385,N_3540);
nand U5049 (N_5049,N_3214,N_2289);
nand U5050 (N_5050,N_3133,N_2426);
or U5051 (N_5051,N_2843,N_2561);
nor U5052 (N_5052,N_2072,N_3768);
and U5053 (N_5053,N_2624,N_2257);
nand U5054 (N_5054,N_2094,N_3484);
nor U5055 (N_5055,N_2641,N_2533);
or U5056 (N_5056,N_2315,N_2778);
nor U5057 (N_5057,N_2325,N_3705);
and U5058 (N_5058,N_2702,N_2016);
or U5059 (N_5059,N_2692,N_2994);
or U5060 (N_5060,N_3636,N_3115);
and U5061 (N_5061,N_2886,N_2432);
nor U5062 (N_5062,N_2718,N_2287);
or U5063 (N_5063,N_2387,N_3829);
or U5064 (N_5064,N_2952,N_3956);
and U5065 (N_5065,N_2047,N_2290);
nand U5066 (N_5066,N_2603,N_2849);
and U5067 (N_5067,N_3130,N_2857);
nor U5068 (N_5068,N_3550,N_2468);
or U5069 (N_5069,N_3390,N_2039);
nand U5070 (N_5070,N_3326,N_2843);
nand U5071 (N_5071,N_3202,N_2741);
or U5072 (N_5072,N_3491,N_3257);
and U5073 (N_5073,N_2618,N_2153);
or U5074 (N_5074,N_3091,N_3230);
or U5075 (N_5075,N_3973,N_2059);
nor U5076 (N_5076,N_2955,N_2653);
nor U5077 (N_5077,N_3422,N_2619);
nand U5078 (N_5078,N_3642,N_3993);
nor U5079 (N_5079,N_2722,N_3336);
and U5080 (N_5080,N_2744,N_3770);
or U5081 (N_5081,N_2986,N_2979);
nor U5082 (N_5082,N_3441,N_2953);
nand U5083 (N_5083,N_3685,N_3642);
and U5084 (N_5084,N_3544,N_3357);
xnor U5085 (N_5085,N_3286,N_3439);
or U5086 (N_5086,N_2728,N_2729);
and U5087 (N_5087,N_2110,N_3897);
nand U5088 (N_5088,N_3018,N_3843);
or U5089 (N_5089,N_2505,N_3028);
and U5090 (N_5090,N_2855,N_3624);
and U5091 (N_5091,N_3294,N_3980);
or U5092 (N_5092,N_2736,N_3014);
nor U5093 (N_5093,N_3988,N_3612);
nor U5094 (N_5094,N_3344,N_3164);
nand U5095 (N_5095,N_2747,N_3373);
nor U5096 (N_5096,N_2965,N_3928);
and U5097 (N_5097,N_3996,N_2468);
nand U5098 (N_5098,N_3249,N_3267);
nand U5099 (N_5099,N_2415,N_3717);
nor U5100 (N_5100,N_2058,N_2086);
nor U5101 (N_5101,N_3119,N_3215);
or U5102 (N_5102,N_3114,N_2646);
xor U5103 (N_5103,N_2306,N_3173);
and U5104 (N_5104,N_3007,N_3682);
and U5105 (N_5105,N_2486,N_2215);
nand U5106 (N_5106,N_2298,N_2418);
and U5107 (N_5107,N_2347,N_3270);
nand U5108 (N_5108,N_3118,N_3082);
nand U5109 (N_5109,N_2011,N_3949);
and U5110 (N_5110,N_2645,N_3347);
and U5111 (N_5111,N_2261,N_2587);
nor U5112 (N_5112,N_2174,N_3863);
nand U5113 (N_5113,N_3748,N_2397);
nor U5114 (N_5114,N_2987,N_2889);
and U5115 (N_5115,N_2345,N_2418);
and U5116 (N_5116,N_2915,N_2039);
nor U5117 (N_5117,N_2765,N_2724);
and U5118 (N_5118,N_3922,N_2280);
nand U5119 (N_5119,N_3919,N_2367);
nand U5120 (N_5120,N_2151,N_2765);
nand U5121 (N_5121,N_2204,N_3761);
xnor U5122 (N_5122,N_2786,N_2149);
or U5123 (N_5123,N_3016,N_2694);
and U5124 (N_5124,N_2531,N_2342);
and U5125 (N_5125,N_3898,N_2611);
or U5126 (N_5126,N_3118,N_2425);
and U5127 (N_5127,N_2680,N_2480);
and U5128 (N_5128,N_2211,N_2085);
and U5129 (N_5129,N_2919,N_3650);
nand U5130 (N_5130,N_2877,N_2592);
or U5131 (N_5131,N_2593,N_2529);
nand U5132 (N_5132,N_2146,N_3234);
nand U5133 (N_5133,N_2492,N_2713);
or U5134 (N_5134,N_2193,N_2163);
nand U5135 (N_5135,N_3074,N_2997);
nand U5136 (N_5136,N_2161,N_3005);
nor U5137 (N_5137,N_2552,N_2251);
and U5138 (N_5138,N_2481,N_3574);
nand U5139 (N_5139,N_2170,N_2461);
nand U5140 (N_5140,N_2733,N_2929);
and U5141 (N_5141,N_2939,N_3387);
nand U5142 (N_5142,N_3961,N_2545);
nand U5143 (N_5143,N_3755,N_3185);
nor U5144 (N_5144,N_3410,N_3988);
nor U5145 (N_5145,N_3604,N_2159);
nand U5146 (N_5146,N_3224,N_3482);
and U5147 (N_5147,N_3102,N_2570);
nand U5148 (N_5148,N_3088,N_2427);
or U5149 (N_5149,N_3018,N_2025);
or U5150 (N_5150,N_2133,N_3453);
nand U5151 (N_5151,N_3868,N_3467);
nand U5152 (N_5152,N_3498,N_3590);
and U5153 (N_5153,N_2969,N_3991);
or U5154 (N_5154,N_3223,N_2206);
nor U5155 (N_5155,N_3199,N_3948);
nor U5156 (N_5156,N_3510,N_2905);
and U5157 (N_5157,N_2998,N_3213);
nand U5158 (N_5158,N_3773,N_3138);
nor U5159 (N_5159,N_2310,N_2108);
nand U5160 (N_5160,N_3556,N_3340);
nand U5161 (N_5161,N_2221,N_3444);
and U5162 (N_5162,N_3202,N_3674);
and U5163 (N_5163,N_2380,N_2686);
nor U5164 (N_5164,N_2551,N_2055);
or U5165 (N_5165,N_3724,N_2387);
and U5166 (N_5166,N_3226,N_3507);
nor U5167 (N_5167,N_2003,N_2424);
nand U5168 (N_5168,N_3527,N_2210);
nor U5169 (N_5169,N_2290,N_2173);
nand U5170 (N_5170,N_3126,N_2703);
or U5171 (N_5171,N_3222,N_3789);
or U5172 (N_5172,N_3326,N_2105);
nor U5173 (N_5173,N_2072,N_2624);
and U5174 (N_5174,N_2695,N_2064);
nor U5175 (N_5175,N_3973,N_3819);
xnor U5176 (N_5176,N_3857,N_3259);
or U5177 (N_5177,N_2760,N_3513);
and U5178 (N_5178,N_3781,N_2506);
nor U5179 (N_5179,N_3255,N_2203);
or U5180 (N_5180,N_2876,N_2960);
or U5181 (N_5181,N_3008,N_2854);
and U5182 (N_5182,N_2815,N_3956);
nor U5183 (N_5183,N_2899,N_3257);
nand U5184 (N_5184,N_2836,N_3965);
nor U5185 (N_5185,N_3252,N_3329);
and U5186 (N_5186,N_3442,N_2170);
and U5187 (N_5187,N_3349,N_3814);
nor U5188 (N_5188,N_2624,N_3314);
and U5189 (N_5189,N_2680,N_3628);
or U5190 (N_5190,N_3996,N_3176);
and U5191 (N_5191,N_2150,N_3536);
nand U5192 (N_5192,N_3861,N_2266);
and U5193 (N_5193,N_2349,N_2460);
or U5194 (N_5194,N_2985,N_3876);
nand U5195 (N_5195,N_2219,N_3297);
nor U5196 (N_5196,N_2760,N_2546);
or U5197 (N_5197,N_3624,N_3967);
and U5198 (N_5198,N_3734,N_3798);
or U5199 (N_5199,N_2860,N_3263);
nand U5200 (N_5200,N_2342,N_3378);
nor U5201 (N_5201,N_2737,N_2504);
and U5202 (N_5202,N_3111,N_3198);
nand U5203 (N_5203,N_3181,N_3014);
and U5204 (N_5204,N_2777,N_3391);
nor U5205 (N_5205,N_2863,N_3272);
nand U5206 (N_5206,N_2079,N_3414);
or U5207 (N_5207,N_2462,N_3316);
or U5208 (N_5208,N_3137,N_3220);
or U5209 (N_5209,N_3438,N_3384);
or U5210 (N_5210,N_3369,N_3743);
and U5211 (N_5211,N_2461,N_3052);
nand U5212 (N_5212,N_2346,N_2449);
nor U5213 (N_5213,N_3140,N_3921);
xnor U5214 (N_5214,N_2073,N_2860);
and U5215 (N_5215,N_3341,N_3584);
nand U5216 (N_5216,N_3349,N_2716);
or U5217 (N_5217,N_2229,N_2793);
nor U5218 (N_5218,N_3814,N_3913);
or U5219 (N_5219,N_2858,N_2848);
or U5220 (N_5220,N_3683,N_3612);
nor U5221 (N_5221,N_2306,N_3910);
nor U5222 (N_5222,N_3006,N_2653);
nor U5223 (N_5223,N_3840,N_2310);
xnor U5224 (N_5224,N_3748,N_3011);
or U5225 (N_5225,N_3023,N_3668);
nor U5226 (N_5226,N_3435,N_3750);
and U5227 (N_5227,N_3037,N_2582);
nor U5228 (N_5228,N_3747,N_2002);
and U5229 (N_5229,N_3766,N_2976);
and U5230 (N_5230,N_3933,N_3159);
nand U5231 (N_5231,N_3744,N_2474);
and U5232 (N_5232,N_3701,N_2023);
nand U5233 (N_5233,N_2658,N_2696);
or U5234 (N_5234,N_3669,N_3021);
or U5235 (N_5235,N_2696,N_3451);
and U5236 (N_5236,N_2235,N_3393);
nor U5237 (N_5237,N_2500,N_3816);
nor U5238 (N_5238,N_3638,N_2806);
nand U5239 (N_5239,N_2042,N_3927);
and U5240 (N_5240,N_2000,N_2463);
or U5241 (N_5241,N_2125,N_3965);
nor U5242 (N_5242,N_2421,N_3707);
xor U5243 (N_5243,N_3536,N_2306);
nand U5244 (N_5244,N_2942,N_2414);
and U5245 (N_5245,N_2569,N_2874);
and U5246 (N_5246,N_2853,N_3027);
and U5247 (N_5247,N_3238,N_2611);
nand U5248 (N_5248,N_2385,N_3924);
or U5249 (N_5249,N_3493,N_3479);
nand U5250 (N_5250,N_2933,N_2676);
nor U5251 (N_5251,N_3500,N_2501);
nand U5252 (N_5252,N_2384,N_3605);
and U5253 (N_5253,N_3213,N_2624);
nor U5254 (N_5254,N_2385,N_3579);
nor U5255 (N_5255,N_2985,N_3154);
nand U5256 (N_5256,N_2170,N_2029);
nand U5257 (N_5257,N_2729,N_3675);
and U5258 (N_5258,N_2849,N_2720);
and U5259 (N_5259,N_2926,N_3146);
nor U5260 (N_5260,N_3169,N_3599);
and U5261 (N_5261,N_2016,N_2448);
nand U5262 (N_5262,N_2684,N_2351);
nor U5263 (N_5263,N_3335,N_2082);
nor U5264 (N_5264,N_2163,N_3261);
xnor U5265 (N_5265,N_3212,N_3694);
or U5266 (N_5266,N_2287,N_2072);
and U5267 (N_5267,N_2792,N_3091);
and U5268 (N_5268,N_2398,N_3634);
or U5269 (N_5269,N_3509,N_3844);
nand U5270 (N_5270,N_2435,N_3047);
nand U5271 (N_5271,N_2522,N_2085);
or U5272 (N_5272,N_2089,N_3372);
or U5273 (N_5273,N_2824,N_3610);
nand U5274 (N_5274,N_3343,N_2844);
or U5275 (N_5275,N_2804,N_3851);
and U5276 (N_5276,N_2043,N_2091);
nor U5277 (N_5277,N_3865,N_3378);
nor U5278 (N_5278,N_2198,N_2878);
or U5279 (N_5279,N_2882,N_2212);
and U5280 (N_5280,N_2620,N_2213);
and U5281 (N_5281,N_2882,N_2631);
nor U5282 (N_5282,N_3049,N_2756);
and U5283 (N_5283,N_3468,N_2698);
and U5284 (N_5284,N_3251,N_2218);
nand U5285 (N_5285,N_2836,N_3103);
nand U5286 (N_5286,N_2055,N_2489);
nand U5287 (N_5287,N_3301,N_3097);
or U5288 (N_5288,N_3325,N_2015);
and U5289 (N_5289,N_3534,N_2278);
nor U5290 (N_5290,N_2356,N_2311);
or U5291 (N_5291,N_2059,N_2850);
or U5292 (N_5292,N_2871,N_2663);
nor U5293 (N_5293,N_3929,N_3795);
and U5294 (N_5294,N_3342,N_3842);
and U5295 (N_5295,N_2716,N_2648);
or U5296 (N_5296,N_2492,N_2284);
or U5297 (N_5297,N_2740,N_2372);
nor U5298 (N_5298,N_2195,N_2273);
or U5299 (N_5299,N_2608,N_3336);
and U5300 (N_5300,N_3631,N_2615);
and U5301 (N_5301,N_3422,N_3295);
or U5302 (N_5302,N_3533,N_2238);
nand U5303 (N_5303,N_2938,N_3361);
and U5304 (N_5304,N_3627,N_2816);
nor U5305 (N_5305,N_2022,N_2049);
nand U5306 (N_5306,N_2475,N_3889);
xor U5307 (N_5307,N_3218,N_2032);
nand U5308 (N_5308,N_2491,N_2742);
nor U5309 (N_5309,N_3762,N_2215);
and U5310 (N_5310,N_3429,N_3363);
nand U5311 (N_5311,N_2144,N_3292);
and U5312 (N_5312,N_3061,N_2193);
xor U5313 (N_5313,N_2115,N_3198);
nor U5314 (N_5314,N_2546,N_2356);
nor U5315 (N_5315,N_3485,N_3799);
and U5316 (N_5316,N_2451,N_2972);
xor U5317 (N_5317,N_2002,N_3337);
and U5318 (N_5318,N_2343,N_3109);
and U5319 (N_5319,N_3847,N_2724);
nand U5320 (N_5320,N_2598,N_2829);
nand U5321 (N_5321,N_3398,N_3425);
or U5322 (N_5322,N_2208,N_3422);
nor U5323 (N_5323,N_2971,N_2991);
nand U5324 (N_5324,N_2078,N_3456);
or U5325 (N_5325,N_2504,N_2976);
or U5326 (N_5326,N_3312,N_3890);
and U5327 (N_5327,N_3643,N_2983);
and U5328 (N_5328,N_2388,N_3345);
nand U5329 (N_5329,N_2423,N_3597);
and U5330 (N_5330,N_2191,N_2199);
xor U5331 (N_5331,N_2881,N_2936);
nand U5332 (N_5332,N_2482,N_2962);
or U5333 (N_5333,N_2385,N_3747);
or U5334 (N_5334,N_3754,N_3846);
or U5335 (N_5335,N_2048,N_3126);
nor U5336 (N_5336,N_3075,N_2004);
nor U5337 (N_5337,N_3349,N_3489);
nor U5338 (N_5338,N_3074,N_3261);
nor U5339 (N_5339,N_3521,N_3232);
or U5340 (N_5340,N_3552,N_2465);
nand U5341 (N_5341,N_2253,N_2303);
and U5342 (N_5342,N_3201,N_2089);
nand U5343 (N_5343,N_3904,N_2994);
nor U5344 (N_5344,N_3234,N_3094);
and U5345 (N_5345,N_3067,N_3473);
nor U5346 (N_5346,N_3345,N_2118);
or U5347 (N_5347,N_3042,N_2188);
nand U5348 (N_5348,N_3720,N_3090);
and U5349 (N_5349,N_3351,N_3635);
and U5350 (N_5350,N_2009,N_3294);
and U5351 (N_5351,N_3667,N_3943);
and U5352 (N_5352,N_3498,N_2316);
nand U5353 (N_5353,N_3229,N_2047);
and U5354 (N_5354,N_3602,N_2945);
nand U5355 (N_5355,N_3884,N_2730);
or U5356 (N_5356,N_3377,N_2567);
and U5357 (N_5357,N_3158,N_2734);
nor U5358 (N_5358,N_2129,N_3537);
and U5359 (N_5359,N_2176,N_3321);
and U5360 (N_5360,N_2024,N_2101);
and U5361 (N_5361,N_2707,N_2999);
nand U5362 (N_5362,N_2559,N_3451);
nand U5363 (N_5363,N_3406,N_3017);
xor U5364 (N_5364,N_3946,N_2918);
or U5365 (N_5365,N_3232,N_2740);
or U5366 (N_5366,N_2906,N_2084);
xor U5367 (N_5367,N_2993,N_2042);
nand U5368 (N_5368,N_2406,N_2277);
and U5369 (N_5369,N_2494,N_3379);
nor U5370 (N_5370,N_2274,N_2183);
and U5371 (N_5371,N_3777,N_3820);
xnor U5372 (N_5372,N_2521,N_2725);
nand U5373 (N_5373,N_2261,N_2523);
nand U5374 (N_5374,N_3398,N_3150);
nand U5375 (N_5375,N_2340,N_2754);
nand U5376 (N_5376,N_2207,N_3136);
or U5377 (N_5377,N_3242,N_3517);
and U5378 (N_5378,N_3239,N_3187);
or U5379 (N_5379,N_3638,N_2927);
or U5380 (N_5380,N_3825,N_2408);
nor U5381 (N_5381,N_2252,N_2103);
nand U5382 (N_5382,N_3677,N_3165);
or U5383 (N_5383,N_3670,N_2046);
and U5384 (N_5384,N_3918,N_3674);
and U5385 (N_5385,N_2332,N_2013);
and U5386 (N_5386,N_3709,N_2605);
nor U5387 (N_5387,N_3253,N_3502);
nor U5388 (N_5388,N_3794,N_3008);
and U5389 (N_5389,N_2389,N_3946);
or U5390 (N_5390,N_3126,N_3546);
nor U5391 (N_5391,N_3668,N_2958);
nand U5392 (N_5392,N_2046,N_3931);
and U5393 (N_5393,N_2408,N_2529);
and U5394 (N_5394,N_2619,N_2579);
or U5395 (N_5395,N_3903,N_3751);
and U5396 (N_5396,N_2394,N_3376);
nor U5397 (N_5397,N_2953,N_3557);
nand U5398 (N_5398,N_3221,N_3565);
nand U5399 (N_5399,N_2380,N_2715);
nand U5400 (N_5400,N_2308,N_3363);
nor U5401 (N_5401,N_2237,N_3414);
nor U5402 (N_5402,N_2131,N_3847);
or U5403 (N_5403,N_2327,N_2460);
and U5404 (N_5404,N_2774,N_3750);
nand U5405 (N_5405,N_3361,N_3358);
nor U5406 (N_5406,N_3330,N_3275);
nand U5407 (N_5407,N_2481,N_2092);
nor U5408 (N_5408,N_3642,N_3422);
nand U5409 (N_5409,N_2176,N_2242);
nand U5410 (N_5410,N_3992,N_2304);
or U5411 (N_5411,N_3146,N_2960);
or U5412 (N_5412,N_2162,N_2958);
nand U5413 (N_5413,N_3568,N_2605);
nand U5414 (N_5414,N_2902,N_3693);
or U5415 (N_5415,N_3905,N_2888);
xor U5416 (N_5416,N_3108,N_3599);
and U5417 (N_5417,N_3326,N_3737);
nand U5418 (N_5418,N_2401,N_2413);
nor U5419 (N_5419,N_2648,N_3038);
or U5420 (N_5420,N_2905,N_2108);
and U5421 (N_5421,N_2368,N_2479);
nand U5422 (N_5422,N_3763,N_3074);
nand U5423 (N_5423,N_3496,N_3103);
or U5424 (N_5424,N_3836,N_3355);
and U5425 (N_5425,N_3123,N_2603);
and U5426 (N_5426,N_3099,N_3155);
nand U5427 (N_5427,N_2429,N_2693);
or U5428 (N_5428,N_3712,N_2854);
nor U5429 (N_5429,N_2536,N_2377);
or U5430 (N_5430,N_3044,N_3264);
and U5431 (N_5431,N_2942,N_2929);
or U5432 (N_5432,N_2063,N_3795);
nor U5433 (N_5433,N_3179,N_3709);
nor U5434 (N_5434,N_3303,N_2233);
nor U5435 (N_5435,N_3483,N_2019);
or U5436 (N_5436,N_3044,N_3737);
nand U5437 (N_5437,N_2288,N_2763);
nand U5438 (N_5438,N_2912,N_3692);
nor U5439 (N_5439,N_2392,N_2490);
or U5440 (N_5440,N_3103,N_2702);
and U5441 (N_5441,N_3502,N_3263);
or U5442 (N_5442,N_2737,N_3321);
nand U5443 (N_5443,N_2259,N_3824);
or U5444 (N_5444,N_2245,N_2859);
and U5445 (N_5445,N_2599,N_3333);
nand U5446 (N_5446,N_2594,N_3788);
or U5447 (N_5447,N_2748,N_2455);
or U5448 (N_5448,N_3264,N_2228);
nor U5449 (N_5449,N_3328,N_2555);
nor U5450 (N_5450,N_2714,N_2000);
nand U5451 (N_5451,N_2176,N_2746);
nand U5452 (N_5452,N_2042,N_3793);
nor U5453 (N_5453,N_3667,N_2055);
nand U5454 (N_5454,N_3973,N_3031);
and U5455 (N_5455,N_3753,N_3776);
and U5456 (N_5456,N_2777,N_3995);
nand U5457 (N_5457,N_2997,N_2247);
and U5458 (N_5458,N_2558,N_3191);
or U5459 (N_5459,N_2679,N_3152);
or U5460 (N_5460,N_2294,N_2453);
nor U5461 (N_5461,N_3879,N_3734);
or U5462 (N_5462,N_3775,N_2892);
and U5463 (N_5463,N_3176,N_2380);
and U5464 (N_5464,N_3147,N_3789);
nor U5465 (N_5465,N_3699,N_2735);
and U5466 (N_5466,N_3667,N_3570);
nand U5467 (N_5467,N_3653,N_3662);
or U5468 (N_5468,N_3819,N_3701);
nor U5469 (N_5469,N_2950,N_2527);
nand U5470 (N_5470,N_2617,N_3990);
and U5471 (N_5471,N_2632,N_3392);
and U5472 (N_5472,N_2582,N_3636);
and U5473 (N_5473,N_3892,N_3782);
or U5474 (N_5474,N_3110,N_3849);
or U5475 (N_5475,N_2218,N_3206);
and U5476 (N_5476,N_3822,N_3616);
or U5477 (N_5477,N_2520,N_3062);
and U5478 (N_5478,N_2031,N_3363);
or U5479 (N_5479,N_3573,N_3870);
nor U5480 (N_5480,N_2486,N_2870);
nand U5481 (N_5481,N_3062,N_2758);
nand U5482 (N_5482,N_3206,N_2626);
nor U5483 (N_5483,N_2755,N_3343);
or U5484 (N_5484,N_3224,N_2402);
nor U5485 (N_5485,N_3706,N_3270);
or U5486 (N_5486,N_3937,N_3430);
and U5487 (N_5487,N_3374,N_3905);
nand U5488 (N_5488,N_2322,N_3541);
nor U5489 (N_5489,N_2351,N_2368);
and U5490 (N_5490,N_2230,N_2066);
and U5491 (N_5491,N_3196,N_3176);
nand U5492 (N_5492,N_2401,N_3577);
nand U5493 (N_5493,N_2555,N_2970);
and U5494 (N_5494,N_2909,N_2099);
nor U5495 (N_5495,N_2403,N_3922);
nor U5496 (N_5496,N_2770,N_3505);
or U5497 (N_5497,N_2335,N_2435);
and U5498 (N_5498,N_2663,N_2661);
nand U5499 (N_5499,N_3602,N_2683);
nor U5500 (N_5500,N_3706,N_3212);
or U5501 (N_5501,N_3426,N_3375);
and U5502 (N_5502,N_2004,N_3924);
nor U5503 (N_5503,N_3754,N_3658);
nand U5504 (N_5504,N_3535,N_2288);
and U5505 (N_5505,N_2722,N_3648);
and U5506 (N_5506,N_3214,N_2173);
and U5507 (N_5507,N_2087,N_2025);
or U5508 (N_5508,N_2746,N_2204);
or U5509 (N_5509,N_3124,N_2575);
or U5510 (N_5510,N_2786,N_2268);
nor U5511 (N_5511,N_3715,N_3029);
nand U5512 (N_5512,N_3317,N_3706);
and U5513 (N_5513,N_3771,N_3572);
and U5514 (N_5514,N_2416,N_2985);
nand U5515 (N_5515,N_3132,N_3176);
nor U5516 (N_5516,N_3817,N_3482);
nor U5517 (N_5517,N_2437,N_3304);
and U5518 (N_5518,N_3431,N_2111);
or U5519 (N_5519,N_2692,N_3422);
nand U5520 (N_5520,N_2937,N_3255);
or U5521 (N_5521,N_2759,N_3036);
and U5522 (N_5522,N_2786,N_3618);
nand U5523 (N_5523,N_3147,N_3994);
nand U5524 (N_5524,N_3568,N_3880);
or U5525 (N_5525,N_2279,N_2842);
and U5526 (N_5526,N_3986,N_2458);
nor U5527 (N_5527,N_3091,N_2454);
and U5528 (N_5528,N_3662,N_3142);
nand U5529 (N_5529,N_3643,N_2504);
or U5530 (N_5530,N_3352,N_2704);
nor U5531 (N_5531,N_2947,N_2389);
and U5532 (N_5532,N_2561,N_2373);
and U5533 (N_5533,N_2464,N_3024);
nand U5534 (N_5534,N_2051,N_2319);
nand U5535 (N_5535,N_3967,N_2193);
nand U5536 (N_5536,N_2160,N_3108);
nand U5537 (N_5537,N_3345,N_2004);
nand U5538 (N_5538,N_2740,N_3982);
nor U5539 (N_5539,N_2146,N_3878);
nor U5540 (N_5540,N_2985,N_2930);
and U5541 (N_5541,N_2323,N_3111);
nand U5542 (N_5542,N_2567,N_2212);
nand U5543 (N_5543,N_2249,N_3673);
and U5544 (N_5544,N_2781,N_3314);
or U5545 (N_5545,N_3518,N_2601);
nand U5546 (N_5546,N_3883,N_2857);
and U5547 (N_5547,N_3390,N_2920);
and U5548 (N_5548,N_2859,N_2026);
or U5549 (N_5549,N_2152,N_2713);
nor U5550 (N_5550,N_2288,N_2692);
or U5551 (N_5551,N_3705,N_3961);
nand U5552 (N_5552,N_2693,N_2588);
nand U5553 (N_5553,N_3144,N_2934);
nand U5554 (N_5554,N_2706,N_3911);
nand U5555 (N_5555,N_3082,N_3979);
nand U5556 (N_5556,N_3817,N_2794);
or U5557 (N_5557,N_3987,N_3171);
and U5558 (N_5558,N_3827,N_3139);
and U5559 (N_5559,N_2030,N_3761);
or U5560 (N_5560,N_2350,N_2715);
nand U5561 (N_5561,N_2027,N_3009);
or U5562 (N_5562,N_3094,N_2419);
or U5563 (N_5563,N_2812,N_3421);
xnor U5564 (N_5564,N_3670,N_2847);
or U5565 (N_5565,N_2294,N_2852);
or U5566 (N_5566,N_2835,N_3643);
nand U5567 (N_5567,N_3311,N_3624);
or U5568 (N_5568,N_3113,N_3778);
nor U5569 (N_5569,N_3240,N_2055);
nand U5570 (N_5570,N_3624,N_3022);
or U5571 (N_5571,N_2342,N_3048);
nand U5572 (N_5572,N_2946,N_3415);
nor U5573 (N_5573,N_3621,N_2758);
nand U5574 (N_5574,N_3379,N_2626);
nand U5575 (N_5575,N_2137,N_3234);
nor U5576 (N_5576,N_3262,N_2953);
or U5577 (N_5577,N_2519,N_2309);
xor U5578 (N_5578,N_2779,N_2464);
xor U5579 (N_5579,N_2860,N_3330);
nand U5580 (N_5580,N_2280,N_3229);
nand U5581 (N_5581,N_3121,N_3609);
nor U5582 (N_5582,N_2189,N_2248);
nor U5583 (N_5583,N_2201,N_2799);
or U5584 (N_5584,N_3826,N_3609);
or U5585 (N_5585,N_2118,N_2117);
and U5586 (N_5586,N_2366,N_3836);
nand U5587 (N_5587,N_2045,N_3700);
nor U5588 (N_5588,N_3882,N_2491);
or U5589 (N_5589,N_2637,N_3514);
or U5590 (N_5590,N_2404,N_3430);
and U5591 (N_5591,N_2182,N_2125);
nor U5592 (N_5592,N_3027,N_2747);
nor U5593 (N_5593,N_3212,N_3553);
nor U5594 (N_5594,N_2569,N_2941);
or U5595 (N_5595,N_2343,N_2102);
nor U5596 (N_5596,N_3239,N_3211);
nand U5597 (N_5597,N_3636,N_3536);
or U5598 (N_5598,N_2007,N_2806);
or U5599 (N_5599,N_2912,N_3514);
nor U5600 (N_5600,N_2813,N_3781);
nor U5601 (N_5601,N_3372,N_3816);
or U5602 (N_5602,N_3446,N_2808);
and U5603 (N_5603,N_3147,N_2917);
and U5604 (N_5604,N_2963,N_2551);
and U5605 (N_5605,N_2816,N_2383);
and U5606 (N_5606,N_2490,N_2887);
and U5607 (N_5607,N_3568,N_2824);
and U5608 (N_5608,N_3608,N_2604);
and U5609 (N_5609,N_3962,N_2847);
nand U5610 (N_5610,N_3606,N_2425);
nor U5611 (N_5611,N_2825,N_3739);
or U5612 (N_5612,N_2987,N_2649);
nor U5613 (N_5613,N_3488,N_2088);
xor U5614 (N_5614,N_3744,N_3996);
or U5615 (N_5615,N_2880,N_2664);
and U5616 (N_5616,N_3575,N_3988);
or U5617 (N_5617,N_2110,N_3324);
nand U5618 (N_5618,N_2366,N_3714);
and U5619 (N_5619,N_2389,N_3554);
and U5620 (N_5620,N_2165,N_3188);
nand U5621 (N_5621,N_3511,N_2381);
nor U5622 (N_5622,N_3258,N_2469);
nand U5623 (N_5623,N_2951,N_3550);
nand U5624 (N_5624,N_3541,N_3599);
or U5625 (N_5625,N_2465,N_3011);
nand U5626 (N_5626,N_3452,N_2250);
and U5627 (N_5627,N_3759,N_2638);
nand U5628 (N_5628,N_2758,N_2850);
nor U5629 (N_5629,N_3979,N_2662);
nor U5630 (N_5630,N_2662,N_2019);
nand U5631 (N_5631,N_2983,N_3025);
nand U5632 (N_5632,N_3414,N_3344);
nand U5633 (N_5633,N_3272,N_2336);
or U5634 (N_5634,N_3303,N_2875);
and U5635 (N_5635,N_3603,N_3361);
and U5636 (N_5636,N_3444,N_2040);
nand U5637 (N_5637,N_3527,N_3120);
nand U5638 (N_5638,N_3139,N_2208);
or U5639 (N_5639,N_2815,N_2573);
and U5640 (N_5640,N_3200,N_3386);
nand U5641 (N_5641,N_2965,N_2156);
or U5642 (N_5642,N_2849,N_3333);
and U5643 (N_5643,N_3015,N_2800);
and U5644 (N_5644,N_2864,N_3017);
nand U5645 (N_5645,N_2655,N_3342);
and U5646 (N_5646,N_3863,N_3858);
or U5647 (N_5647,N_3918,N_2680);
and U5648 (N_5648,N_3291,N_2527);
nor U5649 (N_5649,N_3012,N_2288);
nand U5650 (N_5650,N_2116,N_3698);
or U5651 (N_5651,N_2729,N_3078);
and U5652 (N_5652,N_3363,N_3244);
and U5653 (N_5653,N_2039,N_2527);
and U5654 (N_5654,N_2875,N_2028);
nand U5655 (N_5655,N_3729,N_2281);
or U5656 (N_5656,N_3212,N_3504);
nand U5657 (N_5657,N_2961,N_2535);
nand U5658 (N_5658,N_3734,N_2970);
and U5659 (N_5659,N_3330,N_2790);
nand U5660 (N_5660,N_2379,N_3732);
and U5661 (N_5661,N_3017,N_3559);
nand U5662 (N_5662,N_3973,N_3307);
nor U5663 (N_5663,N_3624,N_3308);
or U5664 (N_5664,N_3088,N_3998);
and U5665 (N_5665,N_3560,N_3054);
nor U5666 (N_5666,N_3394,N_3051);
and U5667 (N_5667,N_2197,N_3376);
or U5668 (N_5668,N_2988,N_3716);
and U5669 (N_5669,N_3004,N_3709);
and U5670 (N_5670,N_2037,N_2812);
nor U5671 (N_5671,N_2791,N_2283);
nor U5672 (N_5672,N_2537,N_2656);
or U5673 (N_5673,N_3572,N_2294);
nand U5674 (N_5674,N_2104,N_2491);
nand U5675 (N_5675,N_2994,N_2364);
and U5676 (N_5676,N_2880,N_2262);
or U5677 (N_5677,N_2299,N_2332);
and U5678 (N_5678,N_3640,N_2307);
nand U5679 (N_5679,N_2742,N_3108);
and U5680 (N_5680,N_2463,N_2523);
and U5681 (N_5681,N_3462,N_2885);
nor U5682 (N_5682,N_2980,N_3587);
and U5683 (N_5683,N_2194,N_3718);
nand U5684 (N_5684,N_2282,N_2575);
nand U5685 (N_5685,N_2548,N_2928);
and U5686 (N_5686,N_2931,N_2546);
and U5687 (N_5687,N_2239,N_2517);
or U5688 (N_5688,N_3572,N_2362);
or U5689 (N_5689,N_2681,N_3496);
or U5690 (N_5690,N_3771,N_2734);
or U5691 (N_5691,N_2509,N_3644);
nor U5692 (N_5692,N_3399,N_3461);
nand U5693 (N_5693,N_2017,N_3569);
nand U5694 (N_5694,N_2502,N_2336);
or U5695 (N_5695,N_2029,N_3624);
and U5696 (N_5696,N_3878,N_2225);
nor U5697 (N_5697,N_3152,N_3421);
and U5698 (N_5698,N_3276,N_3792);
nor U5699 (N_5699,N_3891,N_2773);
nor U5700 (N_5700,N_3486,N_2316);
nor U5701 (N_5701,N_2430,N_2067);
and U5702 (N_5702,N_3974,N_3350);
nor U5703 (N_5703,N_2886,N_3909);
and U5704 (N_5704,N_2721,N_2436);
nor U5705 (N_5705,N_2885,N_2298);
xor U5706 (N_5706,N_3360,N_2257);
nand U5707 (N_5707,N_3870,N_2945);
and U5708 (N_5708,N_2439,N_2152);
nor U5709 (N_5709,N_3323,N_3157);
and U5710 (N_5710,N_2269,N_3586);
or U5711 (N_5711,N_3779,N_3523);
nor U5712 (N_5712,N_2642,N_3619);
or U5713 (N_5713,N_3965,N_3757);
nand U5714 (N_5714,N_2407,N_2844);
nor U5715 (N_5715,N_2900,N_3131);
or U5716 (N_5716,N_3894,N_2092);
nor U5717 (N_5717,N_2254,N_3413);
or U5718 (N_5718,N_3168,N_3156);
nor U5719 (N_5719,N_3048,N_3129);
and U5720 (N_5720,N_2465,N_2021);
nand U5721 (N_5721,N_3334,N_2298);
or U5722 (N_5722,N_2143,N_2505);
or U5723 (N_5723,N_3996,N_2827);
nor U5724 (N_5724,N_2374,N_3320);
and U5725 (N_5725,N_3495,N_2746);
or U5726 (N_5726,N_2499,N_3794);
nand U5727 (N_5727,N_3869,N_2825);
nor U5728 (N_5728,N_3151,N_2511);
or U5729 (N_5729,N_3262,N_3949);
nand U5730 (N_5730,N_2522,N_2415);
or U5731 (N_5731,N_2569,N_3888);
nor U5732 (N_5732,N_2230,N_2830);
nand U5733 (N_5733,N_3303,N_3731);
and U5734 (N_5734,N_2678,N_3632);
or U5735 (N_5735,N_3160,N_3285);
nor U5736 (N_5736,N_2478,N_2511);
and U5737 (N_5737,N_3324,N_3801);
nor U5738 (N_5738,N_3230,N_2320);
nand U5739 (N_5739,N_2245,N_2839);
or U5740 (N_5740,N_3726,N_2316);
and U5741 (N_5741,N_2290,N_3552);
xnor U5742 (N_5742,N_3128,N_3072);
or U5743 (N_5743,N_3213,N_3793);
or U5744 (N_5744,N_2241,N_3537);
nand U5745 (N_5745,N_2434,N_2056);
and U5746 (N_5746,N_2903,N_3560);
or U5747 (N_5747,N_2580,N_2098);
nand U5748 (N_5748,N_3249,N_2696);
and U5749 (N_5749,N_2479,N_2186);
nand U5750 (N_5750,N_3111,N_2531);
nor U5751 (N_5751,N_3475,N_2728);
and U5752 (N_5752,N_3657,N_3818);
nand U5753 (N_5753,N_2520,N_2337);
and U5754 (N_5754,N_2429,N_2655);
nor U5755 (N_5755,N_2982,N_3018);
nand U5756 (N_5756,N_2387,N_2382);
and U5757 (N_5757,N_3210,N_3752);
and U5758 (N_5758,N_2067,N_3145);
nor U5759 (N_5759,N_3716,N_2042);
and U5760 (N_5760,N_3832,N_3908);
nand U5761 (N_5761,N_3917,N_3898);
nand U5762 (N_5762,N_3117,N_2431);
nand U5763 (N_5763,N_2593,N_2187);
nand U5764 (N_5764,N_3959,N_2474);
and U5765 (N_5765,N_2783,N_3791);
nand U5766 (N_5766,N_3716,N_3727);
nand U5767 (N_5767,N_2372,N_3071);
or U5768 (N_5768,N_3030,N_2047);
nand U5769 (N_5769,N_2087,N_2259);
and U5770 (N_5770,N_2718,N_2663);
nor U5771 (N_5771,N_3311,N_2665);
or U5772 (N_5772,N_3513,N_2914);
nor U5773 (N_5773,N_3721,N_3964);
nor U5774 (N_5774,N_2073,N_3287);
nand U5775 (N_5775,N_2642,N_3187);
or U5776 (N_5776,N_3491,N_3700);
nand U5777 (N_5777,N_3483,N_3475);
and U5778 (N_5778,N_3831,N_2812);
or U5779 (N_5779,N_3015,N_2367);
nand U5780 (N_5780,N_2574,N_3422);
nand U5781 (N_5781,N_2513,N_3157);
nand U5782 (N_5782,N_2150,N_3017);
and U5783 (N_5783,N_3386,N_2346);
and U5784 (N_5784,N_3463,N_3292);
or U5785 (N_5785,N_3433,N_3266);
or U5786 (N_5786,N_2508,N_2812);
nor U5787 (N_5787,N_2724,N_2251);
or U5788 (N_5788,N_3204,N_2357);
or U5789 (N_5789,N_3999,N_3633);
or U5790 (N_5790,N_2850,N_3333);
nand U5791 (N_5791,N_2027,N_3707);
nand U5792 (N_5792,N_3766,N_2591);
or U5793 (N_5793,N_2936,N_2885);
and U5794 (N_5794,N_2261,N_3832);
or U5795 (N_5795,N_2142,N_3584);
or U5796 (N_5796,N_3020,N_3044);
or U5797 (N_5797,N_2632,N_3808);
or U5798 (N_5798,N_3659,N_3929);
and U5799 (N_5799,N_3505,N_2420);
nor U5800 (N_5800,N_3986,N_2363);
nor U5801 (N_5801,N_2609,N_3419);
or U5802 (N_5802,N_2123,N_3650);
and U5803 (N_5803,N_3731,N_3546);
or U5804 (N_5804,N_3276,N_3502);
or U5805 (N_5805,N_3560,N_2683);
and U5806 (N_5806,N_3412,N_2849);
or U5807 (N_5807,N_2526,N_2112);
nor U5808 (N_5808,N_2987,N_2590);
nand U5809 (N_5809,N_2290,N_2612);
or U5810 (N_5810,N_3319,N_2076);
or U5811 (N_5811,N_2404,N_3052);
nor U5812 (N_5812,N_3426,N_3658);
and U5813 (N_5813,N_3542,N_2480);
or U5814 (N_5814,N_2940,N_3374);
or U5815 (N_5815,N_2886,N_3192);
nand U5816 (N_5816,N_3515,N_2011);
xor U5817 (N_5817,N_3849,N_2714);
and U5818 (N_5818,N_3818,N_2524);
nand U5819 (N_5819,N_2911,N_3029);
nand U5820 (N_5820,N_3010,N_2843);
or U5821 (N_5821,N_3120,N_3224);
nand U5822 (N_5822,N_2092,N_2734);
nor U5823 (N_5823,N_2616,N_2832);
and U5824 (N_5824,N_3243,N_3553);
nand U5825 (N_5825,N_2746,N_3585);
nor U5826 (N_5826,N_2563,N_3080);
nor U5827 (N_5827,N_2758,N_3973);
xor U5828 (N_5828,N_2092,N_2559);
nor U5829 (N_5829,N_2315,N_2523);
nor U5830 (N_5830,N_2249,N_2310);
or U5831 (N_5831,N_3888,N_2289);
nor U5832 (N_5832,N_3855,N_2253);
and U5833 (N_5833,N_2020,N_2949);
nand U5834 (N_5834,N_2439,N_2441);
nand U5835 (N_5835,N_3708,N_2571);
or U5836 (N_5836,N_2041,N_2919);
nand U5837 (N_5837,N_2398,N_3012);
or U5838 (N_5838,N_3147,N_2637);
and U5839 (N_5839,N_3239,N_3829);
nand U5840 (N_5840,N_3610,N_3433);
or U5841 (N_5841,N_3073,N_3540);
and U5842 (N_5842,N_2096,N_2868);
nor U5843 (N_5843,N_2250,N_3217);
and U5844 (N_5844,N_3455,N_3257);
or U5845 (N_5845,N_2337,N_3975);
and U5846 (N_5846,N_2175,N_2447);
nor U5847 (N_5847,N_2206,N_2117);
and U5848 (N_5848,N_3612,N_2021);
and U5849 (N_5849,N_2728,N_2025);
or U5850 (N_5850,N_2362,N_3369);
xnor U5851 (N_5851,N_2401,N_3548);
nand U5852 (N_5852,N_3536,N_2342);
or U5853 (N_5853,N_3311,N_2291);
nor U5854 (N_5854,N_2947,N_3940);
nand U5855 (N_5855,N_3627,N_3451);
nand U5856 (N_5856,N_2946,N_2544);
nor U5857 (N_5857,N_2552,N_3364);
or U5858 (N_5858,N_2848,N_3725);
nor U5859 (N_5859,N_3984,N_3655);
or U5860 (N_5860,N_3857,N_2374);
nand U5861 (N_5861,N_3403,N_3072);
or U5862 (N_5862,N_2412,N_3341);
and U5863 (N_5863,N_3908,N_3089);
nand U5864 (N_5864,N_2721,N_3188);
nor U5865 (N_5865,N_2682,N_3516);
or U5866 (N_5866,N_3254,N_2923);
and U5867 (N_5867,N_2386,N_2162);
nor U5868 (N_5868,N_2693,N_3900);
nor U5869 (N_5869,N_3643,N_2077);
and U5870 (N_5870,N_2531,N_3379);
nand U5871 (N_5871,N_3432,N_2795);
nor U5872 (N_5872,N_2228,N_3426);
and U5873 (N_5873,N_2259,N_2849);
nor U5874 (N_5874,N_3072,N_3284);
or U5875 (N_5875,N_2947,N_2593);
nor U5876 (N_5876,N_3965,N_3516);
and U5877 (N_5877,N_3124,N_3560);
and U5878 (N_5878,N_3626,N_3956);
or U5879 (N_5879,N_3584,N_3583);
nor U5880 (N_5880,N_2394,N_3195);
or U5881 (N_5881,N_2760,N_2036);
nor U5882 (N_5882,N_2707,N_3783);
and U5883 (N_5883,N_3769,N_3680);
or U5884 (N_5884,N_2360,N_3025);
and U5885 (N_5885,N_2717,N_2249);
nor U5886 (N_5886,N_2896,N_2546);
and U5887 (N_5887,N_2148,N_2361);
nor U5888 (N_5888,N_3130,N_2300);
and U5889 (N_5889,N_2702,N_3836);
nand U5890 (N_5890,N_3611,N_3654);
nor U5891 (N_5891,N_2853,N_3333);
and U5892 (N_5892,N_3597,N_2395);
and U5893 (N_5893,N_2099,N_2104);
or U5894 (N_5894,N_3957,N_3390);
or U5895 (N_5895,N_2086,N_3973);
nand U5896 (N_5896,N_2083,N_2398);
or U5897 (N_5897,N_3466,N_2355);
and U5898 (N_5898,N_2638,N_2355);
or U5899 (N_5899,N_2414,N_2506);
nor U5900 (N_5900,N_3794,N_2668);
xor U5901 (N_5901,N_3093,N_3037);
nand U5902 (N_5902,N_3965,N_3934);
and U5903 (N_5903,N_2917,N_2302);
nor U5904 (N_5904,N_2155,N_2306);
nand U5905 (N_5905,N_2503,N_3233);
nor U5906 (N_5906,N_2817,N_2631);
nand U5907 (N_5907,N_3874,N_2219);
nand U5908 (N_5908,N_2970,N_2585);
nand U5909 (N_5909,N_3728,N_2164);
nand U5910 (N_5910,N_3695,N_2772);
nor U5911 (N_5911,N_3912,N_2354);
or U5912 (N_5912,N_3583,N_2679);
nor U5913 (N_5913,N_3852,N_3600);
nor U5914 (N_5914,N_2632,N_3370);
or U5915 (N_5915,N_2900,N_2971);
nand U5916 (N_5916,N_2203,N_3411);
nor U5917 (N_5917,N_2201,N_2726);
nor U5918 (N_5918,N_2201,N_3659);
nor U5919 (N_5919,N_3248,N_2528);
nand U5920 (N_5920,N_2011,N_3656);
xnor U5921 (N_5921,N_2906,N_2705);
and U5922 (N_5922,N_3901,N_3501);
nand U5923 (N_5923,N_3345,N_2538);
and U5924 (N_5924,N_2076,N_3044);
nand U5925 (N_5925,N_3068,N_3732);
or U5926 (N_5926,N_3709,N_2835);
or U5927 (N_5927,N_3714,N_2357);
and U5928 (N_5928,N_3498,N_2559);
and U5929 (N_5929,N_2182,N_2586);
or U5930 (N_5930,N_2593,N_3112);
xnor U5931 (N_5931,N_2529,N_3303);
nand U5932 (N_5932,N_3143,N_3825);
or U5933 (N_5933,N_2772,N_3904);
or U5934 (N_5934,N_3171,N_3231);
nand U5935 (N_5935,N_3430,N_3700);
nand U5936 (N_5936,N_3406,N_3469);
or U5937 (N_5937,N_3150,N_3445);
or U5938 (N_5938,N_2805,N_2194);
or U5939 (N_5939,N_2195,N_2342);
nand U5940 (N_5940,N_3281,N_2112);
nand U5941 (N_5941,N_3121,N_3665);
and U5942 (N_5942,N_3924,N_3074);
nor U5943 (N_5943,N_3663,N_3828);
and U5944 (N_5944,N_2322,N_2169);
or U5945 (N_5945,N_2129,N_2254);
nand U5946 (N_5946,N_2153,N_3802);
and U5947 (N_5947,N_3577,N_2105);
nand U5948 (N_5948,N_2673,N_2364);
nand U5949 (N_5949,N_3104,N_2428);
nor U5950 (N_5950,N_2991,N_2550);
or U5951 (N_5951,N_3583,N_2736);
xor U5952 (N_5952,N_3126,N_2434);
and U5953 (N_5953,N_2071,N_3942);
nand U5954 (N_5954,N_3141,N_3816);
and U5955 (N_5955,N_3463,N_3863);
nor U5956 (N_5956,N_3416,N_2866);
nand U5957 (N_5957,N_3041,N_2835);
nand U5958 (N_5958,N_3552,N_3240);
nand U5959 (N_5959,N_2758,N_2143);
nor U5960 (N_5960,N_3666,N_3286);
or U5961 (N_5961,N_2524,N_3009);
or U5962 (N_5962,N_3440,N_2250);
nor U5963 (N_5963,N_2267,N_2740);
and U5964 (N_5964,N_3402,N_3462);
or U5965 (N_5965,N_3732,N_3677);
nand U5966 (N_5966,N_3220,N_3853);
or U5967 (N_5967,N_2758,N_3072);
nand U5968 (N_5968,N_3229,N_3813);
nor U5969 (N_5969,N_2813,N_2275);
nor U5970 (N_5970,N_3389,N_3393);
and U5971 (N_5971,N_3536,N_3974);
or U5972 (N_5972,N_2886,N_2851);
nand U5973 (N_5973,N_3976,N_3798);
or U5974 (N_5974,N_3245,N_2488);
and U5975 (N_5975,N_3230,N_2570);
or U5976 (N_5976,N_3403,N_2648);
and U5977 (N_5977,N_2028,N_2826);
or U5978 (N_5978,N_3407,N_3011);
nand U5979 (N_5979,N_2100,N_3962);
nand U5980 (N_5980,N_3117,N_3017);
nor U5981 (N_5981,N_3173,N_2489);
or U5982 (N_5982,N_2528,N_3313);
or U5983 (N_5983,N_2200,N_3589);
or U5984 (N_5984,N_3796,N_2507);
and U5985 (N_5985,N_3695,N_3645);
or U5986 (N_5986,N_3946,N_3987);
and U5987 (N_5987,N_2329,N_2994);
nand U5988 (N_5988,N_3479,N_2509);
nand U5989 (N_5989,N_2272,N_3192);
and U5990 (N_5990,N_2497,N_2323);
and U5991 (N_5991,N_2477,N_3541);
nand U5992 (N_5992,N_2209,N_3239);
nor U5993 (N_5993,N_2597,N_3780);
or U5994 (N_5994,N_2652,N_3196);
and U5995 (N_5995,N_3355,N_3295);
xor U5996 (N_5996,N_3112,N_2089);
and U5997 (N_5997,N_3574,N_2883);
nand U5998 (N_5998,N_2386,N_3771);
nor U5999 (N_5999,N_2480,N_2608);
nand U6000 (N_6000,N_4316,N_5591);
or U6001 (N_6001,N_4664,N_5632);
or U6002 (N_6002,N_5972,N_4264);
nor U6003 (N_6003,N_5141,N_5287);
nor U6004 (N_6004,N_5703,N_5328);
nor U6005 (N_6005,N_4943,N_4928);
nor U6006 (N_6006,N_5037,N_5534);
nor U6007 (N_6007,N_5362,N_5096);
nor U6008 (N_6008,N_4606,N_5842);
nand U6009 (N_6009,N_5340,N_5263);
nand U6010 (N_6010,N_4378,N_5638);
and U6011 (N_6011,N_4573,N_4416);
and U6012 (N_6012,N_5272,N_5518);
and U6013 (N_6013,N_4476,N_4530);
and U6014 (N_6014,N_4022,N_4569);
and U6015 (N_6015,N_5704,N_5385);
nand U6016 (N_6016,N_4953,N_5364);
or U6017 (N_6017,N_4949,N_5475);
and U6018 (N_6018,N_5554,N_4802);
nor U6019 (N_6019,N_5708,N_4309);
or U6020 (N_6020,N_4874,N_4241);
nor U6021 (N_6021,N_5964,N_5885);
xor U6022 (N_6022,N_4858,N_5610);
or U6023 (N_6023,N_5240,N_5281);
and U6024 (N_6024,N_4009,N_5180);
and U6025 (N_6025,N_4366,N_4691);
and U6026 (N_6026,N_4390,N_4137);
or U6027 (N_6027,N_5779,N_5493);
nand U6028 (N_6028,N_4076,N_5877);
and U6029 (N_6029,N_5365,N_4421);
or U6030 (N_6030,N_4932,N_4427);
nand U6031 (N_6031,N_5593,N_5191);
nand U6032 (N_6032,N_4217,N_4966);
nor U6033 (N_6033,N_4417,N_4302);
and U6034 (N_6034,N_4831,N_4806);
and U6035 (N_6035,N_5501,N_4038);
nor U6036 (N_6036,N_4864,N_5932);
and U6037 (N_6037,N_4556,N_4197);
nand U6038 (N_6038,N_5067,N_5587);
nor U6039 (N_6039,N_4150,N_5622);
nor U6040 (N_6040,N_4653,N_4654);
nand U6041 (N_6041,N_4042,N_5312);
and U6042 (N_6042,N_4168,N_5358);
nor U6043 (N_6043,N_4733,N_5884);
nor U6044 (N_6044,N_5774,N_5941);
nor U6045 (N_6045,N_4105,N_5742);
nor U6046 (N_6046,N_5503,N_5125);
nand U6047 (N_6047,N_4532,N_5929);
or U6048 (N_6048,N_4234,N_4717);
nand U6049 (N_6049,N_4647,N_4188);
and U6050 (N_6050,N_5149,N_4068);
nand U6051 (N_6051,N_4274,N_5369);
nand U6052 (N_6052,N_4273,N_5996);
or U6053 (N_6053,N_5173,N_4946);
nor U6054 (N_6054,N_4290,N_4753);
or U6055 (N_6055,N_4792,N_4616);
or U6056 (N_6056,N_5831,N_5537);
or U6057 (N_6057,N_4544,N_4767);
or U6058 (N_6058,N_4441,N_5854);
and U6059 (N_6059,N_4724,N_4298);
and U6060 (N_6060,N_5551,N_5271);
and U6061 (N_6061,N_4325,N_4773);
and U6062 (N_6062,N_5888,N_4511);
or U6063 (N_6063,N_4071,N_4395);
nand U6064 (N_6064,N_4043,N_4382);
or U6065 (N_6065,N_4936,N_5239);
or U6066 (N_6066,N_5601,N_4013);
or U6067 (N_6067,N_5048,N_5778);
nand U6068 (N_6068,N_5781,N_5716);
nor U6069 (N_6069,N_5089,N_5303);
and U6070 (N_6070,N_5266,N_4296);
nor U6071 (N_6071,N_5504,N_5282);
nand U6072 (N_6072,N_4490,N_4089);
or U6073 (N_6073,N_4930,N_4574);
nand U6074 (N_6074,N_5336,N_5101);
nor U6075 (N_6075,N_5939,N_5615);
and U6076 (N_6076,N_4189,N_4442);
and U6077 (N_6077,N_5562,N_4791);
nor U6078 (N_6078,N_5712,N_4412);
nor U6079 (N_6079,N_5404,N_5407);
nand U6080 (N_6080,N_4823,N_5414);
nand U6081 (N_6081,N_5606,N_4207);
xnor U6082 (N_6082,N_4221,N_4705);
or U6083 (N_6083,N_5944,N_4784);
nand U6084 (N_6084,N_4214,N_5027);
or U6085 (N_6085,N_5188,N_4136);
nand U6086 (N_6086,N_4989,N_5729);
or U6087 (N_6087,N_5157,N_4344);
nand U6088 (N_6088,N_5725,N_4644);
nand U6089 (N_6089,N_5231,N_4045);
or U6090 (N_6090,N_4685,N_5649);
nand U6091 (N_6091,N_4563,N_4340);
nor U6092 (N_6092,N_5249,N_4015);
or U6093 (N_6093,N_5953,N_5875);
and U6094 (N_6094,N_4092,N_5359);
or U6095 (N_6095,N_5900,N_4151);
or U6096 (N_6096,N_5979,N_4121);
nand U6097 (N_6097,N_5498,N_4058);
and U6098 (N_6098,N_5543,N_5317);
nor U6099 (N_6099,N_5784,N_4585);
and U6100 (N_6100,N_5765,N_5019);
and U6101 (N_6101,N_5612,N_4001);
nor U6102 (N_6102,N_4583,N_4553);
nand U6103 (N_6103,N_5442,N_5525);
nor U6104 (N_6104,N_4628,N_4896);
or U6105 (N_6105,N_4633,N_5776);
and U6106 (N_6106,N_5536,N_4179);
or U6107 (N_6107,N_4283,N_4426);
nor U6108 (N_6108,N_5009,N_4999);
or U6109 (N_6109,N_5576,N_5791);
nor U6110 (N_6110,N_5608,N_5481);
nor U6111 (N_6111,N_4997,N_5070);
or U6112 (N_6112,N_5017,N_4438);
nand U6113 (N_6113,N_5627,N_5920);
nor U6114 (N_6114,N_4976,N_4921);
and U6115 (N_6115,N_4774,N_4561);
or U6116 (N_6116,N_4166,N_5198);
nor U6117 (N_6117,N_4675,N_4629);
nor U6118 (N_6118,N_4358,N_4070);
nand U6119 (N_6119,N_5313,N_5144);
or U6120 (N_6120,N_5768,N_5849);
nand U6121 (N_6121,N_5694,N_4782);
nand U6122 (N_6122,N_5243,N_4566);
nand U6123 (N_6123,N_4992,N_4794);
nand U6124 (N_6124,N_4252,N_4766);
and U6125 (N_6125,N_5321,N_4034);
and U6126 (N_6126,N_4762,N_5653);
or U6127 (N_6127,N_5706,N_4745);
and U6128 (N_6128,N_5117,N_4580);
nor U6129 (N_6129,N_5441,N_5203);
nand U6130 (N_6130,N_4429,N_4600);
or U6131 (N_6131,N_4819,N_4191);
nor U6132 (N_6132,N_5458,N_5182);
or U6133 (N_6133,N_5511,N_5128);
nand U6134 (N_6134,N_5547,N_4025);
nand U6135 (N_6135,N_4777,N_4318);
and U6136 (N_6136,N_5714,N_4879);
nor U6137 (N_6137,N_5288,N_5646);
nor U6138 (N_6138,N_4560,N_5056);
nand U6139 (N_6139,N_4176,N_5541);
nand U6140 (N_6140,N_5436,N_4697);
xnor U6141 (N_6141,N_4293,N_5630);
and U6142 (N_6142,N_4353,N_4280);
nand U6143 (N_6143,N_4959,N_5479);
nand U6144 (N_6144,N_4597,N_5254);
nor U6145 (N_6145,N_4641,N_5346);
and U6146 (N_6146,N_4827,N_5566);
nand U6147 (N_6147,N_4002,N_5528);
nand U6148 (N_6148,N_4672,N_5057);
or U6149 (N_6149,N_5812,N_5813);
and U6150 (N_6150,N_5891,N_5505);
nor U6151 (N_6151,N_4699,N_4394);
or U6152 (N_6152,N_5538,N_4251);
nor U6153 (N_6153,N_4098,N_5178);
or U6154 (N_6154,N_5739,N_5931);
and U6155 (N_6155,N_5108,N_4361);
and U6156 (N_6156,N_5119,N_4747);
nor U6157 (N_6157,N_4096,N_5991);
or U6158 (N_6158,N_5145,N_4180);
or U6159 (N_6159,N_5348,N_4165);
nand U6160 (N_6160,N_5667,N_5753);
or U6161 (N_6161,N_5533,N_4099);
or U6162 (N_6162,N_4886,N_4565);
or U6163 (N_6163,N_4452,N_4196);
or U6164 (N_6164,N_4898,N_5754);
and U6165 (N_6165,N_5146,N_4117);
or U6166 (N_6166,N_5561,N_5075);
or U6167 (N_6167,N_5572,N_5611);
and U6168 (N_6168,N_4796,N_4446);
nor U6169 (N_6169,N_4319,N_5982);
or U6170 (N_6170,N_4577,N_4797);
nand U6171 (N_6171,N_5951,N_4080);
and U6172 (N_6172,N_5123,N_4228);
nand U6173 (N_6173,N_5315,N_5843);
nand U6174 (N_6174,N_4760,N_5007);
nand U6175 (N_6175,N_5970,N_5887);
and U6176 (N_6176,N_5351,N_4613);
nor U6177 (N_6177,N_5023,N_4499);
nor U6178 (N_6178,N_4330,N_5598);
and U6179 (N_6179,N_4019,N_4006);
and U6180 (N_6180,N_4748,N_5265);
or U6181 (N_6181,N_4030,N_5786);
or U6182 (N_6182,N_5581,N_5223);
or U6183 (N_6183,N_4938,N_5296);
and U6184 (N_6184,N_4904,N_5219);
nand U6185 (N_6185,N_4739,N_5634);
nand U6186 (N_6186,N_5025,N_4036);
nand U6187 (N_6187,N_4589,N_4356);
or U6188 (N_6188,N_5967,N_4210);
nor U6189 (N_6189,N_4870,N_5499);
or U6190 (N_6190,N_5341,N_5815);
nor U6191 (N_6191,N_4125,N_5868);
and U6192 (N_6192,N_4333,N_5406);
nor U6193 (N_6193,N_5535,N_5163);
and U6194 (N_6194,N_5741,N_5790);
or U6195 (N_6195,N_4581,N_4104);
nor U6196 (N_6196,N_4850,N_5827);
nor U6197 (N_6197,N_5497,N_5839);
nor U6198 (N_6198,N_4882,N_5797);
and U6199 (N_6199,N_5297,N_5420);
nand U6200 (N_6200,N_4867,N_5801);
nand U6201 (N_6201,N_4537,N_4260);
and U6202 (N_6202,N_5308,N_4279);
nand U6203 (N_6203,N_4843,N_5564);
nor U6204 (N_6204,N_5422,N_4934);
nand U6205 (N_6205,N_4348,N_5053);
nand U6206 (N_6206,N_5241,N_4551);
or U6207 (N_6207,N_4538,N_4505);
xor U6208 (N_6208,N_5521,N_4562);
and U6209 (N_6209,N_5910,N_5417);
xor U6210 (N_6210,N_5122,N_4063);
and U6211 (N_6211,N_5386,N_4849);
nand U6212 (N_6212,N_5413,N_4391);
and U6213 (N_6213,N_5865,N_4219);
xnor U6214 (N_6214,N_4231,N_4051);
and U6215 (N_6215,N_4247,N_4536);
nand U6216 (N_6216,N_5999,N_5992);
and U6217 (N_6217,N_5002,N_5391);
nand U6218 (N_6218,N_4550,N_4984);
or U6219 (N_6219,N_5726,N_4558);
nor U6220 (N_6220,N_4278,N_5105);
and U6221 (N_6221,N_4525,N_5942);
or U6222 (N_6222,N_4479,N_5927);
nand U6223 (N_6223,N_5283,N_4688);
nand U6224 (N_6224,N_4229,N_5645);
and U6225 (N_6225,N_4508,N_5763);
and U6226 (N_6226,N_4775,N_5862);
or U6227 (N_6227,N_4790,N_5816);
or U6228 (N_6228,N_5803,N_5337);
nand U6229 (N_6229,N_5585,N_5730);
nand U6230 (N_6230,N_4039,N_5175);
or U6231 (N_6231,N_4181,N_4658);
nor U6232 (N_6232,N_4594,N_4257);
and U6233 (N_6233,N_4056,N_5912);
or U6234 (N_6234,N_5016,N_4779);
nor U6235 (N_6235,N_4546,N_5770);
xor U6236 (N_6236,N_4582,N_5990);
nor U6237 (N_6237,N_4910,N_5863);
xor U6238 (N_6238,N_4440,N_4963);
or U6239 (N_6239,N_5492,N_4507);
or U6240 (N_6240,N_4239,N_4408);
and U6241 (N_6241,N_4222,N_5455);
nand U6242 (N_6242,N_4751,N_5902);
nand U6243 (N_6243,N_5270,N_5683);
nor U6244 (N_6244,N_5295,N_5655);
or U6245 (N_6245,N_4712,N_4095);
and U6246 (N_6246,N_4029,N_5660);
and U6247 (N_6247,N_5293,N_4914);
and U6248 (N_6248,N_4884,N_5450);
nor U6249 (N_6249,N_5448,N_4110);
nand U6250 (N_6250,N_5988,N_5568);
nand U6251 (N_6251,N_5305,N_4424);
or U6252 (N_6252,N_5514,N_4346);
and U6253 (N_6253,N_5717,N_4669);
and U6254 (N_6254,N_5680,N_5956);
or U6255 (N_6255,N_4411,N_4998);
or U6256 (N_6256,N_4897,N_4113);
and U6257 (N_6257,N_5233,N_4160);
and U6258 (N_6258,N_4272,N_5738);
nand U6259 (N_6259,N_5751,N_5966);
nand U6260 (N_6260,N_5673,N_5284);
nand U6261 (N_6261,N_5949,N_4385);
and U6262 (N_6262,N_4803,N_5059);
nand U6263 (N_6263,N_5054,N_4467);
nor U6264 (N_6264,N_4847,N_5744);
nor U6265 (N_6265,N_5477,N_5179);
or U6266 (N_6266,N_5926,N_4549);
nor U6267 (N_6267,N_5733,N_4944);
nor U6268 (N_6268,N_5226,N_5845);
nand U6269 (N_6269,N_5976,N_5482);
and U6270 (N_6270,N_4568,N_4103);
and U6271 (N_6271,N_5050,N_4083);
or U6272 (N_6272,N_4266,N_5411);
nor U6273 (N_6273,N_4457,N_4830);
nand U6274 (N_6274,N_5405,N_4519);
or U6275 (N_6275,N_5039,N_5275);
or U6276 (N_6276,N_4488,N_5946);
nand U6277 (N_6277,N_5734,N_4235);
nand U6278 (N_6278,N_4367,N_5427);
nand U6279 (N_6279,N_4050,N_4543);
nand U6280 (N_6280,N_5174,N_4592);
nor U6281 (N_6281,N_4259,N_5962);
and U6282 (N_6282,N_4734,N_5429);
nand U6283 (N_6283,N_4640,N_4971);
nand U6284 (N_6284,N_5819,N_4988);
or U6285 (N_6285,N_4665,N_4254);
or U6286 (N_6286,N_4297,N_5935);
or U6287 (N_6287,N_4539,N_4526);
nor U6288 (N_6288,N_5508,N_4130);
and U6289 (N_6289,N_5506,N_5661);
and U6290 (N_6290,N_4267,N_4958);
nand U6291 (N_6291,N_5262,N_5516);
nor U6292 (N_6292,N_5339,N_4715);
and U6293 (N_6293,N_4555,N_4768);
and U6294 (N_6294,N_5924,N_5727);
nor U6295 (N_6295,N_5724,N_5189);
and U6296 (N_6296,N_5257,N_5036);
and U6297 (N_6297,N_5390,N_5836);
nand U6298 (N_6298,N_4987,N_5780);
nor U6299 (N_6299,N_5913,N_4572);
and U6300 (N_6300,N_5186,N_4624);
nand U6301 (N_6301,N_4376,N_4469);
and U6302 (N_6302,N_5928,N_5998);
nor U6303 (N_6303,N_4848,N_4808);
nor U6304 (N_6304,N_5138,N_5291);
nand U6305 (N_6305,N_4876,N_5237);
nand U6306 (N_6306,N_5892,N_5032);
or U6307 (N_6307,N_4660,N_5987);
or U6308 (N_6308,N_5250,N_4805);
or U6309 (N_6309,N_5033,N_5908);
and U6310 (N_6310,N_5620,N_5158);
and U6311 (N_6311,N_5044,N_4500);
nand U6312 (N_6312,N_5006,N_5452);
nand U6313 (N_6313,N_4945,N_5682);
or U6314 (N_6314,N_4195,N_4182);
xor U6315 (N_6315,N_5818,N_4852);
nor U6316 (N_6316,N_4406,N_5626);
or U6317 (N_6317,N_5151,N_5005);
and U6318 (N_6318,N_5214,N_4486);
and U6319 (N_6319,N_4547,N_4492);
or U6320 (N_6320,N_4617,N_4483);
and U6321 (N_6321,N_4835,N_4147);
nand U6322 (N_6322,N_4609,N_4673);
or U6323 (N_6323,N_4088,N_5771);
nor U6324 (N_6324,N_5721,N_5896);
or U6325 (N_6325,N_4595,N_5467);
nor U6326 (N_6326,N_5360,N_5584);
and U6327 (N_6327,N_5599,N_5332);
and U6328 (N_6328,N_5309,N_5752);
or U6329 (N_6329,N_4212,N_5212);
nand U6330 (N_6330,N_5382,N_4037);
nand U6331 (N_6331,N_5331,N_4332);
nand U6332 (N_6332,N_5258,N_5355);
and U6333 (N_6333,N_5740,N_5997);
and U6334 (N_6334,N_4205,N_4846);
nor U6335 (N_6335,N_5397,N_5433);
and U6336 (N_6336,N_4470,N_5873);
or U6337 (N_6337,N_4980,N_4596);
nand U6338 (N_6338,N_5077,N_5616);
nand U6339 (N_6339,N_5124,N_4170);
nand U6340 (N_6340,N_5995,N_5921);
and U6341 (N_6341,N_4650,N_5793);
and U6342 (N_6342,N_4889,N_4708);
and U6343 (N_6343,N_4593,N_5367);
nor U6344 (N_6344,N_4389,N_5648);
nor U6345 (N_6345,N_5289,N_4501);
and U6346 (N_6346,N_5183,N_5869);
and U6347 (N_6347,N_5209,N_5761);
nor U6348 (N_6348,N_4220,N_5945);
nor U6349 (N_6349,N_5166,N_5480);
nand U6350 (N_6350,N_5669,N_5500);
and U6351 (N_6351,N_4855,N_5256);
xor U6352 (N_6352,N_4078,N_4927);
or U6353 (N_6353,N_4211,N_4466);
xor U6354 (N_6354,N_5416,N_5253);
nor U6355 (N_6355,N_4695,N_4605);
nand U6356 (N_6356,N_5353,N_4461);
nand U6357 (N_6357,N_5856,N_4793);
nor U6358 (N_6358,N_5658,N_5760);
and U6359 (N_6359,N_5623,N_4528);
nor U6360 (N_6360,N_5890,N_4781);
nand U6361 (N_6361,N_5603,N_4303);
or U6362 (N_6362,N_4474,N_4623);
nand U6363 (N_6363,N_4430,N_4292);
or U6364 (N_6364,N_4370,N_5692);
nor U6365 (N_6365,N_4496,N_5832);
and U6366 (N_6366,N_4075,N_5925);
xnor U6367 (N_6367,N_4354,N_5532);
nand U6368 (N_6368,N_4262,N_4880);
xor U6369 (N_6369,N_5745,N_5379);
or U6370 (N_6370,N_4437,N_5294);
or U6371 (N_6371,N_5720,N_5918);
nor U6372 (N_6372,N_5034,N_4010);
nor U6373 (N_6373,N_4060,N_5483);
or U6374 (N_6374,N_4527,N_4116);
nand U6375 (N_6375,N_5657,N_4215);
nand U6376 (N_6376,N_5624,N_4402);
or U6377 (N_6377,N_5981,N_5546);
nor U6378 (N_6378,N_4670,N_5762);
nand U6379 (N_6379,N_5277,N_4809);
and U6380 (N_6380,N_4872,N_4698);
nand U6381 (N_6381,N_4504,N_5469);
or U6382 (N_6382,N_4514,N_4337);
nor U6383 (N_6383,N_4680,N_4815);
nor U6384 (N_6384,N_4729,N_5852);
nand U6385 (N_6385,N_5631,N_5133);
nand U6386 (N_6386,N_5193,N_5343);
nor U6387 (N_6387,N_4769,N_5232);
xnor U6388 (N_6388,N_5361,N_5043);
nor U6389 (N_6389,N_5311,N_4903);
and U6390 (N_6390,N_4304,N_5605);
nor U6391 (N_6391,N_4783,N_5989);
nor U6392 (N_6392,N_4190,N_5540);
and U6393 (N_6393,N_5526,N_5224);
or U6394 (N_6394,N_5798,N_4342);
and U6395 (N_6395,N_5659,N_5398);
or U6396 (N_6396,N_4143,N_4193);
nor U6397 (N_6397,N_5447,N_5063);
nand U6398 (N_6398,N_4232,N_4684);
nand U6399 (N_6399,N_4907,N_4895);
nand U6400 (N_6400,N_5026,N_5808);
nand U6401 (N_6401,N_4571,N_4863);
or U6402 (N_6402,N_4295,N_4869);
or U6403 (N_6403,N_5102,N_5424);
or U6404 (N_6404,N_5306,N_4834);
xnor U6405 (N_6405,N_5381,N_4651);
nor U6406 (N_6406,N_5236,N_5396);
and U6407 (N_6407,N_5809,N_5074);
nand U6408 (N_6408,N_5855,N_4842);
and U6409 (N_6409,N_4749,N_4048);
and U6410 (N_6410,N_4393,N_4053);
or U6411 (N_6411,N_4314,N_5894);
and U6412 (N_6412,N_5268,N_4347);
nor U6413 (N_6413,N_4719,N_4881);
nand U6414 (N_6414,N_4587,N_5983);
nand U6415 (N_6415,N_5523,N_4401);
nand U6416 (N_6416,N_5380,N_5218);
and U6417 (N_6417,N_5449,N_4383);
and U6418 (N_6418,N_5319,N_5795);
and U6419 (N_6419,N_4822,N_5177);
nor U6420 (N_6420,N_4862,N_5375);
or U6421 (N_6421,N_4240,N_5642);
or U6422 (N_6422,N_5874,N_5707);
and U6423 (N_6423,N_5985,N_4503);
nor U6424 (N_6424,N_4961,N_5008);
and U6425 (N_6425,N_5020,N_4860);
nand U6426 (N_6426,N_5371,N_5440);
or U6427 (N_6427,N_4327,N_5161);
or U6428 (N_6428,N_4114,N_5825);
and U6429 (N_6429,N_4091,N_4710);
or U6430 (N_6430,N_5216,N_4696);
and U6431 (N_6431,N_4156,N_5000);
nor U6432 (N_6432,N_5094,N_4662);
or U6433 (N_6433,N_4746,N_5461);
nor U6434 (N_6434,N_5168,N_4618);
and U6435 (N_6435,N_5853,N_4288);
nand U6436 (N_6436,N_4687,N_5357);
xor U6437 (N_6437,N_5399,N_4704);
or U6438 (N_6438,N_4396,N_4957);
nor U6439 (N_6439,N_4064,N_4326);
or U6440 (N_6440,N_5732,N_4909);
nand U6441 (N_6441,N_5677,N_4755);
nor U6442 (N_6442,N_5678,N_4329);
or U6443 (N_6443,N_5022,N_4552);
and U6444 (N_6444,N_4177,N_5049);
and U6445 (N_6445,N_5335,N_4933);
nor U6446 (N_6446,N_5899,N_4243);
and U6447 (N_6447,N_4919,N_4345);
or U6448 (N_6448,N_5933,N_5069);
xor U6449 (N_6449,N_4887,N_4172);
nand U6450 (N_6450,N_4681,N_4159);
nor U6451 (N_6451,N_4493,N_5590);
and U6452 (N_6452,N_4225,N_5345);
or U6453 (N_6453,N_5943,N_5093);
nor U6454 (N_6454,N_4097,N_4630);
nor U6455 (N_6455,N_4542,N_5114);
or U6456 (N_6456,N_4472,N_4634);
nand U6457 (N_6457,N_4576,N_4227);
nand U6458 (N_6458,N_5604,N_4054);
nor U6459 (N_6459,N_4692,N_5208);
and U6460 (N_6460,N_5507,N_4915);
nand U6461 (N_6461,N_5686,N_5290);
xor U6462 (N_6462,N_4981,N_4663);
and U6463 (N_6463,N_4460,N_4780);
nor U6464 (N_6464,N_4677,N_5403);
nand U6465 (N_6465,N_5081,N_5571);
and U6466 (N_6466,N_5097,N_4885);
or U6467 (N_6467,N_4028,N_4026);
nand U6468 (N_6468,N_4646,N_4811);
nand U6469 (N_6469,N_5327,N_4497);
and U6470 (N_6470,N_4727,N_5794);
nor U6471 (N_6471,N_4102,N_5635);
nor U6472 (N_6472,N_4711,N_4584);
nor U6473 (N_6473,N_5650,N_5906);
nand U6474 (N_6474,N_4828,N_4204);
and U6475 (N_6475,N_5679,N_5066);
and U6476 (N_6476,N_4632,N_4865);
nand U6477 (N_6477,N_4816,N_5594);
nand U6478 (N_6478,N_4422,N_5675);
nor U6479 (N_6479,N_4604,N_4564);
and U6480 (N_6480,N_5264,N_4061);
nor U6481 (N_6481,N_4798,N_4206);
nand U6482 (N_6482,N_4638,N_4155);
nor U6483 (N_6483,N_5463,N_4163);
nand U6484 (N_6484,N_4778,N_5746);
nand U6485 (N_6485,N_4818,N_5338);
and U6486 (N_6486,N_5860,N_4129);
nand U6487 (N_6487,N_5126,N_5881);
nand U6488 (N_6488,N_4982,N_5750);
nor U6489 (N_6489,N_5120,N_4305);
or U6490 (N_6490,N_4548,N_4157);
nor U6491 (N_6491,N_4923,N_5113);
nand U6492 (N_6492,N_4433,N_5222);
nand U6493 (N_6493,N_5848,N_5324);
xor U6494 (N_6494,N_5937,N_5065);
or U6495 (N_6495,N_5950,N_4245);
and U6496 (N_6496,N_5374,N_5110);
and U6497 (N_6497,N_4055,N_4403);
xor U6498 (N_6498,N_4369,N_5435);
or U6499 (N_6499,N_5235,N_5969);
nor U6500 (N_6500,N_4198,N_4451);
and U6501 (N_6501,N_5109,N_4668);
or U6502 (N_6502,N_4964,N_4986);
nor U6503 (N_6503,N_4161,N_4737);
nand U6504 (N_6504,N_5495,N_5804);
nand U6505 (N_6505,N_5476,N_4913);
and U6506 (N_6506,N_4033,N_5973);
nor U6507 (N_6507,N_4567,N_4454);
nand U6508 (N_6508,N_5021,N_4268);
nor U6509 (N_6509,N_5676,N_4014);
nand U6510 (N_6510,N_5274,N_5445);
nor U6511 (N_6511,N_5116,N_4335);
xor U6512 (N_6512,N_4301,N_5115);
xnor U6513 (N_6513,N_5715,N_4534);
or U6514 (N_6514,N_4032,N_5559);
nor U6515 (N_6515,N_4223,N_4464);
and U6516 (N_6516,N_5392,N_5478);
nor U6517 (N_6517,N_4602,N_5889);
xor U6518 (N_6518,N_5814,N_5106);
or U6519 (N_6519,N_4445,N_5828);
nor U6520 (N_6520,N_4679,N_4917);
or U6521 (N_6521,N_5688,N_4832);
or U6522 (N_6522,N_5759,N_4883);
xor U6523 (N_6523,N_5773,N_4703);
nor U6524 (N_6524,N_5723,N_4607);
nand U6525 (N_6525,N_5938,N_5958);
or U6526 (N_6526,N_4306,N_5895);
xnor U6527 (N_6527,N_5152,N_4066);
nor U6528 (N_6528,N_4141,N_5971);
and U6529 (N_6529,N_4480,N_5563);
nand U6530 (N_6530,N_5073,N_5273);
and U6531 (N_6531,N_5234,N_4952);
and U6532 (N_6532,N_5302,N_5330);
or U6533 (N_6533,N_4926,N_5666);
or U6534 (N_6534,N_4627,N_4120);
or U6535 (N_6535,N_4740,N_4512);
nand U6536 (N_6536,N_4892,N_5911);
and U6537 (N_6537,N_5531,N_4473);
or U6538 (N_6538,N_5799,N_4559);
nand U6539 (N_6539,N_4786,N_4052);
nor U6540 (N_6540,N_5489,N_5041);
nand U6541 (N_6541,N_4676,N_4761);
nor U6542 (N_6542,N_5292,N_5702);
or U6543 (N_6543,N_5127,N_4743);
nor U6544 (N_6544,N_5045,N_5550);
or U6545 (N_6545,N_4731,N_4750);
and U6546 (N_6546,N_5766,N_4046);
nor U6547 (N_6547,N_4965,N_5304);
nand U6548 (N_6548,N_4286,N_5555);
nor U6549 (N_6549,N_5468,N_5586);
or U6550 (N_6550,N_4639,N_4845);
or U6551 (N_6551,N_4771,N_4355);
nor U6552 (N_6552,N_5530,N_4968);
or U6553 (N_6553,N_4044,N_5090);
or U6554 (N_6554,N_4233,N_5431);
and U6555 (N_6555,N_4901,N_4645);
nand U6556 (N_6556,N_5084,N_5394);
nand U6557 (N_6557,N_4833,N_4837);
and U6558 (N_6558,N_4049,N_5613);
nor U6559 (N_6559,N_4381,N_4414);
nand U6560 (N_6560,N_5851,N_4224);
or U6561 (N_6561,N_4588,N_5718);
nand U6562 (N_6562,N_5965,N_4173);
or U6563 (N_6563,N_5276,N_5207);
nor U6564 (N_6564,N_5164,N_5269);
and U6565 (N_6565,N_4132,N_4249);
or U6566 (N_6566,N_4840,N_4894);
and U6567 (N_6567,N_5662,N_4434);
nand U6568 (N_6568,N_5652,N_5434);
nor U6569 (N_6569,N_4929,N_4657);
nand U6570 (N_6570,N_4443,N_4311);
nand U6571 (N_6571,N_4610,N_4021);
and U6572 (N_6572,N_4397,N_5215);
nand U6573 (N_6573,N_4967,N_4270);
or U6574 (N_6574,N_4122,N_4040);
or U6575 (N_6575,N_4238,N_5464);
nor U6576 (N_6576,N_5960,N_4018);
nand U6577 (N_6577,N_4167,N_5062);
or U6578 (N_6578,N_4515,N_5260);
nand U6579 (N_6579,N_5663,N_5112);
nor U6580 (N_6580,N_5035,N_4090);
nand U6581 (N_6581,N_5060,N_4948);
or U6582 (N_6582,N_5637,N_5904);
and U6583 (N_6583,N_5570,N_4377);
and U6584 (N_6584,N_5542,N_4360);
nand U6585 (N_6585,N_5061,N_5857);
nand U6586 (N_6586,N_4388,N_5131);
nand U6587 (N_6587,N_4922,N_4924);
xor U6588 (N_6588,N_5111,N_4435);
and U6589 (N_6589,N_5879,N_4659);
nand U6590 (N_6590,N_5897,N_4518);
or U6591 (N_6591,N_5737,N_4742);
and U6592 (N_6592,N_5165,N_4334);
and U6593 (N_6593,N_4017,N_4586);
and U6594 (N_6594,N_4144,N_4598);
nand U6595 (N_6595,N_5693,N_5085);
and U6596 (N_6596,N_4995,N_5457);
nand U6597 (N_6597,N_5202,N_5196);
nor U6598 (N_6598,N_4918,N_4825);
nor U6599 (N_6599,N_4960,N_4707);
or U6600 (N_6600,N_4005,N_5975);
or U6601 (N_6601,N_5419,N_5807);
nand U6602 (N_6602,N_4368,N_4899);
or U6603 (N_6603,N_4859,N_5366);
and U6604 (N_6604,N_4082,N_4950);
nand U6605 (N_6605,N_4643,N_4619);
or U6606 (N_6606,N_5647,N_5470);
or U6607 (N_6607,N_5764,N_4701);
and U6608 (N_6608,N_4317,N_5245);
or U6609 (N_6609,N_4202,N_4185);
or U6610 (N_6610,N_4248,N_5015);
or U6611 (N_6611,N_5156,N_5699);
and U6612 (N_6612,N_5004,N_5047);
or U6613 (N_6613,N_4625,N_4615);
nand U6614 (N_6614,N_5589,N_5228);
nand U6615 (N_6615,N_4149,N_4873);
or U6616 (N_6616,N_5580,N_4718);
and U6617 (N_6617,N_4826,N_5858);
nand U6618 (N_6618,N_5388,N_4265);
and U6619 (N_6619,N_5984,N_4153);
nor U6620 (N_6620,N_5545,N_4714);
and U6621 (N_6621,N_4343,N_5040);
and U6622 (N_6622,N_4057,N_5651);
nand U6623 (N_6623,N_4820,N_5206);
nor U6624 (N_6624,N_5596,N_4404);
or U6625 (N_6625,N_5588,N_5329);
or U6626 (N_6626,N_4621,N_5252);
nor U6627 (N_6627,N_4799,N_4575);
and U6628 (N_6628,N_4184,N_4674);
nand U6629 (N_6629,N_5914,N_4978);
nand U6630 (N_6630,N_5130,N_4972);
and U6631 (N_6631,N_5255,N_4656);
nand U6632 (N_6632,N_5671,N_4208);
nor U6633 (N_6633,N_4287,N_4118);
and U6634 (N_6634,N_5389,N_5841);
nand U6635 (N_6635,N_5512,N_5363);
nand U6636 (N_6636,N_5395,N_4759);
nand U6637 (N_6637,N_5082,N_4994);
and U6638 (N_6638,N_5087,N_5552);
and U6639 (N_6639,N_5710,N_5267);
or U6640 (N_6640,N_5068,N_5577);
nor U6641 (N_6641,N_5031,N_5701);
xnor U6642 (N_6642,N_4947,N_4313);
nor U6643 (N_6643,N_5432,N_5028);
xor U6644 (N_6644,N_4213,N_5200);
nor U6645 (N_6645,N_5354,N_4599);
nor U6646 (N_6646,N_4336,N_5154);
and U6647 (N_6647,N_4787,N_5187);
and U6648 (N_6648,N_5412,N_4448);
and U6649 (N_6649,N_5583,N_4509);
nor U6650 (N_6650,N_5952,N_4468);
xor U6651 (N_6651,N_4041,N_4236);
nor U6652 (N_6652,N_5453,N_5840);
and U6653 (N_6653,N_5439,N_5749);
nand U6654 (N_6654,N_5861,N_5010);
and U6655 (N_6655,N_5640,N_4541);
nor U6656 (N_6656,N_5711,N_5847);
and U6657 (N_6657,N_4912,N_5205);
nand U6658 (N_6658,N_4893,N_4359);
or U6659 (N_6659,N_4631,N_4256);
nand U6660 (N_6660,N_5426,N_4124);
and U6661 (N_6661,N_4285,N_5811);
nand U6662 (N_6662,N_5286,N_5557);
and U6663 (N_6663,N_5172,N_5248);
nand U6664 (N_6664,N_5529,N_4517);
nor U6665 (N_6665,N_4073,N_4186);
nand U6666 (N_6666,N_5544,N_5697);
and U6667 (N_6667,N_4209,N_4682);
nor U6668 (N_6668,N_5118,N_5519);
nand U6669 (N_6669,N_4813,N_4425);
and U6670 (N_6670,N_5046,N_5947);
and U6671 (N_6671,N_4142,N_4494);
nand U6672 (N_6672,N_5103,N_5872);
nor U6673 (N_6673,N_5242,N_4169);
nor U6674 (N_6674,N_5190,N_5575);
nand U6675 (N_6675,N_4557,N_4413);
and U6676 (N_6676,N_5788,N_4463);
nand U6677 (N_6677,N_4072,N_4127);
nor U6678 (N_6678,N_5592,N_4216);
and U6679 (N_6679,N_5684,N_4996);
nand U6680 (N_6680,N_5802,N_5408);
and U6681 (N_6681,N_5574,N_5247);
nand U6682 (N_6682,N_5473,N_4477);
nor U6683 (N_6683,N_5672,N_4062);
and U6684 (N_6684,N_4744,N_5994);
or U6685 (N_6685,N_5155,N_4611);
and U6686 (N_6686,N_4770,N_5769);
nand U6687 (N_6687,N_5080,N_4139);
or U6688 (N_6688,N_5549,N_4735);
nor U6689 (N_6689,N_4275,N_5916);
and U6690 (N_6690,N_4709,N_5052);
or U6691 (N_6691,N_5013,N_4752);
nand U6692 (N_6692,N_5901,N_4671);
nand U6693 (N_6693,N_4400,N_4320);
nand U6694 (N_6694,N_5129,N_5978);
and U6695 (N_6695,N_5917,N_4531);
nand U6696 (N_6696,N_4841,N_5644);
nor U6697 (N_6697,N_5757,N_5472);
or U6698 (N_6698,N_4016,N_4379);
xor U6699 (N_6699,N_5278,N_4294);
nand U6700 (N_6700,N_5822,N_5377);
xor U6701 (N_6701,N_4603,N_5690);
nor U6702 (N_6702,N_4878,N_4276);
or U6703 (N_6703,N_5018,N_5486);
and U6704 (N_6704,N_5515,N_4908);
xor U6705 (N_6705,N_5930,N_4844);
nand U6706 (N_6706,N_4171,N_4447);
and U6707 (N_6707,N_5213,N_5344);
nand U6708 (N_6708,N_4008,N_4974);
nor U6709 (N_6709,N_4069,N_5384);
nor U6710 (N_6710,N_4854,N_5934);
and U6711 (N_6711,N_5368,N_5079);
or U6712 (N_6712,N_5051,N_5091);
nor U6713 (N_6713,N_4281,N_4554);
nand U6714 (N_6714,N_5490,N_4364);
or U6715 (N_6715,N_5167,N_4758);
or U6716 (N_6716,N_5474,N_4678);
and U6717 (N_6717,N_5821,N_4513);
nand U6718 (N_6718,N_5600,N_5322);
nand U6719 (N_6719,N_4824,N_4800);
and U6720 (N_6720,N_4626,N_4321);
or U6721 (N_6721,N_4817,N_4084);
or U6722 (N_6722,N_4375,N_5373);
nand U6723 (N_6723,N_5092,N_5909);
and U6724 (N_6724,N_5443,N_4119);
nor U6725 (N_6725,N_5940,N_5488);
and U6726 (N_6726,N_4810,N_4935);
or U6727 (N_6727,N_4094,N_4789);
nor U6728 (N_6728,N_5221,N_4200);
or U6729 (N_6729,N_4444,N_5347);
nand U6730 (N_6730,N_4642,N_5880);
nor U6731 (N_6731,N_4449,N_4535);
or U6732 (N_6732,N_5014,N_5220);
or U6733 (N_6733,N_5326,N_4516);
nor U6734 (N_6734,N_4175,N_4284);
nor U6735 (N_6735,N_4812,N_4436);
or U6736 (N_6736,N_5496,N_5083);
and U6737 (N_6737,N_5665,N_5418);
nor U6738 (N_6738,N_5628,N_5722);
or U6739 (N_6739,N_4776,N_4123);
nand U6740 (N_6740,N_4242,N_4991);
nor U6741 (N_6741,N_4533,N_4906);
nor U6742 (N_6742,N_5558,N_4420);
or U6743 (N_6743,N_5055,N_5636);
nand U6744 (N_6744,N_4720,N_5184);
or U6745 (N_6745,N_4601,N_5517);
or U6746 (N_6746,N_5893,N_4357);
and U6747 (N_6747,N_4489,N_4888);
or U6748 (N_6748,N_4969,N_5334);
nor U6749 (N_6749,N_5001,N_5919);
nor U6750 (N_6750,N_5639,N_5758);
or U6751 (N_6751,N_5176,N_4324);
and U6752 (N_6752,N_4218,N_5227);
and U6753 (N_6753,N_5963,N_5980);
nor U6754 (N_6754,N_5882,N_5307);
or U6755 (N_6755,N_4937,N_5350);
and U6756 (N_6756,N_4418,N_4482);
or U6757 (N_6757,N_4877,N_4351);
nand U6758 (N_6758,N_4409,N_5823);
or U6759 (N_6759,N_5444,N_4866);
xnor U6760 (N_6760,N_5838,N_5030);
nand U6761 (N_6761,N_5719,N_4620);
nand U6762 (N_6762,N_4352,N_5003);
and U6763 (N_6763,N_5829,N_4829);
or U6764 (N_6764,N_4419,N_5955);
and U6765 (N_6765,N_4721,N_4801);
nand U6766 (N_6766,N_5185,N_4203);
nor U6767 (N_6767,N_4890,N_4956);
or U6768 (N_6768,N_4187,N_4023);
nor U6769 (N_6769,N_5668,N_4007);
or U6770 (N_6770,N_5509,N_5747);
nor U6771 (N_6771,N_5314,N_5817);
nor U6772 (N_6772,N_5835,N_4074);
or U6773 (N_6773,N_5423,N_5743);
nand U6774 (N_6774,N_5421,N_5148);
nand U6775 (N_6775,N_4648,N_5664);
and U6776 (N_6776,N_5098,N_4133);
or U6777 (N_6777,N_5820,N_4201);
and U6778 (N_6778,N_5687,N_5135);
and U6779 (N_6779,N_5194,N_5830);
nand U6780 (N_6780,N_5280,N_4322);
or U6781 (N_6781,N_5078,N_5602);
or U6782 (N_6782,N_4821,N_5783);
or U6783 (N_6783,N_4713,N_4521);
or U6784 (N_6784,N_4458,N_4655);
nor U6785 (N_6785,N_4579,N_5805);
nand U6786 (N_6786,N_4856,N_5012);
and U6787 (N_6787,N_4093,N_4131);
nor U6788 (N_6788,N_5844,N_4226);
nand U6789 (N_6789,N_5225,N_5767);
nand U6790 (N_6790,N_5867,N_5957);
nand U6791 (N_6791,N_5905,N_4520);
nand U6792 (N_6792,N_4975,N_4012);
nor U6793 (N_6793,N_5451,N_5731);
nand U6794 (N_6794,N_4111,N_5736);
and U6795 (N_6795,N_4853,N_5132);
or U6796 (N_6796,N_4951,N_4481);
nor U6797 (N_6797,N_5735,N_5777);
nand U6798 (N_6798,N_5787,N_4135);
nand U6799 (N_6799,N_5204,N_4067);
and U6800 (N_6800,N_5136,N_4410);
and U6801 (N_6801,N_4085,N_4814);
and U6802 (N_6802,N_4341,N_4148);
or U6803 (N_6803,N_5378,N_4106);
or U6804 (N_6804,N_5772,N_5824);
nor U6805 (N_6805,N_4128,N_5459);
or U6806 (N_6806,N_5621,N_4134);
and U6807 (N_6807,N_4983,N_4471);
and U6808 (N_6808,N_4307,N_5597);
and U6809 (N_6809,N_4459,N_4077);
and U6810 (N_6810,N_5936,N_4962);
nor U6811 (N_6811,N_4456,N_5674);
and U6812 (N_6812,N_4732,N_5058);
nor U6813 (N_6813,N_4384,N_5883);
xnor U6814 (N_6814,N_5088,N_5140);
and U6815 (N_6815,N_4255,N_5866);
and U6816 (N_6816,N_4689,N_4861);
nand U6817 (N_6817,N_5104,N_5565);
nor U6818 (N_6818,N_4900,N_5556);
or U6819 (N_6819,N_4079,N_5099);
nand U6820 (N_6820,N_5695,N_5460);
nand U6821 (N_6821,N_5974,N_4387);
and U6822 (N_6822,N_5279,N_5510);
or U6823 (N_6823,N_4230,N_5864);
and U6824 (N_6824,N_4902,N_5024);
nor U6825 (N_6825,N_5850,N_5261);
or U6826 (N_6826,N_5134,N_5323);
nor U6827 (N_6827,N_4373,N_5430);
nand U6828 (N_6828,N_4694,N_4916);
nor U6829 (N_6829,N_5670,N_5870);
and U6830 (N_6830,N_5539,N_4020);
nand U6831 (N_6831,N_5494,N_5150);
and U6832 (N_6832,N_4524,N_5629);
nand U6833 (N_6833,N_5071,N_4857);
nand U6834 (N_6834,N_4868,N_5318);
nand U6835 (N_6835,N_4365,N_5800);
or U6836 (N_6836,N_5961,N_4453);
nand U6837 (N_6837,N_4363,N_5171);
or U6838 (N_6838,N_5211,N_5513);
and U6839 (N_6839,N_4591,N_4282);
or U6840 (N_6840,N_4392,N_5876);
and U6841 (N_6841,N_5349,N_4785);
nor U6842 (N_6842,N_5201,N_5402);
nand U6843 (N_6843,N_5029,N_5573);
nor U6844 (N_6844,N_4109,N_4300);
and U6845 (N_6845,N_4570,N_5199);
or U6846 (N_6846,N_4126,N_4350);
nor U6847 (N_6847,N_4940,N_5153);
xnor U6848 (N_6848,N_5299,N_4269);
nand U6849 (N_6849,N_5502,N_5310);
and U6850 (N_6850,N_4484,N_5789);
nand U6851 (N_6851,N_4690,N_5244);
nor U6852 (N_6852,N_5410,N_5372);
nor U6853 (N_6853,N_4237,N_5246);
or U6854 (N_6854,N_4905,N_4004);
nor U6855 (N_6855,N_4722,N_5833);
or U6856 (N_6856,N_5527,N_5560);
nor U6857 (N_6857,N_5238,N_5285);
and U6858 (N_6858,N_5181,N_5197);
nor U6859 (N_6859,N_5871,N_5011);
and U6860 (N_6860,N_5230,N_5462);
nor U6861 (N_6861,N_4246,N_5595);
and U6862 (N_6862,N_4310,N_4183);
and U6863 (N_6863,N_4772,N_5923);
and U6864 (N_6864,N_5792,N_4158);
and U6865 (N_6865,N_4891,N_4289);
or U6866 (N_6866,N_5162,N_4087);
nor U6867 (N_6867,N_4031,N_4545);
nand U6868 (N_6868,N_5785,N_4065);
nor U6869 (N_6869,N_4108,N_4941);
nor U6870 (N_6870,N_5959,N_5456);
nor U6871 (N_6871,N_4635,N_4192);
and U6872 (N_6872,N_5485,N_4725);
or U6873 (N_6873,N_5301,N_4349);
nand U6874 (N_6874,N_5681,N_5617);
nand U6875 (N_6875,N_4328,N_5782);
nor U6876 (N_6876,N_4736,N_4271);
or U6877 (N_6877,N_5147,N_5837);
or U6878 (N_6878,N_4024,N_4431);
or U6879 (N_6879,N_4107,N_5685);
nor U6880 (N_6880,N_4485,N_5210);
or U6881 (N_6881,N_5229,N_4398);
nand U6882 (N_6882,N_5400,N_5886);
nand U6883 (N_6883,N_5619,N_4730);
nand U6884 (N_6884,N_4942,N_4174);
nor U6885 (N_6885,N_4686,N_5948);
or U6886 (N_6886,N_4702,N_4985);
nor U6887 (N_6887,N_5471,N_4716);
or U6888 (N_6888,N_4851,N_5756);
nor U6889 (N_6889,N_5325,N_5393);
and U6890 (N_6890,N_5139,N_4807);
nand U6891 (N_6891,N_5356,N_5748);
nor U6892 (N_6892,N_5487,N_4495);
nor U6893 (N_6893,N_5095,N_4428);
xor U6894 (N_6894,N_5076,N_4112);
nand U6895 (N_6895,N_5100,N_4700);
nand U6896 (N_6896,N_5465,N_4178);
or U6897 (N_6897,N_4081,N_4529);
nand U6898 (N_6898,N_5437,N_4498);
nand U6899 (N_6899,N_5072,N_5143);
and U6900 (N_6900,N_4000,N_5705);
or U6901 (N_6901,N_5654,N_4380);
nand U6902 (N_6902,N_5169,N_5300);
or U6903 (N_6903,N_4027,N_5915);
and U6904 (N_6904,N_4920,N_5859);
or U6905 (N_6905,N_5567,N_4612);
nand U6906 (N_6906,N_5409,N_4931);
and U6907 (N_6907,N_4939,N_4754);
nand U6908 (N_6908,N_4804,N_4506);
and U6909 (N_6909,N_4706,N_4836);
nand U6910 (N_6910,N_4331,N_5383);
or U6911 (N_6911,N_5810,N_5259);
and U6912 (N_6912,N_4261,N_5320);
nor U6913 (N_6913,N_5387,N_4491);
nor U6914 (N_6914,N_5582,N_4199);
nand U6915 (N_6915,N_5691,N_4086);
nor U6916 (N_6916,N_5454,N_4374);
and U6917 (N_6917,N_5713,N_4723);
or U6918 (N_6918,N_4540,N_4145);
and U6919 (N_6919,N_4763,N_4407);
and U6920 (N_6920,N_5846,N_5251);
nor U6921 (N_6921,N_4839,N_4578);
nand U6922 (N_6922,N_4649,N_4990);
and U6923 (N_6923,N_4003,N_5643);
nor U6924 (N_6924,N_4146,N_5579);
nand U6925 (N_6925,N_4667,N_5826);
or U6926 (N_6926,N_5159,N_5796);
nand U6927 (N_6927,N_5625,N_4487);
nor U6928 (N_6928,N_4652,N_4415);
or U6929 (N_6929,N_5415,N_4308);
nand U6930 (N_6930,N_5993,N_5728);
and U6931 (N_6931,N_5038,N_4622);
nor U6932 (N_6932,N_5954,N_4115);
or U6933 (N_6933,N_5878,N_5342);
and U6934 (N_6934,N_4608,N_5121);
nor U6935 (N_6935,N_5922,N_4250);
or U6936 (N_6936,N_5142,N_5370);
and U6937 (N_6937,N_4590,N_5755);
nor U6938 (N_6938,N_5352,N_4795);
xor U6939 (N_6939,N_4726,N_5775);
nand U6940 (N_6940,N_4362,N_5709);
and U6941 (N_6941,N_4970,N_5086);
and U6942 (N_6942,N_4788,N_5064);
nand U6943 (N_6943,N_4728,N_4683);
nand U6944 (N_6944,N_5903,N_5160);
nor U6945 (N_6945,N_4455,N_5446);
nor U6946 (N_6946,N_5298,N_4194);
nor U6947 (N_6947,N_4399,N_5607);
or U6948 (N_6948,N_4439,N_4299);
and U6949 (N_6949,N_4450,N_4101);
nor U6950 (N_6950,N_4138,N_5401);
or U6951 (N_6951,N_4765,N_4973);
nor U6952 (N_6952,N_5898,N_5333);
and U6953 (N_6953,N_4979,N_4423);
or U6954 (N_6954,N_5641,N_4315);
xor U6955 (N_6955,N_4738,N_5107);
nor U6956 (N_6956,N_4741,N_4338);
or U6957 (N_6957,N_5137,N_4405);
or U6958 (N_6958,N_5316,N_5170);
or U6959 (N_6959,N_5548,N_5438);
nor U6960 (N_6960,N_5614,N_4100);
nor U6961 (N_6961,N_4154,N_4140);
and U6962 (N_6962,N_4666,N_4871);
or U6963 (N_6963,N_5491,N_4502);
or U6964 (N_6964,N_4757,N_4522);
and U6965 (N_6965,N_4386,N_5578);
or U6966 (N_6966,N_4371,N_5907);
nand U6967 (N_6967,N_4462,N_4756);
nand U6968 (N_6968,N_5042,N_4475);
and U6969 (N_6969,N_4636,N_4312);
and U6970 (N_6970,N_5428,N_4661);
and U6971 (N_6971,N_4323,N_5696);
nor U6972 (N_6972,N_4263,N_5217);
nand U6973 (N_6973,N_5977,N_5689);
or U6974 (N_6974,N_5522,N_5195);
nor U6975 (N_6975,N_4432,N_5484);
or U6976 (N_6976,N_4925,N_4465);
and U6977 (N_6977,N_4523,N_5553);
and U6978 (N_6978,N_5466,N_5834);
and U6979 (N_6979,N_4277,N_4253);
xnor U6980 (N_6980,N_5609,N_4764);
and U6981 (N_6981,N_4693,N_4162);
nand U6982 (N_6982,N_4955,N_5425);
nand U6983 (N_6983,N_4152,N_5698);
and U6984 (N_6984,N_4035,N_5524);
or U6985 (N_6985,N_4059,N_4954);
and U6986 (N_6986,N_4838,N_5520);
nor U6987 (N_6987,N_4911,N_5618);
nand U6988 (N_6988,N_5968,N_4977);
or U6989 (N_6989,N_4164,N_4875);
or U6990 (N_6990,N_4339,N_4510);
nor U6991 (N_6991,N_4478,N_4614);
nor U6992 (N_6992,N_4993,N_5700);
or U6993 (N_6993,N_5656,N_4372);
and U6994 (N_6994,N_5192,N_4244);
or U6995 (N_6995,N_5569,N_4637);
nand U6996 (N_6996,N_4258,N_4047);
or U6997 (N_6997,N_5986,N_5806);
nand U6998 (N_6998,N_5633,N_4291);
or U6999 (N_6999,N_4011,N_5376);
and U7000 (N_7000,N_4022,N_5366);
and U7001 (N_7001,N_5784,N_4077);
or U7002 (N_7002,N_5091,N_4926);
nand U7003 (N_7003,N_5627,N_5448);
nand U7004 (N_7004,N_5295,N_5348);
or U7005 (N_7005,N_4146,N_5534);
nor U7006 (N_7006,N_4368,N_4788);
or U7007 (N_7007,N_5538,N_4440);
nand U7008 (N_7008,N_5837,N_5430);
or U7009 (N_7009,N_5932,N_4268);
nand U7010 (N_7010,N_5695,N_4224);
or U7011 (N_7011,N_5773,N_4693);
nor U7012 (N_7012,N_5402,N_4071);
nand U7013 (N_7013,N_4060,N_4669);
or U7014 (N_7014,N_5600,N_5807);
xor U7015 (N_7015,N_5557,N_4798);
nor U7016 (N_7016,N_4839,N_5551);
or U7017 (N_7017,N_4896,N_5441);
or U7018 (N_7018,N_5474,N_5340);
nor U7019 (N_7019,N_4041,N_5473);
and U7020 (N_7020,N_5653,N_5435);
nor U7021 (N_7021,N_5245,N_5468);
and U7022 (N_7022,N_5059,N_4191);
nand U7023 (N_7023,N_5022,N_4633);
nand U7024 (N_7024,N_4809,N_5284);
nand U7025 (N_7025,N_5582,N_4485);
or U7026 (N_7026,N_5708,N_4615);
nor U7027 (N_7027,N_5038,N_5410);
nand U7028 (N_7028,N_5640,N_5674);
nand U7029 (N_7029,N_5276,N_4858);
nand U7030 (N_7030,N_4731,N_5114);
or U7031 (N_7031,N_5495,N_4588);
and U7032 (N_7032,N_4467,N_4197);
and U7033 (N_7033,N_4450,N_4193);
nor U7034 (N_7034,N_4807,N_5697);
nand U7035 (N_7035,N_5054,N_5487);
nand U7036 (N_7036,N_4248,N_5385);
nand U7037 (N_7037,N_5322,N_4802);
and U7038 (N_7038,N_5536,N_4841);
nand U7039 (N_7039,N_5234,N_4427);
and U7040 (N_7040,N_4180,N_5257);
or U7041 (N_7041,N_5823,N_5221);
and U7042 (N_7042,N_4048,N_5657);
and U7043 (N_7043,N_4836,N_5915);
xor U7044 (N_7044,N_5156,N_4316);
and U7045 (N_7045,N_5693,N_4465);
nand U7046 (N_7046,N_4912,N_4826);
and U7047 (N_7047,N_4708,N_4571);
xnor U7048 (N_7048,N_4439,N_4894);
and U7049 (N_7049,N_5813,N_4319);
and U7050 (N_7050,N_5189,N_5318);
nor U7051 (N_7051,N_5754,N_5014);
and U7052 (N_7052,N_4367,N_5722);
nor U7053 (N_7053,N_5049,N_4377);
nand U7054 (N_7054,N_4346,N_5596);
nand U7055 (N_7055,N_5743,N_5719);
nand U7056 (N_7056,N_4600,N_5852);
nand U7057 (N_7057,N_4579,N_5750);
xnor U7058 (N_7058,N_4377,N_5481);
nand U7059 (N_7059,N_4269,N_4722);
and U7060 (N_7060,N_5639,N_5793);
nor U7061 (N_7061,N_4418,N_5359);
and U7062 (N_7062,N_4661,N_5964);
nand U7063 (N_7063,N_5979,N_5706);
nor U7064 (N_7064,N_5667,N_4489);
nor U7065 (N_7065,N_5620,N_4936);
and U7066 (N_7066,N_5745,N_5257);
and U7067 (N_7067,N_4561,N_5104);
and U7068 (N_7068,N_5102,N_4529);
and U7069 (N_7069,N_4280,N_4161);
or U7070 (N_7070,N_4256,N_4276);
or U7071 (N_7071,N_5024,N_5583);
xnor U7072 (N_7072,N_5169,N_4401);
nor U7073 (N_7073,N_4548,N_5551);
or U7074 (N_7074,N_5846,N_5575);
nor U7075 (N_7075,N_4390,N_5385);
or U7076 (N_7076,N_5266,N_4275);
nor U7077 (N_7077,N_4206,N_5819);
nand U7078 (N_7078,N_4205,N_5294);
or U7079 (N_7079,N_5559,N_4990);
nand U7080 (N_7080,N_4118,N_5568);
nand U7081 (N_7081,N_4358,N_5392);
and U7082 (N_7082,N_4477,N_4305);
or U7083 (N_7083,N_4647,N_4931);
xor U7084 (N_7084,N_5785,N_4538);
and U7085 (N_7085,N_5122,N_5739);
nor U7086 (N_7086,N_5277,N_4430);
nor U7087 (N_7087,N_4355,N_5184);
and U7088 (N_7088,N_5910,N_5621);
xor U7089 (N_7089,N_4081,N_4927);
nor U7090 (N_7090,N_4238,N_5198);
and U7091 (N_7091,N_5523,N_5954);
or U7092 (N_7092,N_4716,N_4720);
nor U7093 (N_7093,N_4058,N_5656);
xor U7094 (N_7094,N_4458,N_4790);
and U7095 (N_7095,N_4271,N_5043);
and U7096 (N_7096,N_4378,N_5785);
nor U7097 (N_7097,N_4758,N_4802);
nand U7098 (N_7098,N_4764,N_5087);
or U7099 (N_7099,N_4910,N_5790);
nand U7100 (N_7100,N_5352,N_4813);
xnor U7101 (N_7101,N_4196,N_4797);
or U7102 (N_7102,N_5372,N_5172);
or U7103 (N_7103,N_4299,N_4171);
nor U7104 (N_7104,N_4614,N_5259);
nor U7105 (N_7105,N_4244,N_5061);
nor U7106 (N_7106,N_4271,N_5656);
nor U7107 (N_7107,N_4837,N_5841);
nand U7108 (N_7108,N_4444,N_5483);
and U7109 (N_7109,N_4370,N_4369);
and U7110 (N_7110,N_5177,N_5258);
or U7111 (N_7111,N_5152,N_5082);
nand U7112 (N_7112,N_4453,N_4000);
nor U7113 (N_7113,N_5922,N_5275);
nand U7114 (N_7114,N_4855,N_5878);
nor U7115 (N_7115,N_5703,N_5050);
and U7116 (N_7116,N_4661,N_4357);
nand U7117 (N_7117,N_5389,N_4488);
and U7118 (N_7118,N_4623,N_4909);
and U7119 (N_7119,N_5115,N_4538);
and U7120 (N_7120,N_4719,N_4576);
and U7121 (N_7121,N_5500,N_5992);
or U7122 (N_7122,N_5091,N_5993);
nor U7123 (N_7123,N_5554,N_5908);
nor U7124 (N_7124,N_5198,N_4660);
or U7125 (N_7125,N_5895,N_5693);
and U7126 (N_7126,N_5009,N_4457);
nor U7127 (N_7127,N_5370,N_4828);
nand U7128 (N_7128,N_5288,N_5680);
nand U7129 (N_7129,N_5330,N_5528);
xnor U7130 (N_7130,N_4934,N_4549);
and U7131 (N_7131,N_5780,N_5954);
nand U7132 (N_7132,N_4127,N_5292);
and U7133 (N_7133,N_5491,N_4551);
or U7134 (N_7134,N_5097,N_4368);
xor U7135 (N_7135,N_5017,N_5026);
or U7136 (N_7136,N_5659,N_4629);
nor U7137 (N_7137,N_4101,N_4247);
nor U7138 (N_7138,N_5325,N_5704);
nand U7139 (N_7139,N_5146,N_5689);
or U7140 (N_7140,N_5860,N_4664);
nand U7141 (N_7141,N_4481,N_5503);
and U7142 (N_7142,N_5948,N_4547);
and U7143 (N_7143,N_5734,N_4416);
nand U7144 (N_7144,N_4256,N_5161);
nand U7145 (N_7145,N_5285,N_5774);
or U7146 (N_7146,N_4044,N_5801);
nor U7147 (N_7147,N_5142,N_4642);
and U7148 (N_7148,N_5473,N_5458);
nand U7149 (N_7149,N_4160,N_4679);
and U7150 (N_7150,N_5584,N_4255);
or U7151 (N_7151,N_5787,N_5591);
or U7152 (N_7152,N_4125,N_5980);
nand U7153 (N_7153,N_4437,N_4340);
or U7154 (N_7154,N_4758,N_4906);
nor U7155 (N_7155,N_4892,N_4594);
nand U7156 (N_7156,N_5325,N_5395);
nand U7157 (N_7157,N_4301,N_5724);
nand U7158 (N_7158,N_4003,N_5667);
and U7159 (N_7159,N_5478,N_4895);
nand U7160 (N_7160,N_5625,N_5401);
and U7161 (N_7161,N_5969,N_5740);
nand U7162 (N_7162,N_4639,N_4541);
nor U7163 (N_7163,N_5380,N_4973);
xor U7164 (N_7164,N_4205,N_5978);
or U7165 (N_7165,N_4261,N_5013);
or U7166 (N_7166,N_5422,N_5878);
xor U7167 (N_7167,N_5154,N_4306);
and U7168 (N_7168,N_5491,N_5788);
or U7169 (N_7169,N_4423,N_4024);
or U7170 (N_7170,N_4753,N_5165);
and U7171 (N_7171,N_4896,N_5473);
and U7172 (N_7172,N_4498,N_4214);
nor U7173 (N_7173,N_4914,N_5598);
and U7174 (N_7174,N_4745,N_4408);
nor U7175 (N_7175,N_5581,N_4539);
xor U7176 (N_7176,N_5852,N_4359);
or U7177 (N_7177,N_4958,N_4080);
or U7178 (N_7178,N_4016,N_5095);
and U7179 (N_7179,N_5795,N_5346);
nor U7180 (N_7180,N_5195,N_4270);
nor U7181 (N_7181,N_5466,N_4856);
and U7182 (N_7182,N_5794,N_5816);
nand U7183 (N_7183,N_5316,N_4872);
nand U7184 (N_7184,N_4632,N_5632);
nor U7185 (N_7185,N_5042,N_5050);
nor U7186 (N_7186,N_5893,N_4625);
nand U7187 (N_7187,N_4492,N_5251);
nand U7188 (N_7188,N_5368,N_4970);
and U7189 (N_7189,N_5646,N_5796);
nand U7190 (N_7190,N_4967,N_5690);
nor U7191 (N_7191,N_4977,N_5027);
or U7192 (N_7192,N_4902,N_5560);
or U7193 (N_7193,N_4921,N_5621);
nor U7194 (N_7194,N_4676,N_4604);
or U7195 (N_7195,N_5575,N_4775);
nor U7196 (N_7196,N_4026,N_4038);
nand U7197 (N_7197,N_5218,N_5372);
or U7198 (N_7198,N_4812,N_5621);
nor U7199 (N_7199,N_4251,N_5534);
and U7200 (N_7200,N_5738,N_4637);
or U7201 (N_7201,N_4925,N_4946);
nand U7202 (N_7202,N_5238,N_5203);
or U7203 (N_7203,N_5277,N_4180);
nand U7204 (N_7204,N_4370,N_5655);
and U7205 (N_7205,N_5231,N_4750);
nor U7206 (N_7206,N_5289,N_4350);
nor U7207 (N_7207,N_5505,N_4144);
nor U7208 (N_7208,N_5960,N_4987);
nand U7209 (N_7209,N_4903,N_4593);
or U7210 (N_7210,N_5505,N_5222);
or U7211 (N_7211,N_5138,N_4719);
nand U7212 (N_7212,N_4112,N_5025);
nand U7213 (N_7213,N_5457,N_5594);
or U7214 (N_7214,N_5006,N_5787);
nor U7215 (N_7215,N_4747,N_5809);
nand U7216 (N_7216,N_4289,N_5243);
or U7217 (N_7217,N_5182,N_5467);
nand U7218 (N_7218,N_4476,N_4996);
or U7219 (N_7219,N_5721,N_4799);
nor U7220 (N_7220,N_4117,N_4687);
and U7221 (N_7221,N_5460,N_4502);
or U7222 (N_7222,N_5292,N_5134);
and U7223 (N_7223,N_5316,N_4810);
or U7224 (N_7224,N_5904,N_5054);
nor U7225 (N_7225,N_4963,N_5214);
and U7226 (N_7226,N_5842,N_5099);
nor U7227 (N_7227,N_4112,N_5430);
nor U7228 (N_7228,N_5861,N_5023);
or U7229 (N_7229,N_4960,N_4385);
xor U7230 (N_7230,N_5027,N_4274);
or U7231 (N_7231,N_4187,N_4348);
nor U7232 (N_7232,N_4305,N_4779);
nor U7233 (N_7233,N_4744,N_5749);
and U7234 (N_7234,N_5106,N_4242);
nand U7235 (N_7235,N_4325,N_5183);
nor U7236 (N_7236,N_5567,N_4756);
nand U7237 (N_7237,N_4006,N_5749);
and U7238 (N_7238,N_5650,N_5534);
or U7239 (N_7239,N_5852,N_4756);
nor U7240 (N_7240,N_5178,N_4252);
or U7241 (N_7241,N_4649,N_5728);
nor U7242 (N_7242,N_4508,N_4028);
or U7243 (N_7243,N_4825,N_5567);
or U7244 (N_7244,N_5074,N_4758);
nor U7245 (N_7245,N_5231,N_4263);
and U7246 (N_7246,N_5843,N_5887);
and U7247 (N_7247,N_4281,N_4241);
nor U7248 (N_7248,N_4298,N_4771);
or U7249 (N_7249,N_4758,N_4563);
nor U7250 (N_7250,N_5220,N_4796);
or U7251 (N_7251,N_4262,N_5836);
or U7252 (N_7252,N_5900,N_5507);
nor U7253 (N_7253,N_5669,N_4187);
and U7254 (N_7254,N_5059,N_5844);
nand U7255 (N_7255,N_5481,N_4539);
and U7256 (N_7256,N_5007,N_5706);
nand U7257 (N_7257,N_4075,N_5595);
or U7258 (N_7258,N_5901,N_5368);
or U7259 (N_7259,N_4434,N_4371);
or U7260 (N_7260,N_5129,N_4194);
and U7261 (N_7261,N_4435,N_4858);
or U7262 (N_7262,N_4051,N_5318);
nor U7263 (N_7263,N_4762,N_5152);
nand U7264 (N_7264,N_4523,N_4616);
and U7265 (N_7265,N_5166,N_4021);
nand U7266 (N_7266,N_4122,N_4113);
xnor U7267 (N_7267,N_4205,N_4968);
or U7268 (N_7268,N_4342,N_5212);
and U7269 (N_7269,N_4492,N_4652);
and U7270 (N_7270,N_4471,N_4241);
or U7271 (N_7271,N_4488,N_4504);
or U7272 (N_7272,N_5516,N_5549);
and U7273 (N_7273,N_5125,N_5497);
nand U7274 (N_7274,N_4805,N_4822);
or U7275 (N_7275,N_4520,N_4645);
nand U7276 (N_7276,N_4111,N_4012);
nand U7277 (N_7277,N_5325,N_4324);
and U7278 (N_7278,N_5200,N_5580);
and U7279 (N_7279,N_5889,N_5794);
nor U7280 (N_7280,N_5773,N_5205);
nand U7281 (N_7281,N_4547,N_5735);
nor U7282 (N_7282,N_4156,N_4493);
nor U7283 (N_7283,N_4606,N_4644);
nor U7284 (N_7284,N_4759,N_4942);
or U7285 (N_7285,N_4362,N_5556);
nor U7286 (N_7286,N_5247,N_5786);
or U7287 (N_7287,N_4744,N_5668);
nand U7288 (N_7288,N_4892,N_5588);
and U7289 (N_7289,N_4472,N_4272);
or U7290 (N_7290,N_4738,N_5184);
nand U7291 (N_7291,N_5633,N_4813);
or U7292 (N_7292,N_5011,N_5064);
nand U7293 (N_7293,N_4307,N_5802);
xor U7294 (N_7294,N_5301,N_5792);
and U7295 (N_7295,N_4213,N_5470);
nor U7296 (N_7296,N_4600,N_4742);
and U7297 (N_7297,N_5168,N_5494);
or U7298 (N_7298,N_4963,N_5201);
nand U7299 (N_7299,N_4424,N_5388);
nand U7300 (N_7300,N_5766,N_5324);
nand U7301 (N_7301,N_4830,N_4577);
nor U7302 (N_7302,N_5391,N_5385);
nor U7303 (N_7303,N_5175,N_4371);
nand U7304 (N_7304,N_4325,N_5822);
nand U7305 (N_7305,N_4561,N_4599);
nor U7306 (N_7306,N_4245,N_5928);
and U7307 (N_7307,N_4754,N_4664);
and U7308 (N_7308,N_4416,N_4245);
nor U7309 (N_7309,N_4358,N_5513);
nor U7310 (N_7310,N_4931,N_5091);
and U7311 (N_7311,N_4471,N_4375);
or U7312 (N_7312,N_5823,N_5816);
nor U7313 (N_7313,N_4164,N_4194);
or U7314 (N_7314,N_5815,N_4004);
nand U7315 (N_7315,N_4199,N_5483);
or U7316 (N_7316,N_5614,N_5454);
or U7317 (N_7317,N_4865,N_5676);
or U7318 (N_7318,N_4686,N_5453);
and U7319 (N_7319,N_5662,N_4332);
and U7320 (N_7320,N_4883,N_4184);
nand U7321 (N_7321,N_4151,N_4304);
and U7322 (N_7322,N_4323,N_4808);
nand U7323 (N_7323,N_5297,N_5550);
and U7324 (N_7324,N_5154,N_5791);
or U7325 (N_7325,N_4953,N_5676);
nor U7326 (N_7326,N_5500,N_4431);
nand U7327 (N_7327,N_4001,N_5233);
nand U7328 (N_7328,N_4399,N_5587);
nor U7329 (N_7329,N_5421,N_5397);
nand U7330 (N_7330,N_5571,N_5962);
nor U7331 (N_7331,N_5609,N_4794);
nor U7332 (N_7332,N_4043,N_4061);
nand U7333 (N_7333,N_4557,N_5290);
or U7334 (N_7334,N_4983,N_4527);
and U7335 (N_7335,N_5170,N_5454);
nand U7336 (N_7336,N_4323,N_5099);
nor U7337 (N_7337,N_4831,N_4547);
nor U7338 (N_7338,N_4418,N_5622);
and U7339 (N_7339,N_5218,N_4835);
nor U7340 (N_7340,N_4098,N_4461);
and U7341 (N_7341,N_4072,N_4823);
nor U7342 (N_7342,N_5471,N_4056);
nor U7343 (N_7343,N_4125,N_4499);
nand U7344 (N_7344,N_4483,N_4858);
nand U7345 (N_7345,N_4275,N_5248);
or U7346 (N_7346,N_4266,N_5758);
nor U7347 (N_7347,N_5394,N_4977);
nor U7348 (N_7348,N_4739,N_4591);
nand U7349 (N_7349,N_4013,N_4390);
nor U7350 (N_7350,N_4162,N_5012);
nor U7351 (N_7351,N_5914,N_4424);
or U7352 (N_7352,N_4269,N_5783);
nor U7353 (N_7353,N_5413,N_4025);
nor U7354 (N_7354,N_5040,N_4684);
and U7355 (N_7355,N_5936,N_4164);
nand U7356 (N_7356,N_5775,N_5177);
nand U7357 (N_7357,N_5973,N_4380);
and U7358 (N_7358,N_5104,N_4116);
or U7359 (N_7359,N_5080,N_5981);
nor U7360 (N_7360,N_5064,N_4376);
or U7361 (N_7361,N_5518,N_5115);
nand U7362 (N_7362,N_4500,N_5594);
nand U7363 (N_7363,N_4470,N_5943);
xor U7364 (N_7364,N_4816,N_5877);
nor U7365 (N_7365,N_5372,N_5726);
and U7366 (N_7366,N_5384,N_4299);
and U7367 (N_7367,N_5236,N_4670);
and U7368 (N_7368,N_4132,N_5381);
and U7369 (N_7369,N_5377,N_5998);
and U7370 (N_7370,N_4863,N_4031);
and U7371 (N_7371,N_4602,N_4269);
nand U7372 (N_7372,N_4039,N_5498);
nor U7373 (N_7373,N_5470,N_5394);
nor U7374 (N_7374,N_5449,N_4873);
and U7375 (N_7375,N_5557,N_4447);
xnor U7376 (N_7376,N_5252,N_5164);
nor U7377 (N_7377,N_4086,N_4397);
and U7378 (N_7378,N_5172,N_5320);
or U7379 (N_7379,N_4191,N_5873);
or U7380 (N_7380,N_4026,N_5812);
and U7381 (N_7381,N_5054,N_4169);
or U7382 (N_7382,N_4318,N_5639);
nand U7383 (N_7383,N_4413,N_5204);
and U7384 (N_7384,N_4429,N_4089);
nand U7385 (N_7385,N_5935,N_5625);
nor U7386 (N_7386,N_5822,N_5131);
and U7387 (N_7387,N_5027,N_5033);
and U7388 (N_7388,N_5278,N_5175);
and U7389 (N_7389,N_5743,N_4924);
and U7390 (N_7390,N_4711,N_4351);
or U7391 (N_7391,N_4766,N_5231);
and U7392 (N_7392,N_5423,N_5210);
nand U7393 (N_7393,N_5904,N_5853);
nor U7394 (N_7394,N_4232,N_4675);
nand U7395 (N_7395,N_4722,N_4200);
and U7396 (N_7396,N_5078,N_4016);
nand U7397 (N_7397,N_5138,N_4571);
nor U7398 (N_7398,N_5068,N_5136);
nor U7399 (N_7399,N_4850,N_4127);
nor U7400 (N_7400,N_5017,N_4652);
or U7401 (N_7401,N_5326,N_4775);
and U7402 (N_7402,N_4273,N_5908);
and U7403 (N_7403,N_4486,N_4518);
or U7404 (N_7404,N_5973,N_4705);
nor U7405 (N_7405,N_5884,N_4648);
and U7406 (N_7406,N_4714,N_4347);
or U7407 (N_7407,N_4031,N_4063);
and U7408 (N_7408,N_4637,N_4160);
nor U7409 (N_7409,N_5984,N_4772);
or U7410 (N_7410,N_5698,N_4065);
nor U7411 (N_7411,N_4469,N_5391);
or U7412 (N_7412,N_4036,N_4249);
or U7413 (N_7413,N_4590,N_5254);
nand U7414 (N_7414,N_4061,N_4553);
nor U7415 (N_7415,N_4612,N_5840);
nor U7416 (N_7416,N_5274,N_4468);
or U7417 (N_7417,N_5702,N_5039);
nand U7418 (N_7418,N_5452,N_4074);
or U7419 (N_7419,N_5689,N_4157);
or U7420 (N_7420,N_4587,N_5371);
nor U7421 (N_7421,N_4432,N_4298);
nand U7422 (N_7422,N_5814,N_4509);
nor U7423 (N_7423,N_5242,N_4493);
or U7424 (N_7424,N_5011,N_4708);
nor U7425 (N_7425,N_5623,N_5943);
nor U7426 (N_7426,N_5192,N_5218);
nand U7427 (N_7427,N_5784,N_5912);
or U7428 (N_7428,N_5580,N_5655);
and U7429 (N_7429,N_4976,N_5327);
or U7430 (N_7430,N_5250,N_5139);
or U7431 (N_7431,N_5865,N_5568);
or U7432 (N_7432,N_4380,N_5800);
nor U7433 (N_7433,N_5908,N_4181);
nor U7434 (N_7434,N_5620,N_5062);
nand U7435 (N_7435,N_5863,N_4245);
nand U7436 (N_7436,N_5617,N_4347);
and U7437 (N_7437,N_5497,N_4705);
and U7438 (N_7438,N_4567,N_5719);
and U7439 (N_7439,N_4490,N_4364);
nor U7440 (N_7440,N_5995,N_5907);
nand U7441 (N_7441,N_4487,N_5803);
nor U7442 (N_7442,N_4722,N_4487);
nor U7443 (N_7443,N_5448,N_5903);
and U7444 (N_7444,N_5518,N_5330);
or U7445 (N_7445,N_4920,N_5946);
and U7446 (N_7446,N_5167,N_4137);
xor U7447 (N_7447,N_5750,N_4857);
nand U7448 (N_7448,N_5746,N_5046);
or U7449 (N_7449,N_4450,N_4539);
and U7450 (N_7450,N_5152,N_4266);
and U7451 (N_7451,N_4067,N_4995);
and U7452 (N_7452,N_5586,N_5227);
nand U7453 (N_7453,N_5775,N_5503);
nor U7454 (N_7454,N_4408,N_5150);
nor U7455 (N_7455,N_5478,N_4022);
or U7456 (N_7456,N_5956,N_4114);
or U7457 (N_7457,N_4183,N_4616);
or U7458 (N_7458,N_4281,N_4077);
and U7459 (N_7459,N_4870,N_4423);
nand U7460 (N_7460,N_4854,N_5895);
or U7461 (N_7461,N_4828,N_4759);
nand U7462 (N_7462,N_5304,N_4723);
or U7463 (N_7463,N_4642,N_4230);
nand U7464 (N_7464,N_5416,N_4169);
nand U7465 (N_7465,N_5886,N_5980);
and U7466 (N_7466,N_4244,N_4902);
nand U7467 (N_7467,N_4153,N_5603);
nor U7468 (N_7468,N_4205,N_5085);
or U7469 (N_7469,N_4536,N_4631);
nor U7470 (N_7470,N_4446,N_5351);
nor U7471 (N_7471,N_5732,N_4631);
or U7472 (N_7472,N_4398,N_5162);
nor U7473 (N_7473,N_5029,N_4426);
and U7474 (N_7474,N_5868,N_5511);
nand U7475 (N_7475,N_4589,N_4744);
xnor U7476 (N_7476,N_5500,N_5490);
nand U7477 (N_7477,N_4441,N_5628);
xor U7478 (N_7478,N_5537,N_4363);
and U7479 (N_7479,N_5413,N_4932);
and U7480 (N_7480,N_5288,N_4674);
or U7481 (N_7481,N_5388,N_5043);
nor U7482 (N_7482,N_4223,N_5191);
or U7483 (N_7483,N_4137,N_5800);
or U7484 (N_7484,N_4460,N_4934);
nor U7485 (N_7485,N_5710,N_5648);
nand U7486 (N_7486,N_4665,N_5144);
and U7487 (N_7487,N_4961,N_5591);
and U7488 (N_7488,N_5894,N_4717);
and U7489 (N_7489,N_5894,N_4081);
and U7490 (N_7490,N_5263,N_4810);
and U7491 (N_7491,N_4471,N_5051);
nand U7492 (N_7492,N_4924,N_4611);
and U7493 (N_7493,N_5535,N_4816);
nor U7494 (N_7494,N_5269,N_4139);
nand U7495 (N_7495,N_5289,N_5932);
nand U7496 (N_7496,N_4471,N_5204);
nor U7497 (N_7497,N_5756,N_4510);
nand U7498 (N_7498,N_5029,N_4410);
nor U7499 (N_7499,N_4239,N_5113);
or U7500 (N_7500,N_4262,N_4026);
nor U7501 (N_7501,N_4679,N_4193);
or U7502 (N_7502,N_5528,N_5191);
and U7503 (N_7503,N_5493,N_4192);
nor U7504 (N_7504,N_5737,N_5750);
or U7505 (N_7505,N_4144,N_4909);
and U7506 (N_7506,N_4523,N_4706);
nand U7507 (N_7507,N_5692,N_4669);
or U7508 (N_7508,N_5803,N_5841);
nor U7509 (N_7509,N_5510,N_4489);
or U7510 (N_7510,N_4875,N_5728);
or U7511 (N_7511,N_4450,N_4158);
and U7512 (N_7512,N_5758,N_4089);
and U7513 (N_7513,N_5659,N_5638);
and U7514 (N_7514,N_4337,N_5702);
nand U7515 (N_7515,N_4234,N_5731);
nor U7516 (N_7516,N_5966,N_4935);
and U7517 (N_7517,N_5601,N_5320);
xnor U7518 (N_7518,N_5751,N_5623);
nand U7519 (N_7519,N_4476,N_4744);
nand U7520 (N_7520,N_4751,N_4445);
nand U7521 (N_7521,N_4289,N_5700);
and U7522 (N_7522,N_4050,N_4268);
nand U7523 (N_7523,N_4988,N_4121);
or U7524 (N_7524,N_5876,N_5987);
nand U7525 (N_7525,N_5339,N_5030);
or U7526 (N_7526,N_5037,N_4677);
and U7527 (N_7527,N_4749,N_4198);
nor U7528 (N_7528,N_4813,N_5198);
or U7529 (N_7529,N_5218,N_5202);
nor U7530 (N_7530,N_4111,N_4314);
nor U7531 (N_7531,N_5835,N_5363);
or U7532 (N_7532,N_4309,N_4912);
nand U7533 (N_7533,N_5503,N_5078);
nor U7534 (N_7534,N_5958,N_4769);
nand U7535 (N_7535,N_4169,N_5658);
nand U7536 (N_7536,N_5494,N_4409);
xnor U7537 (N_7537,N_4108,N_5297);
nand U7538 (N_7538,N_5578,N_4596);
nand U7539 (N_7539,N_5471,N_5934);
nand U7540 (N_7540,N_5130,N_4669);
and U7541 (N_7541,N_5370,N_4845);
nor U7542 (N_7542,N_5559,N_4437);
and U7543 (N_7543,N_5568,N_5545);
and U7544 (N_7544,N_5229,N_5748);
and U7545 (N_7545,N_4962,N_4963);
and U7546 (N_7546,N_5145,N_5388);
or U7547 (N_7547,N_5419,N_4608);
nor U7548 (N_7548,N_5350,N_4886);
nor U7549 (N_7549,N_4969,N_4482);
or U7550 (N_7550,N_5334,N_5487);
nand U7551 (N_7551,N_5825,N_5919);
nand U7552 (N_7552,N_5563,N_5744);
and U7553 (N_7553,N_4230,N_4444);
nand U7554 (N_7554,N_4008,N_4998);
nand U7555 (N_7555,N_5232,N_5684);
and U7556 (N_7556,N_4926,N_4339);
nor U7557 (N_7557,N_4433,N_5726);
and U7558 (N_7558,N_5773,N_5449);
xnor U7559 (N_7559,N_5836,N_4697);
nor U7560 (N_7560,N_5922,N_4780);
nor U7561 (N_7561,N_4678,N_4645);
or U7562 (N_7562,N_4264,N_4958);
and U7563 (N_7563,N_4073,N_4387);
or U7564 (N_7564,N_5905,N_5093);
or U7565 (N_7565,N_5069,N_5642);
or U7566 (N_7566,N_4331,N_5102);
nor U7567 (N_7567,N_5109,N_5148);
nand U7568 (N_7568,N_4022,N_4389);
and U7569 (N_7569,N_4325,N_5545);
or U7570 (N_7570,N_4662,N_4638);
or U7571 (N_7571,N_5704,N_4404);
and U7572 (N_7572,N_5554,N_5102);
nand U7573 (N_7573,N_4600,N_4503);
nor U7574 (N_7574,N_4281,N_5424);
nand U7575 (N_7575,N_4158,N_5928);
and U7576 (N_7576,N_5138,N_5755);
or U7577 (N_7577,N_4445,N_5815);
and U7578 (N_7578,N_5098,N_5726);
or U7579 (N_7579,N_5567,N_4990);
or U7580 (N_7580,N_5981,N_5732);
nand U7581 (N_7581,N_4899,N_5645);
or U7582 (N_7582,N_4831,N_4797);
nor U7583 (N_7583,N_4806,N_5688);
nor U7584 (N_7584,N_5060,N_4054);
and U7585 (N_7585,N_4656,N_4236);
nand U7586 (N_7586,N_4146,N_5554);
or U7587 (N_7587,N_4030,N_5257);
or U7588 (N_7588,N_5956,N_4100);
nor U7589 (N_7589,N_5306,N_5678);
nor U7590 (N_7590,N_5034,N_5470);
or U7591 (N_7591,N_4253,N_5938);
xor U7592 (N_7592,N_5157,N_4743);
or U7593 (N_7593,N_4507,N_4475);
nor U7594 (N_7594,N_4392,N_5174);
nand U7595 (N_7595,N_5916,N_5042);
nand U7596 (N_7596,N_4029,N_4709);
nor U7597 (N_7597,N_5322,N_5970);
or U7598 (N_7598,N_4475,N_5583);
nor U7599 (N_7599,N_4113,N_4133);
nor U7600 (N_7600,N_5974,N_5038);
or U7601 (N_7601,N_4860,N_4146);
nand U7602 (N_7602,N_4142,N_4814);
nor U7603 (N_7603,N_5660,N_4230);
and U7604 (N_7604,N_4192,N_4400);
nand U7605 (N_7605,N_4422,N_4646);
or U7606 (N_7606,N_5380,N_5060);
nor U7607 (N_7607,N_4257,N_4821);
and U7608 (N_7608,N_4408,N_5524);
nor U7609 (N_7609,N_5539,N_4325);
nand U7610 (N_7610,N_4574,N_4856);
and U7611 (N_7611,N_5551,N_5991);
nand U7612 (N_7612,N_4510,N_5371);
or U7613 (N_7613,N_4553,N_5785);
or U7614 (N_7614,N_5623,N_4631);
nand U7615 (N_7615,N_5739,N_4500);
nor U7616 (N_7616,N_5114,N_4497);
or U7617 (N_7617,N_4422,N_5427);
nor U7618 (N_7618,N_5877,N_5849);
nand U7619 (N_7619,N_4221,N_4569);
nand U7620 (N_7620,N_4827,N_5336);
and U7621 (N_7621,N_4476,N_5024);
nand U7622 (N_7622,N_4573,N_4157);
nor U7623 (N_7623,N_5247,N_4538);
nand U7624 (N_7624,N_4379,N_5200);
nor U7625 (N_7625,N_5505,N_5135);
and U7626 (N_7626,N_4900,N_4643);
nor U7627 (N_7627,N_4996,N_5360);
and U7628 (N_7628,N_4033,N_5895);
nor U7629 (N_7629,N_5854,N_5131);
nand U7630 (N_7630,N_5971,N_4754);
nor U7631 (N_7631,N_4927,N_4891);
and U7632 (N_7632,N_4715,N_5248);
and U7633 (N_7633,N_5892,N_4325);
nand U7634 (N_7634,N_5005,N_5735);
or U7635 (N_7635,N_5680,N_4711);
nand U7636 (N_7636,N_5907,N_4870);
or U7637 (N_7637,N_4129,N_5702);
and U7638 (N_7638,N_5863,N_5233);
or U7639 (N_7639,N_4491,N_4807);
or U7640 (N_7640,N_5325,N_4042);
or U7641 (N_7641,N_4116,N_5015);
nor U7642 (N_7642,N_4650,N_5624);
and U7643 (N_7643,N_5754,N_5574);
nand U7644 (N_7644,N_5789,N_5691);
nor U7645 (N_7645,N_4146,N_4686);
nand U7646 (N_7646,N_4273,N_5465);
or U7647 (N_7647,N_4405,N_4512);
or U7648 (N_7648,N_5332,N_5252);
nor U7649 (N_7649,N_5990,N_4298);
or U7650 (N_7650,N_4413,N_4486);
or U7651 (N_7651,N_5865,N_5883);
or U7652 (N_7652,N_4581,N_4787);
or U7653 (N_7653,N_4368,N_5876);
nor U7654 (N_7654,N_4903,N_4932);
and U7655 (N_7655,N_5353,N_5206);
and U7656 (N_7656,N_4711,N_5132);
or U7657 (N_7657,N_4478,N_5107);
nand U7658 (N_7658,N_4212,N_4944);
nor U7659 (N_7659,N_4370,N_4676);
nand U7660 (N_7660,N_5470,N_4859);
or U7661 (N_7661,N_5070,N_4720);
nand U7662 (N_7662,N_5695,N_4801);
or U7663 (N_7663,N_4872,N_5285);
or U7664 (N_7664,N_5144,N_4051);
nor U7665 (N_7665,N_5875,N_5464);
and U7666 (N_7666,N_5213,N_4972);
and U7667 (N_7667,N_4222,N_4706);
and U7668 (N_7668,N_5175,N_4926);
and U7669 (N_7669,N_4555,N_5106);
or U7670 (N_7670,N_5691,N_4730);
xnor U7671 (N_7671,N_5492,N_4660);
or U7672 (N_7672,N_5038,N_4519);
nor U7673 (N_7673,N_4443,N_4342);
nand U7674 (N_7674,N_4658,N_4107);
nor U7675 (N_7675,N_5709,N_5453);
nand U7676 (N_7676,N_5033,N_5900);
or U7677 (N_7677,N_5076,N_4016);
and U7678 (N_7678,N_5390,N_4151);
or U7679 (N_7679,N_5268,N_4809);
nor U7680 (N_7680,N_5704,N_4652);
and U7681 (N_7681,N_5073,N_5435);
and U7682 (N_7682,N_5692,N_4107);
nor U7683 (N_7683,N_4285,N_4361);
or U7684 (N_7684,N_4710,N_5499);
and U7685 (N_7685,N_4210,N_4226);
or U7686 (N_7686,N_5932,N_4986);
and U7687 (N_7687,N_4489,N_4096);
nand U7688 (N_7688,N_5124,N_4481);
nor U7689 (N_7689,N_5646,N_5043);
nand U7690 (N_7690,N_5534,N_4459);
nand U7691 (N_7691,N_5408,N_5829);
nand U7692 (N_7692,N_4132,N_5206);
nor U7693 (N_7693,N_5077,N_5398);
or U7694 (N_7694,N_5880,N_5113);
or U7695 (N_7695,N_4769,N_4582);
and U7696 (N_7696,N_5953,N_4146);
or U7697 (N_7697,N_4322,N_4512);
nand U7698 (N_7698,N_4052,N_5665);
nand U7699 (N_7699,N_4914,N_4461);
nand U7700 (N_7700,N_5725,N_5769);
or U7701 (N_7701,N_4764,N_4818);
or U7702 (N_7702,N_5022,N_5895);
and U7703 (N_7703,N_4597,N_5430);
nor U7704 (N_7704,N_5073,N_4621);
nand U7705 (N_7705,N_5230,N_5867);
or U7706 (N_7706,N_4274,N_4362);
nor U7707 (N_7707,N_4275,N_5879);
or U7708 (N_7708,N_4729,N_4870);
and U7709 (N_7709,N_5827,N_5251);
nand U7710 (N_7710,N_5993,N_4763);
or U7711 (N_7711,N_4588,N_5242);
nand U7712 (N_7712,N_5842,N_5609);
nand U7713 (N_7713,N_4995,N_5476);
and U7714 (N_7714,N_5805,N_4458);
or U7715 (N_7715,N_4316,N_4865);
and U7716 (N_7716,N_5598,N_5626);
nand U7717 (N_7717,N_4119,N_5066);
or U7718 (N_7718,N_4887,N_4162);
or U7719 (N_7719,N_5054,N_5485);
and U7720 (N_7720,N_5236,N_5338);
and U7721 (N_7721,N_4004,N_5482);
nand U7722 (N_7722,N_5883,N_4049);
nand U7723 (N_7723,N_5009,N_5537);
xnor U7724 (N_7724,N_4511,N_4345);
nand U7725 (N_7725,N_5389,N_4126);
and U7726 (N_7726,N_4863,N_5217);
and U7727 (N_7727,N_4979,N_4997);
nand U7728 (N_7728,N_4739,N_5255);
nand U7729 (N_7729,N_4842,N_4278);
or U7730 (N_7730,N_5468,N_5983);
nand U7731 (N_7731,N_4958,N_4564);
and U7732 (N_7732,N_5628,N_4170);
xnor U7733 (N_7733,N_4059,N_5913);
nor U7734 (N_7734,N_5062,N_5560);
or U7735 (N_7735,N_5674,N_4011);
nand U7736 (N_7736,N_5960,N_5585);
nand U7737 (N_7737,N_5752,N_4834);
nor U7738 (N_7738,N_5736,N_4800);
or U7739 (N_7739,N_5256,N_5088);
and U7740 (N_7740,N_5235,N_5021);
and U7741 (N_7741,N_5353,N_5327);
nor U7742 (N_7742,N_5814,N_5672);
nand U7743 (N_7743,N_5728,N_4707);
or U7744 (N_7744,N_4732,N_5209);
and U7745 (N_7745,N_4548,N_4211);
or U7746 (N_7746,N_4946,N_5300);
or U7747 (N_7747,N_4009,N_4561);
nand U7748 (N_7748,N_5655,N_5726);
or U7749 (N_7749,N_5511,N_4252);
nand U7750 (N_7750,N_4778,N_5421);
or U7751 (N_7751,N_4760,N_5373);
nand U7752 (N_7752,N_5053,N_5273);
and U7753 (N_7753,N_5059,N_4867);
or U7754 (N_7754,N_4149,N_5543);
nand U7755 (N_7755,N_4784,N_5066);
nand U7756 (N_7756,N_5393,N_5825);
and U7757 (N_7757,N_5594,N_4491);
or U7758 (N_7758,N_4306,N_4508);
nor U7759 (N_7759,N_5456,N_5136);
and U7760 (N_7760,N_4508,N_4842);
xor U7761 (N_7761,N_4805,N_5949);
nor U7762 (N_7762,N_5223,N_4441);
and U7763 (N_7763,N_5161,N_4364);
and U7764 (N_7764,N_5662,N_5746);
and U7765 (N_7765,N_5054,N_5311);
and U7766 (N_7766,N_4867,N_4451);
nand U7767 (N_7767,N_4375,N_4932);
and U7768 (N_7768,N_4914,N_5856);
nor U7769 (N_7769,N_5909,N_4068);
nand U7770 (N_7770,N_4661,N_5996);
nand U7771 (N_7771,N_5021,N_4949);
nand U7772 (N_7772,N_4272,N_4415);
nand U7773 (N_7773,N_5686,N_5100);
and U7774 (N_7774,N_5564,N_4719);
and U7775 (N_7775,N_4730,N_5819);
and U7776 (N_7776,N_5736,N_5701);
and U7777 (N_7777,N_4203,N_4153);
and U7778 (N_7778,N_4726,N_5398);
and U7779 (N_7779,N_4412,N_5194);
nor U7780 (N_7780,N_5103,N_4488);
nand U7781 (N_7781,N_5951,N_4439);
nor U7782 (N_7782,N_4541,N_4494);
nand U7783 (N_7783,N_4983,N_4164);
nor U7784 (N_7784,N_5423,N_4421);
nor U7785 (N_7785,N_4814,N_5300);
nor U7786 (N_7786,N_4559,N_4674);
nor U7787 (N_7787,N_5250,N_5358);
xnor U7788 (N_7788,N_5112,N_5142);
and U7789 (N_7789,N_5809,N_5384);
and U7790 (N_7790,N_5554,N_5896);
or U7791 (N_7791,N_4813,N_5041);
nand U7792 (N_7792,N_4621,N_4520);
and U7793 (N_7793,N_5714,N_4895);
xnor U7794 (N_7794,N_5428,N_5386);
nand U7795 (N_7795,N_4225,N_4697);
and U7796 (N_7796,N_5838,N_4920);
nor U7797 (N_7797,N_5154,N_4684);
xnor U7798 (N_7798,N_4697,N_5461);
nand U7799 (N_7799,N_4530,N_4302);
nor U7800 (N_7800,N_5766,N_4923);
nand U7801 (N_7801,N_5954,N_5862);
nor U7802 (N_7802,N_5747,N_5485);
xor U7803 (N_7803,N_4628,N_4564);
or U7804 (N_7804,N_4184,N_4906);
or U7805 (N_7805,N_5501,N_4812);
or U7806 (N_7806,N_5905,N_4041);
nand U7807 (N_7807,N_4287,N_4266);
nor U7808 (N_7808,N_4300,N_4579);
and U7809 (N_7809,N_4395,N_4418);
and U7810 (N_7810,N_4678,N_4975);
nor U7811 (N_7811,N_4731,N_4391);
or U7812 (N_7812,N_5629,N_4005);
nand U7813 (N_7813,N_4518,N_5062);
nor U7814 (N_7814,N_4862,N_5618);
xnor U7815 (N_7815,N_4793,N_4896);
nand U7816 (N_7816,N_5270,N_4483);
nor U7817 (N_7817,N_4911,N_5867);
nand U7818 (N_7818,N_4365,N_4714);
nor U7819 (N_7819,N_5770,N_4578);
nor U7820 (N_7820,N_5781,N_4109);
nor U7821 (N_7821,N_4501,N_5615);
nand U7822 (N_7822,N_5711,N_4456);
or U7823 (N_7823,N_4793,N_4346);
or U7824 (N_7824,N_5076,N_5572);
and U7825 (N_7825,N_5565,N_4266);
nor U7826 (N_7826,N_4860,N_4612);
nand U7827 (N_7827,N_4782,N_4585);
or U7828 (N_7828,N_4560,N_5824);
and U7829 (N_7829,N_4402,N_4434);
and U7830 (N_7830,N_4340,N_5866);
nand U7831 (N_7831,N_4163,N_5737);
nand U7832 (N_7832,N_4890,N_4519);
and U7833 (N_7833,N_4577,N_5522);
nor U7834 (N_7834,N_4825,N_5633);
nor U7835 (N_7835,N_4789,N_5000);
nand U7836 (N_7836,N_4734,N_5196);
nand U7837 (N_7837,N_5001,N_4645);
nand U7838 (N_7838,N_5297,N_5764);
nand U7839 (N_7839,N_5539,N_5913);
and U7840 (N_7840,N_5132,N_4113);
or U7841 (N_7841,N_5983,N_5803);
or U7842 (N_7842,N_5701,N_5901);
nand U7843 (N_7843,N_4063,N_4794);
or U7844 (N_7844,N_4617,N_5746);
or U7845 (N_7845,N_5945,N_4219);
nand U7846 (N_7846,N_4017,N_4038);
nor U7847 (N_7847,N_5489,N_5171);
or U7848 (N_7848,N_4651,N_4185);
nand U7849 (N_7849,N_4582,N_5904);
or U7850 (N_7850,N_4617,N_4046);
and U7851 (N_7851,N_4812,N_5032);
nand U7852 (N_7852,N_5623,N_5739);
nand U7853 (N_7853,N_4160,N_5288);
nand U7854 (N_7854,N_5392,N_5497);
nand U7855 (N_7855,N_5983,N_4787);
or U7856 (N_7856,N_4759,N_5834);
or U7857 (N_7857,N_4825,N_4504);
nor U7858 (N_7858,N_5148,N_4323);
or U7859 (N_7859,N_5474,N_4262);
and U7860 (N_7860,N_4440,N_5107);
and U7861 (N_7861,N_5313,N_4153);
nor U7862 (N_7862,N_5296,N_4411);
nand U7863 (N_7863,N_5053,N_4552);
or U7864 (N_7864,N_5700,N_4533);
nand U7865 (N_7865,N_4736,N_5997);
or U7866 (N_7866,N_5684,N_5754);
nor U7867 (N_7867,N_4198,N_4454);
or U7868 (N_7868,N_5985,N_4434);
nand U7869 (N_7869,N_4391,N_5853);
nand U7870 (N_7870,N_5334,N_5802);
and U7871 (N_7871,N_4152,N_4801);
and U7872 (N_7872,N_5960,N_5063);
nand U7873 (N_7873,N_4752,N_5214);
nor U7874 (N_7874,N_5317,N_5991);
or U7875 (N_7875,N_4289,N_5454);
or U7876 (N_7876,N_4122,N_5069);
xor U7877 (N_7877,N_4462,N_5449);
or U7878 (N_7878,N_4748,N_4811);
nor U7879 (N_7879,N_4338,N_4217);
and U7880 (N_7880,N_4113,N_4203);
or U7881 (N_7881,N_4137,N_5405);
nand U7882 (N_7882,N_5282,N_4550);
nor U7883 (N_7883,N_5973,N_5460);
or U7884 (N_7884,N_4836,N_4194);
nor U7885 (N_7885,N_5808,N_4350);
or U7886 (N_7886,N_5450,N_4970);
xnor U7887 (N_7887,N_5536,N_5127);
nand U7888 (N_7888,N_5520,N_5594);
nand U7889 (N_7889,N_4595,N_5496);
nor U7890 (N_7890,N_4033,N_4131);
or U7891 (N_7891,N_4084,N_4888);
and U7892 (N_7892,N_5611,N_5017);
and U7893 (N_7893,N_4230,N_4214);
or U7894 (N_7894,N_4726,N_5593);
nor U7895 (N_7895,N_4693,N_4498);
and U7896 (N_7896,N_4861,N_4828);
nor U7897 (N_7897,N_5570,N_5212);
nand U7898 (N_7898,N_5253,N_5412);
or U7899 (N_7899,N_5893,N_5865);
nor U7900 (N_7900,N_5243,N_4122);
and U7901 (N_7901,N_5392,N_4835);
and U7902 (N_7902,N_5989,N_4738);
nand U7903 (N_7903,N_4375,N_5009);
and U7904 (N_7904,N_4639,N_5889);
or U7905 (N_7905,N_5436,N_5832);
nand U7906 (N_7906,N_4732,N_5737);
nand U7907 (N_7907,N_4488,N_4982);
and U7908 (N_7908,N_5810,N_4263);
nand U7909 (N_7909,N_4078,N_5688);
or U7910 (N_7910,N_5091,N_4351);
nand U7911 (N_7911,N_4365,N_5294);
nand U7912 (N_7912,N_4202,N_5129);
nand U7913 (N_7913,N_5530,N_4800);
xor U7914 (N_7914,N_4538,N_4629);
or U7915 (N_7915,N_4789,N_5498);
nor U7916 (N_7916,N_4390,N_4811);
nand U7917 (N_7917,N_4010,N_5739);
and U7918 (N_7918,N_5966,N_5048);
nand U7919 (N_7919,N_5538,N_4513);
and U7920 (N_7920,N_5812,N_4658);
nor U7921 (N_7921,N_4956,N_4050);
and U7922 (N_7922,N_5480,N_4376);
nand U7923 (N_7923,N_4701,N_4787);
and U7924 (N_7924,N_4051,N_4538);
or U7925 (N_7925,N_4515,N_4151);
and U7926 (N_7926,N_4976,N_4932);
or U7927 (N_7927,N_5232,N_5001);
or U7928 (N_7928,N_4033,N_5027);
nor U7929 (N_7929,N_5582,N_4723);
nor U7930 (N_7930,N_5194,N_4938);
nand U7931 (N_7931,N_5148,N_4719);
and U7932 (N_7932,N_4218,N_5343);
nand U7933 (N_7933,N_4827,N_5611);
or U7934 (N_7934,N_4086,N_5464);
and U7935 (N_7935,N_4118,N_5285);
nand U7936 (N_7936,N_5909,N_5995);
and U7937 (N_7937,N_5252,N_5351);
or U7938 (N_7938,N_4850,N_5230);
nand U7939 (N_7939,N_5265,N_5228);
nand U7940 (N_7940,N_4147,N_4379);
nor U7941 (N_7941,N_4802,N_4947);
or U7942 (N_7942,N_5818,N_5543);
nand U7943 (N_7943,N_4299,N_4343);
nand U7944 (N_7944,N_5196,N_4067);
and U7945 (N_7945,N_4271,N_5526);
nand U7946 (N_7946,N_5964,N_5729);
or U7947 (N_7947,N_5385,N_5969);
nor U7948 (N_7948,N_5567,N_4047);
nand U7949 (N_7949,N_5111,N_5062);
and U7950 (N_7950,N_4530,N_5850);
or U7951 (N_7951,N_5866,N_4402);
or U7952 (N_7952,N_4688,N_4159);
nand U7953 (N_7953,N_5889,N_5470);
nor U7954 (N_7954,N_5821,N_4904);
and U7955 (N_7955,N_5686,N_5404);
and U7956 (N_7956,N_5672,N_4560);
nand U7957 (N_7957,N_5042,N_4211);
nor U7958 (N_7958,N_5623,N_5368);
and U7959 (N_7959,N_5225,N_5328);
or U7960 (N_7960,N_4575,N_4483);
or U7961 (N_7961,N_4680,N_4105);
nor U7962 (N_7962,N_5264,N_4192);
nand U7963 (N_7963,N_4391,N_4315);
nor U7964 (N_7964,N_5842,N_4120);
and U7965 (N_7965,N_5560,N_5170);
or U7966 (N_7966,N_5621,N_5692);
or U7967 (N_7967,N_4751,N_4697);
or U7968 (N_7968,N_4424,N_4209);
and U7969 (N_7969,N_4279,N_5404);
and U7970 (N_7970,N_4391,N_5762);
or U7971 (N_7971,N_5847,N_5482);
nor U7972 (N_7972,N_4081,N_4461);
nand U7973 (N_7973,N_4101,N_4228);
nand U7974 (N_7974,N_5964,N_5198);
nor U7975 (N_7975,N_4983,N_4218);
nand U7976 (N_7976,N_5885,N_4166);
nor U7977 (N_7977,N_4833,N_5490);
or U7978 (N_7978,N_5841,N_4797);
and U7979 (N_7979,N_4531,N_5484);
or U7980 (N_7980,N_4668,N_4045);
xnor U7981 (N_7981,N_4466,N_5584);
nand U7982 (N_7982,N_4470,N_4996);
nand U7983 (N_7983,N_5820,N_4242);
and U7984 (N_7984,N_5614,N_5162);
and U7985 (N_7985,N_5007,N_4617);
or U7986 (N_7986,N_5551,N_4025);
and U7987 (N_7987,N_4324,N_5951);
or U7988 (N_7988,N_4256,N_5675);
or U7989 (N_7989,N_5354,N_4808);
nor U7990 (N_7990,N_4115,N_4364);
nand U7991 (N_7991,N_5544,N_4340);
nand U7992 (N_7992,N_4761,N_5648);
or U7993 (N_7993,N_4249,N_5332);
and U7994 (N_7994,N_4539,N_5097);
and U7995 (N_7995,N_5676,N_5432);
nor U7996 (N_7996,N_5573,N_4879);
nand U7997 (N_7997,N_5810,N_5464);
and U7998 (N_7998,N_4092,N_4255);
nor U7999 (N_7999,N_5707,N_4762);
or U8000 (N_8000,N_7417,N_7745);
nor U8001 (N_8001,N_7561,N_6097);
nand U8002 (N_8002,N_7785,N_7201);
nand U8003 (N_8003,N_7864,N_7845);
or U8004 (N_8004,N_6144,N_7323);
nand U8005 (N_8005,N_6584,N_7582);
nor U8006 (N_8006,N_6905,N_7757);
or U8007 (N_8007,N_6673,N_6727);
nand U8008 (N_8008,N_7709,N_7381);
or U8009 (N_8009,N_7400,N_6525);
and U8010 (N_8010,N_6627,N_6265);
or U8011 (N_8011,N_7355,N_6964);
and U8012 (N_8012,N_6882,N_6483);
xnor U8013 (N_8013,N_7199,N_6052);
nand U8014 (N_8014,N_6022,N_6896);
nor U8015 (N_8015,N_6261,N_6467);
nand U8016 (N_8016,N_6623,N_6900);
xor U8017 (N_8017,N_7444,N_6972);
or U8018 (N_8018,N_7200,N_7500);
nor U8019 (N_8019,N_6657,N_6267);
and U8020 (N_8020,N_6037,N_6557);
or U8021 (N_8021,N_6262,N_7599);
nand U8022 (N_8022,N_6899,N_6162);
and U8023 (N_8023,N_7795,N_6835);
or U8024 (N_8024,N_6621,N_7643);
or U8025 (N_8025,N_6614,N_7061);
and U8026 (N_8026,N_6661,N_6952);
xor U8027 (N_8027,N_6149,N_7779);
and U8028 (N_8028,N_7882,N_7507);
nand U8029 (N_8029,N_7235,N_6638);
nor U8030 (N_8030,N_7985,N_6220);
nor U8031 (N_8031,N_7987,N_6289);
and U8032 (N_8032,N_6444,N_7628);
and U8033 (N_8033,N_7145,N_7418);
or U8034 (N_8034,N_6577,N_7948);
nand U8035 (N_8035,N_7842,N_6868);
or U8036 (N_8036,N_7627,N_6282);
nor U8037 (N_8037,N_7176,N_7376);
and U8038 (N_8038,N_7256,N_7563);
nand U8039 (N_8039,N_7642,N_6030);
nand U8040 (N_8040,N_6885,N_6237);
and U8041 (N_8041,N_7553,N_7036);
and U8042 (N_8042,N_6151,N_6356);
nor U8043 (N_8043,N_7679,N_7680);
nand U8044 (N_8044,N_6758,N_6836);
or U8045 (N_8045,N_6302,N_6363);
nand U8046 (N_8046,N_6183,N_6209);
or U8047 (N_8047,N_7339,N_6537);
nor U8048 (N_8048,N_6995,N_6344);
nand U8049 (N_8049,N_7285,N_6333);
xnor U8050 (N_8050,N_6231,N_7347);
and U8051 (N_8051,N_7524,N_6032);
and U8052 (N_8052,N_7597,N_7241);
and U8053 (N_8053,N_6509,N_7917);
nor U8054 (N_8054,N_6970,N_7633);
nand U8055 (N_8055,N_6328,N_6874);
and U8056 (N_8056,N_6786,N_6315);
or U8057 (N_8057,N_7548,N_7172);
nor U8058 (N_8058,N_6240,N_6119);
nor U8059 (N_8059,N_6877,N_7203);
and U8060 (N_8060,N_6770,N_7932);
xnor U8061 (N_8061,N_6660,N_7844);
and U8062 (N_8062,N_6530,N_7452);
nand U8063 (N_8063,N_6454,N_6041);
and U8064 (N_8064,N_6983,N_7545);
or U8065 (N_8065,N_7294,N_6671);
nand U8066 (N_8066,N_7449,N_6646);
and U8067 (N_8067,N_6188,N_6173);
and U8068 (N_8068,N_6129,N_7622);
and U8069 (N_8069,N_7170,N_6539);
or U8070 (N_8070,N_6012,N_7330);
nand U8071 (N_8071,N_7003,N_7430);
nand U8072 (N_8072,N_7888,N_6494);
nand U8073 (N_8073,N_7740,N_6999);
nand U8074 (N_8074,N_6244,N_7856);
nand U8075 (N_8075,N_7445,N_7952);
or U8076 (N_8076,N_6980,N_6100);
nand U8077 (N_8077,N_7051,N_6820);
nor U8078 (N_8078,N_7152,N_7059);
and U8079 (N_8079,N_6171,N_7863);
xor U8080 (N_8080,N_7057,N_6146);
nor U8081 (N_8081,N_6784,N_6890);
nand U8082 (N_8082,N_6107,N_7154);
or U8083 (N_8083,N_7492,N_6611);
nand U8084 (N_8084,N_6926,N_6626);
or U8085 (N_8085,N_6254,N_7363);
nor U8086 (N_8086,N_7109,N_7988);
and U8087 (N_8087,N_6743,N_7615);
or U8088 (N_8088,N_7989,N_7516);
and U8089 (N_8089,N_6607,N_6834);
nor U8090 (N_8090,N_6086,N_7828);
or U8091 (N_8091,N_7189,N_6840);
nand U8092 (N_8092,N_6182,N_6250);
nand U8093 (N_8093,N_6515,N_6823);
or U8094 (N_8094,N_7926,N_6070);
nor U8095 (N_8095,N_7242,N_6213);
nand U8096 (N_8096,N_7192,N_6181);
nand U8097 (N_8097,N_6243,N_7372);
and U8098 (N_8098,N_6915,N_6347);
nor U8099 (N_8099,N_7941,N_7425);
or U8100 (N_8100,N_7881,N_7078);
or U8101 (N_8101,N_7494,N_6929);
and U8102 (N_8102,N_7832,N_6618);
and U8103 (N_8103,N_7664,N_6426);
or U8104 (N_8104,N_7440,N_7651);
xnor U8105 (N_8105,N_6637,N_7438);
xor U8106 (N_8106,N_7139,N_7861);
or U8107 (N_8107,N_6534,N_7065);
nor U8108 (N_8108,N_6585,N_6355);
nor U8109 (N_8109,N_6116,N_6691);
nor U8110 (N_8110,N_7284,N_7612);
nor U8111 (N_8111,N_6203,N_6844);
nor U8112 (N_8112,N_7132,N_6062);
nor U8113 (N_8113,N_7944,N_6536);
nand U8114 (N_8114,N_7534,N_6105);
or U8115 (N_8115,N_7510,N_6450);
nand U8116 (N_8116,N_7018,N_6441);
and U8117 (N_8117,N_7148,N_7860);
nor U8118 (N_8118,N_7117,N_7282);
and U8119 (N_8119,N_6471,N_7266);
nor U8120 (N_8120,N_7819,N_7865);
nor U8121 (N_8121,N_6279,N_6043);
or U8122 (N_8122,N_7685,N_7224);
or U8123 (N_8123,N_6291,N_6342);
or U8124 (N_8124,N_6791,N_6420);
nand U8125 (N_8125,N_6196,N_6520);
nor U8126 (N_8126,N_6879,N_7193);
or U8127 (N_8127,N_7435,N_6837);
nand U8128 (N_8128,N_6402,N_7890);
or U8129 (N_8129,N_7232,N_6438);
nand U8130 (N_8130,N_7055,N_7726);
nor U8131 (N_8131,N_7485,N_7105);
nand U8132 (N_8132,N_6499,N_6810);
or U8133 (N_8133,N_6506,N_6619);
nand U8134 (N_8134,N_7039,N_6772);
and U8135 (N_8135,N_7639,N_6424);
or U8136 (N_8136,N_6697,N_7473);
nor U8137 (N_8137,N_7806,N_6378);
nor U8138 (N_8138,N_6393,N_7854);
and U8139 (N_8139,N_7823,N_6716);
and U8140 (N_8140,N_7874,N_7370);
nand U8141 (N_8141,N_7060,N_6535);
or U8142 (N_8142,N_7840,N_6801);
and U8143 (N_8143,N_6689,N_6602);
nor U8144 (N_8144,N_7670,N_7312);
nand U8145 (N_8145,N_7401,N_6479);
nor U8146 (N_8146,N_7799,N_7541);
or U8147 (N_8147,N_6869,N_6497);
nand U8148 (N_8148,N_7737,N_7436);
and U8149 (N_8149,N_7990,N_6137);
nand U8150 (N_8150,N_7222,N_7247);
or U8151 (N_8151,N_6034,N_6398);
nor U8152 (N_8152,N_7134,N_6386);
nor U8153 (N_8153,N_7593,N_6551);
xnor U8154 (N_8154,N_7610,N_6913);
and U8155 (N_8155,N_7921,N_7912);
nor U8156 (N_8156,N_7489,N_6409);
nand U8157 (N_8157,N_6392,N_7813);
nor U8158 (N_8158,N_7653,N_6061);
nand U8159 (N_8159,N_6276,N_6475);
and U8160 (N_8160,N_6635,N_7246);
and U8161 (N_8161,N_7557,N_7163);
or U8162 (N_8162,N_6712,N_6897);
nand U8163 (N_8163,N_6531,N_7182);
or U8164 (N_8164,N_6588,N_6466);
and U8165 (N_8165,N_7778,N_7178);
nand U8166 (N_8166,N_6094,N_7868);
or U8167 (N_8167,N_7621,N_7136);
xor U8168 (N_8168,N_6726,N_7279);
nor U8169 (N_8169,N_7517,N_7578);
nor U8170 (N_8170,N_7360,N_7971);
nor U8171 (N_8171,N_6719,N_6808);
nor U8172 (N_8172,N_6396,N_7220);
or U8173 (N_8173,N_6527,N_6412);
nor U8174 (N_8174,N_6491,N_6880);
nand U8175 (N_8175,N_7515,N_7388);
and U8176 (N_8176,N_6616,N_7259);
nor U8177 (N_8177,N_6803,N_6851);
and U8178 (N_8178,N_6023,N_7816);
nand U8179 (N_8179,N_6709,N_7686);
or U8180 (N_8180,N_6361,N_6266);
nor U8181 (N_8181,N_7533,N_6906);
and U8182 (N_8182,N_7008,N_6039);
nor U8183 (N_8183,N_6961,N_7354);
nand U8184 (N_8184,N_6048,N_7433);
or U8185 (N_8185,N_7369,N_7329);
nand U8186 (N_8186,N_6457,N_6024);
xnor U8187 (N_8187,N_7466,N_7551);
and U8188 (N_8188,N_6156,N_7663);
and U8189 (N_8189,N_6830,N_6437);
and U8190 (N_8190,N_7001,N_6806);
and U8191 (N_8191,N_7684,N_6507);
nand U8192 (N_8192,N_6252,N_6035);
or U8193 (N_8193,N_6544,N_6538);
nand U8194 (N_8194,N_7103,N_6473);
and U8195 (N_8195,N_7211,N_6090);
nor U8196 (N_8196,N_6827,N_6902);
and U8197 (N_8197,N_6884,N_7245);
or U8198 (N_8198,N_6305,N_7046);
or U8199 (N_8199,N_7408,N_6297);
or U8200 (N_8200,N_7866,N_7565);
and U8201 (N_8201,N_6757,N_7775);
and U8202 (N_8202,N_7571,N_6284);
nand U8203 (N_8203,N_7817,N_6692);
nand U8204 (N_8204,N_7280,N_6793);
and U8205 (N_8205,N_6128,N_7542);
and U8206 (N_8206,N_6978,N_7287);
xnor U8207 (N_8207,N_6766,N_6994);
nand U8208 (N_8208,N_6925,N_6047);
nand U8209 (N_8209,N_7106,N_7601);
and U8210 (N_8210,N_6656,N_7855);
nand U8211 (N_8211,N_6389,N_6292);
and U8212 (N_8212,N_6528,N_6423);
and U8213 (N_8213,N_6664,N_6283);
nand U8214 (N_8214,N_7258,N_6492);
and U8215 (N_8215,N_7451,N_6632);
or U8216 (N_8216,N_7850,N_7594);
or U8217 (N_8217,N_7198,N_7315);
or U8218 (N_8218,N_6463,N_7755);
and U8219 (N_8219,N_6841,N_7085);
xor U8220 (N_8220,N_6734,N_7566);
nor U8221 (N_8221,N_7419,N_6434);
nor U8222 (N_8222,N_7540,N_7289);
and U8223 (N_8223,N_6891,N_7471);
and U8224 (N_8224,N_6832,N_7756);
nor U8225 (N_8225,N_7829,N_6595);
and U8226 (N_8226,N_7476,N_7646);
nand U8227 (N_8227,N_7420,N_6629);
nor U8228 (N_8228,N_6460,N_6735);
and U8229 (N_8229,N_6287,N_7387);
and U8230 (N_8230,N_6101,N_7288);
nor U8231 (N_8231,N_6374,N_6590);
nand U8232 (N_8232,N_7807,N_7093);
nor U8233 (N_8233,N_6911,N_6746);
nand U8234 (N_8234,N_7669,N_6939);
or U8235 (N_8235,N_7123,N_7486);
and U8236 (N_8236,N_7160,N_6802);
nor U8237 (N_8237,N_6390,N_7296);
or U8238 (N_8238,N_6990,N_7635);
or U8239 (N_8239,N_6833,N_6221);
xor U8240 (N_8240,N_6087,N_6521);
or U8241 (N_8241,N_6207,N_7812);
nor U8242 (N_8242,N_6445,N_7411);
or U8243 (N_8243,N_7527,N_7316);
nor U8244 (N_8244,N_7194,N_6927);
nor U8245 (N_8245,N_7503,N_6217);
or U8246 (N_8246,N_6367,N_6968);
and U8247 (N_8247,N_6433,N_7945);
and U8248 (N_8248,N_7512,N_6234);
and U8249 (N_8249,N_6651,N_6717);
and U8250 (N_8250,N_6280,N_6501);
nand U8251 (N_8251,N_6576,N_6688);
nand U8252 (N_8252,N_6916,N_7618);
nor U8253 (N_8253,N_6871,N_6125);
and U8254 (N_8254,N_7104,N_7272);
nand U8255 (N_8255,N_7069,N_7184);
nand U8256 (N_8256,N_6042,N_6788);
or U8257 (N_8257,N_6179,N_7760);
or U8258 (N_8258,N_7365,N_6225);
nand U8259 (N_8259,N_7770,N_7270);
or U8260 (N_8260,N_7777,N_6967);
or U8261 (N_8261,N_7077,N_7513);
or U8262 (N_8262,N_6776,N_6411);
and U8263 (N_8263,N_6326,N_6847);
nor U8264 (N_8264,N_7437,N_6645);
and U8265 (N_8265,N_7504,N_7919);
nor U8266 (N_8266,N_6824,N_7432);
and U8267 (N_8267,N_6351,N_7206);
nand U8268 (N_8268,N_7313,N_6379);
nor U8269 (N_8269,N_7402,N_6235);
or U8270 (N_8270,N_7787,N_7448);
nand U8271 (N_8271,N_6729,N_6942);
nand U8272 (N_8272,N_7037,N_7100);
or U8273 (N_8273,N_7719,N_7970);
and U8274 (N_8274,N_6920,N_6498);
and U8275 (N_8275,N_6761,N_7124);
or U8276 (N_8276,N_6003,N_6644);
nand U8277 (N_8277,N_6133,N_7058);
nand U8278 (N_8278,N_7028,N_6751);
and U8279 (N_8279,N_6931,N_7252);
or U8280 (N_8280,N_7386,N_7947);
and U8281 (N_8281,N_6640,N_6804);
nand U8282 (N_8282,N_7954,N_6436);
nor U8283 (N_8283,N_6831,N_6301);
and U8284 (N_8284,N_7572,N_7140);
nand U8285 (N_8285,N_7262,N_6598);
and U8286 (N_8286,N_7341,N_6192);
and U8287 (N_8287,N_6979,N_6600);
nor U8288 (N_8288,N_6860,N_6381);
and U8289 (N_8289,N_7962,N_6126);
nand U8290 (N_8290,N_7113,N_7422);
nor U8291 (N_8291,N_6687,N_6591);
nor U8292 (N_8292,N_7015,N_6084);
or U8293 (N_8293,N_7528,N_6033);
xnor U8294 (N_8294,N_7800,N_7676);
nor U8295 (N_8295,N_6069,N_7630);
nor U8296 (N_8296,N_6440,N_7324);
or U8297 (N_8297,N_7427,N_7293);
or U8298 (N_8298,N_6306,N_7616);
and U8299 (N_8299,N_6257,N_7478);
and U8300 (N_8300,N_7147,N_6345);
xor U8301 (N_8301,N_6936,N_7304);
nand U8302 (N_8302,N_6794,N_7054);
nand U8303 (N_8303,N_7302,N_7586);
nor U8304 (N_8304,N_6186,N_7543);
xnor U8305 (N_8305,N_7584,N_7730);
nor U8306 (N_8306,N_7733,N_7405);
nand U8307 (N_8307,N_6077,N_7887);
or U8308 (N_8308,N_6901,N_7218);
nor U8309 (N_8309,N_7407,N_7005);
and U8310 (N_8310,N_6655,N_6238);
xnor U8311 (N_8311,N_7116,N_7870);
and U8312 (N_8312,N_6988,N_6678);
nor U8313 (N_8313,N_7805,N_6917);
and U8314 (N_8314,N_7502,N_6731);
or U8315 (N_8315,N_7166,N_7072);
nand U8316 (N_8316,N_7511,N_6148);
or U8317 (N_8317,N_7763,N_7927);
nor U8318 (N_8318,N_6912,N_7464);
nor U8319 (N_8319,N_6013,N_7202);
nor U8320 (N_8320,N_6718,N_7552);
nor U8321 (N_8321,N_7849,N_7343);
or U8322 (N_8322,N_7276,N_7950);
and U8323 (N_8323,N_6405,N_7358);
nand U8324 (N_8324,N_6323,N_7942);
nor U8325 (N_8325,N_7644,N_6613);
nand U8326 (N_8326,N_7753,N_7858);
nor U8327 (N_8327,N_7403,N_6680);
or U8328 (N_8328,N_6856,N_6992);
nand U8329 (N_8329,N_6343,N_6317);
nor U8330 (N_8330,N_7914,N_7021);
xor U8331 (N_8331,N_6665,N_7221);
and U8332 (N_8332,N_6928,N_6248);
nor U8333 (N_8333,N_7080,N_6549);
and U8334 (N_8334,N_7611,N_7920);
nor U8335 (N_8335,N_6312,N_7275);
nor U8336 (N_8336,N_6063,N_7196);
or U8337 (N_8337,N_6058,N_7231);
or U8338 (N_8338,N_7470,N_7576);
and U8339 (N_8339,N_6937,N_6563);
nand U8340 (N_8340,N_7071,N_6040);
nand U8341 (N_8341,N_6511,N_7661);
nor U8342 (N_8342,N_6067,N_7838);
nor U8343 (N_8343,N_7993,N_7749);
and U8344 (N_8344,N_6908,N_7447);
nor U8345 (N_8345,N_6121,N_6950);
nor U8346 (N_8346,N_7050,N_7453);
or U8347 (N_8347,N_7596,N_7660);
and U8348 (N_8348,N_6857,N_7859);
nand U8349 (N_8349,N_6736,N_6522);
nor U8350 (N_8350,N_6303,N_7063);
or U8351 (N_8351,N_6459,N_6559);
or U8352 (N_8352,N_7769,N_7146);
nor U8353 (N_8353,N_7562,N_6117);
nand U8354 (N_8354,N_7320,N_6587);
nor U8355 (N_8355,N_7434,N_7450);
or U8356 (N_8356,N_6079,N_6747);
xnor U8357 (N_8357,N_6150,N_6956);
and U8358 (N_8358,N_7555,N_7857);
nand U8359 (N_8359,N_6449,N_7034);
or U8360 (N_8360,N_7558,N_7481);
nand U8361 (N_8361,N_7906,N_6469);
and U8362 (N_8362,N_7508,N_7340);
nand U8363 (N_8363,N_6997,N_7797);
or U8364 (N_8364,N_7491,N_7690);
nand U8365 (N_8365,N_7532,N_7269);
nor U8366 (N_8366,N_7695,N_7151);
nor U8367 (N_8367,N_6989,N_7301);
nand U8368 (N_8368,N_6304,N_7937);
or U8369 (N_8369,N_7271,N_6982);
and U8370 (N_8370,N_7815,N_7705);
or U8371 (N_8371,N_7094,N_6706);
and U8372 (N_8372,N_6206,N_6255);
nor U8373 (N_8373,N_7546,N_6603);
and U8374 (N_8374,N_7371,N_6205);
nand U8375 (N_8375,N_6812,N_7761);
and U8376 (N_8376,N_6199,N_6059);
nand U8377 (N_8377,N_6650,N_7885);
or U8378 (N_8378,N_7168,N_6858);
nor U8379 (N_8379,N_6759,N_7803);
xor U8380 (N_8380,N_7683,N_6892);
or U8381 (N_8381,N_7595,N_7722);
nor U8382 (N_8382,N_7591,N_7898);
nor U8383 (N_8383,N_7000,N_7424);
or U8384 (N_8384,N_6427,N_7847);
and U8385 (N_8385,N_6431,N_7326);
nor U8386 (N_8386,N_6211,N_7260);
or U8387 (N_8387,N_6329,N_7455);
nand U8388 (N_8388,N_7253,N_7714);
or U8389 (N_8389,N_6865,N_6241);
nand U8390 (N_8390,N_6115,N_6592);
or U8391 (N_8391,N_6748,N_6029);
or U8392 (N_8392,N_6031,N_7480);
nor U8393 (N_8393,N_7577,N_7299);
or U8394 (N_8394,N_6785,N_6822);
xor U8395 (N_8395,N_7580,N_7767);
and U8396 (N_8396,N_7096,N_7164);
or U8397 (N_8397,N_7910,N_7111);
nor U8398 (N_8398,N_7645,N_6078);
and U8399 (N_8399,N_6309,N_6318);
nand U8400 (N_8400,N_7338,N_6174);
nand U8401 (N_8401,N_6679,N_6051);
or U8402 (N_8402,N_7234,N_7590);
and U8403 (N_8403,N_6458,N_6991);
xor U8404 (N_8404,N_7053,N_6310);
nor U8405 (N_8405,N_6057,N_6876);
and U8406 (N_8406,N_6742,N_6705);
or U8407 (N_8407,N_7081,N_6930);
nand U8408 (N_8408,N_6505,N_7297);
nor U8409 (N_8409,N_6272,N_6286);
nand U8410 (N_8410,N_7531,N_7834);
and U8411 (N_8411,N_6099,N_6750);
and U8412 (N_8412,N_6805,N_6008);
and U8413 (N_8413,N_6773,N_7413);
and U8414 (N_8414,N_6014,N_6973);
xor U8415 (N_8415,N_7641,N_7752);
xnor U8416 (N_8416,N_6954,N_6215);
and U8417 (N_8417,N_6089,N_6778);
nand U8418 (N_8418,N_7088,N_6177);
or U8419 (N_8419,N_7782,N_7776);
or U8420 (N_8420,N_6566,N_7687);
and U8421 (N_8421,N_7658,N_7357);
or U8422 (N_8422,N_6634,N_6666);
nor U8423 (N_8423,N_6038,N_6532);
nand U8424 (N_8424,N_7802,N_6468);
or U8425 (N_8425,N_6581,N_6704);
or U8426 (N_8426,N_7934,N_7348);
and U8427 (N_8427,N_6797,N_6852);
nand U8428 (N_8428,N_7602,N_6648);
nand U8429 (N_8429,N_6569,N_6212);
or U8430 (N_8430,N_6339,N_6189);
nor U8431 (N_8431,N_7128,N_6922);
nor U8432 (N_8432,N_6417,N_6546);
or U8433 (N_8433,N_7579,N_6092);
nand U8434 (N_8434,N_6571,N_6826);
nand U8435 (N_8435,N_7022,N_7043);
nand U8436 (N_8436,N_6715,N_7366);
nor U8437 (N_8437,N_6518,N_7711);
or U8438 (N_8438,N_7723,N_7300);
nor U8439 (N_8439,N_6825,N_7846);
nor U8440 (N_8440,N_7309,N_7879);
nand U8441 (N_8441,N_7399,N_6075);
and U8442 (N_8442,N_7717,N_7165);
or U8443 (N_8443,N_7655,N_6543);
nand U8444 (N_8444,N_7613,N_7955);
and U8445 (N_8445,N_7237,N_6524);
nand U8446 (N_8446,N_6245,N_7463);
nand U8447 (N_8447,N_6288,N_6958);
and U8448 (N_8448,N_6932,N_7625);
or U8449 (N_8449,N_7731,N_6472);
and U8450 (N_8450,N_7998,N_7848);
nand U8451 (N_8451,N_7349,N_6817);
and U8452 (N_8452,N_7581,N_7040);
nor U8453 (N_8453,N_6914,N_6486);
or U8454 (N_8454,N_6085,N_7836);
nor U8455 (N_8455,N_6533,N_7689);
and U8456 (N_8456,N_7044,N_7662);
xnor U8457 (N_8457,N_6819,N_6728);
or U8458 (N_8458,N_6560,N_6815);
nand U8459 (N_8459,N_6300,N_7678);
nand U8460 (N_8460,N_7648,N_6790);
nor U8461 (N_8461,N_6098,N_6222);
or U8462 (N_8462,N_7283,N_7984);
or U8463 (N_8463,N_6275,N_6554);
or U8464 (N_8464,N_6110,N_6798);
nand U8465 (N_8465,N_6428,N_6768);
and U8466 (N_8466,N_7550,N_7383);
nand U8467 (N_8467,N_7897,N_7956);
and U8468 (N_8468,N_7791,N_6570);
or U8469 (N_8469,N_7536,N_6455);
nand U8470 (N_8470,N_6368,N_6017);
or U8471 (N_8471,N_6765,N_6385);
nand U8472 (N_8472,N_7671,N_6781);
or U8473 (N_8473,N_6432,N_7209);
nand U8474 (N_8474,N_7675,N_7390);
and U8475 (N_8475,N_7107,N_7479);
and U8476 (N_8476,N_7605,N_7102);
nand U8477 (N_8477,N_7014,N_7634);
or U8478 (N_8478,N_6382,N_7236);
or U8479 (N_8479,N_6160,N_6227);
and U8480 (N_8480,N_7310,N_7744);
and U8481 (N_8481,N_6131,N_6337);
nor U8482 (N_8482,N_7525,N_6552);
or U8483 (N_8483,N_7995,N_7238);
nor U8484 (N_8484,N_7949,N_7368);
nand U8485 (N_8485,N_6401,N_6404);
nor U8486 (N_8486,N_6375,N_7951);
nor U8487 (N_8487,N_6429,N_7725);
or U8488 (N_8488,N_6701,N_7395);
nand U8489 (N_8489,N_6631,N_7827);
nor U8490 (N_8490,N_6864,N_6529);
and U8491 (N_8491,N_6451,N_6608);
or U8492 (N_8492,N_6625,N_7682);
nor U8493 (N_8493,N_7484,N_7461);
and U8494 (N_8494,N_6465,N_6548);
and U8495 (N_8495,N_6482,N_6775);
nand U8496 (N_8496,N_7214,N_6955);
nor U8497 (N_8497,N_7378,N_6000);
nand U8498 (N_8498,N_6264,N_7361);
xor U8499 (N_8499,N_7045,N_6745);
nand U8500 (N_8500,N_7841,N_6753);
nand U8501 (N_8501,N_6159,N_6881);
or U8502 (N_8502,N_7911,N_6200);
and U8503 (N_8503,N_6064,N_7862);
nand U8504 (N_8504,N_6813,N_6145);
or U8505 (N_8505,N_7925,N_7884);
or U8506 (N_8506,N_6596,N_7090);
xnor U8507 (N_8507,N_7794,N_6060);
or U8508 (N_8508,N_6331,N_7367);
or U8509 (N_8509,N_6796,N_6346);
and U8510 (N_8510,N_6512,N_6088);
nand U8511 (N_8511,N_6258,N_7588);
and U8512 (N_8512,N_7308,N_6377);
nor U8513 (N_8513,N_7933,N_6456);
nand U8514 (N_8514,N_6523,N_6091);
nor U8515 (N_8515,N_7768,N_6723);
nand U8516 (N_8516,N_6582,N_7903);
nand U8517 (N_8517,N_6740,N_6232);
or U8518 (N_8518,N_7373,N_6943);
and U8519 (N_8519,N_6782,N_7344);
and U8520 (N_8520,N_7654,N_6178);
and U8521 (N_8521,N_6442,N_7598);
and U8522 (N_8522,N_7498,N_6792);
or U8523 (N_8523,N_6464,N_7924);
and U8524 (N_8524,N_7495,N_6859);
nor U8525 (N_8525,N_6118,N_7638);
nand U8526 (N_8526,N_6340,N_7943);
or U8527 (N_8527,N_7886,N_6918);
or U8528 (N_8528,N_7161,N_7788);
or U8529 (N_8529,N_6470,N_7587);
xor U8530 (N_8530,N_6136,N_6578);
nor U8531 (N_8531,N_6677,N_7624);
or U8532 (N_8532,N_7392,N_7334);
and U8533 (N_8533,N_6684,N_7936);
nand U8534 (N_8534,N_7734,N_6066);
nand U8535 (N_8535,N_6861,N_7465);
or U8536 (N_8536,N_6550,N_7889);
nor U8537 (N_8537,N_7336,N_6358);
nand U8538 (N_8538,N_7851,N_6488);
or U8539 (N_8539,N_7974,N_7243);
nor U8540 (N_8540,N_7292,N_6756);
and U8541 (N_8541,N_6606,N_6562);
nand U8542 (N_8542,N_7567,N_7380);
or U8543 (N_8543,N_6072,N_7204);
and U8544 (N_8544,N_7409,N_7820);
nor U8545 (N_8545,N_6223,N_7359);
nor U8546 (N_8546,N_7391,N_6294);
and U8547 (N_8547,N_7030,N_6821);
or U8548 (N_8548,N_7833,N_7674);
and U8549 (N_8549,N_7114,N_7712);
and U8550 (N_8550,N_6575,N_7207);
and U8551 (N_8551,N_6620,N_7426);
or U8552 (N_8552,N_6517,N_7773);
nand U8553 (N_8553,N_6026,N_6015);
and U8554 (N_8554,N_6081,N_7629);
or U8555 (N_8555,N_6744,N_6504);
nor U8556 (N_8556,N_7314,N_6839);
and U8557 (N_8557,N_6141,N_7322);
nor U8558 (N_8558,N_6185,N_7986);
nor U8559 (N_8559,N_7938,N_7876);
and U8560 (N_8560,N_7143,N_7458);
nor U8561 (N_8561,N_7382,N_6965);
and U8562 (N_8562,N_6953,N_6184);
and U8563 (N_8563,N_6829,N_7169);
nand U8564 (N_8564,N_7127,N_7319);
nor U8565 (N_8565,N_6319,N_7181);
nand U8566 (N_8566,N_7721,N_6711);
or U8567 (N_8567,N_7667,N_6695);
nor U8568 (N_8568,N_7261,N_6945);
or U8569 (N_8569,N_7122,N_6109);
and U8570 (N_8570,N_7278,N_7394);
nor U8571 (N_8571,N_6610,N_6663);
nor U8572 (N_8572,N_7101,N_6249);
nand U8573 (N_8573,N_7544,N_7443);
nand U8574 (N_8574,N_7979,N_7233);
or U8575 (N_8575,N_6210,N_7089);
nand U8576 (N_8576,N_7454,N_6332);
nand U8577 (N_8577,N_6894,N_6422);
nor U8578 (N_8578,N_7583,N_6269);
or U8579 (N_8579,N_6049,N_6721);
nand U8580 (N_8580,N_6573,N_6866);
nand U8581 (N_8581,N_6397,N_7575);
nor U8582 (N_8582,N_6561,N_7377);
nor U8583 (N_8583,N_7681,N_6541);
xor U8584 (N_8584,N_7083,N_7907);
nor U8585 (N_8585,N_6850,N_6435);
or U8586 (N_8586,N_7706,N_6124);
nand U8587 (N_8587,N_7404,N_6166);
nand U8588 (N_8588,N_6971,N_7569);
nor U8589 (N_8589,N_6594,N_6354);
or U8590 (N_8590,N_7529,N_6580);
or U8591 (N_8591,N_6986,N_7493);
and U8592 (N_8592,N_6046,N_6006);
and U8593 (N_8593,N_7537,N_7764);
or U8594 (N_8594,N_6845,N_6855);
and U8595 (N_8595,N_6251,N_6246);
nor U8596 (N_8596,N_6838,N_7969);
or U8597 (N_8597,N_6690,N_6807);
nor U8598 (N_8598,N_7789,N_7939);
and U8599 (N_8599,N_6263,N_6686);
nand U8600 (N_8600,N_6011,N_7904);
or U8601 (N_8601,N_6617,N_6242);
xnor U8602 (N_8602,N_6419,N_6018);
and U8603 (N_8603,N_6350,N_6353);
or U8604 (N_8604,N_6224,N_6702);
nor U8605 (N_8605,N_7830,N_7215);
nor U8606 (N_8606,N_7429,N_6553);
nor U8607 (N_8607,N_6233,N_7564);
and U8608 (N_8608,N_7843,N_7186);
or U8609 (N_8609,N_6313,N_7125);
and U8610 (N_8610,N_6642,N_7759);
nand U8611 (N_8611,N_7702,N_7032);
nor U8612 (N_8612,N_7477,N_6158);
nand U8613 (N_8613,N_7414,N_7307);
nor U8614 (N_8614,N_6140,N_6724);
or U8615 (N_8615,N_7728,N_7839);
nor U8616 (N_8616,N_7291,N_7707);
nor U8617 (N_8617,N_7968,N_7156);
or U8618 (N_8618,N_6583,N_6050);
and U8619 (N_8619,N_7724,N_6703);
or U8620 (N_8620,N_6643,N_7758);
or U8621 (N_8621,N_7345,N_7317);
nand U8622 (N_8622,N_6430,N_7428);
or U8623 (N_8623,N_6558,N_6338);
and U8624 (N_8624,N_6407,N_6814);
or U8625 (N_8625,N_7708,N_7356);
and U8626 (N_8626,N_6867,N_6762);
nor U8627 (N_8627,N_7880,N_7568);
and U8628 (N_8628,N_7474,N_7967);
nand U8629 (N_8629,N_6474,N_7902);
nor U8630 (N_8630,N_6854,N_6307);
and U8631 (N_8631,N_6846,N_7657);
nand U8632 (N_8632,N_7872,N_6828);
nor U8633 (N_8633,N_6247,N_6080);
and U8634 (N_8634,N_7126,N_6783);
and U8635 (N_8635,N_7157,N_7727);
xor U8636 (N_8636,N_6139,N_7002);
nor U8637 (N_8637,N_6947,N_6568);
nand U8638 (N_8638,N_6933,N_7075);
and U8639 (N_8639,N_6226,N_6780);
and U8640 (N_8640,N_6966,N_7523);
or U8641 (N_8641,N_7688,N_6779);
nand U8642 (N_8642,N_6487,N_7191);
or U8643 (N_8643,N_6019,N_7213);
or U8644 (N_8644,N_7891,N_7099);
and U8645 (N_8645,N_6764,N_7973);
or U8646 (N_8646,N_6659,N_7701);
and U8647 (N_8647,N_6274,N_7062);
or U8648 (N_8648,N_7738,N_6984);
nand U8649 (N_8649,N_6628,N_6114);
nand U8650 (N_8650,N_6230,N_6395);
nand U8651 (N_8651,N_6732,N_6599);
nand U8652 (N_8652,N_6708,N_7087);
or U8653 (N_8653,N_6669,N_6103);
nor U8654 (N_8654,N_7521,N_7487);
nand U8655 (N_8655,N_7327,N_6106);
nand U8656 (N_8656,N_6959,N_6510);
and U8657 (N_8657,N_6720,N_7007);
nor U8658 (N_8658,N_6478,N_6004);
and U8659 (N_8659,N_7423,N_7929);
and U8660 (N_8660,N_7374,N_7592);
nor U8661 (N_8661,N_7735,N_6229);
or U8662 (N_8662,N_6769,N_6073);
nor U8663 (N_8663,N_7064,N_7931);
or U8664 (N_8664,N_7389,N_6448);
and U8665 (N_8665,N_7765,N_7619);
nand U8666 (N_8666,N_7490,N_7264);
nor U8667 (N_8667,N_6285,N_6811);
or U8668 (N_8668,N_6681,N_7068);
nor U8669 (N_8669,N_7208,N_7048);
nand U8670 (N_8670,N_7636,N_7539);
nor U8671 (N_8671,N_7716,N_6002);
nor U8672 (N_8672,N_6239,N_6555);
and U8673 (N_8673,N_7350,N_7824);
and U8674 (N_8674,N_7137,N_6167);
nand U8675 (N_8675,N_7303,N_6887);
nor U8676 (N_8676,N_6924,N_7751);
nor U8677 (N_8677,N_6143,N_7940);
and U8678 (N_8678,N_7052,N_7640);
nor U8679 (N_8679,N_6904,N_7692);
nor U8680 (N_8680,N_6134,N_7780);
nor U8681 (N_8681,N_7809,N_7609);
xnor U8682 (N_8682,N_6169,N_6739);
nand U8683 (N_8683,N_7342,N_7187);
or U8684 (N_8684,N_7185,N_7456);
and U8685 (N_8685,N_6484,N_7649);
nor U8686 (N_8686,N_7556,N_6653);
xnor U8687 (N_8687,N_7346,N_6082);
and U8688 (N_8688,N_6612,N_7108);
nand U8689 (N_8689,N_7038,N_6104);
or U8690 (N_8690,N_6909,N_6093);
or U8691 (N_8691,N_6586,N_7098);
or U8692 (N_8692,N_7469,N_7110);
nor U8693 (N_8693,N_6308,N_7650);
nand U8694 (N_8694,N_7739,N_7010);
and U8695 (N_8695,N_7025,N_6574);
nor U8696 (N_8696,N_7410,N_7741);
and U8697 (N_8697,N_6699,N_7149);
and U8698 (N_8698,N_6074,N_7869);
or U8699 (N_8699,N_6195,N_6589);
nand U8700 (N_8700,N_6667,N_6025);
nand U8701 (N_8701,N_6204,N_6652);
nor U8702 (N_8702,N_7538,N_7697);
xor U8703 (N_8703,N_6198,N_7462);
nor U8704 (N_8704,N_7696,N_7808);
xnor U8705 (N_8705,N_6987,N_7781);
nand U8706 (N_8706,N_7996,N_6944);
nand U8707 (N_8707,N_7223,N_7875);
and U8708 (N_8708,N_6001,N_7549);
or U8709 (N_8709,N_6672,N_7167);
or U8710 (N_8710,N_6694,N_7659);
and U8711 (N_8711,N_7935,N_7029);
and U8712 (N_8712,N_6760,N_7626);
nor U8713 (N_8713,N_6311,N_6477);
and U8714 (N_8714,N_6502,N_7024);
or U8715 (N_8715,N_6883,N_7743);
and U8716 (N_8716,N_7180,N_7277);
or U8717 (N_8717,N_7699,N_7318);
nor U8718 (N_8718,N_7337,N_6675);
nor U8719 (N_8719,N_7905,N_7774);
nor U8720 (N_8720,N_6053,N_7239);
xnor U8721 (N_8721,N_6197,N_7131);
and U8722 (N_8722,N_7818,N_7026);
xnor U8723 (N_8723,N_7082,N_7923);
nor U8724 (N_8724,N_7519,N_6654);
nand U8725 (N_8725,N_6055,N_6028);
nor U8726 (N_8726,N_7506,N_6878);
or U8727 (N_8727,N_6508,N_7286);
or U8728 (N_8728,N_6996,N_7173);
and U8729 (N_8729,N_6767,N_6384);
or U8730 (N_8730,N_7518,N_6676);
nor U8731 (N_8731,N_6630,N_6934);
nand U8732 (N_8732,N_6165,N_7153);
and U8733 (N_8733,N_7019,N_6045);
nand U8734 (N_8734,N_6540,N_7608);
nor U8735 (N_8735,N_6376,N_7255);
nand U8736 (N_8736,N_6371,N_6636);
nand U8737 (N_8737,N_7793,N_7514);
nor U8738 (N_8738,N_6777,N_7188);
or U8739 (N_8739,N_7614,N_7023);
nor U8740 (N_8740,N_7130,N_7115);
nand U8741 (N_8741,N_6076,N_7992);
nand U8742 (N_8742,N_6774,N_7159);
and U8743 (N_8743,N_7631,N_7496);
or U8744 (N_8744,N_6674,N_6170);
nand U8745 (N_8745,N_7693,N_6519);
nor U8746 (N_8746,N_6495,N_6113);
or U8747 (N_8747,N_6010,N_6190);
and U8748 (N_8748,N_7305,N_7333);
or U8749 (N_8749,N_6919,N_6601);
or U8750 (N_8750,N_7240,N_6493);
and U8751 (N_8751,N_7306,N_6888);
or U8752 (N_8752,N_6341,N_6132);
nor U8753 (N_8753,N_6633,N_7617);
nand U8754 (N_8754,N_7746,N_7522);
nand U8755 (N_8755,N_7412,N_7195);
and U8756 (N_8756,N_7710,N_7831);
and U8757 (N_8757,N_6005,N_7298);
or U8758 (N_8758,N_7899,N_6921);
nor U8759 (N_8759,N_7754,N_7482);
nor U8760 (N_8760,N_7607,N_7011);
or U8761 (N_8761,N_6352,N_7908);
and U8762 (N_8762,N_6698,N_7895);
nand U8763 (N_8763,N_6490,N_6572);
or U8764 (N_8764,N_7766,N_6259);
and U8765 (N_8765,N_6216,N_7825);
nor U8766 (N_8766,N_7263,N_6175);
nand U8767 (N_8767,N_7406,N_6314);
nand U8768 (N_8768,N_7547,N_6324);
and U8769 (N_8769,N_7811,N_7585);
nand U8770 (N_8770,N_7467,N_7822);
nand U8771 (N_8771,N_7790,N_6949);
nand U8772 (N_8772,N_6579,N_6278);
or U8773 (N_8773,N_6281,N_7991);
nand U8774 (N_8774,N_6935,N_6157);
nor U8775 (N_8775,N_7729,N_7120);
or U8776 (N_8776,N_7017,N_7852);
or U8777 (N_8777,N_6903,N_7736);
and U8778 (N_8778,N_7249,N_7229);
nor U8779 (N_8779,N_6647,N_6154);
or U8780 (N_8780,N_6122,N_6842);
nand U8781 (N_8781,N_6977,N_7499);
or U8782 (N_8782,N_6180,N_7074);
nand U8783 (N_8783,N_6941,N_6176);
and U8784 (N_8784,N_6564,N_7798);
nor U8785 (N_8785,N_7248,N_7047);
or U8786 (N_8786,N_6208,N_6683);
nor U8787 (N_8787,N_7035,N_6380);
nor U8788 (N_8788,N_6293,N_7656);
nand U8789 (N_8789,N_7837,N_6071);
or U8790 (N_8790,N_7013,N_7994);
nor U8791 (N_8791,N_6714,N_6875);
or U8792 (N_8792,N_6489,N_6298);
nor U8793 (N_8793,N_7972,N_7073);
or U8794 (N_8794,N_6387,N_6271);
or U8795 (N_8795,N_7554,N_6795);
or U8796 (N_8796,N_6809,N_6056);
nand U8797 (N_8797,N_7980,N_7652);
or U8798 (N_8798,N_6268,N_7873);
nor U8799 (N_8799,N_6923,N_7632);
nand U8800 (N_8800,N_6481,N_6771);
nor U8801 (N_8801,N_6443,N_7027);
nand U8802 (N_8802,N_7623,N_7070);
or U8803 (N_8803,N_6526,N_6480);
xor U8804 (N_8804,N_7016,N_7530);
or U8805 (N_8805,N_7250,N_7677);
nor U8806 (N_8806,N_7953,N_6615);
or U8807 (N_8807,N_7928,N_6725);
and U8808 (N_8808,N_7505,N_7004);
nand U8809 (N_8809,N_6330,N_6334);
and U8810 (N_8810,N_7877,N_6439);
nand U8811 (N_8811,N_7698,N_7916);
nand U8812 (N_8812,N_7431,N_6194);
or U8813 (N_8813,N_7118,N_7909);
and U8814 (N_8814,N_6399,N_7265);
nand U8815 (N_8815,N_6083,N_7460);
and U8816 (N_8816,N_7396,N_7216);
and U8817 (N_8817,N_6009,N_6408);
or U8818 (N_8818,N_7210,N_6741);
nand U8819 (N_8819,N_7472,N_7978);
nor U8820 (N_8820,N_6191,N_7913);
and U8821 (N_8821,N_7574,N_6730);
or U8822 (N_8822,N_6693,N_6556);
and U8823 (N_8823,N_6976,N_6065);
or U8824 (N_8824,N_7012,N_6985);
nor U8825 (N_8825,N_7867,N_6322);
nor U8826 (N_8826,N_6641,N_7900);
and U8827 (N_8827,N_6737,N_6299);
and U8828 (N_8828,N_6296,N_6886);
or U8829 (N_8829,N_7079,N_7982);
nand U8830 (N_8830,N_7520,N_7295);
nand U8831 (N_8831,N_6516,N_6123);
and U8832 (N_8832,N_7896,N_7457);
or U8833 (N_8833,N_6135,N_7397);
or U8834 (N_8834,N_7031,N_7416);
nor U8835 (N_8835,N_7930,N_7804);
and U8836 (N_8836,N_6755,N_6605);
or U8837 (N_8837,N_7918,N_6138);
nand U8838 (N_8838,N_6400,N_6547);
nand U8839 (N_8839,N_7826,N_7006);
nor U8840 (N_8840,N_6670,N_6366);
nor U8841 (N_8841,N_7600,N_6889);
and U8842 (N_8842,N_7228,N_7589);
nor U8843 (N_8843,N_7393,N_6545);
nor U8844 (N_8844,N_7853,N_6446);
nor U8845 (N_8845,N_6410,N_7020);
or U8846 (N_8846,N_6349,N_6295);
and U8847 (N_8847,N_6848,N_7129);
nand U8848 (N_8848,N_6787,N_6102);
and U8849 (N_8849,N_6369,N_7475);
or U8850 (N_8850,N_7335,N_6290);
nand U8851 (N_8851,N_7049,N_7041);
and U8852 (N_8852,N_6496,N_7704);
nor U8853 (N_8853,N_6394,N_7121);
and U8854 (N_8854,N_7713,N_7810);
nor U8855 (N_8855,N_7442,N_6096);
and U8856 (N_8856,N_6108,N_6476);
nand U8857 (N_8857,N_7033,N_7999);
and U8858 (N_8858,N_7915,N_6068);
nor U8859 (N_8859,N_6843,N_7009);
nand U8860 (N_8860,N_6219,N_7133);
and U8861 (N_8861,N_6696,N_6253);
and U8862 (N_8862,N_6622,N_6201);
nand U8863 (N_8863,N_7997,N_7961);
nor U8864 (N_8864,N_7742,N_7981);
or U8865 (N_8865,N_7963,N_6975);
and U8866 (N_8866,N_6940,N_6713);
and U8867 (N_8867,N_7092,N_7175);
or U8868 (N_8868,N_6514,N_7227);
or U8869 (N_8869,N_7497,N_6749);
nor U8870 (N_8870,N_7703,N_6799);
xor U8871 (N_8871,N_7353,N_6960);
nor U8872 (N_8872,N_7792,N_6542);
nand U8873 (N_8873,N_7446,N_7274);
nand U8874 (N_8874,N_7964,N_7892);
or U8875 (N_8875,N_7468,N_7084);
or U8876 (N_8876,N_7976,N_6816);
or U8877 (N_8877,N_6752,N_6127);
nor U8878 (N_8878,N_6365,N_6270);
nand U8879 (N_8879,N_7977,N_7604);
or U8880 (N_8880,N_6421,N_7067);
nand U8881 (N_8881,N_7119,N_7720);
nor U8882 (N_8882,N_6624,N_7526);
nand U8883 (N_8883,N_6155,N_7673);
nand U8884 (N_8884,N_6336,N_7441);
xor U8885 (N_8885,N_7732,N_6658);
xnor U8886 (N_8886,N_7351,N_6016);
and U8887 (N_8887,N_7573,N_6320);
and U8888 (N_8888,N_7691,N_7325);
or U8889 (N_8889,N_6370,N_7205);
and U8890 (N_8890,N_6951,N_6218);
or U8891 (N_8891,N_6316,N_7959);
nor U8892 (N_8892,N_6948,N_6403);
and U8893 (N_8893,N_6710,N_7966);
nor U8894 (N_8894,N_7281,N_6112);
or U8895 (N_8895,N_7385,N_6722);
nand U8896 (N_8896,N_7922,N_7273);
nand U8897 (N_8897,N_7190,N_6981);
and U8898 (N_8898,N_6565,N_6021);
and U8899 (N_8899,N_7066,N_7603);
nand U8900 (N_8900,N_7694,N_6153);
and U8901 (N_8901,N_7668,N_6391);
nor U8902 (N_8902,N_7150,N_6325);
nand U8903 (N_8903,N_6020,N_6228);
nor U8904 (N_8904,N_7217,N_6172);
nor U8905 (N_8905,N_6870,N_6388);
nor U8906 (N_8906,N_7251,N_6513);
nand U8907 (N_8907,N_7142,N_6962);
and U8908 (N_8908,N_6789,N_7056);
nor U8909 (N_8909,N_6872,N_7509);
or U8910 (N_8910,N_7946,N_6130);
and U8911 (N_8911,N_7748,N_6873);
and U8912 (N_8912,N_6853,N_7715);
or U8913 (N_8913,N_6327,N_6597);
nor U8914 (N_8914,N_7212,N_6974);
nand U8915 (N_8915,N_6256,N_6373);
nand U8916 (N_8916,N_7871,N_7975);
and U8917 (N_8917,N_7086,N_6500);
nand U8918 (N_8918,N_7267,N_6609);
or U8919 (N_8919,N_6733,N_6418);
nand U8920 (N_8920,N_7375,N_7535);
and U8921 (N_8921,N_6406,N_7112);
and U8922 (N_8922,N_7097,N_7364);
or U8923 (N_8923,N_6360,N_7700);
and U8924 (N_8924,N_6161,N_7162);
nor U8925 (N_8925,N_7901,N_7177);
nor U8926 (N_8926,N_7958,N_6036);
or U8927 (N_8927,N_6800,N_6277);
or U8928 (N_8928,N_7957,N_6593);
nor U8929 (N_8929,N_6054,N_7091);
and U8930 (N_8930,N_6447,N_6461);
nor U8931 (N_8931,N_6969,N_6946);
nand U8932 (N_8932,N_7762,N_7814);
nor U8933 (N_8933,N_6120,N_6818);
or U8934 (N_8934,N_6763,N_6357);
nand U8935 (N_8935,N_7620,N_6372);
or U8936 (N_8936,N_7771,N_7783);
or U8937 (N_8937,N_7328,N_7570);
or U8938 (N_8938,N_7894,N_7672);
or U8939 (N_8939,N_6898,N_6462);
and U8940 (N_8940,N_7488,N_7772);
and U8941 (N_8941,N_6998,N_7257);
nand U8942 (N_8942,N_6700,N_7362);
and U8943 (N_8943,N_6147,N_7747);
or U8944 (N_8944,N_6604,N_7784);
nand U8945 (N_8945,N_6754,N_6383);
and U8946 (N_8946,N_7415,N_7501);
nand U8947 (N_8947,N_6415,N_7197);
nand U8948 (N_8948,N_7560,N_7219);
nor U8949 (N_8949,N_7439,N_7384);
and U8950 (N_8950,N_7230,N_6993);
nor U8951 (N_8951,N_6202,N_6044);
and U8952 (N_8952,N_7801,N_6273);
and U8953 (N_8953,N_7421,N_6425);
nand U8954 (N_8954,N_6348,N_7965);
or U8955 (N_8955,N_7786,N_6187);
or U8956 (N_8956,N_6111,N_7483);
or U8957 (N_8957,N_7379,N_6685);
and U8958 (N_8958,N_7647,N_6863);
or U8959 (N_8959,N_7135,N_6142);
or U8960 (N_8960,N_7244,N_6662);
nor U8961 (N_8961,N_7352,N_6152);
nand U8962 (N_8962,N_7179,N_7559);
xnor U8963 (N_8963,N_6862,N_6214);
nand U8964 (N_8964,N_7331,N_7141);
and U8965 (N_8965,N_7138,N_6668);
and U8966 (N_8966,N_6163,N_6963);
xor U8967 (N_8967,N_6164,N_7332);
and U8968 (N_8968,N_7606,N_7796);
nand U8969 (N_8969,N_7878,N_6649);
nor U8970 (N_8970,N_6639,N_7718);
or U8971 (N_8971,N_7459,N_6359);
nor U8972 (N_8972,N_6193,N_7226);
and U8973 (N_8973,N_6567,N_6938);
nand U8974 (N_8974,N_7666,N_6452);
nor U8975 (N_8975,N_7155,N_6260);
and U8976 (N_8976,N_7290,N_7821);
and U8977 (N_8977,N_7076,N_6907);
nand U8978 (N_8978,N_7835,N_7171);
and U8979 (N_8979,N_7665,N_7398);
and U8980 (N_8980,N_7158,N_6335);
nand U8981 (N_8981,N_7225,N_6095);
nand U8982 (N_8982,N_6007,N_6682);
or U8983 (N_8983,N_6485,N_6416);
and U8984 (N_8984,N_7960,N_6414);
nor U8985 (N_8985,N_6707,N_6413);
nor U8986 (N_8986,N_7883,N_7254);
nor U8987 (N_8987,N_6168,N_7095);
and U8988 (N_8988,N_6027,N_6503);
or U8989 (N_8989,N_7042,N_6895);
nand U8990 (N_8990,N_7893,N_6453);
nor U8991 (N_8991,N_7311,N_6910);
nor U8992 (N_8992,N_7183,N_7144);
or U8993 (N_8993,N_7983,N_7268);
and U8994 (N_8994,N_6364,N_6738);
or U8995 (N_8995,N_6957,N_6362);
nand U8996 (N_8996,N_7637,N_7321);
nor U8997 (N_8997,N_6849,N_7750);
and U8998 (N_8998,N_6321,N_7174);
nor U8999 (N_8999,N_6236,N_6893);
and U9000 (N_9000,N_7877,N_6020);
nor U9001 (N_9001,N_7946,N_6306);
or U9002 (N_9002,N_6383,N_7039);
nor U9003 (N_9003,N_6632,N_6124);
nor U9004 (N_9004,N_6096,N_6019);
and U9005 (N_9005,N_6467,N_6192);
or U9006 (N_9006,N_7268,N_6051);
nand U9007 (N_9007,N_6696,N_6331);
nor U9008 (N_9008,N_7294,N_6980);
or U9009 (N_9009,N_7926,N_7612);
nand U9010 (N_9010,N_6937,N_7627);
and U9011 (N_9011,N_7703,N_7520);
and U9012 (N_9012,N_6424,N_7579);
nor U9013 (N_9013,N_7694,N_6595);
nor U9014 (N_9014,N_6641,N_6383);
and U9015 (N_9015,N_6017,N_7079);
or U9016 (N_9016,N_7921,N_6720);
and U9017 (N_9017,N_7621,N_6347);
nand U9018 (N_9018,N_7664,N_7318);
nand U9019 (N_9019,N_6230,N_7044);
and U9020 (N_9020,N_6371,N_6227);
nand U9021 (N_9021,N_6113,N_7001);
and U9022 (N_9022,N_7625,N_7703);
and U9023 (N_9023,N_7932,N_7519);
nor U9024 (N_9024,N_7791,N_7473);
nor U9025 (N_9025,N_7877,N_7739);
or U9026 (N_9026,N_7127,N_6344);
or U9027 (N_9027,N_6098,N_6131);
and U9028 (N_9028,N_6345,N_7721);
and U9029 (N_9029,N_7585,N_6870);
or U9030 (N_9030,N_6234,N_7550);
nor U9031 (N_9031,N_7475,N_6813);
nand U9032 (N_9032,N_6609,N_7981);
or U9033 (N_9033,N_6562,N_6051);
nand U9034 (N_9034,N_7036,N_6688);
and U9035 (N_9035,N_6151,N_7591);
or U9036 (N_9036,N_6761,N_7043);
or U9037 (N_9037,N_7736,N_7977);
nand U9038 (N_9038,N_6852,N_6137);
and U9039 (N_9039,N_6896,N_6593);
and U9040 (N_9040,N_7797,N_7828);
or U9041 (N_9041,N_6447,N_7638);
and U9042 (N_9042,N_7113,N_6839);
or U9043 (N_9043,N_7291,N_6600);
nor U9044 (N_9044,N_6712,N_7947);
nor U9045 (N_9045,N_7169,N_6211);
nand U9046 (N_9046,N_6187,N_7309);
and U9047 (N_9047,N_6522,N_6052);
xor U9048 (N_9048,N_7770,N_7744);
nor U9049 (N_9049,N_7726,N_6407);
nor U9050 (N_9050,N_7730,N_6046);
or U9051 (N_9051,N_7957,N_6553);
and U9052 (N_9052,N_6137,N_7148);
or U9053 (N_9053,N_6420,N_7180);
nor U9054 (N_9054,N_6001,N_6452);
nand U9055 (N_9055,N_6373,N_6007);
nand U9056 (N_9056,N_6505,N_7061);
or U9057 (N_9057,N_6463,N_6659);
and U9058 (N_9058,N_7005,N_6507);
nor U9059 (N_9059,N_7788,N_6850);
nand U9060 (N_9060,N_7086,N_7216);
nand U9061 (N_9061,N_7916,N_6451);
nand U9062 (N_9062,N_6334,N_6465);
and U9063 (N_9063,N_6304,N_7764);
nor U9064 (N_9064,N_6690,N_7723);
nor U9065 (N_9065,N_7250,N_6520);
nor U9066 (N_9066,N_6181,N_7584);
nor U9067 (N_9067,N_6666,N_7776);
nand U9068 (N_9068,N_6448,N_6477);
xor U9069 (N_9069,N_6030,N_7518);
and U9070 (N_9070,N_7227,N_7659);
nand U9071 (N_9071,N_6416,N_6564);
nand U9072 (N_9072,N_7584,N_6953);
and U9073 (N_9073,N_6913,N_6984);
nor U9074 (N_9074,N_6588,N_7778);
and U9075 (N_9075,N_6415,N_6463);
and U9076 (N_9076,N_7152,N_6759);
or U9077 (N_9077,N_7825,N_7836);
or U9078 (N_9078,N_7727,N_6782);
or U9079 (N_9079,N_6435,N_6534);
nor U9080 (N_9080,N_7067,N_7724);
and U9081 (N_9081,N_6344,N_7867);
nand U9082 (N_9082,N_7243,N_6248);
and U9083 (N_9083,N_7261,N_7489);
xor U9084 (N_9084,N_7676,N_7851);
nor U9085 (N_9085,N_7234,N_6384);
and U9086 (N_9086,N_7075,N_6614);
nor U9087 (N_9087,N_7109,N_7108);
and U9088 (N_9088,N_7414,N_7280);
and U9089 (N_9089,N_6806,N_7141);
or U9090 (N_9090,N_6124,N_7382);
nand U9091 (N_9091,N_6702,N_6326);
and U9092 (N_9092,N_6931,N_7802);
nand U9093 (N_9093,N_7672,N_6079);
or U9094 (N_9094,N_7839,N_6829);
nor U9095 (N_9095,N_7826,N_6620);
or U9096 (N_9096,N_6237,N_7450);
nor U9097 (N_9097,N_7573,N_7030);
nor U9098 (N_9098,N_7693,N_6346);
and U9099 (N_9099,N_7443,N_6333);
nand U9100 (N_9100,N_6980,N_6296);
nor U9101 (N_9101,N_6289,N_7664);
and U9102 (N_9102,N_6743,N_6846);
nor U9103 (N_9103,N_6030,N_7461);
nor U9104 (N_9104,N_6607,N_6516);
and U9105 (N_9105,N_7206,N_7197);
and U9106 (N_9106,N_6722,N_7659);
nand U9107 (N_9107,N_6979,N_6210);
nor U9108 (N_9108,N_7902,N_7596);
nor U9109 (N_9109,N_6702,N_7757);
nor U9110 (N_9110,N_7475,N_7970);
nor U9111 (N_9111,N_6695,N_7465);
nor U9112 (N_9112,N_7611,N_6679);
and U9113 (N_9113,N_7014,N_7466);
or U9114 (N_9114,N_7111,N_7309);
and U9115 (N_9115,N_6402,N_6715);
and U9116 (N_9116,N_6892,N_6500);
nand U9117 (N_9117,N_6481,N_7356);
nor U9118 (N_9118,N_7391,N_6431);
or U9119 (N_9119,N_7043,N_6751);
nor U9120 (N_9120,N_7913,N_7627);
and U9121 (N_9121,N_7041,N_7565);
nand U9122 (N_9122,N_6981,N_7435);
xnor U9123 (N_9123,N_7932,N_7498);
nand U9124 (N_9124,N_6346,N_7184);
or U9125 (N_9125,N_7821,N_6071);
or U9126 (N_9126,N_6477,N_7891);
and U9127 (N_9127,N_7705,N_7378);
nand U9128 (N_9128,N_6315,N_6435);
and U9129 (N_9129,N_7125,N_7983);
and U9130 (N_9130,N_6144,N_7356);
and U9131 (N_9131,N_6623,N_6086);
nor U9132 (N_9132,N_7198,N_7065);
nand U9133 (N_9133,N_6994,N_6899);
and U9134 (N_9134,N_7661,N_6927);
nor U9135 (N_9135,N_6721,N_6626);
nor U9136 (N_9136,N_7407,N_7263);
nand U9137 (N_9137,N_7381,N_7858);
nor U9138 (N_9138,N_6372,N_7349);
and U9139 (N_9139,N_7737,N_6536);
nor U9140 (N_9140,N_7160,N_7245);
or U9141 (N_9141,N_7621,N_7240);
nand U9142 (N_9142,N_7750,N_6176);
and U9143 (N_9143,N_7967,N_6325);
and U9144 (N_9144,N_7117,N_6135);
nand U9145 (N_9145,N_7267,N_6998);
nor U9146 (N_9146,N_6745,N_6471);
nor U9147 (N_9147,N_6997,N_7867);
and U9148 (N_9148,N_6144,N_6099);
and U9149 (N_9149,N_7782,N_6783);
and U9150 (N_9150,N_6724,N_6119);
or U9151 (N_9151,N_7131,N_7377);
and U9152 (N_9152,N_6375,N_6535);
nand U9153 (N_9153,N_7522,N_7806);
nor U9154 (N_9154,N_7223,N_7156);
or U9155 (N_9155,N_6989,N_7763);
nand U9156 (N_9156,N_7961,N_7655);
and U9157 (N_9157,N_7596,N_6473);
and U9158 (N_9158,N_7597,N_7486);
nand U9159 (N_9159,N_7894,N_7354);
nand U9160 (N_9160,N_7167,N_7816);
nand U9161 (N_9161,N_6360,N_6135);
and U9162 (N_9162,N_6953,N_7704);
nand U9163 (N_9163,N_7126,N_7607);
nor U9164 (N_9164,N_7549,N_7310);
or U9165 (N_9165,N_7478,N_6663);
or U9166 (N_9166,N_7385,N_7127);
and U9167 (N_9167,N_7374,N_7411);
nand U9168 (N_9168,N_7115,N_6709);
and U9169 (N_9169,N_7874,N_6263);
xor U9170 (N_9170,N_7140,N_6368);
or U9171 (N_9171,N_6596,N_6962);
nor U9172 (N_9172,N_7691,N_6906);
nand U9173 (N_9173,N_7354,N_7529);
nand U9174 (N_9174,N_6399,N_7410);
or U9175 (N_9175,N_7377,N_6202);
or U9176 (N_9176,N_7686,N_6186);
nor U9177 (N_9177,N_7878,N_6696);
and U9178 (N_9178,N_6673,N_7796);
nor U9179 (N_9179,N_6683,N_7375);
or U9180 (N_9180,N_7779,N_7990);
and U9181 (N_9181,N_7880,N_7918);
and U9182 (N_9182,N_7255,N_6273);
nand U9183 (N_9183,N_7169,N_7691);
and U9184 (N_9184,N_7292,N_7180);
and U9185 (N_9185,N_7088,N_6611);
nand U9186 (N_9186,N_6617,N_7687);
nor U9187 (N_9187,N_7452,N_7490);
and U9188 (N_9188,N_7883,N_7197);
and U9189 (N_9189,N_6594,N_6988);
nor U9190 (N_9190,N_7615,N_7763);
nor U9191 (N_9191,N_6592,N_7402);
nor U9192 (N_9192,N_6640,N_7371);
nor U9193 (N_9193,N_7381,N_7729);
nor U9194 (N_9194,N_6556,N_7000);
nand U9195 (N_9195,N_6093,N_7044);
nand U9196 (N_9196,N_6674,N_6533);
nand U9197 (N_9197,N_6654,N_7415);
or U9198 (N_9198,N_6170,N_6843);
and U9199 (N_9199,N_7013,N_7965);
or U9200 (N_9200,N_7367,N_6650);
nand U9201 (N_9201,N_6168,N_7455);
nor U9202 (N_9202,N_7608,N_7370);
or U9203 (N_9203,N_7981,N_7532);
nand U9204 (N_9204,N_6372,N_7859);
and U9205 (N_9205,N_6162,N_7220);
and U9206 (N_9206,N_7456,N_7554);
nor U9207 (N_9207,N_7537,N_7718);
and U9208 (N_9208,N_6249,N_7729);
and U9209 (N_9209,N_6313,N_6200);
and U9210 (N_9210,N_7783,N_6378);
nand U9211 (N_9211,N_6112,N_6198);
or U9212 (N_9212,N_7797,N_7590);
and U9213 (N_9213,N_7182,N_7436);
and U9214 (N_9214,N_7428,N_6290);
nand U9215 (N_9215,N_6520,N_7283);
or U9216 (N_9216,N_6009,N_7989);
and U9217 (N_9217,N_6210,N_6617);
and U9218 (N_9218,N_6231,N_7405);
nor U9219 (N_9219,N_6735,N_6744);
or U9220 (N_9220,N_7598,N_6050);
nand U9221 (N_9221,N_7817,N_7331);
nand U9222 (N_9222,N_7993,N_6491);
and U9223 (N_9223,N_6479,N_7399);
and U9224 (N_9224,N_6273,N_7814);
nand U9225 (N_9225,N_7907,N_6861);
and U9226 (N_9226,N_7270,N_6759);
nor U9227 (N_9227,N_7565,N_6004);
or U9228 (N_9228,N_6231,N_7978);
xnor U9229 (N_9229,N_7344,N_7302);
or U9230 (N_9230,N_7762,N_7765);
or U9231 (N_9231,N_6457,N_6545);
and U9232 (N_9232,N_6974,N_6537);
nor U9233 (N_9233,N_7528,N_6006);
nand U9234 (N_9234,N_6237,N_6451);
nand U9235 (N_9235,N_6551,N_7176);
or U9236 (N_9236,N_7952,N_7428);
nand U9237 (N_9237,N_6729,N_6420);
or U9238 (N_9238,N_7377,N_7361);
and U9239 (N_9239,N_6798,N_6643);
nand U9240 (N_9240,N_7586,N_6493);
nor U9241 (N_9241,N_6616,N_7891);
xnor U9242 (N_9242,N_6669,N_7946);
and U9243 (N_9243,N_6828,N_6609);
nor U9244 (N_9244,N_7021,N_7196);
nor U9245 (N_9245,N_6152,N_7809);
nor U9246 (N_9246,N_7521,N_7836);
or U9247 (N_9247,N_6621,N_6877);
nand U9248 (N_9248,N_7726,N_7215);
xor U9249 (N_9249,N_6995,N_7681);
and U9250 (N_9250,N_6604,N_7635);
nor U9251 (N_9251,N_7310,N_6094);
and U9252 (N_9252,N_7209,N_6639);
nor U9253 (N_9253,N_6426,N_6433);
and U9254 (N_9254,N_6896,N_7989);
nand U9255 (N_9255,N_7204,N_7814);
nor U9256 (N_9256,N_6267,N_6856);
and U9257 (N_9257,N_6743,N_7344);
nor U9258 (N_9258,N_6605,N_7485);
nor U9259 (N_9259,N_7483,N_7338);
or U9260 (N_9260,N_7459,N_6171);
and U9261 (N_9261,N_6871,N_6352);
or U9262 (N_9262,N_7890,N_7539);
and U9263 (N_9263,N_7207,N_6545);
nand U9264 (N_9264,N_6771,N_6748);
and U9265 (N_9265,N_7040,N_6114);
nor U9266 (N_9266,N_6518,N_6873);
nand U9267 (N_9267,N_7452,N_6375);
and U9268 (N_9268,N_7179,N_7870);
xnor U9269 (N_9269,N_6010,N_7510);
nor U9270 (N_9270,N_7125,N_7432);
nor U9271 (N_9271,N_6725,N_6087);
or U9272 (N_9272,N_7482,N_6441);
or U9273 (N_9273,N_7815,N_6273);
nand U9274 (N_9274,N_6934,N_6454);
or U9275 (N_9275,N_7108,N_7238);
or U9276 (N_9276,N_6967,N_6835);
or U9277 (N_9277,N_7207,N_7221);
nor U9278 (N_9278,N_6132,N_7021);
and U9279 (N_9279,N_6588,N_6133);
and U9280 (N_9280,N_6142,N_6605);
and U9281 (N_9281,N_6742,N_6633);
nand U9282 (N_9282,N_7958,N_6083);
and U9283 (N_9283,N_6739,N_6120);
or U9284 (N_9284,N_7265,N_6406);
and U9285 (N_9285,N_7435,N_6820);
nor U9286 (N_9286,N_6353,N_6765);
nand U9287 (N_9287,N_7078,N_7076);
xor U9288 (N_9288,N_6158,N_7210);
or U9289 (N_9289,N_7320,N_6354);
or U9290 (N_9290,N_7811,N_6762);
or U9291 (N_9291,N_6719,N_6205);
or U9292 (N_9292,N_7520,N_7963);
nand U9293 (N_9293,N_7197,N_7257);
nor U9294 (N_9294,N_6909,N_7764);
or U9295 (N_9295,N_6257,N_7574);
or U9296 (N_9296,N_7736,N_6652);
and U9297 (N_9297,N_7739,N_6106);
nand U9298 (N_9298,N_6588,N_6193);
nor U9299 (N_9299,N_6435,N_6536);
nor U9300 (N_9300,N_6279,N_7761);
or U9301 (N_9301,N_6181,N_6953);
nand U9302 (N_9302,N_7161,N_7814);
nor U9303 (N_9303,N_7186,N_6833);
nor U9304 (N_9304,N_7296,N_7952);
xor U9305 (N_9305,N_7600,N_6135);
nor U9306 (N_9306,N_6092,N_6325);
nor U9307 (N_9307,N_7671,N_7595);
or U9308 (N_9308,N_7245,N_7519);
or U9309 (N_9309,N_6054,N_6359);
nor U9310 (N_9310,N_7302,N_6003);
or U9311 (N_9311,N_6039,N_6566);
nand U9312 (N_9312,N_7462,N_7212);
nand U9313 (N_9313,N_7930,N_7634);
xnor U9314 (N_9314,N_6482,N_7337);
nand U9315 (N_9315,N_6378,N_6450);
or U9316 (N_9316,N_7010,N_7565);
and U9317 (N_9317,N_7443,N_7189);
or U9318 (N_9318,N_7580,N_7221);
or U9319 (N_9319,N_7270,N_6804);
nor U9320 (N_9320,N_6655,N_6572);
and U9321 (N_9321,N_7525,N_7250);
nand U9322 (N_9322,N_6300,N_7923);
nor U9323 (N_9323,N_6486,N_7242);
nand U9324 (N_9324,N_6279,N_6304);
and U9325 (N_9325,N_6845,N_7179);
and U9326 (N_9326,N_7579,N_6775);
or U9327 (N_9327,N_7475,N_6087);
and U9328 (N_9328,N_6416,N_7362);
and U9329 (N_9329,N_6160,N_6889);
nand U9330 (N_9330,N_6368,N_7716);
and U9331 (N_9331,N_7400,N_7468);
and U9332 (N_9332,N_7602,N_6257);
and U9333 (N_9333,N_6584,N_6302);
nor U9334 (N_9334,N_7324,N_7850);
nand U9335 (N_9335,N_7143,N_6722);
nand U9336 (N_9336,N_7862,N_7661);
nand U9337 (N_9337,N_6356,N_7520);
nand U9338 (N_9338,N_7300,N_6373);
and U9339 (N_9339,N_6425,N_7619);
nand U9340 (N_9340,N_6591,N_6043);
or U9341 (N_9341,N_6436,N_6671);
or U9342 (N_9342,N_6139,N_6091);
nand U9343 (N_9343,N_6419,N_7986);
or U9344 (N_9344,N_6935,N_7318);
or U9345 (N_9345,N_7792,N_7322);
or U9346 (N_9346,N_7771,N_6954);
and U9347 (N_9347,N_7074,N_6330);
nand U9348 (N_9348,N_6416,N_7749);
or U9349 (N_9349,N_7168,N_7266);
nor U9350 (N_9350,N_7523,N_6584);
and U9351 (N_9351,N_7322,N_7969);
nor U9352 (N_9352,N_6606,N_7293);
and U9353 (N_9353,N_6702,N_6420);
or U9354 (N_9354,N_6579,N_6244);
and U9355 (N_9355,N_7643,N_6114);
nor U9356 (N_9356,N_6259,N_6269);
nor U9357 (N_9357,N_6512,N_6288);
xor U9358 (N_9358,N_6855,N_6269);
and U9359 (N_9359,N_6033,N_6290);
or U9360 (N_9360,N_7687,N_6984);
or U9361 (N_9361,N_7584,N_7454);
nor U9362 (N_9362,N_6194,N_6515);
and U9363 (N_9363,N_6956,N_7911);
nor U9364 (N_9364,N_6300,N_7421);
nand U9365 (N_9365,N_6837,N_7460);
nor U9366 (N_9366,N_7875,N_7122);
nor U9367 (N_9367,N_7178,N_7543);
nand U9368 (N_9368,N_7741,N_6966);
nor U9369 (N_9369,N_7664,N_7180);
nand U9370 (N_9370,N_6280,N_6357);
and U9371 (N_9371,N_6250,N_7359);
and U9372 (N_9372,N_7550,N_6109);
nand U9373 (N_9373,N_7897,N_6633);
and U9374 (N_9374,N_7413,N_6501);
nand U9375 (N_9375,N_6964,N_6061);
and U9376 (N_9376,N_7792,N_6613);
or U9377 (N_9377,N_7544,N_7845);
or U9378 (N_9378,N_7132,N_6034);
or U9379 (N_9379,N_7756,N_6947);
nor U9380 (N_9380,N_7761,N_6648);
xnor U9381 (N_9381,N_6508,N_7963);
or U9382 (N_9382,N_6299,N_6684);
nand U9383 (N_9383,N_7741,N_6750);
xor U9384 (N_9384,N_7692,N_7919);
or U9385 (N_9385,N_7189,N_7008);
nor U9386 (N_9386,N_7940,N_6008);
or U9387 (N_9387,N_6143,N_6931);
and U9388 (N_9388,N_6007,N_7001);
or U9389 (N_9389,N_6395,N_7669);
nor U9390 (N_9390,N_7082,N_6887);
xor U9391 (N_9391,N_6924,N_6436);
and U9392 (N_9392,N_6630,N_7644);
and U9393 (N_9393,N_7952,N_7145);
and U9394 (N_9394,N_6914,N_7562);
nand U9395 (N_9395,N_6116,N_7355);
nor U9396 (N_9396,N_6311,N_6403);
nor U9397 (N_9397,N_7324,N_6676);
nor U9398 (N_9398,N_6949,N_6319);
and U9399 (N_9399,N_6508,N_6716);
or U9400 (N_9400,N_7517,N_6078);
or U9401 (N_9401,N_6045,N_7004);
nand U9402 (N_9402,N_6703,N_7109);
nor U9403 (N_9403,N_7340,N_6417);
or U9404 (N_9404,N_7686,N_6653);
nand U9405 (N_9405,N_6900,N_7878);
or U9406 (N_9406,N_7893,N_6225);
xnor U9407 (N_9407,N_6549,N_7381);
nor U9408 (N_9408,N_6985,N_7706);
nor U9409 (N_9409,N_7595,N_6041);
nor U9410 (N_9410,N_7132,N_7090);
and U9411 (N_9411,N_7232,N_6207);
and U9412 (N_9412,N_6324,N_7960);
or U9413 (N_9413,N_7296,N_7190);
xor U9414 (N_9414,N_6418,N_6833);
nor U9415 (N_9415,N_7707,N_6864);
nand U9416 (N_9416,N_6716,N_6091);
nand U9417 (N_9417,N_6115,N_7855);
and U9418 (N_9418,N_6330,N_6888);
nand U9419 (N_9419,N_7027,N_6971);
and U9420 (N_9420,N_6406,N_6991);
and U9421 (N_9421,N_7360,N_7052);
nor U9422 (N_9422,N_6422,N_6565);
or U9423 (N_9423,N_7583,N_6978);
nor U9424 (N_9424,N_7829,N_6912);
or U9425 (N_9425,N_6326,N_7590);
xor U9426 (N_9426,N_6528,N_7144);
or U9427 (N_9427,N_6951,N_7106);
nand U9428 (N_9428,N_7189,N_7992);
nand U9429 (N_9429,N_6077,N_6416);
and U9430 (N_9430,N_7316,N_6373);
xnor U9431 (N_9431,N_7703,N_7600);
or U9432 (N_9432,N_6199,N_6556);
nor U9433 (N_9433,N_7513,N_6462);
nand U9434 (N_9434,N_7112,N_6443);
or U9435 (N_9435,N_6636,N_6094);
or U9436 (N_9436,N_7934,N_6989);
nand U9437 (N_9437,N_7372,N_6835);
nand U9438 (N_9438,N_7029,N_6825);
nor U9439 (N_9439,N_7463,N_7341);
nor U9440 (N_9440,N_7088,N_6008);
nand U9441 (N_9441,N_6224,N_6237);
or U9442 (N_9442,N_6430,N_6813);
or U9443 (N_9443,N_7788,N_6653);
or U9444 (N_9444,N_6959,N_6347);
and U9445 (N_9445,N_6070,N_7451);
nand U9446 (N_9446,N_6194,N_6872);
nand U9447 (N_9447,N_7833,N_7108);
and U9448 (N_9448,N_6905,N_6263);
or U9449 (N_9449,N_6768,N_7704);
nor U9450 (N_9450,N_6671,N_7203);
and U9451 (N_9451,N_6612,N_6762);
or U9452 (N_9452,N_7519,N_7112);
or U9453 (N_9453,N_6919,N_7801);
or U9454 (N_9454,N_7383,N_6184);
or U9455 (N_9455,N_6588,N_6832);
and U9456 (N_9456,N_6701,N_6347);
nor U9457 (N_9457,N_7499,N_6318);
and U9458 (N_9458,N_7149,N_6007);
nand U9459 (N_9459,N_7427,N_7637);
nor U9460 (N_9460,N_6970,N_7702);
or U9461 (N_9461,N_6242,N_7263);
or U9462 (N_9462,N_6407,N_7956);
nor U9463 (N_9463,N_7113,N_7356);
and U9464 (N_9464,N_7888,N_6006);
nor U9465 (N_9465,N_7718,N_6055);
and U9466 (N_9466,N_6409,N_6515);
nor U9467 (N_9467,N_6519,N_7188);
and U9468 (N_9468,N_6551,N_6112);
nor U9469 (N_9469,N_7711,N_6760);
nor U9470 (N_9470,N_6691,N_7224);
or U9471 (N_9471,N_6793,N_6079);
nand U9472 (N_9472,N_7188,N_6549);
and U9473 (N_9473,N_7262,N_6955);
or U9474 (N_9474,N_6899,N_6276);
and U9475 (N_9475,N_7598,N_7795);
nand U9476 (N_9476,N_6068,N_6611);
or U9477 (N_9477,N_6278,N_7283);
nand U9478 (N_9478,N_6805,N_7948);
nor U9479 (N_9479,N_6056,N_6757);
or U9480 (N_9480,N_7782,N_7344);
and U9481 (N_9481,N_7260,N_7706);
nor U9482 (N_9482,N_7308,N_7254);
or U9483 (N_9483,N_7554,N_7689);
nor U9484 (N_9484,N_6907,N_6743);
or U9485 (N_9485,N_6458,N_6073);
or U9486 (N_9486,N_6130,N_7270);
nor U9487 (N_9487,N_7203,N_6436);
nor U9488 (N_9488,N_7383,N_6156);
nand U9489 (N_9489,N_6741,N_6066);
nand U9490 (N_9490,N_7617,N_6244);
or U9491 (N_9491,N_6962,N_7667);
and U9492 (N_9492,N_7242,N_7324);
nand U9493 (N_9493,N_6738,N_6513);
or U9494 (N_9494,N_6498,N_7504);
or U9495 (N_9495,N_6336,N_6840);
or U9496 (N_9496,N_7650,N_7416);
and U9497 (N_9497,N_6938,N_7097);
nor U9498 (N_9498,N_7862,N_7473);
nor U9499 (N_9499,N_6614,N_6865);
or U9500 (N_9500,N_7012,N_6863);
or U9501 (N_9501,N_6811,N_7027);
nand U9502 (N_9502,N_7664,N_7156);
nand U9503 (N_9503,N_6080,N_6297);
xor U9504 (N_9504,N_7859,N_7183);
and U9505 (N_9505,N_7543,N_6719);
and U9506 (N_9506,N_7318,N_6613);
nor U9507 (N_9507,N_7173,N_6976);
nor U9508 (N_9508,N_6878,N_7395);
or U9509 (N_9509,N_7642,N_6786);
nand U9510 (N_9510,N_7797,N_6095);
or U9511 (N_9511,N_6851,N_7512);
nor U9512 (N_9512,N_6905,N_6398);
and U9513 (N_9513,N_7554,N_6770);
nor U9514 (N_9514,N_7686,N_6006);
and U9515 (N_9515,N_7784,N_6561);
and U9516 (N_9516,N_6205,N_7241);
nor U9517 (N_9517,N_6086,N_7695);
nand U9518 (N_9518,N_7432,N_7630);
or U9519 (N_9519,N_7725,N_6340);
or U9520 (N_9520,N_6450,N_7532);
and U9521 (N_9521,N_7636,N_7993);
nor U9522 (N_9522,N_6669,N_7381);
nand U9523 (N_9523,N_6322,N_6525);
and U9524 (N_9524,N_7404,N_6725);
nor U9525 (N_9525,N_6007,N_7924);
nand U9526 (N_9526,N_7945,N_7674);
or U9527 (N_9527,N_7077,N_6018);
nand U9528 (N_9528,N_6854,N_6153);
nand U9529 (N_9529,N_6403,N_6911);
nor U9530 (N_9530,N_7627,N_7663);
or U9531 (N_9531,N_7832,N_6376);
nand U9532 (N_9532,N_7583,N_6099);
nor U9533 (N_9533,N_6096,N_7901);
or U9534 (N_9534,N_7820,N_6034);
nand U9535 (N_9535,N_7110,N_6796);
nor U9536 (N_9536,N_7548,N_7174);
or U9537 (N_9537,N_7638,N_7941);
nor U9538 (N_9538,N_6632,N_6508);
nand U9539 (N_9539,N_6358,N_7558);
xnor U9540 (N_9540,N_7219,N_7908);
nor U9541 (N_9541,N_6101,N_6700);
or U9542 (N_9542,N_7354,N_6055);
nor U9543 (N_9543,N_6704,N_6433);
nor U9544 (N_9544,N_6483,N_6800);
nor U9545 (N_9545,N_6565,N_7804);
and U9546 (N_9546,N_7425,N_7785);
or U9547 (N_9547,N_7066,N_7921);
and U9548 (N_9548,N_7660,N_6704);
or U9549 (N_9549,N_7890,N_7991);
nor U9550 (N_9550,N_7322,N_7351);
or U9551 (N_9551,N_6715,N_6775);
nand U9552 (N_9552,N_7571,N_6432);
nor U9553 (N_9553,N_7329,N_6203);
nand U9554 (N_9554,N_7676,N_7106);
nor U9555 (N_9555,N_6068,N_6935);
nor U9556 (N_9556,N_7843,N_7279);
nand U9557 (N_9557,N_6479,N_6100);
and U9558 (N_9558,N_7916,N_7768);
nor U9559 (N_9559,N_7656,N_6391);
and U9560 (N_9560,N_7538,N_7212);
nand U9561 (N_9561,N_6873,N_7055);
nor U9562 (N_9562,N_6539,N_6828);
nor U9563 (N_9563,N_6368,N_6414);
nor U9564 (N_9564,N_7671,N_7144);
or U9565 (N_9565,N_6714,N_7784);
and U9566 (N_9566,N_7752,N_6086);
nand U9567 (N_9567,N_7703,N_6384);
and U9568 (N_9568,N_6636,N_7575);
and U9569 (N_9569,N_7375,N_6992);
nor U9570 (N_9570,N_7403,N_6060);
nand U9571 (N_9571,N_7112,N_7371);
nor U9572 (N_9572,N_6072,N_7220);
nand U9573 (N_9573,N_7163,N_6854);
nand U9574 (N_9574,N_7457,N_7128);
or U9575 (N_9575,N_6351,N_7667);
or U9576 (N_9576,N_7397,N_7868);
nor U9577 (N_9577,N_7534,N_6217);
nand U9578 (N_9578,N_7914,N_7217);
or U9579 (N_9579,N_7173,N_7666);
nand U9580 (N_9580,N_7513,N_6654);
and U9581 (N_9581,N_7501,N_7689);
nor U9582 (N_9582,N_6130,N_7751);
nor U9583 (N_9583,N_6488,N_7832);
and U9584 (N_9584,N_6483,N_7787);
nor U9585 (N_9585,N_6008,N_6906);
xor U9586 (N_9586,N_7389,N_6677);
xnor U9587 (N_9587,N_6197,N_6230);
or U9588 (N_9588,N_7056,N_7843);
or U9589 (N_9589,N_6309,N_6760);
xnor U9590 (N_9590,N_6059,N_6782);
and U9591 (N_9591,N_6417,N_7345);
nor U9592 (N_9592,N_6647,N_7036);
xnor U9593 (N_9593,N_7929,N_7760);
and U9594 (N_9594,N_6929,N_7197);
and U9595 (N_9595,N_6748,N_6933);
or U9596 (N_9596,N_6006,N_7480);
nand U9597 (N_9597,N_6746,N_6088);
or U9598 (N_9598,N_7156,N_6160);
and U9599 (N_9599,N_7151,N_7769);
or U9600 (N_9600,N_6886,N_7087);
nand U9601 (N_9601,N_6685,N_6835);
nand U9602 (N_9602,N_7000,N_7799);
and U9603 (N_9603,N_6807,N_7622);
nand U9604 (N_9604,N_7449,N_7112);
or U9605 (N_9605,N_6850,N_6398);
and U9606 (N_9606,N_6375,N_6295);
nand U9607 (N_9607,N_7080,N_6087);
or U9608 (N_9608,N_6502,N_6573);
xnor U9609 (N_9609,N_6531,N_6747);
nor U9610 (N_9610,N_7589,N_7676);
nor U9611 (N_9611,N_7069,N_7901);
xor U9612 (N_9612,N_7884,N_7127);
nor U9613 (N_9613,N_7296,N_6115);
or U9614 (N_9614,N_7337,N_7678);
nor U9615 (N_9615,N_7926,N_6708);
nand U9616 (N_9616,N_6186,N_7914);
xor U9617 (N_9617,N_6574,N_6566);
nor U9618 (N_9618,N_6830,N_6097);
and U9619 (N_9619,N_6733,N_6460);
nand U9620 (N_9620,N_7836,N_7190);
and U9621 (N_9621,N_6556,N_6622);
and U9622 (N_9622,N_7080,N_7917);
nor U9623 (N_9623,N_6298,N_7023);
nor U9624 (N_9624,N_6151,N_7667);
and U9625 (N_9625,N_7807,N_7515);
and U9626 (N_9626,N_7084,N_7603);
and U9627 (N_9627,N_7143,N_7124);
nand U9628 (N_9628,N_6281,N_6704);
nand U9629 (N_9629,N_7172,N_6447);
or U9630 (N_9630,N_6195,N_7494);
nor U9631 (N_9631,N_6783,N_6731);
and U9632 (N_9632,N_6113,N_6923);
nor U9633 (N_9633,N_7887,N_6565);
nand U9634 (N_9634,N_6068,N_7751);
nor U9635 (N_9635,N_6179,N_7211);
or U9636 (N_9636,N_6458,N_6483);
and U9637 (N_9637,N_7611,N_7139);
or U9638 (N_9638,N_6548,N_6769);
nor U9639 (N_9639,N_7273,N_6928);
and U9640 (N_9640,N_6127,N_7285);
nor U9641 (N_9641,N_6992,N_7134);
nand U9642 (N_9642,N_6275,N_7621);
and U9643 (N_9643,N_6569,N_7477);
and U9644 (N_9644,N_7188,N_6153);
and U9645 (N_9645,N_7895,N_6130);
and U9646 (N_9646,N_6016,N_7681);
or U9647 (N_9647,N_6779,N_6248);
or U9648 (N_9648,N_7873,N_6057);
nor U9649 (N_9649,N_7879,N_6946);
or U9650 (N_9650,N_7218,N_7571);
nand U9651 (N_9651,N_7413,N_6420);
or U9652 (N_9652,N_7028,N_6234);
and U9653 (N_9653,N_7988,N_7770);
and U9654 (N_9654,N_7036,N_6405);
nand U9655 (N_9655,N_7016,N_7937);
nand U9656 (N_9656,N_7935,N_7390);
or U9657 (N_9657,N_7803,N_7870);
and U9658 (N_9658,N_7985,N_7766);
xor U9659 (N_9659,N_7784,N_7748);
nor U9660 (N_9660,N_6554,N_7744);
nor U9661 (N_9661,N_6977,N_7609);
nor U9662 (N_9662,N_6016,N_7419);
xnor U9663 (N_9663,N_7098,N_7716);
and U9664 (N_9664,N_7589,N_6380);
and U9665 (N_9665,N_6946,N_7962);
nor U9666 (N_9666,N_7869,N_6145);
or U9667 (N_9667,N_7390,N_6198);
or U9668 (N_9668,N_6042,N_7415);
and U9669 (N_9669,N_6675,N_7006);
xnor U9670 (N_9670,N_6875,N_6840);
nor U9671 (N_9671,N_6817,N_6393);
or U9672 (N_9672,N_7666,N_6751);
or U9673 (N_9673,N_6233,N_6186);
nand U9674 (N_9674,N_7234,N_6067);
and U9675 (N_9675,N_7336,N_7368);
nand U9676 (N_9676,N_7758,N_6211);
or U9677 (N_9677,N_6623,N_6168);
nor U9678 (N_9678,N_7903,N_6585);
and U9679 (N_9679,N_6640,N_7543);
nor U9680 (N_9680,N_6265,N_6750);
or U9681 (N_9681,N_6623,N_7378);
and U9682 (N_9682,N_7510,N_7670);
nand U9683 (N_9683,N_6016,N_7701);
nand U9684 (N_9684,N_6129,N_6326);
nor U9685 (N_9685,N_7857,N_6238);
and U9686 (N_9686,N_6853,N_7894);
or U9687 (N_9687,N_6701,N_6526);
nand U9688 (N_9688,N_6599,N_7000);
nand U9689 (N_9689,N_6173,N_7818);
and U9690 (N_9690,N_6219,N_6501);
and U9691 (N_9691,N_6801,N_7114);
or U9692 (N_9692,N_7771,N_7237);
nand U9693 (N_9693,N_6458,N_6469);
nor U9694 (N_9694,N_7479,N_6348);
nor U9695 (N_9695,N_6873,N_7997);
and U9696 (N_9696,N_7710,N_7524);
nand U9697 (N_9697,N_6948,N_6062);
and U9698 (N_9698,N_6742,N_7581);
and U9699 (N_9699,N_6517,N_7764);
and U9700 (N_9700,N_6336,N_7643);
nand U9701 (N_9701,N_6705,N_6028);
nor U9702 (N_9702,N_7744,N_7184);
nor U9703 (N_9703,N_6842,N_6136);
or U9704 (N_9704,N_7769,N_6925);
nand U9705 (N_9705,N_7385,N_7538);
and U9706 (N_9706,N_7325,N_6904);
or U9707 (N_9707,N_6499,N_7065);
xor U9708 (N_9708,N_6535,N_7800);
and U9709 (N_9709,N_6000,N_6309);
and U9710 (N_9710,N_6090,N_7959);
and U9711 (N_9711,N_7155,N_7826);
nor U9712 (N_9712,N_7705,N_7080);
or U9713 (N_9713,N_6742,N_6806);
nand U9714 (N_9714,N_7302,N_6197);
nor U9715 (N_9715,N_6593,N_6338);
nor U9716 (N_9716,N_7411,N_6529);
nand U9717 (N_9717,N_7597,N_7491);
xnor U9718 (N_9718,N_6168,N_6435);
or U9719 (N_9719,N_7167,N_7985);
or U9720 (N_9720,N_6008,N_7472);
nand U9721 (N_9721,N_6848,N_6940);
and U9722 (N_9722,N_6172,N_7143);
and U9723 (N_9723,N_7958,N_7138);
nand U9724 (N_9724,N_6392,N_7938);
and U9725 (N_9725,N_6336,N_6479);
nand U9726 (N_9726,N_6435,N_6982);
or U9727 (N_9727,N_7937,N_6163);
nand U9728 (N_9728,N_6463,N_7388);
nor U9729 (N_9729,N_6500,N_7626);
nor U9730 (N_9730,N_6764,N_7776);
nand U9731 (N_9731,N_6389,N_7209);
and U9732 (N_9732,N_6286,N_6442);
nor U9733 (N_9733,N_6452,N_6039);
nor U9734 (N_9734,N_7596,N_6526);
nor U9735 (N_9735,N_6511,N_6284);
or U9736 (N_9736,N_6488,N_7806);
xnor U9737 (N_9737,N_6167,N_7415);
and U9738 (N_9738,N_7974,N_6974);
or U9739 (N_9739,N_6952,N_6619);
or U9740 (N_9740,N_6924,N_6288);
or U9741 (N_9741,N_6165,N_6322);
nor U9742 (N_9742,N_7450,N_6395);
or U9743 (N_9743,N_6532,N_7523);
nand U9744 (N_9744,N_6926,N_7477);
nand U9745 (N_9745,N_7920,N_6548);
and U9746 (N_9746,N_6830,N_6650);
and U9747 (N_9747,N_7831,N_7378);
and U9748 (N_9748,N_6874,N_6555);
or U9749 (N_9749,N_6707,N_6699);
nand U9750 (N_9750,N_7035,N_7105);
or U9751 (N_9751,N_6986,N_6865);
xor U9752 (N_9752,N_6729,N_7273);
nor U9753 (N_9753,N_7722,N_7525);
or U9754 (N_9754,N_7534,N_7981);
nand U9755 (N_9755,N_6113,N_7019);
nor U9756 (N_9756,N_6953,N_6984);
nor U9757 (N_9757,N_7332,N_6669);
nor U9758 (N_9758,N_7956,N_7136);
and U9759 (N_9759,N_6904,N_6567);
and U9760 (N_9760,N_7618,N_7899);
and U9761 (N_9761,N_6299,N_6092);
and U9762 (N_9762,N_7401,N_7339);
and U9763 (N_9763,N_7901,N_6694);
or U9764 (N_9764,N_7317,N_6903);
nor U9765 (N_9765,N_7747,N_6872);
and U9766 (N_9766,N_7270,N_7272);
nor U9767 (N_9767,N_7437,N_6483);
nand U9768 (N_9768,N_7546,N_6017);
xnor U9769 (N_9769,N_7470,N_7775);
nor U9770 (N_9770,N_6973,N_6337);
or U9771 (N_9771,N_6315,N_7253);
or U9772 (N_9772,N_7204,N_7594);
or U9773 (N_9773,N_6764,N_6100);
nand U9774 (N_9774,N_7275,N_6038);
nor U9775 (N_9775,N_7342,N_7311);
and U9776 (N_9776,N_7823,N_6995);
or U9777 (N_9777,N_7894,N_7341);
xor U9778 (N_9778,N_7694,N_6462);
and U9779 (N_9779,N_6128,N_6720);
or U9780 (N_9780,N_7536,N_7401);
nand U9781 (N_9781,N_7967,N_7608);
nand U9782 (N_9782,N_6113,N_6210);
or U9783 (N_9783,N_6605,N_7516);
and U9784 (N_9784,N_7913,N_6082);
and U9785 (N_9785,N_6181,N_7439);
nor U9786 (N_9786,N_6731,N_7491);
nand U9787 (N_9787,N_7364,N_6987);
nand U9788 (N_9788,N_6490,N_6383);
nor U9789 (N_9789,N_6165,N_6053);
and U9790 (N_9790,N_6813,N_6403);
nand U9791 (N_9791,N_7708,N_7903);
or U9792 (N_9792,N_7451,N_6407);
and U9793 (N_9793,N_7577,N_7513);
or U9794 (N_9794,N_7681,N_7761);
and U9795 (N_9795,N_6098,N_6977);
and U9796 (N_9796,N_7171,N_6341);
or U9797 (N_9797,N_6438,N_6729);
xor U9798 (N_9798,N_6783,N_7079);
nor U9799 (N_9799,N_7892,N_6781);
nand U9800 (N_9800,N_6048,N_6813);
xnor U9801 (N_9801,N_6206,N_7336);
or U9802 (N_9802,N_6231,N_6419);
nor U9803 (N_9803,N_6857,N_6167);
nor U9804 (N_9804,N_6813,N_6142);
or U9805 (N_9805,N_7399,N_6942);
nor U9806 (N_9806,N_6973,N_6573);
nor U9807 (N_9807,N_6537,N_6332);
or U9808 (N_9808,N_7504,N_7961);
xnor U9809 (N_9809,N_7918,N_6297);
and U9810 (N_9810,N_7419,N_7971);
nand U9811 (N_9811,N_7825,N_6413);
or U9812 (N_9812,N_6141,N_6062);
nor U9813 (N_9813,N_7949,N_7612);
xnor U9814 (N_9814,N_6895,N_6597);
nor U9815 (N_9815,N_6667,N_6391);
nand U9816 (N_9816,N_7619,N_6749);
nor U9817 (N_9817,N_6468,N_6805);
or U9818 (N_9818,N_6503,N_6386);
or U9819 (N_9819,N_7818,N_6683);
nand U9820 (N_9820,N_6011,N_6105);
nand U9821 (N_9821,N_7962,N_7164);
and U9822 (N_9822,N_6797,N_7916);
or U9823 (N_9823,N_6410,N_6366);
nand U9824 (N_9824,N_7966,N_6994);
or U9825 (N_9825,N_6169,N_6844);
or U9826 (N_9826,N_6832,N_6382);
or U9827 (N_9827,N_6212,N_6635);
nor U9828 (N_9828,N_7062,N_7365);
nor U9829 (N_9829,N_7378,N_6643);
and U9830 (N_9830,N_6280,N_6676);
nand U9831 (N_9831,N_6293,N_7658);
nor U9832 (N_9832,N_6961,N_6640);
nand U9833 (N_9833,N_6658,N_6141);
and U9834 (N_9834,N_6368,N_7757);
xnor U9835 (N_9835,N_6015,N_7249);
and U9836 (N_9836,N_7206,N_7813);
nor U9837 (N_9837,N_7671,N_6094);
and U9838 (N_9838,N_7786,N_7792);
or U9839 (N_9839,N_6500,N_6023);
or U9840 (N_9840,N_7236,N_6346);
and U9841 (N_9841,N_7904,N_7909);
and U9842 (N_9842,N_7237,N_7429);
nand U9843 (N_9843,N_6987,N_6195);
and U9844 (N_9844,N_6305,N_6511);
nor U9845 (N_9845,N_7651,N_7674);
or U9846 (N_9846,N_6709,N_6930);
nor U9847 (N_9847,N_7641,N_6075);
xor U9848 (N_9848,N_6350,N_7471);
or U9849 (N_9849,N_7846,N_7385);
and U9850 (N_9850,N_7844,N_7551);
or U9851 (N_9851,N_7107,N_6860);
nor U9852 (N_9852,N_6479,N_7623);
or U9853 (N_9853,N_7312,N_7282);
nand U9854 (N_9854,N_6595,N_7430);
and U9855 (N_9855,N_7409,N_7286);
and U9856 (N_9856,N_6295,N_7021);
nor U9857 (N_9857,N_7884,N_6302);
and U9858 (N_9858,N_7442,N_7912);
and U9859 (N_9859,N_7328,N_7159);
nand U9860 (N_9860,N_6657,N_6769);
nand U9861 (N_9861,N_7970,N_7301);
and U9862 (N_9862,N_6592,N_6797);
nor U9863 (N_9863,N_7731,N_6827);
or U9864 (N_9864,N_6429,N_7392);
and U9865 (N_9865,N_7540,N_7839);
nor U9866 (N_9866,N_7504,N_6911);
or U9867 (N_9867,N_6235,N_6763);
and U9868 (N_9868,N_7027,N_6164);
nor U9869 (N_9869,N_6786,N_6964);
xor U9870 (N_9870,N_6859,N_6469);
nor U9871 (N_9871,N_7094,N_6588);
or U9872 (N_9872,N_7946,N_7380);
nor U9873 (N_9873,N_6674,N_6235);
nor U9874 (N_9874,N_6696,N_6881);
nand U9875 (N_9875,N_7963,N_6942);
nand U9876 (N_9876,N_7972,N_6419);
nand U9877 (N_9877,N_7639,N_6892);
nor U9878 (N_9878,N_6945,N_6174);
or U9879 (N_9879,N_7289,N_6130);
nor U9880 (N_9880,N_7746,N_6402);
or U9881 (N_9881,N_6531,N_6392);
nand U9882 (N_9882,N_6260,N_7708);
or U9883 (N_9883,N_7613,N_6886);
nor U9884 (N_9884,N_7130,N_7863);
nor U9885 (N_9885,N_7398,N_6865);
and U9886 (N_9886,N_7381,N_6089);
and U9887 (N_9887,N_6860,N_6786);
and U9888 (N_9888,N_6799,N_6896);
or U9889 (N_9889,N_6664,N_6428);
nand U9890 (N_9890,N_6160,N_7397);
and U9891 (N_9891,N_6972,N_6461);
and U9892 (N_9892,N_6006,N_6493);
xor U9893 (N_9893,N_7510,N_6397);
nand U9894 (N_9894,N_7097,N_6187);
nor U9895 (N_9895,N_6679,N_6507);
and U9896 (N_9896,N_7853,N_7003);
nand U9897 (N_9897,N_6435,N_7746);
or U9898 (N_9898,N_7717,N_7287);
nor U9899 (N_9899,N_7526,N_7322);
or U9900 (N_9900,N_6030,N_7024);
nand U9901 (N_9901,N_6121,N_6643);
or U9902 (N_9902,N_6357,N_6099);
and U9903 (N_9903,N_7290,N_7636);
nor U9904 (N_9904,N_7852,N_6016);
nor U9905 (N_9905,N_7489,N_7000);
nor U9906 (N_9906,N_7607,N_7478);
nor U9907 (N_9907,N_7384,N_7984);
and U9908 (N_9908,N_7442,N_7979);
or U9909 (N_9909,N_7785,N_6976);
or U9910 (N_9910,N_6238,N_6868);
nand U9911 (N_9911,N_7097,N_6376);
nand U9912 (N_9912,N_7445,N_6660);
or U9913 (N_9913,N_7986,N_7651);
or U9914 (N_9914,N_6942,N_6956);
and U9915 (N_9915,N_6590,N_6865);
nor U9916 (N_9916,N_6931,N_7441);
and U9917 (N_9917,N_6898,N_6625);
and U9918 (N_9918,N_6329,N_7869);
nand U9919 (N_9919,N_7057,N_6179);
nand U9920 (N_9920,N_6949,N_7830);
or U9921 (N_9921,N_6486,N_7887);
nand U9922 (N_9922,N_7111,N_6018);
nand U9923 (N_9923,N_7516,N_7403);
or U9924 (N_9924,N_7954,N_7421);
nor U9925 (N_9925,N_6761,N_6399);
and U9926 (N_9926,N_6687,N_6578);
nor U9927 (N_9927,N_6025,N_6805);
nor U9928 (N_9928,N_7621,N_6699);
nand U9929 (N_9929,N_7673,N_7967);
and U9930 (N_9930,N_6654,N_7126);
or U9931 (N_9931,N_6390,N_7659);
and U9932 (N_9932,N_6160,N_7425);
nor U9933 (N_9933,N_6541,N_6253);
or U9934 (N_9934,N_7205,N_6185);
and U9935 (N_9935,N_6020,N_7572);
or U9936 (N_9936,N_6306,N_7154);
nand U9937 (N_9937,N_7174,N_6566);
xnor U9938 (N_9938,N_7306,N_7778);
or U9939 (N_9939,N_6909,N_6715);
or U9940 (N_9940,N_6129,N_7707);
and U9941 (N_9941,N_6550,N_6618);
or U9942 (N_9942,N_7301,N_7527);
nand U9943 (N_9943,N_7848,N_6153);
nor U9944 (N_9944,N_6076,N_7002);
nand U9945 (N_9945,N_7407,N_7620);
nand U9946 (N_9946,N_6794,N_7757);
or U9947 (N_9947,N_7025,N_7681);
nor U9948 (N_9948,N_7366,N_6468);
nor U9949 (N_9949,N_7293,N_6810);
and U9950 (N_9950,N_6291,N_7147);
and U9951 (N_9951,N_7363,N_6058);
nor U9952 (N_9952,N_7404,N_6105);
nor U9953 (N_9953,N_6878,N_6038);
nor U9954 (N_9954,N_6083,N_7088);
nand U9955 (N_9955,N_7982,N_6197);
nand U9956 (N_9956,N_7742,N_6902);
nor U9957 (N_9957,N_6065,N_7874);
and U9958 (N_9958,N_7801,N_7177);
and U9959 (N_9959,N_6129,N_7559);
or U9960 (N_9960,N_6673,N_6892);
or U9961 (N_9961,N_7955,N_7414);
nor U9962 (N_9962,N_7924,N_7279);
or U9963 (N_9963,N_7543,N_7132);
xnor U9964 (N_9964,N_6475,N_7124);
or U9965 (N_9965,N_7143,N_6670);
nand U9966 (N_9966,N_6593,N_7738);
and U9967 (N_9967,N_7207,N_6450);
or U9968 (N_9968,N_6869,N_7012);
nand U9969 (N_9969,N_6355,N_6192);
xnor U9970 (N_9970,N_7818,N_6120);
or U9971 (N_9971,N_7035,N_6892);
or U9972 (N_9972,N_7323,N_6188);
nand U9973 (N_9973,N_7416,N_6861);
nand U9974 (N_9974,N_6130,N_7462);
nand U9975 (N_9975,N_7299,N_6441);
or U9976 (N_9976,N_7526,N_6109);
nor U9977 (N_9977,N_7728,N_6727);
nor U9978 (N_9978,N_7328,N_7721);
or U9979 (N_9979,N_7825,N_6367);
or U9980 (N_9980,N_6978,N_7862);
and U9981 (N_9981,N_6179,N_6694);
nor U9982 (N_9982,N_7267,N_7812);
or U9983 (N_9983,N_6632,N_7017);
or U9984 (N_9984,N_6203,N_6515);
nand U9985 (N_9985,N_7469,N_6528);
or U9986 (N_9986,N_7904,N_6357);
or U9987 (N_9987,N_7948,N_6010);
or U9988 (N_9988,N_7609,N_7095);
or U9989 (N_9989,N_7145,N_6743);
or U9990 (N_9990,N_7963,N_7596);
or U9991 (N_9991,N_7008,N_6451);
or U9992 (N_9992,N_7322,N_7602);
nor U9993 (N_9993,N_7262,N_6977);
nand U9994 (N_9994,N_6600,N_6407);
nand U9995 (N_9995,N_6502,N_7650);
nand U9996 (N_9996,N_6387,N_7251);
nor U9997 (N_9997,N_6298,N_6660);
and U9998 (N_9998,N_6795,N_6305);
or U9999 (N_9999,N_7124,N_6220);
nor UO_0 (O_0,N_9994,N_8420);
xor UO_1 (O_1,N_9563,N_9643);
nand UO_2 (O_2,N_9763,N_9996);
and UO_3 (O_3,N_8092,N_8142);
and UO_4 (O_4,N_9377,N_8994);
nor UO_5 (O_5,N_9389,N_9308);
nor UO_6 (O_6,N_8862,N_8450);
nand UO_7 (O_7,N_8835,N_8687);
nand UO_8 (O_8,N_8488,N_9885);
and UO_9 (O_9,N_9372,N_8303);
nand UO_10 (O_10,N_9082,N_8341);
nor UO_11 (O_11,N_8894,N_8383);
and UO_12 (O_12,N_9892,N_8164);
or UO_13 (O_13,N_9819,N_8436);
nor UO_14 (O_14,N_8710,N_8745);
nand UO_15 (O_15,N_9070,N_8019);
or UO_16 (O_16,N_8509,N_8136);
or UO_17 (O_17,N_8767,N_8929);
xor UO_18 (O_18,N_8864,N_9453);
nor UO_19 (O_19,N_9973,N_9380);
nand UO_20 (O_20,N_9486,N_9790);
or UO_21 (O_21,N_9426,N_8001);
and UO_22 (O_22,N_8721,N_8099);
and UO_23 (O_23,N_8524,N_8597);
nor UO_24 (O_24,N_9371,N_8080);
and UO_25 (O_25,N_8014,N_8065);
nor UO_26 (O_26,N_8210,N_8596);
nor UO_27 (O_27,N_9013,N_8343);
nand UO_28 (O_28,N_9495,N_9835);
nand UO_29 (O_29,N_8367,N_8669);
nand UO_30 (O_30,N_8474,N_9206);
nand UO_31 (O_31,N_9855,N_8585);
nor UO_32 (O_32,N_9154,N_8733);
nand UO_33 (O_33,N_8174,N_9174);
and UO_34 (O_34,N_9960,N_8555);
nand UO_35 (O_35,N_8643,N_8476);
or UO_36 (O_36,N_8677,N_9759);
or UO_37 (O_37,N_9703,N_9040);
or UO_38 (O_38,N_9633,N_9877);
and UO_39 (O_39,N_9535,N_8969);
or UO_40 (O_40,N_9564,N_8196);
and UO_41 (O_41,N_9198,N_8141);
or UO_42 (O_42,N_8814,N_8253);
and UO_43 (O_43,N_8340,N_8122);
and UO_44 (O_44,N_8078,N_9700);
nor UO_45 (O_45,N_9044,N_9692);
or UO_46 (O_46,N_8858,N_9567);
nand UO_47 (O_47,N_9727,N_9108);
nor UO_48 (O_48,N_8836,N_9625);
and UO_49 (O_49,N_8696,N_9736);
nand UO_50 (O_50,N_9497,N_9755);
nor UO_51 (O_51,N_8030,N_9830);
or UO_52 (O_52,N_9420,N_9899);
nand UO_53 (O_53,N_8096,N_9777);
nor UO_54 (O_54,N_9851,N_8849);
or UO_55 (O_55,N_9459,N_8888);
nor UO_56 (O_56,N_8149,N_9365);
nor UO_57 (O_57,N_8156,N_9800);
nor UO_58 (O_58,N_9775,N_9391);
nand UO_59 (O_59,N_9615,N_8647);
or UO_60 (O_60,N_8651,N_9510);
and UO_61 (O_61,N_9518,N_8565);
nand UO_62 (O_62,N_8130,N_9549);
nand UO_63 (O_63,N_8955,N_9509);
or UO_64 (O_64,N_8923,N_9618);
nor UO_65 (O_65,N_8649,N_9020);
nand UO_66 (O_66,N_9418,N_9005);
nor UO_67 (O_67,N_9017,N_9092);
or UO_68 (O_68,N_8103,N_8478);
nand UO_69 (O_69,N_8886,N_8339);
or UO_70 (O_70,N_9268,N_9061);
nand UO_71 (O_71,N_8757,N_8514);
and UO_72 (O_72,N_8935,N_8055);
and UO_73 (O_73,N_8244,N_8069);
and UO_74 (O_74,N_9592,N_8828);
and UO_75 (O_75,N_9989,N_8451);
nand UO_76 (O_76,N_9544,N_9281);
nor UO_77 (O_77,N_9728,N_9995);
or UO_78 (O_78,N_9100,N_9347);
nand UO_79 (O_79,N_9300,N_8521);
nand UO_80 (O_80,N_8952,N_9744);
nand UO_81 (O_81,N_9332,N_8200);
and UO_82 (O_82,N_8638,N_8542);
or UO_83 (O_83,N_9758,N_8553);
nor UO_84 (O_84,N_9208,N_9649);
and UO_85 (O_85,N_9911,N_8538);
nor UO_86 (O_86,N_9712,N_8440);
nand UO_87 (O_87,N_9571,N_8694);
xnor UO_88 (O_88,N_9203,N_8586);
nor UO_89 (O_89,N_8667,N_9757);
nand UO_90 (O_90,N_8225,N_8079);
and UO_91 (O_91,N_9555,N_9417);
or UO_92 (O_92,N_8199,N_8104);
and UO_93 (O_93,N_9504,N_8355);
or UO_94 (O_94,N_8872,N_9796);
nor UO_95 (O_95,N_8530,N_9328);
and UO_96 (O_96,N_9167,N_9578);
or UO_97 (O_97,N_9138,N_8140);
or UO_98 (O_98,N_9536,N_9547);
nor UO_99 (O_99,N_8531,N_8921);
and UO_100 (O_100,N_8959,N_8874);
or UO_101 (O_101,N_8985,N_8443);
nor UO_102 (O_102,N_8599,N_8422);
or UO_103 (O_103,N_9752,N_9980);
nor UO_104 (O_104,N_8656,N_9805);
or UO_105 (O_105,N_8241,N_9500);
nor UO_106 (O_106,N_9290,N_9277);
nor UO_107 (O_107,N_8240,N_8685);
or UO_108 (O_108,N_9694,N_8077);
or UO_109 (O_109,N_9140,N_8941);
or UO_110 (O_110,N_8447,N_8363);
nand UO_111 (O_111,N_8012,N_9530);
and UO_112 (O_112,N_9697,N_8485);
nor UO_113 (O_113,N_8909,N_9818);
and UO_114 (O_114,N_8526,N_8356);
or UO_115 (O_115,N_8507,N_8646);
nor UO_116 (O_116,N_8829,N_8912);
or UO_117 (O_117,N_9968,N_9238);
and UO_118 (O_118,N_9784,N_9189);
or UO_119 (O_119,N_8574,N_8071);
nand UO_120 (O_120,N_8106,N_8911);
nor UO_121 (O_121,N_8152,N_9452);
nor UO_122 (O_122,N_8382,N_8287);
nand UO_123 (O_123,N_8897,N_8505);
nor UO_124 (O_124,N_9127,N_8237);
nor UO_125 (O_125,N_9858,N_8998);
and UO_126 (O_126,N_8026,N_9442);
nor UO_127 (O_127,N_8029,N_9230);
and UO_128 (O_128,N_9396,N_9056);
and UO_129 (O_129,N_8310,N_8841);
or UO_130 (O_130,N_9713,N_8431);
nand UO_131 (O_131,N_8228,N_8748);
and UO_132 (O_132,N_8725,N_8401);
or UO_133 (O_133,N_9693,N_8458);
and UO_134 (O_134,N_8933,N_8259);
or UO_135 (O_135,N_8127,N_9927);
nand UO_136 (O_136,N_8492,N_9445);
nand UO_137 (O_137,N_8540,N_9836);
and UO_138 (O_138,N_9646,N_8977);
nand UO_139 (O_139,N_9856,N_9373);
or UO_140 (O_140,N_9579,N_9887);
nand UO_141 (O_141,N_9981,N_8881);
and UO_142 (O_142,N_9089,N_8290);
or UO_143 (O_143,N_8100,N_9684);
and UO_144 (O_144,N_9745,N_8593);
nand UO_145 (O_145,N_8523,N_9209);
nor UO_146 (O_146,N_9833,N_8203);
and UO_147 (O_147,N_8020,N_9264);
nand UO_148 (O_148,N_9000,N_9589);
nand UO_149 (O_149,N_8332,N_9998);
and UO_150 (O_150,N_8190,N_9113);
and UO_151 (O_151,N_8416,N_9216);
nor UO_152 (O_152,N_9423,N_9030);
or UO_153 (O_153,N_8711,N_8282);
and UO_154 (O_154,N_8758,N_8094);
or UO_155 (O_155,N_9948,N_9025);
nor UO_156 (O_156,N_9144,N_9593);
nor UO_157 (O_157,N_9999,N_8000);
nand UO_158 (O_158,N_8257,N_9492);
nand UO_159 (O_159,N_9468,N_8954);
nand UO_160 (O_160,N_9952,N_9135);
and UO_161 (O_161,N_8723,N_9997);
nor UO_162 (O_162,N_8482,N_8668);
nand UO_163 (O_163,N_9457,N_9085);
nor UO_164 (O_164,N_8256,N_9880);
and UO_165 (O_165,N_9881,N_8306);
nand UO_166 (O_166,N_9449,N_8729);
and UO_167 (O_167,N_9982,N_8213);
and UO_168 (O_168,N_8805,N_9515);
and UO_169 (O_169,N_8792,N_9165);
or UO_170 (O_170,N_9185,N_8085);
xor UO_171 (O_171,N_9307,N_9447);
and UO_172 (O_172,N_8622,N_9966);
or UO_173 (O_173,N_9145,N_9782);
nand UO_174 (O_174,N_8176,N_9047);
nand UO_175 (O_175,N_9793,N_8610);
and UO_176 (O_176,N_8800,N_9699);
and UO_177 (O_177,N_8993,N_8129);
xor UO_178 (O_178,N_9111,N_8479);
nor UO_179 (O_179,N_8279,N_8231);
or UO_180 (O_180,N_9481,N_9679);
or UO_181 (O_181,N_9430,N_9730);
nand UO_182 (O_182,N_9237,N_9034);
or UO_183 (O_183,N_8703,N_9944);
nor UO_184 (O_184,N_8762,N_9936);
or UO_185 (O_185,N_8188,N_8430);
nand UO_186 (O_186,N_9031,N_8301);
nand UO_187 (O_187,N_9916,N_8915);
and UO_188 (O_188,N_9067,N_8317);
or UO_189 (O_189,N_8081,N_9037);
nor UO_190 (O_190,N_8371,N_9149);
nor UO_191 (O_191,N_8624,N_9156);
nand UO_192 (O_192,N_9732,N_9598);
or UO_193 (O_193,N_8330,N_9639);
nor UO_194 (O_194,N_9946,N_8611);
or UO_195 (O_195,N_8751,N_9751);
or UO_196 (O_196,N_8868,N_9245);
and UO_197 (O_197,N_9942,N_8720);
or UO_198 (O_198,N_8676,N_8054);
and UO_199 (O_199,N_8865,N_8808);
nand UO_200 (O_200,N_8090,N_8381);
or UO_201 (O_201,N_8486,N_9807);
or UO_202 (O_202,N_9719,N_9408);
or UO_203 (O_203,N_8937,N_8544);
nand UO_204 (O_204,N_8847,N_9940);
nor UO_205 (O_205,N_8175,N_9152);
and UO_206 (O_206,N_9403,N_8033);
nand UO_207 (O_207,N_8121,N_8691);
nor UO_208 (O_208,N_8499,N_9514);
nand UO_209 (O_209,N_9496,N_9436);
nor UO_210 (O_210,N_8158,N_9770);
nor UO_211 (O_211,N_9412,N_9619);
or UO_212 (O_212,N_9319,N_8101);
nand UO_213 (O_213,N_9783,N_9358);
or UO_214 (O_214,N_9705,N_8641);
and UO_215 (O_215,N_9912,N_9124);
or UO_216 (O_216,N_8334,N_8600);
nor UO_217 (O_217,N_9863,N_8853);
nand UO_218 (O_218,N_9055,N_8229);
and UO_219 (O_219,N_8892,N_8148);
and UO_220 (O_220,N_9658,N_8927);
or UO_221 (O_221,N_9121,N_9614);
or UO_222 (O_222,N_8144,N_8324);
nor UO_223 (O_223,N_9428,N_9769);
and UO_224 (O_224,N_9572,N_9594);
or UO_225 (O_225,N_9018,N_9345);
and UO_226 (O_226,N_9621,N_8556);
nor UO_227 (O_227,N_9126,N_8885);
nand UO_228 (O_228,N_8021,N_8365);
nor UO_229 (O_229,N_8198,N_9406);
or UO_230 (O_230,N_8126,N_8770);
or UO_231 (O_231,N_9803,N_9181);
or UO_232 (O_232,N_8945,N_9150);
or UO_233 (O_233,N_8672,N_8801);
or UO_234 (O_234,N_9582,N_8250);
or UO_235 (O_235,N_8347,N_9976);
or UO_236 (O_236,N_8645,N_9943);
nand UO_237 (O_237,N_8326,N_8208);
or UO_238 (O_238,N_8863,N_9218);
nor UO_239 (O_239,N_9467,N_8372);
nor UO_240 (O_240,N_9708,N_9580);
or UO_241 (O_241,N_8702,N_9917);
or UO_242 (O_242,N_8248,N_9227);
and UO_243 (O_243,N_8296,N_9071);
nor UO_244 (O_244,N_8617,N_9099);
xnor UO_245 (O_245,N_8695,N_9626);
or UO_246 (O_246,N_8370,N_9463);
and UO_247 (O_247,N_8235,N_9460);
or UO_248 (O_248,N_9969,N_9860);
nor UO_249 (O_249,N_8761,N_8234);
nor UO_250 (O_250,N_8582,N_9725);
and UO_251 (O_251,N_8781,N_8648);
nand UO_252 (O_252,N_9933,N_9513);
xor UO_253 (O_253,N_8150,N_9301);
nand UO_254 (O_254,N_8034,N_9664);
or UO_255 (O_255,N_8666,N_9006);
or UO_256 (O_256,N_9740,N_9250);
nand UO_257 (O_257,N_9850,N_8878);
and UO_258 (O_258,N_9147,N_8266);
or UO_259 (O_259,N_8067,N_9584);
nand UO_260 (O_260,N_8780,N_9213);
nand UO_261 (O_261,N_8169,N_9722);
nand UO_262 (O_262,N_9098,N_8918);
nand UO_263 (O_263,N_9284,N_8448);
nand UO_264 (O_264,N_8336,N_9359);
and UO_265 (O_265,N_8528,N_9327);
nand UO_266 (O_266,N_9975,N_8895);
or UO_267 (O_267,N_8851,N_8245);
and UO_268 (O_268,N_9087,N_8764);
and UO_269 (O_269,N_9704,N_9489);
nand UO_270 (O_270,N_9680,N_9634);
nand UO_271 (O_271,N_8454,N_8453);
and UO_272 (O_272,N_8378,N_8261);
or UO_273 (O_273,N_9988,N_8024);
nor UO_274 (O_274,N_9962,N_9004);
nor UO_275 (O_275,N_8418,N_8061);
and UO_276 (O_276,N_9168,N_9438);
or UO_277 (O_277,N_8982,N_8637);
nor UO_278 (O_278,N_8202,N_9552);
nor UO_279 (O_279,N_9945,N_8232);
nor UO_280 (O_280,N_8389,N_8840);
or UO_281 (O_281,N_9874,N_9632);
or UO_282 (O_282,N_8525,N_9691);
and UO_283 (O_283,N_9723,N_9026);
nand UO_284 (O_284,N_8491,N_9240);
or UO_285 (O_285,N_8821,N_9529);
and UO_286 (O_286,N_9627,N_9687);
nand UO_287 (O_287,N_8084,N_8284);
xor UO_288 (O_288,N_8551,N_8115);
nand UO_289 (O_289,N_9059,N_8006);
and UO_290 (O_290,N_9690,N_9231);
nor UO_291 (O_291,N_8449,N_9654);
nor UO_292 (O_292,N_9748,N_9681);
or UO_293 (O_293,N_9970,N_8763);
xor UO_294 (O_294,N_8335,N_9622);
nor UO_295 (O_295,N_9788,N_9974);
or UO_296 (O_296,N_8446,N_9461);
or UO_297 (O_297,N_9348,N_9586);
or UO_298 (O_298,N_9370,N_8437);
or UO_299 (O_299,N_9729,N_9407);
nor UO_300 (O_300,N_9817,N_8297);
nor UO_301 (O_301,N_9665,N_9562);
xnor UO_302 (O_302,N_9631,N_8965);
and UO_303 (O_303,N_9717,N_9379);
or UO_304 (O_304,N_8706,N_9585);
and UO_305 (O_305,N_8193,N_8182);
nand UO_306 (O_306,N_8162,N_8359);
and UO_307 (O_307,N_8390,N_9754);
and UO_308 (O_308,N_8050,N_8419);
or UO_309 (O_309,N_9484,N_8896);
or UO_310 (O_310,N_8777,N_8036);
and UO_311 (O_311,N_8796,N_9282);
nor UO_312 (O_312,N_9058,N_8423);
nor UO_313 (O_313,N_8620,N_9908);
nand UO_314 (O_314,N_8086,N_9792);
nand UO_315 (O_315,N_9199,N_8861);
and UO_316 (O_316,N_8690,N_9338);
nand UO_317 (O_317,N_9223,N_9279);
or UO_318 (O_318,N_9958,N_8361);
or UO_319 (O_319,N_9870,N_9425);
nor UO_320 (O_320,N_9068,N_9656);
xor UO_321 (O_321,N_9638,N_9322);
or UO_322 (O_322,N_9252,N_9450);
nor UO_323 (O_323,N_9288,N_9630);
and UO_324 (O_324,N_8260,N_8673);
and UO_325 (O_325,N_9283,N_8817);
and UO_326 (O_326,N_8124,N_9304);
nor UO_327 (O_327,N_8072,N_9939);
xor UO_328 (O_328,N_9129,N_9077);
nand UO_329 (O_329,N_9239,N_9711);
and UO_330 (O_330,N_9392,N_8117);
nor UO_331 (O_331,N_9689,N_8961);
nand UO_332 (O_332,N_9191,N_9900);
nor UO_333 (O_333,N_8346,N_9846);
nor UO_334 (O_334,N_8910,N_8215);
or UO_335 (O_335,N_9767,N_8212);
and UO_336 (O_336,N_8899,N_8833);
nand UO_337 (O_337,N_8960,N_9873);
and UO_338 (O_338,N_8110,N_9494);
nand UO_339 (O_339,N_8754,N_8409);
and UO_340 (O_340,N_8223,N_8516);
and UO_341 (O_341,N_8769,N_9977);
nor UO_342 (O_342,N_9965,N_9286);
or UO_343 (O_343,N_9172,N_8964);
and UO_344 (O_344,N_9201,N_8151);
nor UO_345 (O_345,N_8995,N_9232);
and UO_346 (O_346,N_9123,N_8013);
or UO_347 (O_347,N_8661,N_8172);
and UO_348 (O_348,N_8983,N_8327);
nor UO_349 (O_349,N_9561,N_8549);
or UO_350 (O_350,N_8047,N_9568);
or UO_351 (O_351,N_8380,N_9390);
nor UO_352 (O_352,N_8893,N_8404);
or UO_353 (O_353,N_8716,N_8291);
and UO_354 (O_354,N_9932,N_9531);
or UO_355 (O_355,N_9636,N_9062);
or UO_356 (O_356,N_9118,N_9961);
nand UO_357 (O_357,N_9289,N_8902);
and UO_358 (O_358,N_9048,N_8709);
nor UO_359 (O_359,N_9242,N_9101);
nand UO_360 (O_360,N_9413,N_9224);
nand UO_361 (O_361,N_8119,N_8795);
or UO_362 (O_362,N_9901,N_8988);
nand UO_363 (O_363,N_9909,N_9720);
and UO_364 (O_364,N_9204,N_9612);
nand UO_365 (O_365,N_8719,N_9707);
nor UO_366 (O_366,N_9688,N_9212);
or UO_367 (O_367,N_9117,N_8602);
or UO_368 (O_368,N_9387,N_8268);
nor UO_369 (O_369,N_9173,N_8300);
nand UO_370 (O_370,N_8932,N_9344);
xor UO_371 (O_371,N_8262,N_8743);
nand UO_372 (O_372,N_8642,N_8045);
nand UO_373 (O_373,N_8475,N_9251);
nand UO_374 (O_374,N_8870,N_9075);
nand UO_375 (O_375,N_9355,N_9762);
nor UO_376 (O_376,N_9110,N_9641);
or UO_377 (O_377,N_8975,N_8537);
nor UO_378 (O_378,N_9749,N_9141);
and UO_379 (O_379,N_8305,N_9724);
nand UO_380 (O_380,N_8322,N_8541);
and UO_381 (O_381,N_8576,N_9941);
nor UO_382 (O_382,N_8277,N_8527);
nor UO_383 (O_383,N_9565,N_8774);
or UO_384 (O_384,N_8570,N_8128);
or UO_385 (O_385,N_9434,N_9336);
nor UO_386 (O_386,N_8986,N_9405);
or UO_387 (O_387,N_9035,N_9928);
nor UO_388 (O_388,N_8846,N_9669);
and UO_389 (O_389,N_9158,N_8292);
and UO_390 (O_390,N_8396,N_9001);
nand UO_391 (O_391,N_8548,N_9214);
and UO_392 (O_392,N_9195,N_8068);
or UO_393 (O_393,N_8819,N_9811);
and UO_394 (O_394,N_8967,N_9306);
and UO_395 (O_395,N_8934,N_8472);
and UO_396 (O_396,N_8506,N_9263);
or UO_397 (O_397,N_8759,N_9255);
or UO_398 (O_398,N_8276,N_8035);
nor UO_399 (O_399,N_8740,N_8686);
or UO_400 (O_400,N_9764,N_9808);
nand UO_401 (O_401,N_8073,N_9768);
nor UO_402 (O_402,N_8640,N_8884);
or UO_403 (O_403,N_9647,N_9871);
and UO_404 (O_404,N_8270,N_9169);
nor UO_405 (O_405,N_8907,N_8023);
nor UO_406 (O_406,N_8603,N_8496);
and UO_407 (O_407,N_9441,N_8704);
nor UO_408 (O_408,N_9221,N_8319);
nand UO_409 (O_409,N_8015,N_9454);
nand UO_410 (O_410,N_9959,N_9291);
or UO_411 (O_411,N_8621,N_8220);
nand UO_412 (O_412,N_9175,N_9820);
or UO_413 (O_413,N_9029,N_9628);
nand UO_414 (O_414,N_8105,N_9521);
nand UO_415 (O_415,N_8939,N_9051);
and UO_416 (O_416,N_9303,N_8468);
nand UO_417 (O_417,N_9350,N_9604);
or UO_418 (O_418,N_8924,N_9011);
xnor UO_419 (O_419,N_8804,N_8314);
nor UO_420 (O_420,N_8304,N_9993);
nor UO_421 (O_421,N_9057,N_8098);
or UO_422 (O_422,N_9566,N_8568);
nand UO_423 (O_423,N_8946,N_9046);
or UO_424 (O_424,N_8739,N_9802);
nor UO_425 (O_425,N_9439,N_8456);
nand UO_426 (O_426,N_9043,N_8867);
or UO_427 (O_427,N_9456,N_8414);
nor UO_428 (O_428,N_9597,N_8753);
or UO_429 (O_429,N_9534,N_9922);
nor UO_430 (O_430,N_9161,N_9073);
nand UO_431 (O_431,N_8387,N_8815);
and UO_432 (O_432,N_9527,N_9196);
xnor UO_433 (O_433,N_9414,N_9272);
or UO_434 (O_434,N_8772,N_9148);
nor UO_435 (O_435,N_8187,N_8353);
xor UO_436 (O_436,N_8628,N_8908);
and UO_437 (O_437,N_9891,N_9543);
and UO_438 (O_438,N_9421,N_8170);
and UO_439 (O_439,N_8980,N_9466);
nand UO_440 (O_440,N_8424,N_8498);
nor UO_441 (O_441,N_8991,N_8818);
or UO_442 (O_442,N_9812,N_9889);
nor UO_443 (O_443,N_8922,N_8145);
nor UO_444 (O_444,N_8614,N_9813);
nor UO_445 (O_445,N_9587,N_9155);
nor UO_446 (O_446,N_9794,N_9483);
nor UO_447 (O_447,N_8254,N_9064);
nand UO_448 (O_448,N_9557,N_8584);
nor UO_449 (O_449,N_9366,N_9674);
nor UO_450 (O_450,N_8374,N_8675);
nor UO_451 (O_451,N_8062,N_9926);
nor UO_452 (O_452,N_9311,N_8415);
and UO_453 (O_453,N_8670,N_8109);
and UO_454 (O_454,N_8052,N_8368);
xnor UO_455 (O_455,N_9078,N_8615);
or UO_456 (O_456,N_8500,N_8825);
or UO_457 (O_457,N_8629,N_9278);
nor UO_458 (O_458,N_8504,N_9330);
nor UO_459 (O_459,N_9197,N_9596);
or UO_460 (O_460,N_8632,N_9894);
or UO_461 (O_461,N_8749,N_8143);
and UO_462 (O_462,N_9829,N_8512);
nor UO_463 (O_463,N_8807,N_8812);
and UO_464 (O_464,N_9109,N_9316);
and UO_465 (O_465,N_9930,N_8567);
xor UO_466 (O_466,N_8421,N_9847);
nor UO_467 (O_467,N_9655,N_9581);
and UO_468 (O_468,N_9134,N_9088);
nor UO_469 (O_469,N_8776,N_9798);
nand UO_470 (O_470,N_8683,N_9244);
or UO_471 (O_471,N_9991,N_9353);
nand UO_472 (O_472,N_9498,N_8583);
and UO_473 (O_473,N_9600,N_8604);
nor UO_474 (O_474,N_8274,N_8138);
nand UO_475 (O_475,N_9919,N_8756);
and UO_476 (O_476,N_8331,N_9538);
and UO_477 (O_477,N_8022,N_9507);
xnor UO_478 (O_478,N_8226,N_8219);
nor UO_479 (O_479,N_9560,N_9735);
nor UO_480 (O_480,N_9367,N_9617);
or UO_481 (O_481,N_8592,N_8883);
and UO_482 (O_482,N_8222,N_9816);
nand UO_483 (O_483,N_8956,N_9393);
and UO_484 (O_484,N_9743,N_9222);
and UO_485 (O_485,N_8605,N_9551);
and UO_486 (O_486,N_9346,N_8650);
nor UO_487 (O_487,N_8075,N_9937);
and UO_488 (O_488,N_9002,N_8309);
or UO_489 (O_489,N_9292,N_8411);
or UO_490 (O_490,N_9682,N_9676);
or UO_491 (O_491,N_8207,N_9128);
nor UO_492 (O_492,N_8837,N_8184);
nor UO_493 (O_493,N_9478,N_9956);
nor UO_494 (O_494,N_9947,N_8247);
nor UO_495 (O_495,N_9045,N_9095);
nand UO_496 (O_496,N_9652,N_8700);
nor UO_497 (O_497,N_8613,N_9177);
nand UO_498 (O_498,N_8216,N_8786);
nor UO_499 (O_499,N_9384,N_9731);
or UO_500 (O_500,N_9119,N_9361);
or UO_501 (O_501,N_9388,N_9234);
nand UO_502 (O_502,N_8060,N_8242);
and UO_503 (O_503,N_9235,N_9716);
or UO_504 (O_504,N_9821,N_8120);
or UO_505 (O_505,N_8375,N_9363);
nor UO_506 (O_506,N_8787,N_8255);
nand UO_507 (O_507,N_9200,N_9202);
and UO_508 (O_508,N_8606,N_9060);
nand UO_509 (O_509,N_9666,N_9341);
or UO_510 (O_510,N_8183,N_8779);
and UO_511 (O_511,N_8679,N_8480);
nand UO_512 (O_512,N_8027,N_9801);
and UO_513 (O_513,N_8272,N_8007);
nor UO_514 (O_514,N_9603,N_9667);
and UO_515 (O_515,N_9102,N_8822);
and UO_516 (O_516,N_8070,N_9971);
and UO_517 (O_517,N_9799,N_9153);
or UO_518 (O_518,N_8470,N_9166);
xnor UO_519 (O_519,N_8827,N_8325);
nand UO_520 (O_520,N_8264,N_9399);
nor UO_521 (O_521,N_8206,N_9033);
nor UO_522 (O_522,N_8728,N_8236);
or UO_523 (O_523,N_9081,N_8963);
nor UO_524 (O_524,N_8429,N_8118);
or UO_525 (O_525,N_9010,N_9957);
or UO_526 (O_526,N_9331,N_9826);
or UO_527 (O_527,N_9410,N_9843);
or UO_528 (O_528,N_9182,N_8803);
or UO_529 (O_529,N_9038,N_8705);
nand UO_530 (O_530,N_9827,N_9210);
nor UO_531 (O_531,N_8376,N_8379);
nand UO_532 (O_532,N_8366,N_9789);
or UO_533 (O_533,N_8968,N_9476);
nor UO_534 (O_534,N_9787,N_9493);
nor UO_535 (O_535,N_9375,N_9257);
nand UO_536 (O_536,N_8636,N_9575);
or UO_537 (O_537,N_8928,N_8191);
or UO_538 (O_538,N_8298,N_9186);
and UO_539 (O_539,N_9660,N_8323);
or UO_540 (O_540,N_9511,N_8752);
or UO_541 (O_541,N_8947,N_9296);
nor UO_542 (O_542,N_8407,N_8095);
nor UO_543 (O_543,N_8385,N_9395);
nand UO_544 (O_544,N_8996,N_9670);
and UO_545 (O_545,N_9437,N_9313);
nor UO_546 (O_546,N_9502,N_8302);
or UO_547 (O_547,N_8205,N_9648);
or UO_548 (O_548,N_8587,N_9400);
or UO_549 (O_549,N_8898,N_8736);
or UO_550 (O_550,N_9685,N_8778);
and UO_551 (O_551,N_8469,N_8249);
or UO_552 (O_552,N_8852,N_8635);
nor UO_553 (O_553,N_9394,N_8395);
or UO_554 (O_554,N_8623,N_8563);
and UO_555 (O_555,N_8942,N_8125);
or UO_556 (O_556,N_9839,N_8295);
nor UO_557 (O_557,N_8560,N_9845);
nor UO_558 (O_558,N_9955,N_8662);
or UO_559 (O_559,N_9368,N_8048);
xnor UO_560 (O_560,N_9474,N_8904);
nor UO_561 (O_561,N_9323,N_9312);
nor UO_562 (O_562,N_9599,N_9335);
nor UO_563 (O_563,N_9890,N_8388);
nand UO_564 (O_564,N_9672,N_8616);
nand UO_565 (O_565,N_8654,N_9271);
or UO_566 (O_566,N_9416,N_8750);
and UO_567 (O_567,N_8283,N_8281);
and UO_568 (O_568,N_9815,N_9096);
nand UO_569 (O_569,N_8003,N_8316);
and UO_570 (O_570,N_9159,N_9104);
nand UO_571 (O_571,N_8441,N_8522);
nor UO_572 (O_572,N_9009,N_8830);
and UO_573 (O_573,N_8495,N_9315);
nand UO_574 (O_574,N_8688,N_8294);
or UO_575 (O_575,N_8882,N_8503);
or UO_576 (O_576,N_9309,N_8186);
or UO_577 (O_577,N_9205,N_9920);
and UO_578 (O_578,N_8832,N_8278);
or UO_579 (O_579,N_8806,N_8246);
nor UO_580 (O_580,N_8214,N_9837);
or UO_581 (O_581,N_8040,N_9422);
nand UO_582 (O_582,N_8848,N_9983);
nand UO_583 (O_583,N_8948,N_8731);
nand UO_584 (O_584,N_9726,N_8233);
and UO_585 (O_585,N_9383,N_9738);
nand UO_586 (O_586,N_9823,N_9640);
or UO_587 (O_587,N_9832,N_8477);
nor UO_588 (O_588,N_8655,N_8552);
nor UO_589 (O_589,N_9903,N_9083);
or UO_590 (O_590,N_9683,N_8397);
nor UO_591 (O_591,N_8701,N_8391);
nand UO_592 (O_592,N_8288,N_8455);
nor UO_593 (O_593,N_9217,N_9872);
nor UO_594 (O_594,N_8513,N_8618);
or UO_595 (O_595,N_8398,N_8227);
nand UO_596 (O_596,N_8426,N_8859);
nor UO_597 (O_597,N_9678,N_8970);
and UO_598 (O_598,N_8217,N_8345);
or UO_599 (O_599,N_9523,N_8195);
and UO_600 (O_600,N_8850,N_8011);
or UO_601 (O_601,N_9022,N_9607);
nor UO_602 (O_602,N_8463,N_9532);
and UO_603 (O_603,N_9179,N_9157);
or UO_604 (O_604,N_9986,N_9776);
nor UO_605 (O_605,N_9008,N_8664);
nand UO_606 (O_606,N_9241,N_8639);
or UO_607 (O_607,N_9696,N_8951);
or UO_608 (O_608,N_8979,N_8887);
and UO_609 (O_609,N_9116,N_9838);
nor UO_610 (O_610,N_8520,N_8357);
nand UO_611 (O_611,N_9027,N_8880);
nand UO_612 (O_612,N_8854,N_9298);
nor UO_613 (O_613,N_9074,N_9935);
nor UO_614 (O_614,N_9151,N_8313);
xor UO_615 (O_615,N_9253,N_9326);
nor UO_616 (O_616,N_8788,N_9354);
or UO_617 (O_617,N_9243,N_8181);
and UO_618 (O_618,N_8031,N_9883);
or UO_619 (O_619,N_8032,N_8626);
and UO_620 (O_620,N_8925,N_8177);
nor UO_621 (O_621,N_8783,N_8674);
nor UO_622 (O_622,N_8487,N_9508);
nand UO_623 (O_623,N_8722,N_8766);
xor UO_624 (O_624,N_8609,N_9162);
and UO_625 (O_625,N_8533,N_8285);
and UO_626 (O_626,N_9541,N_8267);
nor UO_627 (O_627,N_9810,N_8575);
nor UO_628 (O_628,N_8218,N_9554);
and UO_629 (O_629,N_8442,N_9910);
nor UO_630 (O_630,N_8147,N_8133);
or UO_631 (O_631,N_8746,N_9480);
and UO_632 (O_632,N_8417,N_8569);
and UO_633 (O_633,N_8265,N_9023);
nor UO_634 (O_634,N_8773,N_8992);
or UO_635 (O_635,N_9954,N_8461);
or UO_636 (O_636,N_9718,N_8793);
nand UO_637 (O_637,N_9661,N_8434);
nor UO_638 (O_638,N_8204,N_8311);
or UO_639 (O_639,N_9702,N_9834);
nand UO_640 (O_640,N_8039,N_9487);
nor UO_641 (O_641,N_9273,N_8271);
and UO_642 (O_642,N_9475,N_8730);
nand UO_643 (O_643,N_9533,N_9220);
or UO_644 (O_644,N_8564,N_9886);
nor UO_645 (O_645,N_9090,N_8352);
nor UO_646 (O_646,N_9859,N_9978);
nand UO_647 (O_647,N_9967,N_8408);
and UO_648 (O_648,N_8348,N_8529);
or UO_649 (O_649,N_9143,N_9374);
nand UO_650 (O_650,N_8936,N_9583);
or UO_651 (O_651,N_9710,N_8165);
and UO_652 (O_652,N_8579,N_8789);
nor UO_653 (O_653,N_9343,N_8990);
and UO_654 (O_654,N_9042,N_8926);
nor UO_655 (O_655,N_8707,N_9194);
nor UO_656 (O_656,N_8855,N_8269);
nand UO_657 (O_657,N_8930,N_9797);
or UO_658 (O_658,N_9876,N_9695);
or UO_659 (O_659,N_8433,N_9170);
or UO_660 (O_660,N_9314,N_9706);
and UO_661 (O_661,N_9686,N_8741);
nor UO_662 (O_662,N_8004,N_8550);
nand UO_663 (O_663,N_8916,N_9215);
xnor UO_664 (O_664,N_9385,N_9258);
and UO_665 (O_665,N_8824,N_8562);
nand UO_666 (O_666,N_8799,N_8742);
and UO_667 (O_667,N_8906,N_8547);
nand UO_668 (O_668,N_8876,N_9325);
nand UO_669 (O_669,N_8644,N_9613);
nor UO_670 (O_670,N_9275,N_9028);
and UO_671 (O_671,N_9985,N_8438);
and UO_672 (O_672,N_9352,N_8091);
and UO_673 (O_673,N_8905,N_9559);
or UO_674 (O_674,N_9302,N_9795);
nand UO_675 (O_675,N_8230,N_9602);
nor UO_676 (O_676,N_9115,N_9791);
and UO_677 (O_677,N_8405,N_8943);
and UO_678 (O_678,N_8009,N_8684);
nor UO_679 (O_679,N_9036,N_9854);
or UO_680 (O_680,N_9831,N_9505);
nor UO_681 (O_681,N_9558,N_9471);
nor UO_682 (O_682,N_8810,N_8412);
or UO_683 (O_683,N_9317,N_9756);
or UO_684 (O_684,N_8425,N_8194);
nand UO_685 (O_685,N_9984,N_9435);
or UO_686 (O_686,N_9804,N_8873);
nand UO_687 (O_687,N_9785,N_8619);
nor UO_688 (O_688,N_8997,N_8360);
or UO_689 (O_689,N_9990,N_9574);
and UO_690 (O_690,N_8258,N_9193);
or UO_691 (O_691,N_8539,N_9779);
nand UO_692 (O_692,N_9409,N_9485);
and UO_693 (O_693,N_8497,N_9569);
xnor UO_694 (O_694,N_8351,N_9211);
nor UO_695 (O_695,N_9781,N_9766);
nor UO_696 (O_696,N_8517,N_8580);
or UO_697 (O_697,N_8342,N_8116);
and UO_698 (O_698,N_9825,N_9576);
and UO_699 (O_699,N_8146,N_9556);
nand UO_700 (O_700,N_9786,N_9753);
nor UO_701 (O_701,N_9267,N_8601);
xor UO_702 (O_702,N_8718,N_8180);
and UO_703 (O_703,N_8798,N_8074);
nor UO_704 (O_704,N_8088,N_8166);
nor UO_705 (O_705,N_8251,N_9249);
nor UO_706 (O_706,N_8543,N_9105);
nand UO_707 (O_707,N_9130,N_9473);
nor UO_708 (O_708,N_8765,N_9921);
or UO_709 (O_709,N_8775,N_8008);
nand UO_710 (O_710,N_9472,N_8532);
nand UO_711 (O_711,N_8839,N_8112);
or UO_712 (O_712,N_9019,N_8981);
nor UO_713 (O_713,N_9133,N_8439);
nand UO_714 (O_714,N_8481,N_8591);
or UO_715 (O_715,N_9925,N_9849);
or UO_716 (O_716,N_9362,N_9236);
nand UO_717 (O_717,N_9924,N_9882);
nand UO_718 (O_718,N_8826,N_8123);
nand UO_719 (O_719,N_8350,N_8735);
and UO_720 (O_720,N_9844,N_8820);
nor UO_721 (O_721,N_9260,N_8329);
nor UO_722 (O_722,N_8178,N_8598);
xnor UO_723 (O_723,N_9553,N_8784);
or UO_724 (O_724,N_9972,N_9021);
xor UO_725 (O_725,N_9715,N_8049);
or UO_726 (O_726,N_9321,N_8653);
nor UO_727 (O_727,N_8811,N_8466);
and UO_728 (O_728,N_8944,N_9178);
nor UO_729 (O_729,N_9424,N_8554);
nor UO_730 (O_730,N_9188,N_9444);
nor UO_731 (O_731,N_8354,N_8364);
nand UO_732 (O_732,N_8063,N_8534);
and UO_733 (O_733,N_9709,N_9106);
nand UO_734 (O_734,N_8831,N_9107);
and UO_735 (O_735,N_9645,N_8413);
nor UO_736 (O_736,N_9853,N_9084);
nor UO_737 (O_737,N_9120,N_8155);
or UO_738 (O_738,N_9176,N_9773);
nor UO_739 (O_739,N_9651,N_8771);
or UO_740 (O_740,N_9132,N_8866);
nor UO_741 (O_741,N_8844,N_9139);
nor UO_742 (O_742,N_8699,N_8875);
or UO_743 (O_743,N_9356,N_9861);
nand UO_744 (O_744,N_8660,N_8280);
or UO_745 (O_745,N_8665,N_8010);
nand UO_746 (O_746,N_9698,N_9979);
nor UO_747 (O_747,N_8018,N_9601);
nor UO_748 (O_748,N_8891,N_9896);
or UO_749 (O_749,N_8558,N_9131);
or UO_750 (O_750,N_8871,N_8681);
nand UO_751 (O_751,N_8263,N_9470);
and UO_752 (O_752,N_9914,N_8102);
nor UO_753 (O_753,N_8794,N_8410);
nand UO_754 (O_754,N_9905,N_8917);
or UO_755 (O_755,N_8134,N_9867);
or UO_756 (O_756,N_9668,N_9427);
or UO_757 (O_757,N_9878,N_9397);
nor UO_758 (O_758,N_8652,N_8860);
nor UO_759 (O_759,N_9653,N_9079);
nand UO_760 (O_760,N_8594,N_9310);
and UO_761 (O_761,N_9809,N_9122);
nor UO_762 (O_762,N_8161,N_9254);
and UO_763 (O_763,N_8273,N_9016);
nand UO_764 (O_764,N_8462,N_9987);
nand UO_765 (O_765,N_8153,N_9761);
nor UO_766 (O_766,N_9464,N_9065);
and UO_767 (O_767,N_9458,N_8337);
and UO_768 (O_768,N_8163,N_8135);
or UO_769 (O_769,N_9570,N_9915);
or UO_770 (O_770,N_9824,N_9114);
and UO_771 (O_771,N_9893,N_9517);
nand UO_772 (O_772,N_9907,N_9526);
and UO_773 (O_773,N_8760,N_8192);
nand UO_774 (O_774,N_8344,N_8561);
nand UO_775 (O_775,N_8394,N_9063);
nand UO_776 (O_776,N_8400,N_8919);
or UO_777 (O_777,N_9771,N_9269);
nor UO_778 (O_778,N_8321,N_9737);
nor UO_779 (O_779,N_9746,N_9611);
nor UO_780 (O_780,N_8842,N_8132);
or UO_781 (O_781,N_8483,N_8471);
nand UO_782 (O_782,N_8239,N_8633);
and UO_783 (O_783,N_8179,N_8920);
nor UO_784 (O_784,N_9136,N_8914);
nand UO_785 (O_785,N_9072,N_9086);
and UO_786 (O_786,N_9190,N_9446);
and UO_787 (O_787,N_9659,N_9265);
and UO_788 (O_788,N_9163,N_8111);
or UO_789 (O_789,N_8484,N_8578);
and UO_790 (O_790,N_8999,N_8209);
or UO_791 (O_791,N_8051,N_9137);
nor UO_792 (O_792,N_9879,N_9953);
nor UO_793 (O_793,N_9923,N_9841);
and UO_794 (O_794,N_8518,N_9050);
and UO_795 (O_795,N_8738,N_8889);
or UO_796 (O_796,N_8712,N_9520);
or UO_797 (O_797,N_9415,N_8962);
nand UO_798 (O_798,N_8971,N_9462);
xnor UO_799 (O_799,N_8717,N_9525);
and UO_800 (O_800,N_9624,N_9324);
or UO_801 (O_801,N_8590,N_9964);
nand UO_802 (O_802,N_9864,N_9259);
nor UO_803 (O_803,N_8189,N_8082);
or UO_804 (O_804,N_9285,N_8221);
or UO_805 (O_805,N_9357,N_8038);
nand UO_806 (O_806,N_8173,N_9432);
or UO_807 (O_807,N_9411,N_8066);
nand UO_808 (O_808,N_8559,N_8490);
or UO_809 (O_809,N_8393,N_9814);
nor UO_810 (O_810,N_8566,N_9992);
or UO_811 (O_811,N_8510,N_8958);
and UO_812 (O_812,N_8406,N_9125);
nor UO_813 (O_813,N_8747,N_9588);
nand UO_814 (O_814,N_8467,N_9577);
or UO_815 (O_815,N_8693,N_8627);
nor UO_816 (O_816,N_9546,N_8473);
nand UO_817 (O_817,N_8349,N_9491);
nand UO_818 (O_818,N_9750,N_9610);
nand UO_819 (O_819,N_9828,N_8535);
nor UO_820 (O_820,N_8445,N_9431);
and UO_821 (O_821,N_8949,N_9184);
or UO_822 (O_822,N_8976,N_9404);
nand UO_823 (O_823,N_9293,N_8252);
xnor UO_824 (O_824,N_8224,N_8557);
or UO_825 (O_825,N_8900,N_8502);
nand UO_826 (O_826,N_9440,N_9866);
or UO_827 (O_827,N_9595,N_9180);
nand UO_828 (O_828,N_9642,N_9041);
nand UO_829 (O_829,N_9053,N_8058);
and UO_830 (O_830,N_8682,N_8511);
nand UO_831 (O_831,N_9340,N_9225);
and UO_832 (O_832,N_8658,N_9765);
nand UO_833 (O_833,N_8869,N_9774);
nand UO_834 (O_834,N_9857,N_8972);
or UO_835 (O_835,N_8713,N_9376);
or UO_836 (O_836,N_8076,N_8002);
or UO_837 (O_837,N_8457,N_9320);
nor UO_838 (O_838,N_8243,N_8715);
nor UO_839 (O_839,N_9918,N_8737);
nor UO_840 (O_840,N_8328,N_9305);
nand UO_841 (O_841,N_8108,N_8698);
and UO_842 (O_842,N_8046,N_9512);
and UO_843 (O_843,N_8432,N_8931);
or UO_844 (O_844,N_8634,N_9929);
and UO_845 (O_845,N_8427,N_9902);
and UO_846 (O_846,N_9840,N_9852);
nor UO_847 (O_847,N_9545,N_8857);
and UO_848 (O_848,N_8494,N_9294);
and UO_849 (O_849,N_9052,N_8913);
or UO_850 (O_850,N_9386,N_9219);
or UO_851 (O_851,N_9318,N_9297);
or UO_852 (O_852,N_8384,N_8680);
nand UO_853 (O_853,N_9503,N_8171);
nor UO_854 (O_854,N_8338,N_9931);
or UO_855 (O_855,N_9112,N_8107);
nand UO_856 (O_856,N_8160,N_8501);
nor UO_857 (O_857,N_8137,N_9247);
or UO_858 (O_858,N_9039,N_8044);
or UO_859 (O_859,N_8984,N_9299);
or UO_860 (O_860,N_9049,N_8312);
nand UO_861 (O_861,N_8659,N_8573);
or UO_862 (O_862,N_8139,N_8016);
or UO_863 (O_863,N_8987,N_8059);
nand UO_864 (O_864,N_9433,N_8809);
or UO_865 (O_865,N_9160,N_9778);
and UO_866 (O_866,N_8546,N_9479);
nor UO_867 (O_867,N_8315,N_8041);
and UO_868 (O_868,N_9671,N_9522);
and UO_869 (O_869,N_8813,N_8790);
and UO_870 (O_870,N_8097,N_8362);
or UO_871 (O_871,N_8157,N_9949);
nand UO_872 (O_872,N_8843,N_8028);
nand UO_873 (O_873,N_9663,N_8978);
or UO_874 (O_874,N_8877,N_9443);
or UO_875 (O_875,N_8755,N_8938);
nand UO_876 (O_876,N_9261,N_9142);
or UO_877 (O_877,N_9499,N_9806);
nor UO_878 (O_878,N_9351,N_9934);
or UO_879 (O_879,N_9003,N_9455);
nand UO_880 (O_880,N_9747,N_9032);
nor UO_881 (O_881,N_8373,N_9537);
nand UO_882 (O_882,N_9963,N_8973);
nand UO_883 (O_883,N_8289,N_9229);
and UO_884 (O_884,N_9256,N_8588);
xor UO_885 (O_885,N_9714,N_9146);
nor UO_886 (O_886,N_9207,N_8589);
and UO_887 (O_887,N_9637,N_8154);
nand UO_888 (O_888,N_9266,N_8087);
or UO_889 (O_889,N_9635,N_9865);
nor UO_890 (O_890,N_8697,N_9287);
nand UO_891 (O_891,N_8043,N_9262);
nand UO_892 (O_892,N_8056,N_8093);
nor UO_893 (O_893,N_9054,N_9477);
nand UO_894 (O_894,N_8064,N_8744);
nand UO_895 (O_895,N_9103,N_8042);
nor UO_896 (O_896,N_8989,N_8089);
and UO_897 (O_897,N_8689,N_9506);
or UO_898 (O_898,N_8318,N_8734);
nor UO_899 (O_899,N_9951,N_8519);
or UO_900 (O_900,N_9280,N_9419);
nand UO_901 (O_901,N_9429,N_8333);
and UO_902 (O_902,N_9904,N_8131);
nor UO_903 (O_903,N_9528,N_9246);
nand UO_904 (O_904,N_8663,N_9469);
nand UO_905 (O_905,N_9869,N_9378);
and UO_906 (O_906,N_9233,N_9015);
nand UO_907 (O_907,N_9024,N_9524);
or UO_908 (O_908,N_8966,N_9868);
or UO_909 (O_909,N_8435,N_9675);
nand UO_910 (O_910,N_8607,N_9733);
nand UO_911 (O_911,N_8612,N_9516);
nand UO_912 (O_912,N_8608,N_9780);
or UO_913 (O_913,N_8785,N_9677);
nor UO_914 (O_914,N_8536,N_9629);
nand UO_915 (O_915,N_8838,N_9342);
nor UO_916 (O_916,N_8197,N_9884);
xnor UO_917 (O_917,N_8823,N_8377);
nand UO_918 (O_918,N_9465,N_8678);
nand UO_919 (O_919,N_8901,N_9228);
nor UO_920 (O_920,N_9334,N_9012);
and UO_921 (O_921,N_9606,N_9734);
nand UO_922 (O_922,N_9183,N_9364);
or UO_923 (O_923,N_8724,N_9623);
nand UO_924 (O_924,N_8545,N_8572);
nor UO_925 (O_925,N_9620,N_8159);
nand UO_926 (O_926,N_9274,N_8299);
xnor UO_927 (O_927,N_8508,N_9448);
nor UO_928 (O_928,N_8489,N_9772);
and UO_929 (O_929,N_8890,N_9605);
nand UO_930 (O_930,N_9739,N_9270);
xnor UO_931 (O_931,N_8444,N_8708);
and UO_932 (O_932,N_8845,N_9888);
xnor UO_933 (O_933,N_8802,N_9398);
and UO_934 (O_934,N_9381,N_9091);
nor UO_935 (O_935,N_9519,N_9490);
nand UO_936 (O_936,N_9573,N_8369);
and UO_937 (O_937,N_9295,N_9760);
nand UO_938 (O_938,N_9895,N_9337);
nor UO_939 (O_939,N_9590,N_9451);
nor UO_940 (O_940,N_8402,N_9898);
nor UO_941 (O_941,N_9360,N_8386);
and UO_942 (O_942,N_8392,N_9842);
nor UO_943 (O_943,N_9488,N_9097);
xor UO_944 (O_944,N_9862,N_8275);
nor UO_945 (O_945,N_9192,N_8465);
nand UO_946 (O_946,N_8293,N_9662);
and UO_947 (O_947,N_9913,N_9349);
and UO_948 (O_948,N_8974,N_8493);
xnor UO_949 (O_949,N_8782,N_8053);
and UO_950 (O_950,N_9822,N_9550);
nand UO_951 (O_951,N_8950,N_8714);
nor UO_952 (O_952,N_8571,N_8017);
nor UO_953 (O_953,N_8726,N_9848);
nor UO_954 (O_954,N_8577,N_9226);
and UO_955 (O_955,N_8595,N_8308);
nor UO_956 (O_956,N_9093,N_8727);
nand UO_957 (O_957,N_9608,N_8399);
and UO_958 (O_958,N_8238,N_9721);
and UO_959 (O_959,N_9094,N_9673);
nor UO_960 (O_960,N_9591,N_8957);
or UO_961 (O_961,N_8201,N_8460);
nor UO_962 (O_962,N_9369,N_9501);
nand UO_963 (O_963,N_9875,N_8037);
nand UO_964 (O_964,N_9339,N_9069);
nand UO_965 (O_965,N_9382,N_8692);
nand UO_966 (O_966,N_8797,N_9248);
nand UO_967 (O_967,N_9329,N_8057);
and UO_968 (O_968,N_9609,N_9950);
and UO_969 (O_969,N_9333,N_8732);
and UO_970 (O_970,N_9539,N_9066);
and UO_971 (O_971,N_8856,N_8630);
nor UO_972 (O_972,N_9007,N_9657);
or UO_973 (O_973,N_8025,N_8113);
nand UO_974 (O_974,N_8953,N_8185);
or UO_975 (O_975,N_9701,N_8464);
nand UO_976 (O_976,N_8114,N_8005);
or UO_977 (O_977,N_9897,N_8320);
nand UO_978 (O_978,N_9906,N_8631);
or UO_979 (O_979,N_8167,N_9276);
or UO_980 (O_980,N_8816,N_8903);
or UO_981 (O_981,N_8307,N_9650);
and UO_982 (O_982,N_8657,N_8671);
or UO_983 (O_983,N_9540,N_8358);
or UO_984 (O_984,N_8581,N_9644);
and UO_985 (O_985,N_8879,N_8168);
nand UO_986 (O_986,N_8625,N_9014);
and UO_987 (O_987,N_9482,N_8286);
and UO_988 (O_988,N_8515,N_8403);
or UO_989 (O_989,N_8834,N_9402);
nor UO_990 (O_990,N_9742,N_9187);
nand UO_991 (O_991,N_9164,N_8768);
or UO_992 (O_992,N_8083,N_8459);
nand UO_993 (O_993,N_9616,N_8791);
or UO_994 (O_994,N_8940,N_9548);
nor UO_995 (O_995,N_9542,N_8452);
or UO_996 (O_996,N_9171,N_9741);
or UO_997 (O_997,N_9401,N_8211);
xnor UO_998 (O_998,N_9076,N_9080);
or UO_999 (O_999,N_9938,N_8428);
nor UO_1000 (O_1000,N_9886,N_9280);
nor UO_1001 (O_1001,N_8185,N_8353);
nand UO_1002 (O_1002,N_9286,N_8906);
or UO_1003 (O_1003,N_9896,N_8799);
and UO_1004 (O_1004,N_8657,N_9292);
and UO_1005 (O_1005,N_9159,N_9506);
or UO_1006 (O_1006,N_8484,N_9689);
nor UO_1007 (O_1007,N_9755,N_9838);
nor UO_1008 (O_1008,N_8854,N_8504);
or UO_1009 (O_1009,N_9790,N_8425);
and UO_1010 (O_1010,N_9984,N_8228);
nand UO_1011 (O_1011,N_8485,N_9015);
nor UO_1012 (O_1012,N_9068,N_9100);
or UO_1013 (O_1013,N_8597,N_9497);
and UO_1014 (O_1014,N_8002,N_9606);
and UO_1015 (O_1015,N_9729,N_9171);
nor UO_1016 (O_1016,N_9588,N_8062);
nand UO_1017 (O_1017,N_9144,N_9122);
and UO_1018 (O_1018,N_8037,N_9378);
nor UO_1019 (O_1019,N_8146,N_9828);
nor UO_1020 (O_1020,N_8749,N_9295);
nand UO_1021 (O_1021,N_9991,N_9416);
nand UO_1022 (O_1022,N_9696,N_8474);
and UO_1023 (O_1023,N_9096,N_9826);
xnor UO_1024 (O_1024,N_8052,N_9838);
or UO_1025 (O_1025,N_9000,N_9339);
and UO_1026 (O_1026,N_8969,N_9707);
nor UO_1027 (O_1027,N_8621,N_9184);
nand UO_1028 (O_1028,N_8637,N_9823);
xnor UO_1029 (O_1029,N_8085,N_9138);
nand UO_1030 (O_1030,N_8873,N_8664);
or UO_1031 (O_1031,N_9202,N_9743);
or UO_1032 (O_1032,N_9949,N_9338);
or UO_1033 (O_1033,N_9624,N_8474);
or UO_1034 (O_1034,N_8351,N_9101);
nor UO_1035 (O_1035,N_8890,N_8251);
and UO_1036 (O_1036,N_9669,N_8918);
nand UO_1037 (O_1037,N_9047,N_9212);
and UO_1038 (O_1038,N_9436,N_8322);
and UO_1039 (O_1039,N_8315,N_8310);
and UO_1040 (O_1040,N_9642,N_9308);
nor UO_1041 (O_1041,N_9932,N_8804);
or UO_1042 (O_1042,N_9770,N_9166);
and UO_1043 (O_1043,N_9012,N_8509);
and UO_1044 (O_1044,N_9444,N_8151);
and UO_1045 (O_1045,N_8219,N_9163);
or UO_1046 (O_1046,N_8279,N_8265);
nand UO_1047 (O_1047,N_8585,N_8188);
and UO_1048 (O_1048,N_8152,N_9715);
nand UO_1049 (O_1049,N_9651,N_9084);
and UO_1050 (O_1050,N_8702,N_9387);
nand UO_1051 (O_1051,N_8584,N_9226);
nand UO_1052 (O_1052,N_9910,N_9655);
and UO_1053 (O_1053,N_9201,N_8747);
nor UO_1054 (O_1054,N_9986,N_8939);
and UO_1055 (O_1055,N_9365,N_8796);
or UO_1056 (O_1056,N_9899,N_9369);
and UO_1057 (O_1057,N_8089,N_8211);
and UO_1058 (O_1058,N_9457,N_9911);
xor UO_1059 (O_1059,N_8867,N_9811);
nand UO_1060 (O_1060,N_8470,N_8634);
and UO_1061 (O_1061,N_8401,N_8870);
or UO_1062 (O_1062,N_9132,N_9829);
and UO_1063 (O_1063,N_9040,N_9426);
xnor UO_1064 (O_1064,N_8848,N_9438);
nor UO_1065 (O_1065,N_9166,N_9163);
and UO_1066 (O_1066,N_9330,N_9623);
nor UO_1067 (O_1067,N_8798,N_8147);
or UO_1068 (O_1068,N_9154,N_8414);
and UO_1069 (O_1069,N_9055,N_8307);
and UO_1070 (O_1070,N_9212,N_8724);
nor UO_1071 (O_1071,N_8985,N_8877);
xnor UO_1072 (O_1072,N_8058,N_8605);
and UO_1073 (O_1073,N_9020,N_9809);
nor UO_1074 (O_1074,N_8728,N_9937);
nand UO_1075 (O_1075,N_8399,N_8238);
or UO_1076 (O_1076,N_9745,N_8321);
and UO_1077 (O_1077,N_8225,N_8510);
or UO_1078 (O_1078,N_9299,N_8261);
nand UO_1079 (O_1079,N_9806,N_9442);
nor UO_1080 (O_1080,N_9303,N_9985);
nor UO_1081 (O_1081,N_8795,N_8909);
and UO_1082 (O_1082,N_9189,N_9047);
nand UO_1083 (O_1083,N_9497,N_8024);
nand UO_1084 (O_1084,N_8117,N_8869);
and UO_1085 (O_1085,N_8619,N_9486);
and UO_1086 (O_1086,N_8233,N_9021);
nand UO_1087 (O_1087,N_9236,N_9574);
xor UO_1088 (O_1088,N_9602,N_9045);
nor UO_1089 (O_1089,N_9404,N_8026);
and UO_1090 (O_1090,N_9923,N_9043);
nand UO_1091 (O_1091,N_8552,N_9653);
nand UO_1092 (O_1092,N_8248,N_9353);
nand UO_1093 (O_1093,N_8394,N_9709);
and UO_1094 (O_1094,N_8995,N_8242);
xor UO_1095 (O_1095,N_8572,N_9491);
nor UO_1096 (O_1096,N_8744,N_8222);
and UO_1097 (O_1097,N_9878,N_9966);
or UO_1098 (O_1098,N_8579,N_9763);
nor UO_1099 (O_1099,N_8462,N_9090);
or UO_1100 (O_1100,N_8209,N_9062);
nand UO_1101 (O_1101,N_9467,N_9970);
nor UO_1102 (O_1102,N_9779,N_8082);
and UO_1103 (O_1103,N_9419,N_8999);
nor UO_1104 (O_1104,N_9339,N_9643);
or UO_1105 (O_1105,N_9990,N_8372);
and UO_1106 (O_1106,N_9519,N_8137);
nor UO_1107 (O_1107,N_9714,N_8720);
xnor UO_1108 (O_1108,N_8289,N_9702);
or UO_1109 (O_1109,N_9664,N_8714);
and UO_1110 (O_1110,N_8483,N_9724);
nor UO_1111 (O_1111,N_8393,N_8062);
and UO_1112 (O_1112,N_8980,N_9514);
nand UO_1113 (O_1113,N_8615,N_8414);
and UO_1114 (O_1114,N_8680,N_9277);
and UO_1115 (O_1115,N_9413,N_8020);
nand UO_1116 (O_1116,N_8426,N_8358);
and UO_1117 (O_1117,N_9825,N_9188);
or UO_1118 (O_1118,N_8591,N_9045);
xnor UO_1119 (O_1119,N_8703,N_9804);
nor UO_1120 (O_1120,N_9803,N_8939);
nand UO_1121 (O_1121,N_9299,N_8969);
nand UO_1122 (O_1122,N_8708,N_8908);
nand UO_1123 (O_1123,N_8921,N_8711);
nand UO_1124 (O_1124,N_9972,N_9775);
and UO_1125 (O_1125,N_8089,N_9704);
nand UO_1126 (O_1126,N_8214,N_8131);
nand UO_1127 (O_1127,N_9272,N_9267);
and UO_1128 (O_1128,N_9246,N_9033);
or UO_1129 (O_1129,N_9445,N_9200);
or UO_1130 (O_1130,N_9211,N_8516);
or UO_1131 (O_1131,N_9925,N_9142);
nor UO_1132 (O_1132,N_9799,N_8406);
nor UO_1133 (O_1133,N_9517,N_9080);
nor UO_1134 (O_1134,N_8699,N_8199);
nand UO_1135 (O_1135,N_8731,N_9982);
and UO_1136 (O_1136,N_9542,N_9811);
or UO_1137 (O_1137,N_8082,N_8322);
and UO_1138 (O_1138,N_8471,N_9173);
nand UO_1139 (O_1139,N_8210,N_8851);
or UO_1140 (O_1140,N_9102,N_8546);
nor UO_1141 (O_1141,N_8261,N_8523);
or UO_1142 (O_1142,N_9459,N_8610);
nor UO_1143 (O_1143,N_8459,N_9816);
and UO_1144 (O_1144,N_9279,N_9077);
and UO_1145 (O_1145,N_9608,N_9122);
or UO_1146 (O_1146,N_8057,N_9170);
nand UO_1147 (O_1147,N_9082,N_9038);
and UO_1148 (O_1148,N_9117,N_8607);
or UO_1149 (O_1149,N_8159,N_8580);
or UO_1150 (O_1150,N_8590,N_9880);
nand UO_1151 (O_1151,N_9997,N_8306);
nand UO_1152 (O_1152,N_9392,N_9491);
nor UO_1153 (O_1153,N_9404,N_9301);
or UO_1154 (O_1154,N_9389,N_9547);
nand UO_1155 (O_1155,N_9564,N_8847);
nor UO_1156 (O_1156,N_8972,N_9021);
nand UO_1157 (O_1157,N_9059,N_8128);
and UO_1158 (O_1158,N_8669,N_8290);
or UO_1159 (O_1159,N_8921,N_8419);
and UO_1160 (O_1160,N_8168,N_8288);
and UO_1161 (O_1161,N_8947,N_8188);
or UO_1162 (O_1162,N_8463,N_8661);
xor UO_1163 (O_1163,N_9609,N_8828);
nor UO_1164 (O_1164,N_8206,N_9448);
and UO_1165 (O_1165,N_8543,N_9993);
and UO_1166 (O_1166,N_8147,N_9144);
and UO_1167 (O_1167,N_8346,N_9383);
or UO_1168 (O_1168,N_9764,N_8620);
and UO_1169 (O_1169,N_9361,N_8643);
nand UO_1170 (O_1170,N_8527,N_9617);
or UO_1171 (O_1171,N_9668,N_9056);
nand UO_1172 (O_1172,N_8267,N_8613);
nor UO_1173 (O_1173,N_8027,N_8707);
and UO_1174 (O_1174,N_9651,N_8136);
nand UO_1175 (O_1175,N_9946,N_9613);
nor UO_1176 (O_1176,N_9952,N_9886);
and UO_1177 (O_1177,N_8995,N_9028);
nor UO_1178 (O_1178,N_8144,N_9985);
and UO_1179 (O_1179,N_8783,N_9089);
nand UO_1180 (O_1180,N_8532,N_8721);
nor UO_1181 (O_1181,N_8817,N_9626);
nand UO_1182 (O_1182,N_8978,N_8121);
nand UO_1183 (O_1183,N_8024,N_9578);
or UO_1184 (O_1184,N_9509,N_8099);
nand UO_1185 (O_1185,N_8688,N_9876);
or UO_1186 (O_1186,N_9452,N_9551);
nand UO_1187 (O_1187,N_8906,N_8709);
or UO_1188 (O_1188,N_8068,N_9712);
nand UO_1189 (O_1189,N_9260,N_9248);
nor UO_1190 (O_1190,N_8447,N_9244);
nand UO_1191 (O_1191,N_9887,N_9328);
and UO_1192 (O_1192,N_8799,N_8829);
nor UO_1193 (O_1193,N_9448,N_8226);
nor UO_1194 (O_1194,N_8626,N_9633);
nor UO_1195 (O_1195,N_9486,N_9006);
nand UO_1196 (O_1196,N_9198,N_9277);
nand UO_1197 (O_1197,N_9993,N_8154);
and UO_1198 (O_1198,N_9758,N_8285);
xor UO_1199 (O_1199,N_9912,N_8573);
or UO_1200 (O_1200,N_8114,N_9155);
nand UO_1201 (O_1201,N_8459,N_8524);
and UO_1202 (O_1202,N_9162,N_9664);
and UO_1203 (O_1203,N_9156,N_8257);
or UO_1204 (O_1204,N_8564,N_9851);
or UO_1205 (O_1205,N_8095,N_8887);
xor UO_1206 (O_1206,N_8292,N_9209);
nand UO_1207 (O_1207,N_9341,N_9831);
nor UO_1208 (O_1208,N_8957,N_8439);
or UO_1209 (O_1209,N_9543,N_9555);
and UO_1210 (O_1210,N_8439,N_8518);
or UO_1211 (O_1211,N_9264,N_9478);
nand UO_1212 (O_1212,N_8353,N_9417);
or UO_1213 (O_1213,N_8815,N_9857);
and UO_1214 (O_1214,N_9561,N_8278);
or UO_1215 (O_1215,N_9114,N_8680);
and UO_1216 (O_1216,N_8580,N_9754);
nor UO_1217 (O_1217,N_8046,N_9392);
nor UO_1218 (O_1218,N_8912,N_9770);
or UO_1219 (O_1219,N_9416,N_8449);
nor UO_1220 (O_1220,N_8093,N_8414);
nor UO_1221 (O_1221,N_9606,N_9799);
and UO_1222 (O_1222,N_9796,N_8529);
and UO_1223 (O_1223,N_8101,N_9923);
or UO_1224 (O_1224,N_9780,N_8754);
or UO_1225 (O_1225,N_9166,N_8468);
nand UO_1226 (O_1226,N_9910,N_8799);
or UO_1227 (O_1227,N_8122,N_8322);
and UO_1228 (O_1228,N_9848,N_9414);
nor UO_1229 (O_1229,N_9082,N_8539);
or UO_1230 (O_1230,N_8194,N_9842);
nand UO_1231 (O_1231,N_9168,N_8711);
nand UO_1232 (O_1232,N_8827,N_9422);
and UO_1233 (O_1233,N_8595,N_8147);
nor UO_1234 (O_1234,N_8741,N_8284);
nor UO_1235 (O_1235,N_8606,N_9802);
nor UO_1236 (O_1236,N_8804,N_9048);
nor UO_1237 (O_1237,N_9743,N_9791);
nand UO_1238 (O_1238,N_8621,N_8662);
and UO_1239 (O_1239,N_9415,N_8654);
and UO_1240 (O_1240,N_9868,N_8824);
nand UO_1241 (O_1241,N_8732,N_8005);
nor UO_1242 (O_1242,N_8843,N_8239);
xor UO_1243 (O_1243,N_8268,N_8596);
nand UO_1244 (O_1244,N_9327,N_8364);
nor UO_1245 (O_1245,N_8767,N_8653);
nand UO_1246 (O_1246,N_8190,N_9124);
or UO_1247 (O_1247,N_9001,N_9035);
nor UO_1248 (O_1248,N_8605,N_8855);
xor UO_1249 (O_1249,N_8120,N_8708);
nor UO_1250 (O_1250,N_9269,N_8346);
and UO_1251 (O_1251,N_8727,N_8416);
and UO_1252 (O_1252,N_9613,N_8495);
nor UO_1253 (O_1253,N_9510,N_9290);
nor UO_1254 (O_1254,N_9493,N_8846);
nor UO_1255 (O_1255,N_9034,N_9529);
or UO_1256 (O_1256,N_8164,N_8215);
or UO_1257 (O_1257,N_9119,N_8136);
nand UO_1258 (O_1258,N_8201,N_9848);
nor UO_1259 (O_1259,N_8891,N_8510);
nand UO_1260 (O_1260,N_8393,N_8561);
or UO_1261 (O_1261,N_9805,N_9413);
or UO_1262 (O_1262,N_8366,N_8958);
xnor UO_1263 (O_1263,N_9062,N_9406);
and UO_1264 (O_1264,N_9175,N_9517);
and UO_1265 (O_1265,N_8392,N_8784);
and UO_1266 (O_1266,N_9989,N_8769);
nand UO_1267 (O_1267,N_9609,N_8074);
or UO_1268 (O_1268,N_8450,N_8934);
and UO_1269 (O_1269,N_8491,N_9607);
nor UO_1270 (O_1270,N_8566,N_8520);
or UO_1271 (O_1271,N_9279,N_8410);
or UO_1272 (O_1272,N_8914,N_9788);
nand UO_1273 (O_1273,N_8311,N_9529);
nor UO_1274 (O_1274,N_9122,N_8819);
nand UO_1275 (O_1275,N_8450,N_9604);
and UO_1276 (O_1276,N_8431,N_9589);
or UO_1277 (O_1277,N_9474,N_9405);
nor UO_1278 (O_1278,N_8120,N_9565);
nand UO_1279 (O_1279,N_9603,N_9611);
nor UO_1280 (O_1280,N_8518,N_9618);
or UO_1281 (O_1281,N_8276,N_8204);
nand UO_1282 (O_1282,N_8926,N_8580);
nor UO_1283 (O_1283,N_9787,N_9008);
or UO_1284 (O_1284,N_8023,N_9922);
xor UO_1285 (O_1285,N_9016,N_9445);
and UO_1286 (O_1286,N_9669,N_8275);
nand UO_1287 (O_1287,N_8318,N_9599);
and UO_1288 (O_1288,N_9609,N_8696);
or UO_1289 (O_1289,N_8874,N_9952);
or UO_1290 (O_1290,N_8885,N_9994);
and UO_1291 (O_1291,N_9831,N_8613);
nand UO_1292 (O_1292,N_8644,N_9612);
nand UO_1293 (O_1293,N_9623,N_9239);
xor UO_1294 (O_1294,N_8189,N_9938);
and UO_1295 (O_1295,N_9902,N_8609);
and UO_1296 (O_1296,N_9547,N_9548);
or UO_1297 (O_1297,N_9641,N_8510);
or UO_1298 (O_1298,N_8851,N_8035);
and UO_1299 (O_1299,N_9436,N_8814);
or UO_1300 (O_1300,N_9305,N_8285);
nand UO_1301 (O_1301,N_9590,N_8124);
nor UO_1302 (O_1302,N_8477,N_9836);
and UO_1303 (O_1303,N_8472,N_9781);
and UO_1304 (O_1304,N_8924,N_9913);
and UO_1305 (O_1305,N_8907,N_9801);
nand UO_1306 (O_1306,N_8126,N_8362);
and UO_1307 (O_1307,N_9173,N_8124);
nand UO_1308 (O_1308,N_9653,N_9643);
and UO_1309 (O_1309,N_8615,N_8195);
nand UO_1310 (O_1310,N_8942,N_8832);
nand UO_1311 (O_1311,N_9023,N_9185);
or UO_1312 (O_1312,N_8449,N_9767);
nand UO_1313 (O_1313,N_9991,N_9474);
nand UO_1314 (O_1314,N_8879,N_9776);
or UO_1315 (O_1315,N_8293,N_8917);
nor UO_1316 (O_1316,N_8915,N_8318);
or UO_1317 (O_1317,N_9653,N_9827);
or UO_1318 (O_1318,N_9429,N_8260);
nand UO_1319 (O_1319,N_8908,N_8029);
nor UO_1320 (O_1320,N_9809,N_9437);
and UO_1321 (O_1321,N_8819,N_8443);
and UO_1322 (O_1322,N_9237,N_8246);
or UO_1323 (O_1323,N_9234,N_9158);
and UO_1324 (O_1324,N_9431,N_9605);
nand UO_1325 (O_1325,N_8764,N_8251);
nor UO_1326 (O_1326,N_8519,N_8454);
nand UO_1327 (O_1327,N_9535,N_9762);
nand UO_1328 (O_1328,N_9059,N_8500);
and UO_1329 (O_1329,N_8995,N_8418);
or UO_1330 (O_1330,N_8952,N_8853);
and UO_1331 (O_1331,N_8569,N_8536);
nand UO_1332 (O_1332,N_9468,N_9751);
and UO_1333 (O_1333,N_9000,N_9848);
or UO_1334 (O_1334,N_8123,N_8906);
or UO_1335 (O_1335,N_9207,N_8816);
and UO_1336 (O_1336,N_8231,N_8683);
and UO_1337 (O_1337,N_9996,N_8141);
and UO_1338 (O_1338,N_9692,N_8692);
or UO_1339 (O_1339,N_9958,N_9052);
nand UO_1340 (O_1340,N_8416,N_8438);
or UO_1341 (O_1341,N_9762,N_8406);
nor UO_1342 (O_1342,N_8395,N_9081);
and UO_1343 (O_1343,N_9634,N_9423);
nor UO_1344 (O_1344,N_9630,N_8436);
nand UO_1345 (O_1345,N_8035,N_9695);
nand UO_1346 (O_1346,N_9713,N_9474);
or UO_1347 (O_1347,N_8816,N_9287);
or UO_1348 (O_1348,N_8118,N_9923);
and UO_1349 (O_1349,N_9588,N_8272);
nand UO_1350 (O_1350,N_8087,N_8475);
and UO_1351 (O_1351,N_9558,N_9130);
or UO_1352 (O_1352,N_9273,N_8809);
nand UO_1353 (O_1353,N_9907,N_8143);
or UO_1354 (O_1354,N_8106,N_8772);
or UO_1355 (O_1355,N_9102,N_9358);
xnor UO_1356 (O_1356,N_9434,N_9177);
nor UO_1357 (O_1357,N_9620,N_9023);
nor UO_1358 (O_1358,N_9943,N_9189);
nand UO_1359 (O_1359,N_9647,N_9048);
nor UO_1360 (O_1360,N_8149,N_9736);
nand UO_1361 (O_1361,N_9473,N_8149);
and UO_1362 (O_1362,N_9877,N_8896);
or UO_1363 (O_1363,N_9022,N_8978);
nor UO_1364 (O_1364,N_9924,N_8444);
nand UO_1365 (O_1365,N_9610,N_8121);
or UO_1366 (O_1366,N_9360,N_8660);
or UO_1367 (O_1367,N_9966,N_9208);
or UO_1368 (O_1368,N_8924,N_8637);
or UO_1369 (O_1369,N_8063,N_8869);
nand UO_1370 (O_1370,N_9812,N_9484);
xor UO_1371 (O_1371,N_9709,N_9357);
nand UO_1372 (O_1372,N_9724,N_8082);
and UO_1373 (O_1373,N_9654,N_8556);
and UO_1374 (O_1374,N_8132,N_9199);
and UO_1375 (O_1375,N_8688,N_8926);
nand UO_1376 (O_1376,N_8929,N_9973);
or UO_1377 (O_1377,N_9080,N_8876);
or UO_1378 (O_1378,N_8798,N_8709);
nor UO_1379 (O_1379,N_8767,N_8473);
nor UO_1380 (O_1380,N_9444,N_9317);
and UO_1381 (O_1381,N_9273,N_8106);
nand UO_1382 (O_1382,N_8313,N_9450);
xor UO_1383 (O_1383,N_9907,N_9462);
nor UO_1384 (O_1384,N_9654,N_8864);
and UO_1385 (O_1385,N_8355,N_8341);
nand UO_1386 (O_1386,N_8785,N_9168);
and UO_1387 (O_1387,N_9730,N_9372);
nor UO_1388 (O_1388,N_8757,N_9153);
or UO_1389 (O_1389,N_9500,N_8089);
or UO_1390 (O_1390,N_8636,N_8795);
xor UO_1391 (O_1391,N_9431,N_9365);
or UO_1392 (O_1392,N_9024,N_9704);
nand UO_1393 (O_1393,N_8924,N_9548);
or UO_1394 (O_1394,N_9231,N_8982);
or UO_1395 (O_1395,N_9841,N_9314);
and UO_1396 (O_1396,N_8654,N_8674);
nor UO_1397 (O_1397,N_9332,N_9824);
or UO_1398 (O_1398,N_9322,N_8322);
or UO_1399 (O_1399,N_8156,N_9297);
nand UO_1400 (O_1400,N_9569,N_9938);
nand UO_1401 (O_1401,N_9983,N_8858);
and UO_1402 (O_1402,N_9542,N_8759);
or UO_1403 (O_1403,N_9959,N_8464);
nor UO_1404 (O_1404,N_9231,N_9517);
or UO_1405 (O_1405,N_8860,N_9337);
or UO_1406 (O_1406,N_9318,N_8396);
nand UO_1407 (O_1407,N_8092,N_8157);
and UO_1408 (O_1408,N_8073,N_9618);
or UO_1409 (O_1409,N_9598,N_9719);
and UO_1410 (O_1410,N_9685,N_8434);
nor UO_1411 (O_1411,N_8384,N_8301);
and UO_1412 (O_1412,N_9538,N_9457);
xor UO_1413 (O_1413,N_9325,N_9901);
nor UO_1414 (O_1414,N_9303,N_8755);
nand UO_1415 (O_1415,N_9872,N_8210);
or UO_1416 (O_1416,N_8058,N_9478);
and UO_1417 (O_1417,N_9026,N_9523);
and UO_1418 (O_1418,N_8053,N_8568);
nand UO_1419 (O_1419,N_8523,N_8406);
nand UO_1420 (O_1420,N_8686,N_8623);
nand UO_1421 (O_1421,N_8753,N_9678);
or UO_1422 (O_1422,N_8707,N_8008);
nor UO_1423 (O_1423,N_8749,N_9885);
or UO_1424 (O_1424,N_8313,N_8853);
nor UO_1425 (O_1425,N_8877,N_8476);
nor UO_1426 (O_1426,N_9361,N_8503);
nor UO_1427 (O_1427,N_8189,N_9795);
nand UO_1428 (O_1428,N_8174,N_9516);
or UO_1429 (O_1429,N_9015,N_8282);
or UO_1430 (O_1430,N_8682,N_9738);
or UO_1431 (O_1431,N_9301,N_8122);
nand UO_1432 (O_1432,N_8582,N_8381);
or UO_1433 (O_1433,N_8940,N_9031);
or UO_1434 (O_1434,N_8752,N_8584);
xor UO_1435 (O_1435,N_9090,N_8217);
or UO_1436 (O_1436,N_8281,N_8602);
and UO_1437 (O_1437,N_9181,N_9358);
and UO_1438 (O_1438,N_9404,N_9400);
nand UO_1439 (O_1439,N_8972,N_9625);
xor UO_1440 (O_1440,N_8484,N_8189);
or UO_1441 (O_1441,N_9367,N_8774);
nand UO_1442 (O_1442,N_9922,N_9871);
or UO_1443 (O_1443,N_8892,N_8033);
and UO_1444 (O_1444,N_8688,N_9126);
nand UO_1445 (O_1445,N_9967,N_8141);
xor UO_1446 (O_1446,N_9792,N_8703);
nand UO_1447 (O_1447,N_9281,N_9478);
or UO_1448 (O_1448,N_8162,N_8762);
or UO_1449 (O_1449,N_9674,N_8716);
and UO_1450 (O_1450,N_8688,N_8100);
and UO_1451 (O_1451,N_8854,N_8074);
nor UO_1452 (O_1452,N_8315,N_9671);
nand UO_1453 (O_1453,N_8587,N_9397);
and UO_1454 (O_1454,N_8216,N_8164);
nand UO_1455 (O_1455,N_8845,N_9476);
or UO_1456 (O_1456,N_9334,N_9862);
and UO_1457 (O_1457,N_9734,N_8504);
nand UO_1458 (O_1458,N_9151,N_9207);
nor UO_1459 (O_1459,N_9045,N_9443);
or UO_1460 (O_1460,N_9620,N_8437);
and UO_1461 (O_1461,N_9619,N_8189);
and UO_1462 (O_1462,N_9621,N_8697);
nand UO_1463 (O_1463,N_8068,N_8012);
nor UO_1464 (O_1464,N_9525,N_8066);
nor UO_1465 (O_1465,N_9477,N_9597);
and UO_1466 (O_1466,N_9896,N_8190);
or UO_1467 (O_1467,N_8798,N_9267);
xnor UO_1468 (O_1468,N_8721,N_8701);
nor UO_1469 (O_1469,N_9739,N_9756);
or UO_1470 (O_1470,N_9407,N_9286);
nand UO_1471 (O_1471,N_9947,N_9584);
nor UO_1472 (O_1472,N_8773,N_9117);
nor UO_1473 (O_1473,N_9240,N_9329);
nand UO_1474 (O_1474,N_8805,N_8139);
and UO_1475 (O_1475,N_9919,N_9925);
and UO_1476 (O_1476,N_9550,N_9676);
and UO_1477 (O_1477,N_8092,N_8417);
or UO_1478 (O_1478,N_9586,N_8707);
nand UO_1479 (O_1479,N_9902,N_9487);
and UO_1480 (O_1480,N_8900,N_9754);
nand UO_1481 (O_1481,N_9462,N_9981);
xor UO_1482 (O_1482,N_8584,N_8883);
nand UO_1483 (O_1483,N_9286,N_9019);
nor UO_1484 (O_1484,N_9276,N_9589);
and UO_1485 (O_1485,N_8263,N_8953);
nand UO_1486 (O_1486,N_9423,N_8561);
or UO_1487 (O_1487,N_9456,N_9606);
or UO_1488 (O_1488,N_9610,N_8058);
nand UO_1489 (O_1489,N_8453,N_8707);
nand UO_1490 (O_1490,N_8481,N_8145);
nand UO_1491 (O_1491,N_8236,N_8624);
or UO_1492 (O_1492,N_8386,N_8564);
or UO_1493 (O_1493,N_9982,N_8550);
or UO_1494 (O_1494,N_8478,N_9895);
and UO_1495 (O_1495,N_9229,N_9801);
nand UO_1496 (O_1496,N_9929,N_9892);
or UO_1497 (O_1497,N_8212,N_8388);
nand UO_1498 (O_1498,N_9718,N_8189);
or UO_1499 (O_1499,N_8793,N_8667);
endmodule