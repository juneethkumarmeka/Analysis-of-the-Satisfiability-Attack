module basic_1000_10000_1500_5_levels_1xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_154,In_970);
or U1 (N_1,In_799,In_727);
nand U2 (N_2,In_233,In_926);
nand U3 (N_3,In_895,In_356);
and U4 (N_4,In_656,In_928);
nand U5 (N_5,In_107,In_355);
or U6 (N_6,In_674,In_683);
and U7 (N_7,In_743,In_574);
nor U8 (N_8,In_870,In_399);
and U9 (N_9,In_698,In_680);
or U10 (N_10,In_330,In_246);
or U11 (N_11,In_802,In_830);
nor U12 (N_12,In_263,In_883);
and U13 (N_13,In_591,In_853);
nand U14 (N_14,In_358,In_441);
or U15 (N_15,In_253,In_824);
nand U16 (N_16,In_639,In_160);
or U17 (N_17,In_22,In_368);
and U18 (N_18,In_181,In_527);
and U19 (N_19,In_859,In_347);
nor U20 (N_20,In_619,In_620);
or U21 (N_21,In_127,In_573);
or U22 (N_22,In_696,In_538);
nand U23 (N_23,In_18,In_403);
or U24 (N_24,In_924,In_159);
and U25 (N_25,In_633,In_820);
nor U26 (N_26,In_545,In_226);
nor U27 (N_27,In_668,In_670);
nor U28 (N_28,In_459,In_855);
or U29 (N_29,In_690,In_420);
nand U30 (N_30,In_319,In_148);
or U31 (N_31,In_842,In_204);
nor U32 (N_32,In_846,In_925);
nand U33 (N_33,In_558,In_961);
or U34 (N_34,In_50,In_406);
nor U35 (N_35,In_327,In_718);
nand U36 (N_36,In_348,In_292);
or U37 (N_37,In_264,In_163);
nor U38 (N_38,In_713,In_199);
nand U39 (N_39,In_845,In_207);
or U40 (N_40,In_222,In_386);
and U41 (N_41,In_528,In_273);
nand U42 (N_42,In_446,In_776);
and U43 (N_43,In_570,In_251);
and U44 (N_44,In_468,In_200);
nor U45 (N_45,In_499,In_655);
nor U46 (N_46,In_818,In_907);
or U47 (N_47,In_188,In_442);
xnor U48 (N_48,In_681,In_186);
or U49 (N_49,In_508,In_794);
nor U50 (N_50,In_290,In_274);
nor U51 (N_51,In_407,In_878);
or U52 (N_52,In_986,In_708);
nor U53 (N_53,In_989,In_647);
and U54 (N_54,In_83,In_85);
nand U55 (N_55,In_317,In_711);
nor U56 (N_56,In_152,In_780);
or U57 (N_57,In_534,In_79);
and U58 (N_58,In_267,In_487);
and U59 (N_59,In_360,In_749);
or U60 (N_60,In_493,In_747);
nor U61 (N_61,In_481,In_104);
nand U62 (N_62,In_387,In_774);
nor U63 (N_63,In_165,In_426);
or U64 (N_64,In_17,In_724);
or U65 (N_65,In_431,In_131);
nor U66 (N_66,In_423,In_645);
nor U67 (N_67,In_262,In_567);
and U68 (N_68,In_616,In_600);
nor U69 (N_69,In_722,In_583);
or U70 (N_70,In_192,In_930);
or U71 (N_71,In_587,In_404);
or U72 (N_72,In_359,In_892);
nand U73 (N_73,In_491,In_478);
nor U74 (N_74,In_754,In_427);
nor U75 (N_75,In_714,In_950);
or U76 (N_76,In_693,In_94);
xnor U77 (N_77,In_919,In_179);
or U78 (N_78,In_490,In_477);
nor U79 (N_79,In_784,In_444);
nand U80 (N_80,In_612,In_240);
nor U81 (N_81,In_585,In_161);
nand U82 (N_82,In_278,In_514);
nor U83 (N_83,In_972,In_133);
or U84 (N_84,In_617,In_45);
or U85 (N_85,In_461,In_332);
or U86 (N_86,In_309,In_544);
nand U87 (N_87,In_933,In_532);
nand U88 (N_88,In_298,In_5);
nor U89 (N_89,In_433,In_848);
or U90 (N_90,In_409,In_353);
nand U91 (N_91,In_429,In_949);
nor U92 (N_92,In_788,In_969);
nor U93 (N_93,In_768,In_962);
and U94 (N_94,In_266,In_6);
and U95 (N_95,In_627,In_125);
nor U96 (N_96,In_70,In_64);
nor U97 (N_97,In_737,In_502);
and U98 (N_98,In_384,In_470);
and U99 (N_99,In_213,In_957);
nand U100 (N_100,In_98,In_852);
and U101 (N_101,In_648,In_900);
nor U102 (N_102,In_95,In_629);
nor U103 (N_103,In_786,In_275);
or U104 (N_104,In_564,In_288);
and U105 (N_105,In_48,In_413);
or U106 (N_106,In_307,In_603);
or U107 (N_107,In_187,In_33);
and U108 (N_108,In_537,In_773);
nand U109 (N_109,In_568,In_334);
or U110 (N_110,In_157,In_847);
or U111 (N_111,In_272,In_843);
and U112 (N_112,In_15,In_868);
nor U113 (N_113,In_143,In_21);
nor U114 (N_114,In_31,In_662);
and U115 (N_115,In_116,In_676);
nand U116 (N_116,In_610,In_917);
nor U117 (N_117,In_497,In_471);
or U118 (N_118,In_74,In_227);
or U119 (N_119,In_942,In_230);
nor U120 (N_120,In_947,In_644);
and U121 (N_121,In_533,In_220);
and U122 (N_122,In_254,In_707);
nor U123 (N_123,In_341,In_577);
nor U124 (N_124,In_53,In_742);
nor U125 (N_125,In_910,In_88);
nor U126 (N_126,In_710,In_377);
nor U127 (N_127,In_554,In_229);
or U128 (N_128,In_876,In_828);
nor U129 (N_129,In_91,In_604);
or U130 (N_130,In_896,In_864);
nor U131 (N_131,In_315,In_785);
nand U132 (N_132,In_621,In_308);
or U133 (N_133,In_897,In_183);
nor U134 (N_134,In_92,In_775);
nor U135 (N_135,In_484,In_500);
nand U136 (N_136,In_256,In_260);
or U137 (N_137,In_185,In_173);
nand U138 (N_138,In_9,In_608);
nor U139 (N_139,In_951,In_29);
nor U140 (N_140,In_976,In_840);
nand U141 (N_141,In_232,In_562);
nor U142 (N_142,In_289,In_509);
and U143 (N_143,In_465,In_285);
or U144 (N_144,In_927,In_47);
or U145 (N_145,In_362,In_394);
and U146 (N_146,In_526,In_539);
nor U147 (N_147,In_905,In_988);
nand U148 (N_148,In_862,In_995);
nor U149 (N_149,In_849,In_993);
or U150 (N_150,In_419,In_808);
or U151 (N_151,In_501,In_357);
nand U152 (N_152,In_238,In_129);
or U153 (N_153,In_144,In_760);
and U154 (N_154,In_687,In_661);
nor U155 (N_155,In_956,In_39);
nand U156 (N_156,In_814,In_871);
nor U157 (N_157,In_964,In_126);
nand U158 (N_158,In_34,In_0);
nand U159 (N_159,In_496,In_176);
and U160 (N_160,In_36,In_618);
nor U161 (N_161,In_692,In_646);
nor U162 (N_162,In_219,In_415);
nor U163 (N_163,In_664,In_221);
or U164 (N_164,In_114,In_740);
nand U165 (N_165,In_863,In_520);
nand U166 (N_166,In_398,In_452);
nor U167 (N_167,In_703,In_4);
nand U168 (N_168,In_640,In_943);
nor U169 (N_169,In_807,In_110);
or U170 (N_170,In_42,In_944);
and U171 (N_171,In_804,In_198);
and U172 (N_172,In_803,In_738);
or U173 (N_173,In_825,In_450);
or U174 (N_174,In_1,In_689);
nand U175 (N_175,In_966,In_725);
or U176 (N_176,In_325,In_741);
or U177 (N_177,In_312,In_283);
and U178 (N_178,In_196,In_504);
or U179 (N_179,In_155,In_89);
nand U180 (N_180,In_886,In_35);
or U181 (N_181,In_417,In_375);
or U182 (N_182,In_873,In_867);
nand U183 (N_183,In_58,In_8);
or U184 (N_184,In_777,In_598);
or U185 (N_185,In_182,In_349);
nor U186 (N_186,In_701,In_581);
nor U187 (N_187,In_354,In_250);
nand U188 (N_188,In_593,In_630);
or U189 (N_189,In_702,In_236);
nand U190 (N_190,In_565,In_482);
nand U191 (N_191,In_904,In_920);
nor U192 (N_192,In_396,In_479);
or U193 (N_193,In_601,In_819);
and U194 (N_194,In_153,In_958);
nand U195 (N_195,In_467,In_584);
nand U196 (N_196,In_314,In_649);
or U197 (N_197,In_49,In_38);
and U198 (N_198,In_60,In_978);
and U199 (N_199,In_765,In_247);
nor U200 (N_200,In_424,In_832);
nand U201 (N_201,In_699,In_512);
or U202 (N_202,In_335,In_296);
nor U203 (N_203,In_26,In_323);
and U204 (N_204,In_136,In_68);
nor U205 (N_205,In_342,In_135);
nand U206 (N_206,In_453,In_967);
and U207 (N_207,In_752,In_899);
nand U208 (N_208,In_389,In_736);
nand U209 (N_209,In_180,In_77);
or U210 (N_210,In_968,In_320);
or U211 (N_211,In_469,In_178);
nand U212 (N_212,In_757,In_599);
nor U213 (N_213,In_810,In_297);
or U214 (N_214,In_37,In_430);
nand U215 (N_215,In_659,In_102);
nand U216 (N_216,In_709,In_936);
or U217 (N_217,In_428,In_145);
or U218 (N_218,In_498,In_548);
nand U219 (N_219,In_826,In_658);
and U220 (N_220,In_965,In_311);
and U221 (N_221,In_28,In_632);
and U222 (N_222,In_945,In_190);
and U223 (N_223,In_124,In_660);
or U224 (N_224,In_953,In_171);
nor U225 (N_225,In_522,In_553);
and U226 (N_226,In_540,In_797);
nor U227 (N_227,In_11,In_174);
nor U228 (N_228,In_184,In_997);
or U229 (N_229,In_51,In_130);
nand U230 (N_230,In_800,In_435);
or U231 (N_231,In_700,In_378);
nor U232 (N_232,In_322,In_25);
and U233 (N_233,In_231,In_705);
or U234 (N_234,In_913,In_594);
or U235 (N_235,In_975,In_437);
and U236 (N_236,In_379,In_759);
or U237 (N_237,In_418,In_438);
and U238 (N_238,In_669,In_510);
nand U239 (N_239,In_856,In_416);
nor U240 (N_240,In_78,In_328);
nor U241 (N_241,In_530,In_985);
nand U242 (N_242,In_929,In_898);
or U243 (N_243,In_373,In_269);
and U244 (N_244,In_255,In_475);
and U245 (N_245,In_352,In_571);
or U246 (N_246,In_141,In_909);
nor U247 (N_247,In_367,In_483);
nor U248 (N_248,In_866,In_869);
and U249 (N_249,In_243,In_998);
nand U250 (N_250,In_139,In_881);
or U251 (N_251,In_414,In_745);
and U252 (N_252,In_223,In_806);
nor U253 (N_253,In_434,In_813);
nand U254 (N_254,In_480,In_635);
or U255 (N_255,In_836,In_829);
and U256 (N_256,In_388,In_344);
nor U257 (N_257,In_979,In_57);
or U258 (N_258,In_282,In_789);
and U259 (N_259,In_889,In_903);
nor U260 (N_260,In_715,In_994);
nor U261 (N_261,In_542,In_63);
or U262 (N_262,In_147,In_579);
or U263 (N_263,In_506,In_474);
and U264 (N_264,In_756,In_884);
nor U265 (N_265,In_217,In_729);
nor U266 (N_266,In_887,In_425);
nor U267 (N_267,In_202,In_121);
nor U268 (N_268,In_167,In_287);
nor U269 (N_269,In_476,In_634);
nand U270 (N_270,In_891,In_981);
nand U271 (N_271,In_592,In_605);
nor U272 (N_272,In_411,In_595);
or U273 (N_273,In_191,In_128);
or U274 (N_274,In_578,In_370);
nand U275 (N_275,In_326,In_208);
or U276 (N_276,In_666,In_712);
nand U277 (N_277,In_543,In_796);
xnor U278 (N_278,In_303,In_206);
nor U279 (N_279,In_572,In_291);
nor U280 (N_280,In_313,In_665);
and U281 (N_281,In_732,In_463);
and U282 (N_282,In_694,In_305);
nor U283 (N_283,In_455,In_987);
nor U284 (N_284,In_921,In_963);
nand U285 (N_285,In_293,In_460);
nor U286 (N_286,In_383,In_150);
nor U287 (N_287,In_258,In_436);
or U288 (N_288,In_730,In_338);
or U289 (N_289,In_960,In_234);
and U290 (N_290,In_138,In_935);
or U291 (N_291,In_653,In_20);
xor U292 (N_292,In_324,In_955);
nand U293 (N_293,In_623,In_402);
or U294 (N_294,In_893,In_13);
nand U295 (N_295,In_902,In_170);
nand U296 (N_296,In_105,In_901);
nor U297 (N_297,In_582,In_652);
or U298 (N_298,In_778,In_525);
nand U299 (N_299,In_552,In_946);
nor U300 (N_300,In_811,In_62);
xor U301 (N_301,In_122,In_973);
and U302 (N_302,In_458,In_717);
or U303 (N_303,In_590,In_657);
or U304 (N_304,In_637,In_888);
or U305 (N_305,In_120,In_688);
nand U306 (N_306,In_654,In_23);
and U307 (N_307,In_164,In_90);
nor U308 (N_308,In_906,In_489);
nand U309 (N_309,In_763,In_959);
xnor U310 (N_310,In_753,In_492);
or U311 (N_311,In_97,In_823);
nand U312 (N_312,In_265,In_261);
nand U313 (N_313,In_52,In_546);
nor U314 (N_314,In_76,In_3);
nor U315 (N_315,In_462,In_445);
or U316 (N_316,In_268,In_835);
nor U317 (N_317,In_641,In_611);
and U318 (N_318,In_331,In_365);
nand U319 (N_319,In_563,In_551);
or U320 (N_320,In_890,In_142);
nor U321 (N_321,In_954,In_162);
and U322 (N_322,In_447,In_624);
and U323 (N_323,In_61,In_195);
and U324 (N_324,In_815,In_505);
or U325 (N_325,In_391,In_918);
or U326 (N_326,In_519,In_912);
nand U327 (N_327,In_783,In_941);
and U328 (N_328,In_100,In_614);
or U329 (N_329,In_735,In_12);
or U330 (N_330,In_16,In_343);
nor U331 (N_331,In_914,In_822);
nand U332 (N_332,In_561,In_932);
nand U333 (N_333,In_252,In_81);
nand U334 (N_334,In_597,In_201);
and U335 (N_335,In_177,In_249);
nand U336 (N_336,In_939,In_96);
and U337 (N_337,In_395,In_771);
or U338 (N_338,In_879,In_382);
nand U339 (N_339,In_750,In_675);
or U340 (N_340,In_118,In_137);
nor U341 (N_341,In_874,In_706);
nand U342 (N_342,In_682,In_559);
nand U343 (N_343,In_557,In_10);
or U344 (N_344,In_586,In_697);
or U345 (N_345,In_831,In_755);
and U346 (N_346,In_726,In_472);
or U347 (N_347,In_99,In_731);
and U348 (N_348,In_333,In_795);
or U349 (N_349,In_410,In_218);
nand U350 (N_350,In_41,In_259);
nor U351 (N_351,In_751,In_517);
nand U352 (N_352,In_916,In_106);
nor U353 (N_353,In_764,In_566);
nor U354 (N_354,In_279,In_511);
or U355 (N_355,In_366,In_390);
or U356 (N_356,In_734,In_7);
or U357 (N_357,In_875,In_704);
or U358 (N_358,In_767,In_860);
nand U359 (N_359,In_638,In_371);
nor U360 (N_360,In_55,In_271);
or U361 (N_361,In_790,In_369);
or U362 (N_362,In_245,In_672);
nand U363 (N_363,In_982,In_340);
or U364 (N_364,In_169,In_801);
and U365 (N_365,In_346,In_224);
nor U366 (N_366,In_345,In_515);
nor U367 (N_367,In_915,In_400);
nor U368 (N_368,In_865,In_295);
and U369 (N_369,In_556,In_321);
nand U370 (N_370,In_739,In_488);
and U371 (N_371,In_643,In_555);
nand U372 (N_372,In_82,In_938);
and U373 (N_373,In_772,In_19);
nor U374 (N_374,In_172,In_523);
or U375 (N_375,In_922,In_277);
nand U376 (N_376,In_280,In_923);
nand U377 (N_377,In_350,In_93);
nor U378 (N_378,In_242,In_123);
or U379 (N_379,In_529,In_787);
and U380 (N_380,In_550,In_27);
or U381 (N_381,In_209,In_983);
or U382 (N_382,In_650,In_113);
nand U383 (N_383,In_882,In_72);
and U384 (N_384,In_134,In_408);
nor U385 (N_385,In_766,In_575);
and U386 (N_386,In_834,In_677);
or U387 (N_387,In_156,In_215);
or U388 (N_388,In_651,In_239);
and U389 (N_389,In_588,In_996);
xor U390 (N_390,In_844,In_422);
or U391 (N_391,In_746,In_663);
nor U392 (N_392,In_103,In_301);
nor U393 (N_393,In_984,In_992);
or U394 (N_394,In_374,In_980);
and U395 (N_395,In_908,In_80);
and U396 (N_396,In_769,In_329);
or U397 (N_397,In_166,In_999);
and U398 (N_398,In_851,In_503);
and U399 (N_399,In_381,In_494);
or U400 (N_400,In_798,In_149);
nor U401 (N_401,In_337,In_894);
or U402 (N_402,In_560,In_791);
nand U403 (N_403,In_168,In_440);
or U404 (N_404,In_513,In_781);
nand U405 (N_405,In_609,In_65);
nor U406 (N_406,In_339,In_214);
nor U407 (N_407,In_432,In_940);
nor U408 (N_408,In_310,In_880);
nor U409 (N_409,In_971,In_576);
nor U410 (N_410,In_286,In_151);
and U411 (N_411,In_686,In_32);
or U412 (N_412,In_839,In_454);
nor U413 (N_413,In_306,In_46);
nor U414 (N_414,In_54,In_606);
nand U415 (N_415,In_535,In_235);
and U416 (N_416,In_507,In_678);
nor U417 (N_417,In_67,In_43);
nand U418 (N_418,In_631,In_937);
nand U419 (N_419,In_974,In_257);
nand U420 (N_420,In_281,In_376);
and U421 (N_421,In_580,In_112);
nand U422 (N_422,In_372,In_456);
or U423 (N_423,In_642,In_613);
nand U424 (N_424,In_158,In_516);
nand U425 (N_425,In_723,In_782);
and U426 (N_426,In_119,In_473);
nand U427 (N_427,In_952,In_841);
nor U428 (N_428,In_380,In_2);
and U429 (N_429,In_132,In_948);
and U430 (N_430,In_748,In_602);
and U431 (N_431,In_762,In_194);
nand U432 (N_432,In_607,In_486);
nor U433 (N_433,In_684,In_495);
and U434 (N_434,In_991,In_336);
nor U435 (N_435,In_837,In_237);
and U436 (N_436,In_596,In_363);
nand U437 (N_437,In_421,In_812);
or U438 (N_438,In_248,In_225);
nor U439 (N_439,In_877,In_30);
or U440 (N_440,In_75,In_84);
or U441 (N_441,In_569,In_86);
nand U442 (N_442,In_193,In_758);
and U443 (N_443,In_857,In_24);
and U444 (N_444,In_216,In_719);
or U445 (N_445,In_761,In_671);
and U446 (N_446,In_716,In_626);
or U447 (N_447,In_56,In_443);
and U448 (N_448,In_679,In_109);
and U449 (N_449,In_793,In_464);
and U450 (N_450,In_385,In_779);
nand U451 (N_451,In_549,In_304);
and U452 (N_452,In_721,In_361);
or U453 (N_453,In_547,In_451);
nand U454 (N_454,In_728,In_270);
nand U455 (N_455,In_197,In_589);
nand U456 (N_456,In_205,In_977);
or U457 (N_457,In_885,In_838);
nand U458 (N_458,In_827,In_111);
nor U459 (N_459,In_212,In_140);
and U460 (N_460,In_625,In_770);
and U461 (N_461,In_294,In_541);
nor U462 (N_462,In_189,In_397);
nor U463 (N_463,In_175,In_792);
nor U464 (N_464,In_816,In_817);
nor U465 (N_465,In_861,In_691);
nor U466 (N_466,In_720,In_733);
and U467 (N_467,In_44,In_615);
and U468 (N_468,In_87,In_59);
or U469 (N_469,In_316,In_524);
or U470 (N_470,In_66,In_628);
or U471 (N_471,In_805,In_673);
or U472 (N_472,In_115,In_401);
nor U473 (N_473,In_101,In_364);
and U474 (N_474,In_931,In_858);
nand U475 (N_475,In_521,In_318);
nand U476 (N_476,In_466,In_392);
and U477 (N_477,In_73,In_244);
and U478 (N_478,In_302,In_911);
nand U479 (N_479,In_531,In_854);
nor U480 (N_480,In_636,In_485);
nand U481 (N_481,In_351,In_536);
nor U482 (N_482,In_934,In_211);
nand U483 (N_483,In_412,In_228);
and U484 (N_484,In_108,In_821);
and U485 (N_485,In_117,In_518);
nand U486 (N_486,In_695,In_276);
or U487 (N_487,In_667,In_69);
or U488 (N_488,In_457,In_439);
or U489 (N_489,In_40,In_203);
and U490 (N_490,In_833,In_449);
xor U491 (N_491,In_299,In_146);
and U492 (N_492,In_685,In_14);
or U493 (N_493,In_241,In_990);
and U494 (N_494,In_210,In_622);
and U495 (N_495,In_405,In_809);
or U496 (N_496,In_71,In_284);
and U497 (N_497,In_744,In_872);
nand U498 (N_498,In_448,In_300);
nand U499 (N_499,In_850,In_393);
nor U500 (N_500,In_570,In_343);
or U501 (N_501,In_596,In_226);
nand U502 (N_502,In_972,In_720);
or U503 (N_503,In_411,In_645);
nand U504 (N_504,In_734,In_611);
nand U505 (N_505,In_80,In_891);
nor U506 (N_506,In_479,In_749);
nand U507 (N_507,In_686,In_272);
nor U508 (N_508,In_803,In_11);
nor U509 (N_509,In_27,In_938);
nor U510 (N_510,In_402,In_104);
nand U511 (N_511,In_999,In_718);
nand U512 (N_512,In_151,In_567);
and U513 (N_513,In_877,In_147);
and U514 (N_514,In_276,In_125);
nand U515 (N_515,In_741,In_806);
or U516 (N_516,In_497,In_565);
and U517 (N_517,In_233,In_576);
and U518 (N_518,In_983,In_562);
or U519 (N_519,In_976,In_159);
and U520 (N_520,In_919,In_272);
nor U521 (N_521,In_475,In_974);
or U522 (N_522,In_69,In_378);
nand U523 (N_523,In_523,In_535);
or U524 (N_524,In_138,In_721);
and U525 (N_525,In_823,In_651);
or U526 (N_526,In_22,In_735);
nand U527 (N_527,In_384,In_959);
and U528 (N_528,In_493,In_7);
nor U529 (N_529,In_665,In_174);
nand U530 (N_530,In_262,In_929);
or U531 (N_531,In_812,In_518);
or U532 (N_532,In_63,In_136);
nor U533 (N_533,In_30,In_52);
and U534 (N_534,In_536,In_363);
or U535 (N_535,In_538,In_137);
or U536 (N_536,In_250,In_796);
nand U537 (N_537,In_177,In_111);
nor U538 (N_538,In_980,In_144);
and U539 (N_539,In_364,In_760);
nor U540 (N_540,In_432,In_268);
nand U541 (N_541,In_597,In_273);
and U542 (N_542,In_631,In_934);
xnor U543 (N_543,In_733,In_293);
nand U544 (N_544,In_657,In_665);
or U545 (N_545,In_131,In_707);
nand U546 (N_546,In_202,In_546);
nor U547 (N_547,In_532,In_93);
nand U548 (N_548,In_344,In_257);
or U549 (N_549,In_660,In_470);
nor U550 (N_550,In_285,In_853);
and U551 (N_551,In_702,In_462);
or U552 (N_552,In_488,In_856);
nand U553 (N_553,In_403,In_3);
and U554 (N_554,In_800,In_53);
nand U555 (N_555,In_287,In_766);
nor U556 (N_556,In_604,In_376);
or U557 (N_557,In_223,In_776);
nor U558 (N_558,In_425,In_516);
or U559 (N_559,In_682,In_572);
or U560 (N_560,In_661,In_245);
xor U561 (N_561,In_735,In_858);
xor U562 (N_562,In_460,In_25);
and U563 (N_563,In_271,In_453);
or U564 (N_564,In_314,In_463);
nor U565 (N_565,In_130,In_758);
and U566 (N_566,In_439,In_913);
nor U567 (N_567,In_928,In_690);
nor U568 (N_568,In_64,In_463);
or U569 (N_569,In_966,In_864);
nand U570 (N_570,In_232,In_302);
or U571 (N_571,In_702,In_670);
or U572 (N_572,In_491,In_970);
or U573 (N_573,In_135,In_594);
nor U574 (N_574,In_287,In_117);
nand U575 (N_575,In_186,In_653);
nand U576 (N_576,In_481,In_675);
and U577 (N_577,In_112,In_623);
nand U578 (N_578,In_720,In_942);
or U579 (N_579,In_471,In_546);
and U580 (N_580,In_458,In_186);
and U581 (N_581,In_282,In_367);
nand U582 (N_582,In_646,In_401);
or U583 (N_583,In_556,In_620);
or U584 (N_584,In_935,In_429);
and U585 (N_585,In_563,In_520);
nand U586 (N_586,In_992,In_186);
and U587 (N_587,In_690,In_869);
or U588 (N_588,In_26,In_283);
and U589 (N_589,In_274,In_54);
nor U590 (N_590,In_803,In_419);
and U591 (N_591,In_263,In_39);
nand U592 (N_592,In_208,In_904);
and U593 (N_593,In_847,In_134);
nand U594 (N_594,In_350,In_88);
and U595 (N_595,In_722,In_422);
nand U596 (N_596,In_926,In_532);
nor U597 (N_597,In_915,In_175);
or U598 (N_598,In_597,In_866);
nor U599 (N_599,In_800,In_442);
nor U600 (N_600,In_838,In_207);
and U601 (N_601,In_753,In_689);
nor U602 (N_602,In_955,In_479);
and U603 (N_603,In_566,In_442);
nand U604 (N_604,In_968,In_309);
and U605 (N_605,In_239,In_336);
nand U606 (N_606,In_780,In_971);
nor U607 (N_607,In_678,In_211);
nor U608 (N_608,In_489,In_146);
and U609 (N_609,In_833,In_261);
nand U610 (N_610,In_490,In_957);
nor U611 (N_611,In_828,In_113);
nor U612 (N_612,In_416,In_120);
and U613 (N_613,In_79,In_602);
nor U614 (N_614,In_513,In_573);
or U615 (N_615,In_662,In_34);
xor U616 (N_616,In_593,In_480);
or U617 (N_617,In_456,In_894);
and U618 (N_618,In_691,In_396);
and U619 (N_619,In_86,In_410);
and U620 (N_620,In_785,In_74);
nand U621 (N_621,In_683,In_479);
nor U622 (N_622,In_717,In_481);
nor U623 (N_623,In_747,In_271);
or U624 (N_624,In_744,In_345);
nand U625 (N_625,In_551,In_205);
nand U626 (N_626,In_417,In_692);
and U627 (N_627,In_790,In_184);
and U628 (N_628,In_742,In_716);
and U629 (N_629,In_222,In_577);
and U630 (N_630,In_843,In_177);
and U631 (N_631,In_685,In_983);
or U632 (N_632,In_118,In_75);
nor U633 (N_633,In_929,In_341);
nor U634 (N_634,In_285,In_945);
nor U635 (N_635,In_258,In_337);
xnor U636 (N_636,In_32,In_637);
nor U637 (N_637,In_67,In_210);
or U638 (N_638,In_632,In_916);
or U639 (N_639,In_402,In_634);
nand U640 (N_640,In_589,In_923);
nand U641 (N_641,In_120,In_503);
or U642 (N_642,In_820,In_724);
nand U643 (N_643,In_301,In_893);
and U644 (N_644,In_175,In_721);
nor U645 (N_645,In_49,In_407);
or U646 (N_646,In_604,In_994);
and U647 (N_647,In_78,In_488);
nand U648 (N_648,In_848,In_205);
and U649 (N_649,In_280,In_385);
nand U650 (N_650,In_52,In_265);
and U651 (N_651,In_197,In_6);
nor U652 (N_652,In_332,In_37);
nor U653 (N_653,In_241,In_700);
nor U654 (N_654,In_652,In_17);
nand U655 (N_655,In_517,In_898);
or U656 (N_656,In_401,In_375);
nor U657 (N_657,In_371,In_792);
and U658 (N_658,In_873,In_894);
nand U659 (N_659,In_673,In_919);
or U660 (N_660,In_22,In_423);
or U661 (N_661,In_258,In_634);
or U662 (N_662,In_345,In_171);
nand U663 (N_663,In_535,In_445);
and U664 (N_664,In_102,In_382);
and U665 (N_665,In_816,In_366);
nand U666 (N_666,In_748,In_364);
or U667 (N_667,In_899,In_283);
or U668 (N_668,In_118,In_825);
nand U669 (N_669,In_579,In_872);
and U670 (N_670,In_909,In_845);
and U671 (N_671,In_768,In_156);
nand U672 (N_672,In_312,In_31);
nor U673 (N_673,In_856,In_449);
and U674 (N_674,In_401,In_26);
and U675 (N_675,In_957,In_581);
nor U676 (N_676,In_391,In_587);
nor U677 (N_677,In_114,In_885);
nand U678 (N_678,In_460,In_114);
nand U679 (N_679,In_74,In_211);
or U680 (N_680,In_365,In_984);
nand U681 (N_681,In_494,In_68);
nand U682 (N_682,In_363,In_916);
and U683 (N_683,In_146,In_308);
or U684 (N_684,In_288,In_641);
nor U685 (N_685,In_745,In_59);
nand U686 (N_686,In_603,In_65);
and U687 (N_687,In_84,In_762);
nor U688 (N_688,In_853,In_644);
or U689 (N_689,In_186,In_762);
or U690 (N_690,In_161,In_617);
nor U691 (N_691,In_110,In_262);
nand U692 (N_692,In_957,In_761);
nor U693 (N_693,In_851,In_365);
nor U694 (N_694,In_894,In_947);
xnor U695 (N_695,In_323,In_858);
nand U696 (N_696,In_38,In_148);
and U697 (N_697,In_785,In_374);
nand U698 (N_698,In_421,In_847);
and U699 (N_699,In_267,In_763);
nor U700 (N_700,In_773,In_334);
and U701 (N_701,In_110,In_808);
nor U702 (N_702,In_962,In_571);
nor U703 (N_703,In_982,In_434);
or U704 (N_704,In_23,In_848);
nor U705 (N_705,In_289,In_62);
and U706 (N_706,In_744,In_198);
and U707 (N_707,In_165,In_678);
or U708 (N_708,In_615,In_729);
nand U709 (N_709,In_131,In_178);
nand U710 (N_710,In_846,In_93);
and U711 (N_711,In_996,In_231);
nand U712 (N_712,In_946,In_953);
nand U713 (N_713,In_552,In_646);
or U714 (N_714,In_668,In_64);
and U715 (N_715,In_523,In_995);
or U716 (N_716,In_403,In_60);
nand U717 (N_717,In_953,In_330);
or U718 (N_718,In_512,In_146);
and U719 (N_719,In_686,In_186);
nand U720 (N_720,In_635,In_624);
nor U721 (N_721,In_264,In_814);
nand U722 (N_722,In_902,In_13);
nand U723 (N_723,In_532,In_206);
or U724 (N_724,In_749,In_851);
and U725 (N_725,In_744,In_642);
nor U726 (N_726,In_34,In_736);
nand U727 (N_727,In_292,In_476);
nor U728 (N_728,In_859,In_68);
nor U729 (N_729,In_472,In_195);
nand U730 (N_730,In_994,In_635);
nor U731 (N_731,In_535,In_947);
nand U732 (N_732,In_137,In_623);
nand U733 (N_733,In_368,In_571);
nand U734 (N_734,In_701,In_180);
nor U735 (N_735,In_204,In_519);
nor U736 (N_736,In_324,In_534);
nor U737 (N_737,In_496,In_210);
nand U738 (N_738,In_836,In_405);
and U739 (N_739,In_832,In_244);
and U740 (N_740,In_224,In_63);
or U741 (N_741,In_683,In_96);
and U742 (N_742,In_221,In_36);
and U743 (N_743,In_184,In_446);
nor U744 (N_744,In_424,In_103);
or U745 (N_745,In_106,In_325);
and U746 (N_746,In_374,In_574);
nor U747 (N_747,In_445,In_759);
or U748 (N_748,In_607,In_65);
nand U749 (N_749,In_349,In_650);
and U750 (N_750,In_89,In_610);
and U751 (N_751,In_433,In_856);
or U752 (N_752,In_950,In_414);
nand U753 (N_753,In_739,In_979);
and U754 (N_754,In_102,In_807);
and U755 (N_755,In_23,In_98);
or U756 (N_756,In_198,In_576);
and U757 (N_757,In_334,In_126);
nand U758 (N_758,In_212,In_594);
and U759 (N_759,In_589,In_532);
xnor U760 (N_760,In_837,In_763);
or U761 (N_761,In_13,In_132);
nor U762 (N_762,In_822,In_806);
and U763 (N_763,In_539,In_312);
nand U764 (N_764,In_288,In_603);
nand U765 (N_765,In_625,In_952);
nand U766 (N_766,In_17,In_712);
nor U767 (N_767,In_425,In_916);
and U768 (N_768,In_993,In_921);
nand U769 (N_769,In_339,In_446);
nor U770 (N_770,In_435,In_698);
nor U771 (N_771,In_31,In_636);
or U772 (N_772,In_561,In_912);
and U773 (N_773,In_198,In_603);
and U774 (N_774,In_59,In_338);
nand U775 (N_775,In_267,In_408);
nand U776 (N_776,In_306,In_786);
or U777 (N_777,In_179,In_920);
and U778 (N_778,In_296,In_505);
and U779 (N_779,In_401,In_421);
and U780 (N_780,In_219,In_738);
nand U781 (N_781,In_311,In_697);
nand U782 (N_782,In_524,In_145);
and U783 (N_783,In_783,In_991);
or U784 (N_784,In_25,In_95);
and U785 (N_785,In_253,In_126);
or U786 (N_786,In_140,In_348);
nand U787 (N_787,In_52,In_62);
or U788 (N_788,In_655,In_412);
or U789 (N_789,In_890,In_912);
nor U790 (N_790,In_808,In_2);
and U791 (N_791,In_810,In_944);
nor U792 (N_792,In_64,In_983);
and U793 (N_793,In_839,In_933);
or U794 (N_794,In_787,In_605);
nor U795 (N_795,In_356,In_34);
nor U796 (N_796,In_713,In_944);
or U797 (N_797,In_130,In_622);
nand U798 (N_798,In_962,In_825);
nand U799 (N_799,In_390,In_257);
nor U800 (N_800,In_200,In_381);
nor U801 (N_801,In_592,In_546);
or U802 (N_802,In_798,In_83);
nand U803 (N_803,In_37,In_977);
and U804 (N_804,In_154,In_61);
nand U805 (N_805,In_262,In_698);
nand U806 (N_806,In_751,In_202);
nand U807 (N_807,In_400,In_896);
nand U808 (N_808,In_331,In_896);
or U809 (N_809,In_788,In_123);
and U810 (N_810,In_223,In_69);
nand U811 (N_811,In_297,In_961);
or U812 (N_812,In_503,In_665);
nor U813 (N_813,In_981,In_575);
nand U814 (N_814,In_880,In_79);
nor U815 (N_815,In_179,In_88);
nand U816 (N_816,In_530,In_212);
and U817 (N_817,In_78,In_445);
and U818 (N_818,In_369,In_819);
or U819 (N_819,In_173,In_400);
or U820 (N_820,In_495,In_783);
nand U821 (N_821,In_245,In_940);
nand U822 (N_822,In_656,In_846);
and U823 (N_823,In_42,In_633);
or U824 (N_824,In_54,In_639);
nor U825 (N_825,In_889,In_672);
and U826 (N_826,In_941,In_335);
and U827 (N_827,In_917,In_857);
and U828 (N_828,In_913,In_287);
or U829 (N_829,In_785,In_147);
and U830 (N_830,In_595,In_379);
nand U831 (N_831,In_531,In_793);
nand U832 (N_832,In_491,In_396);
nor U833 (N_833,In_313,In_479);
or U834 (N_834,In_322,In_145);
nor U835 (N_835,In_747,In_93);
nor U836 (N_836,In_75,In_217);
and U837 (N_837,In_718,In_359);
nand U838 (N_838,In_402,In_237);
nand U839 (N_839,In_123,In_592);
nor U840 (N_840,In_58,In_599);
nor U841 (N_841,In_678,In_371);
or U842 (N_842,In_419,In_59);
or U843 (N_843,In_273,In_963);
nor U844 (N_844,In_848,In_701);
nor U845 (N_845,In_540,In_765);
nor U846 (N_846,In_791,In_549);
or U847 (N_847,In_645,In_409);
nand U848 (N_848,In_946,In_598);
nand U849 (N_849,In_176,In_618);
or U850 (N_850,In_792,In_747);
nand U851 (N_851,In_663,In_85);
and U852 (N_852,In_107,In_858);
and U853 (N_853,In_215,In_126);
or U854 (N_854,In_248,In_586);
xnor U855 (N_855,In_226,In_541);
nor U856 (N_856,In_851,In_394);
and U857 (N_857,In_320,In_654);
nor U858 (N_858,In_913,In_768);
and U859 (N_859,In_3,In_165);
or U860 (N_860,In_732,In_538);
nand U861 (N_861,In_909,In_28);
nand U862 (N_862,In_969,In_58);
and U863 (N_863,In_319,In_53);
and U864 (N_864,In_699,In_164);
nand U865 (N_865,In_934,In_389);
or U866 (N_866,In_735,In_590);
xor U867 (N_867,In_708,In_879);
nor U868 (N_868,In_897,In_603);
or U869 (N_869,In_166,In_883);
or U870 (N_870,In_867,In_988);
nand U871 (N_871,In_828,In_491);
and U872 (N_872,In_504,In_359);
xor U873 (N_873,In_406,In_685);
and U874 (N_874,In_718,In_140);
or U875 (N_875,In_411,In_507);
nor U876 (N_876,In_268,In_722);
and U877 (N_877,In_987,In_570);
nand U878 (N_878,In_825,In_979);
nor U879 (N_879,In_271,In_464);
or U880 (N_880,In_860,In_123);
nor U881 (N_881,In_277,In_647);
nor U882 (N_882,In_782,In_848);
or U883 (N_883,In_652,In_562);
or U884 (N_884,In_361,In_500);
nor U885 (N_885,In_802,In_289);
or U886 (N_886,In_658,In_611);
or U887 (N_887,In_552,In_165);
and U888 (N_888,In_344,In_54);
or U889 (N_889,In_801,In_851);
and U890 (N_890,In_782,In_525);
nor U891 (N_891,In_414,In_422);
and U892 (N_892,In_93,In_945);
or U893 (N_893,In_85,In_853);
nor U894 (N_894,In_522,In_891);
nand U895 (N_895,In_971,In_422);
nor U896 (N_896,In_485,In_960);
or U897 (N_897,In_851,In_901);
nor U898 (N_898,In_205,In_42);
nand U899 (N_899,In_919,In_948);
or U900 (N_900,In_830,In_678);
and U901 (N_901,In_831,In_73);
or U902 (N_902,In_531,In_859);
and U903 (N_903,In_862,In_997);
nand U904 (N_904,In_259,In_716);
nand U905 (N_905,In_456,In_622);
nor U906 (N_906,In_176,In_987);
nor U907 (N_907,In_152,In_731);
and U908 (N_908,In_64,In_589);
and U909 (N_909,In_911,In_967);
or U910 (N_910,In_765,In_848);
or U911 (N_911,In_135,In_761);
nor U912 (N_912,In_941,In_833);
xor U913 (N_913,In_377,In_796);
or U914 (N_914,In_180,In_28);
or U915 (N_915,In_444,In_655);
nand U916 (N_916,In_909,In_865);
nand U917 (N_917,In_323,In_180);
and U918 (N_918,In_489,In_161);
and U919 (N_919,In_915,In_984);
nand U920 (N_920,In_447,In_569);
nor U921 (N_921,In_214,In_623);
and U922 (N_922,In_876,In_590);
or U923 (N_923,In_139,In_909);
nand U924 (N_924,In_74,In_748);
and U925 (N_925,In_530,In_521);
nor U926 (N_926,In_353,In_510);
or U927 (N_927,In_453,In_46);
or U928 (N_928,In_154,In_604);
nand U929 (N_929,In_46,In_682);
and U930 (N_930,In_43,In_546);
or U931 (N_931,In_495,In_740);
nand U932 (N_932,In_69,In_326);
or U933 (N_933,In_777,In_812);
nand U934 (N_934,In_12,In_794);
xnor U935 (N_935,In_321,In_859);
nor U936 (N_936,In_146,In_691);
or U937 (N_937,In_990,In_107);
and U938 (N_938,In_215,In_319);
nand U939 (N_939,In_21,In_166);
nor U940 (N_940,In_461,In_537);
nor U941 (N_941,In_464,In_803);
or U942 (N_942,In_930,In_568);
nand U943 (N_943,In_273,In_349);
nor U944 (N_944,In_780,In_162);
and U945 (N_945,In_249,In_286);
nor U946 (N_946,In_36,In_477);
or U947 (N_947,In_456,In_388);
nor U948 (N_948,In_983,In_356);
nand U949 (N_949,In_1,In_900);
and U950 (N_950,In_456,In_481);
or U951 (N_951,In_277,In_691);
nand U952 (N_952,In_859,In_588);
nor U953 (N_953,In_144,In_187);
nor U954 (N_954,In_576,In_801);
or U955 (N_955,In_428,In_820);
or U956 (N_956,In_916,In_774);
and U957 (N_957,In_874,In_141);
nand U958 (N_958,In_673,In_348);
nand U959 (N_959,In_47,In_475);
or U960 (N_960,In_286,In_798);
nor U961 (N_961,In_154,In_627);
nor U962 (N_962,In_31,In_672);
or U963 (N_963,In_487,In_418);
nand U964 (N_964,In_723,In_491);
nor U965 (N_965,In_274,In_249);
or U966 (N_966,In_957,In_205);
xor U967 (N_967,In_68,In_217);
and U968 (N_968,In_154,In_789);
or U969 (N_969,In_740,In_93);
or U970 (N_970,In_134,In_523);
and U971 (N_971,In_800,In_661);
or U972 (N_972,In_37,In_641);
nand U973 (N_973,In_783,In_932);
or U974 (N_974,In_807,In_601);
or U975 (N_975,In_953,In_92);
nor U976 (N_976,In_732,In_312);
nand U977 (N_977,In_359,In_502);
nand U978 (N_978,In_205,In_433);
nor U979 (N_979,In_581,In_187);
and U980 (N_980,In_653,In_638);
nand U981 (N_981,In_466,In_158);
nor U982 (N_982,In_4,In_532);
or U983 (N_983,In_644,In_394);
nand U984 (N_984,In_393,In_124);
and U985 (N_985,In_680,In_61);
or U986 (N_986,In_474,In_144);
and U987 (N_987,In_636,In_589);
or U988 (N_988,In_528,In_443);
nand U989 (N_989,In_461,In_204);
and U990 (N_990,In_748,In_48);
nand U991 (N_991,In_792,In_387);
nand U992 (N_992,In_12,In_556);
and U993 (N_993,In_178,In_987);
nor U994 (N_994,In_24,In_116);
nor U995 (N_995,In_699,In_497);
and U996 (N_996,In_227,In_331);
nor U997 (N_997,In_60,In_24);
nand U998 (N_998,In_173,In_704);
nor U999 (N_999,In_825,In_217);
nor U1000 (N_1000,In_557,In_625);
or U1001 (N_1001,In_321,In_663);
nor U1002 (N_1002,In_947,In_185);
nand U1003 (N_1003,In_769,In_653);
nor U1004 (N_1004,In_541,In_949);
nor U1005 (N_1005,In_367,In_612);
and U1006 (N_1006,In_581,In_376);
nand U1007 (N_1007,In_131,In_396);
nand U1008 (N_1008,In_366,In_881);
and U1009 (N_1009,In_896,In_409);
nor U1010 (N_1010,In_659,In_372);
nand U1011 (N_1011,In_170,In_647);
nor U1012 (N_1012,In_397,In_292);
or U1013 (N_1013,In_512,In_326);
nor U1014 (N_1014,In_209,In_907);
and U1015 (N_1015,In_938,In_868);
nor U1016 (N_1016,In_808,In_668);
and U1017 (N_1017,In_519,In_137);
and U1018 (N_1018,In_396,In_438);
and U1019 (N_1019,In_726,In_387);
nor U1020 (N_1020,In_937,In_653);
and U1021 (N_1021,In_359,In_637);
and U1022 (N_1022,In_796,In_552);
nand U1023 (N_1023,In_714,In_443);
nor U1024 (N_1024,In_355,In_211);
and U1025 (N_1025,In_404,In_492);
nand U1026 (N_1026,In_217,In_440);
or U1027 (N_1027,In_927,In_768);
or U1028 (N_1028,In_962,In_351);
or U1029 (N_1029,In_751,In_254);
or U1030 (N_1030,In_754,In_645);
or U1031 (N_1031,In_328,In_584);
nand U1032 (N_1032,In_802,In_755);
nand U1033 (N_1033,In_29,In_757);
nor U1034 (N_1034,In_952,In_350);
nor U1035 (N_1035,In_454,In_986);
nand U1036 (N_1036,In_837,In_710);
and U1037 (N_1037,In_964,In_974);
nand U1038 (N_1038,In_654,In_559);
and U1039 (N_1039,In_828,In_256);
or U1040 (N_1040,In_95,In_928);
xor U1041 (N_1041,In_904,In_136);
and U1042 (N_1042,In_104,In_803);
nand U1043 (N_1043,In_974,In_205);
and U1044 (N_1044,In_571,In_64);
or U1045 (N_1045,In_364,In_643);
nor U1046 (N_1046,In_861,In_490);
nor U1047 (N_1047,In_809,In_64);
nand U1048 (N_1048,In_55,In_962);
nand U1049 (N_1049,In_144,In_116);
and U1050 (N_1050,In_996,In_368);
nor U1051 (N_1051,In_709,In_980);
or U1052 (N_1052,In_616,In_767);
nand U1053 (N_1053,In_955,In_768);
nor U1054 (N_1054,In_299,In_128);
or U1055 (N_1055,In_539,In_615);
nand U1056 (N_1056,In_63,In_845);
nand U1057 (N_1057,In_43,In_481);
nand U1058 (N_1058,In_186,In_382);
nand U1059 (N_1059,In_35,In_872);
nor U1060 (N_1060,In_611,In_364);
nor U1061 (N_1061,In_983,In_7);
and U1062 (N_1062,In_445,In_878);
or U1063 (N_1063,In_618,In_933);
nand U1064 (N_1064,In_478,In_320);
nand U1065 (N_1065,In_530,In_848);
or U1066 (N_1066,In_740,In_285);
nor U1067 (N_1067,In_813,In_846);
nand U1068 (N_1068,In_813,In_180);
and U1069 (N_1069,In_762,In_444);
nand U1070 (N_1070,In_631,In_856);
and U1071 (N_1071,In_444,In_617);
nor U1072 (N_1072,In_605,In_831);
nand U1073 (N_1073,In_954,In_445);
or U1074 (N_1074,In_875,In_482);
and U1075 (N_1075,In_983,In_504);
nand U1076 (N_1076,In_620,In_978);
nand U1077 (N_1077,In_496,In_963);
nor U1078 (N_1078,In_888,In_540);
nand U1079 (N_1079,In_541,In_170);
and U1080 (N_1080,In_232,In_171);
nand U1081 (N_1081,In_827,In_416);
or U1082 (N_1082,In_908,In_486);
nor U1083 (N_1083,In_143,In_827);
nor U1084 (N_1084,In_302,In_43);
nand U1085 (N_1085,In_263,In_962);
and U1086 (N_1086,In_669,In_958);
or U1087 (N_1087,In_497,In_369);
and U1088 (N_1088,In_481,In_786);
nor U1089 (N_1089,In_873,In_471);
nor U1090 (N_1090,In_743,In_423);
or U1091 (N_1091,In_97,In_878);
nand U1092 (N_1092,In_703,In_277);
nand U1093 (N_1093,In_944,In_514);
nor U1094 (N_1094,In_513,In_648);
nor U1095 (N_1095,In_6,In_37);
nand U1096 (N_1096,In_748,In_244);
and U1097 (N_1097,In_562,In_690);
nor U1098 (N_1098,In_319,In_212);
nand U1099 (N_1099,In_23,In_148);
nor U1100 (N_1100,In_734,In_125);
or U1101 (N_1101,In_960,In_181);
nand U1102 (N_1102,In_763,In_431);
or U1103 (N_1103,In_895,In_754);
nand U1104 (N_1104,In_106,In_333);
nor U1105 (N_1105,In_189,In_349);
and U1106 (N_1106,In_619,In_867);
and U1107 (N_1107,In_761,In_266);
or U1108 (N_1108,In_568,In_919);
nand U1109 (N_1109,In_521,In_194);
or U1110 (N_1110,In_917,In_26);
xnor U1111 (N_1111,In_583,In_897);
or U1112 (N_1112,In_348,In_606);
nand U1113 (N_1113,In_495,In_52);
or U1114 (N_1114,In_718,In_125);
or U1115 (N_1115,In_614,In_167);
and U1116 (N_1116,In_173,In_475);
and U1117 (N_1117,In_376,In_561);
and U1118 (N_1118,In_695,In_274);
nand U1119 (N_1119,In_580,In_176);
or U1120 (N_1120,In_788,In_120);
and U1121 (N_1121,In_969,In_132);
nor U1122 (N_1122,In_473,In_56);
or U1123 (N_1123,In_734,In_707);
and U1124 (N_1124,In_972,In_45);
nor U1125 (N_1125,In_338,In_798);
and U1126 (N_1126,In_841,In_365);
or U1127 (N_1127,In_17,In_177);
or U1128 (N_1128,In_494,In_754);
or U1129 (N_1129,In_965,In_476);
and U1130 (N_1130,In_566,In_513);
nor U1131 (N_1131,In_771,In_179);
and U1132 (N_1132,In_486,In_804);
nor U1133 (N_1133,In_383,In_215);
or U1134 (N_1134,In_329,In_372);
and U1135 (N_1135,In_356,In_484);
or U1136 (N_1136,In_334,In_173);
and U1137 (N_1137,In_174,In_774);
or U1138 (N_1138,In_23,In_474);
and U1139 (N_1139,In_495,In_829);
or U1140 (N_1140,In_874,In_450);
or U1141 (N_1141,In_48,In_23);
and U1142 (N_1142,In_144,In_674);
nor U1143 (N_1143,In_728,In_645);
nand U1144 (N_1144,In_310,In_799);
nor U1145 (N_1145,In_835,In_25);
and U1146 (N_1146,In_432,In_705);
or U1147 (N_1147,In_652,In_271);
nand U1148 (N_1148,In_107,In_692);
nand U1149 (N_1149,In_633,In_607);
nand U1150 (N_1150,In_907,In_545);
and U1151 (N_1151,In_893,In_744);
and U1152 (N_1152,In_503,In_782);
and U1153 (N_1153,In_709,In_824);
or U1154 (N_1154,In_898,In_59);
or U1155 (N_1155,In_620,In_640);
nor U1156 (N_1156,In_767,In_575);
or U1157 (N_1157,In_858,In_216);
nor U1158 (N_1158,In_339,In_285);
nor U1159 (N_1159,In_372,In_547);
nor U1160 (N_1160,In_100,In_6);
nor U1161 (N_1161,In_188,In_744);
nand U1162 (N_1162,In_46,In_455);
xor U1163 (N_1163,In_312,In_435);
nand U1164 (N_1164,In_532,In_534);
nor U1165 (N_1165,In_503,In_489);
xor U1166 (N_1166,In_334,In_601);
xor U1167 (N_1167,In_462,In_323);
xor U1168 (N_1168,In_346,In_206);
and U1169 (N_1169,In_784,In_906);
and U1170 (N_1170,In_777,In_612);
or U1171 (N_1171,In_421,In_123);
and U1172 (N_1172,In_499,In_323);
and U1173 (N_1173,In_920,In_953);
or U1174 (N_1174,In_282,In_488);
and U1175 (N_1175,In_624,In_589);
nor U1176 (N_1176,In_988,In_798);
or U1177 (N_1177,In_500,In_58);
xnor U1178 (N_1178,In_96,In_322);
or U1179 (N_1179,In_529,In_775);
or U1180 (N_1180,In_105,In_94);
and U1181 (N_1181,In_184,In_124);
nor U1182 (N_1182,In_338,In_4);
or U1183 (N_1183,In_861,In_157);
nand U1184 (N_1184,In_234,In_838);
or U1185 (N_1185,In_475,In_445);
and U1186 (N_1186,In_61,In_541);
and U1187 (N_1187,In_621,In_168);
xor U1188 (N_1188,In_89,In_786);
nand U1189 (N_1189,In_737,In_356);
nor U1190 (N_1190,In_938,In_688);
nor U1191 (N_1191,In_264,In_935);
nor U1192 (N_1192,In_512,In_727);
or U1193 (N_1193,In_955,In_604);
nor U1194 (N_1194,In_640,In_268);
and U1195 (N_1195,In_945,In_246);
nand U1196 (N_1196,In_849,In_757);
nand U1197 (N_1197,In_14,In_718);
and U1198 (N_1198,In_802,In_180);
or U1199 (N_1199,In_637,In_667);
and U1200 (N_1200,In_423,In_805);
nor U1201 (N_1201,In_106,In_995);
nor U1202 (N_1202,In_974,In_784);
nand U1203 (N_1203,In_575,In_77);
nor U1204 (N_1204,In_382,In_268);
and U1205 (N_1205,In_926,In_807);
nor U1206 (N_1206,In_733,In_26);
nor U1207 (N_1207,In_550,In_857);
nor U1208 (N_1208,In_810,In_321);
nor U1209 (N_1209,In_397,In_446);
or U1210 (N_1210,In_279,In_792);
nand U1211 (N_1211,In_744,In_191);
or U1212 (N_1212,In_803,In_226);
nor U1213 (N_1213,In_44,In_498);
and U1214 (N_1214,In_146,In_531);
nand U1215 (N_1215,In_81,In_489);
nand U1216 (N_1216,In_835,In_402);
and U1217 (N_1217,In_561,In_327);
nand U1218 (N_1218,In_476,In_198);
nor U1219 (N_1219,In_74,In_983);
or U1220 (N_1220,In_393,In_198);
nand U1221 (N_1221,In_656,In_302);
and U1222 (N_1222,In_622,In_9);
nand U1223 (N_1223,In_187,In_802);
or U1224 (N_1224,In_381,In_491);
or U1225 (N_1225,In_911,In_929);
nor U1226 (N_1226,In_196,In_775);
nand U1227 (N_1227,In_447,In_373);
nand U1228 (N_1228,In_585,In_600);
nand U1229 (N_1229,In_175,In_446);
and U1230 (N_1230,In_728,In_211);
and U1231 (N_1231,In_129,In_937);
nand U1232 (N_1232,In_893,In_928);
nor U1233 (N_1233,In_836,In_955);
and U1234 (N_1234,In_799,In_376);
nor U1235 (N_1235,In_554,In_75);
nor U1236 (N_1236,In_606,In_278);
or U1237 (N_1237,In_750,In_462);
and U1238 (N_1238,In_596,In_80);
nand U1239 (N_1239,In_714,In_395);
and U1240 (N_1240,In_849,In_647);
or U1241 (N_1241,In_966,In_897);
or U1242 (N_1242,In_794,In_252);
and U1243 (N_1243,In_560,In_536);
nor U1244 (N_1244,In_33,In_597);
nor U1245 (N_1245,In_28,In_437);
nor U1246 (N_1246,In_807,In_362);
and U1247 (N_1247,In_861,In_181);
nor U1248 (N_1248,In_699,In_663);
or U1249 (N_1249,In_343,In_843);
nor U1250 (N_1250,In_337,In_798);
and U1251 (N_1251,In_696,In_846);
or U1252 (N_1252,In_241,In_653);
or U1253 (N_1253,In_897,In_645);
nand U1254 (N_1254,In_570,In_469);
and U1255 (N_1255,In_587,In_660);
nand U1256 (N_1256,In_833,In_630);
nand U1257 (N_1257,In_677,In_906);
nor U1258 (N_1258,In_140,In_445);
or U1259 (N_1259,In_733,In_477);
nand U1260 (N_1260,In_974,In_669);
nand U1261 (N_1261,In_793,In_903);
and U1262 (N_1262,In_295,In_890);
nand U1263 (N_1263,In_894,In_808);
nand U1264 (N_1264,In_222,In_397);
and U1265 (N_1265,In_211,In_994);
or U1266 (N_1266,In_181,In_436);
nand U1267 (N_1267,In_960,In_211);
nand U1268 (N_1268,In_920,In_2);
nor U1269 (N_1269,In_815,In_173);
and U1270 (N_1270,In_515,In_312);
nand U1271 (N_1271,In_954,In_582);
xor U1272 (N_1272,In_127,In_563);
and U1273 (N_1273,In_97,In_540);
or U1274 (N_1274,In_267,In_706);
and U1275 (N_1275,In_613,In_618);
nor U1276 (N_1276,In_440,In_271);
and U1277 (N_1277,In_358,In_704);
nand U1278 (N_1278,In_567,In_473);
nand U1279 (N_1279,In_68,In_590);
or U1280 (N_1280,In_30,In_605);
nand U1281 (N_1281,In_108,In_204);
or U1282 (N_1282,In_581,In_686);
nand U1283 (N_1283,In_191,In_99);
nand U1284 (N_1284,In_935,In_90);
nor U1285 (N_1285,In_315,In_731);
or U1286 (N_1286,In_108,In_139);
nor U1287 (N_1287,In_510,In_415);
and U1288 (N_1288,In_716,In_913);
and U1289 (N_1289,In_69,In_653);
nand U1290 (N_1290,In_984,In_939);
or U1291 (N_1291,In_705,In_743);
nand U1292 (N_1292,In_520,In_54);
and U1293 (N_1293,In_583,In_429);
nor U1294 (N_1294,In_801,In_629);
nor U1295 (N_1295,In_434,In_381);
and U1296 (N_1296,In_841,In_618);
or U1297 (N_1297,In_123,In_277);
or U1298 (N_1298,In_510,In_371);
or U1299 (N_1299,In_507,In_944);
nor U1300 (N_1300,In_96,In_93);
and U1301 (N_1301,In_773,In_139);
and U1302 (N_1302,In_438,In_741);
nor U1303 (N_1303,In_678,In_953);
or U1304 (N_1304,In_482,In_363);
nor U1305 (N_1305,In_320,In_460);
nor U1306 (N_1306,In_329,In_548);
nor U1307 (N_1307,In_160,In_546);
or U1308 (N_1308,In_83,In_106);
nand U1309 (N_1309,In_252,In_920);
and U1310 (N_1310,In_223,In_344);
or U1311 (N_1311,In_713,In_215);
nor U1312 (N_1312,In_113,In_773);
nand U1313 (N_1313,In_717,In_535);
and U1314 (N_1314,In_240,In_222);
and U1315 (N_1315,In_152,In_633);
nor U1316 (N_1316,In_188,In_61);
nand U1317 (N_1317,In_524,In_602);
or U1318 (N_1318,In_511,In_790);
or U1319 (N_1319,In_186,In_431);
and U1320 (N_1320,In_639,In_35);
and U1321 (N_1321,In_791,In_349);
nand U1322 (N_1322,In_41,In_725);
nor U1323 (N_1323,In_287,In_280);
and U1324 (N_1324,In_679,In_163);
and U1325 (N_1325,In_607,In_549);
nand U1326 (N_1326,In_461,In_498);
or U1327 (N_1327,In_192,In_63);
nor U1328 (N_1328,In_636,In_829);
nand U1329 (N_1329,In_503,In_248);
xnor U1330 (N_1330,In_683,In_384);
or U1331 (N_1331,In_790,In_579);
nand U1332 (N_1332,In_252,In_382);
or U1333 (N_1333,In_506,In_388);
and U1334 (N_1334,In_113,In_973);
nor U1335 (N_1335,In_31,In_432);
nand U1336 (N_1336,In_562,In_31);
and U1337 (N_1337,In_550,In_102);
or U1338 (N_1338,In_221,In_251);
and U1339 (N_1339,In_998,In_198);
nor U1340 (N_1340,In_309,In_603);
nor U1341 (N_1341,In_998,In_324);
nand U1342 (N_1342,In_165,In_438);
and U1343 (N_1343,In_553,In_920);
and U1344 (N_1344,In_201,In_274);
nor U1345 (N_1345,In_131,In_106);
nand U1346 (N_1346,In_252,In_580);
nor U1347 (N_1347,In_682,In_202);
and U1348 (N_1348,In_699,In_261);
and U1349 (N_1349,In_973,In_971);
nand U1350 (N_1350,In_138,In_464);
nor U1351 (N_1351,In_277,In_532);
nor U1352 (N_1352,In_278,In_249);
or U1353 (N_1353,In_582,In_8);
nor U1354 (N_1354,In_419,In_310);
xor U1355 (N_1355,In_615,In_4);
or U1356 (N_1356,In_225,In_733);
nor U1357 (N_1357,In_864,In_887);
and U1358 (N_1358,In_530,In_300);
nand U1359 (N_1359,In_687,In_98);
or U1360 (N_1360,In_644,In_888);
or U1361 (N_1361,In_413,In_162);
and U1362 (N_1362,In_145,In_22);
xnor U1363 (N_1363,In_490,In_175);
and U1364 (N_1364,In_152,In_7);
nand U1365 (N_1365,In_588,In_467);
xnor U1366 (N_1366,In_155,In_768);
nor U1367 (N_1367,In_511,In_58);
nand U1368 (N_1368,In_787,In_120);
nand U1369 (N_1369,In_951,In_416);
or U1370 (N_1370,In_283,In_659);
nor U1371 (N_1371,In_37,In_658);
or U1372 (N_1372,In_12,In_418);
and U1373 (N_1373,In_129,In_740);
or U1374 (N_1374,In_48,In_699);
and U1375 (N_1375,In_0,In_413);
nor U1376 (N_1376,In_852,In_359);
nand U1377 (N_1377,In_894,In_16);
or U1378 (N_1378,In_313,In_836);
or U1379 (N_1379,In_290,In_474);
and U1380 (N_1380,In_519,In_618);
nor U1381 (N_1381,In_638,In_656);
and U1382 (N_1382,In_0,In_961);
nor U1383 (N_1383,In_186,In_463);
or U1384 (N_1384,In_294,In_63);
nand U1385 (N_1385,In_493,In_999);
or U1386 (N_1386,In_167,In_350);
and U1387 (N_1387,In_486,In_158);
and U1388 (N_1388,In_601,In_793);
and U1389 (N_1389,In_756,In_102);
nor U1390 (N_1390,In_871,In_861);
and U1391 (N_1391,In_899,In_48);
or U1392 (N_1392,In_627,In_42);
nand U1393 (N_1393,In_529,In_534);
and U1394 (N_1394,In_339,In_790);
nand U1395 (N_1395,In_984,In_855);
nor U1396 (N_1396,In_336,In_459);
or U1397 (N_1397,In_965,In_101);
or U1398 (N_1398,In_531,In_983);
or U1399 (N_1399,In_102,In_314);
xnor U1400 (N_1400,In_571,In_776);
nand U1401 (N_1401,In_471,In_621);
nand U1402 (N_1402,In_263,In_857);
nor U1403 (N_1403,In_822,In_713);
nor U1404 (N_1404,In_63,In_605);
nand U1405 (N_1405,In_18,In_656);
and U1406 (N_1406,In_107,In_676);
nand U1407 (N_1407,In_823,In_739);
or U1408 (N_1408,In_931,In_488);
nand U1409 (N_1409,In_109,In_385);
nor U1410 (N_1410,In_103,In_794);
nor U1411 (N_1411,In_477,In_752);
and U1412 (N_1412,In_101,In_788);
and U1413 (N_1413,In_182,In_816);
or U1414 (N_1414,In_117,In_133);
or U1415 (N_1415,In_614,In_480);
nand U1416 (N_1416,In_646,In_100);
or U1417 (N_1417,In_87,In_677);
nor U1418 (N_1418,In_28,In_283);
nor U1419 (N_1419,In_211,In_290);
nor U1420 (N_1420,In_697,In_740);
nand U1421 (N_1421,In_63,In_923);
nor U1422 (N_1422,In_134,In_701);
nand U1423 (N_1423,In_352,In_609);
nand U1424 (N_1424,In_247,In_731);
and U1425 (N_1425,In_480,In_741);
xnor U1426 (N_1426,In_950,In_237);
or U1427 (N_1427,In_850,In_371);
nor U1428 (N_1428,In_676,In_545);
nor U1429 (N_1429,In_144,In_433);
and U1430 (N_1430,In_494,In_189);
or U1431 (N_1431,In_323,In_159);
nor U1432 (N_1432,In_215,In_991);
and U1433 (N_1433,In_287,In_697);
nand U1434 (N_1434,In_720,In_886);
nor U1435 (N_1435,In_973,In_237);
or U1436 (N_1436,In_590,In_567);
and U1437 (N_1437,In_598,In_770);
nand U1438 (N_1438,In_525,In_750);
or U1439 (N_1439,In_841,In_536);
nand U1440 (N_1440,In_594,In_855);
nor U1441 (N_1441,In_291,In_294);
nor U1442 (N_1442,In_547,In_287);
or U1443 (N_1443,In_275,In_184);
or U1444 (N_1444,In_806,In_890);
or U1445 (N_1445,In_902,In_464);
nor U1446 (N_1446,In_218,In_448);
or U1447 (N_1447,In_431,In_54);
nand U1448 (N_1448,In_238,In_196);
or U1449 (N_1449,In_68,In_133);
or U1450 (N_1450,In_831,In_866);
and U1451 (N_1451,In_640,In_69);
nand U1452 (N_1452,In_851,In_491);
or U1453 (N_1453,In_736,In_1);
nand U1454 (N_1454,In_58,In_676);
nand U1455 (N_1455,In_907,In_914);
or U1456 (N_1456,In_446,In_363);
nand U1457 (N_1457,In_454,In_393);
and U1458 (N_1458,In_549,In_188);
nand U1459 (N_1459,In_98,In_215);
nand U1460 (N_1460,In_626,In_198);
nand U1461 (N_1461,In_724,In_609);
nor U1462 (N_1462,In_44,In_2);
or U1463 (N_1463,In_552,In_763);
and U1464 (N_1464,In_812,In_169);
nand U1465 (N_1465,In_252,In_110);
and U1466 (N_1466,In_660,In_949);
nand U1467 (N_1467,In_540,In_476);
nor U1468 (N_1468,In_837,In_357);
or U1469 (N_1469,In_294,In_677);
nand U1470 (N_1470,In_949,In_828);
or U1471 (N_1471,In_215,In_231);
nor U1472 (N_1472,In_199,In_180);
and U1473 (N_1473,In_368,In_504);
nand U1474 (N_1474,In_423,In_808);
nor U1475 (N_1475,In_991,In_933);
nor U1476 (N_1476,In_384,In_661);
or U1477 (N_1477,In_374,In_428);
nand U1478 (N_1478,In_773,In_862);
nand U1479 (N_1479,In_56,In_224);
nand U1480 (N_1480,In_800,In_786);
nor U1481 (N_1481,In_486,In_592);
or U1482 (N_1482,In_689,In_545);
or U1483 (N_1483,In_775,In_904);
and U1484 (N_1484,In_853,In_409);
nand U1485 (N_1485,In_772,In_270);
xor U1486 (N_1486,In_150,In_7);
or U1487 (N_1487,In_498,In_285);
nand U1488 (N_1488,In_631,In_682);
nor U1489 (N_1489,In_349,In_121);
or U1490 (N_1490,In_983,In_13);
and U1491 (N_1491,In_643,In_159);
and U1492 (N_1492,In_335,In_321);
and U1493 (N_1493,In_528,In_948);
or U1494 (N_1494,In_479,In_650);
and U1495 (N_1495,In_971,In_532);
nand U1496 (N_1496,In_134,In_413);
nand U1497 (N_1497,In_386,In_938);
and U1498 (N_1498,In_588,In_51);
nand U1499 (N_1499,In_388,In_276);
and U1500 (N_1500,In_125,In_818);
or U1501 (N_1501,In_138,In_714);
or U1502 (N_1502,In_64,In_989);
nor U1503 (N_1503,In_203,In_172);
or U1504 (N_1504,In_630,In_102);
or U1505 (N_1505,In_148,In_519);
or U1506 (N_1506,In_840,In_296);
nor U1507 (N_1507,In_658,In_846);
or U1508 (N_1508,In_132,In_475);
nand U1509 (N_1509,In_210,In_814);
nor U1510 (N_1510,In_812,In_318);
nand U1511 (N_1511,In_133,In_551);
and U1512 (N_1512,In_611,In_300);
nor U1513 (N_1513,In_678,In_186);
nor U1514 (N_1514,In_316,In_37);
and U1515 (N_1515,In_795,In_952);
nor U1516 (N_1516,In_910,In_839);
nand U1517 (N_1517,In_240,In_820);
and U1518 (N_1518,In_576,In_134);
nor U1519 (N_1519,In_982,In_667);
nand U1520 (N_1520,In_665,In_731);
or U1521 (N_1521,In_36,In_569);
and U1522 (N_1522,In_452,In_8);
nor U1523 (N_1523,In_369,In_401);
nor U1524 (N_1524,In_747,In_195);
and U1525 (N_1525,In_270,In_837);
or U1526 (N_1526,In_970,In_60);
nor U1527 (N_1527,In_867,In_657);
and U1528 (N_1528,In_399,In_191);
or U1529 (N_1529,In_65,In_837);
nand U1530 (N_1530,In_843,In_652);
and U1531 (N_1531,In_256,In_173);
nand U1532 (N_1532,In_488,In_555);
nor U1533 (N_1533,In_501,In_132);
or U1534 (N_1534,In_179,In_47);
or U1535 (N_1535,In_668,In_620);
and U1536 (N_1536,In_902,In_452);
nand U1537 (N_1537,In_475,In_576);
nor U1538 (N_1538,In_171,In_571);
and U1539 (N_1539,In_196,In_169);
nand U1540 (N_1540,In_559,In_733);
nor U1541 (N_1541,In_923,In_825);
nand U1542 (N_1542,In_94,In_114);
nand U1543 (N_1543,In_449,In_72);
nand U1544 (N_1544,In_569,In_16);
or U1545 (N_1545,In_694,In_823);
nand U1546 (N_1546,In_573,In_771);
and U1547 (N_1547,In_671,In_80);
nand U1548 (N_1548,In_348,In_264);
nand U1549 (N_1549,In_325,In_965);
or U1550 (N_1550,In_259,In_276);
nand U1551 (N_1551,In_506,In_234);
or U1552 (N_1552,In_724,In_338);
or U1553 (N_1553,In_965,In_517);
nand U1554 (N_1554,In_553,In_832);
and U1555 (N_1555,In_728,In_267);
nor U1556 (N_1556,In_730,In_713);
nor U1557 (N_1557,In_473,In_895);
or U1558 (N_1558,In_529,In_31);
nand U1559 (N_1559,In_528,In_911);
or U1560 (N_1560,In_513,In_783);
or U1561 (N_1561,In_766,In_866);
nor U1562 (N_1562,In_368,In_297);
or U1563 (N_1563,In_508,In_53);
nor U1564 (N_1564,In_444,In_799);
nand U1565 (N_1565,In_179,In_544);
and U1566 (N_1566,In_25,In_257);
xnor U1567 (N_1567,In_981,In_681);
and U1568 (N_1568,In_105,In_753);
nor U1569 (N_1569,In_593,In_2);
and U1570 (N_1570,In_463,In_265);
and U1571 (N_1571,In_771,In_438);
or U1572 (N_1572,In_56,In_145);
and U1573 (N_1573,In_975,In_113);
nor U1574 (N_1574,In_562,In_192);
or U1575 (N_1575,In_628,In_487);
nand U1576 (N_1576,In_463,In_736);
or U1577 (N_1577,In_452,In_335);
and U1578 (N_1578,In_673,In_128);
nand U1579 (N_1579,In_671,In_444);
or U1580 (N_1580,In_203,In_490);
or U1581 (N_1581,In_347,In_715);
nand U1582 (N_1582,In_403,In_539);
xnor U1583 (N_1583,In_860,In_111);
nand U1584 (N_1584,In_34,In_38);
nand U1585 (N_1585,In_721,In_430);
and U1586 (N_1586,In_660,In_30);
or U1587 (N_1587,In_907,In_367);
and U1588 (N_1588,In_910,In_334);
or U1589 (N_1589,In_401,In_863);
nor U1590 (N_1590,In_340,In_503);
and U1591 (N_1591,In_136,In_197);
nand U1592 (N_1592,In_279,In_305);
and U1593 (N_1593,In_436,In_442);
and U1594 (N_1594,In_472,In_763);
and U1595 (N_1595,In_905,In_449);
nor U1596 (N_1596,In_678,In_654);
and U1597 (N_1597,In_568,In_818);
or U1598 (N_1598,In_272,In_278);
nor U1599 (N_1599,In_778,In_917);
or U1600 (N_1600,In_522,In_426);
or U1601 (N_1601,In_124,In_598);
or U1602 (N_1602,In_986,In_195);
nor U1603 (N_1603,In_35,In_829);
nor U1604 (N_1604,In_943,In_5);
and U1605 (N_1605,In_108,In_474);
nand U1606 (N_1606,In_28,In_150);
or U1607 (N_1607,In_800,In_578);
and U1608 (N_1608,In_256,In_195);
or U1609 (N_1609,In_396,In_176);
xnor U1610 (N_1610,In_395,In_710);
or U1611 (N_1611,In_816,In_135);
nand U1612 (N_1612,In_914,In_922);
and U1613 (N_1613,In_815,In_571);
nand U1614 (N_1614,In_745,In_416);
nor U1615 (N_1615,In_984,In_768);
and U1616 (N_1616,In_418,In_338);
nand U1617 (N_1617,In_945,In_48);
nor U1618 (N_1618,In_400,In_634);
or U1619 (N_1619,In_212,In_912);
nand U1620 (N_1620,In_237,In_734);
nand U1621 (N_1621,In_183,In_909);
nand U1622 (N_1622,In_520,In_28);
and U1623 (N_1623,In_215,In_635);
nand U1624 (N_1624,In_286,In_539);
or U1625 (N_1625,In_120,In_319);
or U1626 (N_1626,In_51,In_185);
or U1627 (N_1627,In_642,In_112);
or U1628 (N_1628,In_573,In_522);
and U1629 (N_1629,In_694,In_798);
nor U1630 (N_1630,In_914,In_305);
or U1631 (N_1631,In_799,In_94);
nor U1632 (N_1632,In_359,In_683);
nor U1633 (N_1633,In_235,In_747);
nor U1634 (N_1634,In_562,In_913);
and U1635 (N_1635,In_439,In_645);
nand U1636 (N_1636,In_316,In_938);
nor U1637 (N_1637,In_751,In_965);
nor U1638 (N_1638,In_389,In_17);
and U1639 (N_1639,In_174,In_655);
nand U1640 (N_1640,In_275,In_181);
and U1641 (N_1641,In_921,In_493);
nor U1642 (N_1642,In_47,In_428);
nand U1643 (N_1643,In_922,In_307);
nor U1644 (N_1644,In_595,In_192);
and U1645 (N_1645,In_80,In_763);
or U1646 (N_1646,In_668,In_204);
nor U1647 (N_1647,In_771,In_777);
or U1648 (N_1648,In_887,In_607);
nand U1649 (N_1649,In_21,In_566);
or U1650 (N_1650,In_486,In_344);
nor U1651 (N_1651,In_776,In_21);
or U1652 (N_1652,In_968,In_365);
nand U1653 (N_1653,In_974,In_61);
nand U1654 (N_1654,In_897,In_71);
nand U1655 (N_1655,In_158,In_210);
and U1656 (N_1656,In_713,In_842);
or U1657 (N_1657,In_628,In_723);
nor U1658 (N_1658,In_520,In_934);
nand U1659 (N_1659,In_109,In_101);
and U1660 (N_1660,In_470,In_222);
nand U1661 (N_1661,In_746,In_469);
or U1662 (N_1662,In_347,In_304);
nor U1663 (N_1663,In_410,In_213);
nor U1664 (N_1664,In_454,In_120);
nor U1665 (N_1665,In_889,In_310);
nor U1666 (N_1666,In_308,In_996);
nor U1667 (N_1667,In_110,In_441);
or U1668 (N_1668,In_675,In_632);
nor U1669 (N_1669,In_4,In_473);
nand U1670 (N_1670,In_665,In_411);
nand U1671 (N_1671,In_846,In_432);
nor U1672 (N_1672,In_845,In_252);
nor U1673 (N_1673,In_757,In_121);
nand U1674 (N_1674,In_218,In_320);
nand U1675 (N_1675,In_105,In_893);
and U1676 (N_1676,In_224,In_497);
nand U1677 (N_1677,In_556,In_859);
and U1678 (N_1678,In_539,In_778);
nor U1679 (N_1679,In_253,In_849);
nand U1680 (N_1680,In_133,In_257);
nand U1681 (N_1681,In_191,In_777);
nor U1682 (N_1682,In_588,In_101);
or U1683 (N_1683,In_746,In_489);
nor U1684 (N_1684,In_218,In_659);
nor U1685 (N_1685,In_515,In_859);
or U1686 (N_1686,In_858,In_678);
nor U1687 (N_1687,In_269,In_838);
or U1688 (N_1688,In_527,In_106);
nor U1689 (N_1689,In_145,In_733);
and U1690 (N_1690,In_566,In_386);
nor U1691 (N_1691,In_117,In_252);
and U1692 (N_1692,In_93,In_8);
nor U1693 (N_1693,In_693,In_680);
nand U1694 (N_1694,In_212,In_831);
nor U1695 (N_1695,In_531,In_65);
nor U1696 (N_1696,In_223,In_561);
nor U1697 (N_1697,In_989,In_495);
nor U1698 (N_1698,In_950,In_607);
nand U1699 (N_1699,In_812,In_396);
or U1700 (N_1700,In_248,In_372);
nor U1701 (N_1701,In_436,In_103);
xor U1702 (N_1702,In_55,In_50);
nand U1703 (N_1703,In_699,In_633);
and U1704 (N_1704,In_641,In_680);
or U1705 (N_1705,In_415,In_118);
or U1706 (N_1706,In_64,In_226);
and U1707 (N_1707,In_379,In_101);
nand U1708 (N_1708,In_845,In_902);
nor U1709 (N_1709,In_992,In_558);
nand U1710 (N_1710,In_797,In_341);
nor U1711 (N_1711,In_950,In_584);
nor U1712 (N_1712,In_910,In_918);
nand U1713 (N_1713,In_412,In_253);
and U1714 (N_1714,In_81,In_799);
nor U1715 (N_1715,In_639,In_693);
or U1716 (N_1716,In_250,In_425);
nor U1717 (N_1717,In_612,In_649);
nor U1718 (N_1718,In_137,In_620);
nand U1719 (N_1719,In_668,In_842);
or U1720 (N_1720,In_582,In_39);
or U1721 (N_1721,In_214,In_980);
or U1722 (N_1722,In_63,In_186);
and U1723 (N_1723,In_508,In_842);
nor U1724 (N_1724,In_827,In_925);
nor U1725 (N_1725,In_282,In_294);
or U1726 (N_1726,In_257,In_249);
nor U1727 (N_1727,In_774,In_184);
xnor U1728 (N_1728,In_246,In_404);
or U1729 (N_1729,In_604,In_935);
nor U1730 (N_1730,In_514,In_782);
nand U1731 (N_1731,In_37,In_326);
nand U1732 (N_1732,In_512,In_112);
or U1733 (N_1733,In_518,In_631);
and U1734 (N_1734,In_681,In_42);
nand U1735 (N_1735,In_634,In_893);
and U1736 (N_1736,In_758,In_457);
nor U1737 (N_1737,In_779,In_168);
nand U1738 (N_1738,In_578,In_154);
and U1739 (N_1739,In_607,In_297);
and U1740 (N_1740,In_305,In_598);
nor U1741 (N_1741,In_676,In_236);
xor U1742 (N_1742,In_65,In_867);
nand U1743 (N_1743,In_96,In_532);
nand U1744 (N_1744,In_621,In_710);
nor U1745 (N_1745,In_293,In_503);
or U1746 (N_1746,In_179,In_699);
nand U1747 (N_1747,In_200,In_636);
and U1748 (N_1748,In_904,In_932);
nor U1749 (N_1749,In_44,In_290);
nor U1750 (N_1750,In_531,In_984);
and U1751 (N_1751,In_592,In_695);
or U1752 (N_1752,In_466,In_113);
nor U1753 (N_1753,In_36,In_719);
and U1754 (N_1754,In_860,In_113);
and U1755 (N_1755,In_779,In_264);
nor U1756 (N_1756,In_94,In_954);
nand U1757 (N_1757,In_717,In_396);
nor U1758 (N_1758,In_29,In_858);
nor U1759 (N_1759,In_791,In_501);
or U1760 (N_1760,In_381,In_812);
nor U1761 (N_1761,In_574,In_423);
nor U1762 (N_1762,In_236,In_408);
nand U1763 (N_1763,In_851,In_382);
nor U1764 (N_1764,In_935,In_17);
and U1765 (N_1765,In_633,In_775);
nor U1766 (N_1766,In_914,In_150);
nand U1767 (N_1767,In_168,In_173);
or U1768 (N_1768,In_70,In_78);
nor U1769 (N_1769,In_980,In_404);
or U1770 (N_1770,In_41,In_384);
and U1771 (N_1771,In_437,In_129);
or U1772 (N_1772,In_802,In_937);
and U1773 (N_1773,In_21,In_345);
nand U1774 (N_1774,In_8,In_435);
nand U1775 (N_1775,In_35,In_452);
nand U1776 (N_1776,In_838,In_220);
or U1777 (N_1777,In_890,In_840);
nand U1778 (N_1778,In_746,In_327);
or U1779 (N_1779,In_533,In_981);
nor U1780 (N_1780,In_298,In_521);
nor U1781 (N_1781,In_398,In_759);
nor U1782 (N_1782,In_64,In_918);
or U1783 (N_1783,In_133,In_849);
nand U1784 (N_1784,In_553,In_829);
and U1785 (N_1785,In_405,In_81);
or U1786 (N_1786,In_671,In_650);
or U1787 (N_1787,In_764,In_677);
or U1788 (N_1788,In_328,In_238);
and U1789 (N_1789,In_814,In_661);
nand U1790 (N_1790,In_333,In_841);
nor U1791 (N_1791,In_698,In_658);
nor U1792 (N_1792,In_976,In_620);
nor U1793 (N_1793,In_466,In_778);
or U1794 (N_1794,In_890,In_176);
xor U1795 (N_1795,In_739,In_231);
nor U1796 (N_1796,In_999,In_86);
nor U1797 (N_1797,In_995,In_412);
xnor U1798 (N_1798,In_362,In_977);
or U1799 (N_1799,In_861,In_822);
nand U1800 (N_1800,In_734,In_369);
nor U1801 (N_1801,In_582,In_703);
nand U1802 (N_1802,In_596,In_493);
nor U1803 (N_1803,In_187,In_96);
or U1804 (N_1804,In_197,In_780);
nand U1805 (N_1805,In_40,In_38);
and U1806 (N_1806,In_87,In_953);
or U1807 (N_1807,In_465,In_733);
or U1808 (N_1808,In_560,In_978);
and U1809 (N_1809,In_859,In_630);
nor U1810 (N_1810,In_548,In_689);
nor U1811 (N_1811,In_217,In_268);
nor U1812 (N_1812,In_951,In_696);
nand U1813 (N_1813,In_2,In_321);
and U1814 (N_1814,In_201,In_640);
xor U1815 (N_1815,In_268,In_978);
and U1816 (N_1816,In_89,In_553);
and U1817 (N_1817,In_542,In_290);
and U1818 (N_1818,In_493,In_307);
and U1819 (N_1819,In_800,In_908);
or U1820 (N_1820,In_526,In_122);
and U1821 (N_1821,In_743,In_926);
nand U1822 (N_1822,In_356,In_905);
or U1823 (N_1823,In_14,In_526);
and U1824 (N_1824,In_162,In_745);
nor U1825 (N_1825,In_215,In_327);
and U1826 (N_1826,In_180,In_54);
nand U1827 (N_1827,In_213,In_857);
and U1828 (N_1828,In_816,In_103);
or U1829 (N_1829,In_351,In_286);
nand U1830 (N_1830,In_336,In_641);
nor U1831 (N_1831,In_86,In_109);
nand U1832 (N_1832,In_213,In_733);
and U1833 (N_1833,In_734,In_857);
or U1834 (N_1834,In_596,In_757);
or U1835 (N_1835,In_721,In_775);
nor U1836 (N_1836,In_150,In_262);
and U1837 (N_1837,In_467,In_52);
or U1838 (N_1838,In_82,In_877);
nor U1839 (N_1839,In_576,In_371);
or U1840 (N_1840,In_118,In_807);
or U1841 (N_1841,In_606,In_520);
nand U1842 (N_1842,In_802,In_437);
and U1843 (N_1843,In_317,In_401);
nand U1844 (N_1844,In_617,In_885);
nand U1845 (N_1845,In_349,In_630);
nor U1846 (N_1846,In_343,In_173);
or U1847 (N_1847,In_978,In_791);
nand U1848 (N_1848,In_466,In_323);
or U1849 (N_1849,In_719,In_38);
or U1850 (N_1850,In_668,In_232);
nor U1851 (N_1851,In_236,In_506);
nand U1852 (N_1852,In_906,In_742);
nor U1853 (N_1853,In_195,In_662);
or U1854 (N_1854,In_775,In_739);
nand U1855 (N_1855,In_495,In_678);
and U1856 (N_1856,In_563,In_637);
nand U1857 (N_1857,In_77,In_524);
nand U1858 (N_1858,In_900,In_47);
nor U1859 (N_1859,In_133,In_766);
nor U1860 (N_1860,In_122,In_564);
and U1861 (N_1861,In_207,In_741);
and U1862 (N_1862,In_408,In_275);
and U1863 (N_1863,In_716,In_284);
nor U1864 (N_1864,In_237,In_357);
nor U1865 (N_1865,In_317,In_261);
nand U1866 (N_1866,In_727,In_199);
and U1867 (N_1867,In_209,In_726);
and U1868 (N_1868,In_729,In_706);
nand U1869 (N_1869,In_491,In_126);
and U1870 (N_1870,In_159,In_51);
or U1871 (N_1871,In_434,In_795);
nor U1872 (N_1872,In_63,In_534);
and U1873 (N_1873,In_100,In_573);
nand U1874 (N_1874,In_162,In_62);
and U1875 (N_1875,In_464,In_784);
and U1876 (N_1876,In_356,In_442);
and U1877 (N_1877,In_156,In_974);
or U1878 (N_1878,In_661,In_236);
nand U1879 (N_1879,In_647,In_815);
or U1880 (N_1880,In_66,In_251);
and U1881 (N_1881,In_979,In_836);
and U1882 (N_1882,In_347,In_230);
and U1883 (N_1883,In_174,In_66);
nor U1884 (N_1884,In_465,In_977);
or U1885 (N_1885,In_17,In_242);
and U1886 (N_1886,In_27,In_605);
nor U1887 (N_1887,In_601,In_176);
nand U1888 (N_1888,In_848,In_195);
nor U1889 (N_1889,In_40,In_39);
nand U1890 (N_1890,In_489,In_353);
and U1891 (N_1891,In_203,In_752);
nor U1892 (N_1892,In_768,In_894);
nor U1893 (N_1893,In_22,In_866);
nand U1894 (N_1894,In_335,In_928);
xnor U1895 (N_1895,In_200,In_902);
and U1896 (N_1896,In_933,In_926);
or U1897 (N_1897,In_14,In_469);
nand U1898 (N_1898,In_199,In_702);
nand U1899 (N_1899,In_610,In_643);
and U1900 (N_1900,In_868,In_290);
or U1901 (N_1901,In_718,In_118);
and U1902 (N_1902,In_819,In_920);
or U1903 (N_1903,In_472,In_79);
and U1904 (N_1904,In_237,In_985);
nor U1905 (N_1905,In_678,In_512);
and U1906 (N_1906,In_971,In_167);
nor U1907 (N_1907,In_246,In_356);
and U1908 (N_1908,In_747,In_139);
or U1909 (N_1909,In_720,In_184);
nand U1910 (N_1910,In_11,In_453);
or U1911 (N_1911,In_135,In_966);
xnor U1912 (N_1912,In_731,In_79);
nand U1913 (N_1913,In_473,In_507);
nor U1914 (N_1914,In_642,In_700);
and U1915 (N_1915,In_311,In_290);
or U1916 (N_1916,In_608,In_199);
or U1917 (N_1917,In_332,In_894);
and U1918 (N_1918,In_28,In_763);
or U1919 (N_1919,In_471,In_45);
nor U1920 (N_1920,In_241,In_371);
or U1921 (N_1921,In_457,In_807);
nand U1922 (N_1922,In_70,In_8);
or U1923 (N_1923,In_280,In_249);
or U1924 (N_1924,In_671,In_54);
nand U1925 (N_1925,In_280,In_260);
nand U1926 (N_1926,In_781,In_48);
nor U1927 (N_1927,In_197,In_347);
and U1928 (N_1928,In_190,In_875);
and U1929 (N_1929,In_487,In_262);
or U1930 (N_1930,In_432,In_143);
or U1931 (N_1931,In_881,In_555);
or U1932 (N_1932,In_977,In_592);
or U1933 (N_1933,In_296,In_767);
or U1934 (N_1934,In_463,In_412);
or U1935 (N_1935,In_736,In_147);
or U1936 (N_1936,In_760,In_700);
or U1937 (N_1937,In_383,In_260);
nor U1938 (N_1938,In_357,In_718);
or U1939 (N_1939,In_763,In_98);
and U1940 (N_1940,In_117,In_866);
or U1941 (N_1941,In_331,In_779);
and U1942 (N_1942,In_313,In_35);
nand U1943 (N_1943,In_625,In_914);
nand U1944 (N_1944,In_250,In_529);
nand U1945 (N_1945,In_192,In_83);
nor U1946 (N_1946,In_306,In_870);
nor U1947 (N_1947,In_671,In_777);
and U1948 (N_1948,In_433,In_400);
and U1949 (N_1949,In_821,In_809);
and U1950 (N_1950,In_186,In_209);
and U1951 (N_1951,In_509,In_235);
and U1952 (N_1952,In_948,In_90);
nand U1953 (N_1953,In_721,In_106);
or U1954 (N_1954,In_184,In_174);
nand U1955 (N_1955,In_274,In_845);
nand U1956 (N_1956,In_957,In_817);
nand U1957 (N_1957,In_621,In_501);
nor U1958 (N_1958,In_826,In_346);
or U1959 (N_1959,In_770,In_528);
and U1960 (N_1960,In_353,In_838);
and U1961 (N_1961,In_712,In_312);
nor U1962 (N_1962,In_498,In_473);
and U1963 (N_1963,In_572,In_75);
or U1964 (N_1964,In_787,In_348);
nor U1965 (N_1965,In_144,In_219);
or U1966 (N_1966,In_566,In_841);
and U1967 (N_1967,In_508,In_414);
nand U1968 (N_1968,In_252,In_60);
or U1969 (N_1969,In_202,In_877);
nand U1970 (N_1970,In_945,In_50);
or U1971 (N_1971,In_887,In_348);
and U1972 (N_1972,In_94,In_865);
or U1973 (N_1973,In_85,In_131);
or U1974 (N_1974,In_230,In_248);
or U1975 (N_1975,In_999,In_49);
nor U1976 (N_1976,In_997,In_204);
and U1977 (N_1977,In_988,In_452);
and U1978 (N_1978,In_316,In_812);
or U1979 (N_1979,In_514,In_121);
nor U1980 (N_1980,In_473,In_739);
nor U1981 (N_1981,In_190,In_735);
and U1982 (N_1982,In_546,In_750);
nor U1983 (N_1983,In_432,In_6);
and U1984 (N_1984,In_169,In_604);
nand U1985 (N_1985,In_862,In_189);
nor U1986 (N_1986,In_912,In_704);
nand U1987 (N_1987,In_87,In_560);
nand U1988 (N_1988,In_314,In_356);
and U1989 (N_1989,In_966,In_541);
or U1990 (N_1990,In_461,In_32);
and U1991 (N_1991,In_888,In_294);
nand U1992 (N_1992,In_953,In_742);
nor U1993 (N_1993,In_284,In_517);
and U1994 (N_1994,In_342,In_733);
nor U1995 (N_1995,In_929,In_316);
or U1996 (N_1996,In_281,In_959);
or U1997 (N_1997,In_68,In_382);
nand U1998 (N_1998,In_165,In_246);
or U1999 (N_1999,In_850,In_438);
or U2000 (N_2000,N_1821,N_701);
or U2001 (N_2001,N_1596,N_716);
and U2002 (N_2002,N_1523,N_837);
nand U2003 (N_2003,N_897,N_1293);
nand U2004 (N_2004,N_900,N_936);
and U2005 (N_2005,N_1489,N_46);
and U2006 (N_2006,N_1996,N_221);
nand U2007 (N_2007,N_1599,N_780);
nor U2008 (N_2008,N_770,N_1133);
or U2009 (N_2009,N_1723,N_1294);
nand U2010 (N_2010,N_1032,N_1078);
and U2011 (N_2011,N_1319,N_652);
nor U2012 (N_2012,N_1412,N_366);
nor U2013 (N_2013,N_140,N_1810);
nor U2014 (N_2014,N_1154,N_857);
nor U2015 (N_2015,N_767,N_563);
and U2016 (N_2016,N_487,N_269);
and U2017 (N_2017,N_683,N_1746);
or U2018 (N_2018,N_441,N_911);
nor U2019 (N_2019,N_1117,N_427);
and U2020 (N_2020,N_385,N_822);
nor U2021 (N_2021,N_1218,N_455);
nand U2022 (N_2022,N_242,N_84);
nand U2023 (N_2023,N_821,N_1661);
nor U2024 (N_2024,N_1334,N_682);
nor U2025 (N_2025,N_160,N_1505);
or U2026 (N_2026,N_1688,N_456);
nand U2027 (N_2027,N_162,N_1056);
nor U2028 (N_2028,N_729,N_1331);
or U2029 (N_2029,N_592,N_1935);
nor U2030 (N_2030,N_641,N_1561);
and U2031 (N_2031,N_539,N_1135);
nand U2032 (N_2032,N_352,N_331);
and U2033 (N_2033,N_1955,N_1683);
nand U2034 (N_2034,N_1610,N_89);
nand U2035 (N_2035,N_1164,N_940);
or U2036 (N_2036,N_259,N_1534);
and U2037 (N_2037,N_1809,N_387);
nand U2038 (N_2038,N_1350,N_1073);
and U2039 (N_2039,N_967,N_847);
nor U2040 (N_2040,N_1354,N_58);
or U2041 (N_2041,N_1196,N_396);
nand U2042 (N_2042,N_884,N_1497);
or U2043 (N_2043,N_1581,N_1721);
and U2044 (N_2044,N_856,N_1283);
nand U2045 (N_2045,N_1738,N_1123);
or U2046 (N_2046,N_1940,N_406);
and U2047 (N_2047,N_1081,N_71);
nor U2048 (N_2048,N_654,N_535);
and U2049 (N_2049,N_1941,N_1703);
or U2050 (N_2050,N_42,N_350);
and U2051 (N_2051,N_1097,N_1043);
and U2052 (N_2052,N_1051,N_1156);
and U2053 (N_2053,N_1298,N_183);
nor U2054 (N_2054,N_1911,N_1920);
nor U2055 (N_2055,N_194,N_1449);
and U2056 (N_2056,N_1875,N_1595);
and U2057 (N_2057,N_308,N_19);
and U2058 (N_2058,N_1593,N_1263);
nand U2059 (N_2059,N_843,N_393);
nand U2060 (N_2060,N_964,N_252);
or U2061 (N_2061,N_2,N_1453);
and U2062 (N_2062,N_943,N_1671);
or U2063 (N_2063,N_1356,N_171);
and U2064 (N_2064,N_1716,N_772);
and U2065 (N_2065,N_626,N_31);
or U2066 (N_2066,N_1153,N_203);
and U2067 (N_2067,N_343,N_391);
nand U2068 (N_2068,N_184,N_414);
nand U2069 (N_2069,N_929,N_286);
and U2070 (N_2070,N_1631,N_779);
nor U2071 (N_2071,N_653,N_694);
and U2072 (N_2072,N_1847,N_1734);
nor U2073 (N_2073,N_738,N_1706);
or U2074 (N_2074,N_1205,N_25);
nor U2075 (N_2075,N_714,N_1909);
and U2076 (N_2076,N_602,N_1332);
nand U2077 (N_2077,N_833,N_1029);
nand U2078 (N_2078,N_933,N_1646);
or U2079 (N_2079,N_1256,N_99);
and U2080 (N_2080,N_679,N_497);
nand U2081 (N_2081,N_1755,N_135);
or U2082 (N_2082,N_556,N_1403);
nand U2083 (N_2083,N_390,N_1514);
nand U2084 (N_2084,N_1336,N_1907);
nor U2085 (N_2085,N_672,N_846);
nor U2086 (N_2086,N_1675,N_506);
and U2087 (N_2087,N_154,N_1789);
and U2088 (N_2088,N_1513,N_789);
nand U2089 (N_2089,N_1377,N_1537);
or U2090 (N_2090,N_462,N_1613);
or U2091 (N_2091,N_1224,N_483);
nand U2092 (N_2092,N_213,N_1428);
nand U2093 (N_2093,N_1750,N_1922);
and U2094 (N_2094,N_1348,N_570);
nand U2095 (N_2095,N_1694,N_1228);
nor U2096 (N_2096,N_1141,N_659);
or U2097 (N_2097,N_647,N_1724);
or U2098 (N_2098,N_1492,N_1677);
nand U2099 (N_2099,N_1673,N_1035);
nand U2100 (N_2100,N_1109,N_1824);
or U2101 (N_2101,N_944,N_945);
and U2102 (N_2102,N_394,N_293);
nor U2103 (N_2103,N_412,N_1021);
and U2104 (N_2104,N_1460,N_1663);
xnor U2105 (N_2105,N_155,N_1507);
or U2106 (N_2106,N_485,N_1147);
or U2107 (N_2107,N_1020,N_56);
and U2108 (N_2108,N_256,N_810);
nor U2109 (N_2109,N_1499,N_577);
and U2110 (N_2110,N_158,N_1279);
and U2111 (N_2111,N_1767,N_176);
nand U2112 (N_2112,N_829,N_1168);
nor U2113 (N_2113,N_783,N_1188);
or U2114 (N_2114,N_587,N_1577);
nor U2115 (N_2115,N_369,N_1680);
and U2116 (N_2116,N_284,N_748);
and U2117 (N_2117,N_877,N_955);
nor U2118 (N_2118,N_1430,N_640);
nor U2119 (N_2119,N_54,N_488);
nand U2120 (N_2120,N_410,N_208);
and U2121 (N_2121,N_1819,N_36);
nor U2122 (N_2122,N_334,N_1938);
nor U2123 (N_2123,N_1504,N_190);
or U2124 (N_2124,N_1914,N_823);
and U2125 (N_2125,N_1540,N_1668);
and U2126 (N_2126,N_1539,N_1089);
nand U2127 (N_2127,N_1899,N_472);
or U2128 (N_2128,N_85,N_1628);
nor U2129 (N_2129,N_1187,N_1547);
and U2130 (N_2130,N_1270,N_782);
nor U2131 (N_2131,N_1562,N_542);
and U2132 (N_2132,N_1729,N_1211);
nor U2133 (N_2133,N_508,N_496);
nor U2134 (N_2134,N_603,N_55);
nor U2135 (N_2135,N_1709,N_612);
and U2136 (N_2136,N_826,N_601);
nor U2137 (N_2137,N_188,N_1818);
nor U2138 (N_2138,N_997,N_711);
and U2139 (N_2139,N_1696,N_606);
nor U2140 (N_2140,N_841,N_1500);
or U2141 (N_2141,N_1896,N_1115);
and U2142 (N_2142,N_1287,N_962);
nor U2143 (N_2143,N_632,N_17);
and U2144 (N_2144,N_367,N_1185);
nand U2145 (N_2145,N_1169,N_1972);
and U2146 (N_2146,N_769,N_1225);
nand U2147 (N_2147,N_594,N_1793);
and U2148 (N_2148,N_887,N_1018);
nor U2149 (N_2149,N_1731,N_149);
and U2150 (N_2150,N_105,N_1385);
nand U2151 (N_2151,N_909,N_1105);
nor U2152 (N_2152,N_1095,N_1085);
nor U2153 (N_2153,N_635,N_1766);
nand U2154 (N_2154,N_1083,N_1607);
nand U2155 (N_2155,N_457,N_625);
or U2156 (N_2156,N_72,N_1233);
and U2157 (N_2157,N_1364,N_187);
nor U2158 (N_2158,N_432,N_1897);
nand U2159 (N_2159,N_377,N_1191);
and U2160 (N_2160,N_442,N_464);
or U2161 (N_2161,N_177,N_420);
nor U2162 (N_2162,N_531,N_801);
or U2163 (N_2163,N_1835,N_81);
nand U2164 (N_2164,N_102,N_23);
or U2165 (N_2165,N_1958,N_294);
nor U2166 (N_2166,N_1984,N_82);
nor U2167 (N_2167,N_623,N_673);
nor U2168 (N_2168,N_808,N_1691);
nor U2169 (N_2169,N_1657,N_167);
nand U2170 (N_2170,N_16,N_1199);
and U2171 (N_2171,N_709,N_802);
and U2172 (N_2172,N_1266,N_1867);
or U2173 (N_2173,N_972,N_1892);
nor U2174 (N_2174,N_1010,N_1009);
and U2175 (N_2175,N_584,N_797);
nand U2176 (N_2176,N_565,N_831);
nand U2177 (N_2177,N_206,N_1606);
nor U2178 (N_2178,N_600,N_317);
and U2179 (N_2179,N_1921,N_1391);
nor U2180 (N_2180,N_1349,N_1623);
or U2181 (N_2181,N_1383,N_251);
nor U2182 (N_2182,N_411,N_675);
nand U2183 (N_2183,N_958,N_232);
nor U2184 (N_2184,N_969,N_798);
and U2185 (N_2185,N_1868,N_210);
nand U2186 (N_2186,N_69,N_1936);
and U2187 (N_2187,N_1061,N_216);
or U2188 (N_2188,N_297,N_1007);
and U2189 (N_2189,N_1652,N_1495);
and U2190 (N_2190,N_671,N_1717);
nand U2191 (N_2191,N_1245,N_796);
nand U2192 (N_2192,N_910,N_1327);
nor U2193 (N_2193,N_419,N_1980);
nand U2194 (N_2194,N_1212,N_1380);
nor U2195 (N_2195,N_114,N_503);
nor U2196 (N_2196,N_871,N_460);
or U2197 (N_2197,N_795,N_908);
and U2198 (N_2198,N_749,N_746);
and U2199 (N_2199,N_120,N_1856);
nand U2200 (N_2200,N_1017,N_392);
xor U2201 (N_2201,N_8,N_1172);
or U2202 (N_2202,N_665,N_1440);
nand U2203 (N_2203,N_1590,N_752);
nor U2204 (N_2204,N_916,N_708);
and U2205 (N_2205,N_1536,N_163);
nor U2206 (N_2206,N_1956,N_1857);
and U2207 (N_2207,N_480,N_1137);
and U2208 (N_2208,N_1288,N_1530);
and U2209 (N_2209,N_121,N_7);
nor U2210 (N_2210,N_1426,N_1291);
or U2211 (N_2211,N_863,N_33);
and U2212 (N_2212,N_1761,N_97);
nand U2213 (N_2213,N_1758,N_1392);
or U2214 (N_2214,N_1929,N_1297);
nor U2215 (N_2215,N_1842,N_262);
xnor U2216 (N_2216,N_1053,N_1047);
or U2217 (N_2217,N_1257,N_759);
nand U2218 (N_2218,N_930,N_0);
nor U2219 (N_2219,N_1062,N_891);
nand U2220 (N_2220,N_1214,N_1076);
nand U2221 (N_2221,N_1252,N_1796);
or U2222 (N_2222,N_1317,N_77);
and U2223 (N_2223,N_549,N_1054);
or U2224 (N_2224,N_270,N_15);
nor U2225 (N_2225,N_960,N_47);
or U2226 (N_2226,N_1075,N_133);
nor U2227 (N_2227,N_1894,N_59);
nand U2228 (N_2228,N_1498,N_1414);
or U2229 (N_2229,N_581,N_878);
or U2230 (N_2230,N_1388,N_1630);
or U2231 (N_2231,N_264,N_1854);
and U2232 (N_2232,N_580,N_1699);
nor U2233 (N_2233,N_649,N_1274);
or U2234 (N_2234,N_237,N_399);
and U2235 (N_2235,N_880,N_866);
nor U2236 (N_2236,N_836,N_1210);
nor U2237 (N_2237,N_1950,N_696);
or U2238 (N_2238,N_1251,N_1045);
nor U2239 (N_2239,N_998,N_143);
and U2240 (N_2240,N_951,N_1344);
nor U2241 (N_2241,N_1389,N_1335);
or U2242 (N_2242,N_100,N_784);
and U2243 (N_2243,N_482,N_364);
and U2244 (N_2244,N_678,N_1124);
and U2245 (N_2245,N_235,N_109);
nand U2246 (N_2246,N_1622,N_253);
and U2247 (N_2247,N_854,N_761);
nor U2248 (N_2248,N_1749,N_1116);
nor U2249 (N_2249,N_974,N_1795);
nor U2250 (N_2250,N_1597,N_361);
nand U2251 (N_2251,N_1258,N_423);
nand U2252 (N_2252,N_174,N_115);
or U2253 (N_2253,N_126,N_1379);
nor U2254 (N_2254,N_345,N_1004);
nor U2255 (N_2255,N_1387,N_307);
or U2256 (N_2256,N_1282,N_1551);
and U2257 (N_2257,N_43,N_517);
nor U2258 (N_2258,N_1693,N_1975);
and U2259 (N_2259,N_1496,N_799);
nor U2260 (N_2260,N_359,N_1589);
and U2261 (N_2261,N_1735,N_1741);
nor U2262 (N_2262,N_342,N_1329);
and U2263 (N_2263,N_400,N_1627);
and U2264 (N_2264,N_1374,N_61);
or U2265 (N_2265,N_1890,N_169);
or U2266 (N_2266,N_452,N_1427);
and U2267 (N_2267,N_614,N_1884);
or U2268 (N_2268,N_1429,N_1961);
and U2269 (N_2269,N_1880,N_193);
and U2270 (N_2270,N_1260,N_145);
nor U2271 (N_2271,N_1545,N_40);
nor U2272 (N_2272,N_1158,N_1553);
and U2273 (N_2273,N_80,N_903);
nor U2274 (N_2274,N_996,N_1733);
and U2275 (N_2275,N_1781,N_1674);
nand U2276 (N_2276,N_1844,N_1915);
nor U2277 (N_2277,N_41,N_620);
nor U2278 (N_2278,N_828,N_907);
or U2279 (N_2279,N_1967,N_1368);
nor U2280 (N_2280,N_1194,N_1234);
nand U2281 (N_2281,N_904,N_624);
and U2282 (N_2282,N_1587,N_74);
nand U2283 (N_2283,N_1267,N_1345);
nor U2284 (N_2284,N_323,N_1171);
nand U2285 (N_2285,N_348,N_463);
nand U2286 (N_2286,N_893,N_1373);
nand U2287 (N_2287,N_692,N_1588);
nor U2288 (N_2288,N_1441,N_1447);
and U2289 (N_2289,N_282,N_1338);
nand U2290 (N_2290,N_310,N_575);
or U2291 (N_2291,N_736,N_713);
nand U2292 (N_2292,N_917,N_578);
nand U2293 (N_2293,N_388,N_1908);
and U2294 (N_2294,N_1895,N_1395);
or U2295 (N_2295,N_1157,N_426);
nand U2296 (N_2296,N_876,N_505);
and U2297 (N_2297,N_124,N_1226);
or U2298 (N_2298,N_1058,N_1227);
nand U2299 (N_2299,N_1641,N_1969);
nor U2300 (N_2300,N_1799,N_1946);
or U2301 (N_2301,N_512,N_1285);
nor U2302 (N_2302,N_1409,N_890);
or U2303 (N_2303,N_1617,N_1659);
or U2304 (N_2304,N_451,N_1808);
and U2305 (N_2305,N_1151,N_1456);
nor U2306 (N_2306,N_28,N_1044);
nand U2307 (N_2307,N_319,N_1953);
and U2308 (N_2308,N_1930,N_502);
and U2309 (N_2309,N_638,N_1393);
nand U2310 (N_2310,N_1705,N_1864);
or U2311 (N_2311,N_417,N_1902);
nor U2312 (N_2312,N_1779,N_852);
or U2313 (N_2313,N_582,N_524);
nand U2314 (N_2314,N_750,N_1039);
or U2315 (N_2315,N_278,N_191);
nand U2316 (N_2316,N_1736,N_166);
or U2317 (N_2317,N_379,N_557);
or U2318 (N_2318,N_740,N_1532);
or U2319 (N_2319,N_484,N_428);
and U2320 (N_2320,N_573,N_1202);
nor U2321 (N_2321,N_1748,N_382);
nor U2322 (N_2322,N_848,N_1556);
nor U2323 (N_2323,N_24,N_1598);
nor U2324 (N_2324,N_976,N_101);
or U2325 (N_2325,N_685,N_1110);
nor U2326 (N_2326,N_1104,N_963);
or U2327 (N_2327,N_1023,N_1726);
or U2328 (N_2328,N_421,N_76);
and U2329 (N_2329,N_283,N_687);
and U2330 (N_2330,N_205,N_1524);
or U2331 (N_2331,N_1439,N_1625);
nand U2332 (N_2332,N_337,N_717);
and U2333 (N_2333,N_1250,N_1490);
nand U2334 (N_2334,N_621,N_985);
or U2335 (N_2335,N_1399,N_1422);
nand U2336 (N_2336,N_1351,N_919);
nor U2337 (N_2337,N_1475,N_1365);
nand U2338 (N_2338,N_948,N_988);
nor U2339 (N_2339,N_381,N_465);
or U2340 (N_2340,N_547,N_1415);
or U2341 (N_2341,N_1255,N_536);
or U2342 (N_2342,N_1787,N_725);
nand U2343 (N_2343,N_1792,N_922);
nor U2344 (N_2344,N_1360,N_383);
nand U2345 (N_2345,N_1839,N_1353);
nand U2346 (N_2346,N_1363,N_1670);
nand U2347 (N_2347,N_529,N_481);
nand U2348 (N_2348,N_479,N_1600);
or U2349 (N_2349,N_429,N_1236);
and U2350 (N_2350,N_1114,N_885);
and U2351 (N_2351,N_633,N_537);
and U2352 (N_2352,N_1467,N_1919);
or U2353 (N_2353,N_689,N_1698);
nor U2354 (N_2354,N_138,N_1421);
nand U2355 (N_2355,N_478,N_1684);
nor U2356 (N_2356,N_1965,N_1676);
nor U2357 (N_2357,N_1611,N_1634);
and U2358 (N_2358,N_731,N_946);
nand U2359 (N_2359,N_1650,N_316);
nor U2360 (N_2360,N_413,N_1784);
or U2361 (N_2361,N_574,N_445);
nand U2362 (N_2362,N_1230,N_786);
or U2363 (N_2363,N_1208,N_1770);
nor U2364 (N_2364,N_1247,N_200);
and U2365 (N_2365,N_1027,N_1853);
nor U2366 (N_2366,N_883,N_1015);
or U2367 (N_2367,N_1672,N_680);
nor U2368 (N_2368,N_851,N_1339);
and U2369 (N_2369,N_954,N_1704);
or U2370 (N_2370,N_1849,N_1461);
and U2371 (N_2371,N_1366,N_1813);
nor U2372 (N_2372,N_543,N_766);
nand U2373 (N_2373,N_1292,N_898);
nand U2374 (N_2374,N_443,N_374);
or U2375 (N_2375,N_30,N_991);
nand U2376 (N_2376,N_509,N_1130);
nand U2377 (N_2377,N_1572,N_664);
or U2378 (N_2378,N_199,N_800);
or U2379 (N_2379,N_157,N_613);
or U2380 (N_2380,N_309,N_1923);
nor U2381 (N_2381,N_179,N_516);
xnor U2382 (N_2382,N_1990,N_990);
and U2383 (N_2383,N_1614,N_312);
nor U2384 (N_2384,N_1832,N_1742);
and U2385 (N_2385,N_1402,N_1994);
nor U2386 (N_2386,N_1134,N_583);
and U2387 (N_2387,N_1763,N_1405);
and U2388 (N_2388,N_644,N_1371);
nand U2389 (N_2389,N_1324,N_1246);
and U2390 (N_2390,N_1820,N_1697);
nand U2391 (N_2391,N_1928,N_265);
nand U2392 (N_2392,N_357,N_858);
nor U2393 (N_2393,N_466,N_785);
or U2394 (N_2394,N_1183,N_1471);
and U2395 (N_2395,N_1978,N_775);
and U2396 (N_2396,N_219,N_901);
and U2397 (N_2397,N_520,N_1407);
or U2398 (N_2398,N_1328,N_1443);
or U2399 (N_2399,N_172,N_812);
and U2400 (N_2400,N_1096,N_303);
or U2401 (N_2401,N_341,N_1760);
nor U2402 (N_2402,N_322,N_185);
nor U2403 (N_2403,N_1812,N_131);
nand U2404 (N_2404,N_973,N_1362);
nor U2405 (N_2405,N_311,N_397);
or U2406 (N_2406,N_1048,N_1072);
nand U2407 (N_2407,N_737,N_1785);
nand U2408 (N_2408,N_1432,N_22);
or U2409 (N_2409,N_1942,N_1372);
and U2410 (N_2410,N_241,N_1452);
nor U2411 (N_2411,N_1931,N_528);
nand U2412 (N_2412,N_1913,N_437);
nand U2413 (N_2413,N_1870,N_1991);
or U2414 (N_2414,N_1509,N_1381);
or U2415 (N_2415,N_1038,N_469);
nor U2416 (N_2416,N_500,N_588);
or U2417 (N_2417,N_450,N_1643);
or U2418 (N_2418,N_467,N_1231);
and U2419 (N_2419,N_1797,N_389);
nor U2420 (N_2420,N_1309,N_1531);
or U2421 (N_2421,N_1831,N_132);
xor U2422 (N_2422,N_1311,N_376);
nand U2423 (N_2423,N_939,N_449);
or U2424 (N_2424,N_281,N_363);
nand U2425 (N_2425,N_768,N_850);
or U2426 (N_2426,N_287,N_1976);
or U2427 (N_2427,N_544,N_1491);
nor U2428 (N_2428,N_1346,N_552);
and U2429 (N_2429,N_684,N_926);
nand U2430 (N_2430,N_874,N_153);
nand U2431 (N_2431,N_1070,N_586);
and U2432 (N_2432,N_1128,N_1722);
nor U2433 (N_2433,N_32,N_818);
and U2434 (N_2434,N_223,N_1506);
and U2435 (N_2435,N_471,N_29);
nor U2436 (N_2436,N_1937,N_1800);
and U2437 (N_2437,N_643,N_1322);
nand U2438 (N_2438,N_1046,N_178);
and U2439 (N_2439,N_1034,N_1174);
and U2440 (N_2440,N_1866,N_886);
or U2441 (N_2441,N_372,N_982);
or U2442 (N_2442,N_1526,N_201);
or U2443 (N_2443,N_272,N_1459);
and U2444 (N_2444,N_1057,N_523);
nor U2445 (N_2445,N_1802,N_338);
and U2446 (N_2446,N_1486,N_144);
or U2447 (N_2447,N_627,N_245);
nor U2448 (N_2448,N_1804,N_476);
nand U2449 (N_2449,N_918,N_1626);
nand U2450 (N_2450,N_819,N_541);
nor U2451 (N_2451,N_1619,N_666);
nand U2452 (N_2452,N_1557,N_1290);
nand U2453 (N_2453,N_1026,N_1637);
nor U2454 (N_2454,N_593,N_118);
nor U2455 (N_2455,N_117,N_325);
or U2456 (N_2456,N_824,N_439);
nor U2457 (N_2457,N_1355,N_1451);
or U2458 (N_2458,N_1730,N_68);
nor U2459 (N_2459,N_1063,N_107);
nor U2460 (N_2460,N_195,N_550);
and U2461 (N_2461,N_207,N_518);
and U2462 (N_2462,N_788,N_1586);
nand U2463 (N_2463,N_719,N_710);
nor U2464 (N_2464,N_1759,N_648);
nor U2465 (N_2465,N_1343,N_1240);
nand U2466 (N_2466,N_1340,N_1005);
or U2467 (N_2467,N_650,N_274);
nand U2468 (N_2468,N_569,N_91);
nor U2469 (N_2469,N_244,N_589);
and U2470 (N_2470,N_1357,N_1002);
or U2471 (N_2471,N_365,N_1501);
nand U2472 (N_2472,N_1827,N_1837);
nand U2473 (N_2473,N_526,N_1025);
nor U2474 (N_2474,N_139,N_597);
and U2475 (N_2475,N_1718,N_248);
nand U2476 (N_2476,N_1321,N_1807);
or U2477 (N_2477,N_957,N_1959);
nand U2478 (N_2478,N_560,N_1620);
or U2479 (N_2479,N_743,N_299);
or U2480 (N_2480,N_1872,N_1299);
and U2481 (N_2481,N_1239,N_1905);
nor U2482 (N_2482,N_35,N_1397);
nor U2483 (N_2483,N_1719,N_595);
nor U2484 (N_2484,N_1423,N_1550);
nor U2485 (N_2485,N_1144,N_159);
nor U2486 (N_2486,N_611,N_881);
and U2487 (N_2487,N_546,N_712);
nor U2488 (N_2488,N_123,N_1411);
nand U2489 (N_2489,N_277,N_950);
and U2490 (N_2490,N_180,N_1303);
nor U2491 (N_2491,N_579,N_834);
nor U2492 (N_2492,N_1582,N_431);
or U2493 (N_2493,N_1161,N_1448);
and U2494 (N_2494,N_108,N_1082);
nand U2495 (N_2495,N_57,N_1739);
nor U2496 (N_2496,N_1120,N_1384);
and U2497 (N_2497,N_1314,N_1775);
nand U2498 (N_2498,N_1333,N_1111);
and U2499 (N_2499,N_1149,N_1665);
or U2500 (N_2500,N_1318,N_1544);
or U2501 (N_2501,N_1616,N_1579);
nor U2502 (N_2502,N_228,N_1502);
or U2503 (N_2503,N_707,N_726);
nand U2504 (N_2504,N_667,N_1276);
or U2505 (N_2505,N_1000,N_329);
and U2506 (N_2506,N_639,N_1815);
nand U2507 (N_2507,N_1152,N_840);
nand U2508 (N_2508,N_458,N_1570);
and U2509 (N_2509,N_977,N_739);
and U2510 (N_2510,N_838,N_1019);
nor U2511 (N_2511,N_899,N_688);
or U2512 (N_2512,N_186,N_1067);
and U2513 (N_2513,N_1708,N_1995);
nand U2514 (N_2514,N_1478,N_280);
nand U2515 (N_2515,N_1457,N_953);
and U2516 (N_2516,N_844,N_1179);
and U2517 (N_2517,N_986,N_1580);
or U2518 (N_2518,N_849,N_816);
and U2519 (N_2519,N_161,N_1098);
nand U2520 (N_2520,N_1088,N_634);
or U2521 (N_2521,N_1217,N_324);
nor U2522 (N_2522,N_1139,N_832);
and U2523 (N_2523,N_1347,N_62);
and U2524 (N_2524,N_1418,N_285);
nor U2525 (N_2525,N_1753,N_1484);
nand U2526 (N_2526,N_1645,N_805);
or U2527 (N_2527,N_1223,N_295);
nor U2528 (N_2528,N_1278,N_1369);
nand U2529 (N_2529,N_913,N_106);
nand U2530 (N_2530,N_305,N_418);
or U2531 (N_2531,N_1973,N_288);
nand U2532 (N_2532,N_1181,N_1396);
nand U2533 (N_2533,N_1780,N_1404);
and U2534 (N_2534,N_1235,N_989);
nor U2535 (N_2535,N_1618,N_1003);
nor U2536 (N_2536,N_691,N_1711);
nor U2537 (N_2537,N_39,N_1480);
nand U2538 (N_2538,N_1707,N_1575);
or U2539 (N_2539,N_1916,N_1055);
and U2540 (N_2540,N_495,N_1576);
and U2541 (N_2541,N_1176,N_1757);
nand U2542 (N_2542,N_1101,N_756);
and U2543 (N_2543,N_1681,N_1982);
nand U2544 (N_2544,N_1517,N_254);
or U2545 (N_2545,N_1917,N_1342);
and U2546 (N_2546,N_605,N_378);
nand U2547 (N_2547,N_1803,N_1825);
nand U2548 (N_2548,N_551,N_992);
nor U2549 (N_2549,N_513,N_914);
or U2550 (N_2550,N_1535,N_1566);
and U2551 (N_2551,N_1107,N_1295);
and U2552 (N_2552,N_1814,N_813);
or U2553 (N_2553,N_1822,N_935);
nor U2554 (N_2554,N_1752,N_1898);
and U2555 (N_2555,N_231,N_234);
nor U2556 (N_2556,N_1874,N_1077);
nor U2557 (N_2557,N_1408,N_475);
nand U2558 (N_2558,N_1446,N_1583);
nor U2559 (N_2559,N_1275,N_339);
or U2560 (N_2560,N_1155,N_401);
nor U2561 (N_2561,N_273,N_1603);
nor U2562 (N_2562,N_1743,N_1762);
or U2563 (N_2563,N_733,N_1527);
nor U2564 (N_2564,N_1080,N_1585);
nor U2565 (N_2565,N_1552,N_408);
nor U2566 (N_2566,N_1878,N_226);
nor U2567 (N_2567,N_1173,N_1901);
nor U2568 (N_2568,N_1993,N_522);
or U2569 (N_2569,N_94,N_1184);
nor U2570 (N_2570,N_435,N_1323);
nand U2571 (N_2571,N_386,N_1615);
or U2572 (N_2572,N_1090,N_697);
and U2573 (N_2573,N_825,N_204);
nand U2574 (N_2574,N_576,N_1528);
or U2575 (N_2575,N_1458,N_1483);
nor U2576 (N_2576,N_567,N_229);
or U2577 (N_2577,N_1970,N_1382);
and U2578 (N_2578,N_1728,N_681);
nand U2579 (N_2579,N_1713,N_98);
and U2580 (N_2580,N_146,N_1325);
and U2581 (N_2581,N_468,N_301);
and U2582 (N_2582,N_1269,N_747);
and U2583 (N_2583,N_314,N_1538);
nand U2584 (N_2584,N_1798,N_250);
nor U2585 (N_2585,N_1126,N_1541);
or U2586 (N_2586,N_669,N_300);
or U2587 (N_2587,N_1944,N_1220);
nor U2588 (N_2588,N_1962,N_645);
nor U2589 (N_2589,N_1163,N_1031);
and U2590 (N_2590,N_1050,N_1949);
and U2591 (N_2591,N_787,N_1022);
nand U2592 (N_2592,N_1450,N_239);
or U2593 (N_2593,N_375,N_915);
and U2594 (N_2594,N_1732,N_92);
and U2595 (N_2595,N_744,N_1493);
and U2596 (N_2596,N_1476,N_1776);
and U2597 (N_2597,N_980,N_1910);
and U2598 (N_2598,N_454,N_742);
or U2599 (N_2599,N_1069,N_1011);
nand U2600 (N_2600,N_1992,N_395);
nor U2601 (N_2601,N_1903,N_175);
or U2602 (N_2602,N_1667,N_268);
or U2603 (N_2603,N_773,N_619);
xor U2604 (N_2604,N_263,N_1232);
and U2605 (N_2605,N_1100,N_490);
nand U2606 (N_2606,N_1059,N_757);
nand U2607 (N_2607,N_702,N_1664);
nand U2608 (N_2608,N_212,N_1142);
and U2609 (N_2609,N_1277,N_568);
nand U2610 (N_2610,N_864,N_1981);
nand U2611 (N_2611,N_1131,N_1136);
nand U2612 (N_2612,N_1725,N_3);
and U2613 (N_2613,N_1682,N_1093);
nor U2614 (N_2614,N_1390,N_1999);
nand U2615 (N_2615,N_965,N_921);
nor U2616 (N_2616,N_1466,N_1629);
nor U2617 (N_2617,N_1197,N_1542);
nor U2618 (N_2618,N_18,N_705);
and U2619 (N_2619,N_760,N_1548);
nor U2620 (N_2620,N_447,N_1649);
or U2621 (N_2621,N_211,N_1525);
or U2622 (N_2622,N_905,N_981);
nand U2623 (N_2623,N_1122,N_1444);
or U2624 (N_2624,N_371,N_993);
and U2625 (N_2625,N_1876,N_1014);
nor U2626 (N_2626,N_63,N_1463);
nor U2627 (N_2627,N_1877,N_501);
or U2628 (N_2628,N_141,N_1823);
and U2629 (N_2629,N_1013,N_52);
or U2630 (N_2630,N_995,N_358);
nor U2631 (N_2631,N_1783,N_896);
or U2632 (N_2632,N_50,N_83);
nor U2633 (N_2633,N_1939,N_660);
or U2634 (N_2634,N_86,N_1971);
and U2635 (N_2635,N_370,N_1398);
and U2636 (N_2636,N_923,N_1791);
or U2637 (N_2637,N_865,N_148);
nand U2638 (N_2638,N_781,N_1651);
nand U2639 (N_2639,N_13,N_202);
nor U2640 (N_2640,N_609,N_1655);
and U2641 (N_2641,N_116,N_867);
or U2642 (N_2642,N_630,N_88);
nand U2643 (N_2643,N_1113,N_778);
nand U2644 (N_2644,N_1178,N_486);
and U2645 (N_2645,N_1859,N_10);
nand U2646 (N_2646,N_839,N_734);
or U2647 (N_2647,N_1307,N_1273);
and U2648 (N_2648,N_515,N_1148);
nor U2649 (N_2649,N_1454,N_661);
nand U2650 (N_2650,N_26,N_572);
nand U2651 (N_2651,N_533,N_1112);
nor U2652 (N_2652,N_96,N_1419);
nor U2653 (N_2653,N_723,N_1574);
or U2654 (N_2654,N_1494,N_1033);
and U2655 (N_2655,N_1433,N_835);
or U2656 (N_2656,N_806,N_534);
nand U2657 (N_2657,N_1881,N_93);
or U2658 (N_2658,N_1140,N_1786);
or U2659 (N_2659,N_1715,N_599);
nand U2660 (N_2660,N_1747,N_150);
and U2661 (N_2661,N_1313,N_615);
or U2662 (N_2662,N_1558,N_1656);
and U2663 (N_2663,N_430,N_20);
nor U2664 (N_2664,N_1686,N_1262);
or U2665 (N_2665,N_861,N_440);
xnor U2666 (N_2666,N_349,N_227);
or U2667 (N_2667,N_937,N_1420);
nand U2668 (N_2668,N_1690,N_1639);
nor U2669 (N_2669,N_1243,N_617);
nand U2670 (N_2670,N_1146,N_1253);
and U2671 (N_2671,N_384,N_1653);
nor U2672 (N_2672,N_407,N_815);
nand U2673 (N_2673,N_889,N_398);
and U2674 (N_2674,N_952,N_794);
nand U2675 (N_2675,N_827,N_1662);
nor U2676 (N_2676,N_1,N_218);
nor U2677 (N_2677,N_128,N_1933);
and U2678 (N_2678,N_1094,N_209);
nor U2679 (N_2679,N_1883,N_1108);
or U2680 (N_2680,N_987,N_1840);
and U2681 (N_2681,N_354,N_21);
or U2682 (N_2682,N_347,N_983);
or U2683 (N_2683,N_1028,N_1838);
nand U2684 (N_2684,N_721,N_596);
nor U2685 (N_2685,N_198,N_181);
and U2686 (N_2686,N_296,N_715);
nand U2687 (N_2687,N_862,N_1400);
or U2688 (N_2688,N_978,N_507);
or U2689 (N_2689,N_1102,N_1065);
nor U2690 (N_2690,N_326,N_1367);
nor U2691 (N_2691,N_1904,N_1417);
nor U2692 (N_2692,N_1855,N_1477);
nor U2693 (N_2693,N_275,N_607);
nand U2694 (N_2694,N_330,N_1229);
nand U2695 (N_2695,N_1001,N_1103);
nor U2696 (N_2696,N_564,N_686);
nand U2697 (N_2697,N_971,N_970);
nor U2698 (N_2698,N_1186,N_1869);
or U2699 (N_2699,N_695,N_548);
or U2700 (N_2700,N_636,N_64);
and U2701 (N_2701,N_236,N_931);
and U2702 (N_2702,N_48,N_1636);
nand U2703 (N_2703,N_1985,N_1378);
and U2704 (N_2704,N_1774,N_1455);
nor U2705 (N_2705,N_720,N_755);
nor U2706 (N_2706,N_1359,N_698);
or U2707 (N_2707,N_774,N_753);
nand U2708 (N_2708,N_260,N_1943);
nand U2709 (N_2709,N_1601,N_1464);
or U2710 (N_2710,N_1882,N_732);
and U2711 (N_2711,N_879,N_127);
and U2712 (N_2712,N_11,N_870);
nor U2713 (N_2713,N_894,N_1788);
or U2714 (N_2714,N_845,N_1926);
nor U2715 (N_2715,N_902,N_436);
and U2716 (N_2716,N_598,N_489);
or U2717 (N_2717,N_657,N_1468);
and U2718 (N_2718,N_629,N_540);
and U2719 (N_2719,N_49,N_1308);
and U2720 (N_2720,N_1794,N_809);
or U2721 (N_2721,N_170,N_920);
or U2722 (N_2722,N_959,N_938);
or U2723 (N_2723,N_777,N_95);
nand U2724 (N_2724,N_941,N_906);
and U2725 (N_2725,N_1209,N_368);
nor U2726 (N_2726,N_1469,N_1612);
nor U2727 (N_2727,N_1071,N_642);
or U2728 (N_2728,N_618,N_459);
or U2729 (N_2729,N_1474,N_830);
nor U2730 (N_2730,N_1727,N_1710);
or U2731 (N_2731,N_1963,N_1745);
nor U2732 (N_2732,N_1692,N_1744);
nor U2733 (N_2733,N_70,N_1437);
or U2734 (N_2734,N_853,N_604);
nor U2735 (N_2735,N_924,N_1834);
nand U2736 (N_2736,N_290,N_741);
or U2737 (N_2737,N_60,N_1678);
or U2738 (N_2738,N_1879,N_196);
or U2739 (N_2739,N_1828,N_658);
nand U2740 (N_2740,N_90,N_130);
nand U2741 (N_2741,N_328,N_246);
or U2742 (N_2742,N_289,N_1424);
nor U2743 (N_2743,N_1165,N_882);
nor U2744 (N_2744,N_1060,N_1296);
nor U2745 (N_2745,N_1473,N_585);
and U2746 (N_2746,N_1885,N_1306);
nor U2747 (N_2747,N_735,N_499);
nor U2748 (N_2748,N_1865,N_197);
and U2749 (N_2749,N_1700,N_1648);
and U2750 (N_2750,N_1008,N_1569);
nor U2751 (N_2751,N_1241,N_1036);
and U2752 (N_2752,N_663,N_1138);
nand U2753 (N_2753,N_527,N_1216);
nor U2754 (N_2754,N_1066,N_1951);
and U2755 (N_2755,N_860,N_1932);
nand U2756 (N_2756,N_1442,N_525);
nand U2757 (N_2757,N_790,N_1016);
and U2758 (N_2758,N_1434,N_1954);
and U2759 (N_2759,N_351,N_257);
nor U2760 (N_2760,N_765,N_1167);
nor U2761 (N_2761,N_1635,N_504);
nor U2762 (N_2762,N_1790,N_1326);
and U2763 (N_2763,N_554,N_1605);
and U2764 (N_2764,N_448,N_165);
nand U2765 (N_2765,N_728,N_1559);
nand U2766 (N_2766,N_968,N_1086);
nand U2767 (N_2767,N_1280,N_129);
or U2768 (N_2768,N_1259,N_238);
nand U2769 (N_2769,N_776,N_1305);
and U2770 (N_2770,N_1337,N_332);
nand U2771 (N_2771,N_1886,N_271);
nor U2772 (N_2772,N_151,N_1376);
and U2773 (N_2773,N_1125,N_1121);
or U2774 (N_2774,N_745,N_1851);
nand U2775 (N_2775,N_1522,N_422);
and U2776 (N_2776,N_1150,N_934);
nand U2777 (N_2777,N_1465,N_1772);
nand U2778 (N_2778,N_1470,N_668);
or U2779 (N_2779,N_1040,N_1988);
nand U2780 (N_2780,N_1546,N_1647);
nor U2781 (N_2781,N_1573,N_763);
nor U2782 (N_2782,N_1177,N_1482);
and U2783 (N_2783,N_1079,N_868);
and U2784 (N_2784,N_1567,N_1170);
and U2785 (N_2785,N_1811,N_1462);
or U2786 (N_2786,N_405,N_1301);
or U2787 (N_2787,N_699,N_1289);
or U2788 (N_2788,N_558,N_1068);
nand U2789 (N_2789,N_1413,N_37);
or U2790 (N_2790,N_1817,N_932);
and U2791 (N_2791,N_1265,N_700);
or U2792 (N_2792,N_559,N_1900);
nand U2793 (N_2793,N_444,N_321);
and U2794 (N_2794,N_1948,N_491);
and U2795 (N_2795,N_494,N_1330);
and U2796 (N_2796,N_470,N_1638);
or U2797 (N_2797,N_168,N_1479);
nand U2798 (N_2798,N_1248,N_855);
or U2799 (N_2799,N_631,N_1554);
and U2800 (N_2800,N_1549,N_44);
xor U2801 (N_2801,N_1773,N_1074);
or U2802 (N_2802,N_1632,N_1518);
nor U2803 (N_2803,N_1801,N_1242);
nand U2804 (N_2804,N_1997,N_1564);
nor U2805 (N_2805,N_1621,N_1986);
or U2806 (N_2806,N_807,N_1203);
nand U2807 (N_2807,N_566,N_676);
xor U2808 (N_2808,N_1771,N_928);
nand U2809 (N_2809,N_1833,N_1132);
or U2810 (N_2810,N_136,N_1979);
or U2811 (N_2811,N_1654,N_791);
nand U2812 (N_2812,N_956,N_125);
nand U2813 (N_2813,N_1310,N_1754);
and U2814 (N_2814,N_1852,N_1182);
nand U2815 (N_2815,N_622,N_416);
or U2816 (N_2816,N_892,N_220);
nor U2817 (N_2817,N_1435,N_1889);
or U2818 (N_2818,N_1737,N_637);
nor U2819 (N_2819,N_1642,N_1159);
and U2820 (N_2820,N_1119,N_344);
or U2821 (N_2821,N_1685,N_1037);
nor U2822 (N_2822,N_511,N_703);
nor U2823 (N_2823,N_306,N_1286);
and U2824 (N_2824,N_1515,N_1091);
or U2825 (N_2825,N_1222,N_1826);
nand U2826 (N_2826,N_1633,N_571);
nand U2827 (N_2827,N_1843,N_1431);
nand U2828 (N_2828,N_1543,N_591);
or U2829 (N_2829,N_1983,N_353);
nand U2830 (N_2830,N_142,N_1237);
or U2831 (N_2831,N_1358,N_1200);
or U2832 (N_2832,N_1861,N_1964);
or U2833 (N_2833,N_820,N_1436);
nor U2834 (N_2834,N_561,N_1640);
nor U2835 (N_2835,N_4,N_1268);
and U2836 (N_2836,N_651,N_9);
and U2837 (N_2837,N_403,N_545);
nor U2838 (N_2838,N_793,N_811);
nand U2839 (N_2839,N_1087,N_754);
nor U2840 (N_2840,N_912,N_751);
nor U2841 (N_2841,N_1092,N_1445);
nand U2842 (N_2842,N_1987,N_315);
and U2843 (N_2843,N_304,N_979);
nand U2844 (N_2844,N_1192,N_1571);
nor U2845 (N_2845,N_1190,N_318);
nand U2846 (N_2846,N_1960,N_1945);
and U2847 (N_2847,N_45,N_1578);
and U2848 (N_2848,N_1888,N_1315);
or U2849 (N_2849,N_498,N_1064);
or U2850 (N_2850,N_362,N_5);
and U2851 (N_2851,N_1386,N_727);
or U2852 (N_2852,N_1261,N_1511);
or U2853 (N_2853,N_553,N_1206);
or U2854 (N_2854,N_137,N_1488);
and U2855 (N_2855,N_1472,N_1891);
nor U2856 (N_2856,N_532,N_53);
nand U2857 (N_2857,N_215,N_1906);
or U2858 (N_2858,N_1024,N_1720);
and U2859 (N_2859,N_1846,N_1254);
and U2860 (N_2860,N_704,N_674);
or U2861 (N_2861,N_1106,N_1934);
nor U2862 (N_2862,N_214,N_1485);
nor U2863 (N_2863,N_817,N_233);
and U2864 (N_2864,N_1764,N_461);
or U2865 (N_2865,N_51,N_1830);
nand U2866 (N_2866,N_1201,N_610);
nand U2867 (N_2867,N_562,N_113);
nor U2868 (N_2868,N_152,N_655);
or U2869 (N_2869,N_1042,N_1679);
and U2870 (N_2870,N_1565,N_1519);
or U2871 (N_2871,N_1836,N_1302);
and U2872 (N_2872,N_1560,N_243);
and U2873 (N_2873,N_87,N_313);
and U2874 (N_2874,N_340,N_1160);
or U2875 (N_2875,N_298,N_1394);
nor U2876 (N_2876,N_1213,N_355);
or U2877 (N_2877,N_628,N_1871);
or U2878 (N_2878,N_1320,N_662);
nor U2879 (N_2879,N_415,N_1912);
nor U2880 (N_2880,N_230,N_327);
or U2881 (N_2881,N_927,N_1695);
or U2882 (N_2882,N_771,N_1180);
nor U2883 (N_2883,N_1563,N_1805);
or U2884 (N_2884,N_79,N_1756);
nor U2885 (N_2885,N_1863,N_1998);
and U2886 (N_2886,N_994,N_1778);
or U2887 (N_2887,N_1702,N_164);
nand U2888 (N_2888,N_1052,N_1512);
or U2889 (N_2889,N_373,N_1952);
nor U2890 (N_2890,N_1591,N_1777);
and U2891 (N_2891,N_984,N_722);
and U2892 (N_2892,N_147,N_961);
nand U2893 (N_2893,N_1887,N_1989);
nor U2894 (N_2894,N_1533,N_1714);
and U2895 (N_2895,N_792,N_1272);
nand U2896 (N_2896,N_1221,N_1927);
nor U2897 (N_2897,N_999,N_1041);
nor U2898 (N_2898,N_1204,N_65);
or U2899 (N_2899,N_1816,N_1845);
nand U2900 (N_2900,N_438,N_380);
nor U2901 (N_2901,N_1658,N_1751);
and U2902 (N_2902,N_104,N_519);
nand U2903 (N_2903,N_1352,N_1401);
or U2904 (N_2904,N_656,N_1765);
or U2905 (N_2905,N_134,N_590);
and U2906 (N_2906,N_292,N_1829);
nand U2907 (N_2907,N_335,N_446);
nand U2908 (N_2908,N_872,N_1481);
nand U2909 (N_2909,N_1361,N_1312);
and U2910 (N_2910,N_78,N_266);
or U2911 (N_2911,N_888,N_409);
or U2912 (N_2912,N_261,N_1487);
or U2913 (N_2913,N_616,N_1410);
nand U2914 (N_2914,N_156,N_758);
nor U2915 (N_2915,N_1175,N_975);
and U2916 (N_2916,N_1249,N_646);
nand U2917 (N_2917,N_1555,N_1271);
nand U2918 (N_2918,N_804,N_182);
nor U2919 (N_2919,N_1873,N_1304);
or U2920 (N_2920,N_38,N_1143);
nor U2921 (N_2921,N_693,N_1438);
nor U2922 (N_2922,N_1129,N_1521);
nand U2923 (N_2923,N_1644,N_111);
or U2924 (N_2924,N_103,N_267);
and U2925 (N_2925,N_895,N_1370);
xor U2926 (N_2926,N_225,N_1592);
or U2927 (N_2927,N_1127,N_875);
or U2928 (N_2928,N_1012,N_1195);
nor U2929 (N_2929,N_425,N_1740);
and U2930 (N_2930,N_276,N_173);
or U2931 (N_2931,N_477,N_67);
and U2932 (N_2932,N_1284,N_1893);
nor U2933 (N_2933,N_1516,N_1049);
and U2934 (N_2934,N_1924,N_1375);
nor U2935 (N_2935,N_110,N_1594);
nor U2936 (N_2936,N_189,N_514);
and U2937 (N_2937,N_1712,N_1406);
and U2938 (N_2938,N_255,N_66);
and U2939 (N_2939,N_1219,N_1281);
nor U2940 (N_2940,N_1701,N_1608);
nand U2941 (N_2941,N_404,N_670);
nand U2942 (N_2942,N_336,N_1316);
or U2943 (N_2943,N_966,N_1162);
and U2944 (N_2944,N_1966,N_538);
nor U2945 (N_2945,N_1508,N_333);
or U2946 (N_2946,N_320,N_119);
nor U2947 (N_2947,N_75,N_356);
nor U2948 (N_2948,N_1425,N_1624);
or U2949 (N_2949,N_1244,N_222);
and U2950 (N_2950,N_1660,N_73);
or U2951 (N_2951,N_1862,N_873);
nor U2952 (N_2952,N_12,N_718);
and U2953 (N_2953,N_555,N_608);
nand U2954 (N_2954,N_1860,N_1687);
nor U2955 (N_2955,N_1689,N_346);
nor U2956 (N_2956,N_869,N_1006);
nor U2957 (N_2957,N_1957,N_706);
nor U2958 (N_2958,N_521,N_34);
or U2959 (N_2959,N_192,N_510);
nand U2960 (N_2960,N_258,N_1850);
nor U2961 (N_2961,N_247,N_249);
and U2962 (N_2962,N_493,N_433);
or U2963 (N_2963,N_1947,N_1099);
nor U2964 (N_2964,N_1193,N_1666);
and U2965 (N_2965,N_112,N_1806);
or U2966 (N_2966,N_530,N_360);
xnor U2967 (N_2967,N_1166,N_1145);
nand U2968 (N_2968,N_1215,N_1974);
and U2969 (N_2969,N_1669,N_724);
nor U2970 (N_2970,N_730,N_224);
or U2971 (N_2971,N_1768,N_1604);
nor U2972 (N_2972,N_434,N_122);
or U2973 (N_2973,N_925,N_1782);
or U2974 (N_2974,N_492,N_1841);
nor U2975 (N_2975,N_14,N_27);
or U2976 (N_2976,N_1084,N_1858);
nand U2977 (N_2977,N_1238,N_762);
xor U2978 (N_2978,N_474,N_1118);
nor U2979 (N_2979,N_424,N_1584);
and U2980 (N_2980,N_1520,N_1609);
and U2981 (N_2981,N_473,N_1977);
nor U2982 (N_2982,N_240,N_453);
or U2983 (N_2983,N_6,N_302);
nand U2984 (N_2984,N_1769,N_842);
nor U2985 (N_2985,N_1341,N_1925);
nor U2986 (N_2986,N_1503,N_764);
and U2987 (N_2987,N_1189,N_1568);
nor U2988 (N_2988,N_1602,N_1198);
nor U2989 (N_2989,N_1848,N_677);
and U2990 (N_2990,N_942,N_1416);
nand U2991 (N_2991,N_814,N_803);
nand U2992 (N_2992,N_402,N_279);
nor U2993 (N_2993,N_1030,N_217);
nand U2994 (N_2994,N_1529,N_1300);
and U2995 (N_2995,N_1968,N_1510);
nor U2996 (N_2996,N_291,N_1918);
nand U2997 (N_2997,N_690,N_1207);
and U2998 (N_2998,N_859,N_949);
or U2999 (N_2999,N_947,N_1264);
nor U3000 (N_3000,N_794,N_1095);
or U3001 (N_3001,N_1152,N_619);
and U3002 (N_3002,N_1314,N_374);
and U3003 (N_3003,N_1666,N_1964);
or U3004 (N_3004,N_576,N_509);
nand U3005 (N_3005,N_219,N_1693);
nand U3006 (N_3006,N_871,N_551);
nor U3007 (N_3007,N_1838,N_1066);
nor U3008 (N_3008,N_493,N_808);
and U3009 (N_3009,N_675,N_951);
nand U3010 (N_3010,N_755,N_788);
and U3011 (N_3011,N_549,N_399);
nand U3012 (N_3012,N_724,N_1840);
nor U3013 (N_3013,N_703,N_267);
nor U3014 (N_3014,N_1708,N_578);
or U3015 (N_3015,N_128,N_1425);
nor U3016 (N_3016,N_150,N_719);
nand U3017 (N_3017,N_1477,N_205);
nand U3018 (N_3018,N_1075,N_1423);
nand U3019 (N_3019,N_733,N_237);
nand U3020 (N_3020,N_1406,N_1595);
and U3021 (N_3021,N_512,N_1907);
nor U3022 (N_3022,N_1890,N_420);
nand U3023 (N_3023,N_1273,N_216);
or U3024 (N_3024,N_1391,N_1745);
and U3025 (N_3025,N_1467,N_653);
or U3026 (N_3026,N_1517,N_1762);
and U3027 (N_3027,N_40,N_1803);
or U3028 (N_3028,N_869,N_1576);
or U3029 (N_3029,N_1853,N_1647);
and U3030 (N_3030,N_38,N_683);
and U3031 (N_3031,N_1541,N_271);
and U3032 (N_3032,N_1743,N_1707);
and U3033 (N_3033,N_1617,N_1179);
and U3034 (N_3034,N_1994,N_1040);
nor U3035 (N_3035,N_330,N_1458);
or U3036 (N_3036,N_436,N_1267);
and U3037 (N_3037,N_1085,N_1755);
nand U3038 (N_3038,N_477,N_458);
or U3039 (N_3039,N_1379,N_1138);
nand U3040 (N_3040,N_545,N_260);
and U3041 (N_3041,N_1209,N_1670);
nand U3042 (N_3042,N_1330,N_1912);
nor U3043 (N_3043,N_1726,N_926);
nand U3044 (N_3044,N_1322,N_214);
and U3045 (N_3045,N_1694,N_1360);
or U3046 (N_3046,N_1798,N_91);
or U3047 (N_3047,N_1431,N_1689);
and U3048 (N_3048,N_1653,N_1567);
and U3049 (N_3049,N_1282,N_1058);
nor U3050 (N_3050,N_126,N_123);
or U3051 (N_3051,N_740,N_590);
nand U3052 (N_3052,N_1329,N_994);
and U3053 (N_3053,N_213,N_284);
nand U3054 (N_3054,N_1951,N_1999);
nor U3055 (N_3055,N_840,N_1775);
and U3056 (N_3056,N_963,N_1807);
and U3057 (N_3057,N_1934,N_387);
nand U3058 (N_3058,N_1697,N_1941);
nand U3059 (N_3059,N_1573,N_1731);
nor U3060 (N_3060,N_535,N_1003);
and U3061 (N_3061,N_1777,N_1189);
or U3062 (N_3062,N_1891,N_280);
nand U3063 (N_3063,N_972,N_1743);
nor U3064 (N_3064,N_318,N_1106);
nand U3065 (N_3065,N_376,N_928);
nand U3066 (N_3066,N_1561,N_782);
and U3067 (N_3067,N_1599,N_1673);
nand U3068 (N_3068,N_754,N_1306);
or U3069 (N_3069,N_221,N_1055);
nand U3070 (N_3070,N_1710,N_1438);
and U3071 (N_3071,N_1788,N_1648);
nor U3072 (N_3072,N_166,N_26);
or U3073 (N_3073,N_1562,N_903);
and U3074 (N_3074,N_612,N_485);
and U3075 (N_3075,N_79,N_768);
and U3076 (N_3076,N_466,N_1512);
nand U3077 (N_3077,N_891,N_170);
nand U3078 (N_3078,N_1613,N_967);
nor U3079 (N_3079,N_197,N_1427);
nand U3080 (N_3080,N_1482,N_1024);
and U3081 (N_3081,N_580,N_1869);
or U3082 (N_3082,N_1065,N_1889);
or U3083 (N_3083,N_1711,N_1060);
or U3084 (N_3084,N_1322,N_1367);
and U3085 (N_3085,N_452,N_597);
nor U3086 (N_3086,N_104,N_1440);
nor U3087 (N_3087,N_1819,N_1688);
or U3088 (N_3088,N_896,N_483);
nor U3089 (N_3089,N_1349,N_742);
nand U3090 (N_3090,N_397,N_709);
and U3091 (N_3091,N_988,N_959);
or U3092 (N_3092,N_1474,N_1123);
and U3093 (N_3093,N_335,N_1488);
or U3094 (N_3094,N_959,N_858);
or U3095 (N_3095,N_1499,N_1641);
or U3096 (N_3096,N_1302,N_1562);
nor U3097 (N_3097,N_1250,N_1068);
nor U3098 (N_3098,N_1689,N_1773);
nor U3099 (N_3099,N_1486,N_1424);
nor U3100 (N_3100,N_220,N_450);
nand U3101 (N_3101,N_1190,N_734);
nand U3102 (N_3102,N_971,N_540);
nand U3103 (N_3103,N_418,N_111);
and U3104 (N_3104,N_674,N_62);
nand U3105 (N_3105,N_1386,N_1753);
or U3106 (N_3106,N_1961,N_381);
and U3107 (N_3107,N_362,N_1996);
nand U3108 (N_3108,N_1037,N_685);
or U3109 (N_3109,N_1277,N_1000);
and U3110 (N_3110,N_294,N_1001);
and U3111 (N_3111,N_1796,N_1448);
or U3112 (N_3112,N_1507,N_390);
nand U3113 (N_3113,N_902,N_952);
nand U3114 (N_3114,N_1493,N_1873);
or U3115 (N_3115,N_777,N_1881);
nand U3116 (N_3116,N_1024,N_1017);
or U3117 (N_3117,N_364,N_438);
or U3118 (N_3118,N_1397,N_272);
nand U3119 (N_3119,N_1491,N_1888);
and U3120 (N_3120,N_836,N_1744);
nand U3121 (N_3121,N_418,N_694);
nand U3122 (N_3122,N_1451,N_56);
nand U3123 (N_3123,N_1753,N_1585);
or U3124 (N_3124,N_1344,N_1001);
nand U3125 (N_3125,N_314,N_1785);
or U3126 (N_3126,N_639,N_1198);
and U3127 (N_3127,N_699,N_381);
nor U3128 (N_3128,N_819,N_1450);
nor U3129 (N_3129,N_794,N_1120);
or U3130 (N_3130,N_970,N_862);
or U3131 (N_3131,N_1809,N_1672);
and U3132 (N_3132,N_1745,N_1952);
or U3133 (N_3133,N_988,N_920);
or U3134 (N_3134,N_1211,N_969);
nand U3135 (N_3135,N_813,N_1566);
nand U3136 (N_3136,N_613,N_1025);
or U3137 (N_3137,N_1445,N_339);
xor U3138 (N_3138,N_230,N_1168);
and U3139 (N_3139,N_1495,N_489);
and U3140 (N_3140,N_181,N_1059);
nor U3141 (N_3141,N_352,N_408);
and U3142 (N_3142,N_1956,N_1149);
nand U3143 (N_3143,N_42,N_1027);
nor U3144 (N_3144,N_1071,N_133);
or U3145 (N_3145,N_1127,N_503);
nor U3146 (N_3146,N_787,N_1446);
and U3147 (N_3147,N_1176,N_752);
nor U3148 (N_3148,N_77,N_425);
nor U3149 (N_3149,N_511,N_1217);
nand U3150 (N_3150,N_598,N_1750);
nand U3151 (N_3151,N_1672,N_606);
nor U3152 (N_3152,N_101,N_193);
and U3153 (N_3153,N_978,N_526);
nand U3154 (N_3154,N_167,N_1955);
and U3155 (N_3155,N_1931,N_1253);
nor U3156 (N_3156,N_176,N_962);
nor U3157 (N_3157,N_1201,N_165);
and U3158 (N_3158,N_1431,N_1523);
nor U3159 (N_3159,N_499,N_1218);
nand U3160 (N_3160,N_1953,N_1831);
or U3161 (N_3161,N_557,N_1337);
or U3162 (N_3162,N_57,N_611);
or U3163 (N_3163,N_1851,N_51);
and U3164 (N_3164,N_1448,N_119);
or U3165 (N_3165,N_171,N_1693);
nand U3166 (N_3166,N_1126,N_1124);
and U3167 (N_3167,N_52,N_1795);
or U3168 (N_3168,N_1496,N_1711);
nor U3169 (N_3169,N_38,N_74);
and U3170 (N_3170,N_702,N_159);
nand U3171 (N_3171,N_1295,N_704);
nand U3172 (N_3172,N_324,N_1240);
or U3173 (N_3173,N_605,N_1408);
nor U3174 (N_3174,N_988,N_921);
nand U3175 (N_3175,N_891,N_1707);
nand U3176 (N_3176,N_1597,N_159);
or U3177 (N_3177,N_188,N_1966);
nor U3178 (N_3178,N_1477,N_1256);
or U3179 (N_3179,N_1157,N_1871);
and U3180 (N_3180,N_207,N_642);
nor U3181 (N_3181,N_1142,N_690);
and U3182 (N_3182,N_1159,N_311);
or U3183 (N_3183,N_246,N_1532);
nor U3184 (N_3184,N_436,N_603);
or U3185 (N_3185,N_1691,N_1457);
and U3186 (N_3186,N_307,N_1168);
or U3187 (N_3187,N_622,N_1275);
and U3188 (N_3188,N_1497,N_1366);
or U3189 (N_3189,N_1168,N_1581);
nand U3190 (N_3190,N_832,N_1948);
nand U3191 (N_3191,N_310,N_1381);
nor U3192 (N_3192,N_346,N_433);
nor U3193 (N_3193,N_840,N_584);
or U3194 (N_3194,N_341,N_1172);
or U3195 (N_3195,N_1418,N_1772);
or U3196 (N_3196,N_1547,N_394);
and U3197 (N_3197,N_1391,N_924);
and U3198 (N_3198,N_10,N_891);
nand U3199 (N_3199,N_618,N_1952);
nand U3200 (N_3200,N_1689,N_135);
xnor U3201 (N_3201,N_963,N_511);
nor U3202 (N_3202,N_1549,N_82);
and U3203 (N_3203,N_93,N_1196);
nand U3204 (N_3204,N_457,N_1292);
nand U3205 (N_3205,N_1786,N_1618);
nor U3206 (N_3206,N_1164,N_1391);
and U3207 (N_3207,N_535,N_22);
nor U3208 (N_3208,N_802,N_530);
nor U3209 (N_3209,N_731,N_1735);
or U3210 (N_3210,N_1396,N_1221);
nor U3211 (N_3211,N_1704,N_1468);
or U3212 (N_3212,N_365,N_659);
nor U3213 (N_3213,N_873,N_624);
nor U3214 (N_3214,N_1495,N_1323);
or U3215 (N_3215,N_288,N_610);
and U3216 (N_3216,N_1030,N_1297);
nor U3217 (N_3217,N_1713,N_1943);
or U3218 (N_3218,N_123,N_159);
nor U3219 (N_3219,N_1082,N_1311);
or U3220 (N_3220,N_865,N_357);
and U3221 (N_3221,N_1458,N_704);
nor U3222 (N_3222,N_726,N_244);
and U3223 (N_3223,N_1357,N_1856);
nand U3224 (N_3224,N_409,N_474);
nand U3225 (N_3225,N_1355,N_683);
and U3226 (N_3226,N_1712,N_1751);
and U3227 (N_3227,N_778,N_70);
nor U3228 (N_3228,N_1534,N_1383);
and U3229 (N_3229,N_245,N_580);
nor U3230 (N_3230,N_523,N_519);
nor U3231 (N_3231,N_1974,N_467);
nand U3232 (N_3232,N_377,N_1058);
nand U3233 (N_3233,N_298,N_743);
or U3234 (N_3234,N_1296,N_1568);
nor U3235 (N_3235,N_1130,N_1365);
or U3236 (N_3236,N_909,N_553);
and U3237 (N_3237,N_578,N_712);
nor U3238 (N_3238,N_986,N_811);
nor U3239 (N_3239,N_1612,N_626);
and U3240 (N_3240,N_493,N_60);
and U3241 (N_3241,N_916,N_968);
nand U3242 (N_3242,N_1136,N_250);
xnor U3243 (N_3243,N_96,N_1554);
and U3244 (N_3244,N_809,N_1994);
nand U3245 (N_3245,N_1850,N_536);
nand U3246 (N_3246,N_30,N_764);
nand U3247 (N_3247,N_280,N_647);
and U3248 (N_3248,N_1338,N_489);
and U3249 (N_3249,N_306,N_636);
or U3250 (N_3250,N_449,N_1730);
or U3251 (N_3251,N_1941,N_1026);
nand U3252 (N_3252,N_959,N_846);
and U3253 (N_3253,N_1014,N_435);
nand U3254 (N_3254,N_705,N_1062);
and U3255 (N_3255,N_1149,N_1400);
nand U3256 (N_3256,N_1563,N_1344);
or U3257 (N_3257,N_1668,N_1872);
and U3258 (N_3258,N_1125,N_581);
nand U3259 (N_3259,N_949,N_960);
nand U3260 (N_3260,N_1547,N_838);
nor U3261 (N_3261,N_404,N_740);
nor U3262 (N_3262,N_481,N_748);
nor U3263 (N_3263,N_952,N_469);
nand U3264 (N_3264,N_1461,N_876);
nand U3265 (N_3265,N_1996,N_394);
xnor U3266 (N_3266,N_1848,N_1372);
nand U3267 (N_3267,N_707,N_1655);
or U3268 (N_3268,N_1261,N_1013);
or U3269 (N_3269,N_1963,N_1081);
or U3270 (N_3270,N_558,N_837);
and U3271 (N_3271,N_186,N_474);
nand U3272 (N_3272,N_429,N_28);
nand U3273 (N_3273,N_595,N_842);
nor U3274 (N_3274,N_25,N_1236);
nor U3275 (N_3275,N_266,N_1235);
and U3276 (N_3276,N_903,N_904);
or U3277 (N_3277,N_589,N_1413);
nor U3278 (N_3278,N_1663,N_1815);
or U3279 (N_3279,N_1791,N_298);
nand U3280 (N_3280,N_1375,N_577);
and U3281 (N_3281,N_717,N_929);
nor U3282 (N_3282,N_1037,N_240);
nor U3283 (N_3283,N_1804,N_1348);
nor U3284 (N_3284,N_339,N_1181);
and U3285 (N_3285,N_951,N_1141);
or U3286 (N_3286,N_1446,N_204);
and U3287 (N_3287,N_85,N_747);
and U3288 (N_3288,N_1846,N_823);
nor U3289 (N_3289,N_1060,N_441);
or U3290 (N_3290,N_1154,N_1623);
and U3291 (N_3291,N_1014,N_315);
nor U3292 (N_3292,N_1724,N_19);
nand U3293 (N_3293,N_1764,N_156);
nand U3294 (N_3294,N_592,N_291);
or U3295 (N_3295,N_1504,N_192);
nor U3296 (N_3296,N_1207,N_779);
and U3297 (N_3297,N_1992,N_565);
nor U3298 (N_3298,N_1904,N_1111);
nand U3299 (N_3299,N_1978,N_1475);
nand U3300 (N_3300,N_546,N_1967);
nor U3301 (N_3301,N_567,N_1158);
nand U3302 (N_3302,N_1288,N_1819);
or U3303 (N_3303,N_1948,N_172);
nand U3304 (N_3304,N_566,N_1586);
nand U3305 (N_3305,N_284,N_1989);
nor U3306 (N_3306,N_1129,N_477);
and U3307 (N_3307,N_139,N_788);
nand U3308 (N_3308,N_1075,N_1157);
nand U3309 (N_3309,N_1456,N_414);
nand U3310 (N_3310,N_1306,N_1210);
and U3311 (N_3311,N_123,N_1335);
nand U3312 (N_3312,N_669,N_792);
nor U3313 (N_3313,N_851,N_1537);
or U3314 (N_3314,N_1999,N_16);
xnor U3315 (N_3315,N_541,N_1652);
or U3316 (N_3316,N_375,N_210);
nor U3317 (N_3317,N_1238,N_1429);
nor U3318 (N_3318,N_1604,N_1007);
nand U3319 (N_3319,N_1643,N_1012);
nor U3320 (N_3320,N_1954,N_1694);
and U3321 (N_3321,N_1283,N_236);
and U3322 (N_3322,N_521,N_726);
nor U3323 (N_3323,N_1107,N_444);
and U3324 (N_3324,N_1594,N_1526);
nor U3325 (N_3325,N_270,N_901);
and U3326 (N_3326,N_716,N_1987);
and U3327 (N_3327,N_193,N_1866);
and U3328 (N_3328,N_1650,N_1793);
nand U3329 (N_3329,N_493,N_558);
nor U3330 (N_3330,N_140,N_1934);
and U3331 (N_3331,N_1881,N_171);
and U3332 (N_3332,N_846,N_1210);
nand U3333 (N_3333,N_957,N_578);
nor U3334 (N_3334,N_347,N_831);
nor U3335 (N_3335,N_431,N_57);
or U3336 (N_3336,N_1231,N_1249);
nor U3337 (N_3337,N_255,N_547);
and U3338 (N_3338,N_1994,N_1253);
or U3339 (N_3339,N_1244,N_543);
and U3340 (N_3340,N_615,N_1249);
nor U3341 (N_3341,N_16,N_1037);
nor U3342 (N_3342,N_1942,N_1634);
nand U3343 (N_3343,N_1923,N_109);
nor U3344 (N_3344,N_1063,N_898);
nor U3345 (N_3345,N_1966,N_911);
nor U3346 (N_3346,N_1543,N_1716);
nand U3347 (N_3347,N_471,N_1364);
and U3348 (N_3348,N_1597,N_264);
and U3349 (N_3349,N_1421,N_1850);
nand U3350 (N_3350,N_1522,N_958);
and U3351 (N_3351,N_381,N_512);
nand U3352 (N_3352,N_1780,N_461);
and U3353 (N_3353,N_579,N_363);
and U3354 (N_3354,N_548,N_1022);
nand U3355 (N_3355,N_346,N_1745);
or U3356 (N_3356,N_972,N_1178);
and U3357 (N_3357,N_0,N_131);
and U3358 (N_3358,N_780,N_1291);
or U3359 (N_3359,N_1562,N_1563);
or U3360 (N_3360,N_1132,N_344);
or U3361 (N_3361,N_689,N_796);
or U3362 (N_3362,N_1778,N_1084);
nand U3363 (N_3363,N_59,N_537);
and U3364 (N_3364,N_1368,N_1632);
nand U3365 (N_3365,N_335,N_1245);
or U3366 (N_3366,N_262,N_1234);
or U3367 (N_3367,N_260,N_482);
nand U3368 (N_3368,N_1863,N_824);
nor U3369 (N_3369,N_1468,N_763);
nand U3370 (N_3370,N_1795,N_1958);
nand U3371 (N_3371,N_1458,N_1738);
nand U3372 (N_3372,N_495,N_1503);
nor U3373 (N_3373,N_855,N_1103);
nand U3374 (N_3374,N_1024,N_563);
and U3375 (N_3375,N_1282,N_1016);
and U3376 (N_3376,N_1932,N_1922);
nand U3377 (N_3377,N_613,N_545);
and U3378 (N_3378,N_1527,N_1357);
or U3379 (N_3379,N_563,N_1817);
and U3380 (N_3380,N_269,N_112);
or U3381 (N_3381,N_610,N_1055);
nor U3382 (N_3382,N_1739,N_1193);
nand U3383 (N_3383,N_1928,N_1895);
or U3384 (N_3384,N_373,N_1693);
nor U3385 (N_3385,N_1317,N_1044);
xor U3386 (N_3386,N_1468,N_199);
nor U3387 (N_3387,N_1873,N_1705);
nor U3388 (N_3388,N_247,N_15);
or U3389 (N_3389,N_660,N_1590);
and U3390 (N_3390,N_1818,N_294);
or U3391 (N_3391,N_1148,N_458);
and U3392 (N_3392,N_1575,N_1207);
or U3393 (N_3393,N_1535,N_165);
nor U3394 (N_3394,N_899,N_1766);
nand U3395 (N_3395,N_116,N_1041);
and U3396 (N_3396,N_1397,N_367);
nand U3397 (N_3397,N_1783,N_687);
or U3398 (N_3398,N_631,N_536);
nor U3399 (N_3399,N_406,N_95);
and U3400 (N_3400,N_731,N_457);
and U3401 (N_3401,N_265,N_547);
and U3402 (N_3402,N_1698,N_1618);
nor U3403 (N_3403,N_1365,N_1730);
nand U3404 (N_3404,N_1791,N_569);
nor U3405 (N_3405,N_1477,N_1621);
and U3406 (N_3406,N_1861,N_1041);
nand U3407 (N_3407,N_1582,N_1501);
or U3408 (N_3408,N_1476,N_955);
or U3409 (N_3409,N_543,N_885);
nand U3410 (N_3410,N_1219,N_1564);
or U3411 (N_3411,N_43,N_1300);
and U3412 (N_3412,N_1968,N_1975);
and U3413 (N_3413,N_1229,N_614);
nand U3414 (N_3414,N_103,N_1314);
or U3415 (N_3415,N_1071,N_317);
nand U3416 (N_3416,N_119,N_881);
or U3417 (N_3417,N_903,N_1555);
or U3418 (N_3418,N_1505,N_42);
xnor U3419 (N_3419,N_283,N_392);
nor U3420 (N_3420,N_1768,N_261);
or U3421 (N_3421,N_1953,N_762);
nand U3422 (N_3422,N_1492,N_1083);
and U3423 (N_3423,N_178,N_1537);
nand U3424 (N_3424,N_1337,N_793);
or U3425 (N_3425,N_760,N_747);
nor U3426 (N_3426,N_587,N_466);
nor U3427 (N_3427,N_150,N_403);
nor U3428 (N_3428,N_677,N_1779);
nor U3429 (N_3429,N_162,N_308);
and U3430 (N_3430,N_183,N_824);
nand U3431 (N_3431,N_679,N_1279);
nand U3432 (N_3432,N_358,N_1684);
or U3433 (N_3433,N_1081,N_1087);
nand U3434 (N_3434,N_559,N_1628);
or U3435 (N_3435,N_1983,N_1869);
and U3436 (N_3436,N_1310,N_250);
or U3437 (N_3437,N_111,N_1324);
and U3438 (N_3438,N_1658,N_1856);
and U3439 (N_3439,N_801,N_1651);
nand U3440 (N_3440,N_304,N_864);
nor U3441 (N_3441,N_92,N_199);
nand U3442 (N_3442,N_34,N_1242);
or U3443 (N_3443,N_495,N_888);
or U3444 (N_3444,N_1684,N_619);
or U3445 (N_3445,N_1160,N_1304);
nand U3446 (N_3446,N_1259,N_1135);
or U3447 (N_3447,N_446,N_146);
nor U3448 (N_3448,N_837,N_1083);
or U3449 (N_3449,N_1560,N_1382);
nand U3450 (N_3450,N_1616,N_1597);
xnor U3451 (N_3451,N_1800,N_84);
xnor U3452 (N_3452,N_1449,N_716);
nand U3453 (N_3453,N_1406,N_1737);
and U3454 (N_3454,N_1263,N_1514);
nor U3455 (N_3455,N_380,N_1871);
nor U3456 (N_3456,N_1965,N_143);
and U3457 (N_3457,N_1698,N_186);
and U3458 (N_3458,N_628,N_1263);
or U3459 (N_3459,N_324,N_540);
and U3460 (N_3460,N_1362,N_1825);
nand U3461 (N_3461,N_1874,N_1790);
nand U3462 (N_3462,N_1164,N_340);
or U3463 (N_3463,N_118,N_584);
nor U3464 (N_3464,N_638,N_284);
or U3465 (N_3465,N_683,N_387);
or U3466 (N_3466,N_450,N_1781);
or U3467 (N_3467,N_1708,N_982);
nand U3468 (N_3468,N_890,N_458);
nand U3469 (N_3469,N_124,N_1531);
or U3470 (N_3470,N_1065,N_474);
and U3471 (N_3471,N_193,N_1240);
and U3472 (N_3472,N_1947,N_913);
or U3473 (N_3473,N_1246,N_322);
or U3474 (N_3474,N_67,N_50);
xnor U3475 (N_3475,N_487,N_1219);
and U3476 (N_3476,N_1473,N_596);
and U3477 (N_3477,N_1431,N_1039);
nand U3478 (N_3478,N_1490,N_1882);
and U3479 (N_3479,N_158,N_18);
and U3480 (N_3480,N_1258,N_38);
and U3481 (N_3481,N_801,N_1120);
and U3482 (N_3482,N_271,N_789);
or U3483 (N_3483,N_3,N_1265);
nor U3484 (N_3484,N_1993,N_1408);
and U3485 (N_3485,N_937,N_1355);
nand U3486 (N_3486,N_425,N_316);
nor U3487 (N_3487,N_954,N_1968);
nand U3488 (N_3488,N_1520,N_556);
nor U3489 (N_3489,N_304,N_479);
nand U3490 (N_3490,N_1853,N_1074);
nor U3491 (N_3491,N_150,N_1607);
or U3492 (N_3492,N_131,N_784);
and U3493 (N_3493,N_1400,N_311);
nand U3494 (N_3494,N_510,N_439);
and U3495 (N_3495,N_1441,N_773);
or U3496 (N_3496,N_1983,N_1270);
or U3497 (N_3497,N_14,N_458);
and U3498 (N_3498,N_552,N_1261);
nand U3499 (N_3499,N_1147,N_1702);
nor U3500 (N_3500,N_1853,N_905);
nand U3501 (N_3501,N_1244,N_1439);
nor U3502 (N_3502,N_939,N_6);
nand U3503 (N_3503,N_1736,N_204);
or U3504 (N_3504,N_508,N_872);
nor U3505 (N_3505,N_472,N_1024);
or U3506 (N_3506,N_442,N_1388);
and U3507 (N_3507,N_200,N_360);
nor U3508 (N_3508,N_470,N_778);
or U3509 (N_3509,N_1269,N_1636);
or U3510 (N_3510,N_1785,N_1609);
or U3511 (N_3511,N_1015,N_445);
nand U3512 (N_3512,N_1731,N_1352);
or U3513 (N_3513,N_55,N_1871);
or U3514 (N_3514,N_1526,N_920);
nor U3515 (N_3515,N_377,N_675);
or U3516 (N_3516,N_464,N_599);
nor U3517 (N_3517,N_1741,N_90);
nand U3518 (N_3518,N_593,N_1768);
or U3519 (N_3519,N_799,N_1495);
and U3520 (N_3520,N_1070,N_1863);
and U3521 (N_3521,N_1774,N_1822);
and U3522 (N_3522,N_920,N_1693);
nand U3523 (N_3523,N_1214,N_221);
nor U3524 (N_3524,N_88,N_1202);
or U3525 (N_3525,N_64,N_67);
or U3526 (N_3526,N_1714,N_1581);
or U3527 (N_3527,N_254,N_1825);
nand U3528 (N_3528,N_1493,N_1504);
nor U3529 (N_3529,N_1069,N_1181);
nand U3530 (N_3530,N_678,N_372);
or U3531 (N_3531,N_1174,N_900);
nand U3532 (N_3532,N_1915,N_395);
and U3533 (N_3533,N_1398,N_180);
and U3534 (N_3534,N_1959,N_1659);
or U3535 (N_3535,N_224,N_1110);
nor U3536 (N_3536,N_203,N_1568);
nand U3537 (N_3537,N_1459,N_5);
nand U3538 (N_3538,N_1425,N_766);
nor U3539 (N_3539,N_70,N_1754);
or U3540 (N_3540,N_260,N_1179);
or U3541 (N_3541,N_1273,N_1157);
nor U3542 (N_3542,N_1774,N_797);
or U3543 (N_3543,N_1718,N_180);
and U3544 (N_3544,N_389,N_497);
or U3545 (N_3545,N_1758,N_371);
or U3546 (N_3546,N_1128,N_1224);
or U3547 (N_3547,N_1698,N_1903);
or U3548 (N_3548,N_507,N_1268);
and U3549 (N_3549,N_1735,N_1991);
nor U3550 (N_3550,N_192,N_175);
nor U3551 (N_3551,N_607,N_909);
or U3552 (N_3552,N_1651,N_90);
and U3553 (N_3553,N_588,N_1004);
and U3554 (N_3554,N_359,N_324);
nor U3555 (N_3555,N_870,N_1282);
or U3556 (N_3556,N_1009,N_1973);
or U3557 (N_3557,N_118,N_942);
and U3558 (N_3558,N_1901,N_460);
or U3559 (N_3559,N_1106,N_232);
or U3560 (N_3560,N_607,N_2);
nor U3561 (N_3561,N_1956,N_978);
and U3562 (N_3562,N_1307,N_1123);
nor U3563 (N_3563,N_1081,N_1016);
or U3564 (N_3564,N_135,N_457);
and U3565 (N_3565,N_1815,N_440);
xor U3566 (N_3566,N_1007,N_1073);
and U3567 (N_3567,N_677,N_1430);
or U3568 (N_3568,N_747,N_383);
and U3569 (N_3569,N_1795,N_335);
and U3570 (N_3570,N_911,N_1167);
or U3571 (N_3571,N_220,N_897);
and U3572 (N_3572,N_1982,N_1533);
nand U3573 (N_3573,N_1245,N_1014);
nand U3574 (N_3574,N_208,N_1950);
and U3575 (N_3575,N_1409,N_1410);
or U3576 (N_3576,N_22,N_1396);
nor U3577 (N_3577,N_391,N_571);
or U3578 (N_3578,N_1703,N_77);
or U3579 (N_3579,N_1465,N_591);
or U3580 (N_3580,N_778,N_844);
or U3581 (N_3581,N_1561,N_1882);
nand U3582 (N_3582,N_1814,N_672);
or U3583 (N_3583,N_316,N_629);
or U3584 (N_3584,N_1911,N_1064);
or U3585 (N_3585,N_162,N_178);
nor U3586 (N_3586,N_1370,N_689);
or U3587 (N_3587,N_622,N_519);
nand U3588 (N_3588,N_690,N_432);
nand U3589 (N_3589,N_326,N_401);
nor U3590 (N_3590,N_470,N_369);
nor U3591 (N_3591,N_243,N_393);
or U3592 (N_3592,N_822,N_1280);
nor U3593 (N_3593,N_1881,N_1842);
or U3594 (N_3594,N_20,N_1889);
or U3595 (N_3595,N_1032,N_1565);
and U3596 (N_3596,N_655,N_927);
or U3597 (N_3597,N_361,N_1456);
and U3598 (N_3598,N_1442,N_638);
nand U3599 (N_3599,N_346,N_243);
nand U3600 (N_3600,N_1333,N_476);
nand U3601 (N_3601,N_33,N_1145);
and U3602 (N_3602,N_1575,N_1987);
nand U3603 (N_3603,N_31,N_234);
or U3604 (N_3604,N_526,N_1387);
nand U3605 (N_3605,N_692,N_1371);
or U3606 (N_3606,N_1715,N_1298);
and U3607 (N_3607,N_161,N_618);
nand U3608 (N_3608,N_1736,N_605);
and U3609 (N_3609,N_1270,N_316);
nand U3610 (N_3610,N_415,N_876);
or U3611 (N_3611,N_384,N_140);
or U3612 (N_3612,N_108,N_1963);
and U3613 (N_3613,N_478,N_1127);
or U3614 (N_3614,N_143,N_720);
or U3615 (N_3615,N_795,N_1833);
nand U3616 (N_3616,N_1655,N_198);
nor U3617 (N_3617,N_1747,N_921);
and U3618 (N_3618,N_484,N_1549);
nand U3619 (N_3619,N_255,N_1440);
and U3620 (N_3620,N_543,N_335);
or U3621 (N_3621,N_1197,N_683);
nand U3622 (N_3622,N_927,N_1628);
and U3623 (N_3623,N_1681,N_660);
nor U3624 (N_3624,N_388,N_649);
or U3625 (N_3625,N_702,N_1693);
and U3626 (N_3626,N_1238,N_1675);
and U3627 (N_3627,N_1134,N_483);
nand U3628 (N_3628,N_638,N_1007);
nand U3629 (N_3629,N_432,N_13);
and U3630 (N_3630,N_1393,N_1868);
or U3631 (N_3631,N_1350,N_823);
and U3632 (N_3632,N_725,N_1917);
or U3633 (N_3633,N_1670,N_1001);
and U3634 (N_3634,N_650,N_65);
and U3635 (N_3635,N_1953,N_1127);
nor U3636 (N_3636,N_713,N_1461);
and U3637 (N_3637,N_558,N_1648);
nor U3638 (N_3638,N_1035,N_862);
and U3639 (N_3639,N_1884,N_891);
nor U3640 (N_3640,N_851,N_253);
nor U3641 (N_3641,N_98,N_774);
or U3642 (N_3642,N_1134,N_972);
and U3643 (N_3643,N_1052,N_632);
nand U3644 (N_3644,N_1684,N_1292);
or U3645 (N_3645,N_373,N_1403);
nor U3646 (N_3646,N_1359,N_170);
or U3647 (N_3647,N_1898,N_1357);
nand U3648 (N_3648,N_1650,N_1091);
nand U3649 (N_3649,N_239,N_253);
nand U3650 (N_3650,N_364,N_43);
and U3651 (N_3651,N_1511,N_406);
and U3652 (N_3652,N_1154,N_1905);
nor U3653 (N_3653,N_414,N_1551);
nor U3654 (N_3654,N_1072,N_1580);
xnor U3655 (N_3655,N_394,N_1862);
and U3656 (N_3656,N_861,N_1464);
and U3657 (N_3657,N_1799,N_311);
or U3658 (N_3658,N_247,N_1585);
nand U3659 (N_3659,N_1415,N_73);
and U3660 (N_3660,N_1929,N_560);
and U3661 (N_3661,N_1899,N_783);
nor U3662 (N_3662,N_417,N_645);
nor U3663 (N_3663,N_979,N_1351);
nand U3664 (N_3664,N_826,N_741);
or U3665 (N_3665,N_1041,N_619);
or U3666 (N_3666,N_530,N_1621);
nor U3667 (N_3667,N_1332,N_916);
or U3668 (N_3668,N_1079,N_73);
nand U3669 (N_3669,N_1558,N_1109);
or U3670 (N_3670,N_652,N_1939);
and U3671 (N_3671,N_1542,N_332);
and U3672 (N_3672,N_188,N_1842);
nor U3673 (N_3673,N_442,N_603);
and U3674 (N_3674,N_1856,N_1174);
or U3675 (N_3675,N_1738,N_831);
nor U3676 (N_3676,N_913,N_1417);
nor U3677 (N_3677,N_452,N_1406);
nand U3678 (N_3678,N_518,N_1472);
or U3679 (N_3679,N_1011,N_1317);
and U3680 (N_3680,N_1833,N_510);
nand U3681 (N_3681,N_421,N_1090);
and U3682 (N_3682,N_1720,N_728);
and U3683 (N_3683,N_288,N_1994);
nand U3684 (N_3684,N_1556,N_589);
nand U3685 (N_3685,N_187,N_980);
nor U3686 (N_3686,N_1979,N_220);
and U3687 (N_3687,N_1131,N_336);
or U3688 (N_3688,N_1108,N_104);
nor U3689 (N_3689,N_1266,N_1433);
or U3690 (N_3690,N_718,N_42);
or U3691 (N_3691,N_1982,N_581);
or U3692 (N_3692,N_782,N_809);
nor U3693 (N_3693,N_1574,N_1021);
and U3694 (N_3694,N_127,N_1954);
nor U3695 (N_3695,N_1181,N_570);
nor U3696 (N_3696,N_329,N_1770);
nand U3697 (N_3697,N_984,N_688);
nor U3698 (N_3698,N_1849,N_1131);
and U3699 (N_3699,N_1944,N_655);
nand U3700 (N_3700,N_961,N_788);
and U3701 (N_3701,N_67,N_673);
nand U3702 (N_3702,N_1937,N_511);
nand U3703 (N_3703,N_1720,N_1426);
nor U3704 (N_3704,N_1858,N_1063);
or U3705 (N_3705,N_1802,N_1062);
or U3706 (N_3706,N_1907,N_1376);
nand U3707 (N_3707,N_465,N_1451);
or U3708 (N_3708,N_966,N_1365);
xor U3709 (N_3709,N_82,N_1967);
and U3710 (N_3710,N_269,N_1297);
and U3711 (N_3711,N_1280,N_798);
nand U3712 (N_3712,N_241,N_1652);
nor U3713 (N_3713,N_1509,N_322);
nor U3714 (N_3714,N_1390,N_406);
or U3715 (N_3715,N_1351,N_1626);
and U3716 (N_3716,N_63,N_338);
and U3717 (N_3717,N_337,N_1687);
xor U3718 (N_3718,N_749,N_1206);
nor U3719 (N_3719,N_1988,N_592);
or U3720 (N_3720,N_1247,N_864);
nand U3721 (N_3721,N_1821,N_343);
and U3722 (N_3722,N_735,N_1920);
and U3723 (N_3723,N_659,N_1270);
and U3724 (N_3724,N_710,N_334);
or U3725 (N_3725,N_498,N_1713);
or U3726 (N_3726,N_681,N_886);
nand U3727 (N_3727,N_1807,N_935);
or U3728 (N_3728,N_959,N_1719);
or U3729 (N_3729,N_1990,N_1847);
nand U3730 (N_3730,N_1192,N_542);
and U3731 (N_3731,N_1057,N_1050);
or U3732 (N_3732,N_391,N_1197);
nor U3733 (N_3733,N_1402,N_1770);
and U3734 (N_3734,N_1678,N_1074);
and U3735 (N_3735,N_458,N_1976);
and U3736 (N_3736,N_1995,N_718);
or U3737 (N_3737,N_265,N_1194);
nand U3738 (N_3738,N_1824,N_858);
or U3739 (N_3739,N_435,N_1460);
nand U3740 (N_3740,N_1053,N_13);
or U3741 (N_3741,N_1804,N_1654);
and U3742 (N_3742,N_1403,N_1770);
or U3743 (N_3743,N_1952,N_1149);
nand U3744 (N_3744,N_1507,N_1194);
nor U3745 (N_3745,N_1618,N_1475);
and U3746 (N_3746,N_1866,N_1201);
nand U3747 (N_3747,N_142,N_420);
nand U3748 (N_3748,N_1834,N_911);
nor U3749 (N_3749,N_1187,N_1293);
or U3750 (N_3750,N_1046,N_1880);
or U3751 (N_3751,N_1070,N_243);
and U3752 (N_3752,N_657,N_336);
nand U3753 (N_3753,N_365,N_335);
nand U3754 (N_3754,N_162,N_705);
nand U3755 (N_3755,N_1145,N_67);
and U3756 (N_3756,N_471,N_1796);
nor U3757 (N_3757,N_1062,N_1552);
or U3758 (N_3758,N_1566,N_1463);
and U3759 (N_3759,N_1328,N_1932);
or U3760 (N_3760,N_220,N_704);
nand U3761 (N_3761,N_1348,N_897);
or U3762 (N_3762,N_460,N_914);
nand U3763 (N_3763,N_1621,N_1153);
nand U3764 (N_3764,N_1020,N_7);
nand U3765 (N_3765,N_134,N_807);
nor U3766 (N_3766,N_1552,N_1050);
nand U3767 (N_3767,N_465,N_1101);
nand U3768 (N_3768,N_1370,N_30);
nand U3769 (N_3769,N_1841,N_1174);
or U3770 (N_3770,N_1981,N_505);
nand U3771 (N_3771,N_894,N_924);
and U3772 (N_3772,N_1786,N_475);
nor U3773 (N_3773,N_1080,N_923);
and U3774 (N_3774,N_69,N_1687);
nor U3775 (N_3775,N_761,N_1388);
and U3776 (N_3776,N_1575,N_1100);
or U3777 (N_3777,N_306,N_1684);
or U3778 (N_3778,N_615,N_1818);
nand U3779 (N_3779,N_837,N_1761);
nand U3780 (N_3780,N_1396,N_783);
or U3781 (N_3781,N_1116,N_848);
or U3782 (N_3782,N_30,N_929);
and U3783 (N_3783,N_1288,N_940);
nand U3784 (N_3784,N_1729,N_1912);
or U3785 (N_3785,N_1683,N_327);
nor U3786 (N_3786,N_413,N_946);
and U3787 (N_3787,N_1864,N_276);
or U3788 (N_3788,N_1750,N_1443);
or U3789 (N_3789,N_821,N_1308);
nor U3790 (N_3790,N_896,N_1503);
nor U3791 (N_3791,N_702,N_1603);
and U3792 (N_3792,N_1921,N_64);
nand U3793 (N_3793,N_1172,N_1374);
nor U3794 (N_3794,N_83,N_1376);
and U3795 (N_3795,N_1864,N_1962);
or U3796 (N_3796,N_1013,N_1342);
nand U3797 (N_3797,N_1517,N_1701);
nand U3798 (N_3798,N_32,N_1527);
nor U3799 (N_3799,N_1640,N_1727);
or U3800 (N_3800,N_1376,N_1999);
and U3801 (N_3801,N_716,N_1371);
nor U3802 (N_3802,N_871,N_426);
nor U3803 (N_3803,N_1376,N_1134);
nand U3804 (N_3804,N_1241,N_1570);
or U3805 (N_3805,N_991,N_827);
and U3806 (N_3806,N_176,N_1701);
or U3807 (N_3807,N_995,N_583);
nand U3808 (N_3808,N_1340,N_1216);
or U3809 (N_3809,N_478,N_952);
nor U3810 (N_3810,N_1510,N_1217);
nor U3811 (N_3811,N_1550,N_198);
and U3812 (N_3812,N_1194,N_766);
xor U3813 (N_3813,N_1431,N_1260);
nor U3814 (N_3814,N_1082,N_26);
nand U3815 (N_3815,N_707,N_490);
xor U3816 (N_3816,N_1436,N_613);
or U3817 (N_3817,N_171,N_1484);
nor U3818 (N_3818,N_1741,N_704);
and U3819 (N_3819,N_1105,N_92);
nand U3820 (N_3820,N_273,N_1996);
and U3821 (N_3821,N_975,N_217);
and U3822 (N_3822,N_1284,N_1628);
and U3823 (N_3823,N_1112,N_1104);
or U3824 (N_3824,N_1869,N_1265);
nor U3825 (N_3825,N_578,N_332);
nor U3826 (N_3826,N_1302,N_133);
or U3827 (N_3827,N_699,N_610);
nand U3828 (N_3828,N_537,N_451);
and U3829 (N_3829,N_817,N_1154);
nand U3830 (N_3830,N_885,N_1399);
nand U3831 (N_3831,N_383,N_916);
nand U3832 (N_3832,N_969,N_1787);
nand U3833 (N_3833,N_919,N_796);
nand U3834 (N_3834,N_618,N_1141);
nor U3835 (N_3835,N_1703,N_1618);
nand U3836 (N_3836,N_203,N_1872);
nor U3837 (N_3837,N_1518,N_1252);
nand U3838 (N_3838,N_645,N_731);
or U3839 (N_3839,N_550,N_290);
nor U3840 (N_3840,N_838,N_1120);
and U3841 (N_3841,N_245,N_242);
nor U3842 (N_3842,N_1626,N_150);
nor U3843 (N_3843,N_1091,N_1505);
or U3844 (N_3844,N_1918,N_466);
nand U3845 (N_3845,N_1304,N_1060);
and U3846 (N_3846,N_1585,N_37);
and U3847 (N_3847,N_835,N_705);
and U3848 (N_3848,N_1861,N_1521);
or U3849 (N_3849,N_985,N_585);
xnor U3850 (N_3850,N_806,N_68);
nand U3851 (N_3851,N_1475,N_461);
or U3852 (N_3852,N_1694,N_1965);
and U3853 (N_3853,N_1498,N_485);
xor U3854 (N_3854,N_1351,N_700);
nand U3855 (N_3855,N_1493,N_1169);
or U3856 (N_3856,N_1591,N_1660);
nand U3857 (N_3857,N_718,N_1048);
nand U3858 (N_3858,N_884,N_328);
and U3859 (N_3859,N_449,N_1053);
or U3860 (N_3860,N_918,N_1740);
nor U3861 (N_3861,N_1956,N_518);
or U3862 (N_3862,N_958,N_731);
or U3863 (N_3863,N_319,N_29);
nor U3864 (N_3864,N_686,N_451);
nand U3865 (N_3865,N_1570,N_435);
nand U3866 (N_3866,N_841,N_1273);
nor U3867 (N_3867,N_1456,N_1833);
or U3868 (N_3868,N_450,N_939);
nand U3869 (N_3869,N_718,N_1288);
and U3870 (N_3870,N_482,N_1746);
or U3871 (N_3871,N_1312,N_1497);
nor U3872 (N_3872,N_1069,N_540);
and U3873 (N_3873,N_1279,N_799);
and U3874 (N_3874,N_1561,N_812);
or U3875 (N_3875,N_1748,N_1944);
and U3876 (N_3876,N_1722,N_635);
or U3877 (N_3877,N_1709,N_641);
nand U3878 (N_3878,N_1079,N_126);
and U3879 (N_3879,N_173,N_619);
nand U3880 (N_3880,N_45,N_338);
nor U3881 (N_3881,N_135,N_946);
xor U3882 (N_3882,N_689,N_488);
nor U3883 (N_3883,N_489,N_450);
and U3884 (N_3884,N_1168,N_1534);
nor U3885 (N_3885,N_622,N_1344);
nor U3886 (N_3886,N_1638,N_710);
nor U3887 (N_3887,N_502,N_1993);
nand U3888 (N_3888,N_1399,N_1913);
or U3889 (N_3889,N_1250,N_1032);
nor U3890 (N_3890,N_253,N_1830);
or U3891 (N_3891,N_601,N_1986);
nor U3892 (N_3892,N_1175,N_1567);
nor U3893 (N_3893,N_224,N_877);
nor U3894 (N_3894,N_1767,N_1716);
and U3895 (N_3895,N_1827,N_1017);
and U3896 (N_3896,N_149,N_1049);
nor U3897 (N_3897,N_1686,N_893);
or U3898 (N_3898,N_1321,N_573);
nor U3899 (N_3899,N_1471,N_1952);
nor U3900 (N_3900,N_1557,N_128);
and U3901 (N_3901,N_544,N_1014);
or U3902 (N_3902,N_915,N_374);
nand U3903 (N_3903,N_1337,N_1994);
nand U3904 (N_3904,N_993,N_1232);
and U3905 (N_3905,N_617,N_1875);
or U3906 (N_3906,N_143,N_1398);
nor U3907 (N_3907,N_1979,N_6);
nand U3908 (N_3908,N_1906,N_672);
or U3909 (N_3909,N_12,N_1092);
nor U3910 (N_3910,N_1909,N_173);
and U3911 (N_3911,N_662,N_640);
nor U3912 (N_3912,N_87,N_1427);
nand U3913 (N_3913,N_1223,N_148);
nand U3914 (N_3914,N_155,N_1109);
or U3915 (N_3915,N_1826,N_406);
nor U3916 (N_3916,N_1741,N_129);
nand U3917 (N_3917,N_127,N_685);
or U3918 (N_3918,N_1154,N_71);
nor U3919 (N_3919,N_1142,N_85);
nand U3920 (N_3920,N_1234,N_464);
or U3921 (N_3921,N_1003,N_132);
nor U3922 (N_3922,N_100,N_655);
nand U3923 (N_3923,N_116,N_834);
nor U3924 (N_3924,N_619,N_1036);
nor U3925 (N_3925,N_1023,N_642);
nand U3926 (N_3926,N_1052,N_535);
nor U3927 (N_3927,N_819,N_984);
and U3928 (N_3928,N_677,N_63);
and U3929 (N_3929,N_201,N_1223);
and U3930 (N_3930,N_749,N_1614);
and U3931 (N_3931,N_152,N_486);
and U3932 (N_3932,N_1852,N_281);
and U3933 (N_3933,N_713,N_474);
nand U3934 (N_3934,N_1750,N_1442);
and U3935 (N_3935,N_1610,N_802);
or U3936 (N_3936,N_1344,N_551);
or U3937 (N_3937,N_60,N_268);
or U3938 (N_3938,N_282,N_360);
and U3939 (N_3939,N_340,N_1147);
or U3940 (N_3940,N_1185,N_1363);
nand U3941 (N_3941,N_44,N_1343);
and U3942 (N_3942,N_536,N_400);
or U3943 (N_3943,N_1830,N_257);
nand U3944 (N_3944,N_1521,N_912);
nand U3945 (N_3945,N_1441,N_571);
nor U3946 (N_3946,N_996,N_1450);
and U3947 (N_3947,N_677,N_327);
and U3948 (N_3948,N_1905,N_706);
or U3949 (N_3949,N_1376,N_30);
and U3950 (N_3950,N_1721,N_809);
xor U3951 (N_3951,N_1792,N_1050);
or U3952 (N_3952,N_460,N_125);
and U3953 (N_3953,N_1804,N_1335);
and U3954 (N_3954,N_1357,N_1034);
or U3955 (N_3955,N_538,N_1249);
nor U3956 (N_3956,N_1808,N_289);
and U3957 (N_3957,N_1531,N_1164);
nor U3958 (N_3958,N_1853,N_1977);
or U3959 (N_3959,N_600,N_1899);
and U3960 (N_3960,N_1521,N_1073);
or U3961 (N_3961,N_1655,N_1797);
or U3962 (N_3962,N_1497,N_919);
or U3963 (N_3963,N_835,N_986);
nor U3964 (N_3964,N_1265,N_578);
nand U3965 (N_3965,N_319,N_1174);
nor U3966 (N_3966,N_724,N_1499);
and U3967 (N_3967,N_1182,N_496);
or U3968 (N_3968,N_761,N_1211);
nand U3969 (N_3969,N_1689,N_1836);
or U3970 (N_3970,N_1345,N_923);
or U3971 (N_3971,N_1638,N_1371);
nor U3972 (N_3972,N_148,N_1842);
nand U3973 (N_3973,N_235,N_1239);
nand U3974 (N_3974,N_555,N_196);
nand U3975 (N_3975,N_1086,N_1302);
and U3976 (N_3976,N_62,N_1270);
or U3977 (N_3977,N_1338,N_814);
and U3978 (N_3978,N_1911,N_1110);
or U3979 (N_3979,N_1332,N_1676);
or U3980 (N_3980,N_150,N_137);
and U3981 (N_3981,N_668,N_1283);
and U3982 (N_3982,N_1547,N_172);
or U3983 (N_3983,N_1684,N_9);
nor U3984 (N_3984,N_642,N_1173);
nand U3985 (N_3985,N_33,N_124);
nand U3986 (N_3986,N_1723,N_1454);
or U3987 (N_3987,N_1363,N_1426);
or U3988 (N_3988,N_461,N_992);
or U3989 (N_3989,N_307,N_1595);
nor U3990 (N_3990,N_841,N_341);
nand U3991 (N_3991,N_1398,N_357);
or U3992 (N_3992,N_447,N_955);
nand U3993 (N_3993,N_850,N_1015);
or U3994 (N_3994,N_677,N_1849);
and U3995 (N_3995,N_37,N_1252);
and U3996 (N_3996,N_1552,N_782);
and U3997 (N_3997,N_330,N_85);
nor U3998 (N_3998,N_1714,N_955);
and U3999 (N_3999,N_1125,N_790);
nor U4000 (N_4000,N_2520,N_3273);
or U4001 (N_4001,N_2454,N_3320);
nand U4002 (N_4002,N_2177,N_3722);
nand U4003 (N_4003,N_3743,N_2437);
or U4004 (N_4004,N_3290,N_3905);
and U4005 (N_4005,N_2489,N_2476);
and U4006 (N_4006,N_2978,N_3545);
nand U4007 (N_4007,N_3166,N_2443);
nand U4008 (N_4008,N_2526,N_3081);
nand U4009 (N_4009,N_3440,N_2933);
nor U4010 (N_4010,N_3329,N_2302);
or U4011 (N_4011,N_2672,N_2523);
nor U4012 (N_4012,N_2692,N_3431);
or U4013 (N_4013,N_3910,N_3709);
and U4014 (N_4014,N_3889,N_2707);
or U4015 (N_4015,N_3310,N_2289);
nand U4016 (N_4016,N_2319,N_3209);
or U4017 (N_4017,N_3216,N_2922);
and U4018 (N_4018,N_2369,N_2524);
or U4019 (N_4019,N_3523,N_3227);
or U4020 (N_4020,N_3628,N_2058);
and U4021 (N_4021,N_3085,N_3206);
nand U4022 (N_4022,N_2111,N_2657);
nand U4023 (N_4023,N_2062,N_2774);
nand U4024 (N_4024,N_2766,N_2876);
nor U4025 (N_4025,N_3571,N_3333);
nand U4026 (N_4026,N_3023,N_2728);
or U4027 (N_4027,N_2085,N_2984);
nor U4028 (N_4028,N_3282,N_3336);
nor U4029 (N_4029,N_2482,N_2130);
nor U4030 (N_4030,N_2535,N_3784);
nor U4031 (N_4031,N_3124,N_3991);
and U4032 (N_4032,N_3264,N_2869);
xor U4033 (N_4033,N_3568,N_2293);
and U4034 (N_4034,N_2093,N_2305);
or U4035 (N_4035,N_2034,N_3297);
nor U4036 (N_4036,N_2142,N_2908);
or U4037 (N_4037,N_2798,N_2378);
nand U4038 (N_4038,N_2272,N_3980);
xnor U4039 (N_4039,N_3351,N_3985);
and U4040 (N_4040,N_2945,N_2417);
and U4041 (N_4041,N_2039,N_2871);
nor U4042 (N_4042,N_3367,N_3009);
nor U4043 (N_4043,N_2426,N_2071);
nor U4044 (N_4044,N_3244,N_3446);
or U4045 (N_4045,N_2965,N_3398);
nor U4046 (N_4046,N_2122,N_2837);
nand U4047 (N_4047,N_2867,N_2644);
nor U4048 (N_4048,N_3445,N_2730);
nor U4049 (N_4049,N_2387,N_2303);
or U4050 (N_4050,N_3704,N_2238);
or U4051 (N_4051,N_2446,N_2820);
or U4052 (N_4052,N_3519,N_3886);
or U4053 (N_4053,N_3155,N_2858);
and U4054 (N_4054,N_3470,N_2159);
nor U4055 (N_4055,N_3186,N_2980);
or U4056 (N_4056,N_3218,N_2271);
nand U4057 (N_4057,N_2488,N_2584);
or U4058 (N_4058,N_2220,N_3253);
nand U4059 (N_4059,N_2214,N_2129);
and U4060 (N_4060,N_2023,N_3777);
or U4061 (N_4061,N_3178,N_2184);
nor U4062 (N_4062,N_2300,N_2602);
or U4063 (N_4063,N_3051,N_2567);
and U4064 (N_4064,N_3631,N_3921);
or U4065 (N_4065,N_2118,N_2340);
nor U4066 (N_4066,N_2061,N_2870);
and U4067 (N_4067,N_2912,N_2020);
nand U4068 (N_4068,N_2325,N_3787);
or U4069 (N_4069,N_2823,N_2659);
nor U4070 (N_4070,N_3228,N_2140);
nand U4071 (N_4071,N_2946,N_2780);
or U4072 (N_4072,N_3661,N_2114);
and U4073 (N_4073,N_3971,N_3851);
nand U4074 (N_4074,N_3334,N_3223);
and U4075 (N_4075,N_3198,N_2491);
nand U4076 (N_4076,N_2606,N_2616);
nand U4077 (N_4077,N_2230,N_3861);
nor U4078 (N_4078,N_2828,N_2669);
nor U4079 (N_4079,N_3232,N_2355);
nand U4080 (N_4080,N_3650,N_3745);
and U4081 (N_4081,N_3823,N_2559);
nor U4082 (N_4082,N_2585,N_2102);
nand U4083 (N_4083,N_2879,N_3619);
or U4084 (N_4084,N_3947,N_3959);
nor U4085 (N_4085,N_3029,N_3516);
or U4086 (N_4086,N_3016,N_3790);
nor U4087 (N_4087,N_3912,N_3603);
nor U4088 (N_4088,N_2449,N_2872);
and U4089 (N_4089,N_3202,N_2237);
or U4090 (N_4090,N_2324,N_3587);
or U4091 (N_4091,N_2030,N_2979);
nand U4092 (N_4092,N_3050,N_3832);
nor U4093 (N_4093,N_3167,N_3427);
nor U4094 (N_4094,N_3354,N_2270);
and U4095 (N_4095,N_2065,N_3387);
nor U4096 (N_4096,N_3379,N_3608);
nor U4097 (N_4097,N_3357,N_3879);
and U4098 (N_4098,N_2985,N_2038);
or U4099 (N_4099,N_3199,N_2508);
and U4100 (N_4100,N_2628,N_2041);
nand U4101 (N_4101,N_3239,N_2124);
or U4102 (N_4102,N_3693,N_3042);
and U4103 (N_4103,N_3998,N_2708);
or U4104 (N_4104,N_2537,N_3741);
and U4105 (N_4105,N_2762,N_3688);
nand U4106 (N_4106,N_3047,N_2888);
and U4107 (N_4107,N_3384,N_2295);
nor U4108 (N_4108,N_3696,N_2241);
or U4109 (N_4109,N_3237,N_3936);
nor U4110 (N_4110,N_2274,N_3113);
and U4111 (N_4111,N_3664,N_2347);
nand U4112 (N_4112,N_2789,N_2103);
nand U4113 (N_4113,N_2599,N_3515);
and U4114 (N_4114,N_2283,N_2685);
or U4115 (N_4115,N_3604,N_2648);
nand U4116 (N_4116,N_2626,N_3829);
nand U4117 (N_4117,N_3478,N_3499);
nor U4118 (N_4118,N_2157,N_3818);
or U4119 (N_4119,N_3188,N_3266);
nand U4120 (N_4120,N_2748,N_2250);
or U4121 (N_4121,N_2905,N_3280);
and U4122 (N_4122,N_2558,N_3916);
and U4123 (N_4123,N_2587,N_3540);
and U4124 (N_4124,N_2060,N_2126);
nor U4125 (N_4125,N_3763,N_2649);
and U4126 (N_4126,N_2741,N_3569);
nand U4127 (N_4127,N_3502,N_3040);
and U4128 (N_4128,N_3952,N_3152);
and U4129 (N_4129,N_3512,N_2370);
and U4130 (N_4130,N_3025,N_2952);
or U4131 (N_4131,N_2601,N_2975);
nand U4132 (N_4132,N_2463,N_2646);
and U4133 (N_4133,N_3090,N_2022);
and U4134 (N_4134,N_3672,N_3459);
nand U4135 (N_4135,N_2950,N_3275);
nor U4136 (N_4136,N_2572,N_3945);
nor U4137 (N_4137,N_3321,N_3110);
nor U4138 (N_4138,N_3561,N_3623);
nand U4139 (N_4139,N_3544,N_2090);
and U4140 (N_4140,N_2320,N_3434);
or U4141 (N_4141,N_2703,N_2328);
nor U4142 (N_4142,N_3795,N_2211);
nand U4143 (N_4143,N_3352,N_3620);
nor U4144 (N_4144,N_2439,N_3481);
or U4145 (N_4145,N_2307,N_3324);
nand U4146 (N_4146,N_2120,N_2788);
nor U4147 (N_4147,N_3965,N_2796);
or U4148 (N_4148,N_2835,N_2045);
nor U4149 (N_4149,N_2019,N_3876);
or U4150 (N_4150,N_3156,N_2059);
nand U4151 (N_4151,N_2278,N_2536);
and U4152 (N_4152,N_3003,N_2393);
nor U4153 (N_4153,N_2132,N_3179);
nand U4154 (N_4154,N_2357,N_3014);
or U4155 (N_4155,N_3225,N_3190);
nor U4156 (N_4156,N_2987,N_3150);
nand U4157 (N_4157,N_3299,N_2252);
nand U4158 (N_4158,N_3098,N_3339);
or U4159 (N_4159,N_3432,N_3476);
nor U4160 (N_4160,N_2873,N_2608);
nand U4161 (N_4161,N_3302,N_3695);
or U4162 (N_4162,N_3773,N_3160);
nand U4163 (N_4163,N_2805,N_2406);
or U4164 (N_4164,N_2215,N_2527);
or U4165 (N_4165,N_3376,N_2944);
nand U4166 (N_4166,N_2051,N_2344);
nand U4167 (N_4167,N_3015,N_2073);
or U4168 (N_4168,N_2885,N_3897);
and U4169 (N_4169,N_2679,N_2433);
nand U4170 (N_4170,N_2219,N_3596);
nand U4171 (N_4171,N_2629,N_2410);
and U4172 (N_4172,N_3260,N_2498);
nor U4173 (N_4173,N_3645,N_2256);
nor U4174 (N_4174,N_3941,N_2574);
and U4175 (N_4175,N_3640,N_2963);
nand U4176 (N_4176,N_2191,N_3843);
nand U4177 (N_4177,N_2461,N_2940);
nand U4178 (N_4178,N_2621,N_3183);
nand U4179 (N_4179,N_3443,N_3994);
nand U4180 (N_4180,N_3929,N_2747);
or U4181 (N_4181,N_2395,N_3812);
and U4182 (N_4182,N_3758,N_3801);
nor U4183 (N_4183,N_3347,N_3041);
or U4184 (N_4184,N_3751,N_3141);
and U4185 (N_4185,N_3067,N_3508);
nand U4186 (N_4186,N_3586,N_3838);
and U4187 (N_4187,N_2752,N_2251);
or U4188 (N_4188,N_2533,N_3769);
and U4189 (N_4189,N_3865,N_2939);
and U4190 (N_4190,N_3538,N_3606);
nand U4191 (N_4191,N_2141,N_2545);
and U4192 (N_4192,N_2560,N_2280);
and U4193 (N_4193,N_2654,N_3529);
and U4194 (N_4194,N_2576,N_3691);
nand U4195 (N_4195,N_2702,N_2036);
or U4196 (N_4196,N_3460,N_3144);
or U4197 (N_4197,N_2898,N_2053);
or U4198 (N_4198,N_3423,N_3142);
and U4199 (N_4199,N_2392,N_3442);
nor U4200 (N_4200,N_3580,N_3417);
nor U4201 (N_4201,N_3217,N_2681);
and U4202 (N_4202,N_3669,N_3740);
nand U4203 (N_4203,N_2530,N_3455);
and U4204 (N_4204,N_3289,N_2786);
or U4205 (N_4205,N_2224,N_2091);
nor U4206 (N_4206,N_2301,N_3720);
or U4207 (N_4207,N_3617,N_3969);
or U4208 (N_4208,N_3161,N_2275);
or U4209 (N_4209,N_2326,N_3415);
nor U4210 (N_4210,N_2334,N_2231);
and U4211 (N_4211,N_3957,N_3500);
and U4212 (N_4212,N_2532,N_2983);
nor U4213 (N_4213,N_2098,N_2429);
nor U4214 (N_4214,N_2901,N_3600);
and U4215 (N_4215,N_3318,N_2442);
nand U4216 (N_4216,N_2209,N_2268);
and U4217 (N_4217,N_2299,N_2166);
or U4218 (N_4218,N_3378,N_3477);
nor U4219 (N_4219,N_2399,N_2595);
or U4220 (N_4220,N_3026,N_3024);
or U4221 (N_4221,N_2791,N_2424);
nor U4222 (N_4222,N_3311,N_3982);
nor U4223 (N_4223,N_2338,N_2714);
nor U4224 (N_4224,N_2206,N_3407);
nor U4225 (N_4225,N_3457,N_2726);
and U4226 (N_4226,N_3782,N_2330);
or U4227 (N_4227,N_3277,N_3159);
or U4228 (N_4228,N_3555,N_2064);
or U4229 (N_4229,N_3059,N_2717);
and U4230 (N_4230,N_3621,N_3272);
and U4231 (N_4231,N_2666,N_3942);
and U4232 (N_4232,N_2242,N_3723);
nor U4233 (N_4233,N_3759,N_3552);
or U4234 (N_4234,N_2232,N_3233);
or U4235 (N_4235,N_2731,N_2017);
nand U4236 (N_4236,N_3556,N_2057);
nor U4237 (N_4237,N_2374,N_3993);
nand U4238 (N_4238,N_3493,N_3461);
and U4239 (N_4239,N_3340,N_2686);
nor U4240 (N_4240,N_3953,N_3590);
or U4241 (N_4241,N_2947,N_3060);
and U4242 (N_4242,N_3316,N_2705);
nor U4243 (N_4243,N_2517,N_3899);
nand U4244 (N_4244,N_3256,N_2787);
nand U4245 (N_4245,N_2240,N_3411);
and U4246 (N_4246,N_2597,N_3656);
or U4247 (N_4247,N_3196,N_2164);
and U4248 (N_4248,N_2312,N_3694);
or U4249 (N_4249,N_3674,N_2630);
nor U4250 (N_4250,N_3662,N_3629);
xnor U4251 (N_4251,N_3510,N_3073);
nand U4252 (N_4252,N_2772,N_2138);
or U4253 (N_4253,N_2739,N_3852);
nor U4254 (N_4254,N_2889,N_3514);
or U4255 (N_4255,N_3197,N_3532);
nand U4256 (N_4256,N_2897,N_3083);
nand U4257 (N_4257,N_3563,N_2381);
nand U4258 (N_4258,N_2638,N_3115);
nor U4259 (N_4259,N_2309,N_2856);
or U4260 (N_4260,N_3007,N_2673);
nand U4261 (N_4261,N_2008,N_3658);
or U4262 (N_4262,N_2037,N_2100);
nor U4263 (N_4263,N_2363,N_2382);
or U4264 (N_4264,N_2863,N_2700);
nand U4265 (N_4265,N_2781,N_2564);
nand U4266 (N_4266,N_2627,N_2723);
and U4267 (N_4267,N_2413,N_3101);
nand U4268 (N_4268,N_3097,N_3961);
or U4269 (N_4269,N_3307,N_3308);
and U4270 (N_4270,N_2834,N_3932);
and U4271 (N_4271,N_3973,N_2173);
and U4272 (N_4272,N_3134,N_2265);
or U4273 (N_4273,N_3541,N_3391);
or U4274 (N_4274,N_3574,N_2988);
nor U4275 (N_4275,N_3395,N_3091);
nor U4276 (N_4276,N_3325,N_2081);
or U4277 (N_4277,N_2131,N_2188);
and U4278 (N_4278,N_2956,N_2487);
or U4279 (N_4279,N_2853,N_3451);
nor U4280 (N_4280,N_2423,N_3995);
nand U4281 (N_4281,N_3419,N_3361);
and U4282 (N_4282,N_2304,N_2298);
or U4283 (N_4283,N_2696,N_3518);
nand U4284 (N_4284,N_2936,N_3813);
nand U4285 (N_4285,N_2063,N_2204);
and U4286 (N_4286,N_2507,N_2455);
and U4287 (N_4287,N_3092,N_3844);
nor U4288 (N_4288,N_2208,N_2553);
nand U4289 (N_4289,N_3659,N_2438);
and U4290 (N_4290,N_3667,N_2317);
nand U4291 (N_4291,N_2931,N_3698);
or U4292 (N_4292,N_3082,N_2116);
nand U4293 (N_4293,N_3283,N_2618);
nor U4294 (N_4294,N_3542,N_3862);
and U4295 (N_4295,N_2440,N_3383);
nand U4296 (N_4296,N_3783,N_2884);
and U4297 (N_4297,N_2479,N_2570);
nand U4298 (N_4298,N_2999,N_3189);
nand U4299 (N_4299,N_3803,N_2525);
and U4300 (N_4300,N_3742,N_3401);
nor U4301 (N_4301,N_3975,N_3986);
nor U4302 (N_4302,N_3360,N_2123);
nor U4303 (N_4303,N_3242,N_3655);
and U4304 (N_4304,N_3356,N_2481);
nor U4305 (N_4305,N_3200,N_2636);
and U4306 (N_4306,N_2807,N_3653);
nor U4307 (N_4307,N_3004,N_2735);
or U4308 (N_4308,N_3808,N_3748);
nor U4309 (N_4309,N_2974,N_3885);
nor U4310 (N_4310,N_2868,N_3229);
or U4311 (N_4311,N_2843,N_2937);
nand U4312 (N_4312,N_2712,N_2765);
and U4313 (N_4313,N_2297,N_3444);
nor U4314 (N_4314,N_2949,N_3647);
or U4315 (N_4315,N_2040,N_2682);
nor U4316 (N_4316,N_2764,N_2113);
nand U4317 (N_4317,N_3099,N_3771);
or U4318 (N_4318,N_3607,N_2631);
nand U4319 (N_4319,N_2821,N_2874);
and U4320 (N_4320,N_3250,N_2435);
nor U4321 (N_4321,N_3682,N_3174);
nand U4322 (N_4322,N_3850,N_3774);
nor U4323 (N_4323,N_3609,N_2284);
nand U4324 (N_4324,N_3687,N_3632);
and U4325 (N_4325,N_3671,N_2906);
nand U4326 (N_4326,N_3344,N_3254);
nor U4327 (N_4327,N_3238,N_3298);
and U4328 (N_4328,N_3725,N_2055);
nor U4329 (N_4329,N_2754,N_3927);
nor U4330 (N_4330,N_3924,N_2623);
nor U4331 (N_4331,N_2571,N_2373);
or U4332 (N_4332,N_3317,N_2941);
and U4333 (N_4333,N_2668,N_2082);
and U4334 (N_4334,N_3887,N_3920);
nand U4335 (N_4335,N_2468,N_3950);
nand U4336 (N_4336,N_2183,N_2360);
or U4337 (N_4337,N_2854,N_3996);
and U4338 (N_4338,N_2234,N_2171);
nand U4339 (N_4339,N_2902,N_3909);
or U4340 (N_4340,N_3724,N_2970);
nand U4341 (N_4341,N_2366,N_2942);
nand U4342 (N_4342,N_3805,N_3900);
and U4343 (N_4343,N_2620,N_3992);
or U4344 (N_4344,N_3210,N_2639);
nand U4345 (N_4345,N_2929,N_2550);
or U4346 (N_4346,N_2108,N_3839);
nand U4347 (N_4347,N_2269,N_2699);
nand U4348 (N_4348,N_3331,N_2803);
nand U4349 (N_4349,N_2266,N_2492);
and U4350 (N_4350,N_2400,N_2257);
nand U4351 (N_4351,N_2989,N_2105);
or U4352 (N_4352,N_2444,N_3281);
nor U4353 (N_4353,N_2002,N_2691);
nand U4354 (N_4354,N_2031,N_2313);
nand U4355 (N_4355,N_2695,N_2331);
and U4356 (N_4356,N_3789,N_3894);
nand U4357 (N_4357,N_3473,N_3718);
nand U4358 (N_4358,N_3911,N_2032);
or U4359 (N_4359,N_2362,N_3093);
or U4360 (N_4360,N_3034,N_2751);
xnor U4361 (N_4361,N_3158,N_3441);
nand U4362 (N_4362,N_2494,N_2009);
nor U4363 (N_4363,N_2542,N_2511);
and U4364 (N_4364,N_3578,N_3588);
nor U4365 (N_4365,N_2194,N_3657);
and U4366 (N_4366,N_3488,N_2877);
nand U4367 (N_4367,N_2086,N_2809);
nor U4368 (N_4368,N_3185,N_3880);
nor U4369 (N_4369,N_3028,N_3312);
nor U4370 (N_4370,N_3262,N_3371);
or U4371 (N_4371,N_3856,N_2150);
and U4372 (N_4372,N_2895,N_3130);
nor U4373 (N_4373,N_3868,N_3319);
and U4374 (N_4374,N_3030,N_2568);
nor U4375 (N_4375,N_3454,N_3102);
nand U4376 (N_4376,N_3875,N_2784);
and U4377 (N_4377,N_3435,N_2697);
or U4378 (N_4378,N_2848,N_3364);
nand U4379 (N_4379,N_3668,N_3939);
nand U4380 (N_4380,N_2948,N_3878);
or U4381 (N_4381,N_2480,N_3666);
or U4382 (N_4382,N_2005,N_2917);
nor U4383 (N_4383,N_3903,N_2580);
and U4384 (N_4384,N_2667,N_3456);
or U4385 (N_4385,N_3859,N_3013);
and U4386 (N_4386,N_2645,N_3602);
and U4387 (N_4387,N_2495,N_3230);
or U4388 (N_4388,N_2408,N_3907);
or U4389 (N_4389,N_3153,N_3278);
or U4390 (N_4390,N_3111,N_3012);
or U4391 (N_4391,N_3468,N_3738);
nand U4392 (N_4392,N_3122,N_3702);
xor U4393 (N_4393,N_2306,N_2997);
and U4394 (N_4394,N_2453,N_2198);
nor U4395 (N_4395,N_2716,N_2418);
nand U4396 (N_4396,N_2401,N_2074);
or U4397 (N_4397,N_3639,N_2662);
nand U4398 (N_4398,N_3690,N_3840);
and U4399 (N_4399,N_3926,N_3491);
and U4400 (N_4400,N_2050,N_2153);
nor U4401 (N_4401,N_3560,N_2971);
nor U4402 (N_4402,N_3106,N_2808);
nor U4403 (N_4403,N_3922,N_2029);
nand U4404 (N_4404,N_3279,N_2862);
and U4405 (N_4405,N_3437,N_2499);
nor U4406 (N_4406,N_3970,N_2187);
nand U4407 (N_4407,N_3827,N_2197);
nor U4408 (N_4408,N_3222,N_2335);
or U4409 (N_4409,N_2701,N_3715);
nand U4410 (N_4410,N_2107,N_3554);
nor U4411 (N_4411,N_2955,N_2954);
or U4412 (N_4412,N_2361,N_2115);
or U4413 (N_4413,N_2007,N_3471);
and U4414 (N_4414,N_3616,N_2407);
nor U4415 (N_4415,N_2160,N_2934);
or U4416 (N_4416,N_2539,N_3974);
and U4417 (N_4417,N_2448,N_3643);
and U4418 (N_4418,N_3775,N_3997);
nor U4419 (N_4419,N_3366,N_2549);
and U4420 (N_4420,N_3353,N_2743);
and U4421 (N_4421,N_3891,N_3389);
and U4422 (N_4422,N_2880,N_2859);
and U4423 (N_4423,N_3768,N_3129);
or U4424 (N_4424,N_3143,N_3065);
or U4425 (N_4425,N_3337,N_3268);
or U4426 (N_4426,N_3145,N_2546);
nand U4427 (N_4427,N_2015,N_2785);
nor U4428 (N_4428,N_3521,N_3436);
nand U4429 (N_4429,N_2811,N_2729);
and U4430 (N_4430,N_2044,N_3076);
or U4431 (N_4431,N_2519,N_2416);
and U4432 (N_4432,N_3753,N_3637);
and U4433 (N_4433,N_3358,N_2758);
nor U4434 (N_4434,N_2918,N_3036);
nand U4435 (N_4435,N_2358,N_2277);
or U4436 (N_4436,N_3240,N_2814);
or U4437 (N_4437,N_3125,N_2991);
nor U4438 (N_4438,N_2004,N_3486);
and U4439 (N_4439,N_3562,N_3677);
or U4440 (N_4440,N_2078,N_2593);
and U4441 (N_4441,N_2202,N_2878);
nor U4442 (N_4442,N_3585,N_3053);
or U4443 (N_4443,N_2321,N_2279);
nand U4444 (N_4444,N_3728,N_3313);
nor U4445 (N_4445,N_3817,N_2793);
nand U4446 (N_4446,N_2779,N_2592);
nor U4447 (N_4447,N_2486,N_2430);
nor U4448 (N_4448,N_2671,N_2561);
nor U4449 (N_4449,N_3565,N_3791);
nor U4450 (N_4450,N_3286,N_3480);
nand U4451 (N_4451,N_3804,N_3438);
nand U4452 (N_4452,N_3410,N_3796);
and U4453 (N_4453,N_3537,N_2385);
and U4454 (N_4454,N_3492,N_3372);
nor U4455 (N_4455,N_2386,N_2706);
and U4456 (N_4456,N_3447,N_3303);
and U4457 (N_4457,N_3749,N_2011);
nor U4458 (N_4458,N_2996,N_3126);
nand U4459 (N_4459,N_3701,N_3304);
nand U4460 (N_4460,N_2195,N_2350);
or U4461 (N_4461,N_2588,N_3573);
and U4462 (N_4462,N_3252,N_3306);
or U4463 (N_4463,N_3261,N_3495);
xnor U4464 (N_4464,N_2087,N_2094);
or U4465 (N_4465,N_2199,N_3931);
nand U4466 (N_4466,N_2722,N_3496);
nand U4467 (N_4467,N_2106,N_2860);
xor U4468 (N_4468,N_2249,N_3760);
nand U4469 (N_4469,N_2590,N_3276);
and U4470 (N_4470,N_3735,N_2169);
nand U4471 (N_4471,N_2981,N_3678);
and U4472 (N_4472,N_3413,N_3448);
or U4473 (N_4473,N_3855,N_2172);
and U4474 (N_4474,N_3780,N_3405);
nor U4475 (N_4475,N_2851,N_3895);
or U4476 (N_4476,N_2452,N_3258);
nand U4477 (N_4477,N_2092,N_3084);
and U4478 (N_4478,N_2972,N_2964);
nand U4479 (N_4479,N_3614,N_3902);
nand U4480 (N_4480,N_3467,N_3660);
nand U4481 (N_4481,N_2790,N_3000);
and U4482 (N_4482,N_3806,N_3187);
or U4483 (N_4483,N_2528,N_2168);
nor U4484 (N_4484,N_3032,N_2921);
nand U4485 (N_4485,N_2891,N_3999);
or U4486 (N_4486,N_2773,N_2846);
or U4487 (N_4487,N_3846,N_3341);
and U4488 (N_4488,N_2579,N_2464);
nor U4489 (N_4489,N_2016,N_2583);
and U4490 (N_4490,N_2738,N_2694);
nand U4491 (N_4491,N_2148,N_3820);
nand U4492 (N_4492,N_2824,N_2190);
and U4493 (N_4493,N_3270,N_3412);
nor U4494 (N_4494,N_3121,N_2333);
or U4495 (N_4495,N_2380,N_3716);
and U4496 (N_4496,N_2842,N_2409);
and U4497 (N_4497,N_3874,N_3954);
or U4498 (N_4498,N_3548,N_2913);
or U4499 (N_4499,N_3021,N_3761);
and U4500 (N_4500,N_3754,N_3734);
and U4501 (N_4501,N_3816,N_3207);
nand U4502 (N_4502,N_2683,N_3330);
nand U4503 (N_4503,N_3853,N_2962);
nand U4504 (N_4504,N_3248,N_3326);
nor U4505 (N_4505,N_2581,N_2367);
nor U4506 (N_4506,N_3972,N_2147);
nand U4507 (N_4507,N_3464,N_2403);
xnor U4508 (N_4508,N_2513,N_3663);
nor U4509 (N_4509,N_2228,N_2596);
or U4510 (N_4510,N_2046,N_2474);
nor U4511 (N_4511,N_3002,N_3234);
or U4512 (N_4512,N_3422,N_2900);
nand U4513 (N_4513,N_3546,N_3884);
nor U4514 (N_4514,N_2052,N_2720);
and U4515 (N_4515,N_2145,N_2925);
and U4516 (N_4516,N_3116,N_3536);
or U4517 (N_4517,N_2915,N_2146);
or U4518 (N_4518,N_2575,N_2158);
and U4519 (N_4519,N_3539,N_2881);
nor U4520 (N_4520,N_3689,N_3214);
or U4521 (N_4521,N_3163,N_3140);
or U4522 (N_4522,N_3956,N_3219);
or U4523 (N_4523,N_3683,N_3171);
or U4524 (N_4524,N_3860,N_3914);
or U4525 (N_4525,N_2441,N_2292);
or U4526 (N_4526,N_2457,N_3837);
or U4527 (N_4527,N_3575,N_2677);
nand U4528 (N_4528,N_2043,N_3168);
or U4529 (N_4529,N_3733,N_3831);
nor U4530 (N_4530,N_2072,N_3766);
or U4531 (N_4531,N_3428,N_3685);
nand U4532 (N_4532,N_3064,N_3680);
nand U4533 (N_4533,N_2149,N_3525);
and U4534 (N_4534,N_3181,N_3605);
or U4535 (N_4535,N_3744,N_2260);
and U4536 (N_4536,N_3375,N_2687);
and U4537 (N_4537,N_2084,N_3466);
nor U4538 (N_4538,N_2000,N_3797);
nor U4539 (N_4539,N_3182,N_2247);
nor U4540 (N_4540,N_2770,N_2200);
or U4541 (N_4541,N_2025,N_3388);
nand U4542 (N_4542,N_3547,N_3088);
xnor U4543 (N_4543,N_2315,N_2656);
and U4544 (N_4544,N_2760,N_2818);
nor U4545 (N_4545,N_2816,N_2756);
nand U4546 (N_4546,N_3483,N_3558);
and U4547 (N_4547,N_2336,N_3534);
and U4548 (N_4548,N_3074,N_3119);
nor U4549 (N_4549,N_2839,N_3108);
and U4550 (N_4550,N_3038,N_3906);
nor U4551 (N_4551,N_3008,N_3854);
or U4552 (N_4552,N_2573,N_2127);
nand U4553 (N_4553,N_3589,N_3430);
and U4554 (N_4554,N_2641,N_3251);
and U4555 (N_4555,N_2089,N_2125);
or U4556 (N_4556,N_2831,N_3641);
and U4557 (N_4557,N_2603,N_3342);
or U4558 (N_4558,N_3913,N_3300);
nor U4559 (N_4559,N_3369,N_2740);
nor U4560 (N_4560,N_2329,N_3504);
or U4561 (N_4561,N_2619,N_3027);
and U4562 (N_4562,N_3528,N_2458);
and U4563 (N_4563,N_2893,N_3901);
or U4564 (N_4564,N_3581,N_2734);
and U4565 (N_4565,N_2541,N_2516);
or U4566 (N_4566,N_3713,N_2391);
and U4567 (N_4567,N_3978,N_2502);
nor U4568 (N_4568,N_2995,N_3634);
nor U4569 (N_4569,N_2664,N_2346);
or U4570 (N_4570,N_2676,N_3983);
nand U4571 (N_4571,N_3944,N_3020);
nand U4572 (N_4572,N_2613,N_2021);
and U4573 (N_4573,N_3424,N_3757);
nand U4574 (N_4574,N_2128,N_2343);
or U4575 (N_4575,N_3807,N_2684);
and U4576 (N_4576,N_3146,N_3221);
or U4577 (N_4577,N_2652,N_2822);
nor U4578 (N_4578,N_3535,N_3648);
nor U4579 (N_4579,N_3194,N_2953);
nand U4580 (N_4580,N_2724,N_3295);
nor U4581 (N_4581,N_3915,N_3636);
nor U4582 (N_4582,N_3706,N_2162);
or U4583 (N_4583,N_2104,N_2389);
and U4584 (N_4584,N_2688,N_3904);
nand U4585 (N_4585,N_3224,N_3612);
nor U4586 (N_4586,N_2727,N_3079);
nor U4587 (N_4587,N_3479,N_2026);
or U4588 (N_4588,N_2478,N_2719);
or U4589 (N_4589,N_2510,N_2144);
or U4590 (N_4590,N_3006,N_2514);
nor U4591 (N_4591,N_3567,N_3964);
nor U4592 (N_4592,N_2286,N_3220);
nor U4593 (N_4593,N_3896,N_3137);
and U4594 (N_4594,N_2792,N_3096);
nand U4595 (N_4595,N_3487,N_3877);
or U4596 (N_4596,N_2914,N_2799);
nor U4597 (N_4597,N_2185,N_2951);
xor U4598 (N_4598,N_3873,N_3871);
and U4599 (N_4599,N_3463,N_2001);
and U4600 (N_4600,N_3984,N_2327);
nor U4601 (N_4601,N_2958,N_3673);
and U4602 (N_4602,N_3255,N_2605);
or U4603 (N_4603,N_3595,N_2882);
or U4604 (N_4604,N_2467,N_3292);
and U4605 (N_4605,N_3989,N_3247);
nand U4606 (N_4606,N_3400,N_2422);
nor U4607 (N_4607,N_2432,N_2076);
and U4608 (N_4608,N_3374,N_2841);
nor U4609 (N_4609,N_2244,N_2591);
or U4610 (N_4610,N_3857,N_2924);
or U4611 (N_4611,N_2308,N_2852);
and U4612 (N_4612,N_2529,N_2753);
nand U4613 (N_4613,N_2661,N_2845);
nor U4614 (N_4614,N_2371,N_3165);
nor U4615 (N_4615,N_3314,N_3136);
nor U4616 (N_4616,N_3559,N_2689);
nand U4617 (N_4617,N_2663,N_3919);
nor U4618 (N_4618,N_3385,N_2316);
nor U4619 (N_4619,N_3511,N_2551);
nor U4620 (N_4620,N_3291,N_2028);
or U4621 (N_4621,N_3406,N_2290);
nor U4622 (N_4622,N_3935,N_2855);
and U4623 (N_4623,N_2182,N_3001);
nor U4624 (N_4624,N_3469,N_2285);
nor U4625 (N_4625,N_2243,N_2680);
nor U4626 (N_4626,N_3627,N_3465);
and U4627 (N_4627,N_3699,N_3930);
nor U4628 (N_4628,N_3613,N_2709);
nor U4629 (N_4629,N_2003,N_2693);
or U4630 (N_4630,N_3781,N_2653);
or U4631 (N_4631,N_2776,N_3752);
or U4632 (N_4632,N_2800,N_3475);
nor U4633 (N_4633,N_3138,N_2365);
nand U4634 (N_4634,N_3069,N_2368);
or U4635 (N_4635,N_2456,N_3810);
nor U4636 (N_4636,N_3285,N_3195);
nor U4637 (N_4637,N_2261,N_2068);
nand U4638 (N_4638,N_3584,N_3582);
or U4639 (N_4639,N_2223,N_2555);
nand U4640 (N_4640,N_3819,N_3809);
nor U4641 (N_4641,N_3294,N_3215);
nor U4642 (N_4642,N_3824,N_3649);
nand U4643 (N_4643,N_2604,N_2763);
or U4644 (N_4644,N_2566,N_2769);
nand U4645 (N_4645,N_3800,N_3892);
and U4646 (N_4646,N_3109,N_2675);
and U4647 (N_4647,N_3458,N_2847);
or U4648 (N_4648,N_3045,N_2259);
nand U4649 (N_4649,N_2887,N_2704);
or U4650 (N_4650,N_3592,N_2761);
and U4651 (N_4651,N_3075,N_2797);
and U4652 (N_4652,N_3315,N_2609);
nor U4653 (N_4653,N_2294,N_2175);
nor U4654 (N_4654,N_2069,N_3208);
and U4655 (N_4655,N_3527,N_2012);
nand U4656 (N_4656,N_2794,N_3390);
nand U4657 (N_4657,N_3946,N_3826);
or U4658 (N_4658,N_3033,N_2518);
and U4659 (N_4659,N_2445,N_2377);
nor U4660 (N_4660,N_3164,N_2923);
nor U4661 (N_4661,N_2414,N_2372);
and U4662 (N_4662,N_3533,N_2600);
and U4663 (N_4663,N_3035,N_3201);
nand U4664 (N_4664,N_3958,N_2462);
nor U4665 (N_4665,N_2436,N_3967);
nor U4666 (N_4666,N_3246,N_3131);
nor U4667 (N_4667,N_3403,N_2547);
and U4668 (N_4668,N_3822,N_2179);
nand U4669 (N_4669,N_3731,N_3044);
and U4670 (N_4670,N_2612,N_3462);
nand U4671 (N_4671,N_2339,N_3828);
nor U4672 (N_4672,N_2633,N_3296);
nor U4673 (N_4673,N_2967,N_3363);
and U4674 (N_4674,N_2804,N_2282);
nand U4675 (N_4675,N_2832,N_3593);
or U4676 (N_4676,N_2014,N_3670);
xnor U4677 (N_4677,N_2460,N_2047);
and U4678 (N_4678,N_3979,N_3531);
or U4679 (N_4679,N_3882,N_2018);
or U4680 (N_4680,N_2725,N_2450);
and U4681 (N_4681,N_2783,N_3750);
and U4682 (N_4682,N_2167,N_3162);
nand U4683 (N_4683,N_2557,N_3429);
nand U4684 (N_4684,N_2291,N_3798);
and U4685 (N_4685,N_3157,N_2112);
or U4686 (N_4686,N_2201,N_2332);
or U4687 (N_4687,N_3729,N_3633);
or U4688 (N_4688,N_3553,N_3017);
or U4689 (N_4689,N_3676,N_2755);
and U4690 (N_4690,N_3231,N_3151);
nand U4691 (N_4691,N_3550,N_2109);
nor U4692 (N_4692,N_3095,N_3043);
nor U4693 (N_4693,N_2864,N_2066);
and U4694 (N_4694,N_3746,N_2910);
nor U4695 (N_4695,N_3867,N_2744);
nor U4696 (N_4696,N_2248,N_3583);
xor U4697 (N_4697,N_3408,N_3087);
and U4698 (N_4698,N_3287,N_2152);
nor U4699 (N_4699,N_3046,N_3416);
or U4700 (N_4700,N_2650,N_3977);
or U4701 (N_4701,N_3103,N_3259);
nand U4702 (N_4702,N_3386,N_2957);
or U4703 (N_4703,N_2625,N_3399);
and U4704 (N_4704,N_3503,N_2548);
and U4705 (N_4705,N_3305,N_2986);
nand U4706 (N_4706,N_2233,N_3192);
and U4707 (N_4707,N_3425,N_3094);
nand U4708 (N_4708,N_3123,N_2670);
nor U4709 (N_4709,N_3149,N_2554);
or U4710 (N_4710,N_2749,N_3133);
nor U4711 (N_4711,N_2151,N_2472);
xor U4712 (N_4712,N_2544,N_3938);
nand U4713 (N_4713,N_3811,N_3147);
nor U4714 (N_4714,N_3019,N_2048);
nor U4715 (N_4715,N_2813,N_3309);
nor U4716 (N_4716,N_3509,N_3381);
nor U4717 (N_4717,N_3058,N_2359);
nand U4718 (N_4718,N_3881,N_2212);
and U4719 (N_4719,N_2447,N_2966);
nor U4720 (N_4720,N_3052,N_2836);
nor U4721 (N_4721,N_2176,N_2830);
or U4722 (N_4722,N_2674,N_3684);
and U4723 (N_4723,N_3530,N_2405);
nand U4724 (N_4724,N_2042,N_2634);
xnor U4725 (N_4725,N_3507,N_2412);
or U4726 (N_4726,N_2135,N_2911);
nor U4727 (N_4727,N_2500,N_3526);
nor U4728 (N_4728,N_3883,N_2154);
nor U4729 (N_4729,N_2276,N_3211);
or U4730 (N_4730,N_3736,N_2431);
or U4731 (N_4731,N_2192,N_2501);
nor U4732 (N_4732,N_2771,N_2732);
nand U4733 (N_4733,N_3501,N_2352);
or U4734 (N_4734,N_3071,N_3054);
and U4735 (N_4735,N_2186,N_2647);
nand U4736 (N_4736,N_2239,N_3786);
nor U4737 (N_4737,N_3730,N_2928);
and U4738 (N_4738,N_3365,N_2099);
nand U4739 (N_4739,N_2095,N_3205);
nor U4740 (N_4740,N_2383,N_2982);
or U4741 (N_4741,N_3452,N_2337);
or U4742 (N_4742,N_2205,N_3263);
nor U4743 (N_4743,N_2750,N_2024);
nand U4744 (N_4744,N_2505,N_2170);
nand U4745 (N_4745,N_2598,N_3426);
and U4746 (N_4746,N_3988,N_2565);
nor U4747 (N_4747,N_3794,N_2833);
and U4748 (N_4748,N_2624,N_3732);
nor U4749 (N_4749,N_2376,N_3721);
and U4750 (N_4750,N_3057,N_3890);
nand U4751 (N_4751,N_2883,N_3990);
nand U4752 (N_4752,N_2196,N_3943);
and U4753 (N_4753,N_2534,N_2990);
or U4754 (N_4754,N_2079,N_3170);
nor U4755 (N_4755,N_2777,N_3841);
nand U4756 (N_4756,N_3236,N_3193);
and U4757 (N_4757,N_3870,N_3599);
or U4758 (N_4758,N_2193,N_2101);
and U4759 (N_4759,N_3373,N_3591);
nor U4760 (N_4760,N_2795,N_3987);
nor U4761 (N_4761,N_3086,N_2977);
and U4762 (N_4762,N_2434,N_3453);
or U4763 (N_4763,N_3089,N_2354);
or U4764 (N_4764,N_3293,N_2733);
or U4765 (N_4765,N_3177,N_2033);
and U4766 (N_4766,N_2637,N_3981);
or U4767 (N_4767,N_2993,N_3450);
and U4768 (N_4768,N_2222,N_2746);
nand U4769 (N_4769,N_2227,N_3719);
nor U4770 (N_4770,N_3864,N_3779);
or U4771 (N_4771,N_3711,N_3271);
and U4772 (N_4772,N_2174,N_2504);
nor U4773 (N_4773,N_3707,N_2136);
or U4774 (N_4774,N_3269,N_2210);
nor U4775 (N_4775,N_2427,N_2866);
or U4776 (N_4776,N_3066,N_2419);
and U4777 (N_4777,N_3635,N_2825);
nor U4778 (N_4778,N_2892,N_3642);
nand U4779 (N_4779,N_2512,N_2345);
nor U4780 (N_4780,N_3010,N_2838);
nand U4781 (N_4781,N_2394,N_3638);
nand U4782 (N_4782,N_2819,N_2894);
and U4783 (N_4783,N_3601,N_3834);
nand U4784 (N_4784,N_3472,N_2471);
nand U4785 (N_4785,N_3037,N_3522);
nor U4786 (N_4786,N_3869,N_2757);
nor U4787 (N_4787,N_3940,N_3127);
nand U4788 (N_4788,N_3180,N_3714);
nand U4789 (N_4789,N_2782,N_3404);
nand U4790 (N_4790,N_3439,N_2916);
nand U4791 (N_4791,N_2484,N_2768);
nand U4792 (N_4792,N_2384,N_2710);
nor U4793 (N_4793,N_3105,N_3346);
nand U4794 (N_4794,N_3393,N_3349);
or U4795 (N_4795,N_2767,N_3355);
nor U4796 (N_4796,N_2351,N_2969);
nand U4797 (N_4797,N_3799,N_2245);
and U4798 (N_4798,N_3433,N_2759);
or U4799 (N_4799,N_2577,N_2607);
and U4800 (N_4800,N_3934,N_2556);
and U4801 (N_4801,N_3622,N_3397);
and U4802 (N_4802,N_3078,N_2397);
nand U4803 (N_4803,N_3770,N_3524);
or U4804 (N_4804,N_2165,N_3888);
xnor U4805 (N_4805,N_2428,N_2678);
and U4806 (N_4806,N_2961,N_3203);
nand U4807 (N_4807,N_3708,N_2156);
nor U4808 (N_4808,N_2006,N_3517);
nor U4809 (N_4809,N_2775,N_3679);
and U4810 (N_4810,N_3489,N_2349);
or U4811 (N_4811,N_3257,N_3100);
nand U4812 (N_4812,N_3288,N_3018);
and U4813 (N_4813,N_3778,N_3335);
or U4814 (N_4814,N_2540,N_2815);
nand U4815 (N_4815,N_2080,N_3618);
nor U4816 (N_4816,N_3863,N_2865);
or U4817 (N_4817,N_2133,N_2610);
nand U4818 (N_4818,N_2509,N_3039);
and U4819 (N_4819,N_2379,N_3830);
nand U4820 (N_4820,N_2919,N_3474);
nand U4821 (N_4821,N_2451,N_3727);
nand U4822 (N_4822,N_2909,N_2907);
or U4823 (N_4823,N_2521,N_3343);
and U4824 (N_4824,N_3772,N_2229);
nand U4825 (N_4825,N_3577,N_3368);
nor U4826 (N_4826,N_3549,N_3597);
and U4827 (N_4827,N_2217,N_2810);
or U4828 (N_4828,N_3362,N_3955);
xnor U4829 (N_4829,N_2163,N_3626);
nor U4830 (N_4830,N_2263,N_2035);
nand U4831 (N_4831,N_3594,N_2470);
or U4832 (N_4832,N_3703,N_2935);
nand U4833 (N_4833,N_2221,N_3825);
or U4834 (N_4834,N_3814,N_2404);
nor U4835 (N_4835,N_2829,N_2943);
or U4836 (N_4836,N_3963,N_2976);
nor U4837 (N_4837,N_2253,N_3359);
or U4838 (N_4838,N_2375,N_2415);
nor U4839 (N_4839,N_2490,N_3243);
or U4840 (N_4840,N_3705,N_3063);
or U4841 (N_4841,N_3566,N_2896);
nand U4842 (N_4842,N_3712,N_3976);
nor U4843 (N_4843,N_2651,N_2056);
or U4844 (N_4844,N_3644,N_2992);
nand U4845 (N_4845,N_2827,N_3739);
nor U4846 (N_4846,N_3418,N_2643);
nand U4847 (N_4847,N_2314,N_3172);
or U4848 (N_4848,N_3697,N_2617);
or U4849 (N_4849,N_2589,N_3402);
or U4850 (N_4850,N_3654,N_2552);
nor U4851 (N_4851,N_2802,N_2181);
or U4852 (N_4852,N_3893,N_3148);
nor U4853 (N_4853,N_2310,N_2563);
and U4854 (N_4854,N_2236,N_2388);
and U4855 (N_4855,N_3414,N_2713);
and U4856 (N_4856,N_3396,N_3767);
and U4857 (N_4857,N_3918,N_2258);
and U4858 (N_4858,N_2622,N_2899);
and U4859 (N_4859,N_2658,N_3928);
nand U4860 (N_4860,N_2077,N_2473);
or U4861 (N_4861,N_2903,N_2497);
nand U4862 (N_4862,N_2806,N_3421);
nor U4863 (N_4863,N_3968,N_3345);
nor U4864 (N_4864,N_2812,N_2522);
or U4865 (N_4865,N_2998,N_3765);
nand U4866 (N_4866,N_2844,N_3394);
or U4867 (N_4867,N_3557,N_3494);
nor U4868 (N_4868,N_3241,N_2049);
nand U4869 (N_4869,N_3611,N_2075);
nor U4870 (N_4870,N_2121,N_2218);
nor U4871 (N_4871,N_2013,N_2960);
or U4872 (N_4872,N_3842,N_2904);
and U4873 (N_4873,N_2690,N_3651);
nand U4874 (N_4874,N_3114,N_3776);
nand U4875 (N_4875,N_3551,N_3031);
or U4876 (N_4876,N_2614,N_3338);
nor U4877 (N_4877,N_3948,N_2110);
or U4878 (N_4878,N_3610,N_2496);
nor U4879 (N_4879,N_3380,N_2067);
and U4880 (N_4880,N_2711,N_3966);
and U4881 (N_4881,N_2890,N_2273);
nand U4882 (N_4882,N_2180,N_3788);
or U4883 (N_4883,N_2255,N_3323);
nand U4884 (N_4884,N_3077,N_3482);
and U4885 (N_4885,N_3049,N_3692);
nand U4886 (N_4886,N_2262,N_2097);
and U4887 (N_4887,N_3267,N_2088);
nand U4888 (N_4888,N_3322,N_2635);
and U4889 (N_4889,N_2515,N_2886);
nand U4890 (N_4890,N_2117,N_3184);
nor U4891 (N_4891,N_2483,N_3062);
nand U4892 (N_4892,N_3120,N_2745);
nor U4893 (N_4893,N_3409,N_2254);
or U4894 (N_4894,N_2543,N_2932);
nand U4895 (N_4895,N_3117,N_3128);
nand U4896 (N_4896,N_2850,N_3710);
or U4897 (N_4897,N_3072,N_2493);
nor U4898 (N_4898,N_2538,N_3923);
nor U4899 (N_4899,N_2353,N_3630);
and U4900 (N_4900,N_3048,N_2225);
nor U4901 (N_4901,N_3506,N_2420);
nand U4902 (N_4902,N_2341,N_2840);
or U4903 (N_4903,N_3173,N_2531);
nor U4904 (N_4904,N_2485,N_2615);
nand U4905 (N_4905,N_3700,N_3802);
or U4906 (N_4906,N_3925,N_3833);
xor U4907 (N_4907,N_3917,N_2632);
or U4908 (N_4908,N_3949,N_2396);
and U4909 (N_4909,N_3937,N_2226);
or U4910 (N_4910,N_3792,N_3836);
and U4911 (N_4911,N_2778,N_3070);
and U4912 (N_4912,N_2348,N_3646);
nand U4913 (N_4913,N_2356,N_2469);
and U4914 (N_4914,N_3933,N_3332);
and U4915 (N_4915,N_2938,N_2930);
nand U4916 (N_4916,N_2398,N_3212);
nor U4917 (N_4917,N_3056,N_3061);
and U4918 (N_4918,N_2207,N_2235);
xnor U4919 (N_4919,N_3139,N_3348);
or U4920 (N_4920,N_2322,N_3898);
nand U4921 (N_4921,N_2642,N_3858);
and U4922 (N_4922,N_2155,N_3392);
nand U4923 (N_4923,N_3080,N_3570);
and U4924 (N_4924,N_3132,N_2665);
nand U4925 (N_4925,N_3872,N_2927);
nand U4926 (N_4926,N_2425,N_2161);
nor U4927 (N_4927,N_3821,N_3962);
nor U4928 (N_4928,N_3204,N_3815);
and U4929 (N_4929,N_2503,N_2139);
nand U4930 (N_4930,N_2402,N_3665);
or U4931 (N_4931,N_3675,N_3022);
nand U4932 (N_4932,N_2475,N_3615);
and U4933 (N_4933,N_3175,N_3505);
or U4934 (N_4934,N_2594,N_3301);
and U4935 (N_4935,N_3755,N_2288);
or U4936 (N_4936,N_3284,N_2640);
and U4937 (N_4937,N_3055,N_3579);
nand U4938 (N_4938,N_3847,N_2054);
nor U4939 (N_4939,N_3235,N_2582);
and U4940 (N_4940,N_3572,N_3756);
or U4941 (N_4941,N_2134,N_3449);
nor U4942 (N_4942,N_3213,N_3485);
nor U4943 (N_4943,N_2506,N_2119);
xor U4944 (N_4944,N_2920,N_2611);
or U4945 (N_4945,N_2421,N_3377);
or U4946 (N_4946,N_3382,N_2083);
nor U4947 (N_4947,N_2826,N_3005);
or U4948 (N_4948,N_3370,N_2742);
nand U4949 (N_4949,N_2203,N_2318);
nor U4950 (N_4950,N_3169,N_2926);
or U4951 (N_4951,N_3960,N_2143);
or U4952 (N_4952,N_3866,N_2411);
and U4953 (N_4953,N_2264,N_3327);
nor U4954 (N_4954,N_2246,N_3564);
nand U4955 (N_4955,N_3845,N_2213);
or U4956 (N_4956,N_3726,N_2287);
xnor U4957 (N_4957,N_3598,N_3265);
nand U4958 (N_4958,N_2857,N_3497);
and U4959 (N_4959,N_3011,N_3686);
nand U4960 (N_4960,N_3245,N_2267);
nor U4961 (N_4961,N_2096,N_2296);
nand U4962 (N_4962,N_3176,N_3848);
or U4963 (N_4963,N_2342,N_2027);
and U4964 (N_4964,N_3764,N_2465);
or U4965 (N_4965,N_2390,N_2737);
or U4966 (N_4966,N_3135,N_2364);
or U4967 (N_4967,N_2973,N_3737);
and U4968 (N_4968,N_2968,N_2070);
or U4969 (N_4969,N_2477,N_3951);
nor U4970 (N_4970,N_2817,N_3118);
and U4971 (N_4971,N_3112,N_2801);
and U4972 (N_4972,N_2137,N_2994);
nand U4973 (N_4973,N_3908,N_2466);
or U4974 (N_4974,N_2660,N_3835);
and U4975 (N_4975,N_3490,N_2010);
and U4976 (N_4976,N_2715,N_2586);
and U4977 (N_4977,N_3328,N_3484);
or U4978 (N_4978,N_3762,N_2311);
nand U4979 (N_4979,N_2861,N_2281);
or U4980 (N_4980,N_2875,N_3249);
nor U4981 (N_4981,N_3420,N_3154);
and U4982 (N_4982,N_3625,N_3068);
and U4983 (N_4983,N_3498,N_3104);
and U4984 (N_4984,N_2698,N_2718);
nor U4985 (N_4985,N_3520,N_3350);
and U4986 (N_4986,N_2459,N_3747);
or U4987 (N_4987,N_3576,N_2655);
nand U4988 (N_4988,N_3513,N_2849);
nand U4989 (N_4989,N_3793,N_2562);
nor U4990 (N_4990,N_3274,N_2216);
nor U4991 (N_4991,N_3107,N_3652);
nand U4992 (N_4992,N_2189,N_2721);
and U4993 (N_4993,N_3681,N_2578);
nand U4994 (N_4994,N_2178,N_2569);
nor U4995 (N_4995,N_2323,N_3543);
nand U4996 (N_4996,N_3226,N_3717);
nor U4997 (N_4997,N_3191,N_2959);
nor U4998 (N_4998,N_2736,N_3785);
and U4999 (N_4999,N_3849,N_3624);
or U5000 (N_5000,N_3579,N_3950);
or U5001 (N_5001,N_2580,N_2953);
or U5002 (N_5002,N_2271,N_2193);
or U5003 (N_5003,N_3160,N_3894);
nand U5004 (N_5004,N_3393,N_3379);
nand U5005 (N_5005,N_2465,N_3036);
and U5006 (N_5006,N_3917,N_2272);
and U5007 (N_5007,N_2455,N_2825);
nand U5008 (N_5008,N_2843,N_2957);
nor U5009 (N_5009,N_2763,N_2865);
nand U5010 (N_5010,N_2214,N_3309);
nor U5011 (N_5011,N_2794,N_3880);
nor U5012 (N_5012,N_2550,N_3689);
and U5013 (N_5013,N_3273,N_3912);
nand U5014 (N_5014,N_3710,N_3030);
nor U5015 (N_5015,N_2422,N_3186);
nand U5016 (N_5016,N_3117,N_3699);
nor U5017 (N_5017,N_2633,N_3450);
or U5018 (N_5018,N_2240,N_3622);
or U5019 (N_5019,N_3797,N_2784);
nor U5020 (N_5020,N_3254,N_2747);
or U5021 (N_5021,N_3054,N_3435);
xnor U5022 (N_5022,N_3333,N_3423);
nand U5023 (N_5023,N_3883,N_3500);
or U5024 (N_5024,N_3925,N_2412);
or U5025 (N_5025,N_3762,N_2456);
and U5026 (N_5026,N_3348,N_2519);
or U5027 (N_5027,N_3713,N_3859);
nand U5028 (N_5028,N_3037,N_2208);
or U5029 (N_5029,N_2255,N_3960);
or U5030 (N_5030,N_2115,N_3107);
xnor U5031 (N_5031,N_3772,N_2873);
or U5032 (N_5032,N_3279,N_3730);
or U5033 (N_5033,N_3980,N_3594);
nor U5034 (N_5034,N_2712,N_2521);
nor U5035 (N_5035,N_3731,N_3884);
or U5036 (N_5036,N_2186,N_3707);
nor U5037 (N_5037,N_3014,N_3781);
or U5038 (N_5038,N_2676,N_2159);
and U5039 (N_5039,N_2441,N_3162);
and U5040 (N_5040,N_2533,N_3376);
and U5041 (N_5041,N_3272,N_2571);
nand U5042 (N_5042,N_3814,N_3424);
nor U5043 (N_5043,N_3397,N_2297);
or U5044 (N_5044,N_3337,N_3274);
and U5045 (N_5045,N_3448,N_2703);
and U5046 (N_5046,N_2799,N_2669);
or U5047 (N_5047,N_2911,N_3711);
nand U5048 (N_5048,N_3002,N_2138);
nor U5049 (N_5049,N_2746,N_2295);
or U5050 (N_5050,N_3654,N_3291);
or U5051 (N_5051,N_3547,N_2159);
nand U5052 (N_5052,N_2954,N_2293);
and U5053 (N_5053,N_2001,N_3173);
nor U5054 (N_5054,N_3653,N_3770);
and U5055 (N_5055,N_2867,N_2699);
and U5056 (N_5056,N_3040,N_2744);
nor U5057 (N_5057,N_2940,N_3858);
nor U5058 (N_5058,N_2947,N_3940);
nand U5059 (N_5059,N_3895,N_2039);
and U5060 (N_5060,N_2186,N_3433);
nand U5061 (N_5061,N_3894,N_3685);
and U5062 (N_5062,N_2370,N_2393);
or U5063 (N_5063,N_3772,N_3085);
or U5064 (N_5064,N_2856,N_3470);
and U5065 (N_5065,N_2890,N_2086);
or U5066 (N_5066,N_2272,N_2456);
and U5067 (N_5067,N_3038,N_3380);
nand U5068 (N_5068,N_2784,N_2652);
or U5069 (N_5069,N_2948,N_3855);
nor U5070 (N_5070,N_2178,N_2089);
xor U5071 (N_5071,N_2817,N_2765);
nor U5072 (N_5072,N_2780,N_2510);
or U5073 (N_5073,N_2161,N_2576);
and U5074 (N_5074,N_2296,N_2174);
nor U5075 (N_5075,N_3015,N_3910);
or U5076 (N_5076,N_3201,N_2665);
nor U5077 (N_5077,N_3946,N_2577);
and U5078 (N_5078,N_3215,N_2568);
nand U5079 (N_5079,N_2825,N_3443);
nand U5080 (N_5080,N_2313,N_3095);
nand U5081 (N_5081,N_2032,N_2549);
nand U5082 (N_5082,N_2239,N_2700);
or U5083 (N_5083,N_2761,N_3967);
or U5084 (N_5084,N_3720,N_2252);
and U5085 (N_5085,N_2774,N_3420);
or U5086 (N_5086,N_3744,N_3311);
nor U5087 (N_5087,N_3722,N_2309);
nand U5088 (N_5088,N_2613,N_2863);
nor U5089 (N_5089,N_3979,N_3333);
nor U5090 (N_5090,N_2989,N_2585);
or U5091 (N_5091,N_3950,N_2344);
and U5092 (N_5092,N_3845,N_2743);
nand U5093 (N_5093,N_2183,N_2404);
and U5094 (N_5094,N_2211,N_2925);
and U5095 (N_5095,N_3900,N_3599);
nand U5096 (N_5096,N_3538,N_3036);
nor U5097 (N_5097,N_3292,N_2437);
or U5098 (N_5098,N_3994,N_3084);
nand U5099 (N_5099,N_2450,N_2524);
nor U5100 (N_5100,N_3599,N_3624);
nor U5101 (N_5101,N_3928,N_3707);
nor U5102 (N_5102,N_2874,N_2700);
and U5103 (N_5103,N_3470,N_2702);
and U5104 (N_5104,N_3717,N_2791);
and U5105 (N_5105,N_2869,N_2377);
and U5106 (N_5106,N_2714,N_2227);
nand U5107 (N_5107,N_2871,N_2158);
nand U5108 (N_5108,N_2012,N_2389);
and U5109 (N_5109,N_2652,N_3758);
nand U5110 (N_5110,N_2866,N_3147);
nor U5111 (N_5111,N_3551,N_3949);
and U5112 (N_5112,N_3196,N_2182);
or U5113 (N_5113,N_3796,N_2487);
and U5114 (N_5114,N_2487,N_2406);
or U5115 (N_5115,N_2967,N_3305);
nand U5116 (N_5116,N_2176,N_2097);
or U5117 (N_5117,N_3513,N_3920);
nand U5118 (N_5118,N_3215,N_3372);
and U5119 (N_5119,N_2188,N_2144);
nand U5120 (N_5120,N_2329,N_3229);
or U5121 (N_5121,N_2507,N_2991);
and U5122 (N_5122,N_3949,N_3707);
or U5123 (N_5123,N_3587,N_2431);
nand U5124 (N_5124,N_3390,N_2218);
nand U5125 (N_5125,N_2382,N_3435);
or U5126 (N_5126,N_2688,N_2118);
nor U5127 (N_5127,N_2724,N_3162);
nand U5128 (N_5128,N_2051,N_2389);
and U5129 (N_5129,N_2789,N_2837);
nor U5130 (N_5130,N_2360,N_2274);
or U5131 (N_5131,N_2782,N_3383);
nand U5132 (N_5132,N_3704,N_2848);
or U5133 (N_5133,N_3438,N_3344);
nor U5134 (N_5134,N_2866,N_3288);
and U5135 (N_5135,N_3927,N_3409);
or U5136 (N_5136,N_3741,N_2483);
nand U5137 (N_5137,N_2047,N_2799);
nor U5138 (N_5138,N_3031,N_3847);
or U5139 (N_5139,N_2175,N_3760);
nand U5140 (N_5140,N_2838,N_2712);
nor U5141 (N_5141,N_3616,N_3682);
and U5142 (N_5142,N_2104,N_3096);
or U5143 (N_5143,N_2909,N_3531);
or U5144 (N_5144,N_2300,N_3972);
or U5145 (N_5145,N_3328,N_3186);
or U5146 (N_5146,N_3944,N_2262);
nor U5147 (N_5147,N_3962,N_2686);
or U5148 (N_5148,N_3671,N_3174);
nor U5149 (N_5149,N_2026,N_2470);
nand U5150 (N_5150,N_3208,N_3929);
and U5151 (N_5151,N_2607,N_3270);
nand U5152 (N_5152,N_2724,N_3312);
and U5153 (N_5153,N_2997,N_2965);
or U5154 (N_5154,N_3149,N_2398);
or U5155 (N_5155,N_2982,N_2904);
nor U5156 (N_5156,N_2978,N_3739);
and U5157 (N_5157,N_3668,N_3842);
nand U5158 (N_5158,N_2977,N_2276);
nor U5159 (N_5159,N_2721,N_2524);
and U5160 (N_5160,N_3880,N_2724);
xor U5161 (N_5161,N_3199,N_2858);
nor U5162 (N_5162,N_3485,N_3475);
nand U5163 (N_5163,N_3694,N_3520);
nand U5164 (N_5164,N_3677,N_2281);
or U5165 (N_5165,N_3791,N_2541);
or U5166 (N_5166,N_2587,N_2358);
nor U5167 (N_5167,N_3201,N_2331);
nand U5168 (N_5168,N_3285,N_3889);
and U5169 (N_5169,N_2553,N_3403);
nand U5170 (N_5170,N_2643,N_3774);
nand U5171 (N_5171,N_3675,N_2223);
nand U5172 (N_5172,N_3266,N_3848);
or U5173 (N_5173,N_3119,N_3762);
or U5174 (N_5174,N_3465,N_3598);
or U5175 (N_5175,N_3715,N_2745);
nor U5176 (N_5176,N_2405,N_3107);
and U5177 (N_5177,N_3741,N_2983);
xnor U5178 (N_5178,N_2279,N_2519);
nor U5179 (N_5179,N_3642,N_2792);
and U5180 (N_5180,N_3912,N_2378);
and U5181 (N_5181,N_3082,N_3952);
or U5182 (N_5182,N_3147,N_2935);
and U5183 (N_5183,N_3573,N_3788);
nand U5184 (N_5184,N_2761,N_3120);
nand U5185 (N_5185,N_3473,N_2169);
nand U5186 (N_5186,N_3885,N_3041);
nor U5187 (N_5187,N_3475,N_2499);
or U5188 (N_5188,N_2116,N_2622);
nand U5189 (N_5189,N_3705,N_3156);
nand U5190 (N_5190,N_2172,N_2037);
and U5191 (N_5191,N_3548,N_2963);
nand U5192 (N_5192,N_3219,N_3853);
nor U5193 (N_5193,N_3016,N_3195);
nor U5194 (N_5194,N_2336,N_3661);
nor U5195 (N_5195,N_3762,N_3180);
nor U5196 (N_5196,N_3922,N_3602);
and U5197 (N_5197,N_3759,N_2665);
or U5198 (N_5198,N_3121,N_3190);
nor U5199 (N_5199,N_2589,N_3308);
nor U5200 (N_5200,N_2198,N_3076);
or U5201 (N_5201,N_2325,N_2872);
or U5202 (N_5202,N_2229,N_2180);
and U5203 (N_5203,N_2436,N_3816);
nand U5204 (N_5204,N_3490,N_3360);
and U5205 (N_5205,N_2480,N_3193);
nor U5206 (N_5206,N_2337,N_2360);
and U5207 (N_5207,N_2451,N_2399);
or U5208 (N_5208,N_2905,N_2682);
nand U5209 (N_5209,N_2948,N_3232);
xnor U5210 (N_5210,N_2848,N_2372);
and U5211 (N_5211,N_2465,N_2667);
nor U5212 (N_5212,N_3717,N_2836);
nor U5213 (N_5213,N_3729,N_3850);
xnor U5214 (N_5214,N_2797,N_2495);
or U5215 (N_5215,N_3905,N_3448);
and U5216 (N_5216,N_3459,N_2343);
nor U5217 (N_5217,N_2109,N_3718);
and U5218 (N_5218,N_3479,N_2402);
or U5219 (N_5219,N_2782,N_2698);
nor U5220 (N_5220,N_2486,N_3819);
nor U5221 (N_5221,N_2152,N_2138);
nand U5222 (N_5222,N_3957,N_2539);
and U5223 (N_5223,N_3643,N_3199);
and U5224 (N_5224,N_3715,N_2487);
nor U5225 (N_5225,N_2412,N_2902);
and U5226 (N_5226,N_3115,N_2682);
nand U5227 (N_5227,N_2574,N_2693);
nand U5228 (N_5228,N_2302,N_2370);
nor U5229 (N_5229,N_3337,N_2755);
nand U5230 (N_5230,N_2078,N_2477);
nand U5231 (N_5231,N_2850,N_3986);
nor U5232 (N_5232,N_2593,N_3410);
or U5233 (N_5233,N_2025,N_3282);
and U5234 (N_5234,N_2404,N_3335);
nand U5235 (N_5235,N_3335,N_3282);
nor U5236 (N_5236,N_2311,N_2371);
and U5237 (N_5237,N_3311,N_2748);
or U5238 (N_5238,N_2314,N_3714);
nand U5239 (N_5239,N_3544,N_3986);
nand U5240 (N_5240,N_3969,N_3126);
or U5241 (N_5241,N_2370,N_3034);
and U5242 (N_5242,N_3206,N_3175);
or U5243 (N_5243,N_2532,N_2397);
nor U5244 (N_5244,N_3951,N_2595);
nor U5245 (N_5245,N_2396,N_3633);
or U5246 (N_5246,N_2820,N_2547);
or U5247 (N_5247,N_2175,N_2722);
nand U5248 (N_5248,N_3403,N_2224);
and U5249 (N_5249,N_2538,N_3344);
or U5250 (N_5250,N_3214,N_2694);
nand U5251 (N_5251,N_2531,N_3872);
or U5252 (N_5252,N_2264,N_3311);
nor U5253 (N_5253,N_2917,N_2737);
nand U5254 (N_5254,N_2593,N_3021);
nor U5255 (N_5255,N_2328,N_3100);
nand U5256 (N_5256,N_2789,N_3444);
nand U5257 (N_5257,N_2228,N_3935);
and U5258 (N_5258,N_3263,N_2749);
nor U5259 (N_5259,N_2054,N_2157);
nand U5260 (N_5260,N_3956,N_3512);
nor U5261 (N_5261,N_3638,N_2002);
or U5262 (N_5262,N_2680,N_3289);
and U5263 (N_5263,N_2138,N_2732);
nor U5264 (N_5264,N_3488,N_3639);
nor U5265 (N_5265,N_3037,N_3969);
and U5266 (N_5266,N_3055,N_2338);
and U5267 (N_5267,N_2651,N_2141);
nand U5268 (N_5268,N_2292,N_2020);
nor U5269 (N_5269,N_3598,N_3973);
nand U5270 (N_5270,N_2706,N_3877);
nor U5271 (N_5271,N_2191,N_3418);
nor U5272 (N_5272,N_3755,N_2481);
and U5273 (N_5273,N_2301,N_2481);
nor U5274 (N_5274,N_2624,N_2981);
nand U5275 (N_5275,N_3838,N_3681);
and U5276 (N_5276,N_3685,N_2980);
nand U5277 (N_5277,N_3121,N_2505);
nor U5278 (N_5278,N_2667,N_3023);
and U5279 (N_5279,N_2174,N_3780);
nor U5280 (N_5280,N_2619,N_3313);
or U5281 (N_5281,N_3460,N_2466);
nor U5282 (N_5282,N_2533,N_2098);
nor U5283 (N_5283,N_3982,N_2662);
or U5284 (N_5284,N_2794,N_3840);
nand U5285 (N_5285,N_2028,N_2736);
nand U5286 (N_5286,N_2710,N_2682);
nand U5287 (N_5287,N_2679,N_3566);
nand U5288 (N_5288,N_3516,N_2015);
nor U5289 (N_5289,N_3855,N_3938);
nor U5290 (N_5290,N_2965,N_3490);
nand U5291 (N_5291,N_3196,N_3348);
nand U5292 (N_5292,N_2273,N_3314);
nor U5293 (N_5293,N_2074,N_2152);
and U5294 (N_5294,N_3900,N_2347);
or U5295 (N_5295,N_3884,N_3369);
or U5296 (N_5296,N_2850,N_3263);
or U5297 (N_5297,N_3103,N_3816);
and U5298 (N_5298,N_3358,N_2432);
nor U5299 (N_5299,N_3517,N_2498);
nor U5300 (N_5300,N_3045,N_2798);
nand U5301 (N_5301,N_3477,N_3000);
nand U5302 (N_5302,N_3472,N_3860);
nor U5303 (N_5303,N_3698,N_2153);
nor U5304 (N_5304,N_2438,N_2451);
and U5305 (N_5305,N_2384,N_2859);
nand U5306 (N_5306,N_2669,N_3913);
or U5307 (N_5307,N_3673,N_2786);
nor U5308 (N_5308,N_2455,N_3350);
nand U5309 (N_5309,N_3225,N_2032);
and U5310 (N_5310,N_3723,N_2806);
or U5311 (N_5311,N_2773,N_2104);
or U5312 (N_5312,N_3503,N_3587);
nand U5313 (N_5313,N_3799,N_3395);
or U5314 (N_5314,N_3050,N_2193);
nand U5315 (N_5315,N_2342,N_2207);
or U5316 (N_5316,N_2722,N_2356);
or U5317 (N_5317,N_2271,N_3381);
and U5318 (N_5318,N_3082,N_2768);
nor U5319 (N_5319,N_2184,N_3493);
xnor U5320 (N_5320,N_2206,N_3446);
and U5321 (N_5321,N_2711,N_2961);
nor U5322 (N_5322,N_3655,N_2653);
nor U5323 (N_5323,N_3973,N_3143);
and U5324 (N_5324,N_3778,N_3697);
and U5325 (N_5325,N_2930,N_2142);
or U5326 (N_5326,N_2524,N_2851);
xor U5327 (N_5327,N_3821,N_3031);
nand U5328 (N_5328,N_3473,N_3870);
and U5329 (N_5329,N_3978,N_3329);
or U5330 (N_5330,N_2943,N_2778);
and U5331 (N_5331,N_3391,N_2423);
nand U5332 (N_5332,N_2236,N_2270);
xnor U5333 (N_5333,N_2780,N_2352);
and U5334 (N_5334,N_2411,N_3480);
nor U5335 (N_5335,N_2392,N_3363);
and U5336 (N_5336,N_3032,N_3551);
nor U5337 (N_5337,N_2459,N_2331);
or U5338 (N_5338,N_2544,N_3783);
and U5339 (N_5339,N_3378,N_2924);
nand U5340 (N_5340,N_3155,N_2355);
and U5341 (N_5341,N_2551,N_2509);
nand U5342 (N_5342,N_2577,N_3229);
and U5343 (N_5343,N_3734,N_3406);
or U5344 (N_5344,N_3652,N_2581);
nand U5345 (N_5345,N_2533,N_2715);
nor U5346 (N_5346,N_2039,N_2362);
or U5347 (N_5347,N_3224,N_3588);
nor U5348 (N_5348,N_2766,N_2171);
or U5349 (N_5349,N_3304,N_2811);
and U5350 (N_5350,N_2383,N_3836);
nor U5351 (N_5351,N_3354,N_2314);
nor U5352 (N_5352,N_3211,N_3740);
nand U5353 (N_5353,N_2093,N_3987);
nand U5354 (N_5354,N_3829,N_3630);
nand U5355 (N_5355,N_3717,N_2512);
nor U5356 (N_5356,N_2032,N_3602);
or U5357 (N_5357,N_2865,N_3356);
nand U5358 (N_5358,N_2069,N_3736);
or U5359 (N_5359,N_3198,N_3044);
nor U5360 (N_5360,N_3388,N_2144);
or U5361 (N_5361,N_3814,N_2439);
and U5362 (N_5362,N_3318,N_3368);
and U5363 (N_5363,N_3506,N_3817);
nand U5364 (N_5364,N_3392,N_2256);
xor U5365 (N_5365,N_2815,N_2888);
nand U5366 (N_5366,N_3454,N_3914);
or U5367 (N_5367,N_2308,N_3820);
nor U5368 (N_5368,N_3924,N_3860);
nand U5369 (N_5369,N_3212,N_3078);
nor U5370 (N_5370,N_2245,N_2429);
nor U5371 (N_5371,N_3689,N_2259);
nand U5372 (N_5372,N_2970,N_2905);
or U5373 (N_5373,N_2882,N_2985);
and U5374 (N_5374,N_3365,N_2986);
or U5375 (N_5375,N_3494,N_3338);
or U5376 (N_5376,N_2759,N_2524);
or U5377 (N_5377,N_3149,N_2215);
and U5378 (N_5378,N_3566,N_3431);
or U5379 (N_5379,N_3112,N_3718);
and U5380 (N_5380,N_2490,N_2798);
nor U5381 (N_5381,N_3798,N_3584);
or U5382 (N_5382,N_3892,N_2625);
nand U5383 (N_5383,N_2414,N_2199);
nand U5384 (N_5384,N_2250,N_2420);
and U5385 (N_5385,N_3946,N_3386);
xnor U5386 (N_5386,N_2622,N_3589);
nor U5387 (N_5387,N_2023,N_2406);
or U5388 (N_5388,N_2123,N_3394);
and U5389 (N_5389,N_3189,N_2223);
or U5390 (N_5390,N_2086,N_2401);
or U5391 (N_5391,N_3320,N_3769);
or U5392 (N_5392,N_3837,N_2536);
or U5393 (N_5393,N_3444,N_3910);
and U5394 (N_5394,N_2809,N_2303);
or U5395 (N_5395,N_3495,N_2047);
and U5396 (N_5396,N_2017,N_3726);
nand U5397 (N_5397,N_3954,N_2681);
nand U5398 (N_5398,N_3655,N_3018);
nor U5399 (N_5399,N_3988,N_3529);
or U5400 (N_5400,N_3612,N_2822);
and U5401 (N_5401,N_3424,N_3053);
and U5402 (N_5402,N_2799,N_3704);
or U5403 (N_5403,N_3957,N_2806);
or U5404 (N_5404,N_3105,N_3049);
nand U5405 (N_5405,N_3218,N_3255);
nor U5406 (N_5406,N_2973,N_3328);
or U5407 (N_5407,N_3072,N_2153);
nand U5408 (N_5408,N_2193,N_2386);
nand U5409 (N_5409,N_3060,N_2415);
and U5410 (N_5410,N_3626,N_3667);
and U5411 (N_5411,N_3463,N_2608);
nand U5412 (N_5412,N_2993,N_2715);
nand U5413 (N_5413,N_3119,N_3761);
and U5414 (N_5414,N_2106,N_3278);
or U5415 (N_5415,N_3541,N_3606);
nor U5416 (N_5416,N_2515,N_3853);
nor U5417 (N_5417,N_3066,N_2833);
and U5418 (N_5418,N_2392,N_3205);
nand U5419 (N_5419,N_3580,N_3811);
nor U5420 (N_5420,N_2307,N_2483);
and U5421 (N_5421,N_3129,N_3820);
nor U5422 (N_5422,N_3558,N_2201);
nor U5423 (N_5423,N_2755,N_2977);
nand U5424 (N_5424,N_3036,N_2639);
nand U5425 (N_5425,N_3831,N_3457);
nor U5426 (N_5426,N_3890,N_2018);
nand U5427 (N_5427,N_2485,N_3173);
nor U5428 (N_5428,N_3302,N_3406);
or U5429 (N_5429,N_2527,N_3845);
nand U5430 (N_5430,N_2649,N_3449);
nor U5431 (N_5431,N_3185,N_2255);
or U5432 (N_5432,N_2946,N_2005);
or U5433 (N_5433,N_3639,N_3417);
and U5434 (N_5434,N_3564,N_3870);
or U5435 (N_5435,N_3489,N_2895);
nand U5436 (N_5436,N_3579,N_2443);
nand U5437 (N_5437,N_3731,N_3703);
and U5438 (N_5438,N_3991,N_3598);
nor U5439 (N_5439,N_3256,N_2050);
and U5440 (N_5440,N_2352,N_3381);
nor U5441 (N_5441,N_2540,N_3788);
nor U5442 (N_5442,N_3500,N_2008);
nor U5443 (N_5443,N_3427,N_3209);
and U5444 (N_5444,N_2689,N_3389);
nand U5445 (N_5445,N_2614,N_2676);
nand U5446 (N_5446,N_2834,N_2680);
nor U5447 (N_5447,N_3824,N_2694);
nand U5448 (N_5448,N_2789,N_2449);
nand U5449 (N_5449,N_2451,N_3729);
or U5450 (N_5450,N_3157,N_2949);
or U5451 (N_5451,N_3468,N_2599);
or U5452 (N_5452,N_3820,N_3885);
nor U5453 (N_5453,N_3271,N_2636);
or U5454 (N_5454,N_2711,N_2624);
nor U5455 (N_5455,N_3049,N_2463);
xnor U5456 (N_5456,N_2943,N_3596);
nand U5457 (N_5457,N_3367,N_2051);
or U5458 (N_5458,N_2501,N_2811);
or U5459 (N_5459,N_3303,N_3744);
and U5460 (N_5460,N_3020,N_3804);
and U5461 (N_5461,N_2791,N_2835);
and U5462 (N_5462,N_2249,N_2046);
and U5463 (N_5463,N_2313,N_3968);
nor U5464 (N_5464,N_3612,N_3180);
or U5465 (N_5465,N_3426,N_2850);
or U5466 (N_5466,N_2544,N_2091);
nor U5467 (N_5467,N_2514,N_2421);
or U5468 (N_5468,N_3717,N_3974);
nand U5469 (N_5469,N_3247,N_2788);
nor U5470 (N_5470,N_2309,N_3755);
nand U5471 (N_5471,N_2905,N_2425);
and U5472 (N_5472,N_2306,N_3987);
or U5473 (N_5473,N_3141,N_3799);
nand U5474 (N_5474,N_2747,N_3601);
nand U5475 (N_5475,N_3849,N_2043);
and U5476 (N_5476,N_2394,N_3569);
nor U5477 (N_5477,N_2123,N_3676);
nand U5478 (N_5478,N_3856,N_3036);
and U5479 (N_5479,N_2342,N_2620);
nor U5480 (N_5480,N_2315,N_2304);
and U5481 (N_5481,N_3327,N_2912);
nand U5482 (N_5482,N_3933,N_3129);
nand U5483 (N_5483,N_3980,N_3000);
nand U5484 (N_5484,N_3486,N_3775);
nor U5485 (N_5485,N_2158,N_3732);
nand U5486 (N_5486,N_3506,N_2719);
and U5487 (N_5487,N_3666,N_2921);
nand U5488 (N_5488,N_2221,N_2385);
nand U5489 (N_5489,N_3208,N_3391);
nor U5490 (N_5490,N_2126,N_2033);
nor U5491 (N_5491,N_3915,N_2046);
nor U5492 (N_5492,N_2859,N_3688);
and U5493 (N_5493,N_3039,N_3435);
nor U5494 (N_5494,N_2756,N_3957);
and U5495 (N_5495,N_2721,N_2702);
and U5496 (N_5496,N_2397,N_3657);
and U5497 (N_5497,N_3803,N_2495);
and U5498 (N_5498,N_3227,N_2196);
nor U5499 (N_5499,N_3956,N_2701);
and U5500 (N_5500,N_2126,N_3545);
or U5501 (N_5501,N_3616,N_3113);
or U5502 (N_5502,N_2796,N_2379);
nor U5503 (N_5503,N_2752,N_2464);
or U5504 (N_5504,N_3613,N_3405);
or U5505 (N_5505,N_3217,N_2615);
and U5506 (N_5506,N_2474,N_2033);
and U5507 (N_5507,N_3295,N_2016);
nor U5508 (N_5508,N_3264,N_2988);
and U5509 (N_5509,N_3451,N_2339);
or U5510 (N_5510,N_2100,N_2526);
or U5511 (N_5511,N_3153,N_3121);
and U5512 (N_5512,N_3821,N_2656);
or U5513 (N_5513,N_2187,N_3014);
nor U5514 (N_5514,N_3811,N_2244);
nand U5515 (N_5515,N_2385,N_3741);
and U5516 (N_5516,N_2765,N_3887);
and U5517 (N_5517,N_3585,N_2167);
or U5518 (N_5518,N_2903,N_2217);
and U5519 (N_5519,N_3059,N_2420);
nand U5520 (N_5520,N_3334,N_2289);
or U5521 (N_5521,N_3741,N_3297);
or U5522 (N_5522,N_3217,N_3449);
nor U5523 (N_5523,N_2212,N_3347);
nor U5524 (N_5524,N_2764,N_3679);
nand U5525 (N_5525,N_2481,N_2653);
and U5526 (N_5526,N_2053,N_3741);
nor U5527 (N_5527,N_3103,N_3704);
nand U5528 (N_5528,N_3832,N_3532);
and U5529 (N_5529,N_3785,N_3432);
and U5530 (N_5530,N_3548,N_3991);
and U5531 (N_5531,N_2456,N_3591);
or U5532 (N_5532,N_3734,N_2203);
xnor U5533 (N_5533,N_2217,N_3761);
and U5534 (N_5534,N_3679,N_3862);
nand U5535 (N_5535,N_3778,N_3957);
and U5536 (N_5536,N_3434,N_2261);
nand U5537 (N_5537,N_2317,N_3260);
nand U5538 (N_5538,N_2710,N_2520);
and U5539 (N_5539,N_3142,N_3445);
and U5540 (N_5540,N_2070,N_2311);
nand U5541 (N_5541,N_3743,N_3274);
nand U5542 (N_5542,N_3241,N_3020);
and U5543 (N_5543,N_3053,N_2044);
or U5544 (N_5544,N_3038,N_2067);
and U5545 (N_5545,N_2326,N_3802);
nor U5546 (N_5546,N_2766,N_2796);
or U5547 (N_5547,N_2768,N_2776);
and U5548 (N_5548,N_2634,N_3720);
nor U5549 (N_5549,N_3591,N_3352);
nand U5550 (N_5550,N_2410,N_3736);
and U5551 (N_5551,N_3531,N_3368);
or U5552 (N_5552,N_3212,N_3857);
and U5553 (N_5553,N_3262,N_2035);
or U5554 (N_5554,N_3800,N_3378);
and U5555 (N_5555,N_3522,N_3820);
nand U5556 (N_5556,N_3388,N_3706);
or U5557 (N_5557,N_2755,N_2945);
nand U5558 (N_5558,N_2837,N_3854);
or U5559 (N_5559,N_3865,N_3845);
and U5560 (N_5560,N_2523,N_2245);
nand U5561 (N_5561,N_2321,N_2916);
xor U5562 (N_5562,N_2865,N_2045);
nor U5563 (N_5563,N_2391,N_3771);
nand U5564 (N_5564,N_2342,N_3180);
nor U5565 (N_5565,N_2541,N_2850);
or U5566 (N_5566,N_2062,N_2705);
nand U5567 (N_5567,N_2717,N_2507);
or U5568 (N_5568,N_3155,N_3048);
or U5569 (N_5569,N_2363,N_3538);
nand U5570 (N_5570,N_3811,N_3428);
and U5571 (N_5571,N_2452,N_3079);
nand U5572 (N_5572,N_3740,N_3496);
nand U5573 (N_5573,N_3933,N_2885);
nor U5574 (N_5574,N_2340,N_3460);
nand U5575 (N_5575,N_2477,N_2866);
nor U5576 (N_5576,N_3589,N_2115);
nand U5577 (N_5577,N_2167,N_3664);
nor U5578 (N_5578,N_3299,N_2936);
or U5579 (N_5579,N_2984,N_3980);
and U5580 (N_5580,N_3265,N_2770);
nand U5581 (N_5581,N_2913,N_2524);
nand U5582 (N_5582,N_2816,N_2132);
and U5583 (N_5583,N_2656,N_2030);
and U5584 (N_5584,N_2994,N_3193);
nand U5585 (N_5585,N_3160,N_3029);
and U5586 (N_5586,N_2523,N_2429);
nor U5587 (N_5587,N_3697,N_3093);
or U5588 (N_5588,N_2906,N_2190);
nor U5589 (N_5589,N_3138,N_2191);
nand U5590 (N_5590,N_2741,N_3145);
nand U5591 (N_5591,N_2599,N_3903);
or U5592 (N_5592,N_2914,N_2361);
or U5593 (N_5593,N_2709,N_3670);
nand U5594 (N_5594,N_3208,N_3156);
and U5595 (N_5595,N_2596,N_3660);
nand U5596 (N_5596,N_2488,N_3009);
or U5597 (N_5597,N_2431,N_3801);
or U5598 (N_5598,N_2978,N_2967);
and U5599 (N_5599,N_2464,N_3919);
or U5600 (N_5600,N_3026,N_2786);
xnor U5601 (N_5601,N_2899,N_3941);
or U5602 (N_5602,N_3757,N_3176);
and U5603 (N_5603,N_3440,N_3580);
and U5604 (N_5604,N_3993,N_3551);
or U5605 (N_5605,N_2100,N_3894);
or U5606 (N_5606,N_2834,N_2456);
and U5607 (N_5607,N_3782,N_2745);
or U5608 (N_5608,N_3663,N_2576);
or U5609 (N_5609,N_2924,N_3737);
and U5610 (N_5610,N_2670,N_3591);
or U5611 (N_5611,N_3689,N_3664);
nand U5612 (N_5612,N_2150,N_2905);
nand U5613 (N_5613,N_2056,N_3290);
nor U5614 (N_5614,N_2280,N_2983);
and U5615 (N_5615,N_2771,N_3240);
nand U5616 (N_5616,N_3926,N_2339);
or U5617 (N_5617,N_2387,N_3269);
nand U5618 (N_5618,N_3324,N_3301);
or U5619 (N_5619,N_3829,N_2393);
or U5620 (N_5620,N_3402,N_2563);
and U5621 (N_5621,N_3906,N_2003);
and U5622 (N_5622,N_2417,N_3615);
or U5623 (N_5623,N_3732,N_3917);
and U5624 (N_5624,N_3083,N_2496);
nor U5625 (N_5625,N_3066,N_3381);
nor U5626 (N_5626,N_3469,N_2356);
nor U5627 (N_5627,N_3795,N_2920);
nand U5628 (N_5628,N_2546,N_3836);
and U5629 (N_5629,N_2105,N_2990);
and U5630 (N_5630,N_2923,N_3760);
nand U5631 (N_5631,N_3728,N_3608);
and U5632 (N_5632,N_2165,N_3455);
nor U5633 (N_5633,N_2151,N_3118);
and U5634 (N_5634,N_2629,N_3678);
or U5635 (N_5635,N_3970,N_2510);
nand U5636 (N_5636,N_2966,N_2160);
nand U5637 (N_5637,N_3861,N_2467);
and U5638 (N_5638,N_2896,N_2223);
nand U5639 (N_5639,N_2233,N_3572);
and U5640 (N_5640,N_3116,N_2663);
nor U5641 (N_5641,N_2827,N_3779);
or U5642 (N_5642,N_3445,N_2052);
nor U5643 (N_5643,N_2490,N_3590);
nor U5644 (N_5644,N_3612,N_3395);
and U5645 (N_5645,N_2728,N_3803);
or U5646 (N_5646,N_2147,N_2861);
or U5647 (N_5647,N_3025,N_2405);
nand U5648 (N_5648,N_2486,N_2722);
or U5649 (N_5649,N_3184,N_3101);
nand U5650 (N_5650,N_2216,N_2750);
and U5651 (N_5651,N_3988,N_3170);
and U5652 (N_5652,N_2894,N_2376);
and U5653 (N_5653,N_2096,N_3481);
and U5654 (N_5654,N_3264,N_3870);
or U5655 (N_5655,N_2204,N_2483);
or U5656 (N_5656,N_3794,N_3176);
and U5657 (N_5657,N_3135,N_2969);
nand U5658 (N_5658,N_3634,N_3174);
nor U5659 (N_5659,N_2058,N_2849);
nand U5660 (N_5660,N_3164,N_2031);
nand U5661 (N_5661,N_3438,N_2150);
nor U5662 (N_5662,N_3421,N_3884);
nor U5663 (N_5663,N_2735,N_3510);
or U5664 (N_5664,N_2026,N_3466);
nor U5665 (N_5665,N_2083,N_2422);
or U5666 (N_5666,N_3641,N_3375);
and U5667 (N_5667,N_2952,N_3942);
and U5668 (N_5668,N_2132,N_2642);
or U5669 (N_5669,N_3281,N_2520);
or U5670 (N_5670,N_3385,N_3672);
and U5671 (N_5671,N_3210,N_2789);
or U5672 (N_5672,N_3966,N_3671);
nand U5673 (N_5673,N_2076,N_2868);
nor U5674 (N_5674,N_3366,N_3197);
or U5675 (N_5675,N_3717,N_3086);
nor U5676 (N_5676,N_2794,N_2606);
nor U5677 (N_5677,N_3354,N_2530);
or U5678 (N_5678,N_2053,N_2061);
nand U5679 (N_5679,N_2676,N_3102);
or U5680 (N_5680,N_3604,N_3844);
or U5681 (N_5681,N_2565,N_3677);
nand U5682 (N_5682,N_2775,N_2325);
nand U5683 (N_5683,N_2800,N_2074);
or U5684 (N_5684,N_2569,N_2099);
nor U5685 (N_5685,N_2700,N_2165);
nand U5686 (N_5686,N_2812,N_3078);
and U5687 (N_5687,N_3320,N_2280);
or U5688 (N_5688,N_2092,N_2252);
or U5689 (N_5689,N_2405,N_2299);
or U5690 (N_5690,N_3206,N_3961);
or U5691 (N_5691,N_2288,N_3144);
or U5692 (N_5692,N_2460,N_2866);
nor U5693 (N_5693,N_2399,N_3699);
nor U5694 (N_5694,N_2004,N_3911);
nand U5695 (N_5695,N_3107,N_2208);
and U5696 (N_5696,N_2123,N_3002);
nor U5697 (N_5697,N_2362,N_2942);
nor U5698 (N_5698,N_3916,N_3577);
nor U5699 (N_5699,N_2298,N_3470);
and U5700 (N_5700,N_3538,N_2075);
nor U5701 (N_5701,N_3644,N_3761);
and U5702 (N_5702,N_2178,N_2835);
or U5703 (N_5703,N_3618,N_3994);
and U5704 (N_5704,N_2216,N_2143);
nand U5705 (N_5705,N_2782,N_2675);
and U5706 (N_5706,N_3034,N_3033);
nand U5707 (N_5707,N_2691,N_3477);
nor U5708 (N_5708,N_3014,N_3877);
nand U5709 (N_5709,N_3109,N_2578);
nor U5710 (N_5710,N_3321,N_2534);
or U5711 (N_5711,N_3536,N_2478);
nand U5712 (N_5712,N_2938,N_3557);
and U5713 (N_5713,N_3285,N_3658);
and U5714 (N_5714,N_2294,N_2407);
nor U5715 (N_5715,N_3238,N_3904);
or U5716 (N_5716,N_2585,N_3255);
or U5717 (N_5717,N_3626,N_2628);
and U5718 (N_5718,N_3390,N_2928);
and U5719 (N_5719,N_2066,N_3554);
nor U5720 (N_5720,N_2107,N_3508);
nor U5721 (N_5721,N_2340,N_3772);
nor U5722 (N_5722,N_3201,N_2597);
and U5723 (N_5723,N_2553,N_2782);
and U5724 (N_5724,N_2282,N_2525);
and U5725 (N_5725,N_3415,N_3668);
or U5726 (N_5726,N_3082,N_3574);
nand U5727 (N_5727,N_3485,N_3452);
and U5728 (N_5728,N_2317,N_2060);
or U5729 (N_5729,N_3616,N_2417);
nor U5730 (N_5730,N_3072,N_3851);
xnor U5731 (N_5731,N_3317,N_3746);
nor U5732 (N_5732,N_2196,N_3520);
nand U5733 (N_5733,N_3775,N_2457);
xnor U5734 (N_5734,N_2213,N_3139);
nand U5735 (N_5735,N_2216,N_2310);
or U5736 (N_5736,N_3824,N_2358);
and U5737 (N_5737,N_3820,N_2247);
nand U5738 (N_5738,N_2893,N_2746);
and U5739 (N_5739,N_2747,N_3657);
nor U5740 (N_5740,N_3358,N_3673);
nand U5741 (N_5741,N_2256,N_2668);
nor U5742 (N_5742,N_3903,N_2769);
nor U5743 (N_5743,N_3064,N_3829);
and U5744 (N_5744,N_2821,N_2860);
or U5745 (N_5745,N_3408,N_2309);
nand U5746 (N_5746,N_3718,N_3488);
nand U5747 (N_5747,N_3709,N_3728);
and U5748 (N_5748,N_2691,N_3669);
and U5749 (N_5749,N_2684,N_2137);
and U5750 (N_5750,N_3048,N_2288);
nor U5751 (N_5751,N_3235,N_2270);
nand U5752 (N_5752,N_2351,N_3144);
or U5753 (N_5753,N_2731,N_3686);
and U5754 (N_5754,N_2510,N_3266);
nand U5755 (N_5755,N_2513,N_2733);
or U5756 (N_5756,N_2475,N_3580);
or U5757 (N_5757,N_2266,N_2360);
or U5758 (N_5758,N_3662,N_3835);
nand U5759 (N_5759,N_3806,N_3358);
and U5760 (N_5760,N_2808,N_3272);
nor U5761 (N_5761,N_3037,N_3184);
and U5762 (N_5762,N_2403,N_2456);
nand U5763 (N_5763,N_3105,N_2087);
or U5764 (N_5764,N_2803,N_3727);
and U5765 (N_5765,N_2307,N_3580);
nor U5766 (N_5766,N_3889,N_3980);
and U5767 (N_5767,N_2685,N_3569);
nand U5768 (N_5768,N_3445,N_2200);
nand U5769 (N_5769,N_2580,N_3706);
nor U5770 (N_5770,N_3964,N_3763);
nand U5771 (N_5771,N_3729,N_2466);
nand U5772 (N_5772,N_3773,N_2980);
nor U5773 (N_5773,N_3969,N_2612);
and U5774 (N_5774,N_3033,N_2604);
nand U5775 (N_5775,N_2970,N_2078);
nand U5776 (N_5776,N_2815,N_2757);
and U5777 (N_5777,N_2148,N_3330);
and U5778 (N_5778,N_2673,N_2205);
nand U5779 (N_5779,N_2607,N_3218);
or U5780 (N_5780,N_3288,N_2922);
and U5781 (N_5781,N_3616,N_3666);
nor U5782 (N_5782,N_3059,N_3724);
nand U5783 (N_5783,N_2980,N_3136);
and U5784 (N_5784,N_2213,N_3640);
or U5785 (N_5785,N_2051,N_2870);
nor U5786 (N_5786,N_2174,N_2325);
nand U5787 (N_5787,N_2904,N_3141);
nand U5788 (N_5788,N_3232,N_2900);
nand U5789 (N_5789,N_2610,N_2550);
and U5790 (N_5790,N_3433,N_2112);
or U5791 (N_5791,N_2517,N_2436);
or U5792 (N_5792,N_3795,N_2788);
nand U5793 (N_5793,N_2938,N_3378);
or U5794 (N_5794,N_2583,N_2336);
and U5795 (N_5795,N_2125,N_3086);
nand U5796 (N_5796,N_2113,N_3568);
and U5797 (N_5797,N_2632,N_2327);
and U5798 (N_5798,N_2284,N_2432);
and U5799 (N_5799,N_2895,N_2452);
or U5800 (N_5800,N_2490,N_3710);
and U5801 (N_5801,N_3074,N_2371);
nor U5802 (N_5802,N_3296,N_3111);
nand U5803 (N_5803,N_3128,N_2708);
nand U5804 (N_5804,N_3400,N_3804);
and U5805 (N_5805,N_3411,N_2816);
nor U5806 (N_5806,N_2049,N_2559);
nor U5807 (N_5807,N_2617,N_2812);
or U5808 (N_5808,N_2543,N_2061);
or U5809 (N_5809,N_2115,N_2272);
nor U5810 (N_5810,N_3266,N_3149);
or U5811 (N_5811,N_3914,N_3814);
nor U5812 (N_5812,N_3620,N_3544);
or U5813 (N_5813,N_3678,N_3054);
nor U5814 (N_5814,N_2102,N_3679);
and U5815 (N_5815,N_3795,N_3753);
nor U5816 (N_5816,N_2936,N_2984);
nor U5817 (N_5817,N_2384,N_3577);
and U5818 (N_5818,N_2355,N_3391);
nand U5819 (N_5819,N_2808,N_2642);
nand U5820 (N_5820,N_2765,N_3767);
nor U5821 (N_5821,N_2216,N_2077);
xor U5822 (N_5822,N_3373,N_2582);
nand U5823 (N_5823,N_2561,N_3743);
and U5824 (N_5824,N_3421,N_2636);
or U5825 (N_5825,N_3727,N_2880);
nor U5826 (N_5826,N_2632,N_2868);
nand U5827 (N_5827,N_2155,N_2237);
and U5828 (N_5828,N_3453,N_3171);
or U5829 (N_5829,N_3559,N_3594);
nand U5830 (N_5830,N_3550,N_3504);
nand U5831 (N_5831,N_2049,N_3052);
or U5832 (N_5832,N_2922,N_2269);
and U5833 (N_5833,N_2872,N_3399);
nand U5834 (N_5834,N_2247,N_2182);
and U5835 (N_5835,N_3799,N_3760);
or U5836 (N_5836,N_3388,N_2323);
or U5837 (N_5837,N_2861,N_3252);
and U5838 (N_5838,N_3614,N_2387);
or U5839 (N_5839,N_3948,N_2034);
nand U5840 (N_5840,N_2201,N_3637);
or U5841 (N_5841,N_2283,N_2052);
nor U5842 (N_5842,N_3271,N_2852);
nor U5843 (N_5843,N_3412,N_3779);
nand U5844 (N_5844,N_2079,N_3226);
and U5845 (N_5845,N_2669,N_2596);
nand U5846 (N_5846,N_2513,N_3337);
nand U5847 (N_5847,N_3794,N_3296);
or U5848 (N_5848,N_2312,N_3685);
or U5849 (N_5849,N_2133,N_3526);
or U5850 (N_5850,N_2531,N_2210);
and U5851 (N_5851,N_2023,N_2458);
nor U5852 (N_5852,N_3074,N_3557);
nand U5853 (N_5853,N_3722,N_2936);
and U5854 (N_5854,N_2035,N_2108);
or U5855 (N_5855,N_2385,N_3960);
and U5856 (N_5856,N_3428,N_3241);
and U5857 (N_5857,N_2009,N_2613);
or U5858 (N_5858,N_3414,N_3996);
or U5859 (N_5859,N_2560,N_3620);
nand U5860 (N_5860,N_2248,N_2955);
nand U5861 (N_5861,N_3723,N_2493);
nor U5862 (N_5862,N_3996,N_3454);
or U5863 (N_5863,N_3936,N_3771);
and U5864 (N_5864,N_2404,N_2253);
nor U5865 (N_5865,N_3788,N_3651);
or U5866 (N_5866,N_2985,N_2765);
nand U5867 (N_5867,N_3793,N_2464);
xnor U5868 (N_5868,N_2220,N_3104);
and U5869 (N_5869,N_3875,N_2272);
or U5870 (N_5870,N_2609,N_3952);
nor U5871 (N_5871,N_3678,N_3494);
nor U5872 (N_5872,N_2169,N_3864);
nand U5873 (N_5873,N_2297,N_3840);
or U5874 (N_5874,N_2272,N_3641);
nand U5875 (N_5875,N_3037,N_3089);
nand U5876 (N_5876,N_2158,N_2761);
or U5877 (N_5877,N_2098,N_3674);
nor U5878 (N_5878,N_2493,N_2228);
and U5879 (N_5879,N_2021,N_3333);
and U5880 (N_5880,N_3260,N_2099);
nand U5881 (N_5881,N_2006,N_2851);
nor U5882 (N_5882,N_2282,N_3685);
nor U5883 (N_5883,N_3708,N_3456);
nor U5884 (N_5884,N_3976,N_3219);
and U5885 (N_5885,N_2692,N_2937);
and U5886 (N_5886,N_3817,N_3502);
and U5887 (N_5887,N_2526,N_3752);
nand U5888 (N_5888,N_3361,N_2858);
nor U5889 (N_5889,N_3008,N_2386);
and U5890 (N_5890,N_2103,N_3091);
and U5891 (N_5891,N_3785,N_2762);
nand U5892 (N_5892,N_2365,N_3711);
nand U5893 (N_5893,N_3532,N_2515);
and U5894 (N_5894,N_2842,N_3442);
or U5895 (N_5895,N_3260,N_3381);
nor U5896 (N_5896,N_3235,N_2657);
and U5897 (N_5897,N_3474,N_2714);
and U5898 (N_5898,N_3523,N_2159);
and U5899 (N_5899,N_2713,N_2124);
or U5900 (N_5900,N_3734,N_3930);
nand U5901 (N_5901,N_3914,N_2082);
or U5902 (N_5902,N_2928,N_2082);
or U5903 (N_5903,N_2690,N_2327);
and U5904 (N_5904,N_3925,N_3881);
and U5905 (N_5905,N_2342,N_3947);
nor U5906 (N_5906,N_3463,N_2817);
and U5907 (N_5907,N_2584,N_3369);
nand U5908 (N_5908,N_3863,N_3629);
or U5909 (N_5909,N_3154,N_3604);
nor U5910 (N_5910,N_2099,N_3673);
nand U5911 (N_5911,N_3441,N_3193);
nor U5912 (N_5912,N_2886,N_3745);
nor U5913 (N_5913,N_3599,N_3108);
or U5914 (N_5914,N_2304,N_3922);
nor U5915 (N_5915,N_3528,N_2254);
and U5916 (N_5916,N_3594,N_2859);
nor U5917 (N_5917,N_2481,N_2945);
or U5918 (N_5918,N_2390,N_3839);
and U5919 (N_5919,N_3853,N_2478);
and U5920 (N_5920,N_2600,N_3589);
nand U5921 (N_5921,N_3647,N_2361);
or U5922 (N_5922,N_2436,N_2524);
nand U5923 (N_5923,N_3634,N_2624);
or U5924 (N_5924,N_2816,N_3469);
or U5925 (N_5925,N_3833,N_3976);
and U5926 (N_5926,N_3061,N_2415);
and U5927 (N_5927,N_3832,N_2766);
and U5928 (N_5928,N_2202,N_3636);
or U5929 (N_5929,N_2241,N_2521);
and U5930 (N_5930,N_3380,N_2573);
or U5931 (N_5931,N_2786,N_2015);
or U5932 (N_5932,N_2178,N_3065);
or U5933 (N_5933,N_2515,N_3198);
or U5934 (N_5934,N_2918,N_2103);
or U5935 (N_5935,N_3368,N_2611);
or U5936 (N_5936,N_3806,N_2542);
nor U5937 (N_5937,N_2612,N_3417);
nor U5938 (N_5938,N_3094,N_3358);
and U5939 (N_5939,N_2107,N_3204);
or U5940 (N_5940,N_3221,N_2162);
or U5941 (N_5941,N_3925,N_2184);
and U5942 (N_5942,N_2639,N_2211);
nand U5943 (N_5943,N_2872,N_3898);
xor U5944 (N_5944,N_2414,N_2926);
and U5945 (N_5945,N_2253,N_2523);
nand U5946 (N_5946,N_2032,N_3484);
and U5947 (N_5947,N_3594,N_2680);
or U5948 (N_5948,N_3759,N_2624);
or U5949 (N_5949,N_2628,N_2096);
nand U5950 (N_5950,N_2478,N_3680);
nor U5951 (N_5951,N_3441,N_3003);
and U5952 (N_5952,N_3501,N_2086);
nand U5953 (N_5953,N_2050,N_2927);
or U5954 (N_5954,N_3486,N_3967);
nand U5955 (N_5955,N_2440,N_3249);
and U5956 (N_5956,N_2509,N_2089);
and U5957 (N_5957,N_3203,N_3603);
nand U5958 (N_5958,N_2447,N_2620);
nand U5959 (N_5959,N_2277,N_2828);
and U5960 (N_5960,N_2974,N_3833);
nand U5961 (N_5961,N_3795,N_2109);
and U5962 (N_5962,N_3630,N_3798);
nor U5963 (N_5963,N_2641,N_3585);
nor U5964 (N_5964,N_2235,N_3178);
or U5965 (N_5965,N_2761,N_3260);
or U5966 (N_5966,N_3607,N_3990);
or U5967 (N_5967,N_3503,N_2988);
nand U5968 (N_5968,N_3914,N_2992);
and U5969 (N_5969,N_3818,N_3228);
nand U5970 (N_5970,N_3197,N_2308);
nand U5971 (N_5971,N_3696,N_3283);
or U5972 (N_5972,N_2931,N_3306);
nor U5973 (N_5973,N_3796,N_3456);
or U5974 (N_5974,N_3177,N_3921);
and U5975 (N_5975,N_3194,N_2253);
nand U5976 (N_5976,N_3431,N_3427);
nand U5977 (N_5977,N_3355,N_2643);
nand U5978 (N_5978,N_2561,N_2865);
nor U5979 (N_5979,N_3330,N_3230);
and U5980 (N_5980,N_3681,N_2642);
nand U5981 (N_5981,N_2347,N_2633);
or U5982 (N_5982,N_2941,N_3753);
or U5983 (N_5983,N_3086,N_3212);
nand U5984 (N_5984,N_3203,N_3500);
and U5985 (N_5985,N_2668,N_2683);
nand U5986 (N_5986,N_2184,N_3777);
nor U5987 (N_5987,N_3257,N_2284);
nor U5988 (N_5988,N_3822,N_2395);
or U5989 (N_5989,N_3292,N_3889);
nand U5990 (N_5990,N_3436,N_3573);
or U5991 (N_5991,N_3522,N_3950);
or U5992 (N_5992,N_2824,N_3859);
nor U5993 (N_5993,N_3230,N_3944);
nand U5994 (N_5994,N_2520,N_2916);
or U5995 (N_5995,N_2661,N_3731);
or U5996 (N_5996,N_2468,N_3151);
nand U5997 (N_5997,N_2908,N_2535);
or U5998 (N_5998,N_2259,N_2122);
or U5999 (N_5999,N_3416,N_2817);
and U6000 (N_6000,N_4770,N_4283);
nand U6001 (N_6001,N_5899,N_5195);
or U6002 (N_6002,N_5280,N_5695);
and U6003 (N_6003,N_4158,N_5020);
nand U6004 (N_6004,N_5567,N_4986);
and U6005 (N_6005,N_5309,N_5580);
and U6006 (N_6006,N_5140,N_4887);
or U6007 (N_6007,N_5018,N_4467);
nor U6008 (N_6008,N_5273,N_4666);
or U6009 (N_6009,N_4134,N_4150);
nor U6010 (N_6010,N_4246,N_5628);
nor U6011 (N_6011,N_5855,N_4675);
nor U6012 (N_6012,N_5532,N_4284);
or U6013 (N_6013,N_4978,N_4495);
nand U6014 (N_6014,N_5151,N_5376);
or U6015 (N_6015,N_5978,N_5063);
nor U6016 (N_6016,N_5997,N_4093);
nand U6017 (N_6017,N_5191,N_5279);
nand U6018 (N_6018,N_5683,N_5988);
or U6019 (N_6019,N_5318,N_4631);
nor U6020 (N_6020,N_4724,N_5475);
nand U6021 (N_6021,N_4983,N_4453);
and U6022 (N_6022,N_5930,N_5687);
nor U6023 (N_6023,N_5425,N_5431);
nand U6024 (N_6024,N_4826,N_4152);
nor U6025 (N_6025,N_4113,N_5242);
and U6026 (N_6026,N_4255,N_4911);
nor U6027 (N_6027,N_5918,N_4261);
or U6028 (N_6028,N_5188,N_4046);
or U6029 (N_6029,N_4501,N_5562);
and U6030 (N_6030,N_5255,N_4903);
nor U6031 (N_6031,N_4021,N_4984);
and U6032 (N_6032,N_5497,N_4394);
nor U6033 (N_6033,N_4904,N_5525);
or U6034 (N_6034,N_5471,N_5155);
or U6035 (N_6035,N_4757,N_4247);
nand U6036 (N_6036,N_4872,N_4192);
or U6037 (N_6037,N_4435,N_5378);
nand U6038 (N_6038,N_5516,N_4380);
nand U6039 (N_6039,N_4787,N_5552);
nor U6040 (N_6040,N_5791,N_4964);
nor U6041 (N_6041,N_5075,N_4979);
nand U6042 (N_6042,N_5760,N_4156);
and U6043 (N_6043,N_5247,N_4776);
or U6044 (N_6044,N_5897,N_5780);
and U6045 (N_6045,N_4204,N_5396);
nand U6046 (N_6046,N_4734,N_5873);
xnor U6047 (N_6047,N_4325,N_4934);
and U6048 (N_6048,N_4362,N_5402);
nor U6049 (N_6049,N_5608,N_5544);
nor U6050 (N_6050,N_4174,N_4803);
and U6051 (N_6051,N_4746,N_4017);
and U6052 (N_6052,N_4062,N_5088);
or U6053 (N_6053,N_4109,N_4430);
nand U6054 (N_6054,N_5771,N_5297);
or U6055 (N_6055,N_4310,N_5754);
nand U6056 (N_6056,N_5688,N_4193);
nor U6057 (N_6057,N_5194,N_4267);
or U6058 (N_6058,N_5511,N_5970);
or U6059 (N_6059,N_4483,N_4208);
or U6060 (N_6060,N_4140,N_4167);
nand U6061 (N_6061,N_5727,N_4254);
and U6062 (N_6062,N_5914,N_5428);
or U6063 (N_6063,N_5951,N_5576);
nand U6064 (N_6064,N_4699,N_5631);
or U6065 (N_6065,N_5937,N_5369);
xor U6066 (N_6066,N_5885,N_5905);
or U6067 (N_6067,N_4458,N_5207);
and U6068 (N_6068,N_5572,N_4792);
nand U6069 (N_6069,N_4009,N_4440);
and U6070 (N_6070,N_5617,N_5526);
nand U6071 (N_6071,N_5622,N_4235);
nand U6072 (N_6072,N_4682,N_4993);
nor U6073 (N_6073,N_5149,N_5130);
nand U6074 (N_6074,N_4599,N_5296);
or U6075 (N_6075,N_5841,N_4895);
nand U6076 (N_6076,N_5346,N_4484);
and U6077 (N_6077,N_5190,N_4580);
or U6078 (N_6078,N_4443,N_4120);
and U6079 (N_6079,N_5728,N_4956);
nor U6080 (N_6080,N_4859,N_4361);
or U6081 (N_6081,N_4111,N_5809);
or U6082 (N_6082,N_5457,N_4894);
or U6083 (N_6083,N_4653,N_5927);
and U6084 (N_6084,N_5398,N_5110);
and U6085 (N_6085,N_4236,N_4590);
nor U6086 (N_6086,N_4054,N_5848);
nand U6087 (N_6087,N_4099,N_5454);
or U6088 (N_6088,N_4268,N_4578);
or U6089 (N_6089,N_4239,N_4588);
nor U6090 (N_6090,N_5568,N_5571);
or U6091 (N_6091,N_4926,N_4582);
nand U6092 (N_6092,N_5230,N_5726);
and U6093 (N_6093,N_5104,N_5347);
or U6094 (N_6094,N_5667,N_5514);
or U6095 (N_6095,N_4795,N_5894);
nand U6096 (N_6096,N_5226,N_5636);
nand U6097 (N_6097,N_5417,N_4948);
or U6098 (N_6098,N_5050,N_4216);
or U6099 (N_6099,N_5886,N_5872);
nand U6100 (N_6100,N_5253,N_5258);
or U6101 (N_6101,N_4034,N_4605);
and U6102 (N_6102,N_5249,N_5310);
nor U6103 (N_6103,N_4581,N_5038);
nand U6104 (N_6104,N_5819,N_5351);
or U6105 (N_6105,N_4013,N_4711);
and U6106 (N_6106,N_5118,N_5916);
and U6107 (N_6107,N_4579,N_4504);
or U6108 (N_6108,N_4468,N_4656);
and U6109 (N_6109,N_5477,N_4667);
nor U6110 (N_6110,N_5401,N_5634);
nand U6111 (N_6111,N_5559,N_4908);
nor U6112 (N_6112,N_5181,N_4975);
or U6113 (N_6113,N_5212,N_4873);
nand U6114 (N_6114,N_4808,N_5787);
or U6115 (N_6115,N_4147,N_4418);
or U6116 (N_6116,N_5842,N_5912);
or U6117 (N_6117,N_4555,N_5330);
nand U6118 (N_6118,N_5120,N_5095);
nor U6119 (N_6119,N_4506,N_4011);
nor U6120 (N_6120,N_4498,N_4250);
nand U6121 (N_6121,N_5519,N_4187);
nand U6122 (N_6122,N_5926,N_5876);
and U6123 (N_6123,N_5372,N_5414);
nand U6124 (N_6124,N_5302,N_4971);
and U6125 (N_6125,N_5343,N_4633);
nor U6126 (N_6126,N_5764,N_4355);
xor U6127 (N_6127,N_5633,N_4058);
or U6128 (N_6128,N_5100,N_5768);
nand U6129 (N_6129,N_5956,N_4122);
and U6130 (N_6130,N_4020,N_5850);
and U6131 (N_6131,N_4816,N_5933);
and U6132 (N_6132,N_4996,N_5678);
or U6133 (N_6133,N_5495,N_4118);
nor U6134 (N_6134,N_5411,N_5476);
and U6135 (N_6135,N_5698,N_5071);
nand U6136 (N_6136,N_5136,N_4755);
or U6137 (N_6137,N_4095,N_5959);
or U6138 (N_6138,N_5998,N_5064);
nor U6139 (N_6139,N_4264,N_4562);
nor U6140 (N_6140,N_5700,N_4415);
nand U6141 (N_6141,N_5621,N_4696);
nor U6142 (N_6142,N_5877,N_4447);
nor U6143 (N_6143,N_5804,N_5452);
or U6144 (N_6144,N_4516,N_5157);
and U6145 (N_6145,N_5736,N_5939);
nor U6146 (N_6146,N_5045,N_4995);
or U6147 (N_6147,N_4469,N_4330);
and U6148 (N_6148,N_5512,N_5578);
and U6149 (N_6149,N_4368,N_5394);
nor U6150 (N_6150,N_4847,N_5437);
nor U6151 (N_6151,N_5616,N_5725);
or U6152 (N_6152,N_5052,N_4210);
and U6153 (N_6153,N_4314,N_4742);
nor U6154 (N_6154,N_4545,N_5220);
nand U6155 (N_6155,N_5598,N_5328);
nor U6156 (N_6156,N_5976,N_4870);
nand U6157 (N_6157,N_4388,N_5917);
and U6158 (N_6158,N_4999,N_5947);
and U6159 (N_6159,N_5153,N_4139);
nand U6160 (N_6160,N_4214,N_5421);
and U6161 (N_6161,N_4212,N_4358);
nor U6162 (N_6162,N_5966,N_4220);
and U6163 (N_6163,N_5805,N_5761);
and U6164 (N_6164,N_5252,N_5134);
nor U6165 (N_6165,N_4805,N_5314);
or U6166 (N_6166,N_5419,N_5447);
or U6167 (N_6167,N_4091,N_5023);
and U6168 (N_6168,N_4016,N_4019);
and U6169 (N_6169,N_4177,N_4442);
nand U6170 (N_6170,N_5931,N_4491);
and U6171 (N_6171,N_5440,N_4456);
or U6172 (N_6172,N_4830,N_5671);
nand U6173 (N_6173,N_4481,N_5438);
nor U6174 (N_6174,N_4237,N_5270);
or U6175 (N_6175,N_5464,N_4660);
nand U6176 (N_6176,N_5215,N_4608);
nor U6177 (N_6177,N_5745,N_4138);
nand U6178 (N_6178,N_5932,N_5061);
nand U6179 (N_6179,N_5126,N_5742);
nor U6180 (N_6180,N_5500,N_5265);
nor U6181 (N_6181,N_5166,N_4315);
nand U6182 (N_6182,N_4727,N_4640);
nor U6183 (N_6183,N_5028,N_4129);
nand U6184 (N_6184,N_5847,N_5219);
or U6185 (N_6185,N_5349,N_4086);
nand U6186 (N_6186,N_4142,N_5364);
nor U6187 (N_6187,N_4252,N_4197);
and U6188 (N_6188,N_4061,N_4240);
nor U6189 (N_6189,N_4128,N_4572);
or U6190 (N_6190,N_4914,N_5418);
nor U6191 (N_6191,N_5016,N_4026);
nand U6192 (N_6192,N_5625,N_5743);
and U6193 (N_6193,N_5766,N_5363);
nor U6194 (N_6194,N_5081,N_4836);
nor U6195 (N_6195,N_4701,N_4381);
nand U6196 (N_6196,N_4922,N_5164);
or U6197 (N_6197,N_4326,N_4840);
nand U6198 (N_6198,N_4248,N_4419);
nor U6199 (N_6199,N_4014,N_4117);
or U6200 (N_6200,N_5000,N_4733);
or U6201 (N_6201,N_4613,N_4991);
nor U6202 (N_6202,N_4302,N_4589);
nor U6203 (N_6203,N_5325,N_5554);
or U6204 (N_6204,N_5759,N_4012);
nand U6205 (N_6205,N_5903,N_5090);
and U6206 (N_6206,N_4346,N_5292);
or U6207 (N_6207,N_4750,N_5094);
or U6208 (N_6208,N_4918,N_5575);
and U6209 (N_6209,N_4151,N_4815);
nand U6210 (N_6210,N_5246,N_5596);
xor U6211 (N_6211,N_5360,N_5233);
or U6212 (N_6212,N_4657,N_5680);
and U6213 (N_6213,N_4707,N_4593);
or U6214 (N_6214,N_5439,N_5991);
and U6215 (N_6215,N_4921,N_5611);
and U6216 (N_6216,N_4766,N_4690);
nor U6217 (N_6217,N_5920,N_4577);
nand U6218 (N_6218,N_4981,N_5757);
nor U6219 (N_6219,N_5952,N_5150);
and U6220 (N_6220,N_5869,N_4260);
and U6221 (N_6221,N_4771,N_4751);
nor U6222 (N_6222,N_5125,N_5925);
nand U6223 (N_6223,N_5820,N_4265);
or U6224 (N_6224,N_4327,N_4624);
nor U6225 (N_6225,N_4459,N_4172);
nand U6226 (N_6226,N_5986,N_5665);
nand U6227 (N_6227,N_4632,N_4655);
nand U6228 (N_6228,N_5606,N_5227);
and U6229 (N_6229,N_4731,N_5675);
or U6230 (N_6230,N_5710,N_4723);
or U6231 (N_6231,N_4171,N_5335);
nand U6232 (N_6232,N_4654,N_4909);
and U6233 (N_6233,N_4100,N_4060);
nand U6234 (N_6234,N_4162,N_4671);
or U6235 (N_6235,N_4321,N_4332);
and U6236 (N_6236,N_5109,N_4568);
nand U6237 (N_6237,N_5307,N_5790);
nand U6238 (N_6238,N_4329,N_4460);
nand U6239 (N_6239,N_4040,N_5702);
or U6240 (N_6240,N_5413,N_5668);
or U6241 (N_6241,N_4865,N_4931);
nand U6242 (N_6242,N_5837,N_4420);
and U6243 (N_6243,N_4899,N_5659);
xnor U6244 (N_6244,N_4797,N_5973);
or U6245 (N_6245,N_5672,N_4584);
nor U6246 (N_6246,N_4886,N_4672);
nor U6247 (N_6247,N_5740,N_5216);
nand U6248 (N_6248,N_4681,N_5218);
nor U6249 (N_6249,N_4846,N_4520);
or U6250 (N_6250,N_4548,N_5213);
nand U6251 (N_6251,N_5906,N_4299);
nand U6252 (N_6252,N_5225,N_4901);
xor U6253 (N_6253,N_5479,N_5012);
and U6254 (N_6254,N_5393,N_4271);
or U6255 (N_6255,N_5783,N_5317);
nor U6256 (N_6256,N_4774,N_4612);
nand U6257 (N_6257,N_4647,N_4807);
and U6258 (N_6258,N_4243,N_4068);
and U6259 (N_6259,N_5652,N_5160);
nand U6260 (N_6260,N_4627,N_4287);
or U6261 (N_6261,N_4730,N_5716);
nand U6262 (N_6262,N_4546,N_5241);
or U6263 (N_6263,N_5266,N_4376);
nand U6264 (N_6264,N_5893,N_4607);
and U6265 (N_6265,N_4526,N_4630);
nor U6266 (N_6266,N_5019,N_4360);
and U6267 (N_6267,N_5400,N_5067);
nor U6268 (N_6268,N_5184,N_5733);
nor U6269 (N_6269,N_5456,N_5527);
xnor U6270 (N_6270,N_5092,N_4449);
and U6271 (N_6271,N_5531,N_5251);
or U6272 (N_6272,N_4281,N_5640);
nand U6273 (N_6273,N_4799,N_4888);
and U6274 (N_6274,N_4359,N_5504);
nor U6275 (N_6275,N_4992,N_4475);
nand U6276 (N_6276,N_5984,N_4769);
or U6277 (N_6277,N_4850,N_5713);
nor U6278 (N_6278,N_4432,N_4749);
or U6279 (N_6279,N_5581,N_5046);
nor U6280 (N_6280,N_5538,N_4066);
nand U6281 (N_6281,N_5679,N_5461);
nand U6282 (N_6282,N_4333,N_4476);
and U6283 (N_6283,N_5674,N_4153);
nand U6284 (N_6284,N_5615,N_5523);
nand U6285 (N_6285,N_5256,N_5008);
nor U6286 (N_6286,N_5548,N_4125);
and U6287 (N_6287,N_4241,N_4941);
and U6288 (N_6288,N_5545,N_4636);
or U6289 (N_6289,N_4038,N_4409);
or U6290 (N_6290,N_5792,N_4688);
nand U6291 (N_6291,N_5948,N_4154);
or U6292 (N_6292,N_4573,N_4067);
and U6293 (N_6293,N_4871,N_5676);
nand U6294 (N_6294,N_4963,N_4356);
nand U6295 (N_6295,N_5815,N_4768);
or U6296 (N_6296,N_4375,N_4396);
or U6297 (N_6297,N_4298,N_4905);
and U6298 (N_6298,N_5185,N_4085);
nor U6299 (N_6299,N_5222,N_5732);
or U6300 (N_6300,N_4441,N_4869);
nand U6301 (N_6301,N_5717,N_4189);
nand U6302 (N_6302,N_5515,N_5856);
nor U6303 (N_6303,N_5958,N_4628);
nand U6304 (N_6304,N_4595,N_4124);
and U6305 (N_6305,N_4141,N_5076);
and U6306 (N_6306,N_5410,N_5341);
and U6307 (N_6307,N_5705,N_5096);
nand U6308 (N_6308,N_5186,N_4338);
and U6309 (N_6309,N_4175,N_4301);
nor U6310 (N_6310,N_4446,N_4598);
nand U6311 (N_6311,N_4383,N_4290);
nor U6312 (N_6312,N_4743,N_4411);
or U6313 (N_6313,N_4207,N_4018);
or U6314 (N_6314,N_4079,N_4758);
nor U6315 (N_6315,N_4790,N_5170);
nand U6316 (N_6316,N_5312,N_5189);
or U6317 (N_6317,N_4047,N_5326);
nand U6318 (N_6318,N_4575,N_4933);
nor U6319 (N_6319,N_5604,N_4928);
or U6320 (N_6320,N_5404,N_5874);
or U6321 (N_6321,N_4074,N_4163);
or U6322 (N_6322,N_4245,N_5355);
nand U6323 (N_6323,N_4354,N_5391);
nor U6324 (N_6324,N_5789,N_5786);
and U6325 (N_6325,N_5942,N_5582);
nand U6326 (N_6326,N_4276,N_4937);
nand U6327 (N_6327,N_4434,N_5223);
and U6328 (N_6328,N_5434,N_5272);
and U6329 (N_6329,N_5642,N_4282);
and U6330 (N_6330,N_4146,N_4882);
nand U6331 (N_6331,N_4684,N_4752);
nand U6332 (N_6332,N_5569,N_4164);
or U6333 (N_6333,N_5620,N_4635);
nor U6334 (N_6334,N_5321,N_4834);
and U6335 (N_6335,N_5175,N_4035);
and U6336 (N_6336,N_4412,N_5699);
and U6337 (N_6337,N_5719,N_5880);
nor U6338 (N_6338,N_5972,N_5248);
or U6339 (N_6339,N_5954,N_5735);
nor U6340 (N_6340,N_4883,N_4527);
and U6341 (N_6341,N_4088,N_4715);
nor U6342 (N_6342,N_5980,N_4536);
nor U6343 (N_6343,N_5446,N_5042);
nor U6344 (N_6344,N_4958,N_5843);
and U6345 (N_6345,N_4788,N_4528);
and U6346 (N_6346,N_5051,N_5770);
or U6347 (N_6347,N_5911,N_5802);
or U6348 (N_6348,N_5276,N_5331);
nand U6349 (N_6349,N_5995,N_4233);
nor U6350 (N_6350,N_4370,N_4912);
nand U6351 (N_6351,N_4002,N_5448);
nor U6352 (N_6352,N_5694,N_5558);
or U6353 (N_6353,N_5826,N_4663);
or U6354 (N_6354,N_5977,N_5513);
and U6355 (N_6355,N_4005,N_5922);
or U6356 (N_6356,N_5782,N_4102);
nor U6357 (N_6357,N_5483,N_4274);
and U6358 (N_6358,N_5825,N_4879);
or U6359 (N_6359,N_5221,N_5442);
nand U6360 (N_6360,N_4994,N_4829);
and U6361 (N_6361,N_5180,N_5301);
nand U6362 (N_6362,N_4006,N_4132);
and U6363 (N_6363,N_4404,N_5397);
and U6364 (N_6364,N_5217,N_5585);
nor U6365 (N_6365,N_4509,N_5384);
or U6366 (N_6366,N_5586,N_5648);
nor U6367 (N_6367,N_5143,N_4126);
and U6368 (N_6368,N_5589,N_5473);
nand U6369 (N_6369,N_4385,N_5472);
or U6370 (N_6370,N_5111,N_5953);
nor U6371 (N_6371,N_5741,N_4200);
nor U6372 (N_6372,N_5773,N_4490);
nor U6373 (N_6373,N_5103,N_4223);
nand U6374 (N_6374,N_5853,N_4423);
nor U6375 (N_6375,N_4482,N_4070);
nand U6376 (N_6376,N_5549,N_5451);
and U6377 (N_6377,N_4523,N_5852);
or U6378 (N_6378,N_5281,N_5141);
nand U6379 (N_6379,N_4625,N_5798);
or U6380 (N_6380,N_5300,N_4782);
or U6381 (N_6381,N_4661,N_4463);
nand U6382 (N_6382,N_4538,N_4676);
or U6383 (N_6383,N_4535,N_4553);
and U6384 (N_6384,N_4053,N_5083);
or U6385 (N_6385,N_5767,N_4096);
nor U6386 (N_6386,N_4347,N_5867);
nor U6387 (N_6387,N_5047,N_5860);
nor U6388 (N_6388,N_5555,N_4195);
and U6389 (N_6389,N_5535,N_4897);
and U6390 (N_6390,N_4611,N_5487);
nor U6391 (N_6391,N_5835,N_5910);
xor U6392 (N_6392,N_5929,N_5583);
and U6393 (N_6393,N_5144,N_4566);
nand U6394 (N_6394,N_4953,N_4479);
and U6395 (N_6395,N_5298,N_4709);
nor U6396 (N_6396,N_4306,N_5799);
nand U6397 (N_6397,N_4263,N_5074);
nand U6398 (N_6398,N_4041,N_5229);
nor U6399 (N_6399,N_5563,N_4097);
and U6400 (N_6400,N_5499,N_5817);
nand U6401 (N_6401,N_5750,N_5553);
or U6402 (N_6402,N_4379,N_5938);
nor U6403 (N_6403,N_5490,N_4779);
nand U6404 (N_6404,N_4324,N_4781);
or U6405 (N_6405,N_5123,N_5520);
nor U6406 (N_6406,N_5573,N_4540);
and U6407 (N_6407,N_4397,N_4165);
nor U6408 (N_6408,N_4135,N_4344);
and U6409 (N_6409,N_4051,N_4874);
or U6410 (N_6410,N_4119,N_4371);
and U6411 (N_6411,N_4515,N_4042);
or U6412 (N_6412,N_4462,N_5077);
and U6413 (N_6413,N_4194,N_4902);
nor U6414 (N_6414,N_5202,N_4244);
nand U6415 (N_6415,N_5305,N_5138);
or U6416 (N_6416,N_4960,N_5488);
nand U6417 (N_6417,N_4444,N_4427);
nor U6418 (N_6418,N_4110,N_4763);
and U6419 (N_6419,N_4669,N_4105);
nand U6420 (N_6420,N_5154,N_5163);
or U6421 (N_6421,N_5032,N_4438);
and U6422 (N_6422,N_4203,N_4848);
and U6423 (N_6423,N_4309,N_4739);
or U6424 (N_6424,N_4266,N_5579);
nor U6425 (N_6425,N_4817,N_4689);
nor U6426 (N_6426,N_4155,N_4622);
and U6427 (N_6427,N_5696,N_4576);
nor U6428 (N_6428,N_5387,N_5287);
and U6429 (N_6429,N_4319,N_5999);
nor U6430 (N_6430,N_5338,N_5127);
nand U6431 (N_6431,N_5883,N_4534);
nand U6432 (N_6432,N_4521,N_4962);
nand U6433 (N_6433,N_4496,N_4778);
or U6434 (N_6434,N_4511,N_4721);
and U6435 (N_6435,N_5884,N_5540);
and U6436 (N_6436,N_4278,N_5533);
or U6437 (N_6437,N_5199,N_4679);
or U6438 (N_6438,N_5308,N_4819);
nor U6439 (N_6439,N_5721,N_4036);
nand U6440 (N_6440,N_5715,N_4081);
nand U6441 (N_6441,N_5793,N_5379);
and U6442 (N_6442,N_4982,N_5602);
nand U6443 (N_6443,N_5878,N_5196);
and U6444 (N_6444,N_4304,N_4961);
xnor U6445 (N_6445,N_5594,N_5781);
nand U6446 (N_6446,N_5755,N_5896);
or U6447 (N_6447,N_5902,N_4231);
or U6448 (N_6448,N_4802,N_4917);
or U6449 (N_6449,N_4296,N_5964);
or U6450 (N_6450,N_5101,N_4116);
or U6451 (N_6451,N_4272,N_4533);
nand U6452 (N_6452,N_4114,N_5803);
or U6453 (N_6453,N_4080,N_4289);
nand U6454 (N_6454,N_5591,N_4004);
nor U6455 (N_6455,N_4084,N_5203);
nand U6456 (N_6456,N_4069,N_4487);
nand U6457 (N_6457,N_4227,N_5015);
nand U6458 (N_6458,N_5291,N_5179);
and U6459 (N_6459,N_5963,N_5868);
or U6460 (N_6460,N_4760,N_4753);
and U6461 (N_6461,N_4747,N_5635);
and U6462 (N_6462,N_4785,N_5430);
nand U6463 (N_6463,N_5277,N_5691);
or U6464 (N_6464,N_5231,N_4205);
nor U6465 (N_6465,N_4664,N_5610);
or U6466 (N_6466,N_5650,N_4144);
nand U6467 (N_6467,N_4213,N_4955);
or U6468 (N_6468,N_4809,N_4190);
and U6469 (N_6469,N_5587,N_4065);
and U6470 (N_6470,N_5935,N_4686);
nor U6471 (N_6471,N_4417,N_5168);
nand U6472 (N_6472,N_4644,N_5812);
nand U6473 (N_6473,N_5982,N_5530);
xor U6474 (N_6474,N_5171,N_5971);
and U6475 (N_6475,N_4571,N_5666);
or U6476 (N_6476,N_5827,N_4104);
nor U6477 (N_6477,N_5744,N_5936);
or U6478 (N_6478,N_4225,N_5517);
nand U6479 (N_6479,N_5777,N_5941);
or U6480 (N_6480,N_5366,N_5565);
nor U6481 (N_6481,N_4569,N_5035);
and U6482 (N_6482,N_4551,N_4023);
nor U6483 (N_6483,N_5630,N_5601);
or U6484 (N_6484,N_4854,N_5048);
nor U6485 (N_6485,N_5261,N_5967);
nor U6486 (N_6486,N_4073,N_5173);
nand U6487 (N_6487,N_4188,N_5915);
or U6488 (N_6488,N_4884,N_4930);
nor U6489 (N_6489,N_5373,N_4431);
or U6490 (N_6490,N_4784,N_4615);
and U6491 (N_6491,N_4662,N_5085);
and U6492 (N_6492,N_5521,N_4519);
and U6493 (N_6493,N_4437,N_5463);
nor U6494 (N_6494,N_4032,N_5114);
and U6495 (N_6495,N_5010,N_5528);
nor U6496 (N_6496,N_5731,N_5752);
or U6497 (N_6497,N_5228,N_5994);
nor U6498 (N_6498,N_5089,N_4288);
nand U6499 (N_6499,N_5329,N_5235);
or U6500 (N_6500,N_4651,N_4775);
nand U6501 (N_6501,N_4702,N_5776);
nand U6502 (N_6502,N_5557,N_4334);
and U6503 (N_6503,N_4998,N_5316);
and U6504 (N_6504,N_5858,N_4173);
or U6505 (N_6505,N_4885,N_5361);
and U6506 (N_6506,N_4010,N_4855);
xor U6507 (N_6507,N_4997,N_4765);
nor U6508 (N_6508,N_5639,N_5283);
nand U6509 (N_6509,N_5550,N_5785);
or U6510 (N_6510,N_4604,N_5161);
nor U6511 (N_6511,N_5086,N_4974);
or U6512 (N_6512,N_4337,N_4814);
and U6513 (N_6513,N_4988,N_4098);
nand U6514 (N_6514,N_5993,N_4471);
nand U6515 (N_6515,N_5961,N_4838);
or U6516 (N_6516,N_5737,N_4373);
nand U6517 (N_6517,N_5974,N_5453);
and U6518 (N_6518,N_4094,N_5775);
nor U6519 (N_6519,N_5200,N_5822);
nand U6520 (N_6520,N_4698,N_5823);
and U6521 (N_6521,N_4985,N_5593);
and U6522 (N_6522,N_5165,N_4136);
nor U6523 (N_6523,N_4502,N_4563);
and U6524 (N_6524,N_5263,N_5618);
or U6525 (N_6525,N_4168,N_4421);
and U6526 (N_6526,N_5493,N_5178);
and U6527 (N_6527,N_5443,N_5380);
nand U6528 (N_6528,N_5844,N_4352);
nor U6529 (N_6529,N_5002,N_5132);
nor U6530 (N_6530,N_5353,N_4665);
or U6531 (N_6531,N_5004,N_4294);
nand U6532 (N_6532,N_4101,N_5319);
and U6533 (N_6533,N_5259,N_4391);
nand U6534 (N_6534,N_5091,N_4877);
nand U6535 (N_6535,N_5409,N_4554);
or U6536 (N_6536,N_5108,N_4387);
or U6537 (N_6537,N_4637,N_4783);
or U6538 (N_6538,N_5670,N_4425);
nor U6539 (N_6539,N_5183,N_5892);
nor U6540 (N_6540,N_5232,N_5870);
nand U6541 (N_6541,N_4735,N_5407);
and U6542 (N_6542,N_5801,N_4257);
nand U6543 (N_6543,N_4049,N_5113);
and U6544 (N_6544,N_5315,N_5854);
or U6545 (N_6545,N_4947,N_5128);
xnor U6546 (N_6546,N_4532,N_5365);
and U6547 (N_6547,N_4537,N_5159);
nand U6548 (N_6548,N_4022,N_4372);
or U6549 (N_6549,N_5949,N_5663);
and U6550 (N_6550,N_4279,N_5208);
xor U6551 (N_6551,N_5262,N_4839);
nand U6552 (N_6552,N_4720,N_5098);
and U6553 (N_6553,N_4033,N_5882);
nand U6554 (N_6554,N_4889,N_4827);
nand U6555 (N_6555,N_5368,N_5121);
nor U6556 (N_6556,N_4439,N_5501);
nor U6557 (N_6557,N_5362,N_5058);
nand U6558 (N_6558,N_5901,N_4377);
and U6559 (N_6559,N_4710,N_5043);
and U6560 (N_6560,N_4952,N_5480);
and U6561 (N_6561,N_4629,N_4003);
and U6562 (N_6562,N_5005,N_4044);
nor U6563 (N_6563,N_4180,N_5267);
and U6564 (N_6564,N_4764,N_5838);
nor U6565 (N_6565,N_4063,N_5177);
or U6566 (N_6566,N_5260,N_5322);
nand U6567 (N_6567,N_5286,N_4323);
or U6568 (N_6568,N_5763,N_5257);
and U6569 (N_6569,N_5669,N_5758);
nand U6570 (N_6570,N_4112,N_4619);
nor U6571 (N_6571,N_4585,N_4972);
nand U6572 (N_6572,N_5320,N_5470);
or U6573 (N_6573,N_4382,N_4924);
and U6574 (N_6574,N_5810,N_4031);
nand U6575 (N_6575,N_4363,N_4620);
and U6576 (N_6576,N_4977,N_4277);
or U6577 (N_6577,N_4378,N_5818);
nand U6578 (N_6578,N_5624,N_5137);
and U6579 (N_6579,N_4754,N_4374);
nand U6580 (N_6580,N_4028,N_5234);
and U6581 (N_6581,N_5655,N_5460);
nand U6582 (N_6582,N_4413,N_4348);
nand U6583 (N_6583,N_5778,N_4740);
nor U6584 (N_6584,N_4148,N_4410);
nor U6585 (N_6585,N_5701,N_5429);
nand U6586 (N_6586,N_5522,N_5268);
or U6587 (N_6587,N_5416,N_4072);
or U6588 (N_6588,N_4428,N_4196);
nor U6589 (N_6589,N_4357,N_4253);
or U6590 (N_6590,N_5436,N_5390);
nor U6591 (N_6591,N_4966,N_4039);
and U6592 (N_6592,N_5529,N_5112);
nand U6593 (N_6593,N_5303,N_4641);
and U6594 (N_6594,N_5489,N_4759);
and U6595 (N_6595,N_4617,N_4229);
and U6596 (N_6596,N_5357,N_4891);
or U6597 (N_6597,N_5037,N_5382);
and U6598 (N_6598,N_5657,N_5808);
nor U6599 (N_6599,N_5498,N_5254);
nand U6600 (N_6600,N_4127,N_4861);
and U6601 (N_6601,N_4161,N_4336);
or U6602 (N_6602,N_4959,N_4967);
nor U6603 (N_6603,N_5311,N_5774);
and U6604 (N_6604,N_4531,N_4202);
nor U6605 (N_6605,N_5983,N_5654);
and U6606 (N_6606,N_4567,N_5306);
nor U6607 (N_6607,N_4512,N_4646);
and U6608 (N_6608,N_4693,N_4182);
or U6609 (N_6609,N_5041,N_4293);
nand U6610 (N_6610,N_5632,N_5607);
nand U6611 (N_6611,N_4932,N_5236);
or U6612 (N_6612,N_5969,N_5026);
and U6613 (N_6613,N_5542,N_5433);
nor U6614 (N_6614,N_4549,N_5465);
or U6615 (N_6615,N_5455,N_5795);
nand U6616 (N_6616,N_5211,N_5765);
or U6617 (N_6617,N_4694,N_5800);
and U6618 (N_6618,N_4920,N_4878);
and U6619 (N_6619,N_5560,N_4547);
or U6620 (N_6620,N_4591,N_4414);
nand U6621 (N_6621,N_4791,N_4454);
and U6622 (N_6622,N_5638,N_5068);
or U6623 (N_6623,N_4907,N_4601);
nand U6624 (N_6624,N_5851,N_5697);
nand U6625 (N_6625,N_5375,N_4320);
or U6626 (N_6626,N_4464,N_5206);
nand U6627 (N_6627,N_5950,N_5919);
nand U6628 (N_6628,N_4249,N_4824);
nand U6629 (N_6629,N_4728,N_4489);
nor U6630 (N_6630,N_5739,N_4478);
nand U6631 (N_6631,N_5597,N_4713);
nand U6632 (N_6632,N_4700,N_5299);
or U6633 (N_6633,N_5269,N_4793);
and U6634 (N_6634,N_4322,N_4866);
nand U6635 (N_6635,N_5588,N_5336);
nor U6636 (N_6636,N_4416,N_4570);
nand U6637 (N_6637,N_4825,N_4513);
and U6638 (N_6638,N_5720,N_5313);
and U6639 (N_6639,N_4400,N_5145);
nor U6640 (N_6640,N_4936,N_4228);
nor U6641 (N_6641,N_5749,N_5274);
nor U6642 (N_6642,N_5135,N_4123);
or U6643 (N_6643,N_4366,N_5685);
or U6644 (N_6644,N_5459,N_5332);
nor U6645 (N_6645,N_5139,N_4881);
nand U6646 (N_6646,N_5681,N_5371);
and U6647 (N_6647,N_4317,N_5900);
or U6648 (N_6648,N_5730,N_5981);
nor U6649 (N_6649,N_5466,N_5115);
nand U6650 (N_6650,N_4470,N_5857);
nor U6651 (N_6651,N_4064,N_4349);
and U6652 (N_6652,N_5105,N_4384);
nand U6653 (N_6653,N_4818,N_4219);
and U6654 (N_6654,N_4452,N_5506);
nand U6655 (N_6655,N_4048,N_5192);
nand U6656 (N_6656,N_5482,N_4645);
and U6657 (N_6657,N_5009,N_5612);
or U6658 (N_6658,N_4313,N_5992);
or U6659 (N_6659,N_4224,N_4852);
nand U6660 (N_6660,N_4522,N_5832);
nor U6661 (N_6661,N_4541,N_5239);
or U6662 (N_6662,N_5057,N_5444);
nor U6663 (N_6663,N_5044,N_5592);
and U6664 (N_6664,N_5703,N_5603);
or U6665 (N_6665,N_4341,N_5968);
nand U6666 (N_6666,N_5340,N_5107);
xnor U6667 (N_6667,N_4798,N_4609);
nor U6668 (N_6668,N_4856,N_5469);
nand U6669 (N_6669,N_4445,N_4029);
nor U6670 (N_6670,N_4108,N_5551);
nand U6671 (N_6671,N_4718,N_4007);
and U6672 (N_6672,N_5133,N_4639);
and U6673 (N_6673,N_5831,N_5828);
and U6674 (N_6674,N_4311,N_5069);
nand U6675 (N_6675,N_5129,N_5637);
nor U6676 (N_6676,N_4226,N_4390);
or U6677 (N_6677,N_4910,N_5861);
nor U6678 (N_6678,N_4485,N_4078);
and U6679 (N_6679,N_4056,N_5859);
or U6680 (N_6680,N_4198,N_5946);
or U6681 (N_6681,N_5162,N_4251);
nand U6682 (N_6682,N_5690,N_5093);
or U6683 (N_6683,N_4083,N_4230);
xnor U6684 (N_6684,N_4403,N_4831);
nand U6685 (N_6685,N_4945,N_4340);
nand U6686 (N_6686,N_4238,N_4001);
and U6687 (N_6687,N_5541,N_5955);
nand U6688 (N_6688,N_4143,N_5875);
or U6689 (N_6689,N_4087,N_4801);
nor U6690 (N_6690,N_4990,N_4280);
or U6691 (N_6691,N_4291,N_4369);
nand U6692 (N_6692,N_5746,N_4550);
and U6693 (N_6693,N_5275,N_5122);
and U6694 (N_6694,N_5034,N_4652);
or U6695 (N_6695,N_4557,N_4965);
nand U6696 (N_6696,N_4183,N_4386);
nand U6697 (N_6697,N_5422,N_5412);
nand U6698 (N_6698,N_4744,N_5282);
or U6699 (N_6699,N_4761,N_5237);
and U6700 (N_6700,N_4695,N_4705);
nand U6701 (N_6701,N_4273,N_5662);
or U6702 (N_6702,N_4714,N_5467);
nor U6703 (N_6703,N_4149,N_5358);
nor U6704 (N_6704,N_4166,N_4692);
or U6705 (N_6705,N_4685,N_5940);
nand U6706 (N_6706,N_4729,N_4181);
nand U6707 (N_6707,N_4969,N_5492);
nor U6708 (N_6708,N_4913,N_4050);
nor U6709 (N_6709,N_4179,N_5813);
and U6710 (N_6710,N_4927,N_5865);
nand U6711 (N_6711,N_4473,N_4683);
and U6712 (N_6712,N_4726,N_5027);
nor U6713 (N_6713,N_5288,N_5965);
or U6714 (N_6714,N_4583,N_5866);
nor U6715 (N_6715,N_5904,N_4436);
nand U6716 (N_6716,N_5824,N_5907);
and U6717 (N_6717,N_5619,N_5066);
or U6718 (N_6718,N_5478,N_5863);
or U6719 (N_6719,N_4524,N_4822);
or U6720 (N_6720,N_5600,N_5462);
or U6721 (N_6721,N_4773,N_5943);
nand U6722 (N_6722,N_5889,N_4160);
nor U6723 (N_6723,N_4395,N_5119);
nand U6724 (N_6724,N_4564,N_4343);
and U6725 (N_6725,N_4137,N_4565);
nor U6726 (N_6726,N_5458,N_4145);
or U6727 (N_6727,N_4868,N_5395);
nor U6728 (N_6728,N_4082,N_4804);
and U6729 (N_6729,N_4530,N_5729);
nand U6730 (N_6730,N_4594,N_4133);
nor U6731 (N_6731,N_5647,N_4864);
and U6732 (N_6732,N_4558,N_4275);
nor U6733 (N_6733,N_4242,N_5794);
nand U6734 (N_6734,N_4121,N_5605);
nand U6735 (N_6735,N_5449,N_5036);
and U6736 (N_6736,N_5686,N_4106);
nand U6737 (N_6737,N_5345,N_4398);
nand U6738 (N_6738,N_4935,N_5485);
and U6739 (N_6739,N_4845,N_4429);
nor U6740 (N_6740,N_4486,N_5864);
nor U6741 (N_6741,N_4130,N_4389);
nor U6742 (N_6742,N_4949,N_5209);
nand U6743 (N_6743,N_5833,N_5474);
and U6744 (N_6744,N_4217,N_5484);
nor U6745 (N_6745,N_4716,N_4706);
nor U6746 (N_6746,N_5435,N_4426);
and U6747 (N_6747,N_4722,N_5003);
nand U6748 (N_6748,N_5546,N_5022);
and U6749 (N_6749,N_5881,N_5073);
nand U6750 (N_6750,N_4399,N_4493);
and U6751 (N_6751,N_5339,N_4860);
nor U6752 (N_6752,N_4015,N_5158);
nand U6753 (N_6753,N_4488,N_4043);
nand U6754 (N_6754,N_5264,N_4024);
or U6755 (N_6755,N_4833,N_5830);
or U6756 (N_6756,N_5811,N_4841);
and U6757 (N_6757,N_5862,N_5849);
and U6758 (N_6758,N_5714,N_4185);
nor U6759 (N_6759,N_5087,N_4514);
and U6760 (N_6760,N_5011,N_5644);
nand U6761 (N_6761,N_4221,N_4980);
nand U6762 (N_6762,N_5677,N_4638);
nor U6763 (N_6763,N_4503,N_5609);
nand U6764 (N_6764,N_5350,N_4610);
nand U6765 (N_6765,N_4131,N_5244);
nand U6766 (N_6766,N_4823,N_5284);
nand U6767 (N_6767,N_5945,N_4312);
or U6768 (N_6768,N_4741,N_5403);
or U6769 (N_6769,N_5131,N_5962);
and U6770 (N_6770,N_5734,N_5099);
and U6771 (N_6771,N_5711,N_5543);
or U6772 (N_6772,N_5147,N_4543);
nand U6773 (N_6773,N_4328,N_5079);
nand U6774 (N_6774,N_5420,N_5494);
and U6775 (N_6775,N_4592,N_4480);
and U6776 (N_6776,N_4339,N_5909);
or U6777 (N_6777,N_4364,N_5324);
or U6778 (N_6778,N_5124,N_5626);
nor U6779 (N_6779,N_5359,N_5334);
or U6780 (N_6780,N_4813,N_5682);
nor U6781 (N_6781,N_5293,N_5245);
nand U6782 (N_6782,N_4307,N_5106);
nand U6783 (N_6783,N_4597,N_5039);
and U6784 (N_6784,N_4518,N_5614);
nor U6785 (N_6785,N_4876,N_5738);
or U6786 (N_6786,N_4552,N_5704);
or U6787 (N_6787,N_4806,N_5661);
or U6788 (N_6788,N_5502,N_5834);
nand U6789 (N_6789,N_4505,N_4820);
nor U6790 (N_6790,N_5507,N_4259);
or U6791 (N_6791,N_4925,N_4853);
or U6792 (N_6792,N_5712,N_4670);
nor U6793 (N_6793,N_4059,N_4772);
nand U6794 (N_6794,N_4286,N_4842);
and U6795 (N_6795,N_4450,N_5645);
or U6796 (N_6796,N_5327,N_4351);
nand U6797 (N_6797,N_4262,N_4648);
nand U6798 (N_6798,N_4107,N_4603);
and U6799 (N_6799,N_5846,N_4525);
nand U6800 (N_6800,N_4199,N_4618);
nor U6801 (N_6801,N_5243,N_4812);
nand U6802 (N_6802,N_5148,N_5649);
or U6803 (N_6803,N_4115,N_5062);
or U6804 (N_6804,N_4559,N_4408);
nor U6805 (N_6805,N_5944,N_4596);
or U6806 (N_6806,N_5503,N_5629);
and U6807 (N_6807,N_5250,N_5323);
and U6808 (N_6808,N_5599,N_5664);
and U6809 (N_6809,N_4650,N_5816);
or U6810 (N_6810,N_4756,N_4668);
and U6811 (N_6811,N_5304,N_4737);
nor U6812 (N_6812,N_5102,N_4045);
nor U6813 (N_6813,N_4270,N_4777);
nor U6814 (N_6814,N_5214,N_4191);
and U6815 (N_6815,N_4159,N_5193);
and U6816 (N_6816,N_4392,N_5797);
nand U6817 (N_6817,N_4052,N_5660);
and U6818 (N_6818,N_4600,N_5025);
nor U6819 (N_6819,N_5486,N_4649);
and U6820 (N_6820,N_5623,N_5201);
nand U6821 (N_6821,N_5049,N_4089);
and U6822 (N_6822,N_5895,N_4499);
or U6823 (N_6823,N_4892,N_5070);
nand U6824 (N_6824,N_5751,N_5673);
or U6825 (N_6825,N_5182,N_4712);
nor U6826 (N_6826,N_4076,N_5352);
and U6827 (N_6827,N_4451,N_5021);
nand U6828 (N_6828,N_4494,N_4169);
and U6829 (N_6829,N_5156,N_4606);
and U6830 (N_6830,N_5210,N_5574);
nor U6831 (N_6831,N_4176,N_4422);
nor U6832 (N_6832,N_4968,N_4796);
nor U6833 (N_6833,N_4970,N_4544);
nand U6834 (N_6834,N_4634,N_5367);
or U6835 (N_6835,N_4614,N_4517);
nor U6836 (N_6836,N_5762,N_4973);
and U6837 (N_6837,N_5445,N_4497);
nor U6838 (N_6838,N_5658,N_5060);
and U6839 (N_6839,N_4780,N_4461);
and U6840 (N_6840,N_4184,N_5784);
nand U6841 (N_6841,N_4539,N_5708);
nor U6842 (N_6842,N_4256,N_4673);
or U6843 (N_6843,N_4821,N_5174);
nor U6844 (N_6844,N_4929,N_5080);
nor U6845 (N_6845,N_4939,N_5561);
and U6846 (N_6846,N_4987,N_5383);
nor U6847 (N_6847,N_4455,N_4401);
nand U6848 (N_6848,N_4851,N_5829);
nor U6849 (N_6849,N_4057,N_5116);
nor U6850 (N_6850,N_4335,N_4587);
and U6851 (N_6851,N_4406,N_4642);
nor U6852 (N_6852,N_4616,N_5595);
nand U6853 (N_6853,N_4900,N_4472);
nand U6854 (N_6854,N_5240,N_5374);
nand U6855 (N_6855,N_5570,N_4055);
or U6856 (N_6856,N_4658,N_5536);
and U6857 (N_6857,N_5152,N_4465);
nor U6858 (N_6858,N_4837,N_5198);
nor U6859 (N_6859,N_5923,N_4300);
or U6860 (N_6860,N_4030,N_4474);
nand U6861 (N_6861,N_5975,N_4211);
nor U6862 (N_6862,N_5518,N_4938);
or U6863 (N_6863,N_5342,N_4574);
or U6864 (N_6864,N_4691,N_4875);
and U6865 (N_6865,N_5709,N_4697);
nand U6866 (N_6866,N_4092,N_5566);
nand U6867 (N_6867,N_4736,N_5913);
nor U6868 (N_6868,N_5840,N_5238);
nand U6869 (N_6869,N_5748,N_4946);
or U6870 (N_6870,N_4542,N_5040);
and U6871 (N_6871,N_4075,N_4508);
nor U6872 (N_6872,N_4232,N_4407);
nor U6873 (N_6873,N_4433,N_4234);
nand U6874 (N_6874,N_5510,N_5392);
or U6875 (N_6875,N_4832,N_4602);
or U6876 (N_6876,N_5772,N_5524);
nor U6877 (N_6877,N_4037,N_5887);
nand U6878 (N_6878,N_5271,N_5921);
or U6879 (N_6879,N_4893,N_5788);
nand U6880 (N_6880,N_5405,N_5388);
and U6881 (N_6881,N_4678,N_4507);
or U6882 (N_6882,N_5415,N_5065);
and U6883 (N_6883,N_5505,N_5399);
nor U6884 (N_6884,N_4215,N_4269);
and U6885 (N_6885,N_4027,N_4393);
and U6886 (N_6886,N_5656,N_5960);
nand U6887 (N_6887,N_5481,N_5072);
nand U6888 (N_6888,N_5990,N_5753);
or U6889 (N_6889,N_5779,N_5053);
and U6890 (N_6890,N_5172,N_5646);
or U6891 (N_6891,N_5651,N_5450);
nor U6892 (N_6892,N_5013,N_4767);
or U6893 (N_6893,N_5908,N_5386);
nor U6894 (N_6894,N_5508,N_4170);
nand U6895 (N_6895,N_5871,N_4424);
nand U6896 (N_6896,N_5054,N_5928);
and U6897 (N_6897,N_5724,N_4316);
and U6898 (N_6898,N_4789,N_5957);
nand U6899 (N_6899,N_4318,N_5537);
or U6900 (N_6900,N_4492,N_5722);
nor U6901 (N_6901,N_5564,N_4835);
or U6902 (N_6902,N_5278,N_5290);
and U6903 (N_6903,N_4623,N_4529);
nor U6904 (N_6904,N_5747,N_4556);
and U6905 (N_6905,N_5584,N_4621);
or U6906 (N_6906,N_4951,N_5924);
nor U6907 (N_6907,N_5723,N_5033);
nand U6908 (N_6908,N_4561,N_4303);
and U6909 (N_6909,N_4810,N_5821);
or U6910 (N_6910,N_5839,N_5224);
nor U6911 (N_6911,N_5590,N_5756);
or U6912 (N_6912,N_5423,N_5979);
and U6913 (N_6913,N_5295,N_5001);
or U6914 (N_6914,N_5167,N_4745);
or U6915 (N_6915,N_4862,N_4896);
nor U6916 (N_6916,N_4500,N_5684);
nor U6917 (N_6917,N_4786,N_5692);
xnor U6918 (N_6918,N_4857,N_5989);
nand U6919 (N_6919,N_4295,N_4350);
nor U6920 (N_6920,N_4844,N_5197);
and U6921 (N_6921,N_5006,N_5653);
and U6922 (N_6922,N_4811,N_5348);
nor U6923 (N_6923,N_4725,N_5718);
or U6924 (N_6924,N_5814,N_4738);
nor U6925 (N_6925,N_4976,N_4732);
nand U6926 (N_6926,N_4308,N_4659);
nand U6927 (N_6927,N_4915,N_4367);
and U6928 (N_6928,N_5613,N_5985);
and U6929 (N_6929,N_5491,N_5205);
nor U6930 (N_6930,N_4510,N_4586);
and U6931 (N_6931,N_5059,N_4880);
or U6932 (N_6932,N_5627,N_5879);
and U6933 (N_6933,N_4206,N_5509);
and U6934 (N_6934,N_4025,N_5534);
or U6935 (N_6935,N_5427,N_5169);
nand U6936 (N_6936,N_5556,N_4828);
nor U6937 (N_6937,N_5934,N_5547);
or U6938 (N_6938,N_4923,N_5406);
or U6939 (N_6939,N_4906,N_5030);
nand U6940 (N_6940,N_4687,N_5176);
or U6941 (N_6941,N_4365,N_4626);
nor U6942 (N_6942,N_4762,N_5836);
or U6943 (N_6943,N_4292,N_4201);
nor U6944 (N_6944,N_4957,N_5693);
and U6945 (N_6945,N_4674,N_5204);
or U6946 (N_6946,N_4916,N_4704);
nor U6947 (N_6947,N_5468,N_4178);
nor U6948 (N_6948,N_4940,N_4800);
nor U6949 (N_6949,N_4719,N_4209);
or U6950 (N_6950,N_5441,N_5055);
and U6951 (N_6951,N_4954,N_5891);
nor U6952 (N_6952,N_5796,N_4943);
nand U6953 (N_6953,N_4331,N_5333);
nor U6954 (N_6954,N_4297,N_5017);
or U6955 (N_6955,N_5987,N_5888);
and U6956 (N_6956,N_4186,N_4466);
and U6957 (N_6957,N_4157,N_5432);
and U6958 (N_6958,N_5689,N_4448);
and U6959 (N_6959,N_4863,N_4950);
and U6960 (N_6960,N_5845,N_5187);
or U6961 (N_6961,N_4703,N_5337);
nor U6962 (N_6962,N_5029,N_4708);
nand U6963 (N_6963,N_4305,N_4258);
and U6964 (N_6964,N_4989,N_5377);
or U6965 (N_6965,N_5142,N_5381);
or U6966 (N_6966,N_5344,N_4867);
nor U6967 (N_6967,N_4944,N_4353);
or U6968 (N_6968,N_4849,N_5706);
and U6969 (N_6969,N_5807,N_5146);
or U6970 (N_6970,N_5285,N_4077);
nand U6971 (N_6971,N_4677,N_4794);
or U6972 (N_6972,N_4717,N_4090);
nor U6973 (N_6973,N_4919,N_4342);
and U6974 (N_6974,N_5014,N_4218);
nand U6975 (N_6975,N_4103,N_5643);
nand U6976 (N_6976,N_4858,N_4457);
nand U6977 (N_6977,N_5577,N_4405);
nor U6978 (N_6978,N_4345,N_5356);
nand U6979 (N_6979,N_4000,N_5370);
nand U6980 (N_6980,N_4643,N_5890);
nor U6981 (N_6981,N_4942,N_4071);
or U6982 (N_6982,N_5539,N_5056);
or U6983 (N_6983,N_5289,N_5082);
or U6984 (N_6984,N_5078,N_5641);
or U6985 (N_6985,N_5496,N_5426);
xnor U6986 (N_6986,N_5806,N_4843);
nor U6987 (N_6987,N_5424,N_5084);
nand U6988 (N_6988,N_5769,N_5354);
nand U6989 (N_6989,N_5385,N_5031);
nor U6990 (N_6990,N_5117,N_5007);
nand U6991 (N_6991,N_4008,N_4680);
nor U6992 (N_6992,N_5408,N_5707);
or U6993 (N_6993,N_4285,N_4477);
xnor U6994 (N_6994,N_4402,N_5097);
nor U6995 (N_6995,N_5389,N_4560);
or U6996 (N_6996,N_5294,N_4890);
and U6997 (N_6997,N_4898,N_4222);
nand U6998 (N_6998,N_5898,N_4748);
xnor U6999 (N_6999,N_5996,N_5024);
nor U7000 (N_7000,N_4981,N_5235);
nor U7001 (N_7001,N_5779,N_5613);
and U7002 (N_7002,N_4410,N_4971);
and U7003 (N_7003,N_5961,N_4568);
and U7004 (N_7004,N_4838,N_5162);
and U7005 (N_7005,N_5955,N_4287);
nand U7006 (N_7006,N_4957,N_4462);
nand U7007 (N_7007,N_5574,N_5661);
or U7008 (N_7008,N_5519,N_4263);
nand U7009 (N_7009,N_5762,N_5877);
nand U7010 (N_7010,N_5112,N_5517);
nand U7011 (N_7011,N_5124,N_5582);
or U7012 (N_7012,N_5573,N_5830);
nand U7013 (N_7013,N_5477,N_5149);
nand U7014 (N_7014,N_5601,N_5378);
and U7015 (N_7015,N_4854,N_5300);
or U7016 (N_7016,N_5842,N_5947);
nand U7017 (N_7017,N_4614,N_5994);
nor U7018 (N_7018,N_5573,N_5366);
xor U7019 (N_7019,N_5706,N_4202);
and U7020 (N_7020,N_4308,N_4229);
nor U7021 (N_7021,N_4999,N_5892);
and U7022 (N_7022,N_4570,N_4282);
and U7023 (N_7023,N_4881,N_5588);
nor U7024 (N_7024,N_4478,N_4976);
nand U7025 (N_7025,N_5799,N_5476);
nor U7026 (N_7026,N_5282,N_5544);
and U7027 (N_7027,N_5768,N_5724);
and U7028 (N_7028,N_4310,N_5025);
nand U7029 (N_7029,N_4937,N_4876);
and U7030 (N_7030,N_5468,N_4573);
or U7031 (N_7031,N_5794,N_4407);
nand U7032 (N_7032,N_4636,N_4758);
nor U7033 (N_7033,N_4911,N_4330);
nand U7034 (N_7034,N_4518,N_5179);
nand U7035 (N_7035,N_5499,N_4659);
nand U7036 (N_7036,N_5378,N_4081);
nor U7037 (N_7037,N_4678,N_5188);
and U7038 (N_7038,N_5109,N_4340);
or U7039 (N_7039,N_5283,N_5484);
and U7040 (N_7040,N_5256,N_4776);
nor U7041 (N_7041,N_5047,N_5566);
nand U7042 (N_7042,N_5180,N_4238);
nor U7043 (N_7043,N_5786,N_5616);
nor U7044 (N_7044,N_5624,N_5666);
nor U7045 (N_7045,N_5279,N_4981);
nand U7046 (N_7046,N_5397,N_5691);
and U7047 (N_7047,N_5434,N_4978);
and U7048 (N_7048,N_5564,N_5414);
or U7049 (N_7049,N_5190,N_4506);
nor U7050 (N_7050,N_5287,N_4298);
nor U7051 (N_7051,N_4649,N_4100);
or U7052 (N_7052,N_5203,N_4406);
and U7053 (N_7053,N_5825,N_5336);
nor U7054 (N_7054,N_4502,N_4359);
and U7055 (N_7055,N_4043,N_5175);
nor U7056 (N_7056,N_4824,N_4049);
nand U7057 (N_7057,N_5706,N_5493);
and U7058 (N_7058,N_4678,N_4534);
nor U7059 (N_7059,N_4676,N_5639);
or U7060 (N_7060,N_5993,N_4535);
nand U7061 (N_7061,N_4538,N_5045);
or U7062 (N_7062,N_4635,N_4752);
nor U7063 (N_7063,N_4806,N_5877);
and U7064 (N_7064,N_4599,N_5598);
nand U7065 (N_7065,N_4252,N_4413);
and U7066 (N_7066,N_4362,N_4654);
or U7067 (N_7067,N_4410,N_4146);
nand U7068 (N_7068,N_4663,N_5437);
nor U7069 (N_7069,N_4771,N_5834);
or U7070 (N_7070,N_5007,N_5096);
and U7071 (N_7071,N_4368,N_4702);
nand U7072 (N_7072,N_4597,N_5980);
and U7073 (N_7073,N_4675,N_5113);
and U7074 (N_7074,N_5803,N_5572);
nor U7075 (N_7075,N_5619,N_5961);
or U7076 (N_7076,N_5522,N_5422);
xnor U7077 (N_7077,N_4804,N_4873);
and U7078 (N_7078,N_5372,N_5071);
and U7079 (N_7079,N_4000,N_5706);
nor U7080 (N_7080,N_4747,N_5514);
and U7081 (N_7081,N_5939,N_4119);
nor U7082 (N_7082,N_5381,N_5875);
and U7083 (N_7083,N_5946,N_4611);
nor U7084 (N_7084,N_4363,N_4316);
or U7085 (N_7085,N_5882,N_5497);
or U7086 (N_7086,N_4092,N_5737);
or U7087 (N_7087,N_5782,N_4860);
nor U7088 (N_7088,N_4243,N_4837);
nor U7089 (N_7089,N_4179,N_4290);
nor U7090 (N_7090,N_5926,N_4425);
or U7091 (N_7091,N_4896,N_5512);
nand U7092 (N_7092,N_4158,N_4933);
xor U7093 (N_7093,N_4995,N_5479);
or U7094 (N_7094,N_4178,N_4909);
nor U7095 (N_7095,N_4402,N_4189);
nand U7096 (N_7096,N_5571,N_5797);
or U7097 (N_7097,N_5998,N_5645);
and U7098 (N_7098,N_5264,N_5170);
or U7099 (N_7099,N_5680,N_4881);
and U7100 (N_7100,N_5023,N_5149);
and U7101 (N_7101,N_5499,N_4298);
nor U7102 (N_7102,N_4252,N_5307);
and U7103 (N_7103,N_5350,N_4056);
nor U7104 (N_7104,N_4667,N_4766);
and U7105 (N_7105,N_5624,N_4801);
nand U7106 (N_7106,N_5854,N_4878);
and U7107 (N_7107,N_5173,N_5756);
nand U7108 (N_7108,N_4335,N_5664);
or U7109 (N_7109,N_5623,N_5141);
nor U7110 (N_7110,N_5661,N_5952);
and U7111 (N_7111,N_4551,N_5932);
nor U7112 (N_7112,N_5008,N_4020);
and U7113 (N_7113,N_4982,N_5502);
nor U7114 (N_7114,N_4433,N_4944);
or U7115 (N_7115,N_5612,N_4819);
or U7116 (N_7116,N_5814,N_4626);
nand U7117 (N_7117,N_5550,N_5589);
and U7118 (N_7118,N_4791,N_4476);
nand U7119 (N_7119,N_4982,N_4118);
nand U7120 (N_7120,N_4227,N_5073);
and U7121 (N_7121,N_4785,N_5489);
nand U7122 (N_7122,N_5560,N_4513);
or U7123 (N_7123,N_4004,N_5295);
or U7124 (N_7124,N_5128,N_4812);
and U7125 (N_7125,N_4961,N_5873);
and U7126 (N_7126,N_4458,N_5910);
nor U7127 (N_7127,N_5270,N_5089);
or U7128 (N_7128,N_5572,N_5029);
or U7129 (N_7129,N_4122,N_5858);
nor U7130 (N_7130,N_4546,N_4517);
nand U7131 (N_7131,N_4296,N_4426);
or U7132 (N_7132,N_4129,N_4623);
and U7133 (N_7133,N_5497,N_4694);
nand U7134 (N_7134,N_5641,N_4870);
and U7135 (N_7135,N_5798,N_4989);
and U7136 (N_7136,N_5568,N_5210);
nor U7137 (N_7137,N_5527,N_5084);
and U7138 (N_7138,N_5573,N_5797);
or U7139 (N_7139,N_5797,N_4335);
nand U7140 (N_7140,N_4767,N_5700);
or U7141 (N_7141,N_5780,N_4416);
and U7142 (N_7142,N_4793,N_5143);
nand U7143 (N_7143,N_5498,N_4932);
xnor U7144 (N_7144,N_5594,N_5358);
nand U7145 (N_7145,N_5259,N_5232);
and U7146 (N_7146,N_5367,N_4194);
or U7147 (N_7147,N_5378,N_4579);
nand U7148 (N_7148,N_5659,N_4654);
and U7149 (N_7149,N_4148,N_4314);
nand U7150 (N_7150,N_5095,N_4676);
nor U7151 (N_7151,N_4487,N_4439);
nand U7152 (N_7152,N_4124,N_5296);
or U7153 (N_7153,N_4128,N_5686);
nand U7154 (N_7154,N_4651,N_4086);
or U7155 (N_7155,N_5294,N_5747);
or U7156 (N_7156,N_4582,N_4151);
and U7157 (N_7157,N_4004,N_5990);
nand U7158 (N_7158,N_4411,N_5683);
nor U7159 (N_7159,N_5000,N_5186);
or U7160 (N_7160,N_5916,N_4072);
nand U7161 (N_7161,N_5316,N_5308);
nor U7162 (N_7162,N_4452,N_5245);
or U7163 (N_7163,N_5333,N_4208);
and U7164 (N_7164,N_4202,N_5635);
and U7165 (N_7165,N_5690,N_5888);
nand U7166 (N_7166,N_4228,N_4119);
nand U7167 (N_7167,N_4523,N_4955);
nand U7168 (N_7168,N_4027,N_5008);
and U7169 (N_7169,N_4549,N_5851);
or U7170 (N_7170,N_4862,N_4331);
nor U7171 (N_7171,N_4324,N_5084);
nor U7172 (N_7172,N_5777,N_4026);
nand U7173 (N_7173,N_4607,N_4410);
or U7174 (N_7174,N_4640,N_5726);
nor U7175 (N_7175,N_4585,N_4052);
nand U7176 (N_7176,N_5712,N_5196);
nor U7177 (N_7177,N_5661,N_5967);
and U7178 (N_7178,N_4730,N_4880);
nor U7179 (N_7179,N_4085,N_5017);
nand U7180 (N_7180,N_4895,N_4107);
xnor U7181 (N_7181,N_4795,N_5818);
and U7182 (N_7182,N_5253,N_5493);
and U7183 (N_7183,N_5319,N_5444);
or U7184 (N_7184,N_5529,N_5749);
nor U7185 (N_7185,N_4281,N_4459);
and U7186 (N_7186,N_4120,N_5160);
nor U7187 (N_7187,N_4396,N_4322);
and U7188 (N_7188,N_4108,N_4933);
or U7189 (N_7189,N_4502,N_4813);
or U7190 (N_7190,N_4787,N_4362);
and U7191 (N_7191,N_4947,N_5970);
and U7192 (N_7192,N_4051,N_4882);
nand U7193 (N_7193,N_4254,N_5331);
or U7194 (N_7194,N_4066,N_5586);
nand U7195 (N_7195,N_5201,N_5717);
nor U7196 (N_7196,N_4397,N_5407);
nand U7197 (N_7197,N_4073,N_4362);
and U7198 (N_7198,N_4158,N_4580);
and U7199 (N_7199,N_5299,N_4472);
or U7200 (N_7200,N_5507,N_5974);
or U7201 (N_7201,N_4479,N_5329);
or U7202 (N_7202,N_4993,N_4764);
and U7203 (N_7203,N_5744,N_5404);
or U7204 (N_7204,N_5257,N_4697);
or U7205 (N_7205,N_5976,N_5847);
nor U7206 (N_7206,N_4595,N_4129);
and U7207 (N_7207,N_4772,N_4420);
nor U7208 (N_7208,N_5711,N_4565);
and U7209 (N_7209,N_5811,N_4661);
nand U7210 (N_7210,N_4906,N_4219);
nand U7211 (N_7211,N_5352,N_5971);
and U7212 (N_7212,N_5034,N_5328);
nor U7213 (N_7213,N_4880,N_5812);
or U7214 (N_7214,N_4989,N_4657);
nor U7215 (N_7215,N_4339,N_5779);
nor U7216 (N_7216,N_4085,N_4406);
and U7217 (N_7217,N_4963,N_5192);
nor U7218 (N_7218,N_4221,N_4835);
nand U7219 (N_7219,N_4024,N_5953);
xnor U7220 (N_7220,N_4840,N_4328);
or U7221 (N_7221,N_5364,N_4499);
nand U7222 (N_7222,N_5556,N_5629);
nand U7223 (N_7223,N_5488,N_5652);
and U7224 (N_7224,N_4069,N_4834);
or U7225 (N_7225,N_4500,N_5168);
nor U7226 (N_7226,N_4941,N_5394);
nor U7227 (N_7227,N_4066,N_4480);
nor U7228 (N_7228,N_5736,N_4656);
nor U7229 (N_7229,N_4376,N_4667);
or U7230 (N_7230,N_4041,N_4093);
and U7231 (N_7231,N_5115,N_5403);
nand U7232 (N_7232,N_5049,N_5291);
nor U7233 (N_7233,N_5761,N_5412);
nor U7234 (N_7234,N_4965,N_5260);
or U7235 (N_7235,N_4109,N_5839);
nand U7236 (N_7236,N_4612,N_5831);
nand U7237 (N_7237,N_5326,N_4238);
nor U7238 (N_7238,N_4363,N_5192);
or U7239 (N_7239,N_4986,N_5700);
and U7240 (N_7240,N_5659,N_4330);
or U7241 (N_7241,N_4117,N_4194);
and U7242 (N_7242,N_5193,N_4172);
nand U7243 (N_7243,N_4840,N_5276);
or U7244 (N_7244,N_4591,N_5292);
nand U7245 (N_7245,N_4805,N_4521);
nand U7246 (N_7246,N_4848,N_5108);
or U7247 (N_7247,N_4303,N_4110);
or U7248 (N_7248,N_4500,N_5900);
and U7249 (N_7249,N_5571,N_4720);
nor U7250 (N_7250,N_5008,N_5812);
or U7251 (N_7251,N_4570,N_5772);
and U7252 (N_7252,N_4842,N_4459);
nand U7253 (N_7253,N_4684,N_4260);
xor U7254 (N_7254,N_4908,N_4212);
nor U7255 (N_7255,N_5180,N_5877);
and U7256 (N_7256,N_4226,N_5706);
and U7257 (N_7257,N_4917,N_5621);
nand U7258 (N_7258,N_4369,N_4582);
and U7259 (N_7259,N_4358,N_5858);
nor U7260 (N_7260,N_5326,N_5976);
nand U7261 (N_7261,N_5927,N_5905);
or U7262 (N_7262,N_5632,N_4842);
and U7263 (N_7263,N_4160,N_4178);
or U7264 (N_7264,N_5385,N_5607);
or U7265 (N_7265,N_5389,N_5539);
nor U7266 (N_7266,N_4569,N_5801);
and U7267 (N_7267,N_5068,N_5200);
or U7268 (N_7268,N_4673,N_5397);
or U7269 (N_7269,N_4658,N_4642);
nor U7270 (N_7270,N_5917,N_4886);
nand U7271 (N_7271,N_5387,N_4915);
nor U7272 (N_7272,N_5787,N_4813);
and U7273 (N_7273,N_4881,N_4332);
nor U7274 (N_7274,N_5352,N_5208);
nand U7275 (N_7275,N_4755,N_5283);
and U7276 (N_7276,N_5252,N_4129);
nor U7277 (N_7277,N_4301,N_4359);
and U7278 (N_7278,N_5661,N_4642);
nor U7279 (N_7279,N_4944,N_4587);
nor U7280 (N_7280,N_4759,N_4547);
or U7281 (N_7281,N_5386,N_5682);
nor U7282 (N_7282,N_4668,N_5354);
or U7283 (N_7283,N_4970,N_5995);
nor U7284 (N_7284,N_4915,N_4276);
or U7285 (N_7285,N_5376,N_4083);
nor U7286 (N_7286,N_5157,N_5270);
or U7287 (N_7287,N_4049,N_4466);
nand U7288 (N_7288,N_5990,N_5303);
and U7289 (N_7289,N_4955,N_4091);
and U7290 (N_7290,N_4078,N_5993);
or U7291 (N_7291,N_4900,N_4377);
nor U7292 (N_7292,N_4763,N_4446);
nand U7293 (N_7293,N_5142,N_4709);
and U7294 (N_7294,N_5866,N_5307);
nor U7295 (N_7295,N_4826,N_5609);
nand U7296 (N_7296,N_5683,N_5715);
nand U7297 (N_7297,N_5944,N_4014);
nor U7298 (N_7298,N_5867,N_5907);
or U7299 (N_7299,N_4686,N_5297);
and U7300 (N_7300,N_4770,N_4621);
xor U7301 (N_7301,N_5363,N_4874);
and U7302 (N_7302,N_5583,N_5122);
and U7303 (N_7303,N_4099,N_4852);
and U7304 (N_7304,N_5805,N_5465);
nand U7305 (N_7305,N_5456,N_4216);
and U7306 (N_7306,N_5160,N_4129);
nor U7307 (N_7307,N_4814,N_4603);
or U7308 (N_7308,N_4571,N_4071);
and U7309 (N_7309,N_5186,N_5310);
xor U7310 (N_7310,N_5840,N_4964);
nor U7311 (N_7311,N_5979,N_4106);
and U7312 (N_7312,N_5438,N_5134);
or U7313 (N_7313,N_5652,N_5964);
nand U7314 (N_7314,N_4550,N_5456);
or U7315 (N_7315,N_4811,N_5243);
nand U7316 (N_7316,N_5414,N_5070);
nand U7317 (N_7317,N_5549,N_4096);
nand U7318 (N_7318,N_4208,N_4168);
and U7319 (N_7319,N_5315,N_4714);
nor U7320 (N_7320,N_4833,N_5626);
and U7321 (N_7321,N_4257,N_4720);
and U7322 (N_7322,N_5501,N_4818);
nand U7323 (N_7323,N_4093,N_5549);
or U7324 (N_7324,N_4094,N_5697);
and U7325 (N_7325,N_5053,N_4659);
and U7326 (N_7326,N_5898,N_4445);
nor U7327 (N_7327,N_4883,N_4310);
or U7328 (N_7328,N_5039,N_4594);
and U7329 (N_7329,N_5238,N_5113);
nand U7330 (N_7330,N_5171,N_4235);
nand U7331 (N_7331,N_5236,N_4993);
nand U7332 (N_7332,N_5310,N_4999);
or U7333 (N_7333,N_4987,N_4822);
and U7334 (N_7334,N_5980,N_5100);
or U7335 (N_7335,N_4641,N_4924);
nor U7336 (N_7336,N_5632,N_5332);
and U7337 (N_7337,N_5840,N_4819);
or U7338 (N_7338,N_5409,N_4456);
and U7339 (N_7339,N_5707,N_5497);
nand U7340 (N_7340,N_5195,N_5336);
or U7341 (N_7341,N_5653,N_5801);
nand U7342 (N_7342,N_5737,N_5859);
nand U7343 (N_7343,N_4747,N_5902);
nor U7344 (N_7344,N_4131,N_5281);
nand U7345 (N_7345,N_4286,N_5601);
xor U7346 (N_7346,N_4768,N_4354);
nor U7347 (N_7347,N_5140,N_4374);
or U7348 (N_7348,N_4041,N_5081);
nand U7349 (N_7349,N_5980,N_4804);
and U7350 (N_7350,N_4914,N_4846);
or U7351 (N_7351,N_5820,N_5805);
nor U7352 (N_7352,N_5505,N_4666);
nand U7353 (N_7353,N_4547,N_4373);
nand U7354 (N_7354,N_4448,N_4502);
or U7355 (N_7355,N_4353,N_5981);
nand U7356 (N_7356,N_4072,N_5219);
and U7357 (N_7357,N_5520,N_5794);
or U7358 (N_7358,N_5142,N_4864);
or U7359 (N_7359,N_5095,N_4031);
nand U7360 (N_7360,N_5697,N_4842);
nor U7361 (N_7361,N_5765,N_4120);
and U7362 (N_7362,N_5698,N_4180);
and U7363 (N_7363,N_5115,N_5576);
and U7364 (N_7364,N_4421,N_4963);
or U7365 (N_7365,N_4473,N_5544);
nand U7366 (N_7366,N_5604,N_4883);
or U7367 (N_7367,N_4456,N_4876);
or U7368 (N_7368,N_4973,N_4256);
nor U7369 (N_7369,N_5486,N_5733);
or U7370 (N_7370,N_5138,N_5247);
or U7371 (N_7371,N_5396,N_4047);
and U7372 (N_7372,N_4413,N_4087);
nor U7373 (N_7373,N_5047,N_5804);
or U7374 (N_7374,N_5184,N_5183);
or U7375 (N_7375,N_4268,N_5217);
nor U7376 (N_7376,N_5648,N_5085);
nor U7377 (N_7377,N_5486,N_4074);
or U7378 (N_7378,N_5787,N_5455);
or U7379 (N_7379,N_4326,N_4226);
nor U7380 (N_7380,N_4079,N_5891);
or U7381 (N_7381,N_4035,N_4811);
nand U7382 (N_7382,N_4654,N_5073);
nand U7383 (N_7383,N_4422,N_4756);
nand U7384 (N_7384,N_5481,N_4488);
and U7385 (N_7385,N_5103,N_4157);
and U7386 (N_7386,N_5935,N_4223);
and U7387 (N_7387,N_5490,N_5133);
and U7388 (N_7388,N_5594,N_4747);
nand U7389 (N_7389,N_5923,N_5901);
and U7390 (N_7390,N_5934,N_4867);
and U7391 (N_7391,N_4526,N_4144);
nor U7392 (N_7392,N_5294,N_5718);
or U7393 (N_7393,N_4633,N_5292);
or U7394 (N_7394,N_5954,N_5222);
or U7395 (N_7395,N_5819,N_4816);
nand U7396 (N_7396,N_5702,N_5627);
nor U7397 (N_7397,N_5476,N_4110);
and U7398 (N_7398,N_4899,N_5366);
and U7399 (N_7399,N_4712,N_4963);
nand U7400 (N_7400,N_5685,N_4329);
nor U7401 (N_7401,N_5881,N_4588);
and U7402 (N_7402,N_5390,N_5792);
nor U7403 (N_7403,N_5031,N_5663);
and U7404 (N_7404,N_5452,N_4801);
or U7405 (N_7405,N_4316,N_4528);
nor U7406 (N_7406,N_4865,N_5613);
or U7407 (N_7407,N_5862,N_4509);
nor U7408 (N_7408,N_4033,N_4271);
nand U7409 (N_7409,N_4269,N_5167);
xnor U7410 (N_7410,N_4407,N_4812);
or U7411 (N_7411,N_4425,N_4113);
and U7412 (N_7412,N_5586,N_5169);
and U7413 (N_7413,N_5090,N_5780);
nand U7414 (N_7414,N_5034,N_5340);
and U7415 (N_7415,N_4467,N_5881);
nand U7416 (N_7416,N_4938,N_5446);
and U7417 (N_7417,N_4678,N_4356);
and U7418 (N_7418,N_5548,N_4944);
or U7419 (N_7419,N_4131,N_5317);
and U7420 (N_7420,N_4747,N_4352);
and U7421 (N_7421,N_4667,N_4501);
nor U7422 (N_7422,N_4926,N_5516);
or U7423 (N_7423,N_4328,N_5104);
nand U7424 (N_7424,N_5506,N_5790);
or U7425 (N_7425,N_4708,N_4866);
nor U7426 (N_7426,N_4333,N_4961);
and U7427 (N_7427,N_4783,N_4859);
and U7428 (N_7428,N_4390,N_5972);
and U7429 (N_7429,N_4635,N_5156);
or U7430 (N_7430,N_4772,N_4294);
and U7431 (N_7431,N_4036,N_5428);
and U7432 (N_7432,N_5376,N_4209);
nand U7433 (N_7433,N_5345,N_4790);
nand U7434 (N_7434,N_4850,N_5111);
nor U7435 (N_7435,N_5039,N_4937);
or U7436 (N_7436,N_4872,N_5073);
xor U7437 (N_7437,N_5605,N_4832);
and U7438 (N_7438,N_4349,N_5002);
and U7439 (N_7439,N_4624,N_5046);
and U7440 (N_7440,N_4510,N_4077);
or U7441 (N_7441,N_4732,N_5792);
nand U7442 (N_7442,N_4014,N_5489);
and U7443 (N_7443,N_5024,N_5252);
or U7444 (N_7444,N_5066,N_5796);
and U7445 (N_7445,N_5376,N_5410);
nor U7446 (N_7446,N_5374,N_5917);
nand U7447 (N_7447,N_5494,N_4131);
nand U7448 (N_7448,N_4288,N_4133);
and U7449 (N_7449,N_4977,N_4347);
nor U7450 (N_7450,N_5303,N_4509);
and U7451 (N_7451,N_4014,N_5179);
and U7452 (N_7452,N_5622,N_4069);
nor U7453 (N_7453,N_4109,N_4112);
nand U7454 (N_7454,N_4748,N_4929);
nor U7455 (N_7455,N_5157,N_4845);
nor U7456 (N_7456,N_5940,N_4665);
nand U7457 (N_7457,N_5515,N_5169);
and U7458 (N_7458,N_4192,N_4430);
or U7459 (N_7459,N_4343,N_5970);
and U7460 (N_7460,N_5755,N_5796);
or U7461 (N_7461,N_5664,N_4068);
nor U7462 (N_7462,N_5354,N_5451);
or U7463 (N_7463,N_4224,N_5900);
nor U7464 (N_7464,N_5326,N_4885);
nor U7465 (N_7465,N_4698,N_5436);
nand U7466 (N_7466,N_4018,N_4845);
nor U7467 (N_7467,N_5584,N_4445);
and U7468 (N_7468,N_4007,N_4619);
nand U7469 (N_7469,N_4101,N_5633);
and U7470 (N_7470,N_4095,N_5864);
and U7471 (N_7471,N_4233,N_5807);
xor U7472 (N_7472,N_5609,N_4666);
and U7473 (N_7473,N_5770,N_4803);
and U7474 (N_7474,N_4398,N_5188);
nand U7475 (N_7475,N_5646,N_5109);
and U7476 (N_7476,N_5602,N_5530);
nand U7477 (N_7477,N_5303,N_4663);
nor U7478 (N_7478,N_4504,N_4035);
or U7479 (N_7479,N_4707,N_5149);
nor U7480 (N_7480,N_4512,N_5270);
nor U7481 (N_7481,N_5024,N_5062);
nand U7482 (N_7482,N_5624,N_5937);
nand U7483 (N_7483,N_5225,N_5558);
nor U7484 (N_7484,N_5116,N_5021);
and U7485 (N_7485,N_5458,N_4167);
nand U7486 (N_7486,N_4413,N_4538);
and U7487 (N_7487,N_4041,N_4708);
nor U7488 (N_7488,N_5642,N_4536);
and U7489 (N_7489,N_4725,N_4915);
nand U7490 (N_7490,N_5940,N_4603);
nand U7491 (N_7491,N_5664,N_5613);
nor U7492 (N_7492,N_5291,N_4717);
nor U7493 (N_7493,N_4859,N_4096);
nand U7494 (N_7494,N_4247,N_4174);
nor U7495 (N_7495,N_4694,N_4538);
or U7496 (N_7496,N_5679,N_4737);
nor U7497 (N_7497,N_4138,N_5730);
and U7498 (N_7498,N_5091,N_4838);
nand U7499 (N_7499,N_5629,N_4853);
nor U7500 (N_7500,N_4799,N_4419);
nor U7501 (N_7501,N_4151,N_4737);
or U7502 (N_7502,N_5475,N_4022);
nand U7503 (N_7503,N_5660,N_4492);
nor U7504 (N_7504,N_5332,N_4705);
or U7505 (N_7505,N_4085,N_4225);
and U7506 (N_7506,N_5838,N_4611);
nand U7507 (N_7507,N_4112,N_4749);
nor U7508 (N_7508,N_4397,N_5919);
and U7509 (N_7509,N_4646,N_5507);
and U7510 (N_7510,N_4364,N_5759);
or U7511 (N_7511,N_4873,N_5433);
or U7512 (N_7512,N_5719,N_5704);
nor U7513 (N_7513,N_5556,N_5218);
nor U7514 (N_7514,N_5167,N_4606);
nand U7515 (N_7515,N_4015,N_5815);
or U7516 (N_7516,N_4274,N_4874);
and U7517 (N_7517,N_5692,N_5651);
nand U7518 (N_7518,N_5570,N_4403);
nand U7519 (N_7519,N_5669,N_5503);
or U7520 (N_7520,N_5424,N_4082);
nor U7521 (N_7521,N_4778,N_4634);
nor U7522 (N_7522,N_5043,N_4890);
nor U7523 (N_7523,N_4063,N_5880);
or U7524 (N_7524,N_4512,N_5167);
or U7525 (N_7525,N_4172,N_4153);
and U7526 (N_7526,N_4155,N_5442);
or U7527 (N_7527,N_5168,N_5936);
nand U7528 (N_7528,N_4946,N_4468);
or U7529 (N_7529,N_4226,N_4741);
nand U7530 (N_7530,N_4964,N_4076);
or U7531 (N_7531,N_5380,N_5431);
nand U7532 (N_7532,N_5602,N_4639);
or U7533 (N_7533,N_4230,N_5630);
or U7534 (N_7534,N_5907,N_5008);
nor U7535 (N_7535,N_5036,N_4469);
or U7536 (N_7536,N_5524,N_4277);
or U7537 (N_7537,N_5218,N_4985);
nand U7538 (N_7538,N_5776,N_4349);
and U7539 (N_7539,N_5659,N_5641);
nor U7540 (N_7540,N_5195,N_5289);
and U7541 (N_7541,N_4448,N_5842);
and U7542 (N_7542,N_5760,N_4477);
or U7543 (N_7543,N_5006,N_5707);
or U7544 (N_7544,N_5768,N_4546);
nor U7545 (N_7545,N_4576,N_5353);
nor U7546 (N_7546,N_4865,N_5564);
or U7547 (N_7547,N_4556,N_5847);
nor U7548 (N_7548,N_5580,N_5961);
nor U7549 (N_7549,N_4358,N_5929);
xnor U7550 (N_7550,N_4631,N_5881);
and U7551 (N_7551,N_4861,N_5524);
nor U7552 (N_7552,N_5275,N_4707);
nand U7553 (N_7553,N_4083,N_4394);
nor U7554 (N_7554,N_5179,N_5130);
and U7555 (N_7555,N_4928,N_4755);
and U7556 (N_7556,N_5946,N_5447);
and U7557 (N_7557,N_4167,N_4872);
and U7558 (N_7558,N_4349,N_5712);
and U7559 (N_7559,N_5756,N_4507);
and U7560 (N_7560,N_4766,N_5396);
nor U7561 (N_7561,N_4206,N_5573);
nand U7562 (N_7562,N_4747,N_5349);
nand U7563 (N_7563,N_5429,N_5249);
or U7564 (N_7564,N_5936,N_4803);
and U7565 (N_7565,N_4713,N_4181);
nand U7566 (N_7566,N_4528,N_4312);
and U7567 (N_7567,N_5083,N_4654);
and U7568 (N_7568,N_4010,N_5692);
and U7569 (N_7569,N_5465,N_4518);
nand U7570 (N_7570,N_4736,N_5503);
or U7571 (N_7571,N_4990,N_5563);
and U7572 (N_7572,N_4102,N_5053);
nor U7573 (N_7573,N_5355,N_5991);
and U7574 (N_7574,N_5266,N_5352);
or U7575 (N_7575,N_5612,N_5868);
and U7576 (N_7576,N_5857,N_4010);
nand U7577 (N_7577,N_4498,N_5924);
and U7578 (N_7578,N_4853,N_4542);
or U7579 (N_7579,N_5016,N_5293);
nor U7580 (N_7580,N_4754,N_4755);
or U7581 (N_7581,N_4162,N_4831);
nor U7582 (N_7582,N_4140,N_5847);
and U7583 (N_7583,N_5576,N_4144);
nor U7584 (N_7584,N_5725,N_4889);
or U7585 (N_7585,N_4032,N_4552);
nand U7586 (N_7586,N_5373,N_5588);
nor U7587 (N_7587,N_5841,N_4435);
nand U7588 (N_7588,N_4624,N_5159);
or U7589 (N_7589,N_4414,N_4883);
or U7590 (N_7590,N_5107,N_5989);
nand U7591 (N_7591,N_5125,N_5842);
or U7592 (N_7592,N_5842,N_5932);
and U7593 (N_7593,N_4391,N_4325);
nor U7594 (N_7594,N_4727,N_5002);
or U7595 (N_7595,N_4969,N_4948);
nor U7596 (N_7596,N_4110,N_4748);
or U7597 (N_7597,N_4378,N_4904);
nor U7598 (N_7598,N_5681,N_5502);
and U7599 (N_7599,N_5799,N_4184);
and U7600 (N_7600,N_4940,N_4164);
nor U7601 (N_7601,N_4123,N_5925);
or U7602 (N_7602,N_5049,N_4479);
nand U7603 (N_7603,N_4933,N_4042);
and U7604 (N_7604,N_5602,N_5525);
or U7605 (N_7605,N_4941,N_4745);
nor U7606 (N_7606,N_5060,N_4072);
nand U7607 (N_7607,N_5099,N_4125);
nand U7608 (N_7608,N_4460,N_5366);
or U7609 (N_7609,N_4235,N_5221);
nand U7610 (N_7610,N_5768,N_5075);
and U7611 (N_7611,N_5929,N_5740);
or U7612 (N_7612,N_4511,N_5793);
nor U7613 (N_7613,N_4192,N_5811);
nor U7614 (N_7614,N_4463,N_4839);
and U7615 (N_7615,N_4339,N_5964);
nor U7616 (N_7616,N_5874,N_5830);
or U7617 (N_7617,N_4897,N_5812);
and U7618 (N_7618,N_5867,N_4741);
nor U7619 (N_7619,N_4149,N_5458);
and U7620 (N_7620,N_5071,N_4300);
nor U7621 (N_7621,N_4642,N_5278);
nand U7622 (N_7622,N_5571,N_5501);
or U7623 (N_7623,N_4323,N_4737);
and U7624 (N_7624,N_4377,N_5217);
nand U7625 (N_7625,N_5207,N_5662);
and U7626 (N_7626,N_4805,N_5050);
nor U7627 (N_7627,N_5254,N_5023);
nor U7628 (N_7628,N_4745,N_5969);
and U7629 (N_7629,N_4410,N_4430);
or U7630 (N_7630,N_5421,N_4363);
or U7631 (N_7631,N_5185,N_5706);
nand U7632 (N_7632,N_5982,N_4320);
or U7633 (N_7633,N_4977,N_4733);
nor U7634 (N_7634,N_5670,N_5114);
and U7635 (N_7635,N_5642,N_4083);
nand U7636 (N_7636,N_4063,N_5906);
or U7637 (N_7637,N_5325,N_4996);
and U7638 (N_7638,N_5819,N_5527);
nor U7639 (N_7639,N_5894,N_4974);
nor U7640 (N_7640,N_4434,N_5237);
or U7641 (N_7641,N_5167,N_4818);
and U7642 (N_7642,N_4237,N_4794);
nand U7643 (N_7643,N_5706,N_4928);
or U7644 (N_7644,N_4871,N_5086);
and U7645 (N_7645,N_4352,N_4299);
and U7646 (N_7646,N_4875,N_5463);
or U7647 (N_7647,N_4998,N_4095);
and U7648 (N_7648,N_4576,N_4142);
nor U7649 (N_7649,N_4832,N_4990);
or U7650 (N_7650,N_5477,N_4568);
nand U7651 (N_7651,N_5265,N_4738);
and U7652 (N_7652,N_5812,N_4292);
or U7653 (N_7653,N_4993,N_5944);
nor U7654 (N_7654,N_4834,N_4152);
nand U7655 (N_7655,N_5924,N_5058);
nor U7656 (N_7656,N_5454,N_4041);
nand U7657 (N_7657,N_4746,N_5728);
or U7658 (N_7658,N_4558,N_5045);
nand U7659 (N_7659,N_5776,N_4013);
xnor U7660 (N_7660,N_4613,N_4038);
and U7661 (N_7661,N_4001,N_4572);
nor U7662 (N_7662,N_5055,N_5222);
and U7663 (N_7663,N_4930,N_5559);
nand U7664 (N_7664,N_5088,N_5282);
or U7665 (N_7665,N_5565,N_5073);
nand U7666 (N_7666,N_4075,N_5037);
or U7667 (N_7667,N_4599,N_5645);
or U7668 (N_7668,N_5402,N_5715);
nand U7669 (N_7669,N_5873,N_4592);
or U7670 (N_7670,N_4649,N_4764);
or U7671 (N_7671,N_4435,N_4503);
nand U7672 (N_7672,N_4256,N_4351);
and U7673 (N_7673,N_4172,N_5338);
xor U7674 (N_7674,N_4982,N_5494);
or U7675 (N_7675,N_4467,N_5077);
nand U7676 (N_7676,N_4181,N_5953);
nand U7677 (N_7677,N_4819,N_4663);
nand U7678 (N_7678,N_5577,N_4277);
nand U7679 (N_7679,N_4809,N_4723);
or U7680 (N_7680,N_5734,N_4461);
nand U7681 (N_7681,N_5658,N_5035);
or U7682 (N_7682,N_4991,N_4094);
nor U7683 (N_7683,N_4345,N_4975);
nand U7684 (N_7684,N_5890,N_4802);
and U7685 (N_7685,N_4941,N_5168);
nor U7686 (N_7686,N_5099,N_4396);
or U7687 (N_7687,N_4141,N_5041);
nor U7688 (N_7688,N_5390,N_4921);
nor U7689 (N_7689,N_4810,N_4710);
or U7690 (N_7690,N_5507,N_5382);
and U7691 (N_7691,N_5904,N_4207);
nand U7692 (N_7692,N_4172,N_5407);
and U7693 (N_7693,N_4063,N_5538);
nor U7694 (N_7694,N_4678,N_4187);
nor U7695 (N_7695,N_4111,N_5922);
or U7696 (N_7696,N_5516,N_4896);
nand U7697 (N_7697,N_4932,N_4919);
nor U7698 (N_7698,N_5563,N_5694);
or U7699 (N_7699,N_4435,N_5112);
or U7700 (N_7700,N_5216,N_5458);
or U7701 (N_7701,N_4525,N_4570);
and U7702 (N_7702,N_5066,N_4708);
nor U7703 (N_7703,N_5581,N_5084);
or U7704 (N_7704,N_4321,N_4709);
and U7705 (N_7705,N_5767,N_5811);
nand U7706 (N_7706,N_5151,N_4340);
nand U7707 (N_7707,N_5358,N_4151);
and U7708 (N_7708,N_5598,N_4984);
nand U7709 (N_7709,N_5718,N_5627);
nor U7710 (N_7710,N_4262,N_4872);
nor U7711 (N_7711,N_5242,N_4204);
and U7712 (N_7712,N_4512,N_4531);
and U7713 (N_7713,N_4694,N_5808);
nand U7714 (N_7714,N_5605,N_5246);
and U7715 (N_7715,N_5019,N_5388);
or U7716 (N_7716,N_4201,N_5906);
and U7717 (N_7717,N_4922,N_4873);
nand U7718 (N_7718,N_5774,N_5737);
or U7719 (N_7719,N_5332,N_4850);
and U7720 (N_7720,N_4282,N_4962);
nand U7721 (N_7721,N_4917,N_5489);
nand U7722 (N_7722,N_5465,N_4756);
or U7723 (N_7723,N_5567,N_5962);
or U7724 (N_7724,N_4249,N_5064);
nand U7725 (N_7725,N_4363,N_5838);
nand U7726 (N_7726,N_4987,N_5847);
and U7727 (N_7727,N_4266,N_4225);
or U7728 (N_7728,N_5111,N_4606);
nand U7729 (N_7729,N_5063,N_5458);
or U7730 (N_7730,N_5017,N_5889);
nor U7731 (N_7731,N_5370,N_5726);
nand U7732 (N_7732,N_5800,N_4447);
or U7733 (N_7733,N_4998,N_5717);
nor U7734 (N_7734,N_4518,N_4389);
nand U7735 (N_7735,N_4492,N_5960);
and U7736 (N_7736,N_4262,N_4774);
or U7737 (N_7737,N_5154,N_4467);
or U7738 (N_7738,N_4042,N_5314);
nor U7739 (N_7739,N_4803,N_4435);
or U7740 (N_7740,N_4316,N_5816);
and U7741 (N_7741,N_5257,N_4392);
or U7742 (N_7742,N_4510,N_4859);
and U7743 (N_7743,N_4048,N_4676);
or U7744 (N_7744,N_5346,N_5083);
nor U7745 (N_7745,N_4820,N_5506);
and U7746 (N_7746,N_4436,N_5373);
or U7747 (N_7747,N_5790,N_4143);
or U7748 (N_7748,N_4306,N_5785);
nor U7749 (N_7749,N_5455,N_5481);
nor U7750 (N_7750,N_5108,N_4398);
and U7751 (N_7751,N_4898,N_5054);
nand U7752 (N_7752,N_4510,N_4440);
nand U7753 (N_7753,N_5234,N_5038);
nor U7754 (N_7754,N_5262,N_5835);
or U7755 (N_7755,N_4110,N_5334);
and U7756 (N_7756,N_5656,N_5897);
nor U7757 (N_7757,N_5042,N_5737);
and U7758 (N_7758,N_5732,N_5652);
or U7759 (N_7759,N_4153,N_5425);
nand U7760 (N_7760,N_4467,N_5490);
and U7761 (N_7761,N_5784,N_4858);
nand U7762 (N_7762,N_4255,N_5357);
nor U7763 (N_7763,N_4689,N_4735);
nand U7764 (N_7764,N_5993,N_5851);
nor U7765 (N_7765,N_4158,N_4277);
and U7766 (N_7766,N_5185,N_4917);
nor U7767 (N_7767,N_5653,N_4931);
and U7768 (N_7768,N_5490,N_5246);
or U7769 (N_7769,N_4264,N_5361);
nand U7770 (N_7770,N_5821,N_4512);
or U7771 (N_7771,N_4659,N_4090);
nor U7772 (N_7772,N_5666,N_4909);
nor U7773 (N_7773,N_5942,N_5840);
or U7774 (N_7774,N_5462,N_5092);
nand U7775 (N_7775,N_4321,N_4929);
nand U7776 (N_7776,N_5773,N_4897);
and U7777 (N_7777,N_4707,N_5691);
and U7778 (N_7778,N_4798,N_5822);
or U7779 (N_7779,N_5610,N_4889);
nand U7780 (N_7780,N_4868,N_4369);
and U7781 (N_7781,N_4717,N_5929);
nand U7782 (N_7782,N_4448,N_5536);
nand U7783 (N_7783,N_4392,N_4733);
nor U7784 (N_7784,N_4697,N_5954);
and U7785 (N_7785,N_5496,N_5854);
nor U7786 (N_7786,N_5904,N_5362);
or U7787 (N_7787,N_4122,N_4615);
or U7788 (N_7788,N_5544,N_5157);
nor U7789 (N_7789,N_5185,N_5995);
nand U7790 (N_7790,N_5492,N_4283);
xnor U7791 (N_7791,N_4292,N_5205);
and U7792 (N_7792,N_4615,N_4808);
nor U7793 (N_7793,N_4527,N_5222);
or U7794 (N_7794,N_4618,N_4434);
and U7795 (N_7795,N_4692,N_5940);
nand U7796 (N_7796,N_4631,N_4917);
and U7797 (N_7797,N_4452,N_4956);
nand U7798 (N_7798,N_4205,N_5268);
nand U7799 (N_7799,N_4383,N_4641);
and U7800 (N_7800,N_5669,N_4853);
nor U7801 (N_7801,N_5131,N_4023);
nor U7802 (N_7802,N_5835,N_4124);
nor U7803 (N_7803,N_5293,N_4002);
nand U7804 (N_7804,N_4509,N_5178);
nor U7805 (N_7805,N_4109,N_5432);
or U7806 (N_7806,N_5383,N_4967);
nand U7807 (N_7807,N_5068,N_5874);
and U7808 (N_7808,N_4027,N_5844);
xnor U7809 (N_7809,N_4112,N_4237);
or U7810 (N_7810,N_4821,N_5141);
xnor U7811 (N_7811,N_5555,N_5867);
nand U7812 (N_7812,N_4667,N_4179);
and U7813 (N_7813,N_4370,N_4508);
nor U7814 (N_7814,N_5359,N_5203);
nand U7815 (N_7815,N_4233,N_4320);
and U7816 (N_7816,N_4368,N_4651);
and U7817 (N_7817,N_5462,N_4193);
or U7818 (N_7818,N_5623,N_5589);
nand U7819 (N_7819,N_5911,N_4769);
nand U7820 (N_7820,N_5897,N_5811);
nor U7821 (N_7821,N_5941,N_5470);
nor U7822 (N_7822,N_5235,N_5880);
nand U7823 (N_7823,N_4867,N_4657);
and U7824 (N_7824,N_5143,N_5669);
nor U7825 (N_7825,N_5583,N_5771);
nor U7826 (N_7826,N_4798,N_5357);
nand U7827 (N_7827,N_5549,N_5977);
and U7828 (N_7828,N_5302,N_5691);
nor U7829 (N_7829,N_4994,N_5342);
nor U7830 (N_7830,N_4896,N_4501);
and U7831 (N_7831,N_4412,N_4719);
or U7832 (N_7832,N_4105,N_5500);
nor U7833 (N_7833,N_4658,N_4343);
or U7834 (N_7834,N_5855,N_4118);
nand U7835 (N_7835,N_5044,N_5843);
or U7836 (N_7836,N_4337,N_5666);
nand U7837 (N_7837,N_4652,N_4420);
nand U7838 (N_7838,N_5760,N_5019);
nand U7839 (N_7839,N_5459,N_4228);
or U7840 (N_7840,N_5006,N_4869);
nor U7841 (N_7841,N_4370,N_5382);
and U7842 (N_7842,N_4345,N_5447);
and U7843 (N_7843,N_4556,N_5912);
or U7844 (N_7844,N_5499,N_4674);
or U7845 (N_7845,N_4974,N_4244);
and U7846 (N_7846,N_4336,N_4454);
or U7847 (N_7847,N_5872,N_4004);
and U7848 (N_7848,N_4474,N_5579);
or U7849 (N_7849,N_5997,N_5027);
or U7850 (N_7850,N_5988,N_5010);
nor U7851 (N_7851,N_4554,N_4540);
nand U7852 (N_7852,N_5593,N_5196);
and U7853 (N_7853,N_4407,N_5741);
and U7854 (N_7854,N_5645,N_4098);
or U7855 (N_7855,N_5353,N_4756);
nand U7856 (N_7856,N_4431,N_5796);
and U7857 (N_7857,N_5374,N_5055);
nor U7858 (N_7858,N_4220,N_5955);
or U7859 (N_7859,N_5251,N_5722);
nor U7860 (N_7860,N_4932,N_5410);
or U7861 (N_7861,N_5819,N_4035);
nand U7862 (N_7862,N_4876,N_5436);
and U7863 (N_7863,N_5733,N_4821);
nor U7864 (N_7864,N_5071,N_5095);
and U7865 (N_7865,N_5528,N_5973);
nand U7866 (N_7866,N_5675,N_4654);
nor U7867 (N_7867,N_4778,N_4667);
and U7868 (N_7868,N_4688,N_4147);
or U7869 (N_7869,N_4017,N_5260);
nand U7870 (N_7870,N_4961,N_5544);
and U7871 (N_7871,N_5829,N_4587);
nor U7872 (N_7872,N_5156,N_4713);
and U7873 (N_7873,N_5410,N_5352);
nand U7874 (N_7874,N_4629,N_5358);
nand U7875 (N_7875,N_4705,N_5144);
or U7876 (N_7876,N_5863,N_5710);
and U7877 (N_7877,N_5542,N_4481);
and U7878 (N_7878,N_5406,N_5571);
and U7879 (N_7879,N_4225,N_5285);
nand U7880 (N_7880,N_5071,N_4121);
or U7881 (N_7881,N_5666,N_5891);
or U7882 (N_7882,N_5071,N_4021);
and U7883 (N_7883,N_4551,N_5241);
or U7884 (N_7884,N_5243,N_5358);
or U7885 (N_7885,N_4608,N_4213);
and U7886 (N_7886,N_4445,N_5247);
or U7887 (N_7887,N_4583,N_4208);
nor U7888 (N_7888,N_4445,N_4799);
and U7889 (N_7889,N_5921,N_5395);
and U7890 (N_7890,N_4939,N_4337);
or U7891 (N_7891,N_5199,N_5756);
nor U7892 (N_7892,N_5260,N_4410);
and U7893 (N_7893,N_4312,N_4949);
nand U7894 (N_7894,N_4999,N_5278);
nor U7895 (N_7895,N_5828,N_5621);
nand U7896 (N_7896,N_5090,N_4460);
nand U7897 (N_7897,N_4464,N_4660);
nor U7898 (N_7898,N_5029,N_5463);
xnor U7899 (N_7899,N_5435,N_4385);
nand U7900 (N_7900,N_5431,N_4584);
nand U7901 (N_7901,N_4018,N_5282);
nand U7902 (N_7902,N_4518,N_5720);
and U7903 (N_7903,N_5074,N_5756);
and U7904 (N_7904,N_4342,N_4347);
or U7905 (N_7905,N_5498,N_4165);
and U7906 (N_7906,N_5766,N_5877);
and U7907 (N_7907,N_5164,N_4067);
and U7908 (N_7908,N_4176,N_5863);
and U7909 (N_7909,N_5679,N_4982);
nor U7910 (N_7910,N_5700,N_5016);
nor U7911 (N_7911,N_5843,N_5057);
or U7912 (N_7912,N_5307,N_5660);
nand U7913 (N_7913,N_5799,N_4111);
nor U7914 (N_7914,N_4085,N_4476);
or U7915 (N_7915,N_4299,N_5871);
nand U7916 (N_7916,N_4731,N_4906);
or U7917 (N_7917,N_5536,N_4332);
or U7918 (N_7918,N_5326,N_5248);
nand U7919 (N_7919,N_4582,N_4533);
nor U7920 (N_7920,N_5771,N_5813);
nor U7921 (N_7921,N_5098,N_5555);
nand U7922 (N_7922,N_5161,N_4423);
nor U7923 (N_7923,N_5682,N_5653);
nor U7924 (N_7924,N_5840,N_5447);
nor U7925 (N_7925,N_5164,N_5900);
nand U7926 (N_7926,N_5030,N_4583);
nor U7927 (N_7927,N_4138,N_4498);
and U7928 (N_7928,N_5790,N_4911);
and U7929 (N_7929,N_4578,N_5987);
nor U7930 (N_7930,N_5823,N_4711);
and U7931 (N_7931,N_5251,N_4195);
nand U7932 (N_7932,N_5366,N_5764);
nand U7933 (N_7933,N_4000,N_4088);
nor U7934 (N_7934,N_4023,N_5588);
nor U7935 (N_7935,N_4381,N_5505);
and U7936 (N_7936,N_4743,N_5944);
and U7937 (N_7937,N_5372,N_5882);
or U7938 (N_7938,N_4940,N_4727);
nand U7939 (N_7939,N_4240,N_4524);
and U7940 (N_7940,N_5298,N_4870);
or U7941 (N_7941,N_5298,N_5610);
and U7942 (N_7942,N_5925,N_4872);
or U7943 (N_7943,N_4699,N_4370);
and U7944 (N_7944,N_4429,N_4688);
and U7945 (N_7945,N_4309,N_4405);
or U7946 (N_7946,N_5753,N_4622);
or U7947 (N_7947,N_4628,N_5031);
and U7948 (N_7948,N_5083,N_5093);
nor U7949 (N_7949,N_5981,N_5247);
or U7950 (N_7950,N_4200,N_5858);
nor U7951 (N_7951,N_4106,N_4525);
nor U7952 (N_7952,N_5142,N_4181);
nor U7953 (N_7953,N_4466,N_5507);
nand U7954 (N_7954,N_5208,N_4401);
nand U7955 (N_7955,N_5433,N_4571);
or U7956 (N_7956,N_5341,N_4050);
or U7957 (N_7957,N_5839,N_5968);
nor U7958 (N_7958,N_4999,N_5068);
and U7959 (N_7959,N_4480,N_5164);
or U7960 (N_7960,N_4263,N_4993);
and U7961 (N_7961,N_4020,N_4448);
or U7962 (N_7962,N_4477,N_5045);
and U7963 (N_7963,N_4630,N_4413);
or U7964 (N_7964,N_5899,N_4592);
and U7965 (N_7965,N_4226,N_4135);
or U7966 (N_7966,N_4168,N_5621);
nor U7967 (N_7967,N_4248,N_5745);
xor U7968 (N_7968,N_4828,N_5931);
nand U7969 (N_7969,N_5291,N_5392);
and U7970 (N_7970,N_4046,N_5625);
or U7971 (N_7971,N_5132,N_5020);
nand U7972 (N_7972,N_5652,N_4571);
and U7973 (N_7973,N_5994,N_5704);
or U7974 (N_7974,N_5646,N_5902);
nor U7975 (N_7975,N_4918,N_5437);
and U7976 (N_7976,N_4394,N_5618);
nor U7977 (N_7977,N_5564,N_4448);
nor U7978 (N_7978,N_5079,N_5757);
and U7979 (N_7979,N_5152,N_5812);
or U7980 (N_7980,N_5861,N_5407);
or U7981 (N_7981,N_5775,N_5725);
or U7982 (N_7982,N_5261,N_5630);
or U7983 (N_7983,N_5387,N_5695);
nand U7984 (N_7984,N_4886,N_5666);
and U7985 (N_7985,N_4385,N_5982);
nor U7986 (N_7986,N_4149,N_5487);
nand U7987 (N_7987,N_4467,N_4555);
or U7988 (N_7988,N_4351,N_5132);
nor U7989 (N_7989,N_5959,N_4262);
or U7990 (N_7990,N_5542,N_4189);
and U7991 (N_7991,N_5849,N_4508);
and U7992 (N_7992,N_5141,N_4909);
and U7993 (N_7993,N_4005,N_4374);
and U7994 (N_7994,N_5147,N_4625);
nand U7995 (N_7995,N_4357,N_5750);
or U7996 (N_7996,N_5911,N_4075);
nand U7997 (N_7997,N_5400,N_4508);
and U7998 (N_7998,N_5545,N_4038);
and U7999 (N_7999,N_4638,N_4733);
or U8000 (N_8000,N_6827,N_6982);
and U8001 (N_8001,N_6103,N_6857);
nand U8002 (N_8002,N_6483,N_7719);
nor U8003 (N_8003,N_7410,N_7893);
or U8004 (N_8004,N_6184,N_7199);
nand U8005 (N_8005,N_7048,N_7153);
and U8006 (N_8006,N_6219,N_6462);
or U8007 (N_8007,N_6634,N_6583);
or U8008 (N_8008,N_7497,N_6209);
nand U8009 (N_8009,N_6041,N_6809);
and U8010 (N_8010,N_7094,N_6033);
and U8011 (N_8011,N_7328,N_7091);
xor U8012 (N_8012,N_7227,N_7670);
or U8013 (N_8013,N_7815,N_7068);
or U8014 (N_8014,N_7281,N_7134);
or U8015 (N_8015,N_6735,N_6196);
nor U8016 (N_8016,N_6315,N_6265);
and U8017 (N_8017,N_6683,N_6097);
and U8018 (N_8018,N_7812,N_6118);
nor U8019 (N_8019,N_6451,N_7407);
nor U8020 (N_8020,N_7035,N_7138);
nor U8021 (N_8021,N_7832,N_7366);
and U8022 (N_8022,N_7274,N_7646);
nand U8023 (N_8023,N_6765,N_6043);
nand U8024 (N_8024,N_6040,N_6336);
or U8025 (N_8025,N_6333,N_7548);
and U8026 (N_8026,N_6266,N_7962);
or U8027 (N_8027,N_6142,N_6967);
nand U8028 (N_8028,N_7868,N_6183);
and U8029 (N_8029,N_7530,N_6820);
nand U8030 (N_8030,N_7341,N_6477);
nand U8031 (N_8031,N_6295,N_7899);
nor U8032 (N_8032,N_7985,N_6612);
nor U8033 (N_8033,N_7345,N_6995);
or U8034 (N_8034,N_6861,N_6104);
and U8035 (N_8035,N_7904,N_6302);
nand U8036 (N_8036,N_6567,N_6341);
nor U8037 (N_8037,N_7825,N_6706);
nand U8038 (N_8038,N_7042,N_7754);
and U8039 (N_8039,N_7735,N_7808);
nand U8040 (N_8040,N_6461,N_7222);
or U8041 (N_8041,N_6091,N_6494);
nor U8042 (N_8042,N_7803,N_7124);
and U8043 (N_8043,N_7677,N_7461);
and U8044 (N_8044,N_6695,N_6344);
and U8045 (N_8045,N_6850,N_6356);
nor U8046 (N_8046,N_6999,N_6785);
nor U8047 (N_8047,N_6086,N_6030);
or U8048 (N_8048,N_7974,N_6805);
or U8049 (N_8049,N_7306,N_6597);
nor U8050 (N_8050,N_7896,N_7667);
nand U8051 (N_8051,N_7590,N_6883);
and U8052 (N_8052,N_6403,N_7626);
and U8053 (N_8053,N_6394,N_6591);
nand U8054 (N_8054,N_6289,N_7859);
or U8055 (N_8055,N_6371,N_7304);
nor U8056 (N_8056,N_6505,N_6509);
or U8057 (N_8057,N_6784,N_6538);
nor U8058 (N_8058,N_7598,N_7814);
nor U8059 (N_8059,N_7720,N_6121);
or U8060 (N_8060,N_7044,N_6386);
and U8061 (N_8061,N_6675,N_6790);
nand U8062 (N_8062,N_7241,N_6585);
nand U8063 (N_8063,N_7601,N_7908);
nand U8064 (N_8064,N_6176,N_6520);
nor U8065 (N_8065,N_7840,N_6899);
nand U8066 (N_8066,N_6412,N_6698);
or U8067 (N_8067,N_6846,N_7090);
nor U8068 (N_8068,N_7415,N_6124);
or U8069 (N_8069,N_6946,N_6249);
nor U8070 (N_8070,N_7866,N_6681);
or U8071 (N_8071,N_7665,N_7897);
or U8072 (N_8072,N_7378,N_6450);
nand U8073 (N_8073,N_6770,N_7631);
nand U8074 (N_8074,N_6632,N_6164);
and U8075 (N_8075,N_6794,N_6900);
nor U8076 (N_8076,N_6437,N_7639);
nor U8077 (N_8077,N_7755,N_6831);
or U8078 (N_8078,N_6990,N_6867);
nand U8079 (N_8079,N_6918,N_7202);
nand U8080 (N_8080,N_7903,N_7217);
or U8081 (N_8081,N_7823,N_7089);
or U8082 (N_8082,N_6777,N_6324);
nor U8083 (N_8083,N_7266,N_6102);
and U8084 (N_8084,N_7956,N_7718);
or U8085 (N_8085,N_7422,N_7573);
nor U8086 (N_8086,N_7877,N_7184);
nand U8087 (N_8087,N_7085,N_6185);
nand U8088 (N_8088,N_6711,N_6082);
nand U8089 (N_8089,N_7704,N_6724);
nor U8090 (N_8090,N_6364,N_6804);
or U8091 (N_8091,N_6607,N_7248);
nor U8092 (N_8092,N_7234,N_7565);
xnor U8093 (N_8093,N_6460,N_6865);
and U8094 (N_8094,N_7127,N_6816);
nor U8095 (N_8095,N_7151,N_6439);
nand U8096 (N_8096,N_6405,N_6390);
nand U8097 (N_8097,N_6841,N_7492);
nor U8098 (N_8098,N_6814,N_7087);
and U8099 (N_8099,N_6734,N_7982);
and U8100 (N_8100,N_6313,N_7453);
and U8101 (N_8101,N_6913,N_7233);
nand U8102 (N_8102,N_6125,N_6180);
or U8103 (N_8103,N_7917,N_6068);
nand U8104 (N_8104,N_7243,N_7237);
nand U8105 (N_8105,N_6984,N_7137);
or U8106 (N_8106,N_6113,N_6516);
nand U8107 (N_8107,N_6685,N_7999);
nor U8108 (N_8108,N_6912,N_7521);
nand U8109 (N_8109,N_7249,N_7141);
and U8110 (N_8110,N_7181,N_6376);
nand U8111 (N_8111,N_6745,N_7213);
or U8112 (N_8112,N_7796,N_7173);
nor U8113 (N_8113,N_7169,N_6859);
and U8114 (N_8114,N_7988,N_6329);
or U8115 (N_8115,N_7715,N_6940);
or U8116 (N_8116,N_7552,N_6579);
or U8117 (N_8117,N_7933,N_6666);
nand U8118 (N_8118,N_7978,N_6025);
and U8119 (N_8119,N_6062,N_7011);
and U8120 (N_8120,N_7686,N_6463);
and U8121 (N_8121,N_7675,N_6026);
nand U8122 (N_8122,N_7687,N_7270);
nand U8123 (N_8123,N_7480,N_6932);
nand U8124 (N_8124,N_6527,N_7051);
nand U8125 (N_8125,N_6748,N_7142);
nor U8126 (N_8126,N_6481,N_7721);
or U8127 (N_8127,N_6638,N_6264);
or U8128 (N_8128,N_6544,N_7570);
nor U8129 (N_8129,N_7801,N_6070);
nand U8130 (N_8130,N_6349,N_7285);
or U8131 (N_8131,N_7388,N_6098);
or U8132 (N_8132,N_7693,N_7564);
nand U8133 (N_8133,N_6572,N_7852);
nor U8134 (N_8134,N_7516,N_7887);
and U8135 (N_8135,N_7458,N_7156);
nor U8136 (N_8136,N_7658,N_6957);
nand U8137 (N_8137,N_7283,N_6002);
and U8138 (N_8138,N_7728,N_6452);
nand U8139 (N_8139,N_7514,N_7713);
or U8140 (N_8140,N_7621,N_6599);
or U8141 (N_8141,N_7839,N_7501);
nor U8142 (N_8142,N_7219,N_6127);
nand U8143 (N_8143,N_6747,N_7890);
or U8144 (N_8144,N_6280,N_6725);
nor U8145 (N_8145,N_6168,N_6590);
nand U8146 (N_8146,N_7630,N_6253);
nor U8147 (N_8147,N_7171,N_7060);
and U8148 (N_8148,N_7734,N_7950);
and U8149 (N_8149,N_6073,N_6760);
nor U8150 (N_8150,N_6528,N_7945);
nor U8151 (N_8151,N_7330,N_7816);
nor U8152 (N_8152,N_7723,N_7488);
and U8153 (N_8153,N_7977,N_6881);
xor U8154 (N_8154,N_7117,N_7186);
nor U8155 (N_8155,N_6354,N_6948);
nor U8156 (N_8156,N_7533,N_7440);
or U8157 (N_8157,N_7012,N_7253);
and U8158 (N_8158,N_6928,N_6704);
or U8159 (N_8159,N_7707,N_7826);
nand U8160 (N_8160,N_6262,N_7857);
nand U8161 (N_8161,N_7316,N_7298);
or U8162 (N_8162,N_6239,N_7209);
and U8163 (N_8163,N_7053,N_7017);
and U8164 (N_8164,N_7182,N_7470);
or U8165 (N_8165,N_6971,N_6497);
xor U8166 (N_8166,N_6444,N_6521);
or U8167 (N_8167,N_6015,N_6236);
and U8168 (N_8168,N_6663,N_6863);
and U8169 (N_8169,N_7211,N_6949);
nor U8170 (N_8170,N_7037,N_6631);
nor U8171 (N_8171,N_7997,N_6079);
or U8172 (N_8172,N_7196,N_6966);
and U8173 (N_8173,N_6988,N_6830);
and U8174 (N_8174,N_7534,N_6391);
nor U8175 (N_8175,N_6897,N_7640);
nand U8176 (N_8176,N_7535,N_6480);
nor U8177 (N_8177,N_7411,N_7257);
nand U8178 (N_8178,N_7468,N_6347);
nand U8179 (N_8179,N_6231,N_6757);
and U8180 (N_8180,N_7870,N_6301);
nand U8181 (N_8181,N_7150,N_7439);
nor U8182 (N_8182,N_6036,N_6511);
nor U8183 (N_8183,N_6578,N_7313);
or U8184 (N_8184,N_7240,N_7119);
nor U8185 (N_8185,N_7981,N_6189);
nand U8186 (N_8186,N_6862,N_7389);
and U8187 (N_8187,N_6906,N_6868);
and U8188 (N_8188,N_7296,N_7102);
and U8189 (N_8189,N_7420,N_6673);
nor U8190 (N_8190,N_6429,N_6383);
and U8191 (N_8191,N_7891,N_6751);
nor U8192 (N_8192,N_6998,N_6377);
nor U8193 (N_8193,N_6898,N_6992);
nor U8194 (N_8194,N_7619,N_6517);
or U8195 (N_8195,N_6705,N_7522);
nand U8196 (N_8196,N_7479,N_7070);
nor U8197 (N_8197,N_6308,N_7401);
or U8198 (N_8198,N_7082,N_6114);
nand U8199 (N_8199,N_7584,N_6258);
nor U8200 (N_8200,N_6506,N_6615);
or U8201 (N_8201,N_6909,N_7749);
and U8202 (N_8202,N_7702,N_7600);
nand U8203 (N_8203,N_7284,N_6975);
or U8204 (N_8204,N_7710,N_6738);
nor U8205 (N_8205,N_6016,N_6985);
nand U8206 (N_8206,N_7342,N_6434);
nand U8207 (N_8207,N_7529,N_7556);
and U8208 (N_8208,N_6969,N_6187);
nand U8209 (N_8209,N_7784,N_6422);
and U8210 (N_8210,N_7804,N_7643);
nand U8211 (N_8211,N_7863,N_6340);
or U8212 (N_8212,N_7992,N_7135);
nor U8213 (N_8213,N_6569,N_6312);
nand U8214 (N_8214,N_7419,N_6667);
nand U8215 (N_8215,N_6646,N_7783);
nand U8216 (N_8216,N_7673,N_6260);
nor U8217 (N_8217,N_6054,N_6380);
nand U8218 (N_8218,N_7476,N_6174);
or U8219 (N_8219,N_7958,N_7477);
or U8220 (N_8220,N_6335,N_7813);
or U8221 (N_8221,N_6762,N_7758);
or U8222 (N_8222,N_7023,N_6956);
nor U8223 (N_8223,N_7756,N_7436);
or U8224 (N_8224,N_7180,N_6287);
and U8225 (N_8225,N_7560,N_7036);
and U8226 (N_8226,N_7039,N_6535);
nor U8227 (N_8227,N_7286,N_6603);
nor U8228 (N_8228,N_7581,N_6404);
nand U8229 (N_8229,N_6691,N_6492);
or U8230 (N_8230,N_7375,N_7869);
nor U8231 (N_8231,N_7109,N_7391);
nor U8232 (N_8232,N_6692,N_6873);
nor U8233 (N_8233,N_6580,N_6071);
nand U8234 (N_8234,N_7964,N_6786);
and U8235 (N_8235,N_6779,N_7210);
and U8236 (N_8236,N_7294,N_6093);
nor U8237 (N_8237,N_7688,N_6923);
or U8238 (N_8238,N_6367,N_7768);
nor U8239 (N_8239,N_6801,N_6676);
and U8240 (N_8240,N_7778,N_7575);
and U8241 (N_8241,N_7207,N_7267);
nand U8242 (N_8242,N_7319,N_6508);
or U8243 (N_8243,N_7878,N_6826);
nand U8244 (N_8244,N_6717,N_7500);
xnor U8245 (N_8245,N_6927,N_7973);
nor U8246 (N_8246,N_6924,N_7763);
and U8247 (N_8247,N_6241,N_6929);
or U8248 (N_8248,N_7218,N_6144);
nor U8249 (N_8249,N_7464,N_7197);
and U8250 (N_8250,N_7299,N_7446);
nand U8251 (N_8251,N_6112,N_7926);
nor U8252 (N_8252,N_7520,N_6566);
or U8253 (N_8253,N_6227,N_6962);
nor U8254 (N_8254,N_6600,N_6172);
or U8255 (N_8255,N_6080,N_6067);
or U8256 (N_8256,N_6192,N_7177);
or U8257 (N_8257,N_6773,N_7663);
nand U8258 (N_8258,N_7484,N_6024);
nand U8259 (N_8259,N_6272,N_7699);
nor U8260 (N_8260,N_7849,N_6529);
xor U8261 (N_8261,N_7255,N_7885);
and U8262 (N_8262,N_7547,N_7927);
nand U8263 (N_8263,N_6755,N_7510);
nand U8264 (N_8264,N_6010,N_7147);
nor U8265 (N_8265,N_6800,N_7661);
and U8266 (N_8266,N_6935,N_7200);
or U8267 (N_8267,N_6056,N_7189);
or U8268 (N_8268,N_7224,N_7901);
and U8269 (N_8269,N_7146,N_7059);
and U8270 (N_8270,N_6322,N_7503);
and U8271 (N_8271,N_6120,N_7732);
nand U8272 (N_8272,N_6488,N_6854);
and U8273 (N_8273,N_6148,N_7368);
nor U8274 (N_8274,N_6598,N_6042);
or U8275 (N_8275,N_7416,N_7406);
and U8276 (N_8276,N_7627,N_6359);
and U8277 (N_8277,N_6664,N_7385);
and U8278 (N_8278,N_7539,N_6951);
or U8279 (N_8279,N_7174,N_6563);
nand U8280 (N_8280,N_6983,N_6728);
nand U8281 (N_8281,N_7800,N_6440);
and U8282 (N_8282,N_7122,N_7307);
or U8283 (N_8283,N_6244,N_7472);
nor U8284 (N_8284,N_6836,N_7830);
or U8285 (N_8285,N_7429,N_6166);
nor U8286 (N_8286,N_6531,N_6373);
and U8287 (N_8287,N_6332,N_6296);
nor U8288 (N_8288,N_7604,N_7191);
xor U8289 (N_8289,N_6355,N_6338);
nand U8290 (N_8290,N_6298,N_7622);
and U8291 (N_8291,N_6058,N_6059);
nand U8292 (N_8292,N_6891,N_7265);
nand U8293 (N_8293,N_7157,N_6438);
or U8294 (N_8294,N_7989,N_6533);
nor U8295 (N_8295,N_6447,N_6552);
or U8296 (N_8296,N_6525,N_7690);
or U8297 (N_8297,N_7045,N_7324);
nor U8298 (N_8298,N_7773,N_6661);
nand U8299 (N_8299,N_6345,N_7272);
nand U8300 (N_8300,N_7215,N_7326);
or U8301 (N_8301,N_7340,N_6623);
nand U8302 (N_8302,N_6513,N_6742);
nor U8303 (N_8303,N_7448,N_7460);
or U8304 (N_8304,N_6611,N_7442);
nor U8305 (N_8305,N_6872,N_7443);
nand U8306 (N_8306,N_7187,N_7519);
nor U8307 (N_8307,N_6737,N_6173);
and U8308 (N_8308,N_6620,N_7953);
or U8309 (N_8309,N_6602,N_7551);
nand U8310 (N_8310,N_7128,N_6182);
or U8311 (N_8311,N_7225,N_6108);
and U8312 (N_8312,N_7260,N_7072);
nand U8313 (N_8313,N_7591,N_6261);
nor U8314 (N_8314,N_6369,N_7006);
nand U8315 (N_8315,N_6022,N_6549);
or U8316 (N_8316,N_7795,N_6614);
nand U8317 (N_8317,N_6498,N_6225);
nor U8318 (N_8318,N_6604,N_7923);
or U8319 (N_8319,N_6778,N_7140);
nand U8320 (N_8320,N_7594,N_7921);
and U8321 (N_8321,N_7954,N_7349);
or U8322 (N_8322,N_7049,N_7543);
nand U8323 (N_8323,N_7435,N_6574);
or U8324 (N_8324,N_6635,N_6060);
or U8325 (N_8325,N_7876,N_7913);
nand U8326 (N_8326,N_7861,N_7152);
nand U8327 (N_8327,N_6581,N_7325);
and U8328 (N_8328,N_6720,N_7192);
nor U8329 (N_8329,N_6764,N_7684);
nand U8330 (N_8330,N_7025,N_7165);
nand U8331 (N_8331,N_7761,N_7736);
and U8332 (N_8332,N_6671,N_7015);
nor U8333 (N_8333,N_6639,N_7572);
and U8334 (N_8334,N_6378,N_6084);
or U8335 (N_8335,N_7785,N_6910);
nor U8336 (N_8336,N_7792,N_6892);
nand U8337 (N_8337,N_6920,N_7076);
or U8338 (N_8338,N_7979,N_7297);
nor U8339 (N_8339,N_6979,N_7188);
nand U8340 (N_8340,N_7414,N_7542);
nand U8341 (N_8341,N_7636,N_7567);
nand U8342 (N_8342,N_6637,N_6277);
or U8343 (N_8343,N_7312,N_6464);
nor U8344 (N_8344,N_6372,N_7669);
and U8345 (N_8345,N_7772,N_7562);
or U8346 (N_8346,N_7172,N_7555);
nand U8347 (N_8347,N_7456,N_6561);
nor U8348 (N_8348,N_7935,N_7777);
nor U8349 (N_8349,N_7589,N_6213);
nor U8350 (N_8350,N_7771,N_6076);
and U8351 (N_8351,N_6677,N_6876);
nand U8352 (N_8352,N_6672,N_7568);
or U8353 (N_8353,N_6592,N_6353);
or U8354 (N_8354,N_7379,N_6393);
or U8355 (N_8355,N_6901,N_7327);
and U8356 (N_8356,N_6630,N_6601);
nand U8357 (N_8357,N_7088,N_6388);
nor U8358 (N_8358,N_6582,N_6766);
nor U8359 (N_8359,N_6642,N_7960);
or U8360 (N_8360,N_7236,N_6806);
nor U8361 (N_8361,N_6803,N_7620);
and U8362 (N_8362,N_7104,N_6138);
or U8363 (N_8363,N_7659,N_6278);
nand U8364 (N_8364,N_6240,N_7502);
or U8365 (N_8365,N_7027,N_6221);
nand U8366 (N_8366,N_7867,N_7941);
nor U8367 (N_8367,N_6715,N_6247);
and U8368 (N_8368,N_6293,N_7205);
nor U8369 (N_8369,N_6866,N_7229);
nor U8370 (N_8370,N_6472,N_7805);
nand U8371 (N_8371,N_6772,N_7245);
nor U8372 (N_8372,N_6507,N_6206);
and U8373 (N_8373,N_7158,N_6515);
or U8374 (N_8374,N_6981,N_6000);
nand U8375 (N_8375,N_6584,N_6409);
and U8376 (N_8376,N_7466,N_7374);
and U8377 (N_8377,N_6658,N_6852);
and U8378 (N_8378,N_7990,N_7557);
nand U8379 (N_8379,N_7972,N_7279);
or U8380 (N_8380,N_7132,N_7183);
nor U8381 (N_8381,N_7498,N_7100);
and U8382 (N_8382,N_7616,N_6292);
or U8383 (N_8383,N_6191,N_7062);
nand U8384 (N_8384,N_6586,N_6255);
or U8385 (N_8385,N_6467,N_6047);
nor U8386 (N_8386,N_7709,N_6330);
nand U8387 (N_8387,N_7335,N_6001);
nor U8388 (N_8388,N_6743,N_7524);
or U8389 (N_8389,N_7238,N_6943);
and U8390 (N_8390,N_7216,N_7517);
nand U8391 (N_8391,N_7424,N_7308);
nand U8392 (N_8392,N_7175,N_6471);
or U8393 (N_8393,N_6482,N_6092);
and U8394 (N_8394,N_6453,N_7384);
nand U8395 (N_8395,N_7975,N_7204);
or U8396 (N_8396,N_6305,N_7126);
or U8397 (N_8397,N_6660,N_7275);
and U8398 (N_8398,N_7106,N_7649);
nor U8399 (N_8399,N_6311,N_6346);
nand U8400 (N_8400,N_6065,N_6855);
and U8401 (N_8401,N_6808,N_7741);
xnor U8402 (N_8402,N_6726,N_6035);
nor U8403 (N_8403,N_6775,N_7228);
and U8404 (N_8404,N_7421,N_6413);
nand U8405 (N_8405,N_6887,N_6702);
and U8406 (N_8406,N_7277,N_6514);
or U8407 (N_8407,N_7129,N_6466);
and U8408 (N_8408,N_7776,N_6270);
or U8409 (N_8409,N_6942,N_6541);
nand U8410 (N_8410,N_7322,N_6457);
nand U8411 (N_8411,N_6709,N_6276);
and U8412 (N_8412,N_7028,N_6776);
and U8413 (N_8413,N_7775,N_6141);
nor U8414 (N_8414,N_7121,N_6132);
nand U8415 (N_8415,N_7475,N_7418);
or U8416 (N_8416,N_6589,N_7939);
nand U8417 (N_8417,N_6389,N_7774);
nor U8418 (N_8418,N_7782,N_7613);
nand U8419 (N_8419,N_7525,N_7347);
nand U8420 (N_8420,N_7889,N_6848);
nor U8421 (N_8421,N_7676,N_6813);
nor U8422 (N_8422,N_7559,N_7747);
and U8423 (N_8423,N_6254,N_7337);
nand U8424 (N_8424,N_6003,N_6643);
nor U8425 (N_8425,N_6122,N_7008);
or U8426 (N_8426,N_7398,N_7802);
and U8427 (N_8427,N_6303,N_7080);
and U8428 (N_8428,N_6007,N_7817);
and U8429 (N_8429,N_7133,N_6996);
or U8430 (N_8430,N_7862,N_6245);
and U8431 (N_8431,N_7696,N_7714);
and U8432 (N_8432,N_6028,N_7603);
nor U8433 (N_8433,N_7360,N_7751);
or U8434 (N_8434,N_6847,N_6911);
nor U8435 (N_8435,N_7952,N_7580);
nor U8436 (N_8436,N_7392,N_7226);
nor U8437 (N_8437,N_6947,N_6616);
and U8438 (N_8438,N_6163,N_6880);
nor U8439 (N_8439,N_7336,N_7593);
and U8440 (N_8440,N_6526,N_7352);
nor U8441 (N_8441,N_6570,N_7115);
and U8442 (N_8442,N_6414,N_7427);
nand U8443 (N_8443,N_7261,N_6837);
or U8444 (N_8444,N_7163,N_7526);
nor U8445 (N_8445,N_7907,N_6844);
nand U8446 (N_8446,N_6259,N_6432);
nand U8447 (N_8447,N_7381,N_7550);
nor U8448 (N_8448,N_6135,N_6532);
and U8449 (N_8449,N_7592,N_6411);
nor U8450 (N_8450,N_6860,N_6443);
nor U8451 (N_8451,N_6365,N_7746);
nand U8452 (N_8452,N_6459,N_6449);
or U8453 (N_8453,N_7656,N_6139);
nand U8454 (N_8454,N_7668,N_6564);
or U8455 (N_8455,N_6339,N_7577);
or U8456 (N_8456,N_7871,N_6430);
or U8457 (N_8457,N_7097,N_7101);
and U8458 (N_8458,N_7538,N_6716);
and U8459 (N_8459,N_7949,N_7077);
nand U8460 (N_8460,N_6491,N_7996);
and U8461 (N_8461,N_6694,N_6421);
and U8462 (N_8462,N_6986,N_6636);
and U8463 (N_8463,N_6843,N_7789);
nor U8464 (N_8464,N_6562,N_6408);
nor U8465 (N_8465,N_7936,N_7447);
nor U8466 (N_8466,N_6769,N_6649);
nor U8467 (N_8467,N_6690,N_6781);
nand U8468 (N_8468,N_6707,N_6903);
nor U8469 (N_8469,N_6484,N_6399);
nand U8470 (N_8470,N_6496,N_7932);
and U8471 (N_8471,N_6780,N_7489);
or U8472 (N_8472,N_7483,N_6931);
and U8473 (N_8473,N_6559,N_6271);
and U8474 (N_8474,N_7961,N_6633);
or U8475 (N_8475,N_7518,N_6548);
and U8476 (N_8476,N_7162,N_6152);
and U8477 (N_8477,N_6687,N_6342);
nor U8478 (N_8478,N_7144,N_6651);
or U8479 (N_8479,N_6455,N_7623);
or U8480 (N_8480,N_7810,N_7765);
nor U8481 (N_8481,N_6407,N_6571);
and U8482 (N_8482,N_6368,N_6489);
nor U8483 (N_8483,N_7991,N_6415);
or U8484 (N_8484,N_6933,N_7432);
or U8485 (N_8485,N_6214,N_6744);
or U8486 (N_8486,N_6441,N_6997);
or U8487 (N_8487,N_6953,N_6087);
and U8488 (N_8488,N_7781,N_7905);
nand U8489 (N_8489,N_7739,N_6787);
nor U8490 (N_8490,N_7881,N_6096);
nor U8491 (N_8491,N_7321,N_6107);
or U8492 (N_8492,N_7365,N_6655);
and U8493 (N_8493,N_6023,N_6679);
and U8494 (N_8494,N_7331,N_6834);
nand U8495 (N_8495,N_7452,N_6700);
and U8496 (N_8496,N_7499,N_6090);
and U8497 (N_8497,N_6595,N_7361);
or U8498 (N_8498,N_6479,N_7642);
nand U8499 (N_8499,N_6697,N_6137);
nand U8500 (N_8500,N_7541,N_7726);
or U8501 (N_8501,N_6074,N_6886);
or U8502 (N_8502,N_7853,N_6281);
nand U8503 (N_8503,N_7291,N_6251);
or U8504 (N_8504,N_6829,N_6798);
or U8505 (N_8505,N_6678,N_7041);
nand U8506 (N_8506,N_6487,N_7263);
or U8507 (N_8507,N_7288,N_7323);
or U8508 (N_8508,N_6171,N_7681);
or U8509 (N_8509,N_7882,N_6547);
nand U8510 (N_8510,N_6045,N_7959);
nand U8511 (N_8511,N_6878,N_6545);
or U8512 (N_8512,N_6840,N_6952);
nor U8513 (N_8513,N_7318,N_6626);
and U8514 (N_8514,N_7850,N_7029);
or U8515 (N_8515,N_6625,N_7528);
and U8516 (N_8516,N_6851,N_6162);
and U8517 (N_8517,N_7386,N_6004);
or U8518 (N_8518,N_6713,N_7875);
and U8519 (N_8519,N_7356,N_6314);
and U8520 (N_8520,N_7346,N_7478);
nand U8521 (N_8521,N_7372,N_7929);
and U8522 (N_8522,N_6233,N_7026);
nand U8523 (N_8523,N_6674,N_7376);
or U8524 (N_8524,N_7160,N_7301);
nand U8525 (N_8525,N_7358,N_7176);
nand U8526 (N_8526,N_6445,N_7770);
nand U8527 (N_8527,N_7066,N_6228);
nand U8528 (N_8528,N_7915,N_7258);
nand U8529 (N_8529,N_6657,N_6014);
or U8530 (N_8530,N_6869,N_7231);
nor U8531 (N_8531,N_6970,N_6195);
and U8532 (N_8532,N_6613,N_6767);
nor U8533 (N_8533,N_7009,N_6622);
nor U8534 (N_8534,N_6018,N_7024);
or U8535 (N_8535,N_6044,N_6327);
nand U8536 (N_8536,N_6543,N_7295);
or U8537 (N_8537,N_7983,N_6431);
or U8538 (N_8538,N_7683,N_6011);
nor U8539 (N_8539,N_7485,N_6286);
nand U8540 (N_8540,N_6147,N_6894);
xor U8541 (N_8541,N_6055,N_6199);
nand U8542 (N_8542,N_6750,N_7055);
nor U8543 (N_8543,N_6316,N_7052);
and U8544 (N_8544,N_6210,N_7395);
nor U8545 (N_8545,N_6807,N_7835);
nand U8546 (N_8546,N_7067,N_6617);
nand U8547 (N_8547,N_6237,N_6387);
nor U8548 (N_8548,N_6131,N_6754);
and U8549 (N_8549,N_7431,N_7198);
nand U8550 (N_8550,N_6088,N_6782);
nand U8551 (N_8551,N_6424,N_7113);
or U8552 (N_8552,N_6156,N_6627);
or U8553 (N_8553,N_6536,N_6968);
and U8554 (N_8554,N_7493,N_7947);
nor U8555 (N_8555,N_6588,N_6426);
and U8556 (N_8556,N_7595,N_6619);
or U8557 (N_8557,N_6032,N_7969);
and U8558 (N_8558,N_7164,N_6057);
nand U8559 (N_8559,N_7762,N_6178);
and U8560 (N_8560,N_6401,N_6337);
nor U8561 (N_8561,N_6419,N_7021);
nand U8562 (N_8562,N_7075,N_6965);
nand U8563 (N_8563,N_6703,N_6177);
or U8564 (N_8564,N_7367,N_7433);
nand U8565 (N_8565,N_7383,N_6606);
nor U8566 (N_8566,N_7664,N_7161);
nor U8567 (N_8567,N_6896,N_6160);
nand U8568 (N_8568,N_7032,N_6652);
or U8569 (N_8569,N_7558,N_7845);
and U8570 (N_8570,N_6650,N_6500);
and U8571 (N_8571,N_7531,N_7629);
nand U8572 (N_8572,N_6406,N_7806);
nor U8573 (N_8573,N_7856,N_6291);
or U8574 (N_8574,N_7610,N_6885);
nand U8575 (N_8575,N_7725,N_6038);
or U8576 (N_8576,N_6963,N_6167);
nor U8577 (N_8577,N_6366,N_6628);
and U8578 (N_8578,N_7239,N_7706);
nand U8579 (N_8579,N_7079,N_6741);
nor U8580 (N_8580,N_6425,N_6306);
nor U8581 (N_8581,N_6882,N_6143);
or U8582 (N_8582,N_6476,N_6609);
nor U8583 (N_8583,N_6117,N_7214);
nor U8584 (N_8584,N_7752,N_7976);
or U8585 (N_8585,N_7858,N_7482);
and U8586 (N_8586,N_6550,N_6540);
and U8587 (N_8587,N_6972,N_7865);
nor U8588 (N_8588,N_7571,N_6656);
nor U8589 (N_8589,N_7597,N_6384);
nand U8590 (N_8590,N_7393,N_6012);
and U8591 (N_8591,N_7574,N_6048);
nor U8592 (N_8592,N_6008,N_7689);
or U8593 (N_8593,N_6274,N_6051);
nor U8594 (N_8594,N_7838,N_7276);
nor U8595 (N_8595,N_7438,N_7244);
nor U8596 (N_8596,N_6179,N_6126);
and U8597 (N_8597,N_7018,N_6468);
and U8598 (N_8598,N_7278,N_7167);
nand U8599 (N_8599,N_6853,N_7900);
nor U8600 (N_8600,N_6212,N_7114);
and U8601 (N_8601,N_7148,N_6761);
nand U8602 (N_8602,N_6832,N_7993);
nand U8603 (N_8603,N_6502,N_6864);
nand U8604 (N_8604,N_6792,N_6157);
or U8605 (N_8605,N_6688,N_7201);
or U8606 (N_8606,N_6175,N_6215);
nand U8607 (N_8607,N_6158,N_6037);
or U8608 (N_8608,N_7095,N_6170);
nor U8609 (N_8609,N_7001,N_7057);
nand U8610 (N_8610,N_7451,N_7505);
and U8611 (N_8611,N_6993,N_6653);
or U8612 (N_8612,N_6458,N_7348);
and U8613 (N_8613,N_6534,N_6427);
and U8614 (N_8614,N_7767,N_7944);
nand U8615 (N_8615,N_6629,N_6109);
and U8616 (N_8616,N_6708,N_7578);
nand U8617 (N_8617,N_7963,N_7256);
nor U8618 (N_8618,N_7481,N_6197);
nand U8619 (N_8619,N_7824,N_7462);
or U8620 (N_8620,N_7364,N_6594);
nand U8621 (N_8621,N_6146,N_6955);
or U8622 (N_8622,N_7019,N_7491);
nand U8623 (N_8623,N_6930,N_6052);
nor U8624 (N_8624,N_7911,N_7987);
and U8625 (N_8625,N_6129,N_7705);
and U8626 (N_8626,N_6504,N_7096);
nor U8627 (N_8627,N_6299,N_7682);
nor U8628 (N_8628,N_7957,N_7537);
or U8629 (N_8629,N_7628,N_6351);
nand U8630 (N_8630,N_6648,N_7292);
nand U8631 (N_8631,N_7282,N_7110);
nor U8632 (N_8632,N_7251,N_6478);
and U8633 (N_8633,N_7980,N_7811);
nor U8634 (N_8634,N_6939,N_7879);
nand U8635 (N_8635,N_6907,N_7145);
or U8636 (N_8636,N_7428,N_6269);
nor U8637 (N_8637,N_7408,N_6465);
nand U8638 (N_8638,N_7221,N_6283);
nor U8639 (N_8639,N_6290,N_6682);
nand U8640 (N_8640,N_6925,N_6696);
or U8641 (N_8641,N_6624,N_6753);
or U8642 (N_8642,N_7193,N_6902);
or U8643 (N_8643,N_7844,N_7430);
nand U8644 (N_8644,N_7512,N_7232);
and U8645 (N_8645,N_6811,N_7179);
nand U8646 (N_8646,N_7847,N_7264);
nand U8647 (N_8647,N_7178,N_7599);
or U8648 (N_8648,N_7846,N_7054);
or U8649 (N_8649,N_7515,N_7463);
and U8650 (N_8650,N_7740,N_7737);
nand U8651 (N_8651,N_6774,N_7799);
nor U8652 (N_8652,N_6151,N_6818);
and U8653 (N_8653,N_7925,N_7851);
and U8654 (N_8654,N_7553,N_7536);
or U8655 (N_8655,N_7273,N_6250);
nand U8656 (N_8656,N_6331,N_6207);
or U8657 (N_8657,N_7841,N_6530);
and U8658 (N_8658,N_7371,N_7797);
nor U8659 (N_8659,N_7338,N_6285);
and U8660 (N_8660,N_6822,N_6081);
or U8661 (N_8661,N_6116,N_7078);
nand U8662 (N_8662,N_7250,N_7038);
or U8663 (N_8663,N_6294,N_7827);
and U8664 (N_8664,N_7449,N_7563);
and U8665 (N_8665,N_7654,N_7190);
xnor U8666 (N_8666,N_7780,N_7596);
nor U8667 (N_8667,N_7143,N_7387);
nor U8668 (N_8668,N_7120,N_6684);
nand U8669 (N_8669,N_6326,N_7678);
nor U8670 (N_8670,N_6130,N_6795);
nand U8671 (N_8671,N_7854,N_7764);
nor U8672 (N_8672,N_7016,N_6190);
and U8673 (N_8673,N_6323,N_7587);
or U8674 (N_8674,N_7948,N_6433);
and U8675 (N_8675,N_6789,N_6436);
and U8676 (N_8676,N_7828,N_6382);
and U8677 (N_8677,N_7005,N_7672);
or U8678 (N_8678,N_7602,N_6558);
nand U8679 (N_8679,N_7833,N_7509);
nand U8680 (N_8680,N_6224,N_7745);
and U8681 (N_8681,N_7942,N_6557);
or U8682 (N_8682,N_7195,N_7864);
nand U8683 (N_8683,N_7898,N_6686);
nor U8684 (N_8684,N_7302,N_7561);
nor U8685 (N_8685,N_6473,N_7047);
and U8686 (N_8686,N_7373,N_7081);
or U8687 (N_8687,N_6799,N_6934);
nand U8688 (N_8688,N_7159,N_7695);
nor U8689 (N_8689,N_6680,N_6669);
nand U8690 (N_8690,N_6154,N_6729);
nand U8691 (N_8691,N_6575,N_7607);
nor U8692 (N_8692,N_7545,N_7787);
nand U8693 (N_8693,N_6659,N_6960);
or U8694 (N_8694,N_6718,N_6300);
or U8695 (N_8695,N_6101,N_7698);
and U8696 (N_8696,N_6689,N_6304);
nand U8697 (N_8697,N_7652,N_6325);
nand U8698 (N_8698,N_7994,N_7455);
and U8699 (N_8699,N_7403,N_7662);
nor U8700 (N_8700,N_6363,N_6397);
and U8701 (N_8701,N_6134,N_7657);
and U8702 (N_8702,N_6608,N_6512);
nand U8703 (N_8703,N_7166,N_7708);
and U8704 (N_8704,N_6095,N_7305);
nor U8705 (N_8705,N_7362,N_7700);
or U8706 (N_8706,N_7063,N_7605);
or U8707 (N_8707,N_6736,N_7426);
and U8708 (N_8708,N_7396,N_7909);
nand U8709 (N_8709,N_7744,N_6788);
nor U8710 (N_8710,N_7354,N_7750);
and U8711 (N_8711,N_7400,N_7504);
or U8712 (N_8712,N_7691,N_7692);
and U8713 (N_8713,N_6739,N_7004);
nand U8714 (N_8714,N_6020,N_7742);
and U8715 (N_8715,N_7086,N_7540);
nor U8716 (N_8716,N_7970,N_6937);
nor U8717 (N_8717,N_7259,N_7660);
nor U8718 (N_8718,N_6499,N_6423);
or U8719 (N_8719,N_7280,N_7680);
nand U8720 (N_8720,N_7471,N_6596);
nor U8721 (N_8721,N_6111,N_6922);
and U8722 (N_8722,N_6049,N_6890);
or U8723 (N_8723,N_6796,N_7608);
nor U8724 (N_8724,N_7922,N_6699);
or U8725 (N_8725,N_6398,N_7230);
nand U8726 (N_8726,N_7809,N_7916);
or U8727 (N_8727,N_7269,N_7819);
nand U8728 (N_8728,N_6542,N_6381);
and U8729 (N_8729,N_6064,N_7582);
and U8730 (N_8730,N_7511,N_7467);
nor U8731 (N_8731,N_7829,N_7252);
or U8732 (N_8732,N_7311,N_7353);
nor U8733 (N_8733,N_7290,N_6522);
nor U8734 (N_8734,N_7000,N_7494);
nand U8735 (N_8735,N_6916,N_7412);
nor U8736 (N_8736,N_7423,N_7874);
nor U8737 (N_8737,N_7506,N_6230);
nor U8738 (N_8738,N_6223,N_7583);
nand U8739 (N_8739,N_6587,N_6740);
nor U8740 (N_8740,N_7951,N_6470);
or U8741 (N_8741,N_7995,N_6297);
nor U8742 (N_8742,N_6273,N_6879);
nor U8743 (N_8743,N_6723,N_6085);
nor U8744 (N_8744,N_6229,N_6870);
or U8745 (N_8745,N_6208,N_7549);
xnor U8746 (N_8746,N_7390,N_6964);
nor U8747 (N_8747,N_6746,N_6503);
nor U8748 (N_8748,N_6919,N_6936);
nand U8749 (N_8749,N_7554,N_7003);
and U8750 (N_8750,N_7434,N_6410);
nor U8751 (N_8751,N_7108,N_7786);
or U8752 (N_8752,N_7370,N_6029);
and U8753 (N_8753,N_7585,N_7920);
nand U8754 (N_8754,N_6537,N_7727);
and U8755 (N_8755,N_6670,N_6730);
and U8756 (N_8756,N_6759,N_7287);
nor U8757 (N_8757,N_7892,N_7724);
nand U8758 (N_8758,N_7712,N_6825);
nor U8759 (N_8759,N_6017,N_6454);
nand U8760 (N_8760,N_6647,N_6693);
nand U8761 (N_8761,N_6921,N_6034);
nand U8762 (N_8762,N_6824,N_7711);
nor U8763 (N_8763,N_7655,N_6721);
and U8764 (N_8764,N_7417,N_6733);
and U8765 (N_8765,N_6153,N_6392);
or U8766 (N_8766,N_6418,N_6242);
nand U8767 (N_8767,N_7641,N_6944);
nor U8768 (N_8768,N_7757,N_7030);
nand U8769 (N_8769,N_6379,N_6161);
nand U8770 (N_8770,N_6050,N_6267);
and U8771 (N_8771,N_7617,N_7441);
or U8772 (N_8772,N_6758,N_6288);
nand U8773 (N_8773,N_7355,N_7043);
and U8774 (N_8774,N_6518,N_7943);
or U8775 (N_8775,N_7118,N_6618);
or U8776 (N_8776,N_7332,N_7444);
nor U8777 (N_8777,N_6257,N_7984);
nand U8778 (N_8778,N_6554,N_7930);
nand U8779 (N_8779,N_6875,N_7685);
or U8780 (N_8780,N_6908,N_7399);
nand U8781 (N_8781,N_6605,N_7733);
nand U8782 (N_8782,N_7894,N_7918);
or U8783 (N_8783,N_6812,N_7873);
or U8784 (N_8784,N_6884,N_6063);
and U8785 (N_8785,N_7790,N_7363);
nand U8786 (N_8786,N_7615,N_6094);
and U8787 (N_8787,N_7007,N_7208);
nor U8788 (N_8788,N_6845,N_7940);
and U8789 (N_8789,N_7834,N_6155);
and U8790 (N_8790,N_7624,N_7377);
and U8791 (N_8791,N_7872,N_7527);
nor U8792 (N_8792,N_7459,N_7820);
nand U8793 (N_8793,N_7343,N_7474);
and U8794 (N_8794,N_6645,N_7022);
nor U8795 (N_8795,N_6078,N_6256);
or U8796 (N_8796,N_7638,N_7588);
nand U8797 (N_8797,N_7344,N_6435);
or U8798 (N_8798,N_6714,N_6402);
or U8799 (N_8799,N_6756,N_7883);
nor U8800 (N_8800,N_7469,N_7569);
and U8801 (N_8801,N_6895,N_6334);
nand U8802 (N_8802,N_7650,N_7968);
or U8803 (N_8803,N_7753,N_6823);
or U8804 (N_8804,N_6905,N_6752);
nor U8805 (N_8805,N_6317,N_6976);
and U8806 (N_8806,N_7694,N_7380);
or U8807 (N_8807,N_6819,N_6069);
nand U8808 (N_8808,N_7880,N_7056);
and U8809 (N_8809,N_6701,N_7955);
nand U8810 (N_8810,N_7637,N_6926);
nor U8811 (N_8811,N_6053,N_6849);
nand U8812 (N_8812,N_7566,N_6089);
and U8813 (N_8813,N_7651,N_7223);
and U8814 (N_8814,N_7125,N_7050);
or U8815 (N_8815,N_6874,N_7271);
and U8816 (N_8816,N_7154,N_6428);
and U8817 (N_8817,N_7611,N_6490);
and U8818 (N_8818,N_6802,N_6204);
nor U8819 (N_8819,N_6099,N_6123);
and U8820 (N_8820,N_7092,N_6551);
and U8821 (N_8821,N_6959,N_7033);
nand U8822 (N_8822,N_6193,N_6565);
and U8823 (N_8823,N_7473,N_6348);
or U8824 (N_8824,N_7112,N_7634);
nor U8825 (N_8825,N_7058,N_7579);
and U8826 (N_8826,N_6889,N_7350);
nand U8827 (N_8827,N_7437,N_6201);
or U8828 (N_8828,N_6222,N_6553);
and U8829 (N_8829,N_6105,N_6320);
nand U8830 (N_8830,N_6654,N_6560);
nand U8831 (N_8831,N_7369,N_6954);
and U8832 (N_8832,N_6573,N_6220);
nand U8833 (N_8833,N_7487,N_6362);
and U8834 (N_8834,N_6248,N_7532);
nor U8835 (N_8835,N_6119,N_7716);
or U8836 (N_8836,N_6279,N_6978);
or U8837 (N_8837,N_7648,N_7098);
nand U8838 (N_8838,N_7220,N_6246);
nor U8839 (N_8839,N_7938,N_6039);
or U8840 (N_8840,N_7206,N_7357);
or U8841 (N_8841,N_7262,N_7409);
nand U8842 (N_8842,N_7674,N_7203);
and U8843 (N_8843,N_7759,N_7821);
nand U8844 (N_8844,N_6858,N_6791);
and U8845 (N_8845,N_7103,N_7303);
and U8846 (N_8846,N_7644,N_6833);
nor U8847 (N_8847,N_6749,N_6310);
nor U8848 (N_8848,N_6448,N_7099);
nor U8849 (N_8849,N_7612,N_7465);
or U8850 (N_8850,N_7717,N_7779);
or U8851 (N_8851,N_7314,N_7807);
nand U8852 (N_8852,N_6610,N_6486);
nand U8853 (N_8853,N_6485,N_6350);
nor U8854 (N_8854,N_6941,N_6357);
and U8855 (N_8855,N_7793,N_7065);
nor U8856 (N_8856,N_7123,N_6360);
nor U8857 (N_8857,N_6165,N_7544);
nand U8858 (N_8858,N_6077,N_6731);
and U8859 (N_8859,N_7046,N_7425);
nor U8860 (N_8860,N_7083,N_7130);
or U8861 (N_8861,N_6027,N_6842);
nand U8862 (N_8862,N_6835,N_6046);
nor U8863 (N_8863,N_6817,N_6456);
and U8864 (N_8864,N_7334,N_7293);
or U8865 (N_8865,N_7139,N_6732);
nand U8866 (N_8866,N_6719,N_7843);
or U8867 (N_8867,N_7170,N_7986);
or U8868 (N_8868,N_6005,N_6352);
and U8869 (N_8869,N_7906,N_7729);
nand U8870 (N_8870,N_7788,N_7246);
nor U8871 (N_8871,N_6186,N_7647);
or U8872 (N_8872,N_7315,N_6938);
and U8873 (N_8873,N_6263,N_6973);
and U8874 (N_8874,N_6009,N_6523);
nand U8875 (N_8875,N_7625,N_7185);
xor U8876 (N_8876,N_6977,N_6793);
nand U8877 (N_8877,N_6061,N_7309);
nor U8878 (N_8878,N_7855,N_6668);
or U8879 (N_8879,N_6797,N_6205);
nand U8880 (N_8880,N_6385,N_7212);
and U8881 (N_8881,N_6361,N_6621);
and U8882 (N_8882,N_6577,N_6961);
nor U8883 (N_8883,N_7576,N_6031);
and U8884 (N_8884,N_6915,N_7168);
and U8885 (N_8885,N_7450,N_7766);
or U8886 (N_8886,N_6319,N_7666);
nor U8887 (N_8887,N_7928,N_6169);
nand U8888 (N_8888,N_7822,N_7194);
or U8889 (N_8889,N_7965,N_7946);
nor U8890 (N_8890,N_6128,N_6593);
nor U8891 (N_8891,N_6856,N_6268);
and U8892 (N_8892,N_6358,N_6328);
nor U8893 (N_8893,N_6309,N_7105);
and U8894 (N_8894,N_7842,N_7413);
nor U8895 (N_8895,N_6519,N_7235);
nor U8896 (N_8896,N_7031,N_7798);
and U8897 (N_8897,N_6416,N_6877);
or U8898 (N_8898,N_7074,N_7495);
and U8899 (N_8899,N_7914,N_7760);
nor U8900 (N_8900,N_6469,N_6370);
and U8901 (N_8901,N_7069,N_6275);
or U8902 (N_8902,N_6989,N_6555);
nor U8903 (N_8903,N_7937,N_6149);
and U8904 (N_8904,N_7653,N_6396);
nand U8905 (N_8905,N_7586,N_7402);
nand U8906 (N_8906,N_7919,N_6640);
and U8907 (N_8907,N_7998,N_6202);
and U8908 (N_8908,N_7738,N_7697);
nor U8909 (N_8909,N_6066,N_6644);
nand U8910 (N_8910,N_7912,N_6783);
and U8911 (N_8911,N_6216,N_7339);
nor U8912 (N_8912,N_7486,N_7329);
or U8913 (N_8913,N_7382,N_7404);
or U8914 (N_8914,N_7730,N_6136);
or U8915 (N_8915,N_6318,N_6991);
or U8916 (N_8916,N_6763,N_7116);
or U8917 (N_8917,N_7794,N_6871);
nand U8918 (N_8918,N_7310,N_6474);
and U8919 (N_8919,N_6013,N_6442);
or U8920 (N_8920,N_7242,N_7445);
or U8921 (N_8921,N_6838,N_6100);
and U8922 (N_8922,N_7020,N_6321);
and U8923 (N_8923,N_6106,N_6232);
and U8924 (N_8924,N_6375,N_7254);
or U8925 (N_8925,N_6420,N_7061);
or U8926 (N_8926,N_6282,N_6021);
and U8927 (N_8927,N_7093,N_7010);
nand U8928 (N_8928,N_7333,N_7268);
nor U8929 (N_8929,N_7769,N_6252);
nor U8930 (N_8930,N_6115,N_7722);
nor U8931 (N_8931,N_6495,N_6417);
and U8932 (N_8932,N_7743,N_7836);
nor U8933 (N_8933,N_6211,N_6218);
or U8934 (N_8934,N_6140,N_7397);
nor U8935 (N_8935,N_6501,N_6181);
nand U8936 (N_8936,N_7111,N_6958);
nor U8937 (N_8937,N_7902,N_7457);
nor U8938 (N_8938,N_7895,N_7394);
nand U8939 (N_8939,N_7300,N_7084);
and U8940 (N_8940,N_7837,N_7971);
and U8941 (N_8941,N_7934,N_6641);
nand U8942 (N_8942,N_7633,N_6150);
and U8943 (N_8943,N_6110,N_6235);
and U8944 (N_8944,N_6475,N_7910);
nand U8945 (N_8945,N_7289,N_7073);
nor U8946 (N_8946,N_7034,N_6904);
nor U8947 (N_8947,N_7014,N_7523);
nor U8948 (N_8948,N_6893,N_7791);
nand U8949 (N_8949,N_6839,N_6133);
nor U8950 (N_8950,N_6072,N_7966);
nand U8951 (N_8951,N_6576,N_6395);
and U8952 (N_8952,N_7508,N_7632);
or U8953 (N_8953,N_6710,N_6217);
xor U8954 (N_8954,N_7317,N_6145);
nor U8955 (N_8955,N_6945,N_7931);
nand U8956 (N_8956,N_6284,N_7405);
nand U8957 (N_8957,N_7359,N_7490);
or U8958 (N_8958,N_6888,N_7731);
or U8959 (N_8959,N_6075,N_6243);
and U8960 (N_8960,N_6083,N_6980);
and U8961 (N_8961,N_7860,N_7149);
and U8962 (N_8962,N_7064,N_6768);
nand U8963 (N_8963,N_7703,N_6524);
nor U8964 (N_8964,N_6510,N_7635);
nand U8965 (N_8965,N_7924,N_7606);
or U8966 (N_8966,N_7040,N_7247);
or U8967 (N_8967,N_7131,N_7513);
nand U8968 (N_8968,N_6400,N_6950);
and U8969 (N_8969,N_6188,N_6917);
nor U8970 (N_8970,N_6203,N_6019);
nand U8971 (N_8971,N_6374,N_7320);
nand U8972 (N_8972,N_7671,N_7831);
or U8973 (N_8973,N_7454,N_7679);
nand U8974 (N_8974,N_7848,N_7886);
nand U8975 (N_8975,N_7609,N_6307);
nand U8976 (N_8976,N_7818,N_7748);
nor U8977 (N_8977,N_7618,N_7136);
and U8978 (N_8978,N_6821,N_7507);
nand U8979 (N_8979,N_6539,N_7107);
and U8980 (N_8980,N_6446,N_6006);
or U8981 (N_8981,N_7496,N_6987);
nor U8982 (N_8982,N_6810,N_6712);
nand U8983 (N_8983,N_6194,N_7351);
nand U8984 (N_8984,N_6914,N_7546);
nand U8985 (N_8985,N_6493,N_7013);
and U8986 (N_8986,N_6556,N_6198);
nand U8987 (N_8987,N_6546,N_6200);
or U8988 (N_8988,N_7884,N_6771);
and U8989 (N_8989,N_6974,N_7155);
and U8990 (N_8990,N_6727,N_6815);
and U8991 (N_8991,N_7967,N_7071);
nor U8992 (N_8992,N_6343,N_7614);
nor U8993 (N_8993,N_7701,N_7645);
and U8994 (N_8994,N_6238,N_7888);
nand U8995 (N_8995,N_7002,N_6234);
and U8996 (N_8996,N_6994,N_6722);
and U8997 (N_8997,N_6665,N_6226);
nand U8998 (N_8998,N_6159,N_6568);
nand U8999 (N_8999,N_6828,N_6662);
nand U9000 (N_9000,N_7197,N_7886);
nand U9001 (N_9001,N_6955,N_7623);
nand U9002 (N_9002,N_6569,N_7729);
nand U9003 (N_9003,N_7112,N_7472);
or U9004 (N_9004,N_7785,N_6481);
or U9005 (N_9005,N_6593,N_6781);
xor U9006 (N_9006,N_6199,N_6943);
and U9007 (N_9007,N_6208,N_6396);
nand U9008 (N_9008,N_7321,N_6992);
and U9009 (N_9009,N_6993,N_7195);
nand U9010 (N_9010,N_7062,N_6139);
nor U9011 (N_9011,N_7553,N_7186);
or U9012 (N_9012,N_6034,N_7651);
nand U9013 (N_9013,N_6394,N_7558);
nand U9014 (N_9014,N_6707,N_7089);
nor U9015 (N_9015,N_6438,N_6522);
or U9016 (N_9016,N_7545,N_6155);
xnor U9017 (N_9017,N_6774,N_7674);
or U9018 (N_9018,N_7380,N_7869);
and U9019 (N_9019,N_7770,N_7578);
and U9020 (N_9020,N_6357,N_7775);
nand U9021 (N_9021,N_7313,N_6543);
nor U9022 (N_9022,N_7260,N_7068);
or U9023 (N_9023,N_6780,N_7455);
nand U9024 (N_9024,N_7031,N_7540);
nand U9025 (N_9025,N_6484,N_7809);
or U9026 (N_9026,N_7328,N_7941);
or U9027 (N_9027,N_6317,N_6624);
nand U9028 (N_9028,N_7564,N_6013);
and U9029 (N_9029,N_6418,N_7495);
or U9030 (N_9030,N_7898,N_6897);
or U9031 (N_9031,N_7413,N_6728);
nand U9032 (N_9032,N_6422,N_6721);
nand U9033 (N_9033,N_6751,N_7997);
nor U9034 (N_9034,N_7784,N_7053);
nor U9035 (N_9035,N_6444,N_6566);
or U9036 (N_9036,N_7865,N_7506);
and U9037 (N_9037,N_6952,N_6860);
nand U9038 (N_9038,N_7098,N_7997);
nand U9039 (N_9039,N_7088,N_6060);
nor U9040 (N_9040,N_7053,N_6612);
nor U9041 (N_9041,N_7478,N_7489);
and U9042 (N_9042,N_6841,N_6251);
and U9043 (N_9043,N_7329,N_7141);
and U9044 (N_9044,N_7145,N_7173);
or U9045 (N_9045,N_6249,N_7583);
and U9046 (N_9046,N_7132,N_7770);
nand U9047 (N_9047,N_6237,N_7546);
nor U9048 (N_9048,N_6209,N_6142);
and U9049 (N_9049,N_6893,N_7095);
or U9050 (N_9050,N_7373,N_6322);
or U9051 (N_9051,N_6081,N_7661);
nor U9052 (N_9052,N_7082,N_7308);
nand U9053 (N_9053,N_6087,N_7311);
nand U9054 (N_9054,N_6331,N_6932);
or U9055 (N_9055,N_7958,N_7503);
and U9056 (N_9056,N_6177,N_7823);
nor U9057 (N_9057,N_6161,N_6728);
or U9058 (N_9058,N_6699,N_6607);
or U9059 (N_9059,N_7680,N_7603);
nand U9060 (N_9060,N_7240,N_7039);
nor U9061 (N_9061,N_6778,N_7510);
or U9062 (N_9062,N_7230,N_7832);
and U9063 (N_9063,N_7065,N_7716);
nor U9064 (N_9064,N_6283,N_7395);
nor U9065 (N_9065,N_6930,N_6741);
nor U9066 (N_9066,N_7656,N_6333);
and U9067 (N_9067,N_7818,N_7098);
nand U9068 (N_9068,N_6247,N_6689);
or U9069 (N_9069,N_6281,N_6055);
and U9070 (N_9070,N_6390,N_7893);
or U9071 (N_9071,N_7622,N_6437);
xor U9072 (N_9072,N_7434,N_6456);
nand U9073 (N_9073,N_7966,N_7408);
nand U9074 (N_9074,N_6840,N_7228);
nor U9075 (N_9075,N_6341,N_7847);
nor U9076 (N_9076,N_7233,N_7903);
or U9077 (N_9077,N_7516,N_6780);
nand U9078 (N_9078,N_7705,N_7114);
nor U9079 (N_9079,N_7105,N_6089);
nand U9080 (N_9080,N_7261,N_6893);
or U9081 (N_9081,N_7070,N_6060);
nand U9082 (N_9082,N_7437,N_7498);
or U9083 (N_9083,N_7720,N_7047);
and U9084 (N_9084,N_6042,N_7704);
nand U9085 (N_9085,N_6469,N_7190);
nor U9086 (N_9086,N_6903,N_7558);
nand U9087 (N_9087,N_7617,N_6798);
or U9088 (N_9088,N_7227,N_6982);
nor U9089 (N_9089,N_6353,N_7369);
nand U9090 (N_9090,N_6048,N_6374);
nand U9091 (N_9091,N_6274,N_7243);
or U9092 (N_9092,N_6805,N_7317);
nand U9093 (N_9093,N_6407,N_7855);
and U9094 (N_9094,N_7322,N_7467);
nor U9095 (N_9095,N_6072,N_7183);
nor U9096 (N_9096,N_6635,N_6015);
or U9097 (N_9097,N_7733,N_6755);
nor U9098 (N_9098,N_6819,N_7407);
or U9099 (N_9099,N_7672,N_7074);
and U9100 (N_9100,N_7728,N_6598);
and U9101 (N_9101,N_7334,N_6003);
or U9102 (N_9102,N_7331,N_7349);
and U9103 (N_9103,N_7619,N_6928);
nand U9104 (N_9104,N_6123,N_7426);
or U9105 (N_9105,N_6815,N_7543);
or U9106 (N_9106,N_7470,N_6271);
and U9107 (N_9107,N_6029,N_7998);
nor U9108 (N_9108,N_6090,N_6736);
nor U9109 (N_9109,N_6874,N_6335);
and U9110 (N_9110,N_7973,N_7947);
nand U9111 (N_9111,N_7566,N_6057);
nor U9112 (N_9112,N_7955,N_6564);
and U9113 (N_9113,N_7004,N_7016);
nor U9114 (N_9114,N_6977,N_6444);
nand U9115 (N_9115,N_6880,N_6058);
nor U9116 (N_9116,N_7770,N_6625);
and U9117 (N_9117,N_6864,N_7755);
nand U9118 (N_9118,N_7233,N_7064);
nor U9119 (N_9119,N_6351,N_7107);
nor U9120 (N_9120,N_6283,N_7106);
and U9121 (N_9121,N_6960,N_6724);
nand U9122 (N_9122,N_6723,N_7473);
or U9123 (N_9123,N_7962,N_7414);
nand U9124 (N_9124,N_7032,N_6198);
and U9125 (N_9125,N_7344,N_7045);
nor U9126 (N_9126,N_7094,N_7887);
nor U9127 (N_9127,N_6881,N_6368);
nor U9128 (N_9128,N_7765,N_7365);
and U9129 (N_9129,N_7941,N_6340);
nand U9130 (N_9130,N_7403,N_7539);
nand U9131 (N_9131,N_6310,N_7241);
nor U9132 (N_9132,N_6065,N_7073);
and U9133 (N_9133,N_6700,N_7679);
nor U9134 (N_9134,N_6860,N_6471);
or U9135 (N_9135,N_6262,N_7579);
nand U9136 (N_9136,N_6068,N_6536);
nand U9137 (N_9137,N_7071,N_7864);
or U9138 (N_9138,N_7401,N_7855);
nand U9139 (N_9139,N_7917,N_6857);
nand U9140 (N_9140,N_6190,N_6807);
nand U9141 (N_9141,N_6275,N_7551);
xor U9142 (N_9142,N_6514,N_6552);
nor U9143 (N_9143,N_6761,N_6572);
nand U9144 (N_9144,N_6537,N_6153);
or U9145 (N_9145,N_6287,N_6457);
and U9146 (N_9146,N_7289,N_7221);
nor U9147 (N_9147,N_6536,N_6562);
or U9148 (N_9148,N_7563,N_7744);
and U9149 (N_9149,N_7433,N_7333);
or U9150 (N_9150,N_6690,N_6441);
nand U9151 (N_9151,N_7086,N_7894);
or U9152 (N_9152,N_6614,N_6147);
and U9153 (N_9153,N_7251,N_6857);
nor U9154 (N_9154,N_6001,N_7545);
and U9155 (N_9155,N_7368,N_6250);
and U9156 (N_9156,N_6702,N_6753);
nor U9157 (N_9157,N_6718,N_6566);
and U9158 (N_9158,N_7671,N_6295);
or U9159 (N_9159,N_7440,N_7419);
and U9160 (N_9160,N_7514,N_6040);
and U9161 (N_9161,N_6100,N_7456);
nor U9162 (N_9162,N_6977,N_7981);
xnor U9163 (N_9163,N_7239,N_6930);
or U9164 (N_9164,N_7883,N_6928);
or U9165 (N_9165,N_7329,N_7652);
or U9166 (N_9166,N_6832,N_7248);
and U9167 (N_9167,N_7660,N_7379);
or U9168 (N_9168,N_6073,N_6698);
nand U9169 (N_9169,N_6441,N_6592);
nor U9170 (N_9170,N_6323,N_6306);
and U9171 (N_9171,N_6161,N_7219);
or U9172 (N_9172,N_6011,N_7196);
nand U9173 (N_9173,N_7247,N_6742);
or U9174 (N_9174,N_7823,N_7530);
or U9175 (N_9175,N_7709,N_6324);
nand U9176 (N_9176,N_6157,N_6100);
nand U9177 (N_9177,N_7198,N_6623);
nand U9178 (N_9178,N_6378,N_6459);
and U9179 (N_9179,N_6029,N_7960);
and U9180 (N_9180,N_6764,N_6228);
and U9181 (N_9181,N_7987,N_6832);
nor U9182 (N_9182,N_7687,N_6845);
and U9183 (N_9183,N_6103,N_7944);
and U9184 (N_9184,N_7876,N_6071);
or U9185 (N_9185,N_6021,N_7810);
nor U9186 (N_9186,N_6963,N_7336);
nand U9187 (N_9187,N_6803,N_7298);
and U9188 (N_9188,N_6951,N_6414);
and U9189 (N_9189,N_7846,N_7027);
and U9190 (N_9190,N_6478,N_7015);
and U9191 (N_9191,N_6075,N_7220);
nand U9192 (N_9192,N_7201,N_7045);
nand U9193 (N_9193,N_7251,N_7960);
nand U9194 (N_9194,N_6103,N_6513);
nor U9195 (N_9195,N_7368,N_6785);
and U9196 (N_9196,N_6601,N_7888);
nor U9197 (N_9197,N_7123,N_7898);
nor U9198 (N_9198,N_6415,N_7569);
or U9199 (N_9199,N_7962,N_6654);
nor U9200 (N_9200,N_7893,N_6582);
nor U9201 (N_9201,N_6196,N_6162);
nor U9202 (N_9202,N_7877,N_6934);
nor U9203 (N_9203,N_6189,N_7714);
or U9204 (N_9204,N_7871,N_7518);
or U9205 (N_9205,N_7730,N_7831);
or U9206 (N_9206,N_7236,N_7670);
nor U9207 (N_9207,N_7904,N_6735);
or U9208 (N_9208,N_7149,N_7593);
and U9209 (N_9209,N_6552,N_6500);
or U9210 (N_9210,N_7044,N_7684);
nor U9211 (N_9211,N_7704,N_6009);
nor U9212 (N_9212,N_6811,N_7194);
and U9213 (N_9213,N_6440,N_6423);
nand U9214 (N_9214,N_7425,N_6166);
or U9215 (N_9215,N_6604,N_6889);
nor U9216 (N_9216,N_6711,N_7333);
and U9217 (N_9217,N_7575,N_6780);
or U9218 (N_9218,N_6603,N_7400);
nor U9219 (N_9219,N_7072,N_7682);
and U9220 (N_9220,N_7009,N_7275);
or U9221 (N_9221,N_7735,N_7145);
nor U9222 (N_9222,N_6912,N_6815);
or U9223 (N_9223,N_7872,N_6158);
nor U9224 (N_9224,N_7591,N_7383);
nand U9225 (N_9225,N_7032,N_7556);
nor U9226 (N_9226,N_7599,N_7867);
nor U9227 (N_9227,N_6774,N_7053);
nand U9228 (N_9228,N_7819,N_6873);
nand U9229 (N_9229,N_6948,N_6676);
nand U9230 (N_9230,N_6247,N_6163);
nand U9231 (N_9231,N_7154,N_7866);
xor U9232 (N_9232,N_6177,N_6794);
or U9233 (N_9233,N_6058,N_7041);
or U9234 (N_9234,N_6793,N_7804);
or U9235 (N_9235,N_6734,N_7555);
nor U9236 (N_9236,N_6798,N_6177);
nand U9237 (N_9237,N_7529,N_7316);
or U9238 (N_9238,N_6187,N_7443);
nand U9239 (N_9239,N_7876,N_6785);
and U9240 (N_9240,N_7392,N_6905);
nand U9241 (N_9241,N_7278,N_6315);
nor U9242 (N_9242,N_6172,N_6471);
and U9243 (N_9243,N_7699,N_7830);
and U9244 (N_9244,N_6769,N_6830);
nor U9245 (N_9245,N_6698,N_7512);
or U9246 (N_9246,N_7215,N_7366);
nor U9247 (N_9247,N_6185,N_7438);
or U9248 (N_9248,N_7515,N_6147);
and U9249 (N_9249,N_7542,N_6834);
or U9250 (N_9250,N_7865,N_7768);
or U9251 (N_9251,N_6413,N_6416);
nand U9252 (N_9252,N_6506,N_7008);
or U9253 (N_9253,N_6939,N_6683);
and U9254 (N_9254,N_7810,N_6182);
nand U9255 (N_9255,N_7367,N_7381);
and U9256 (N_9256,N_6604,N_6227);
nand U9257 (N_9257,N_7522,N_6620);
or U9258 (N_9258,N_6140,N_6906);
and U9259 (N_9259,N_7975,N_6380);
or U9260 (N_9260,N_6701,N_7641);
and U9261 (N_9261,N_7315,N_7810);
nor U9262 (N_9262,N_6893,N_7456);
or U9263 (N_9263,N_6928,N_6467);
and U9264 (N_9264,N_6561,N_7364);
and U9265 (N_9265,N_6704,N_7344);
nand U9266 (N_9266,N_6770,N_6877);
and U9267 (N_9267,N_7426,N_6768);
and U9268 (N_9268,N_6255,N_6986);
and U9269 (N_9269,N_6599,N_7334);
or U9270 (N_9270,N_6223,N_6970);
or U9271 (N_9271,N_6060,N_7073);
or U9272 (N_9272,N_7428,N_7765);
xor U9273 (N_9273,N_6266,N_6334);
nand U9274 (N_9274,N_6136,N_6920);
nor U9275 (N_9275,N_6604,N_7579);
or U9276 (N_9276,N_6239,N_6064);
and U9277 (N_9277,N_6357,N_6798);
nand U9278 (N_9278,N_7350,N_6482);
nand U9279 (N_9279,N_6188,N_6390);
or U9280 (N_9280,N_7487,N_7495);
or U9281 (N_9281,N_7643,N_7662);
nand U9282 (N_9282,N_7975,N_6996);
and U9283 (N_9283,N_6165,N_6809);
or U9284 (N_9284,N_7674,N_6018);
nand U9285 (N_9285,N_6061,N_6770);
nand U9286 (N_9286,N_6941,N_7541);
and U9287 (N_9287,N_6226,N_7848);
or U9288 (N_9288,N_6088,N_7619);
nand U9289 (N_9289,N_6454,N_7514);
nor U9290 (N_9290,N_7537,N_7395);
nand U9291 (N_9291,N_6817,N_6345);
and U9292 (N_9292,N_6938,N_6607);
nand U9293 (N_9293,N_7942,N_7906);
nor U9294 (N_9294,N_7592,N_6850);
and U9295 (N_9295,N_6313,N_7729);
and U9296 (N_9296,N_7375,N_7028);
and U9297 (N_9297,N_6186,N_7116);
and U9298 (N_9298,N_6056,N_7809);
xnor U9299 (N_9299,N_7345,N_6705);
or U9300 (N_9300,N_6685,N_7742);
nor U9301 (N_9301,N_7435,N_6054);
nand U9302 (N_9302,N_7425,N_6592);
nand U9303 (N_9303,N_7915,N_6480);
nor U9304 (N_9304,N_6867,N_6660);
or U9305 (N_9305,N_6571,N_6121);
nand U9306 (N_9306,N_7454,N_7137);
nor U9307 (N_9307,N_7613,N_6339);
nand U9308 (N_9308,N_6831,N_7275);
and U9309 (N_9309,N_6507,N_7312);
and U9310 (N_9310,N_6006,N_7493);
nand U9311 (N_9311,N_7014,N_7202);
nor U9312 (N_9312,N_6690,N_7487);
nand U9313 (N_9313,N_6540,N_6196);
nor U9314 (N_9314,N_6355,N_7607);
or U9315 (N_9315,N_6812,N_7185);
nor U9316 (N_9316,N_7953,N_7007);
nor U9317 (N_9317,N_7927,N_7177);
nor U9318 (N_9318,N_6511,N_6860);
or U9319 (N_9319,N_6523,N_7403);
and U9320 (N_9320,N_7693,N_6440);
nor U9321 (N_9321,N_7342,N_7961);
or U9322 (N_9322,N_6986,N_6087);
nor U9323 (N_9323,N_6038,N_6806);
nand U9324 (N_9324,N_6978,N_6920);
nand U9325 (N_9325,N_6867,N_7748);
and U9326 (N_9326,N_7687,N_7013);
and U9327 (N_9327,N_6497,N_7847);
and U9328 (N_9328,N_7499,N_7367);
and U9329 (N_9329,N_7772,N_6819);
xnor U9330 (N_9330,N_6525,N_6631);
nor U9331 (N_9331,N_7385,N_6568);
and U9332 (N_9332,N_6096,N_7158);
nor U9333 (N_9333,N_6375,N_6939);
nand U9334 (N_9334,N_7976,N_7304);
or U9335 (N_9335,N_6515,N_6238);
or U9336 (N_9336,N_6662,N_6281);
nor U9337 (N_9337,N_7884,N_6048);
or U9338 (N_9338,N_7480,N_6977);
and U9339 (N_9339,N_6328,N_7616);
nand U9340 (N_9340,N_7474,N_6623);
nor U9341 (N_9341,N_7112,N_6725);
nand U9342 (N_9342,N_6521,N_6833);
nand U9343 (N_9343,N_6054,N_7238);
nor U9344 (N_9344,N_6375,N_6214);
and U9345 (N_9345,N_6631,N_6188);
or U9346 (N_9346,N_6002,N_7091);
nor U9347 (N_9347,N_7610,N_7273);
nand U9348 (N_9348,N_6593,N_7716);
or U9349 (N_9349,N_6571,N_6164);
and U9350 (N_9350,N_6310,N_6324);
nand U9351 (N_9351,N_6394,N_7051);
and U9352 (N_9352,N_6396,N_7768);
nand U9353 (N_9353,N_7221,N_7741);
and U9354 (N_9354,N_6002,N_7876);
nand U9355 (N_9355,N_7840,N_7843);
nor U9356 (N_9356,N_6088,N_6200);
nand U9357 (N_9357,N_7645,N_7020);
nor U9358 (N_9358,N_7052,N_6459);
or U9359 (N_9359,N_7747,N_6811);
and U9360 (N_9360,N_6880,N_6774);
nand U9361 (N_9361,N_6396,N_7016);
or U9362 (N_9362,N_7858,N_6898);
nand U9363 (N_9363,N_6675,N_6646);
nand U9364 (N_9364,N_6489,N_6504);
nand U9365 (N_9365,N_7570,N_7244);
or U9366 (N_9366,N_7268,N_7610);
or U9367 (N_9367,N_7587,N_6548);
and U9368 (N_9368,N_6743,N_6032);
or U9369 (N_9369,N_6938,N_7507);
or U9370 (N_9370,N_6747,N_6155);
xor U9371 (N_9371,N_7524,N_6961);
or U9372 (N_9372,N_6782,N_6603);
nand U9373 (N_9373,N_6779,N_6180);
or U9374 (N_9374,N_6796,N_7812);
nor U9375 (N_9375,N_6207,N_7920);
or U9376 (N_9376,N_7732,N_6927);
or U9377 (N_9377,N_7028,N_7969);
and U9378 (N_9378,N_7295,N_6172);
nor U9379 (N_9379,N_6540,N_7655);
nor U9380 (N_9380,N_6196,N_7911);
nor U9381 (N_9381,N_7480,N_6961);
or U9382 (N_9382,N_7112,N_6430);
nor U9383 (N_9383,N_6751,N_7066);
nand U9384 (N_9384,N_7305,N_7090);
nand U9385 (N_9385,N_6280,N_7764);
nand U9386 (N_9386,N_7118,N_6747);
nor U9387 (N_9387,N_6226,N_7924);
nor U9388 (N_9388,N_7622,N_7015);
or U9389 (N_9389,N_7881,N_7156);
or U9390 (N_9390,N_6279,N_7920);
or U9391 (N_9391,N_7856,N_6923);
nand U9392 (N_9392,N_6709,N_6148);
and U9393 (N_9393,N_6612,N_6362);
nand U9394 (N_9394,N_7465,N_6378);
or U9395 (N_9395,N_6959,N_6660);
nand U9396 (N_9396,N_6207,N_6473);
nand U9397 (N_9397,N_6760,N_6559);
nor U9398 (N_9398,N_7393,N_7681);
and U9399 (N_9399,N_7726,N_7899);
and U9400 (N_9400,N_7791,N_6868);
or U9401 (N_9401,N_7367,N_6284);
nor U9402 (N_9402,N_7669,N_6263);
nand U9403 (N_9403,N_6613,N_7014);
nand U9404 (N_9404,N_6633,N_6499);
and U9405 (N_9405,N_7536,N_7766);
and U9406 (N_9406,N_7813,N_7303);
nand U9407 (N_9407,N_6884,N_7765);
nor U9408 (N_9408,N_7196,N_7937);
nor U9409 (N_9409,N_7882,N_6687);
nor U9410 (N_9410,N_6285,N_6431);
and U9411 (N_9411,N_6605,N_6563);
and U9412 (N_9412,N_7245,N_7454);
or U9413 (N_9413,N_6321,N_6847);
and U9414 (N_9414,N_7222,N_6116);
nand U9415 (N_9415,N_6821,N_6713);
or U9416 (N_9416,N_6919,N_6025);
or U9417 (N_9417,N_6900,N_6538);
or U9418 (N_9418,N_7620,N_6596);
nand U9419 (N_9419,N_6259,N_6100);
and U9420 (N_9420,N_6373,N_6800);
nor U9421 (N_9421,N_7032,N_7014);
and U9422 (N_9422,N_7721,N_7616);
and U9423 (N_9423,N_7726,N_7919);
nor U9424 (N_9424,N_7092,N_6520);
or U9425 (N_9425,N_7442,N_7691);
and U9426 (N_9426,N_6436,N_6899);
or U9427 (N_9427,N_7439,N_6771);
nor U9428 (N_9428,N_6913,N_7717);
nor U9429 (N_9429,N_6003,N_6252);
nor U9430 (N_9430,N_6997,N_7800);
and U9431 (N_9431,N_6643,N_7567);
xnor U9432 (N_9432,N_7402,N_7156);
nor U9433 (N_9433,N_7609,N_7156);
nor U9434 (N_9434,N_7842,N_7399);
nor U9435 (N_9435,N_7829,N_6328);
nand U9436 (N_9436,N_6463,N_6547);
nor U9437 (N_9437,N_6503,N_6403);
and U9438 (N_9438,N_7585,N_7402);
and U9439 (N_9439,N_6346,N_6525);
or U9440 (N_9440,N_7560,N_7673);
nor U9441 (N_9441,N_6972,N_6264);
or U9442 (N_9442,N_7063,N_7471);
nor U9443 (N_9443,N_6420,N_7875);
nand U9444 (N_9444,N_6384,N_6748);
or U9445 (N_9445,N_7239,N_6630);
or U9446 (N_9446,N_6512,N_7106);
nand U9447 (N_9447,N_6501,N_7851);
and U9448 (N_9448,N_6454,N_6962);
and U9449 (N_9449,N_6983,N_6117);
nor U9450 (N_9450,N_6951,N_7188);
and U9451 (N_9451,N_7356,N_6753);
nand U9452 (N_9452,N_6208,N_7618);
nor U9453 (N_9453,N_6385,N_6168);
or U9454 (N_9454,N_6879,N_6730);
nand U9455 (N_9455,N_7449,N_6691);
nor U9456 (N_9456,N_7231,N_6666);
nor U9457 (N_9457,N_7652,N_6990);
nand U9458 (N_9458,N_6826,N_7495);
or U9459 (N_9459,N_7434,N_6208);
nor U9460 (N_9460,N_7787,N_7720);
or U9461 (N_9461,N_6425,N_7218);
nand U9462 (N_9462,N_7030,N_6874);
or U9463 (N_9463,N_7747,N_6064);
or U9464 (N_9464,N_7858,N_6852);
or U9465 (N_9465,N_7721,N_7011);
and U9466 (N_9466,N_6427,N_6750);
nor U9467 (N_9467,N_7762,N_6238);
nor U9468 (N_9468,N_7929,N_7661);
nor U9469 (N_9469,N_6241,N_6219);
nor U9470 (N_9470,N_7806,N_7564);
nand U9471 (N_9471,N_6409,N_6418);
nor U9472 (N_9472,N_6772,N_6831);
and U9473 (N_9473,N_6624,N_6210);
nand U9474 (N_9474,N_7673,N_6284);
nand U9475 (N_9475,N_7081,N_7476);
nor U9476 (N_9476,N_7382,N_7602);
nor U9477 (N_9477,N_6215,N_7519);
or U9478 (N_9478,N_7727,N_6753);
or U9479 (N_9479,N_7199,N_6565);
xor U9480 (N_9480,N_7814,N_7464);
and U9481 (N_9481,N_7136,N_6292);
nand U9482 (N_9482,N_6566,N_7330);
or U9483 (N_9483,N_7079,N_7315);
nor U9484 (N_9484,N_7954,N_7641);
nor U9485 (N_9485,N_7572,N_7907);
or U9486 (N_9486,N_7127,N_6081);
nand U9487 (N_9487,N_7126,N_6034);
or U9488 (N_9488,N_6944,N_7298);
nor U9489 (N_9489,N_7539,N_7228);
or U9490 (N_9490,N_7792,N_6353);
nor U9491 (N_9491,N_6694,N_6383);
nor U9492 (N_9492,N_6277,N_7507);
nor U9493 (N_9493,N_6002,N_7311);
nand U9494 (N_9494,N_6701,N_6525);
nor U9495 (N_9495,N_7957,N_6967);
nor U9496 (N_9496,N_7916,N_6444);
nor U9497 (N_9497,N_7278,N_7303);
nand U9498 (N_9498,N_7022,N_7454);
nor U9499 (N_9499,N_6869,N_6653);
nand U9500 (N_9500,N_7543,N_7718);
nor U9501 (N_9501,N_6284,N_6876);
nor U9502 (N_9502,N_6936,N_7966);
nand U9503 (N_9503,N_6246,N_7559);
nor U9504 (N_9504,N_6499,N_7743);
and U9505 (N_9505,N_6634,N_6791);
nor U9506 (N_9506,N_6267,N_7943);
nor U9507 (N_9507,N_7143,N_7483);
and U9508 (N_9508,N_6084,N_7604);
nand U9509 (N_9509,N_7033,N_7312);
nand U9510 (N_9510,N_6715,N_6271);
nand U9511 (N_9511,N_6954,N_6223);
nor U9512 (N_9512,N_7486,N_6112);
nand U9513 (N_9513,N_6053,N_6802);
or U9514 (N_9514,N_6184,N_7699);
or U9515 (N_9515,N_6785,N_6598);
and U9516 (N_9516,N_7291,N_7193);
nor U9517 (N_9517,N_7309,N_7302);
nand U9518 (N_9518,N_7689,N_6608);
nand U9519 (N_9519,N_6777,N_7384);
nor U9520 (N_9520,N_6692,N_7250);
nand U9521 (N_9521,N_6247,N_6013);
and U9522 (N_9522,N_7838,N_6416);
or U9523 (N_9523,N_6263,N_6450);
or U9524 (N_9524,N_7786,N_6949);
and U9525 (N_9525,N_7854,N_7922);
nand U9526 (N_9526,N_7775,N_7007);
nand U9527 (N_9527,N_6230,N_6207);
nor U9528 (N_9528,N_7156,N_7034);
and U9529 (N_9529,N_6662,N_6254);
and U9530 (N_9530,N_6980,N_6417);
and U9531 (N_9531,N_6617,N_7693);
or U9532 (N_9532,N_7681,N_6744);
nor U9533 (N_9533,N_6540,N_7456);
or U9534 (N_9534,N_6150,N_7933);
nand U9535 (N_9535,N_6366,N_6523);
nor U9536 (N_9536,N_7322,N_7900);
nand U9537 (N_9537,N_6673,N_6506);
nand U9538 (N_9538,N_6221,N_6179);
nor U9539 (N_9539,N_7661,N_7285);
nor U9540 (N_9540,N_6420,N_6960);
nor U9541 (N_9541,N_7864,N_6119);
nor U9542 (N_9542,N_6293,N_7530);
nand U9543 (N_9543,N_6695,N_7353);
or U9544 (N_9544,N_7094,N_6305);
xnor U9545 (N_9545,N_6761,N_7267);
and U9546 (N_9546,N_7619,N_6076);
or U9547 (N_9547,N_6393,N_7848);
nand U9548 (N_9548,N_7289,N_7608);
or U9549 (N_9549,N_7327,N_6236);
nand U9550 (N_9550,N_6238,N_6730);
and U9551 (N_9551,N_6839,N_6271);
nand U9552 (N_9552,N_7902,N_6556);
and U9553 (N_9553,N_7063,N_6435);
nand U9554 (N_9554,N_7245,N_6120);
nor U9555 (N_9555,N_7063,N_6000);
and U9556 (N_9556,N_6221,N_6778);
nand U9557 (N_9557,N_7811,N_6636);
nor U9558 (N_9558,N_7400,N_7647);
and U9559 (N_9559,N_7776,N_6312);
and U9560 (N_9560,N_6264,N_6732);
nor U9561 (N_9561,N_7619,N_7234);
nand U9562 (N_9562,N_7597,N_7222);
or U9563 (N_9563,N_6593,N_7491);
and U9564 (N_9564,N_7572,N_6995);
nand U9565 (N_9565,N_7305,N_7948);
nand U9566 (N_9566,N_7325,N_7309);
and U9567 (N_9567,N_6425,N_6255);
or U9568 (N_9568,N_6121,N_6339);
nand U9569 (N_9569,N_7222,N_6492);
nor U9570 (N_9570,N_7760,N_6256);
xnor U9571 (N_9571,N_6305,N_7610);
nand U9572 (N_9572,N_7038,N_6309);
nand U9573 (N_9573,N_7447,N_6527);
nand U9574 (N_9574,N_6023,N_6970);
or U9575 (N_9575,N_7090,N_6758);
nor U9576 (N_9576,N_6657,N_7622);
nand U9577 (N_9577,N_7275,N_6077);
nor U9578 (N_9578,N_7305,N_7298);
and U9579 (N_9579,N_6367,N_7992);
or U9580 (N_9580,N_7996,N_6484);
or U9581 (N_9581,N_6698,N_6756);
and U9582 (N_9582,N_7344,N_7144);
nor U9583 (N_9583,N_7368,N_6712);
or U9584 (N_9584,N_7051,N_6402);
xnor U9585 (N_9585,N_7753,N_7563);
nand U9586 (N_9586,N_6180,N_7234);
nand U9587 (N_9587,N_6452,N_6692);
and U9588 (N_9588,N_7247,N_7652);
nand U9589 (N_9589,N_6041,N_6475);
nand U9590 (N_9590,N_6250,N_6283);
nor U9591 (N_9591,N_7573,N_7633);
and U9592 (N_9592,N_6798,N_7601);
nor U9593 (N_9593,N_6331,N_6660);
and U9594 (N_9594,N_6322,N_7242);
or U9595 (N_9595,N_6782,N_7207);
or U9596 (N_9596,N_7901,N_7131);
or U9597 (N_9597,N_7299,N_6658);
or U9598 (N_9598,N_6394,N_7132);
and U9599 (N_9599,N_7967,N_6146);
nand U9600 (N_9600,N_7590,N_7920);
and U9601 (N_9601,N_7330,N_6951);
or U9602 (N_9602,N_7214,N_7659);
nor U9603 (N_9603,N_6149,N_6341);
nand U9604 (N_9604,N_7157,N_6776);
or U9605 (N_9605,N_7434,N_6119);
and U9606 (N_9606,N_6200,N_7034);
nand U9607 (N_9607,N_6480,N_6435);
and U9608 (N_9608,N_6821,N_7066);
and U9609 (N_9609,N_6073,N_7596);
nor U9610 (N_9610,N_6224,N_6295);
xnor U9611 (N_9611,N_7112,N_6720);
nand U9612 (N_9612,N_7349,N_6231);
nor U9613 (N_9613,N_7878,N_7729);
and U9614 (N_9614,N_6066,N_6811);
nand U9615 (N_9615,N_7593,N_7731);
nand U9616 (N_9616,N_6115,N_6821);
or U9617 (N_9617,N_6051,N_6719);
nor U9618 (N_9618,N_6342,N_6066);
nor U9619 (N_9619,N_7346,N_6181);
nor U9620 (N_9620,N_7947,N_6461);
and U9621 (N_9621,N_6084,N_6635);
and U9622 (N_9622,N_6803,N_6572);
or U9623 (N_9623,N_7293,N_7521);
and U9624 (N_9624,N_6487,N_7597);
or U9625 (N_9625,N_7564,N_6633);
nand U9626 (N_9626,N_6178,N_6083);
nor U9627 (N_9627,N_7986,N_7739);
or U9628 (N_9628,N_6977,N_6816);
or U9629 (N_9629,N_6613,N_6371);
nor U9630 (N_9630,N_7631,N_7637);
or U9631 (N_9631,N_7002,N_7906);
nor U9632 (N_9632,N_6322,N_7164);
or U9633 (N_9633,N_7673,N_7428);
and U9634 (N_9634,N_6278,N_6785);
nor U9635 (N_9635,N_6213,N_7764);
or U9636 (N_9636,N_6656,N_7190);
or U9637 (N_9637,N_7368,N_6921);
and U9638 (N_9638,N_6319,N_6896);
or U9639 (N_9639,N_7124,N_6515);
and U9640 (N_9640,N_6523,N_7430);
and U9641 (N_9641,N_7231,N_7585);
nor U9642 (N_9642,N_7837,N_7957);
nor U9643 (N_9643,N_7577,N_7455);
nand U9644 (N_9644,N_6148,N_6615);
nand U9645 (N_9645,N_7206,N_7309);
or U9646 (N_9646,N_6788,N_7565);
and U9647 (N_9647,N_6867,N_7011);
or U9648 (N_9648,N_7920,N_6488);
nand U9649 (N_9649,N_6173,N_7095);
nand U9650 (N_9650,N_7569,N_6465);
nand U9651 (N_9651,N_7507,N_7030);
nor U9652 (N_9652,N_7839,N_6573);
nor U9653 (N_9653,N_6835,N_6264);
nand U9654 (N_9654,N_7958,N_7955);
nand U9655 (N_9655,N_7070,N_7682);
nor U9656 (N_9656,N_7458,N_6722);
nand U9657 (N_9657,N_6913,N_6553);
and U9658 (N_9658,N_7205,N_6247);
and U9659 (N_9659,N_6480,N_6873);
nand U9660 (N_9660,N_7187,N_7396);
or U9661 (N_9661,N_6170,N_6030);
nand U9662 (N_9662,N_7717,N_7860);
or U9663 (N_9663,N_6231,N_6162);
or U9664 (N_9664,N_7830,N_6542);
nand U9665 (N_9665,N_6159,N_6470);
nand U9666 (N_9666,N_7488,N_7582);
or U9667 (N_9667,N_6472,N_7707);
and U9668 (N_9668,N_6291,N_6908);
nand U9669 (N_9669,N_6969,N_7471);
nor U9670 (N_9670,N_6143,N_7422);
nand U9671 (N_9671,N_7281,N_7020);
or U9672 (N_9672,N_6355,N_6829);
nand U9673 (N_9673,N_6000,N_7814);
nor U9674 (N_9674,N_6120,N_7823);
nor U9675 (N_9675,N_7361,N_6883);
xnor U9676 (N_9676,N_7066,N_6776);
and U9677 (N_9677,N_6907,N_6104);
nand U9678 (N_9678,N_7195,N_7604);
nand U9679 (N_9679,N_7129,N_7088);
and U9680 (N_9680,N_6213,N_7367);
nor U9681 (N_9681,N_6093,N_7919);
or U9682 (N_9682,N_6071,N_6216);
nor U9683 (N_9683,N_7861,N_7353);
or U9684 (N_9684,N_6012,N_6917);
or U9685 (N_9685,N_6043,N_7572);
and U9686 (N_9686,N_7285,N_6419);
nand U9687 (N_9687,N_6862,N_6172);
nor U9688 (N_9688,N_7968,N_7012);
or U9689 (N_9689,N_6543,N_6767);
or U9690 (N_9690,N_7291,N_6860);
nor U9691 (N_9691,N_7154,N_7808);
nor U9692 (N_9692,N_6521,N_6103);
nor U9693 (N_9693,N_7834,N_7909);
and U9694 (N_9694,N_7310,N_7555);
or U9695 (N_9695,N_7787,N_6139);
and U9696 (N_9696,N_6140,N_6279);
nand U9697 (N_9697,N_6804,N_6876);
nand U9698 (N_9698,N_7115,N_7053);
nand U9699 (N_9699,N_7218,N_6900);
nor U9700 (N_9700,N_6601,N_7198);
nand U9701 (N_9701,N_7988,N_7147);
nand U9702 (N_9702,N_7451,N_7529);
and U9703 (N_9703,N_7534,N_6469);
nor U9704 (N_9704,N_7431,N_6045);
or U9705 (N_9705,N_6675,N_6248);
or U9706 (N_9706,N_7000,N_6835);
or U9707 (N_9707,N_7418,N_6695);
and U9708 (N_9708,N_7337,N_6353);
or U9709 (N_9709,N_6450,N_7886);
nor U9710 (N_9710,N_6837,N_6250);
nor U9711 (N_9711,N_7592,N_6570);
and U9712 (N_9712,N_7398,N_7787);
nor U9713 (N_9713,N_6688,N_7187);
or U9714 (N_9714,N_7888,N_7556);
and U9715 (N_9715,N_6797,N_7523);
and U9716 (N_9716,N_7700,N_7371);
and U9717 (N_9717,N_6134,N_7379);
xor U9718 (N_9718,N_6472,N_6187);
nor U9719 (N_9719,N_7708,N_7346);
or U9720 (N_9720,N_7496,N_6370);
or U9721 (N_9721,N_6759,N_7810);
nor U9722 (N_9722,N_6793,N_6425);
nor U9723 (N_9723,N_7447,N_6195);
nand U9724 (N_9724,N_7361,N_6504);
nor U9725 (N_9725,N_7289,N_6390);
and U9726 (N_9726,N_6117,N_6302);
and U9727 (N_9727,N_6808,N_6540);
or U9728 (N_9728,N_6850,N_6904);
nand U9729 (N_9729,N_7155,N_7576);
or U9730 (N_9730,N_7808,N_7394);
nor U9731 (N_9731,N_7069,N_7859);
or U9732 (N_9732,N_7054,N_6984);
nor U9733 (N_9733,N_7917,N_6907);
and U9734 (N_9734,N_6846,N_7378);
and U9735 (N_9735,N_6446,N_6950);
nand U9736 (N_9736,N_7595,N_6912);
and U9737 (N_9737,N_7447,N_6510);
nand U9738 (N_9738,N_6211,N_7235);
nor U9739 (N_9739,N_6046,N_6914);
nor U9740 (N_9740,N_7783,N_6674);
and U9741 (N_9741,N_6607,N_7447);
or U9742 (N_9742,N_6323,N_7898);
xnor U9743 (N_9743,N_7522,N_6595);
and U9744 (N_9744,N_6481,N_6907);
and U9745 (N_9745,N_6910,N_7071);
or U9746 (N_9746,N_6516,N_6317);
or U9747 (N_9747,N_7103,N_7606);
nor U9748 (N_9748,N_7124,N_7491);
nand U9749 (N_9749,N_6707,N_7525);
nor U9750 (N_9750,N_6003,N_7444);
or U9751 (N_9751,N_7005,N_7376);
nor U9752 (N_9752,N_6257,N_7856);
nand U9753 (N_9753,N_7886,N_7315);
or U9754 (N_9754,N_7777,N_7319);
or U9755 (N_9755,N_6881,N_6270);
nor U9756 (N_9756,N_6749,N_7638);
or U9757 (N_9757,N_7633,N_6773);
nand U9758 (N_9758,N_7711,N_7099);
and U9759 (N_9759,N_7162,N_7383);
nand U9760 (N_9760,N_6571,N_7932);
nand U9761 (N_9761,N_7349,N_6550);
nand U9762 (N_9762,N_7846,N_7868);
or U9763 (N_9763,N_7378,N_7667);
or U9764 (N_9764,N_7795,N_7065);
nor U9765 (N_9765,N_6220,N_6521);
or U9766 (N_9766,N_7626,N_6797);
nor U9767 (N_9767,N_6706,N_6654);
nand U9768 (N_9768,N_6620,N_7018);
nor U9769 (N_9769,N_6182,N_6572);
nand U9770 (N_9770,N_6566,N_6550);
and U9771 (N_9771,N_6902,N_7747);
and U9772 (N_9772,N_7286,N_6981);
or U9773 (N_9773,N_6213,N_7957);
nand U9774 (N_9774,N_7000,N_6107);
nor U9775 (N_9775,N_7807,N_7990);
nor U9776 (N_9776,N_7731,N_7654);
nor U9777 (N_9777,N_6555,N_6491);
nor U9778 (N_9778,N_7648,N_7935);
or U9779 (N_9779,N_6602,N_6251);
and U9780 (N_9780,N_7285,N_7239);
and U9781 (N_9781,N_6902,N_7654);
or U9782 (N_9782,N_6450,N_6398);
nor U9783 (N_9783,N_7706,N_6958);
nor U9784 (N_9784,N_6483,N_6693);
nand U9785 (N_9785,N_6742,N_6015);
nand U9786 (N_9786,N_6007,N_6660);
or U9787 (N_9787,N_6648,N_7365);
or U9788 (N_9788,N_6470,N_7201);
and U9789 (N_9789,N_6544,N_7396);
nand U9790 (N_9790,N_6334,N_7056);
and U9791 (N_9791,N_7575,N_6281);
or U9792 (N_9792,N_7950,N_6617);
nand U9793 (N_9793,N_7167,N_7808);
or U9794 (N_9794,N_6404,N_7378);
nand U9795 (N_9795,N_7856,N_6598);
nor U9796 (N_9796,N_7593,N_7068);
nand U9797 (N_9797,N_6771,N_6056);
and U9798 (N_9798,N_7535,N_6782);
nand U9799 (N_9799,N_7369,N_6957);
nand U9800 (N_9800,N_7762,N_6294);
or U9801 (N_9801,N_7724,N_6764);
and U9802 (N_9802,N_6246,N_7079);
nand U9803 (N_9803,N_6167,N_6066);
nand U9804 (N_9804,N_7000,N_7742);
nand U9805 (N_9805,N_7421,N_7430);
nand U9806 (N_9806,N_6945,N_7284);
and U9807 (N_9807,N_6827,N_6964);
nand U9808 (N_9808,N_7611,N_6641);
or U9809 (N_9809,N_7545,N_7275);
nand U9810 (N_9810,N_7607,N_6506);
or U9811 (N_9811,N_6861,N_6090);
nand U9812 (N_9812,N_7849,N_6928);
nand U9813 (N_9813,N_7547,N_6552);
or U9814 (N_9814,N_6833,N_6305);
nor U9815 (N_9815,N_7922,N_7734);
nor U9816 (N_9816,N_7959,N_7683);
or U9817 (N_9817,N_7974,N_7695);
nor U9818 (N_9818,N_7000,N_6962);
nand U9819 (N_9819,N_7115,N_7242);
nor U9820 (N_9820,N_6764,N_7526);
nand U9821 (N_9821,N_6071,N_7851);
or U9822 (N_9822,N_7468,N_7506);
and U9823 (N_9823,N_7147,N_6030);
or U9824 (N_9824,N_6179,N_6853);
nand U9825 (N_9825,N_6791,N_6224);
nor U9826 (N_9826,N_7191,N_7619);
nand U9827 (N_9827,N_6247,N_6364);
nand U9828 (N_9828,N_6656,N_7732);
nor U9829 (N_9829,N_7062,N_7603);
and U9830 (N_9830,N_7830,N_7989);
nor U9831 (N_9831,N_7152,N_6821);
or U9832 (N_9832,N_6317,N_7397);
nand U9833 (N_9833,N_6268,N_7454);
or U9834 (N_9834,N_7448,N_6570);
nor U9835 (N_9835,N_7687,N_6253);
nor U9836 (N_9836,N_7481,N_6566);
or U9837 (N_9837,N_6092,N_6120);
nor U9838 (N_9838,N_7994,N_7000);
or U9839 (N_9839,N_6300,N_6587);
or U9840 (N_9840,N_7057,N_6356);
nor U9841 (N_9841,N_7225,N_7038);
or U9842 (N_9842,N_7676,N_6941);
nand U9843 (N_9843,N_7356,N_7884);
nor U9844 (N_9844,N_6343,N_7444);
and U9845 (N_9845,N_7991,N_7405);
nand U9846 (N_9846,N_6114,N_6638);
nor U9847 (N_9847,N_6043,N_7889);
xnor U9848 (N_9848,N_6726,N_7630);
and U9849 (N_9849,N_7446,N_6448);
or U9850 (N_9850,N_6107,N_7520);
nand U9851 (N_9851,N_6553,N_7132);
and U9852 (N_9852,N_6468,N_7493);
or U9853 (N_9853,N_7924,N_7994);
and U9854 (N_9854,N_7859,N_7186);
nor U9855 (N_9855,N_6144,N_6753);
and U9856 (N_9856,N_7817,N_7390);
and U9857 (N_9857,N_7038,N_7674);
nand U9858 (N_9858,N_7792,N_7067);
nor U9859 (N_9859,N_7326,N_7023);
nor U9860 (N_9860,N_6381,N_6322);
nand U9861 (N_9861,N_7594,N_6460);
nand U9862 (N_9862,N_7120,N_6026);
nand U9863 (N_9863,N_7912,N_7695);
and U9864 (N_9864,N_7992,N_6711);
nor U9865 (N_9865,N_6299,N_6646);
and U9866 (N_9866,N_7152,N_7518);
and U9867 (N_9867,N_7058,N_7859);
or U9868 (N_9868,N_6912,N_6927);
and U9869 (N_9869,N_6527,N_7619);
nor U9870 (N_9870,N_7121,N_6412);
and U9871 (N_9871,N_6100,N_7160);
and U9872 (N_9872,N_7765,N_6762);
nand U9873 (N_9873,N_6730,N_7606);
nor U9874 (N_9874,N_7595,N_7266);
and U9875 (N_9875,N_6298,N_7719);
nand U9876 (N_9876,N_6796,N_6762);
and U9877 (N_9877,N_7122,N_7800);
and U9878 (N_9878,N_6064,N_7387);
nand U9879 (N_9879,N_7057,N_7161);
nor U9880 (N_9880,N_6968,N_6191);
or U9881 (N_9881,N_6787,N_6191);
or U9882 (N_9882,N_6647,N_7914);
or U9883 (N_9883,N_7586,N_6891);
nor U9884 (N_9884,N_6321,N_7573);
nand U9885 (N_9885,N_7104,N_6879);
or U9886 (N_9886,N_7194,N_6211);
and U9887 (N_9887,N_7203,N_6918);
nor U9888 (N_9888,N_7377,N_7753);
nor U9889 (N_9889,N_7740,N_7893);
nor U9890 (N_9890,N_7958,N_7670);
or U9891 (N_9891,N_6746,N_7109);
nand U9892 (N_9892,N_6260,N_7028);
nor U9893 (N_9893,N_6028,N_7280);
and U9894 (N_9894,N_6035,N_7452);
and U9895 (N_9895,N_6697,N_6984);
and U9896 (N_9896,N_6534,N_7541);
nor U9897 (N_9897,N_7765,N_7285);
and U9898 (N_9898,N_7874,N_6893);
and U9899 (N_9899,N_6548,N_6857);
or U9900 (N_9900,N_6657,N_6679);
nor U9901 (N_9901,N_7675,N_7979);
nor U9902 (N_9902,N_7154,N_6256);
and U9903 (N_9903,N_7031,N_6018);
and U9904 (N_9904,N_6744,N_7611);
nor U9905 (N_9905,N_6913,N_6483);
nor U9906 (N_9906,N_7765,N_6663);
or U9907 (N_9907,N_6184,N_7296);
or U9908 (N_9908,N_7145,N_7743);
nor U9909 (N_9909,N_6353,N_7992);
and U9910 (N_9910,N_7995,N_7052);
and U9911 (N_9911,N_7517,N_6900);
and U9912 (N_9912,N_7295,N_6047);
or U9913 (N_9913,N_6711,N_7017);
or U9914 (N_9914,N_7921,N_6999);
and U9915 (N_9915,N_6292,N_6572);
and U9916 (N_9916,N_6810,N_7662);
and U9917 (N_9917,N_6029,N_6265);
and U9918 (N_9918,N_7585,N_7563);
nor U9919 (N_9919,N_7183,N_6709);
nand U9920 (N_9920,N_6587,N_6973);
nand U9921 (N_9921,N_6560,N_6746);
nor U9922 (N_9922,N_7324,N_7116);
and U9923 (N_9923,N_7659,N_7966);
or U9924 (N_9924,N_6905,N_7599);
nand U9925 (N_9925,N_7225,N_7136);
nor U9926 (N_9926,N_7162,N_6741);
nor U9927 (N_9927,N_7050,N_6913);
nand U9928 (N_9928,N_7595,N_7611);
or U9929 (N_9929,N_7095,N_7272);
or U9930 (N_9930,N_7666,N_7003);
nand U9931 (N_9931,N_7455,N_6808);
nand U9932 (N_9932,N_7504,N_7766);
or U9933 (N_9933,N_6348,N_7479);
or U9934 (N_9934,N_7131,N_7657);
nand U9935 (N_9935,N_6720,N_7412);
nand U9936 (N_9936,N_7274,N_6762);
and U9937 (N_9937,N_6392,N_6122);
nand U9938 (N_9938,N_6686,N_7930);
nor U9939 (N_9939,N_7142,N_7569);
nor U9940 (N_9940,N_6958,N_7927);
nor U9941 (N_9941,N_7241,N_7951);
nand U9942 (N_9942,N_7588,N_6674);
nor U9943 (N_9943,N_6394,N_6128);
and U9944 (N_9944,N_7202,N_7138);
and U9945 (N_9945,N_7681,N_6413);
nand U9946 (N_9946,N_6633,N_7955);
or U9947 (N_9947,N_7907,N_6822);
nor U9948 (N_9948,N_7242,N_7255);
or U9949 (N_9949,N_6722,N_6221);
nor U9950 (N_9950,N_6598,N_6654);
or U9951 (N_9951,N_6691,N_7428);
or U9952 (N_9952,N_7923,N_6981);
and U9953 (N_9953,N_6967,N_7577);
and U9954 (N_9954,N_7367,N_6280);
or U9955 (N_9955,N_6702,N_6815);
nor U9956 (N_9956,N_7896,N_6658);
and U9957 (N_9957,N_6440,N_7463);
nor U9958 (N_9958,N_6727,N_6761);
or U9959 (N_9959,N_6669,N_7415);
and U9960 (N_9960,N_7671,N_6490);
nor U9961 (N_9961,N_6182,N_6825);
nand U9962 (N_9962,N_6946,N_6580);
nor U9963 (N_9963,N_7695,N_7091);
nand U9964 (N_9964,N_7441,N_6179);
and U9965 (N_9965,N_7993,N_7985);
or U9966 (N_9966,N_7022,N_6654);
nor U9967 (N_9967,N_7243,N_7723);
nand U9968 (N_9968,N_7585,N_7001);
nand U9969 (N_9969,N_7466,N_6695);
nor U9970 (N_9970,N_6561,N_6625);
or U9971 (N_9971,N_6380,N_6956);
nor U9972 (N_9972,N_7531,N_7190);
or U9973 (N_9973,N_7879,N_6037);
or U9974 (N_9974,N_7354,N_7468);
and U9975 (N_9975,N_6549,N_7221);
nor U9976 (N_9976,N_6139,N_6739);
nor U9977 (N_9977,N_7015,N_6022);
nor U9978 (N_9978,N_6657,N_7949);
nand U9979 (N_9979,N_7532,N_7577);
and U9980 (N_9980,N_6652,N_6737);
and U9981 (N_9981,N_6915,N_7063);
nor U9982 (N_9982,N_7661,N_7817);
nor U9983 (N_9983,N_6628,N_7540);
nand U9984 (N_9984,N_7906,N_7281);
or U9985 (N_9985,N_6422,N_7768);
or U9986 (N_9986,N_6179,N_7371);
and U9987 (N_9987,N_7121,N_7715);
nand U9988 (N_9988,N_6037,N_6249);
or U9989 (N_9989,N_7070,N_7458);
or U9990 (N_9990,N_7114,N_7647);
and U9991 (N_9991,N_7933,N_7324);
nand U9992 (N_9992,N_7127,N_7167);
nand U9993 (N_9993,N_6950,N_7686);
nand U9994 (N_9994,N_7565,N_7998);
nor U9995 (N_9995,N_7674,N_6980);
nand U9996 (N_9996,N_6494,N_6090);
and U9997 (N_9997,N_7652,N_7529);
or U9998 (N_9998,N_6232,N_7234);
and U9999 (N_9999,N_7576,N_7001);
and UO_0 (O_0,N_9342,N_9133);
or UO_1 (O_1,N_8424,N_8632);
or UO_2 (O_2,N_9909,N_8415);
nor UO_3 (O_3,N_8299,N_9692);
nand UO_4 (O_4,N_8801,N_8274);
or UO_5 (O_5,N_8828,N_9084);
and UO_6 (O_6,N_9581,N_8396);
nand UO_7 (O_7,N_8595,N_8936);
nand UO_8 (O_8,N_8164,N_9366);
nand UO_9 (O_9,N_9756,N_9644);
or UO_10 (O_10,N_9855,N_8699);
or UO_11 (O_11,N_9596,N_9691);
nand UO_12 (O_12,N_8572,N_8496);
nand UO_13 (O_13,N_9716,N_8811);
and UO_14 (O_14,N_9982,N_9006);
nor UO_15 (O_15,N_9954,N_9584);
nand UO_16 (O_16,N_8513,N_9633);
and UO_17 (O_17,N_9424,N_8069);
nor UO_18 (O_18,N_8093,N_9327);
and UO_19 (O_19,N_9058,N_8590);
or UO_20 (O_20,N_8559,N_8237);
nor UO_21 (O_21,N_9421,N_9773);
and UO_22 (O_22,N_8933,N_9358);
nand UO_23 (O_23,N_9919,N_9175);
or UO_24 (O_24,N_8119,N_8778);
nand UO_25 (O_25,N_9764,N_9190);
and UO_26 (O_26,N_8623,N_8388);
and UO_27 (O_27,N_8710,N_8187);
or UO_28 (O_28,N_8494,N_8667);
and UO_29 (O_29,N_8246,N_9630);
nand UO_30 (O_30,N_9602,N_8136);
and UO_31 (O_31,N_8028,N_8271);
and UO_32 (O_32,N_9997,N_8967);
or UO_33 (O_33,N_8938,N_9635);
and UO_34 (O_34,N_9244,N_9809);
nand UO_35 (O_35,N_9835,N_8498);
nand UO_36 (O_36,N_9607,N_8926);
nand UO_37 (O_37,N_8514,N_9659);
xnor UO_38 (O_38,N_9873,N_9243);
or UO_39 (O_39,N_9878,N_8740);
nand UO_40 (O_40,N_9844,N_8975);
nor UO_41 (O_41,N_8690,N_9286);
nor UO_42 (O_42,N_8642,N_9488);
and UO_43 (O_43,N_9709,N_8989);
nand UO_44 (O_44,N_8780,N_9673);
or UO_45 (O_45,N_8238,N_8333);
and UO_46 (O_46,N_8945,N_9622);
nand UO_47 (O_47,N_9329,N_8914);
nand UO_48 (O_48,N_9300,N_9715);
nor UO_49 (O_49,N_8368,N_8308);
or UO_50 (O_50,N_9128,N_8353);
or UO_51 (O_51,N_8749,N_8488);
nand UO_52 (O_52,N_9034,N_9224);
nand UO_53 (O_53,N_8545,N_9263);
nand UO_54 (O_54,N_8402,N_8501);
nand UO_55 (O_55,N_9568,N_8554);
or UO_56 (O_56,N_8739,N_8586);
or UO_57 (O_57,N_9718,N_8422);
nor UO_58 (O_58,N_8949,N_8864);
nor UO_59 (O_59,N_9428,N_8845);
nor UO_60 (O_60,N_8460,N_9796);
or UO_61 (O_61,N_8820,N_9642);
and UO_62 (O_62,N_9615,N_9432);
nand UO_63 (O_63,N_8678,N_9566);
nor UO_64 (O_64,N_8929,N_8195);
nand UO_65 (O_65,N_9143,N_8796);
nand UO_66 (O_66,N_9879,N_9041);
or UO_67 (O_67,N_9916,N_8003);
nor UO_68 (O_68,N_8986,N_9904);
nand UO_69 (O_69,N_8311,N_8305);
or UO_70 (O_70,N_9524,N_9818);
nor UO_71 (O_71,N_8960,N_9409);
and UO_72 (O_72,N_8483,N_8022);
nand UO_73 (O_73,N_9576,N_9350);
and UO_74 (O_74,N_9441,N_8384);
nand UO_75 (O_75,N_8248,N_8042);
nand UO_76 (O_76,N_8903,N_8024);
nor UO_77 (O_77,N_9407,N_8755);
and UO_78 (O_78,N_9491,N_8371);
or UO_79 (O_79,N_8830,N_8961);
and UO_80 (O_80,N_9532,N_8329);
nor UO_81 (O_81,N_8116,N_9823);
and UO_82 (O_82,N_8529,N_9134);
nand UO_83 (O_83,N_8980,N_9340);
nand UO_84 (O_84,N_9621,N_9341);
and UO_85 (O_85,N_9089,N_8844);
nand UO_86 (O_86,N_8279,N_8681);
nand UO_87 (O_87,N_8410,N_8592);
nand UO_88 (O_88,N_8290,N_9578);
and UO_89 (O_89,N_9755,N_9145);
or UO_90 (O_90,N_9092,N_9708);
or UO_91 (O_91,N_8139,N_8858);
nor UO_92 (O_92,N_9923,N_9198);
nand UO_93 (O_93,N_8197,N_9189);
or UO_94 (O_94,N_8626,N_8800);
nand UO_95 (O_95,N_9192,N_9012);
nand UO_96 (O_96,N_9082,N_9336);
and UO_97 (O_97,N_8480,N_8132);
and UO_98 (O_98,N_9634,N_9011);
xnor UO_99 (O_99,N_9745,N_8898);
nor UO_100 (O_100,N_9298,N_9217);
nand UO_101 (O_101,N_8120,N_9452);
nand UO_102 (O_102,N_9753,N_9639);
and UO_103 (O_103,N_8382,N_9972);
and UO_104 (O_104,N_9683,N_9283);
and UO_105 (O_105,N_9461,N_8807);
nor UO_106 (O_106,N_9023,N_8567);
nand UO_107 (O_107,N_8922,N_8735);
and UO_108 (O_108,N_8923,N_8704);
nand UO_109 (O_109,N_9103,N_9958);
nand UO_110 (O_110,N_9988,N_8231);
or UO_111 (O_111,N_9454,N_9132);
or UO_112 (O_112,N_8066,N_8239);
nor UO_113 (O_113,N_9724,N_8565);
and UO_114 (O_114,N_9876,N_9487);
and UO_115 (O_115,N_9646,N_8478);
nand UO_116 (O_116,N_8365,N_8751);
and UO_117 (O_117,N_9647,N_9155);
nor UO_118 (O_118,N_9557,N_9864);
or UO_119 (O_119,N_9613,N_8385);
nor UO_120 (O_120,N_9901,N_9817);
or UO_121 (O_121,N_8899,N_9881);
nand UO_122 (O_122,N_9885,N_9385);
nand UO_123 (O_123,N_9250,N_8229);
or UO_124 (O_124,N_8953,N_9146);
or UO_125 (O_125,N_9111,N_8769);
nand UO_126 (O_126,N_9404,N_8457);
or UO_127 (O_127,N_8049,N_8935);
nand UO_128 (O_128,N_8890,N_8547);
nor UO_129 (O_129,N_9582,N_8993);
or UO_130 (O_130,N_9882,N_9285);
nor UO_131 (O_131,N_9181,N_9625);
nand UO_132 (O_132,N_9603,N_8319);
xnor UO_133 (O_133,N_8802,N_9321);
nand UO_134 (O_134,N_9542,N_9776);
nor UO_135 (O_135,N_9239,N_8679);
or UO_136 (O_136,N_8915,N_8880);
nor UO_137 (O_137,N_9307,N_9706);
and UO_138 (O_138,N_9938,N_9831);
or UO_139 (O_139,N_9924,N_8249);
or UO_140 (O_140,N_9883,N_8883);
and UO_141 (O_141,N_9860,N_8253);
nor UO_142 (O_142,N_9196,N_8613);
nor UO_143 (O_143,N_8798,N_8100);
and UO_144 (O_144,N_8712,N_9076);
xnor UO_145 (O_145,N_9771,N_8026);
nor UO_146 (O_146,N_9429,N_8439);
nor UO_147 (O_147,N_9124,N_9932);
nor UO_148 (O_148,N_9278,N_9083);
and UO_149 (O_149,N_8436,N_8286);
or UO_150 (O_150,N_8909,N_8325);
or UO_151 (O_151,N_8192,N_9317);
nand UO_152 (O_152,N_8355,N_8487);
or UO_153 (O_153,N_9186,N_8574);
or UO_154 (O_154,N_8320,N_9370);
and UO_155 (O_155,N_8255,N_9178);
nor UO_156 (O_156,N_8448,N_8694);
xor UO_157 (O_157,N_8387,N_9812);
nand UO_158 (O_158,N_9987,N_9100);
nand UO_159 (O_159,N_8427,N_8486);
and UO_160 (O_160,N_8101,N_9721);
or UO_161 (O_161,N_9090,N_8443);
or UO_162 (O_162,N_9609,N_9655);
and UO_163 (O_163,N_9216,N_8757);
nor UO_164 (O_164,N_9523,N_8930);
nand UO_165 (O_165,N_8301,N_9334);
and UO_166 (O_166,N_8548,N_9995);
or UO_167 (O_167,N_9117,N_9526);
or UO_168 (O_168,N_8435,N_9116);
and UO_169 (O_169,N_8153,N_8074);
nor UO_170 (O_170,N_9115,N_8170);
nand UO_171 (O_171,N_8393,N_9159);
or UO_172 (O_172,N_8978,N_8686);
nor UO_173 (O_173,N_8401,N_9797);
nor UO_174 (O_174,N_9269,N_8639);
and UO_175 (O_175,N_8538,N_8045);
and UO_176 (O_176,N_9031,N_9824);
and UO_177 (O_177,N_8596,N_8175);
and UO_178 (O_178,N_9900,N_9547);
or UO_179 (O_179,N_8896,N_8018);
nor UO_180 (O_180,N_8614,N_8150);
or UO_181 (O_181,N_9463,N_9019);
and UO_182 (O_182,N_9983,N_8783);
nand UO_183 (O_183,N_9276,N_9913);
or UO_184 (O_184,N_9308,N_8671);
nor UO_185 (O_185,N_9373,N_8793);
or UO_186 (O_186,N_8672,N_8376);
nand UO_187 (O_187,N_8616,N_8321);
xnor UO_188 (O_188,N_9653,N_9455);
nand UO_189 (O_189,N_8144,N_9238);
or UO_190 (O_190,N_9767,N_9562);
nor UO_191 (O_191,N_9629,N_8797);
and UO_192 (O_192,N_9412,N_9726);
or UO_193 (O_193,N_9788,N_9335);
or UO_194 (O_194,N_9234,N_9548);
or UO_195 (O_195,N_8577,N_9331);
or UO_196 (O_196,N_9142,N_9670);
and UO_197 (O_197,N_8588,N_9386);
and UO_198 (O_198,N_9168,N_9322);
nor UO_199 (O_199,N_9515,N_8799);
nand UO_200 (O_200,N_8726,N_8475);
nand UO_201 (O_201,N_8428,N_8189);
and UO_202 (O_202,N_9471,N_8640);
or UO_203 (O_203,N_8723,N_8736);
or UO_204 (O_204,N_8622,N_9383);
nand UO_205 (O_205,N_9888,N_9390);
and UO_206 (O_206,N_8283,N_8029);
nor UO_207 (O_207,N_8766,N_8416);
nor UO_208 (O_208,N_9606,N_9561);
or UO_209 (O_209,N_9815,N_8179);
and UO_210 (O_210,N_8528,N_9230);
nand UO_211 (O_211,N_9389,N_9554);
nand UO_212 (O_212,N_9467,N_9039);
nand UO_213 (O_213,N_8183,N_9918);
and UO_214 (O_214,N_9460,N_8791);
nand UO_215 (O_215,N_8971,N_9804);
and UO_216 (O_216,N_8708,N_8206);
nor UO_217 (O_217,N_9852,N_9037);
nor UO_218 (O_218,N_9534,N_8937);
nor UO_219 (O_219,N_8234,N_8663);
or UO_220 (O_220,N_9387,N_8096);
or UO_221 (O_221,N_9937,N_8342);
nor UO_222 (O_222,N_9931,N_8805);
and UO_223 (O_223,N_8522,N_8602);
nand UO_224 (O_224,N_8134,N_8142);
nand UO_225 (O_225,N_8364,N_8036);
nor UO_226 (O_226,N_9406,N_9541);
nor UO_227 (O_227,N_9624,N_8784);
nand UO_228 (O_228,N_8223,N_8835);
or UO_229 (O_229,N_9200,N_8138);
nand UO_230 (O_230,N_8445,N_9648);
nor UO_231 (O_231,N_8786,N_8532);
and UO_232 (O_232,N_8979,N_8657);
or UO_233 (O_233,N_8920,N_8169);
nand UO_234 (O_234,N_8982,N_9710);
nand UO_235 (O_235,N_9574,N_9068);
or UO_236 (O_236,N_9097,N_9669);
nor UO_237 (O_237,N_8853,N_8481);
and UO_238 (O_238,N_8997,N_9054);
nand UO_239 (O_239,N_9759,N_8235);
and UO_240 (O_240,N_8098,N_8974);
and UO_241 (O_241,N_8861,N_9301);
nor UO_242 (O_242,N_8412,N_8168);
nand UO_243 (O_243,N_8067,N_9080);
and UO_244 (O_244,N_8050,N_9049);
nand UO_245 (O_245,N_8570,N_9261);
nand UO_246 (O_246,N_8395,N_9908);
nand UO_247 (O_247,N_9065,N_9685);
and UO_248 (O_248,N_9026,N_9204);
nor UO_249 (O_249,N_9245,N_8698);
and UO_250 (O_250,N_9191,N_9912);
or UO_251 (O_251,N_9290,N_9949);
nor UO_252 (O_252,N_8734,N_9637);
nor UO_253 (O_253,N_8220,N_8556);
nand UO_254 (O_254,N_8687,N_8829);
or UO_255 (O_255,N_8897,N_8767);
and UO_256 (O_256,N_9302,N_8400);
or UO_257 (O_257,N_9241,N_8612);
nand UO_258 (O_258,N_8927,N_9246);
xor UO_259 (O_259,N_9205,N_9862);
nand UO_260 (O_260,N_8607,N_9712);
and UO_261 (O_261,N_8135,N_9277);
nand UO_262 (O_262,N_9096,N_9770);
nand UO_263 (O_263,N_9792,N_8877);
or UO_264 (O_264,N_9567,N_9173);
nor UO_265 (O_265,N_9045,N_8347);
nor UO_266 (O_266,N_9846,N_9893);
and UO_267 (O_267,N_8563,N_9868);
or UO_268 (O_268,N_9950,N_9678);
and UO_269 (O_269,N_9154,N_9814);
and UO_270 (O_270,N_8470,N_8888);
or UO_271 (O_271,N_9729,N_9720);
nand UO_272 (O_272,N_8181,N_8437);
nor UO_273 (O_273,N_9686,N_8806);
nand UO_274 (O_274,N_8336,N_8215);
nor UO_275 (O_275,N_9063,N_8288);
or UO_276 (O_276,N_8988,N_8002);
nor UO_277 (O_277,N_9936,N_8046);
xor UO_278 (O_278,N_9351,N_9722);
and UO_279 (O_279,N_9343,N_8852);
and UO_280 (O_280,N_9786,N_9620);
or UO_281 (O_281,N_8326,N_9394);
and UO_282 (O_282,N_9061,N_8031);
or UO_283 (O_283,N_9337,N_8576);
or UO_284 (O_284,N_8847,N_8161);
nand UO_285 (O_285,N_8425,N_9521);
nand UO_286 (O_286,N_8064,N_8591);
and UO_287 (O_287,N_9053,N_8753);
nor UO_288 (O_288,N_8628,N_8203);
or UO_289 (O_289,N_8881,N_8582);
nand UO_290 (O_290,N_8605,N_8531);
nand UO_291 (O_291,N_8313,N_9150);
and UO_292 (O_292,N_9741,N_8789);
and UO_293 (O_293,N_8348,N_9183);
nor UO_294 (O_294,N_9450,N_8863);
nand UO_295 (O_295,N_9088,N_8294);
nand UO_296 (O_296,N_8808,N_9593);
nor UO_297 (O_297,N_9698,N_8104);
nand UO_298 (O_298,N_9886,N_9525);
nor UO_299 (O_299,N_9215,N_9682);
and UO_300 (O_300,N_8893,N_9929);
nand UO_301 (O_301,N_8912,N_8051);
nand UO_302 (O_302,N_9699,N_8972);
or UO_303 (O_303,N_8981,N_8644);
and UO_304 (O_304,N_8824,N_8188);
and UO_305 (O_305,N_8449,N_8597);
nand UO_306 (O_306,N_9687,N_8075);
nor UO_307 (O_307,N_8650,N_8287);
and UO_308 (O_308,N_8059,N_9464);
and UO_309 (O_309,N_8184,N_8198);
nor UO_310 (O_310,N_9651,N_8499);
or UO_311 (O_311,N_8647,N_9472);
nand UO_312 (O_312,N_8095,N_9135);
nor UO_313 (O_313,N_8160,N_9265);
and UO_314 (O_314,N_8831,N_9315);
and UO_315 (O_315,N_8733,N_8842);
and UO_316 (O_316,N_8121,N_8118);
or UO_317 (O_317,N_8334,N_9545);
nand UO_318 (O_318,N_9349,N_8351);
nor UO_319 (O_319,N_9445,N_9312);
and UO_320 (O_320,N_8111,N_9661);
nand UO_321 (O_321,N_9957,N_8341);
nor UO_322 (O_322,N_9035,N_8770);
and UO_323 (O_323,N_8946,N_8080);
or UO_324 (O_324,N_8534,N_8434);
nand UO_325 (O_325,N_8374,N_8213);
nor UO_326 (O_326,N_9305,N_9232);
or UO_327 (O_327,N_8190,N_9287);
or UO_328 (O_328,N_9543,N_8775);
or UO_329 (O_329,N_9850,N_8219);
nand UO_330 (O_330,N_8262,N_8872);
nand UO_331 (O_331,N_8099,N_8030);
nor UO_332 (O_332,N_8916,N_8291);
and UO_333 (O_333,N_9377,N_9257);
nand UO_334 (O_334,N_8833,N_8137);
nand UO_335 (O_335,N_8660,N_9976);
or UO_336 (O_336,N_9255,N_8544);
nand UO_337 (O_337,N_9182,N_9802);
nor UO_338 (O_338,N_9601,N_9573);
nand UO_339 (O_339,N_8955,N_8741);
and UO_340 (O_340,N_9826,N_8633);
or UO_341 (O_341,N_9763,N_8758);
or UO_342 (O_342,N_8816,N_9829);
and UO_343 (O_343,N_9509,N_8875);
and UO_344 (O_344,N_8510,N_9806);
nor UO_345 (O_345,N_9588,N_9253);
nand UO_346 (O_346,N_9689,N_9108);
nand UO_347 (O_347,N_8133,N_9311);
nand UO_348 (O_348,N_9925,N_8408);
nand UO_349 (O_349,N_9619,N_9374);
nor UO_350 (O_350,N_8516,N_9368);
nand UO_351 (O_351,N_8527,N_8041);
nor UO_352 (O_352,N_8432,N_9520);
nor UO_353 (O_353,N_8465,N_8202);
nand UO_354 (O_354,N_8638,N_9905);
or UO_355 (O_355,N_8092,N_8683);
and UO_356 (O_356,N_9798,N_8007);
or UO_357 (O_357,N_9228,N_9013);
or UO_358 (O_358,N_9591,N_9400);
nor UO_359 (O_359,N_9592,N_9998);
nand UO_360 (O_360,N_8076,N_8892);
nor UO_361 (O_361,N_8743,N_9410);
nor UO_362 (O_362,N_9816,N_8942);
and UO_363 (O_363,N_8044,N_8774);
nor UO_364 (O_364,N_9533,N_8837);
nand UO_365 (O_365,N_9990,N_9328);
nor UO_366 (O_366,N_9680,N_9158);
or UO_367 (O_367,N_9608,N_8406);
nor UO_368 (O_368,N_8969,N_8636);
and UO_369 (O_369,N_8484,N_8907);
and UO_370 (O_370,N_9830,N_8210);
nor UO_371 (O_371,N_9967,N_9075);
nand UO_372 (O_372,N_9402,N_9110);
nand UO_373 (O_373,N_9361,N_9740);
nand UO_374 (O_374,N_9364,N_8579);
and UO_375 (O_375,N_9579,N_8970);
and UO_376 (O_376,N_8297,N_8717);
nor UO_377 (O_377,N_8108,N_8079);
or UO_378 (O_378,N_9476,N_9985);
nor UO_379 (O_379,N_9440,N_9784);
or UO_380 (O_380,N_9742,N_8515);
nor UO_381 (O_381,N_8718,N_9782);
and UO_382 (O_382,N_9033,N_8885);
and UO_383 (O_383,N_8241,N_9866);
nand UO_384 (O_384,N_8540,N_9978);
nand UO_385 (O_385,N_9156,N_8000);
nor UO_386 (O_386,N_9892,N_8309);
nand UO_387 (O_387,N_9233,N_9020);
or UO_388 (O_388,N_8839,N_9347);
nand UO_389 (O_389,N_9781,N_8707);
and UO_390 (O_390,N_9112,N_8998);
nor UO_391 (O_391,N_9810,N_9580);
and UO_392 (O_392,N_8558,N_8921);
and UO_393 (O_393,N_9427,N_9165);
nor UO_394 (O_394,N_8207,N_8021);
or UO_395 (O_395,N_9704,N_9027);
nand UO_396 (O_396,N_9185,N_9751);
or UO_397 (O_397,N_9915,N_9731);
nor UO_398 (O_398,N_9992,N_8849);
and UO_399 (O_399,N_9805,N_8430);
or UO_400 (O_400,N_8732,N_8856);
or UO_401 (O_401,N_8211,N_8151);
nand UO_402 (O_402,N_9130,N_9016);
and UO_403 (O_403,N_9338,N_8407);
and UO_404 (O_404,N_9707,N_8176);
and UO_405 (O_405,N_9457,N_9393);
nor UO_406 (O_406,N_9861,N_9093);
and UO_407 (O_407,N_9744,N_8919);
nand UO_408 (O_408,N_9057,N_8155);
nor UO_409 (O_409,N_8372,N_9149);
nand UO_410 (O_410,N_8696,N_9865);
or UO_411 (O_411,N_9705,N_9789);
xor UO_412 (O_412,N_9431,N_8551);
nor UO_413 (O_413,N_8397,N_8016);
and UO_414 (O_414,N_8386,N_8772);
and UO_415 (O_415,N_8505,N_8367);
and UO_416 (O_416,N_9179,N_9227);
and UO_417 (O_417,N_9399,N_8314);
nor UO_418 (O_418,N_9598,N_8598);
or UO_419 (O_419,N_8205,N_9960);
nand UO_420 (O_420,N_8918,N_9360);
nand UO_421 (O_421,N_9681,N_9493);
and UO_422 (O_422,N_9403,N_8661);
and UO_423 (O_423,N_9748,N_9527);
nor UO_424 (O_424,N_9914,N_9951);
nor UO_425 (O_425,N_8366,N_9426);
and UO_426 (O_426,N_8521,N_9005);
nor UO_427 (O_427,N_9184,N_9254);
nand UO_428 (O_428,N_8245,N_9813);
nand UO_429 (O_429,N_8676,N_8379);
nand UO_430 (O_430,N_8296,N_9446);
nand UO_431 (O_431,N_9466,N_9605);
nor UO_432 (O_432,N_9869,N_8746);
nor UO_433 (O_433,N_8167,N_9935);
nand UO_434 (O_434,N_8280,N_9480);
nand UO_435 (O_435,N_8452,N_8617);
nand UO_436 (O_436,N_9743,N_9372);
nor UO_437 (O_437,N_9610,N_8131);
and UO_438 (O_438,N_9760,N_9120);
nor UO_439 (O_439,N_8781,N_9473);
nand UO_440 (O_440,N_8113,N_8862);
and UO_441 (O_441,N_8306,N_8047);
nand UO_442 (O_442,N_9279,N_9242);
and UO_443 (O_443,N_8910,N_8005);
nand UO_444 (O_444,N_8350,N_9894);
and UO_445 (O_445,N_8292,N_8090);
or UO_446 (O_446,N_8212,N_9197);
and UO_447 (O_447,N_8097,N_8900);
and UO_448 (O_448,N_9667,N_8524);
and UO_449 (O_449,N_8608,N_9656);
nand UO_450 (O_450,N_8738,N_9064);
or UO_451 (O_451,N_9123,N_9003);
nor UO_452 (O_452,N_8490,N_8442);
nor UO_453 (O_453,N_8265,N_9435);
and UO_454 (O_454,N_9418,N_9974);
or UO_455 (O_455,N_8268,N_8010);
and UO_456 (O_456,N_8014,N_9762);
nand UO_457 (O_457,N_8418,N_8782);
nor UO_458 (O_458,N_9456,N_8258);
nand UO_459 (O_459,N_9640,N_9222);
or UO_460 (O_460,N_8871,N_9837);
nor UO_461 (O_461,N_8684,N_8485);
or UO_462 (O_462,N_8225,N_9437);
nor UO_463 (O_463,N_9947,N_9036);
nor UO_464 (O_464,N_9102,N_8455);
and UO_465 (O_465,N_8230,N_8284);
or UO_466 (O_466,N_9725,N_9564);
and UO_467 (O_467,N_9210,N_9044);
nand UO_468 (O_468,N_8300,N_9398);
and UO_469 (O_469,N_8182,N_8073);
or UO_470 (O_470,N_9996,N_9470);
nand UO_471 (O_471,N_9519,N_8307);
and UO_472 (O_472,N_9008,N_9696);
nand UO_473 (O_473,N_8232,N_9136);
or UO_474 (O_474,N_9164,N_9326);
nor UO_475 (O_475,N_8670,N_8803);
nand UO_476 (O_476,N_9066,N_9911);
nor UO_477 (O_477,N_8441,N_9749);
and UO_478 (O_478,N_9657,N_8171);
nor UO_479 (O_479,N_9875,N_9654);
or UO_480 (O_480,N_8426,N_8275);
nor UO_481 (O_481,N_9993,N_9193);
or UO_482 (O_482,N_9941,N_8695);
and UO_483 (O_483,N_8724,N_8328);
or UO_484 (O_484,N_9478,N_9959);
or UO_485 (O_485,N_8604,N_9397);
nand UO_486 (O_486,N_9530,N_8312);
nor UO_487 (O_487,N_9055,N_9235);
nand UO_488 (O_488,N_8411,N_9652);
nor UO_489 (O_489,N_8261,N_8804);
nand UO_490 (O_490,N_8019,N_8009);
or UO_491 (O_491,N_8459,N_9040);
nor UO_492 (O_492,N_9702,N_8318);
or UO_493 (O_493,N_8085,N_8295);
nand UO_494 (O_494,N_8731,N_8987);
or UO_495 (O_495,N_8236,N_8107);
or UO_496 (O_496,N_9109,N_9552);
nand UO_497 (O_497,N_8932,N_9114);
and UO_498 (O_498,N_8323,N_8380);
nor UO_499 (O_499,N_8984,N_9733);
nor UO_500 (O_500,N_9980,N_8713);
nand UO_501 (O_501,N_9626,N_9152);
nor UO_502 (O_502,N_8637,N_9223);
or UO_503 (O_503,N_8122,N_8886);
nand UO_504 (O_504,N_9973,N_9979);
or UO_505 (O_505,N_8887,N_9052);
and UO_506 (O_506,N_9144,N_9604);
or UO_507 (O_507,N_9320,N_8533);
or UO_508 (O_508,N_8065,N_9845);
nor UO_509 (O_509,N_9775,N_9795);
or UO_510 (O_510,N_9887,N_8226);
nand UO_511 (O_511,N_8180,N_9294);
nand UO_512 (O_512,N_8788,N_9258);
or UO_513 (O_513,N_9458,N_8391);
or UO_514 (O_514,N_8587,N_8652);
nand UO_515 (O_515,N_9127,N_8869);
and UO_516 (O_516,N_9612,N_8196);
nand UO_517 (O_517,N_9313,N_8266);
and UO_518 (O_518,N_8785,N_9214);
and UO_519 (O_519,N_8941,N_8693);
nand UO_520 (O_520,N_9736,N_9989);
and UO_521 (O_521,N_8573,N_8433);
nor UO_522 (O_522,N_8750,N_8035);
or UO_523 (O_523,N_9528,N_8361);
nor UO_524 (O_524,N_8322,N_8519);
nor UO_525 (O_525,N_9060,N_8583);
nor UO_526 (O_526,N_9765,N_9438);
nor UO_527 (O_527,N_8389,N_8145);
nand UO_528 (O_528,N_8630,N_8310);
nor UO_529 (O_529,N_9636,N_8629);
and UO_530 (O_530,N_9790,N_8615);
nor UO_531 (O_531,N_9325,N_9903);
and UO_532 (O_532,N_9203,N_9703);
nor UO_533 (O_533,N_9001,N_8330);
nor UO_534 (O_534,N_8599,N_9176);
or UO_535 (O_535,N_9969,N_8973);
nand UO_536 (O_536,N_9961,N_9735);
and UO_537 (O_537,N_8939,N_8130);
and UO_538 (O_538,N_8281,N_9046);
and UO_539 (O_539,N_9839,N_9732);
nor UO_540 (O_540,N_8403,N_8752);
nor UO_541 (O_541,N_8078,N_9679);
and UO_542 (O_542,N_8349,N_9162);
nand UO_543 (O_543,N_8648,N_9014);
nor UO_544 (O_544,N_9570,N_9906);
nand UO_545 (O_545,N_8359,N_8469);
nor UO_546 (O_546,N_8508,N_9388);
and UO_547 (O_547,N_8263,N_9379);
and UO_548 (O_548,N_9880,N_8377);
nand UO_549 (O_549,N_9062,N_8846);
nand UO_550 (O_550,N_9536,N_9768);
and UO_551 (O_551,N_8884,N_8620);
nor UO_552 (O_552,N_9448,N_9469);
or UO_553 (O_553,N_8185,N_9838);
or UO_554 (O_554,N_8247,N_9126);
nand UO_555 (O_555,N_8012,N_8222);
nor UO_556 (O_556,N_9737,N_9863);
nand UO_557 (O_557,N_9991,N_8716);
nor UO_558 (O_558,N_9352,N_8048);
or UO_559 (O_559,N_8115,N_9964);
or UO_560 (O_560,N_8354,N_8124);
nor UO_561 (O_561,N_9451,N_9275);
or UO_562 (O_562,N_8257,N_9842);
nor UO_563 (O_563,N_8129,N_8776);
nand UO_564 (O_564,N_8224,N_8204);
or UO_565 (O_565,N_8506,N_8429);
nand UO_566 (O_566,N_9422,N_8553);
nor UO_567 (O_567,N_9094,N_9971);
or UO_568 (O_568,N_9803,N_8697);
nor UO_569 (O_569,N_8889,N_9688);
nor UO_570 (O_570,N_9583,N_9194);
nor UO_571 (O_571,N_9248,N_8904);
and UO_572 (O_572,N_8471,N_9141);
and UO_573 (O_573,N_9411,N_9207);
xnor UO_574 (O_574,N_8561,N_8201);
and UO_575 (O_575,N_8102,N_9077);
nor UO_576 (O_576,N_9252,N_8827);
nand UO_577 (O_577,N_9819,N_8272);
and UO_578 (O_578,N_9867,N_9496);
nor UO_579 (O_579,N_9444,N_9994);
and UO_580 (O_580,N_9664,N_8081);
or UO_581 (O_581,N_8466,N_8913);
nor UO_582 (O_582,N_9433,N_9549);
nand UO_583 (O_583,N_8055,N_9420);
or UO_584 (O_584,N_8339,N_9822);
nor UO_585 (O_585,N_9808,N_9820);
and UO_586 (O_586,N_9714,N_8911);
nor UO_587 (O_587,N_8762,N_9050);
and UO_588 (O_588,N_8303,N_9000);
nor UO_589 (O_589,N_9157,N_8358);
and UO_590 (O_590,N_9025,N_9069);
or UO_591 (O_591,N_9968,N_9498);
nand UO_592 (O_592,N_8362,N_9323);
and UO_593 (O_593,N_9081,N_9188);
nor UO_594 (O_594,N_8259,N_9369);
and UO_595 (O_595,N_9225,N_8209);
or UO_596 (O_596,N_8689,N_8654);
and UO_597 (O_597,N_9153,N_8878);
nand UO_598 (O_598,N_8504,N_8662);
and UO_599 (O_599,N_8825,N_9354);
nor UO_600 (O_600,N_9563,N_8218);
or UO_601 (O_601,N_8502,N_9631);
nand UO_602 (O_602,N_9717,N_9942);
or UO_603 (O_603,N_8568,N_9504);
nand UO_604 (O_604,N_8958,N_9357);
or UO_605 (O_605,N_8453,N_9091);
and UO_606 (O_606,N_9098,N_9890);
nand UO_607 (O_607,N_9791,N_8511);
and UO_608 (O_608,N_9220,N_8621);
nand UO_609 (O_609,N_8240,N_8768);
nor UO_610 (O_610,N_9874,N_8832);
or UO_611 (O_611,N_8902,N_9518);
nor UO_612 (O_612,N_8491,N_9777);
or UO_613 (O_613,N_9981,N_8764);
nor UO_614 (O_614,N_9212,N_9575);
nand UO_615 (O_615,N_8728,N_8575);
and UO_616 (O_616,N_9638,N_9585);
or UO_617 (O_617,N_8655,N_9943);
nor UO_618 (O_618,N_8873,N_8166);
nand UO_619 (O_619,N_9171,N_8834);
or UO_620 (O_620,N_9010,N_9577);
or UO_621 (O_621,N_9674,N_8156);
and UO_622 (O_622,N_8015,N_8779);
or UO_623 (O_623,N_8447,N_9271);
nand UO_624 (O_624,N_9556,N_9209);
nor UO_625 (O_625,N_9072,N_8062);
nand UO_626 (O_626,N_8112,N_9169);
and UO_627 (O_627,N_8070,N_8860);
and UO_628 (O_628,N_9481,N_9529);
nand UO_629 (O_629,N_8464,N_9266);
nand UO_630 (O_630,N_9769,N_8537);
and UO_631 (O_631,N_9928,N_8462);
nor UO_632 (O_632,N_9288,N_8143);
and UO_633 (O_633,N_8244,N_9948);
nand UO_634 (O_634,N_9897,N_8020);
or UO_635 (O_635,N_8995,N_8063);
and UO_636 (O_636,N_8777,N_8669);
nand UO_637 (O_637,N_9870,N_8027);
or UO_638 (O_638,N_9849,N_9774);
nand UO_639 (O_639,N_8054,N_8033);
nand UO_640 (O_640,N_8327,N_9206);
nor UO_641 (O_641,N_9024,N_8818);
and UO_642 (O_642,N_8331,N_9459);
nor UO_643 (O_643,N_9811,N_9256);
nand UO_644 (O_644,N_8634,N_8025);
nor UO_645 (O_645,N_9986,N_8836);
and UO_646 (O_646,N_8580,N_8091);
nor UO_647 (O_647,N_8951,N_8906);
and UO_648 (O_648,N_9772,N_9356);
and UO_649 (O_649,N_8659,N_8087);
or UO_650 (O_650,N_9558,N_9711);
and UO_651 (O_651,N_9611,N_8110);
or UO_652 (O_652,N_8905,N_8420);
nor UO_653 (O_653,N_8352,N_8948);
nand UO_654 (O_654,N_9362,N_8649);
nor UO_655 (O_655,N_8147,N_8454);
nand UO_656 (O_656,N_9787,N_9926);
and UO_657 (O_657,N_8721,N_9043);
and UO_658 (O_658,N_8664,N_9289);
and UO_659 (O_659,N_9627,N_8482);
or UO_660 (O_660,N_9174,N_9199);
or UO_661 (O_661,N_9296,N_9030);
nand UO_662 (O_662,N_8571,N_8158);
nor UO_663 (O_663,N_9505,N_8943);
and UO_664 (O_664,N_8479,N_9794);
or UO_665 (O_665,N_8177,N_8369);
or UO_666 (O_666,N_9380,N_9419);
nor UO_667 (O_667,N_9828,N_9281);
or UO_668 (O_668,N_9268,N_8840);
and UO_669 (O_669,N_8216,N_8477);
or UO_670 (O_670,N_9595,N_8017);
nand UO_671 (O_671,N_8214,N_8578);
or UO_672 (O_672,N_8703,N_8011);
or UO_673 (O_673,N_9734,N_9675);
nand UO_674 (O_674,N_8706,N_8925);
and UO_675 (O_675,N_8023,N_9780);
and UO_676 (O_676,N_8217,N_9375);
or UO_677 (O_677,N_9163,N_8963);
or UO_678 (O_678,N_8821,N_9750);
nand UO_679 (O_679,N_9417,N_8709);
and UO_680 (O_680,N_9694,N_9221);
nand UO_681 (O_681,N_9405,N_8584);
and UO_682 (O_682,N_8635,N_9727);
or UO_683 (O_683,N_9042,N_8039);
nand UO_684 (O_684,N_8826,N_9975);
and UO_685 (O_685,N_9202,N_9078);
or UO_686 (O_686,N_9160,N_9423);
nand UO_687 (O_687,N_8128,N_9310);
or UO_688 (O_688,N_9070,N_9345);
nor UO_689 (O_689,N_8965,N_8264);
nand UO_690 (O_690,N_8125,N_8843);
nor UO_691 (O_691,N_9267,N_8282);
or UO_692 (O_692,N_8154,N_9522);
and UO_693 (O_693,N_8293,N_9022);
or UO_694 (O_694,N_8727,N_9447);
nand UO_695 (O_695,N_8859,N_8609);
nor UO_696 (O_696,N_8536,N_8857);
and UO_697 (O_697,N_9507,N_9939);
and UO_698 (O_698,N_8394,N_8700);
nand UO_699 (O_699,N_8094,N_9872);
nor UO_700 (O_700,N_8152,N_8302);
nand UO_701 (O_701,N_9147,N_8363);
nor UO_702 (O_702,N_8542,N_8497);
and UO_703 (O_703,N_8159,N_9396);
or UO_704 (O_704,N_8186,N_9671);
nor UO_705 (O_705,N_9056,N_9779);
and UO_706 (O_706,N_9272,N_9616);
or UO_707 (O_707,N_9778,N_8277);
and UO_708 (O_708,N_8985,N_8711);
nand UO_709 (O_709,N_8117,N_9161);
xnor UO_710 (O_710,N_9339,N_9324);
and UO_711 (O_711,N_9240,N_9730);
and UO_712 (O_712,N_9208,N_9332);
or UO_713 (O_713,N_8345,N_8141);
or UO_714 (O_714,N_9004,N_9260);
xnor UO_715 (O_715,N_9015,N_9728);
and UO_716 (O_716,N_8618,N_8585);
nand UO_717 (O_717,N_8625,N_9853);
nor UO_718 (O_718,N_8392,N_8966);
and UO_719 (O_719,N_9666,N_8404);
nand UO_720 (O_720,N_8665,N_9319);
or UO_721 (O_721,N_9946,N_8566);
and UO_722 (O_722,N_9506,N_9247);
nand UO_723 (O_723,N_9889,N_9953);
nor UO_724 (O_724,N_8761,N_9840);
nor UO_725 (O_725,N_8968,N_9739);
or UO_726 (O_726,N_9095,N_8760);
or UO_727 (O_727,N_8541,N_8737);
or UO_728 (O_728,N_8867,N_9274);
nor UO_729 (O_729,N_9474,N_8431);
nand UO_730 (O_730,N_8451,N_8564);
or UO_731 (O_731,N_9700,N_8809);
and UO_732 (O_732,N_9392,N_8193);
or UO_733 (O_733,N_9237,N_8178);
and UO_734 (O_734,N_9511,N_9213);
nand UO_735 (O_735,N_9148,N_8123);
nand UO_736 (O_736,N_8172,N_9462);
or UO_737 (O_737,N_9539,N_8243);
or UO_738 (O_738,N_9531,N_8819);
and UO_739 (O_739,N_9482,N_8338);
or UO_740 (O_740,N_8964,N_9952);
nor UO_741 (O_741,N_8756,N_9956);
nor UO_742 (O_742,N_8278,N_9125);
or UO_743 (O_743,N_8084,N_9371);
and UO_744 (O_744,N_8378,N_8603);
nand UO_745 (O_745,N_9516,N_9408);
nand UO_746 (O_746,N_9834,N_8962);
nand UO_747 (O_747,N_9668,N_8068);
nor UO_748 (O_748,N_8109,N_9752);
nand UO_749 (O_749,N_8759,N_8855);
nand UO_750 (O_750,N_8924,N_8032);
or UO_751 (O_751,N_8472,N_8250);
or UO_752 (O_752,N_8344,N_8520);
nor UO_753 (O_753,N_8316,N_9586);
nand UO_754 (O_754,N_8438,N_8815);
or UO_755 (O_755,N_9477,N_9483);
or UO_756 (O_756,N_8200,N_9218);
nor UO_757 (O_757,N_8944,N_9977);
and UO_758 (O_758,N_9945,N_8298);
nand UO_759 (O_759,N_9382,N_9384);
nand UO_760 (O_760,N_8373,N_9047);
nand UO_761 (O_761,N_8866,N_9927);
and UO_762 (O_762,N_9079,N_9701);
or UO_763 (O_763,N_8624,N_9645);
nand UO_764 (O_764,N_9695,N_9934);
nand UO_765 (O_765,N_8658,N_8535);
nand UO_766 (O_766,N_8688,N_9658);
nor UO_767 (O_767,N_9559,N_8653);
nor UO_768 (O_768,N_9413,N_8643);
nor UO_769 (O_769,N_9589,N_8631);
nor UO_770 (O_770,N_8851,N_8901);
or UO_771 (O_771,N_8221,N_9293);
nand UO_772 (O_772,N_8543,N_9121);
nand UO_773 (O_773,N_8646,N_8848);
or UO_774 (O_774,N_8601,N_9270);
or UO_775 (O_775,N_9107,N_9641);
and UO_776 (O_776,N_9663,N_9684);
nand UO_777 (O_777,N_8461,N_9484);
nand UO_778 (O_778,N_8550,N_8089);
nand UO_779 (O_779,N_8467,N_8409);
nor UO_780 (O_780,N_8276,N_9922);
or UO_781 (O_781,N_9259,N_9486);
or UO_782 (O_782,N_9009,N_8006);
and UO_783 (O_783,N_8343,N_8191);
nor UO_784 (O_784,N_8745,N_9236);
and UO_785 (O_785,N_9367,N_8701);
nand UO_786 (O_786,N_9827,N_9757);
and UO_787 (O_787,N_9754,N_9219);
or UO_788 (O_788,N_9309,N_9623);
and UO_789 (O_789,N_8414,N_8763);
or UO_790 (O_790,N_9965,N_9172);
or UO_791 (O_791,N_9572,N_8895);
nand UO_792 (O_792,N_8034,N_8157);
and UO_793 (O_793,N_9333,N_8619);
nor UO_794 (O_794,N_8509,N_9363);
or UO_795 (O_795,N_8560,N_9282);
or UO_796 (O_796,N_8419,N_8725);
nor UO_797 (O_797,N_9799,N_9877);
nor UO_798 (O_798,N_8357,N_9851);
or UO_799 (O_799,N_9201,N_8627);
or UO_800 (O_800,N_8423,N_9344);
nor UO_801 (O_801,N_8383,N_8593);
and UO_802 (O_802,N_9489,N_9059);
nor UO_803 (O_803,N_9565,N_8446);
nand UO_804 (O_804,N_8088,N_8233);
or UO_805 (O_805,N_8952,N_9086);
nor UO_806 (O_806,N_8040,N_8399);
or UO_807 (O_807,N_9550,N_8254);
nor UO_808 (O_808,N_9378,N_8983);
nor UO_809 (O_809,N_8267,N_9415);
nor UO_810 (O_810,N_8489,N_8795);
and UO_811 (O_811,N_9177,N_8127);
and UO_812 (O_812,N_8468,N_8950);
or UO_813 (O_813,N_9920,N_9510);
or UO_814 (O_814,N_9503,N_9513);
nand UO_815 (O_815,N_9571,N_8056);
and UO_816 (O_816,N_9139,N_8114);
nand UO_817 (O_817,N_9537,N_8252);
nor UO_818 (O_818,N_8589,N_9783);
or UO_819 (O_819,N_8037,N_9262);
and UO_820 (O_820,N_8057,N_8251);
nor UO_821 (O_821,N_9944,N_9038);
or UO_822 (O_822,N_9963,N_8814);
or UO_823 (O_823,N_8917,N_8381);
nand UO_824 (O_824,N_8285,N_9436);
nand UO_825 (O_825,N_9443,N_8105);
and UO_826 (O_826,N_9800,N_8340);
nor UO_827 (O_827,N_9758,N_9962);
and UO_828 (O_828,N_8086,N_8606);
and UO_829 (O_829,N_8375,N_9600);
or UO_830 (O_830,N_8823,N_8165);
or UO_831 (O_831,N_8476,N_9414);
nor UO_832 (O_832,N_9843,N_8194);
and UO_833 (O_833,N_8682,N_9761);
nor UO_834 (O_834,N_8894,N_8822);
or UO_835 (O_835,N_9535,N_9871);
or UO_836 (O_836,N_9508,N_9074);
nor UO_837 (O_837,N_9497,N_9587);
nand UO_838 (O_838,N_8517,N_9560);
and UO_839 (O_839,N_9546,N_8581);
or UO_840 (O_840,N_9857,N_9713);
or UO_841 (O_841,N_9825,N_8817);
nor UO_842 (O_842,N_8083,N_9599);
nand UO_843 (O_843,N_8677,N_9676);
nor UO_844 (O_844,N_9719,N_9551);
nand UO_845 (O_845,N_9665,N_8061);
nor UO_846 (O_846,N_9355,N_9101);
and UO_847 (O_847,N_8492,N_9677);
nor UO_848 (O_848,N_8146,N_9048);
nor UO_849 (O_849,N_8940,N_9538);
nor UO_850 (O_850,N_9618,N_8530);
and UO_851 (O_851,N_8413,N_9807);
or UO_852 (O_852,N_8208,N_8242);
nor UO_853 (O_853,N_9021,N_8908);
and UO_854 (O_854,N_8071,N_9318);
and UO_855 (O_855,N_8013,N_9231);
and UO_856 (O_856,N_8947,N_8562);
nor UO_857 (O_857,N_9614,N_9297);
nor UO_858 (O_858,N_9723,N_8523);
or UO_859 (O_859,N_8810,N_8503);
nor UO_860 (O_860,N_9113,N_9821);
nor UO_861 (O_861,N_8594,N_8868);
nor UO_862 (O_862,N_9895,N_8456);
and UO_863 (O_863,N_9499,N_9439);
and UO_864 (O_864,N_9299,N_9211);
nand UO_865 (O_865,N_9848,N_8792);
nand UO_866 (O_866,N_9854,N_8610);
and UO_867 (O_867,N_8256,N_8148);
nand UO_868 (O_868,N_8742,N_8773);
nor UO_869 (O_869,N_9346,N_9747);
or UO_870 (O_870,N_8991,N_9119);
and UO_871 (O_871,N_8850,N_9251);
nor UO_872 (O_872,N_9292,N_8748);
or UO_873 (O_873,N_8956,N_9284);
nand UO_874 (O_874,N_8106,N_8546);
or UO_875 (O_875,N_8390,N_9738);
nor UO_876 (O_876,N_8666,N_8813);
and UO_877 (O_877,N_9494,N_8744);
or UO_878 (O_878,N_9690,N_8552);
and UO_879 (O_879,N_8674,N_8999);
nand UO_880 (O_880,N_9785,N_8103);
or UO_881 (O_881,N_9514,N_9649);
nor UO_882 (O_882,N_9832,N_9468);
and UO_883 (O_883,N_9632,N_8004);
nand UO_884 (O_884,N_9512,N_8854);
xor UO_885 (O_885,N_9195,N_8729);
and UO_886 (O_886,N_8270,N_8289);
nor UO_887 (O_887,N_9007,N_9833);
nor UO_888 (O_888,N_9249,N_9465);
or UO_889 (O_889,N_8173,N_8273);
or UO_890 (O_890,N_9793,N_8685);
nand UO_891 (O_891,N_9672,N_8977);
and UO_892 (O_892,N_8651,N_9891);
nor UO_893 (O_893,N_9597,N_9594);
nand UO_894 (O_894,N_9167,N_9391);
or UO_895 (O_895,N_8227,N_8771);
xnor UO_896 (O_896,N_9801,N_8790);
and UO_897 (O_897,N_8444,N_9430);
or UO_898 (O_898,N_8405,N_9348);
nand UO_899 (O_899,N_9475,N_9118);
and UO_900 (O_900,N_8149,N_8928);
and UO_901 (O_901,N_9381,N_9051);
nor UO_902 (O_902,N_8421,N_9073);
or UO_903 (O_903,N_8199,N_9502);
nand UO_904 (O_904,N_9138,N_9930);
and UO_905 (O_905,N_9099,N_8346);
and UO_906 (O_906,N_9940,N_9359);
or UO_907 (O_907,N_8838,N_9841);
and UO_908 (O_908,N_8876,N_9229);
nor UO_909 (O_909,N_8994,N_9490);
nor UO_910 (O_910,N_9628,N_9590);
nor UO_911 (O_911,N_9955,N_8260);
nor UO_912 (O_912,N_9017,N_8720);
or UO_913 (O_913,N_9907,N_8954);
xnor UO_914 (O_914,N_8645,N_9984);
nor UO_915 (O_915,N_9859,N_8060);
or UO_916 (O_916,N_8549,N_8008);
nand UO_917 (O_917,N_8714,N_9847);
nor UO_918 (O_918,N_9495,N_9314);
nand UO_919 (O_919,N_9970,N_9067);
and UO_920 (O_920,N_9921,N_9226);
or UO_921 (O_921,N_9122,N_8722);
nand UO_922 (O_922,N_8812,N_9273);
nor UO_923 (O_923,N_9140,N_8463);
and UO_924 (O_924,N_8841,N_9187);
and UO_925 (O_925,N_9291,N_8417);
nor UO_926 (O_926,N_8787,N_9650);
or UO_927 (O_927,N_8174,N_8990);
nand UO_928 (O_928,N_8641,N_8611);
nand UO_929 (O_929,N_9365,N_9131);
or UO_930 (O_930,N_9316,N_9966);
or UO_931 (O_931,N_8228,N_8518);
nor UO_932 (O_932,N_9836,N_9264);
nand UO_933 (O_933,N_8337,N_8691);
and UO_934 (O_934,N_8525,N_8730);
or UO_935 (O_935,N_9453,N_9917);
or UO_936 (O_936,N_9104,N_9910);
and UO_937 (O_937,N_8754,N_8957);
nand UO_938 (O_938,N_8715,N_9304);
and UO_939 (O_939,N_8356,N_8976);
and UO_940 (O_940,N_9166,N_8992);
and UO_941 (O_941,N_9856,N_8794);
or UO_942 (O_942,N_9353,N_8934);
nor UO_943 (O_943,N_9899,N_8360);
and UO_944 (O_944,N_9085,N_8526);
nand UO_945 (O_945,N_8569,N_8072);
or UO_946 (O_946,N_8317,N_9306);
nor UO_947 (O_947,N_8680,N_9896);
and UO_948 (O_948,N_8692,N_9151);
or UO_949 (O_949,N_8891,N_9032);
nand UO_950 (O_950,N_8304,N_9540);
or UO_951 (O_951,N_9425,N_8370);
or UO_952 (O_952,N_9517,N_8126);
or UO_953 (O_953,N_8493,N_9697);
nor UO_954 (O_954,N_8931,N_8702);
or UO_955 (O_955,N_9442,N_8082);
and UO_956 (O_956,N_9002,N_8539);
nand UO_957 (O_957,N_8673,N_8440);
nor UO_958 (O_958,N_9555,N_8269);
nor UO_959 (O_959,N_9693,N_8512);
or UO_960 (O_960,N_8163,N_9028);
nand UO_961 (O_961,N_9902,N_8996);
nand UO_962 (O_962,N_9129,N_8600);
nor UO_963 (O_963,N_8668,N_9500);
or UO_964 (O_964,N_8315,N_9106);
or UO_965 (O_965,N_8879,N_8398);
and UO_966 (O_966,N_9137,N_9858);
nand UO_967 (O_967,N_8043,N_9071);
nor UO_968 (O_968,N_8495,N_9330);
or UO_969 (O_969,N_9544,N_9170);
nand UO_970 (O_970,N_8874,N_8675);
nand UO_971 (O_971,N_8458,N_8882);
or UO_972 (O_972,N_9569,N_8053);
nor UO_973 (O_973,N_8719,N_9746);
or UO_974 (O_974,N_9180,N_8656);
nand UO_975 (O_975,N_8450,N_8058);
and UO_976 (O_976,N_9376,N_9660);
and UO_977 (O_977,N_8555,N_8332);
nand UO_978 (O_978,N_9766,N_8324);
nand UO_979 (O_979,N_8038,N_8959);
and UO_980 (O_980,N_9018,N_9485);
nand UO_981 (O_981,N_8162,N_9492);
nor UO_982 (O_982,N_9501,N_8747);
xor UO_983 (O_983,N_9280,N_9434);
or UO_984 (O_984,N_8765,N_9303);
and UO_985 (O_985,N_9553,N_8077);
and UO_986 (O_986,N_9395,N_8865);
or UO_987 (O_987,N_9884,N_9999);
nor UO_988 (O_988,N_9087,N_9898);
nor UO_989 (O_989,N_9416,N_9933);
or UO_990 (O_990,N_8140,N_9401);
nor UO_991 (O_991,N_8500,N_8473);
and UO_992 (O_992,N_8052,N_8507);
nor UO_993 (O_993,N_8557,N_9617);
nand UO_994 (O_994,N_9105,N_9449);
or UO_995 (O_995,N_8474,N_9643);
nand UO_996 (O_996,N_8705,N_8335);
or UO_997 (O_997,N_9479,N_9295);
nand UO_998 (O_998,N_9662,N_8001);
and UO_999 (O_999,N_8870,N_9029);
nor UO_1000 (O_1000,N_8813,N_8537);
nor UO_1001 (O_1001,N_9195,N_8260);
nor UO_1002 (O_1002,N_8516,N_9256);
nor UO_1003 (O_1003,N_8656,N_9004);
nand UO_1004 (O_1004,N_9867,N_8702);
nand UO_1005 (O_1005,N_8786,N_9373);
nand UO_1006 (O_1006,N_9123,N_8715);
nor UO_1007 (O_1007,N_9446,N_8720);
or UO_1008 (O_1008,N_9193,N_8816);
or UO_1009 (O_1009,N_9029,N_8233);
nor UO_1010 (O_1010,N_8777,N_8799);
or UO_1011 (O_1011,N_8155,N_9287);
nand UO_1012 (O_1012,N_8500,N_9735);
and UO_1013 (O_1013,N_8652,N_8288);
or UO_1014 (O_1014,N_8342,N_8593);
nand UO_1015 (O_1015,N_8756,N_9182);
or UO_1016 (O_1016,N_8225,N_8792);
and UO_1017 (O_1017,N_9578,N_8832);
or UO_1018 (O_1018,N_9020,N_8410);
nor UO_1019 (O_1019,N_9789,N_9622);
or UO_1020 (O_1020,N_9046,N_9897);
nand UO_1021 (O_1021,N_9734,N_8028);
nor UO_1022 (O_1022,N_8590,N_8522);
nand UO_1023 (O_1023,N_9624,N_9701);
nor UO_1024 (O_1024,N_8459,N_9626);
or UO_1025 (O_1025,N_9616,N_8943);
nand UO_1026 (O_1026,N_8398,N_8562);
or UO_1027 (O_1027,N_9421,N_8899);
and UO_1028 (O_1028,N_9341,N_8771);
or UO_1029 (O_1029,N_8129,N_9625);
nand UO_1030 (O_1030,N_9404,N_9887);
nand UO_1031 (O_1031,N_8936,N_9790);
nand UO_1032 (O_1032,N_8485,N_8472);
and UO_1033 (O_1033,N_9279,N_9574);
and UO_1034 (O_1034,N_9902,N_8849);
and UO_1035 (O_1035,N_9570,N_9149);
nand UO_1036 (O_1036,N_8356,N_9363);
and UO_1037 (O_1037,N_9303,N_9117);
and UO_1038 (O_1038,N_8311,N_9413);
nand UO_1039 (O_1039,N_8828,N_9755);
nor UO_1040 (O_1040,N_9288,N_9273);
nand UO_1041 (O_1041,N_9091,N_8452);
nor UO_1042 (O_1042,N_9092,N_8698);
nand UO_1043 (O_1043,N_9999,N_8629);
and UO_1044 (O_1044,N_8748,N_9739);
nand UO_1045 (O_1045,N_9062,N_9830);
and UO_1046 (O_1046,N_8313,N_8292);
or UO_1047 (O_1047,N_8364,N_9655);
nand UO_1048 (O_1048,N_9036,N_8847);
and UO_1049 (O_1049,N_8778,N_9148);
and UO_1050 (O_1050,N_8593,N_9136);
or UO_1051 (O_1051,N_8455,N_8509);
nand UO_1052 (O_1052,N_9373,N_9105);
or UO_1053 (O_1053,N_8798,N_8485);
nand UO_1054 (O_1054,N_8552,N_8356);
nand UO_1055 (O_1055,N_8333,N_9752);
or UO_1056 (O_1056,N_8363,N_8599);
nand UO_1057 (O_1057,N_8352,N_9340);
or UO_1058 (O_1058,N_9469,N_9087);
and UO_1059 (O_1059,N_9519,N_8535);
nand UO_1060 (O_1060,N_8546,N_8713);
nand UO_1061 (O_1061,N_9127,N_9424);
nor UO_1062 (O_1062,N_9869,N_8590);
and UO_1063 (O_1063,N_8224,N_9223);
or UO_1064 (O_1064,N_9521,N_9441);
nand UO_1065 (O_1065,N_9463,N_9215);
and UO_1066 (O_1066,N_8015,N_8316);
nor UO_1067 (O_1067,N_8995,N_9055);
nand UO_1068 (O_1068,N_8274,N_8278);
nand UO_1069 (O_1069,N_9468,N_8011);
or UO_1070 (O_1070,N_9749,N_8143);
or UO_1071 (O_1071,N_8228,N_8931);
and UO_1072 (O_1072,N_9330,N_9704);
and UO_1073 (O_1073,N_9020,N_8885);
or UO_1074 (O_1074,N_8855,N_9597);
or UO_1075 (O_1075,N_8582,N_8246);
nor UO_1076 (O_1076,N_8187,N_9063);
or UO_1077 (O_1077,N_8625,N_8755);
or UO_1078 (O_1078,N_9718,N_9445);
nand UO_1079 (O_1079,N_8769,N_8105);
nand UO_1080 (O_1080,N_9920,N_8335);
nor UO_1081 (O_1081,N_9389,N_8485);
xnor UO_1082 (O_1082,N_9217,N_8361);
and UO_1083 (O_1083,N_9731,N_9200);
or UO_1084 (O_1084,N_9753,N_8546);
or UO_1085 (O_1085,N_8694,N_9192);
or UO_1086 (O_1086,N_8440,N_9273);
or UO_1087 (O_1087,N_9381,N_8469);
nor UO_1088 (O_1088,N_8420,N_9642);
nor UO_1089 (O_1089,N_9595,N_9569);
or UO_1090 (O_1090,N_8824,N_9632);
and UO_1091 (O_1091,N_9504,N_8940);
or UO_1092 (O_1092,N_9970,N_9735);
and UO_1093 (O_1093,N_9191,N_8997);
or UO_1094 (O_1094,N_8956,N_8616);
nand UO_1095 (O_1095,N_9290,N_9325);
or UO_1096 (O_1096,N_8162,N_8000);
nand UO_1097 (O_1097,N_8609,N_9616);
nand UO_1098 (O_1098,N_9431,N_8474);
and UO_1099 (O_1099,N_9514,N_9551);
and UO_1100 (O_1100,N_9005,N_8963);
nor UO_1101 (O_1101,N_8961,N_8119);
or UO_1102 (O_1102,N_8100,N_9860);
or UO_1103 (O_1103,N_9247,N_9329);
nand UO_1104 (O_1104,N_9992,N_9331);
or UO_1105 (O_1105,N_9822,N_8189);
nand UO_1106 (O_1106,N_8719,N_9326);
nor UO_1107 (O_1107,N_8807,N_9645);
nor UO_1108 (O_1108,N_9056,N_8698);
and UO_1109 (O_1109,N_9051,N_9493);
or UO_1110 (O_1110,N_9073,N_8862);
nor UO_1111 (O_1111,N_9322,N_9388);
or UO_1112 (O_1112,N_9366,N_8979);
nor UO_1113 (O_1113,N_9491,N_9460);
and UO_1114 (O_1114,N_8311,N_9542);
or UO_1115 (O_1115,N_9338,N_9817);
or UO_1116 (O_1116,N_9166,N_9031);
or UO_1117 (O_1117,N_9994,N_8015);
or UO_1118 (O_1118,N_8184,N_9752);
nand UO_1119 (O_1119,N_9278,N_9067);
and UO_1120 (O_1120,N_8479,N_8795);
or UO_1121 (O_1121,N_9534,N_8181);
nor UO_1122 (O_1122,N_9113,N_8153);
nor UO_1123 (O_1123,N_9118,N_9709);
and UO_1124 (O_1124,N_8488,N_8097);
nor UO_1125 (O_1125,N_9696,N_9832);
or UO_1126 (O_1126,N_8368,N_8913);
nand UO_1127 (O_1127,N_9913,N_8611);
or UO_1128 (O_1128,N_8414,N_8295);
nor UO_1129 (O_1129,N_9404,N_8411);
or UO_1130 (O_1130,N_9997,N_9183);
nand UO_1131 (O_1131,N_8054,N_9478);
or UO_1132 (O_1132,N_9354,N_8112);
nor UO_1133 (O_1133,N_9158,N_8690);
nand UO_1134 (O_1134,N_8317,N_8435);
or UO_1135 (O_1135,N_9681,N_8650);
or UO_1136 (O_1136,N_8224,N_9753);
nand UO_1137 (O_1137,N_9676,N_9842);
nand UO_1138 (O_1138,N_9435,N_9965);
and UO_1139 (O_1139,N_9371,N_8393);
nand UO_1140 (O_1140,N_9676,N_8618);
and UO_1141 (O_1141,N_9350,N_9896);
nand UO_1142 (O_1142,N_8972,N_8049);
and UO_1143 (O_1143,N_8535,N_9003);
nor UO_1144 (O_1144,N_9290,N_9190);
nor UO_1145 (O_1145,N_9534,N_9770);
and UO_1146 (O_1146,N_9479,N_9377);
and UO_1147 (O_1147,N_8889,N_8727);
nor UO_1148 (O_1148,N_9740,N_8466);
nand UO_1149 (O_1149,N_9146,N_9311);
and UO_1150 (O_1150,N_9470,N_8230);
nand UO_1151 (O_1151,N_8429,N_9106);
nor UO_1152 (O_1152,N_8300,N_8474);
or UO_1153 (O_1153,N_9875,N_8307);
nand UO_1154 (O_1154,N_9802,N_9345);
nor UO_1155 (O_1155,N_8857,N_8459);
and UO_1156 (O_1156,N_8794,N_8938);
or UO_1157 (O_1157,N_9066,N_8456);
nand UO_1158 (O_1158,N_9649,N_9707);
nand UO_1159 (O_1159,N_8217,N_8727);
nand UO_1160 (O_1160,N_8847,N_8296);
nor UO_1161 (O_1161,N_9886,N_8953);
nor UO_1162 (O_1162,N_9178,N_9787);
and UO_1163 (O_1163,N_9397,N_8857);
and UO_1164 (O_1164,N_9380,N_9813);
nand UO_1165 (O_1165,N_8142,N_8348);
nand UO_1166 (O_1166,N_8218,N_9962);
or UO_1167 (O_1167,N_9526,N_9345);
nor UO_1168 (O_1168,N_9942,N_8163);
and UO_1169 (O_1169,N_8183,N_9733);
or UO_1170 (O_1170,N_9574,N_8623);
nor UO_1171 (O_1171,N_9952,N_9326);
nand UO_1172 (O_1172,N_8194,N_9826);
or UO_1173 (O_1173,N_9822,N_9273);
and UO_1174 (O_1174,N_9183,N_9110);
and UO_1175 (O_1175,N_9858,N_8112);
and UO_1176 (O_1176,N_9674,N_8281);
nand UO_1177 (O_1177,N_8888,N_8710);
nand UO_1178 (O_1178,N_8350,N_8882);
and UO_1179 (O_1179,N_8366,N_8463);
or UO_1180 (O_1180,N_8097,N_8093);
nand UO_1181 (O_1181,N_8982,N_9143);
and UO_1182 (O_1182,N_9705,N_9008);
xnor UO_1183 (O_1183,N_8592,N_8283);
and UO_1184 (O_1184,N_9485,N_9424);
or UO_1185 (O_1185,N_8187,N_8078);
and UO_1186 (O_1186,N_8320,N_9705);
nand UO_1187 (O_1187,N_9649,N_9162);
nor UO_1188 (O_1188,N_8747,N_8840);
and UO_1189 (O_1189,N_8803,N_9041);
nand UO_1190 (O_1190,N_9344,N_8516);
and UO_1191 (O_1191,N_8810,N_8626);
nand UO_1192 (O_1192,N_9137,N_8554);
or UO_1193 (O_1193,N_9699,N_8141);
or UO_1194 (O_1194,N_9728,N_8602);
nand UO_1195 (O_1195,N_8585,N_8284);
and UO_1196 (O_1196,N_9216,N_8543);
or UO_1197 (O_1197,N_9665,N_8663);
nand UO_1198 (O_1198,N_9627,N_8302);
nor UO_1199 (O_1199,N_9211,N_8194);
and UO_1200 (O_1200,N_9663,N_9362);
xor UO_1201 (O_1201,N_8056,N_9265);
and UO_1202 (O_1202,N_8239,N_8481);
and UO_1203 (O_1203,N_9527,N_9105);
or UO_1204 (O_1204,N_9963,N_9477);
nor UO_1205 (O_1205,N_8539,N_8509);
and UO_1206 (O_1206,N_8791,N_9395);
and UO_1207 (O_1207,N_8736,N_8999);
or UO_1208 (O_1208,N_9272,N_9262);
nor UO_1209 (O_1209,N_8027,N_8967);
or UO_1210 (O_1210,N_8800,N_9850);
nand UO_1211 (O_1211,N_8246,N_8776);
or UO_1212 (O_1212,N_9207,N_9855);
or UO_1213 (O_1213,N_8001,N_9418);
or UO_1214 (O_1214,N_8915,N_9246);
nand UO_1215 (O_1215,N_9656,N_8906);
nor UO_1216 (O_1216,N_8409,N_8898);
nor UO_1217 (O_1217,N_8652,N_9371);
nor UO_1218 (O_1218,N_8635,N_8901);
or UO_1219 (O_1219,N_8665,N_9061);
or UO_1220 (O_1220,N_9612,N_8246);
or UO_1221 (O_1221,N_8522,N_8303);
nand UO_1222 (O_1222,N_9746,N_9166);
nor UO_1223 (O_1223,N_9062,N_9455);
or UO_1224 (O_1224,N_9562,N_9993);
nor UO_1225 (O_1225,N_9449,N_9672);
nand UO_1226 (O_1226,N_9128,N_9463);
nand UO_1227 (O_1227,N_9011,N_8252);
and UO_1228 (O_1228,N_8045,N_8473);
nand UO_1229 (O_1229,N_9206,N_9634);
nor UO_1230 (O_1230,N_9307,N_9045);
nor UO_1231 (O_1231,N_9918,N_9830);
nor UO_1232 (O_1232,N_8283,N_8124);
nor UO_1233 (O_1233,N_8541,N_9212);
and UO_1234 (O_1234,N_9343,N_9546);
or UO_1235 (O_1235,N_9490,N_8063);
nor UO_1236 (O_1236,N_9555,N_8000);
nor UO_1237 (O_1237,N_9172,N_8735);
and UO_1238 (O_1238,N_9912,N_8465);
and UO_1239 (O_1239,N_9728,N_9378);
nor UO_1240 (O_1240,N_8931,N_9304);
or UO_1241 (O_1241,N_8062,N_9253);
nand UO_1242 (O_1242,N_8131,N_8124);
nand UO_1243 (O_1243,N_8739,N_8243);
and UO_1244 (O_1244,N_8403,N_9922);
and UO_1245 (O_1245,N_9970,N_8267);
and UO_1246 (O_1246,N_9903,N_9420);
nand UO_1247 (O_1247,N_8801,N_8536);
or UO_1248 (O_1248,N_8155,N_8855);
and UO_1249 (O_1249,N_9521,N_9246);
or UO_1250 (O_1250,N_9421,N_8479);
nor UO_1251 (O_1251,N_8498,N_9869);
or UO_1252 (O_1252,N_9644,N_8844);
and UO_1253 (O_1253,N_9296,N_9071);
nor UO_1254 (O_1254,N_9280,N_9632);
nand UO_1255 (O_1255,N_9413,N_8603);
nand UO_1256 (O_1256,N_9594,N_9122);
or UO_1257 (O_1257,N_9849,N_8800);
or UO_1258 (O_1258,N_8629,N_9693);
nor UO_1259 (O_1259,N_9789,N_9801);
or UO_1260 (O_1260,N_8185,N_9746);
or UO_1261 (O_1261,N_9515,N_9692);
or UO_1262 (O_1262,N_8277,N_8613);
nand UO_1263 (O_1263,N_9379,N_8589);
or UO_1264 (O_1264,N_9286,N_9668);
nand UO_1265 (O_1265,N_9105,N_9753);
nand UO_1266 (O_1266,N_8987,N_8365);
nor UO_1267 (O_1267,N_8118,N_9616);
nor UO_1268 (O_1268,N_9676,N_9521);
or UO_1269 (O_1269,N_8588,N_8891);
and UO_1270 (O_1270,N_9040,N_8483);
or UO_1271 (O_1271,N_8650,N_8043);
nor UO_1272 (O_1272,N_8291,N_8193);
or UO_1273 (O_1273,N_9690,N_9442);
nand UO_1274 (O_1274,N_8061,N_9965);
nand UO_1275 (O_1275,N_9773,N_9572);
nor UO_1276 (O_1276,N_8120,N_8379);
or UO_1277 (O_1277,N_8396,N_8379);
nand UO_1278 (O_1278,N_8692,N_9941);
or UO_1279 (O_1279,N_8910,N_8804);
and UO_1280 (O_1280,N_8447,N_9409);
and UO_1281 (O_1281,N_9325,N_8809);
or UO_1282 (O_1282,N_8601,N_9827);
nand UO_1283 (O_1283,N_8694,N_9139);
or UO_1284 (O_1284,N_8196,N_8166);
nor UO_1285 (O_1285,N_8991,N_8225);
nand UO_1286 (O_1286,N_9596,N_9345);
nor UO_1287 (O_1287,N_8184,N_9734);
and UO_1288 (O_1288,N_8395,N_8495);
or UO_1289 (O_1289,N_8063,N_9544);
nor UO_1290 (O_1290,N_8660,N_9388);
and UO_1291 (O_1291,N_8162,N_9830);
nor UO_1292 (O_1292,N_8002,N_9345);
and UO_1293 (O_1293,N_8508,N_8983);
or UO_1294 (O_1294,N_8280,N_8348);
and UO_1295 (O_1295,N_9469,N_9253);
nand UO_1296 (O_1296,N_9881,N_9044);
nor UO_1297 (O_1297,N_8745,N_9718);
nand UO_1298 (O_1298,N_9900,N_9855);
or UO_1299 (O_1299,N_8323,N_8447);
nand UO_1300 (O_1300,N_9836,N_8970);
and UO_1301 (O_1301,N_9489,N_8054);
and UO_1302 (O_1302,N_9406,N_9063);
nand UO_1303 (O_1303,N_8772,N_8535);
or UO_1304 (O_1304,N_8384,N_8254);
nand UO_1305 (O_1305,N_8326,N_9771);
or UO_1306 (O_1306,N_9041,N_9249);
and UO_1307 (O_1307,N_8606,N_9798);
or UO_1308 (O_1308,N_8534,N_8106);
nor UO_1309 (O_1309,N_8741,N_9433);
and UO_1310 (O_1310,N_8992,N_9948);
or UO_1311 (O_1311,N_8777,N_9742);
nand UO_1312 (O_1312,N_8587,N_9484);
nor UO_1313 (O_1313,N_8770,N_8069);
nor UO_1314 (O_1314,N_9766,N_9167);
nand UO_1315 (O_1315,N_9568,N_8026);
nor UO_1316 (O_1316,N_9049,N_8644);
nor UO_1317 (O_1317,N_9003,N_8241);
and UO_1318 (O_1318,N_9906,N_8075);
and UO_1319 (O_1319,N_8882,N_9708);
xor UO_1320 (O_1320,N_8023,N_8434);
and UO_1321 (O_1321,N_9642,N_9048);
or UO_1322 (O_1322,N_9477,N_9482);
and UO_1323 (O_1323,N_8746,N_9954);
nor UO_1324 (O_1324,N_9714,N_8775);
nand UO_1325 (O_1325,N_9186,N_9735);
and UO_1326 (O_1326,N_9106,N_8445);
or UO_1327 (O_1327,N_9851,N_9354);
nor UO_1328 (O_1328,N_8203,N_8909);
and UO_1329 (O_1329,N_8960,N_8681);
or UO_1330 (O_1330,N_9387,N_9742);
and UO_1331 (O_1331,N_9810,N_8694);
or UO_1332 (O_1332,N_9529,N_9988);
and UO_1333 (O_1333,N_8626,N_9913);
and UO_1334 (O_1334,N_8234,N_8204);
nor UO_1335 (O_1335,N_9893,N_8937);
nor UO_1336 (O_1336,N_9021,N_9417);
or UO_1337 (O_1337,N_8453,N_8692);
or UO_1338 (O_1338,N_8636,N_9924);
nor UO_1339 (O_1339,N_9694,N_9537);
nor UO_1340 (O_1340,N_8343,N_9699);
nor UO_1341 (O_1341,N_8290,N_9053);
or UO_1342 (O_1342,N_9359,N_9184);
nand UO_1343 (O_1343,N_8755,N_9951);
nor UO_1344 (O_1344,N_9516,N_8178);
nand UO_1345 (O_1345,N_9331,N_9881);
nand UO_1346 (O_1346,N_8461,N_9992);
and UO_1347 (O_1347,N_8722,N_9746);
nor UO_1348 (O_1348,N_8346,N_9451);
and UO_1349 (O_1349,N_9807,N_9464);
nand UO_1350 (O_1350,N_8542,N_9750);
and UO_1351 (O_1351,N_9811,N_8286);
nor UO_1352 (O_1352,N_8613,N_8712);
nor UO_1353 (O_1353,N_8025,N_9862);
nand UO_1354 (O_1354,N_9138,N_8495);
or UO_1355 (O_1355,N_8542,N_8169);
and UO_1356 (O_1356,N_9549,N_9365);
or UO_1357 (O_1357,N_8052,N_8604);
and UO_1358 (O_1358,N_9666,N_8401);
nand UO_1359 (O_1359,N_9775,N_9115);
and UO_1360 (O_1360,N_9356,N_9993);
and UO_1361 (O_1361,N_8120,N_8038);
or UO_1362 (O_1362,N_9404,N_9872);
nor UO_1363 (O_1363,N_8510,N_9411);
nor UO_1364 (O_1364,N_8214,N_8614);
nand UO_1365 (O_1365,N_8647,N_8920);
or UO_1366 (O_1366,N_8853,N_9747);
nand UO_1367 (O_1367,N_9293,N_9213);
and UO_1368 (O_1368,N_9370,N_9014);
nand UO_1369 (O_1369,N_9791,N_9506);
and UO_1370 (O_1370,N_9012,N_8138);
and UO_1371 (O_1371,N_9320,N_9605);
nand UO_1372 (O_1372,N_9691,N_9316);
or UO_1373 (O_1373,N_8896,N_8778);
nand UO_1374 (O_1374,N_9716,N_9510);
and UO_1375 (O_1375,N_8526,N_8167);
nor UO_1376 (O_1376,N_8245,N_9792);
and UO_1377 (O_1377,N_8859,N_8952);
and UO_1378 (O_1378,N_9149,N_9890);
or UO_1379 (O_1379,N_9702,N_8999);
nand UO_1380 (O_1380,N_8024,N_8490);
and UO_1381 (O_1381,N_9945,N_9081);
and UO_1382 (O_1382,N_9494,N_8996);
nand UO_1383 (O_1383,N_9375,N_8866);
or UO_1384 (O_1384,N_9602,N_8759);
nor UO_1385 (O_1385,N_8430,N_8577);
and UO_1386 (O_1386,N_8060,N_8586);
nor UO_1387 (O_1387,N_8462,N_8737);
and UO_1388 (O_1388,N_8206,N_9822);
xnor UO_1389 (O_1389,N_9265,N_9627);
or UO_1390 (O_1390,N_9356,N_8355);
nand UO_1391 (O_1391,N_8293,N_9904);
nor UO_1392 (O_1392,N_8550,N_9668);
or UO_1393 (O_1393,N_9739,N_9647);
nor UO_1394 (O_1394,N_9249,N_8125);
nand UO_1395 (O_1395,N_8406,N_8795);
and UO_1396 (O_1396,N_9735,N_8947);
nor UO_1397 (O_1397,N_9470,N_9258);
nand UO_1398 (O_1398,N_9612,N_9736);
and UO_1399 (O_1399,N_9669,N_8326);
or UO_1400 (O_1400,N_8727,N_9374);
xor UO_1401 (O_1401,N_8787,N_9472);
nand UO_1402 (O_1402,N_8002,N_9616);
or UO_1403 (O_1403,N_9843,N_8119);
and UO_1404 (O_1404,N_8483,N_8788);
nand UO_1405 (O_1405,N_9378,N_8357);
nand UO_1406 (O_1406,N_9293,N_9394);
or UO_1407 (O_1407,N_9165,N_8473);
nand UO_1408 (O_1408,N_8569,N_8477);
or UO_1409 (O_1409,N_8217,N_9547);
or UO_1410 (O_1410,N_8938,N_8916);
nand UO_1411 (O_1411,N_8754,N_9467);
nand UO_1412 (O_1412,N_8332,N_9006);
nor UO_1413 (O_1413,N_8226,N_9204);
nand UO_1414 (O_1414,N_9670,N_8303);
and UO_1415 (O_1415,N_9286,N_8730);
nand UO_1416 (O_1416,N_9805,N_8647);
nand UO_1417 (O_1417,N_9294,N_8405);
nand UO_1418 (O_1418,N_8696,N_9205);
nor UO_1419 (O_1419,N_8714,N_8767);
nand UO_1420 (O_1420,N_9652,N_8373);
nand UO_1421 (O_1421,N_8241,N_8502);
and UO_1422 (O_1422,N_8217,N_8920);
or UO_1423 (O_1423,N_9176,N_9705);
nor UO_1424 (O_1424,N_9019,N_8117);
or UO_1425 (O_1425,N_9104,N_9661);
nor UO_1426 (O_1426,N_8759,N_9311);
nor UO_1427 (O_1427,N_9644,N_8546);
nor UO_1428 (O_1428,N_9194,N_8463);
and UO_1429 (O_1429,N_8246,N_9253);
nand UO_1430 (O_1430,N_9632,N_9390);
nand UO_1431 (O_1431,N_8610,N_9372);
nand UO_1432 (O_1432,N_8711,N_9528);
and UO_1433 (O_1433,N_8856,N_9140);
and UO_1434 (O_1434,N_9427,N_8927);
or UO_1435 (O_1435,N_9212,N_9808);
and UO_1436 (O_1436,N_8265,N_9272);
nor UO_1437 (O_1437,N_9503,N_9701);
or UO_1438 (O_1438,N_9331,N_9702);
and UO_1439 (O_1439,N_8753,N_9893);
nor UO_1440 (O_1440,N_8723,N_9990);
nand UO_1441 (O_1441,N_8590,N_9224);
nand UO_1442 (O_1442,N_9248,N_9796);
and UO_1443 (O_1443,N_8621,N_9665);
nand UO_1444 (O_1444,N_8575,N_8335);
nor UO_1445 (O_1445,N_8649,N_9492);
nor UO_1446 (O_1446,N_8992,N_8249);
nand UO_1447 (O_1447,N_9780,N_9606);
nor UO_1448 (O_1448,N_9764,N_9654);
nand UO_1449 (O_1449,N_9767,N_8149);
nor UO_1450 (O_1450,N_8902,N_8365);
nand UO_1451 (O_1451,N_9482,N_9581);
nand UO_1452 (O_1452,N_8611,N_9995);
nor UO_1453 (O_1453,N_8073,N_8705);
nor UO_1454 (O_1454,N_8589,N_8190);
nor UO_1455 (O_1455,N_9138,N_9054);
nand UO_1456 (O_1456,N_9661,N_9483);
nor UO_1457 (O_1457,N_9733,N_8694);
and UO_1458 (O_1458,N_9779,N_9416);
or UO_1459 (O_1459,N_9367,N_8037);
and UO_1460 (O_1460,N_8738,N_8009);
or UO_1461 (O_1461,N_8436,N_8325);
nand UO_1462 (O_1462,N_9519,N_8631);
and UO_1463 (O_1463,N_9496,N_8201);
and UO_1464 (O_1464,N_9991,N_8081);
nand UO_1465 (O_1465,N_8170,N_9208);
and UO_1466 (O_1466,N_9368,N_9791);
and UO_1467 (O_1467,N_8711,N_8769);
nand UO_1468 (O_1468,N_8118,N_9400);
nand UO_1469 (O_1469,N_8727,N_9065);
nand UO_1470 (O_1470,N_8009,N_8395);
and UO_1471 (O_1471,N_9171,N_8450);
or UO_1472 (O_1472,N_8569,N_9970);
nor UO_1473 (O_1473,N_8595,N_8991);
nand UO_1474 (O_1474,N_8935,N_9890);
and UO_1475 (O_1475,N_9102,N_9230);
nand UO_1476 (O_1476,N_9840,N_9005);
nand UO_1477 (O_1477,N_8688,N_8271);
or UO_1478 (O_1478,N_8985,N_8273);
or UO_1479 (O_1479,N_8109,N_9932);
nand UO_1480 (O_1480,N_8827,N_9802);
and UO_1481 (O_1481,N_9691,N_8977);
and UO_1482 (O_1482,N_8312,N_8081);
and UO_1483 (O_1483,N_9558,N_8745);
or UO_1484 (O_1484,N_8745,N_8035);
or UO_1485 (O_1485,N_8661,N_9813);
xor UO_1486 (O_1486,N_9098,N_8601);
nand UO_1487 (O_1487,N_8685,N_8299);
nand UO_1488 (O_1488,N_8158,N_8959);
or UO_1489 (O_1489,N_8483,N_9525);
or UO_1490 (O_1490,N_9903,N_9453);
nand UO_1491 (O_1491,N_8626,N_8522);
or UO_1492 (O_1492,N_9952,N_9611);
or UO_1493 (O_1493,N_8803,N_9826);
and UO_1494 (O_1494,N_9269,N_8805);
nand UO_1495 (O_1495,N_9226,N_9704);
or UO_1496 (O_1496,N_9426,N_8667);
nor UO_1497 (O_1497,N_8006,N_8985);
nand UO_1498 (O_1498,N_8871,N_8486);
nand UO_1499 (O_1499,N_9531,N_8875);
endmodule