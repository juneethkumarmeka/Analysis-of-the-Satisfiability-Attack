module basic_500_3000_500_15_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_21,In_396);
nor U1 (N_1,In_297,In_270);
nand U2 (N_2,In_435,In_97);
nand U3 (N_3,In_43,In_398);
or U4 (N_4,In_261,In_351);
nor U5 (N_5,In_402,In_285);
and U6 (N_6,In_315,In_366);
or U7 (N_7,In_240,In_277);
or U8 (N_8,In_168,In_30);
and U9 (N_9,In_9,In_459);
nor U10 (N_10,In_468,In_188);
or U11 (N_11,In_385,In_195);
and U12 (N_12,In_37,In_72);
and U13 (N_13,In_289,In_146);
nor U14 (N_14,In_492,In_498);
or U15 (N_15,In_104,In_122);
and U16 (N_16,In_99,In_475);
nand U17 (N_17,In_437,In_292);
or U18 (N_18,In_455,In_25);
and U19 (N_19,In_324,In_451);
and U20 (N_20,In_28,In_323);
nor U21 (N_21,In_346,In_259);
nand U22 (N_22,In_153,In_87);
or U23 (N_23,In_6,In_51);
and U24 (N_24,In_283,In_453);
xor U25 (N_25,In_284,In_372);
and U26 (N_26,In_441,In_477);
nand U27 (N_27,In_249,In_295);
or U28 (N_28,In_290,In_313);
nand U29 (N_29,In_410,In_52);
and U30 (N_30,In_348,In_312);
nor U31 (N_31,In_35,In_219);
or U32 (N_32,In_210,In_144);
or U33 (N_33,In_326,In_182);
or U34 (N_34,In_361,In_258);
nor U35 (N_35,In_349,In_68);
or U36 (N_36,In_484,In_470);
or U37 (N_37,In_273,In_243);
or U38 (N_38,In_14,In_76);
xor U39 (N_39,In_169,In_389);
nor U40 (N_40,In_424,In_34);
or U41 (N_41,In_159,In_449);
nand U42 (N_42,In_208,In_364);
nand U43 (N_43,In_119,In_16);
and U44 (N_44,In_73,In_335);
xor U45 (N_45,In_417,In_151);
or U46 (N_46,In_124,In_338);
nor U47 (N_47,In_170,In_408);
nor U48 (N_48,In_90,In_46);
nand U49 (N_49,In_67,In_118);
and U50 (N_50,In_352,In_345);
nor U51 (N_51,In_264,In_212);
and U52 (N_52,In_379,In_71);
nor U53 (N_53,In_452,In_306);
or U54 (N_54,In_458,In_232);
or U55 (N_55,In_370,In_29);
or U56 (N_56,In_216,In_185);
nand U57 (N_57,In_127,In_95);
nor U58 (N_58,In_155,In_248);
nor U59 (N_59,In_101,In_450);
and U60 (N_60,In_462,In_448);
and U61 (N_61,In_89,In_412);
nand U62 (N_62,In_461,In_1);
nor U63 (N_63,In_332,In_262);
and U64 (N_64,In_365,In_150);
nand U65 (N_65,In_291,In_12);
or U66 (N_66,In_91,In_422);
nand U67 (N_67,In_478,In_126);
nor U68 (N_68,In_180,In_282);
nand U69 (N_69,In_84,In_486);
nand U70 (N_70,In_5,In_110);
nand U71 (N_71,In_148,In_142);
or U72 (N_72,In_154,In_111);
and U73 (N_73,In_79,In_54);
or U74 (N_74,In_114,In_303);
and U75 (N_75,In_265,In_247);
nor U76 (N_76,In_483,In_328);
or U77 (N_77,In_239,In_56);
nand U78 (N_78,In_339,In_171);
or U79 (N_79,In_260,In_405);
nor U80 (N_80,In_438,In_304);
or U81 (N_81,In_288,In_128);
or U82 (N_82,In_436,In_309);
nor U83 (N_83,In_369,In_255);
nand U84 (N_84,In_416,In_471);
and U85 (N_85,In_112,In_428);
nor U86 (N_86,In_152,In_480);
and U87 (N_87,In_414,In_238);
and U88 (N_88,In_399,In_341);
and U89 (N_89,In_74,In_161);
nand U90 (N_90,In_359,In_447);
nor U91 (N_91,In_77,In_286);
nand U92 (N_92,In_93,In_454);
nor U93 (N_93,In_141,In_116);
nand U94 (N_94,In_225,In_164);
and U95 (N_95,In_465,In_439);
nand U96 (N_96,In_57,In_446);
or U97 (N_97,In_443,In_373);
or U98 (N_98,In_157,In_226);
and U99 (N_99,In_163,In_469);
or U100 (N_100,In_299,In_65);
nand U101 (N_101,In_125,In_251);
and U102 (N_102,In_136,In_497);
nor U103 (N_103,In_493,In_460);
nor U104 (N_104,In_482,In_98);
or U105 (N_105,In_204,In_381);
nor U106 (N_106,In_472,In_392);
or U107 (N_107,In_367,In_172);
nor U108 (N_108,In_429,In_7);
nor U109 (N_109,In_203,In_213);
nor U110 (N_110,In_8,In_268);
and U111 (N_111,In_318,In_222);
or U112 (N_112,In_69,In_401);
and U113 (N_113,In_147,In_134);
and U114 (N_114,In_106,In_187);
nand U115 (N_115,In_131,In_227);
or U116 (N_116,In_194,In_426);
or U117 (N_117,In_193,In_357);
and U118 (N_118,In_209,In_235);
nand U119 (N_119,In_186,In_221);
and U120 (N_120,In_19,In_121);
nor U121 (N_121,In_63,In_44);
xor U122 (N_122,In_167,In_388);
nand U123 (N_123,In_409,In_61);
xnor U124 (N_124,In_275,In_181);
nor U125 (N_125,In_499,In_330);
nand U126 (N_126,In_189,In_397);
nor U127 (N_127,In_109,In_229);
nor U128 (N_128,In_241,In_419);
or U129 (N_129,In_53,In_390);
or U130 (N_130,In_246,In_430);
and U131 (N_131,In_266,In_256);
nand U132 (N_132,In_343,In_257);
nor U133 (N_133,In_192,In_269);
or U134 (N_134,In_415,In_179);
nand U135 (N_135,In_10,In_380);
xor U136 (N_136,In_433,In_231);
nor U137 (N_137,In_327,In_94);
nor U138 (N_138,In_431,In_383);
or U139 (N_139,In_418,In_342);
nand U140 (N_140,In_376,In_245);
and U141 (N_141,In_120,In_133);
and U142 (N_142,In_336,In_4);
nor U143 (N_143,In_220,In_78);
nand U144 (N_144,In_325,In_233);
nor U145 (N_145,In_23,In_50);
and U146 (N_146,In_496,In_82);
nand U147 (N_147,In_344,In_407);
and U148 (N_148,In_242,In_384);
or U149 (N_149,In_363,In_374);
nand U150 (N_150,In_276,In_442);
nor U151 (N_151,In_22,In_317);
nand U152 (N_152,In_314,In_293);
xor U153 (N_153,In_107,In_413);
and U154 (N_154,In_244,In_355);
nand U155 (N_155,In_39,In_196);
or U156 (N_156,In_178,In_113);
nor U157 (N_157,In_27,In_26);
nor U158 (N_158,In_271,In_20);
and U159 (N_159,In_234,In_400);
and U160 (N_160,In_250,In_137);
nand U161 (N_161,In_377,In_337);
xnor U162 (N_162,In_404,In_356);
nand U163 (N_163,In_81,In_387);
nand U164 (N_164,In_253,In_481);
or U165 (N_165,In_165,In_183);
and U166 (N_166,In_427,In_375);
and U167 (N_167,In_228,In_139);
or U168 (N_168,In_279,In_130);
and U169 (N_169,In_103,In_162);
or U170 (N_170,In_202,In_135);
or U171 (N_171,In_300,In_393);
nand U172 (N_172,In_100,In_92);
nand U173 (N_173,In_15,In_96);
nand U174 (N_174,In_190,In_287);
and U175 (N_175,In_411,In_218);
nand U176 (N_176,In_425,In_47);
nor U177 (N_177,In_174,In_80);
nor U178 (N_178,In_310,In_13);
nand U179 (N_179,In_457,In_340);
or U180 (N_180,In_173,In_490);
or U181 (N_181,In_421,In_254);
nand U182 (N_182,In_440,In_205);
nor U183 (N_183,In_32,In_354);
nor U184 (N_184,In_444,In_214);
nor U185 (N_185,In_191,In_463);
and U186 (N_186,In_322,In_143);
nor U187 (N_187,In_487,In_347);
or U188 (N_188,In_382,In_156);
nand U189 (N_189,In_358,In_467);
nand U190 (N_190,In_108,In_115);
and U191 (N_191,In_434,In_302);
or U192 (N_192,In_488,In_368);
nor U193 (N_193,In_224,In_184);
nand U194 (N_194,In_31,In_237);
or U195 (N_195,In_305,In_298);
or U196 (N_196,In_296,In_223);
nor U197 (N_197,In_105,In_489);
and U198 (N_198,In_132,In_17);
and U199 (N_199,In_70,In_272);
or U200 (N_200,N_15,In_175);
and U201 (N_201,N_167,N_108);
and U202 (N_202,N_104,N_128);
nor U203 (N_203,N_26,N_90);
nor U204 (N_204,N_74,In_38);
nor U205 (N_205,In_406,N_193);
nor U206 (N_206,N_134,N_160);
or U207 (N_207,N_184,N_157);
nor U208 (N_208,N_51,In_329);
and U209 (N_209,N_119,In_420);
nor U210 (N_210,N_140,N_66);
or U211 (N_211,In_308,N_54);
nor U212 (N_212,N_122,N_99);
nor U213 (N_213,N_35,N_114);
or U214 (N_214,In_360,N_52);
nor U215 (N_215,In_40,In_267);
or U216 (N_216,N_153,N_73);
and U217 (N_217,N_97,In_177);
nand U218 (N_218,N_154,In_394);
or U219 (N_219,In_350,In_476);
and U220 (N_220,N_3,In_252);
and U221 (N_221,In_371,N_22);
or U222 (N_222,In_386,N_100);
or U223 (N_223,In_211,N_48);
or U224 (N_224,In_55,In_274);
nor U225 (N_225,In_2,N_111);
and U226 (N_226,N_64,In_311);
and U227 (N_227,N_103,N_162);
and U228 (N_228,N_101,N_170);
or U229 (N_229,N_40,N_163);
or U230 (N_230,In_198,N_152);
nand U231 (N_231,In_41,N_6);
xor U232 (N_232,In_86,N_199);
or U233 (N_233,N_20,N_164);
nor U234 (N_234,N_24,N_25);
nor U235 (N_235,N_8,N_41);
or U236 (N_236,N_180,N_4);
nand U237 (N_237,N_185,In_117);
nor U238 (N_238,N_196,N_145);
nand U239 (N_239,N_9,N_197);
nand U240 (N_240,N_106,N_188);
or U241 (N_241,N_43,N_85);
or U242 (N_242,In_319,In_160);
nand U243 (N_243,N_171,N_34);
or U244 (N_244,In_176,N_33);
or U245 (N_245,In_464,N_65);
nor U246 (N_246,N_146,N_189);
or U247 (N_247,N_50,N_137);
nor U248 (N_248,N_95,N_27);
nand U249 (N_249,N_53,In_200);
and U250 (N_250,N_29,N_182);
nor U251 (N_251,In_432,N_38);
nor U252 (N_252,N_174,N_39);
nor U253 (N_253,N_102,N_7);
and U254 (N_254,N_172,In_199);
and U255 (N_255,N_138,In_145);
xor U256 (N_256,N_118,In_333);
nand U257 (N_257,N_112,N_135);
and U258 (N_258,N_136,N_142);
nor U259 (N_259,In_485,N_71);
nand U260 (N_260,N_28,N_126);
or U261 (N_261,N_63,In_280);
and U262 (N_262,N_23,N_32);
and U263 (N_263,In_321,N_195);
nand U264 (N_264,N_123,N_79);
and U265 (N_265,In_391,N_30);
or U266 (N_266,N_91,In_85);
and U267 (N_267,N_84,N_31);
nand U268 (N_268,In_445,N_143);
or U269 (N_269,In_378,In_24);
nor U270 (N_270,N_49,N_16);
or U271 (N_271,In_158,N_5);
or U272 (N_272,N_67,N_82);
nand U273 (N_273,In_66,In_201);
and U274 (N_274,In_11,N_47);
and U275 (N_275,N_61,N_125);
nor U276 (N_276,N_80,N_62);
nand U277 (N_277,N_173,N_113);
and U278 (N_278,In_362,N_149);
nand U279 (N_279,N_155,In_149);
nor U280 (N_280,In_395,N_141);
or U281 (N_281,N_161,N_148);
and U282 (N_282,N_192,In_217);
and U283 (N_283,N_186,N_19);
and U284 (N_284,In_316,N_198);
or U285 (N_285,In_301,N_77);
nand U286 (N_286,N_131,N_55);
nand U287 (N_287,N_169,N_46);
nand U288 (N_288,N_133,N_87);
or U289 (N_289,In_18,In_281);
or U290 (N_290,N_92,N_165);
or U291 (N_291,N_57,In_215);
and U292 (N_292,In_474,In_60);
and U293 (N_293,In_263,N_86);
and U294 (N_294,N_18,N_88);
and U295 (N_295,N_132,N_2);
nor U296 (N_296,N_56,N_127);
nor U297 (N_297,N_0,In_138);
nand U298 (N_298,N_181,N_81);
nand U299 (N_299,In_331,N_14);
nand U300 (N_300,In_88,N_11);
nor U301 (N_301,N_107,N_98);
nor U302 (N_302,In_278,N_176);
nor U303 (N_303,In_166,N_89);
and U304 (N_304,In_479,In_320);
or U305 (N_305,N_121,In_230);
nand U306 (N_306,N_58,In_59);
and U307 (N_307,N_194,N_156);
or U308 (N_308,N_179,In_495);
nor U309 (N_309,N_120,In_140);
and U310 (N_310,N_110,N_183);
or U311 (N_311,N_96,N_168);
nand U312 (N_312,In_466,N_191);
nand U313 (N_313,In_123,N_37);
and U314 (N_314,In_64,N_60);
or U315 (N_315,N_68,In_294);
or U316 (N_316,N_109,N_76);
or U317 (N_317,N_10,In_75);
or U318 (N_318,N_69,N_59);
and U319 (N_319,In_3,N_21);
nand U320 (N_320,In_45,N_93);
and U321 (N_321,In_42,In_48);
nor U322 (N_322,N_75,In_102);
and U323 (N_323,In_62,In_353);
nand U324 (N_324,N_177,In_36);
and U325 (N_325,In_403,N_175);
nand U326 (N_326,N_151,In_83);
nand U327 (N_327,N_166,N_124);
or U328 (N_328,N_187,N_12);
or U329 (N_329,In_58,In_236);
or U330 (N_330,N_158,In_307);
and U331 (N_331,N_139,In_207);
and U332 (N_332,In_456,N_72);
and U333 (N_333,N_44,N_36);
and U334 (N_334,N_129,In_129);
nand U335 (N_335,N_105,In_494);
or U336 (N_336,N_83,N_78);
and U337 (N_337,N_147,N_178);
and U338 (N_338,In_334,N_190);
and U339 (N_339,N_1,N_70);
and U340 (N_340,N_17,N_150);
nor U341 (N_341,In_423,N_45);
or U342 (N_342,In_197,In_206);
or U343 (N_343,N_42,In_33);
nand U344 (N_344,In_473,N_130);
xnor U345 (N_345,N_116,In_0);
and U346 (N_346,N_117,N_144);
nand U347 (N_347,N_13,In_49);
and U348 (N_348,In_491,N_115);
nand U349 (N_349,N_94,N_159);
nand U350 (N_350,N_127,N_162);
xor U351 (N_351,N_173,In_11);
or U352 (N_352,N_115,N_108);
and U353 (N_353,N_132,N_72);
nor U354 (N_354,N_33,In_494);
and U355 (N_355,N_100,N_141);
nand U356 (N_356,N_44,N_51);
nor U357 (N_357,N_70,N_111);
and U358 (N_358,In_117,N_138);
or U359 (N_359,N_125,N_96);
nor U360 (N_360,N_80,In_334);
nor U361 (N_361,N_139,N_162);
nor U362 (N_362,In_211,In_75);
and U363 (N_363,In_491,In_267);
nor U364 (N_364,N_112,N_77);
nor U365 (N_365,N_12,N_7);
or U366 (N_366,N_54,In_485);
or U367 (N_367,N_93,N_163);
nand U368 (N_368,N_16,N_130);
nor U369 (N_369,N_101,N_32);
and U370 (N_370,N_122,In_177);
nor U371 (N_371,In_432,N_115);
xnor U372 (N_372,N_93,In_42);
nand U373 (N_373,In_491,In_40);
nor U374 (N_374,In_86,N_95);
nor U375 (N_375,N_8,N_116);
nor U376 (N_376,N_134,In_395);
and U377 (N_377,N_73,N_157);
nor U378 (N_378,N_9,N_188);
or U379 (N_379,N_51,In_215);
nand U380 (N_380,N_97,N_143);
nand U381 (N_381,In_476,In_311);
xnor U382 (N_382,In_66,N_65);
or U383 (N_383,N_170,N_120);
nor U384 (N_384,N_131,In_307);
or U385 (N_385,N_86,N_91);
nor U386 (N_386,In_145,N_158);
and U387 (N_387,N_130,N_152);
and U388 (N_388,In_474,In_316);
and U389 (N_389,In_479,N_29);
and U390 (N_390,In_123,N_47);
and U391 (N_391,In_473,In_294);
or U392 (N_392,In_123,N_49);
nor U393 (N_393,N_85,In_88);
nand U394 (N_394,N_162,N_144);
nor U395 (N_395,N_60,N_87);
xnor U396 (N_396,In_456,N_169);
nor U397 (N_397,N_165,In_206);
nor U398 (N_398,In_18,N_89);
nor U399 (N_399,In_55,In_0);
or U400 (N_400,N_303,N_202);
nand U401 (N_401,N_356,N_214);
nor U402 (N_402,N_355,N_353);
or U403 (N_403,N_359,N_322);
nor U404 (N_404,N_235,N_250);
and U405 (N_405,N_247,N_251);
nor U406 (N_406,N_352,N_278);
or U407 (N_407,N_351,N_215);
nor U408 (N_408,N_369,N_349);
or U409 (N_409,N_286,N_365);
xnor U410 (N_410,N_336,N_208);
and U411 (N_411,N_234,N_261);
or U412 (N_412,N_258,N_361);
nand U413 (N_413,N_209,N_375);
and U414 (N_414,N_330,N_255);
nand U415 (N_415,N_344,N_378);
and U416 (N_416,N_331,N_296);
or U417 (N_417,N_343,N_253);
and U418 (N_418,N_364,N_212);
and U419 (N_419,N_300,N_268);
nor U420 (N_420,N_285,N_233);
or U421 (N_421,N_216,N_370);
xor U422 (N_422,N_210,N_313);
or U423 (N_423,N_318,N_211);
nor U424 (N_424,N_305,N_223);
nand U425 (N_425,N_382,N_307);
nor U426 (N_426,N_267,N_315);
and U427 (N_427,N_326,N_269);
or U428 (N_428,N_227,N_327);
and U429 (N_429,N_304,N_289);
nand U430 (N_430,N_309,N_265);
and U431 (N_431,N_266,N_236);
nor U432 (N_432,N_317,N_246);
xnor U433 (N_433,N_218,N_340);
and U434 (N_434,N_276,N_206);
and U435 (N_435,N_393,N_379);
and U436 (N_436,N_363,N_252);
nor U437 (N_437,N_282,N_345);
nor U438 (N_438,N_243,N_231);
or U439 (N_439,N_368,N_395);
nor U440 (N_440,N_244,N_341);
nor U441 (N_441,N_389,N_271);
or U442 (N_442,N_298,N_354);
and U443 (N_443,N_362,N_275);
nand U444 (N_444,N_387,N_337);
or U445 (N_445,N_347,N_397);
or U446 (N_446,N_302,N_335);
nor U447 (N_447,N_238,N_371);
nand U448 (N_448,N_241,N_294);
nand U449 (N_449,N_372,N_346);
and U450 (N_450,N_385,N_219);
and U451 (N_451,N_383,N_220);
or U452 (N_452,N_325,N_260);
and U453 (N_453,N_259,N_273);
nor U454 (N_454,N_301,N_329);
nand U455 (N_455,N_339,N_320);
or U456 (N_456,N_229,N_237);
or U457 (N_457,N_348,N_270);
nand U458 (N_458,N_399,N_213);
or U459 (N_459,N_367,N_328);
or U460 (N_460,N_277,N_299);
or U461 (N_461,N_332,N_388);
nor U462 (N_462,N_308,N_323);
nor U463 (N_463,N_207,N_377);
or U464 (N_464,N_274,N_358);
and U465 (N_465,N_287,N_357);
nand U466 (N_466,N_312,N_263);
nor U467 (N_467,N_314,N_230);
nand U468 (N_468,N_217,N_222);
and U469 (N_469,N_295,N_293);
or U470 (N_470,N_381,N_200);
nor U471 (N_471,N_224,N_394);
or U472 (N_472,N_334,N_386);
nor U473 (N_473,N_232,N_306);
nor U474 (N_474,N_392,N_342);
nand U475 (N_475,N_254,N_272);
and U476 (N_476,N_291,N_390);
and U477 (N_477,N_221,N_225);
nand U478 (N_478,N_280,N_373);
xor U479 (N_479,N_249,N_248);
or U480 (N_480,N_316,N_350);
or U481 (N_481,N_205,N_366);
and U482 (N_482,N_360,N_283);
nand U483 (N_483,N_384,N_374);
nand U484 (N_484,N_240,N_324);
or U485 (N_485,N_311,N_242);
or U486 (N_486,N_333,N_321);
and U487 (N_487,N_279,N_290);
and U488 (N_488,N_201,N_310);
nor U489 (N_489,N_391,N_264);
or U490 (N_490,N_297,N_262);
or U491 (N_491,N_396,N_319);
nand U492 (N_492,N_228,N_256);
nand U493 (N_493,N_284,N_281);
nand U494 (N_494,N_288,N_292);
nor U495 (N_495,N_376,N_226);
nand U496 (N_496,N_239,N_245);
nand U497 (N_497,N_203,N_338);
nor U498 (N_498,N_398,N_380);
or U499 (N_499,N_204,N_257);
nand U500 (N_500,N_329,N_339);
or U501 (N_501,N_394,N_293);
nor U502 (N_502,N_236,N_377);
xnor U503 (N_503,N_213,N_257);
nand U504 (N_504,N_288,N_387);
or U505 (N_505,N_231,N_248);
nand U506 (N_506,N_300,N_233);
nand U507 (N_507,N_340,N_203);
and U508 (N_508,N_276,N_284);
nor U509 (N_509,N_260,N_245);
or U510 (N_510,N_298,N_328);
and U511 (N_511,N_267,N_376);
and U512 (N_512,N_214,N_328);
and U513 (N_513,N_295,N_389);
nor U514 (N_514,N_227,N_292);
or U515 (N_515,N_306,N_319);
nand U516 (N_516,N_204,N_221);
and U517 (N_517,N_254,N_390);
nor U518 (N_518,N_210,N_290);
nand U519 (N_519,N_253,N_277);
xor U520 (N_520,N_396,N_347);
and U521 (N_521,N_252,N_345);
nor U522 (N_522,N_289,N_357);
nor U523 (N_523,N_328,N_345);
or U524 (N_524,N_286,N_315);
nand U525 (N_525,N_296,N_329);
and U526 (N_526,N_359,N_396);
nor U527 (N_527,N_329,N_324);
nor U528 (N_528,N_377,N_308);
or U529 (N_529,N_266,N_368);
or U530 (N_530,N_298,N_396);
or U531 (N_531,N_239,N_377);
or U532 (N_532,N_274,N_350);
and U533 (N_533,N_327,N_297);
nor U534 (N_534,N_290,N_284);
or U535 (N_535,N_219,N_232);
nor U536 (N_536,N_382,N_350);
or U537 (N_537,N_206,N_328);
and U538 (N_538,N_216,N_251);
nor U539 (N_539,N_262,N_279);
nand U540 (N_540,N_377,N_373);
and U541 (N_541,N_219,N_371);
or U542 (N_542,N_365,N_252);
nor U543 (N_543,N_325,N_278);
nor U544 (N_544,N_284,N_389);
nor U545 (N_545,N_268,N_319);
or U546 (N_546,N_206,N_323);
and U547 (N_547,N_354,N_203);
or U548 (N_548,N_218,N_319);
nor U549 (N_549,N_323,N_378);
and U550 (N_550,N_387,N_362);
nand U551 (N_551,N_325,N_330);
or U552 (N_552,N_273,N_386);
nand U553 (N_553,N_294,N_344);
or U554 (N_554,N_377,N_399);
or U555 (N_555,N_326,N_392);
or U556 (N_556,N_247,N_322);
nand U557 (N_557,N_218,N_265);
and U558 (N_558,N_233,N_246);
nor U559 (N_559,N_351,N_370);
and U560 (N_560,N_272,N_337);
and U561 (N_561,N_340,N_349);
or U562 (N_562,N_236,N_206);
nand U563 (N_563,N_230,N_335);
or U564 (N_564,N_317,N_399);
nor U565 (N_565,N_307,N_236);
nor U566 (N_566,N_329,N_258);
or U567 (N_567,N_314,N_227);
nor U568 (N_568,N_219,N_214);
nor U569 (N_569,N_329,N_328);
or U570 (N_570,N_239,N_319);
and U571 (N_571,N_354,N_376);
nand U572 (N_572,N_362,N_238);
nor U573 (N_573,N_353,N_227);
and U574 (N_574,N_395,N_293);
and U575 (N_575,N_390,N_270);
nor U576 (N_576,N_346,N_263);
or U577 (N_577,N_292,N_373);
or U578 (N_578,N_290,N_375);
xnor U579 (N_579,N_263,N_334);
and U580 (N_580,N_311,N_280);
and U581 (N_581,N_247,N_270);
or U582 (N_582,N_211,N_248);
or U583 (N_583,N_317,N_350);
or U584 (N_584,N_230,N_252);
nand U585 (N_585,N_285,N_379);
and U586 (N_586,N_260,N_248);
nor U587 (N_587,N_343,N_377);
nand U588 (N_588,N_209,N_216);
nor U589 (N_589,N_289,N_259);
nor U590 (N_590,N_333,N_360);
nand U591 (N_591,N_350,N_237);
nor U592 (N_592,N_254,N_208);
nand U593 (N_593,N_278,N_329);
nand U594 (N_594,N_344,N_287);
nor U595 (N_595,N_350,N_345);
xnor U596 (N_596,N_398,N_249);
xnor U597 (N_597,N_271,N_222);
or U598 (N_598,N_360,N_399);
nor U599 (N_599,N_370,N_373);
nor U600 (N_600,N_535,N_415);
and U601 (N_601,N_482,N_597);
nor U602 (N_602,N_528,N_476);
nor U603 (N_603,N_548,N_445);
nand U604 (N_604,N_582,N_418);
and U605 (N_605,N_449,N_561);
nor U606 (N_606,N_439,N_587);
nand U607 (N_607,N_573,N_401);
and U608 (N_608,N_450,N_579);
or U609 (N_609,N_454,N_531);
and U610 (N_610,N_478,N_409);
and U611 (N_611,N_514,N_524);
nor U612 (N_612,N_596,N_511);
nor U613 (N_613,N_461,N_487);
nand U614 (N_614,N_571,N_431);
or U615 (N_615,N_414,N_529);
or U616 (N_616,N_441,N_468);
and U617 (N_617,N_540,N_448);
nand U618 (N_618,N_547,N_570);
nor U619 (N_619,N_544,N_501);
nor U620 (N_620,N_477,N_552);
and U621 (N_621,N_444,N_568);
nor U622 (N_622,N_519,N_527);
or U623 (N_623,N_575,N_405);
and U624 (N_624,N_443,N_594);
nor U625 (N_625,N_475,N_518);
and U626 (N_626,N_536,N_435);
or U627 (N_627,N_410,N_549);
and U628 (N_628,N_492,N_526);
or U629 (N_629,N_403,N_442);
nand U630 (N_630,N_499,N_498);
nor U631 (N_631,N_555,N_564);
nand U632 (N_632,N_543,N_598);
nand U633 (N_633,N_473,N_497);
and U634 (N_634,N_457,N_485);
nor U635 (N_635,N_469,N_590);
or U636 (N_636,N_400,N_577);
and U637 (N_637,N_480,N_560);
nand U638 (N_638,N_525,N_488);
and U639 (N_639,N_495,N_422);
or U640 (N_640,N_533,N_586);
and U641 (N_641,N_496,N_592);
or U642 (N_642,N_412,N_486);
nor U643 (N_643,N_509,N_563);
nor U644 (N_644,N_411,N_433);
or U645 (N_645,N_506,N_578);
or U646 (N_646,N_532,N_589);
or U647 (N_647,N_440,N_446);
or U648 (N_648,N_407,N_430);
nor U649 (N_649,N_432,N_484);
nand U650 (N_650,N_416,N_503);
nor U651 (N_651,N_417,N_510);
and U652 (N_652,N_539,N_436);
or U653 (N_653,N_434,N_451);
and U654 (N_654,N_565,N_580);
nor U655 (N_655,N_413,N_456);
and U656 (N_656,N_493,N_467);
and U657 (N_657,N_479,N_470);
nor U658 (N_658,N_554,N_491);
or U659 (N_659,N_438,N_566);
or U660 (N_660,N_428,N_585);
and U661 (N_661,N_502,N_483);
or U662 (N_662,N_545,N_569);
or U663 (N_663,N_576,N_419);
or U664 (N_664,N_542,N_481);
nand U665 (N_665,N_558,N_462);
nand U666 (N_666,N_460,N_588);
and U667 (N_667,N_516,N_474);
and U668 (N_668,N_466,N_447);
nor U669 (N_669,N_472,N_504);
and U670 (N_670,N_530,N_595);
nand U671 (N_671,N_522,N_452);
nand U672 (N_672,N_562,N_515);
nand U673 (N_673,N_546,N_437);
or U674 (N_674,N_559,N_567);
and U675 (N_675,N_581,N_574);
and U676 (N_676,N_420,N_427);
nand U677 (N_677,N_507,N_424);
xnor U678 (N_678,N_517,N_538);
nand U679 (N_679,N_404,N_556);
nand U680 (N_680,N_593,N_408);
nor U681 (N_681,N_551,N_572);
and U682 (N_682,N_550,N_425);
and U683 (N_683,N_500,N_458);
or U684 (N_684,N_523,N_406);
or U685 (N_685,N_490,N_505);
and U686 (N_686,N_508,N_421);
or U687 (N_687,N_537,N_557);
nand U688 (N_688,N_520,N_463);
or U689 (N_689,N_494,N_426);
and U690 (N_690,N_591,N_553);
or U691 (N_691,N_429,N_584);
nor U692 (N_692,N_489,N_512);
nand U693 (N_693,N_402,N_583);
nand U694 (N_694,N_423,N_541);
or U695 (N_695,N_459,N_534);
nand U696 (N_696,N_453,N_521);
or U697 (N_697,N_599,N_513);
or U698 (N_698,N_465,N_455);
nor U699 (N_699,N_464,N_471);
nand U700 (N_700,N_459,N_558);
or U701 (N_701,N_575,N_595);
nor U702 (N_702,N_480,N_569);
and U703 (N_703,N_420,N_571);
nor U704 (N_704,N_483,N_509);
nand U705 (N_705,N_439,N_572);
or U706 (N_706,N_425,N_462);
or U707 (N_707,N_541,N_540);
and U708 (N_708,N_549,N_453);
or U709 (N_709,N_557,N_496);
nor U710 (N_710,N_476,N_434);
xnor U711 (N_711,N_400,N_498);
nand U712 (N_712,N_435,N_402);
nand U713 (N_713,N_535,N_598);
or U714 (N_714,N_408,N_480);
nand U715 (N_715,N_514,N_474);
or U716 (N_716,N_555,N_504);
nand U717 (N_717,N_536,N_526);
and U718 (N_718,N_592,N_545);
xor U719 (N_719,N_460,N_545);
or U720 (N_720,N_595,N_579);
or U721 (N_721,N_422,N_411);
and U722 (N_722,N_428,N_512);
xor U723 (N_723,N_490,N_404);
and U724 (N_724,N_552,N_439);
or U725 (N_725,N_540,N_426);
and U726 (N_726,N_500,N_518);
or U727 (N_727,N_447,N_457);
nand U728 (N_728,N_589,N_433);
or U729 (N_729,N_488,N_528);
nor U730 (N_730,N_510,N_524);
or U731 (N_731,N_453,N_487);
nor U732 (N_732,N_469,N_464);
or U733 (N_733,N_455,N_469);
nand U734 (N_734,N_401,N_486);
and U735 (N_735,N_591,N_559);
nand U736 (N_736,N_546,N_459);
and U737 (N_737,N_510,N_444);
and U738 (N_738,N_428,N_409);
and U739 (N_739,N_516,N_563);
or U740 (N_740,N_547,N_456);
or U741 (N_741,N_520,N_499);
nand U742 (N_742,N_542,N_549);
nand U743 (N_743,N_553,N_503);
nor U744 (N_744,N_425,N_421);
nor U745 (N_745,N_562,N_434);
or U746 (N_746,N_455,N_433);
and U747 (N_747,N_522,N_585);
or U748 (N_748,N_495,N_406);
and U749 (N_749,N_449,N_445);
nor U750 (N_750,N_489,N_485);
xor U751 (N_751,N_472,N_465);
and U752 (N_752,N_464,N_443);
nand U753 (N_753,N_438,N_475);
xor U754 (N_754,N_560,N_413);
and U755 (N_755,N_519,N_532);
and U756 (N_756,N_565,N_526);
nor U757 (N_757,N_407,N_501);
nor U758 (N_758,N_550,N_413);
or U759 (N_759,N_539,N_564);
nor U760 (N_760,N_408,N_443);
nor U761 (N_761,N_579,N_541);
nor U762 (N_762,N_486,N_510);
nor U763 (N_763,N_445,N_584);
or U764 (N_764,N_469,N_466);
and U765 (N_765,N_411,N_416);
nor U766 (N_766,N_422,N_547);
and U767 (N_767,N_457,N_412);
or U768 (N_768,N_580,N_475);
nand U769 (N_769,N_589,N_580);
nand U770 (N_770,N_440,N_565);
or U771 (N_771,N_462,N_482);
nor U772 (N_772,N_554,N_512);
or U773 (N_773,N_441,N_582);
nor U774 (N_774,N_437,N_480);
and U775 (N_775,N_456,N_540);
nand U776 (N_776,N_450,N_591);
xor U777 (N_777,N_577,N_425);
and U778 (N_778,N_559,N_420);
nor U779 (N_779,N_579,N_571);
and U780 (N_780,N_588,N_585);
nand U781 (N_781,N_503,N_424);
or U782 (N_782,N_534,N_435);
nand U783 (N_783,N_545,N_405);
nand U784 (N_784,N_570,N_443);
nor U785 (N_785,N_566,N_497);
and U786 (N_786,N_413,N_488);
nand U787 (N_787,N_476,N_549);
or U788 (N_788,N_517,N_597);
and U789 (N_789,N_460,N_487);
nand U790 (N_790,N_565,N_547);
and U791 (N_791,N_476,N_433);
nor U792 (N_792,N_550,N_597);
or U793 (N_793,N_478,N_575);
or U794 (N_794,N_458,N_594);
and U795 (N_795,N_451,N_448);
and U796 (N_796,N_560,N_582);
and U797 (N_797,N_401,N_419);
xor U798 (N_798,N_583,N_448);
and U799 (N_799,N_495,N_438);
nor U800 (N_800,N_753,N_725);
and U801 (N_801,N_617,N_793);
and U802 (N_802,N_769,N_749);
and U803 (N_803,N_676,N_646);
nand U804 (N_804,N_746,N_663);
nand U805 (N_805,N_779,N_667);
and U806 (N_806,N_620,N_628);
or U807 (N_807,N_641,N_665);
or U808 (N_808,N_684,N_739);
nor U809 (N_809,N_724,N_696);
nand U810 (N_810,N_709,N_629);
and U811 (N_811,N_690,N_758);
nand U812 (N_812,N_650,N_736);
or U813 (N_813,N_695,N_777);
and U814 (N_814,N_612,N_608);
or U815 (N_815,N_773,N_688);
nor U816 (N_816,N_619,N_697);
or U817 (N_817,N_780,N_673);
or U818 (N_818,N_607,N_674);
or U819 (N_819,N_655,N_741);
nor U820 (N_820,N_601,N_718);
nor U821 (N_821,N_638,N_711);
nor U822 (N_822,N_727,N_630);
and U823 (N_823,N_679,N_645);
nand U824 (N_824,N_759,N_634);
or U825 (N_825,N_687,N_657);
nand U826 (N_826,N_656,N_751);
nand U827 (N_827,N_770,N_635);
and U828 (N_828,N_787,N_776);
nand U829 (N_829,N_774,N_745);
nand U830 (N_830,N_721,N_636);
nand U831 (N_831,N_671,N_789);
nand U832 (N_832,N_742,N_798);
nor U833 (N_833,N_784,N_642);
and U834 (N_834,N_735,N_706);
nand U835 (N_835,N_639,N_707);
and U836 (N_836,N_717,N_654);
or U837 (N_837,N_653,N_720);
nor U838 (N_838,N_652,N_783);
nor U839 (N_839,N_734,N_614);
and U840 (N_840,N_765,N_730);
nor U841 (N_841,N_791,N_748);
and U842 (N_842,N_767,N_691);
and U843 (N_843,N_775,N_731);
nand U844 (N_844,N_703,N_668);
nor U845 (N_845,N_604,N_627);
and U846 (N_846,N_708,N_719);
or U847 (N_847,N_738,N_678);
and U848 (N_848,N_651,N_796);
or U849 (N_849,N_752,N_714);
xor U850 (N_850,N_682,N_611);
and U851 (N_851,N_672,N_680);
and U852 (N_852,N_771,N_768);
and U853 (N_853,N_686,N_700);
nor U854 (N_854,N_747,N_615);
or U855 (N_855,N_681,N_694);
and U856 (N_856,N_755,N_754);
and U857 (N_857,N_609,N_795);
and U858 (N_858,N_662,N_623);
and U859 (N_859,N_649,N_661);
nor U860 (N_860,N_733,N_766);
or U861 (N_861,N_797,N_701);
nand U862 (N_862,N_762,N_713);
nand U863 (N_863,N_764,N_772);
nor U864 (N_864,N_723,N_610);
or U865 (N_865,N_613,N_632);
or U866 (N_866,N_737,N_750);
and U867 (N_867,N_740,N_716);
nand U868 (N_868,N_626,N_643);
or U869 (N_869,N_644,N_677);
nor U870 (N_870,N_647,N_685);
xor U871 (N_871,N_603,N_616);
and U872 (N_872,N_778,N_618);
nand U873 (N_873,N_799,N_658);
nor U874 (N_874,N_785,N_683);
or U875 (N_875,N_743,N_689);
nor U876 (N_876,N_622,N_666);
nor U877 (N_877,N_637,N_664);
nand U878 (N_878,N_794,N_704);
nand U879 (N_879,N_669,N_763);
nor U880 (N_880,N_782,N_786);
or U881 (N_881,N_790,N_631);
nor U882 (N_882,N_624,N_659);
and U883 (N_883,N_675,N_640);
or U884 (N_884,N_744,N_699);
and U885 (N_885,N_698,N_625);
and U886 (N_886,N_792,N_761);
or U887 (N_887,N_760,N_722);
nand U888 (N_888,N_602,N_660);
or U889 (N_889,N_693,N_621);
nand U890 (N_890,N_726,N_712);
nor U891 (N_891,N_729,N_605);
or U892 (N_892,N_648,N_788);
nand U893 (N_893,N_710,N_781);
nor U894 (N_894,N_702,N_728);
or U895 (N_895,N_606,N_670);
or U896 (N_896,N_732,N_633);
or U897 (N_897,N_600,N_692);
nand U898 (N_898,N_715,N_756);
and U899 (N_899,N_705,N_757);
and U900 (N_900,N_794,N_685);
nor U901 (N_901,N_745,N_710);
or U902 (N_902,N_783,N_654);
nand U903 (N_903,N_647,N_728);
or U904 (N_904,N_764,N_769);
xor U905 (N_905,N_676,N_776);
xnor U906 (N_906,N_772,N_680);
nor U907 (N_907,N_667,N_735);
nand U908 (N_908,N_608,N_681);
nand U909 (N_909,N_663,N_789);
nor U910 (N_910,N_675,N_799);
nand U911 (N_911,N_787,N_627);
and U912 (N_912,N_756,N_675);
or U913 (N_913,N_787,N_767);
nand U914 (N_914,N_748,N_756);
nand U915 (N_915,N_772,N_768);
nor U916 (N_916,N_704,N_750);
nand U917 (N_917,N_719,N_705);
nand U918 (N_918,N_733,N_760);
and U919 (N_919,N_603,N_670);
and U920 (N_920,N_727,N_650);
nor U921 (N_921,N_630,N_759);
nor U922 (N_922,N_683,N_676);
or U923 (N_923,N_771,N_773);
and U924 (N_924,N_765,N_677);
and U925 (N_925,N_631,N_782);
or U926 (N_926,N_741,N_650);
or U927 (N_927,N_642,N_756);
nand U928 (N_928,N_750,N_606);
and U929 (N_929,N_653,N_680);
and U930 (N_930,N_687,N_797);
or U931 (N_931,N_773,N_646);
nor U932 (N_932,N_680,N_645);
nand U933 (N_933,N_655,N_601);
or U934 (N_934,N_760,N_723);
and U935 (N_935,N_747,N_676);
nor U936 (N_936,N_719,N_611);
and U937 (N_937,N_790,N_768);
nor U938 (N_938,N_750,N_720);
nor U939 (N_939,N_659,N_723);
and U940 (N_940,N_684,N_738);
nand U941 (N_941,N_640,N_626);
and U942 (N_942,N_608,N_724);
nor U943 (N_943,N_644,N_619);
nand U944 (N_944,N_682,N_650);
nor U945 (N_945,N_794,N_668);
and U946 (N_946,N_734,N_654);
nand U947 (N_947,N_739,N_726);
xor U948 (N_948,N_674,N_629);
nand U949 (N_949,N_612,N_630);
and U950 (N_950,N_764,N_646);
or U951 (N_951,N_675,N_791);
nand U952 (N_952,N_676,N_605);
nor U953 (N_953,N_672,N_633);
nor U954 (N_954,N_680,N_789);
nand U955 (N_955,N_711,N_672);
or U956 (N_956,N_663,N_734);
or U957 (N_957,N_683,N_617);
or U958 (N_958,N_655,N_636);
nand U959 (N_959,N_717,N_643);
nor U960 (N_960,N_652,N_666);
or U961 (N_961,N_778,N_627);
or U962 (N_962,N_774,N_632);
or U963 (N_963,N_600,N_798);
nor U964 (N_964,N_761,N_781);
nor U965 (N_965,N_686,N_781);
and U966 (N_966,N_606,N_705);
or U967 (N_967,N_647,N_775);
and U968 (N_968,N_610,N_645);
or U969 (N_969,N_609,N_771);
nor U970 (N_970,N_769,N_779);
or U971 (N_971,N_650,N_754);
or U972 (N_972,N_604,N_647);
nand U973 (N_973,N_643,N_699);
and U974 (N_974,N_744,N_618);
and U975 (N_975,N_655,N_628);
nor U976 (N_976,N_746,N_763);
nor U977 (N_977,N_718,N_668);
nor U978 (N_978,N_689,N_719);
nand U979 (N_979,N_668,N_749);
nor U980 (N_980,N_621,N_692);
or U981 (N_981,N_601,N_636);
nor U982 (N_982,N_795,N_682);
nand U983 (N_983,N_667,N_659);
and U984 (N_984,N_611,N_776);
nor U985 (N_985,N_661,N_701);
nor U986 (N_986,N_704,N_666);
nor U987 (N_987,N_649,N_751);
nor U988 (N_988,N_692,N_795);
and U989 (N_989,N_639,N_628);
or U990 (N_990,N_728,N_686);
xnor U991 (N_991,N_732,N_757);
nor U992 (N_992,N_681,N_656);
and U993 (N_993,N_776,N_644);
nand U994 (N_994,N_783,N_693);
and U995 (N_995,N_754,N_664);
nand U996 (N_996,N_660,N_656);
or U997 (N_997,N_724,N_600);
and U998 (N_998,N_786,N_677);
or U999 (N_999,N_783,N_793);
or U1000 (N_1000,N_849,N_838);
nor U1001 (N_1001,N_847,N_927);
nand U1002 (N_1002,N_971,N_974);
or U1003 (N_1003,N_985,N_900);
or U1004 (N_1004,N_889,N_960);
and U1005 (N_1005,N_888,N_873);
nor U1006 (N_1006,N_866,N_980);
and U1007 (N_1007,N_881,N_916);
nand U1008 (N_1008,N_904,N_989);
and U1009 (N_1009,N_879,N_958);
nor U1010 (N_1010,N_902,N_996);
or U1011 (N_1011,N_874,N_869);
nor U1012 (N_1012,N_997,N_875);
and U1013 (N_1013,N_969,N_843);
nor U1014 (N_1014,N_801,N_800);
nand U1015 (N_1015,N_906,N_912);
or U1016 (N_1016,N_820,N_984);
or U1017 (N_1017,N_844,N_898);
and U1018 (N_1018,N_831,N_834);
or U1019 (N_1019,N_911,N_872);
nor U1020 (N_1020,N_812,N_821);
and U1021 (N_1021,N_810,N_817);
and U1022 (N_1022,N_860,N_840);
nor U1023 (N_1023,N_887,N_924);
nand U1024 (N_1024,N_992,N_846);
xor U1025 (N_1025,N_982,N_963);
nand U1026 (N_1026,N_948,N_914);
nor U1027 (N_1027,N_897,N_936);
and U1028 (N_1028,N_962,N_892);
xor U1029 (N_1029,N_908,N_944);
and U1030 (N_1030,N_933,N_921);
or U1031 (N_1031,N_907,N_991);
nor U1032 (N_1032,N_839,N_825);
nor U1033 (N_1033,N_853,N_932);
or U1034 (N_1034,N_951,N_885);
nor U1035 (N_1035,N_949,N_998);
or U1036 (N_1036,N_965,N_895);
nor U1037 (N_1037,N_942,N_999);
nand U1038 (N_1038,N_935,N_857);
nand U1039 (N_1039,N_808,N_976);
nor U1040 (N_1040,N_905,N_882);
or U1041 (N_1041,N_957,N_811);
or U1042 (N_1042,N_883,N_913);
nor U1043 (N_1043,N_993,N_804);
and U1044 (N_1044,N_823,N_862);
nor U1045 (N_1045,N_918,N_878);
nand U1046 (N_1046,N_954,N_937);
nand U1047 (N_1047,N_864,N_972);
xor U1048 (N_1048,N_922,N_968);
nor U1049 (N_1049,N_995,N_929);
or U1050 (N_1050,N_930,N_955);
and U1051 (N_1051,N_870,N_822);
nor U1052 (N_1052,N_893,N_863);
and U1053 (N_1053,N_966,N_832);
and U1054 (N_1054,N_826,N_842);
nor U1055 (N_1055,N_950,N_915);
nand U1056 (N_1056,N_824,N_837);
and U1057 (N_1057,N_871,N_865);
and U1058 (N_1058,N_956,N_977);
and U1059 (N_1059,N_833,N_959);
nor U1060 (N_1060,N_880,N_941);
and U1061 (N_1061,N_926,N_939);
and U1062 (N_1062,N_859,N_836);
nor U1063 (N_1063,N_981,N_986);
nand U1064 (N_1064,N_815,N_901);
or U1065 (N_1065,N_945,N_920);
nand U1066 (N_1066,N_899,N_953);
nand U1067 (N_1067,N_827,N_970);
and U1068 (N_1068,N_946,N_814);
and U1069 (N_1069,N_990,N_877);
nand U1070 (N_1070,N_983,N_919);
and U1071 (N_1071,N_829,N_923);
and U1072 (N_1072,N_876,N_975);
nor U1073 (N_1073,N_909,N_848);
and U1074 (N_1074,N_818,N_994);
nand U1075 (N_1075,N_884,N_841);
or U1076 (N_1076,N_861,N_819);
nor U1077 (N_1077,N_979,N_978);
and U1078 (N_1078,N_903,N_855);
nor U1079 (N_1079,N_910,N_828);
nand U1080 (N_1080,N_987,N_940);
nand U1081 (N_1081,N_947,N_813);
nand U1082 (N_1082,N_925,N_917);
and U1083 (N_1083,N_886,N_890);
nor U1084 (N_1084,N_896,N_802);
and U1085 (N_1085,N_805,N_807);
and U1086 (N_1086,N_894,N_967);
and U1087 (N_1087,N_830,N_891);
nand U1088 (N_1088,N_851,N_854);
and U1089 (N_1089,N_931,N_835);
nand U1090 (N_1090,N_868,N_852);
and U1091 (N_1091,N_850,N_938);
and U1092 (N_1092,N_961,N_845);
and U1093 (N_1093,N_803,N_867);
and U1094 (N_1094,N_973,N_952);
and U1095 (N_1095,N_928,N_964);
nor U1096 (N_1096,N_934,N_816);
and U1097 (N_1097,N_943,N_809);
or U1098 (N_1098,N_858,N_856);
nor U1099 (N_1099,N_806,N_988);
and U1100 (N_1100,N_989,N_951);
and U1101 (N_1101,N_897,N_996);
and U1102 (N_1102,N_861,N_803);
nand U1103 (N_1103,N_838,N_993);
and U1104 (N_1104,N_984,N_959);
and U1105 (N_1105,N_818,N_868);
or U1106 (N_1106,N_875,N_882);
and U1107 (N_1107,N_943,N_808);
nor U1108 (N_1108,N_897,N_985);
or U1109 (N_1109,N_858,N_829);
nand U1110 (N_1110,N_968,N_943);
and U1111 (N_1111,N_805,N_925);
and U1112 (N_1112,N_847,N_991);
or U1113 (N_1113,N_910,N_958);
and U1114 (N_1114,N_835,N_847);
nor U1115 (N_1115,N_800,N_960);
nand U1116 (N_1116,N_981,N_893);
nor U1117 (N_1117,N_938,N_919);
nor U1118 (N_1118,N_832,N_860);
nand U1119 (N_1119,N_983,N_857);
and U1120 (N_1120,N_996,N_893);
or U1121 (N_1121,N_824,N_907);
or U1122 (N_1122,N_947,N_833);
xnor U1123 (N_1123,N_977,N_806);
nor U1124 (N_1124,N_815,N_846);
nor U1125 (N_1125,N_813,N_838);
nor U1126 (N_1126,N_842,N_990);
nor U1127 (N_1127,N_823,N_892);
and U1128 (N_1128,N_900,N_802);
or U1129 (N_1129,N_828,N_942);
and U1130 (N_1130,N_801,N_854);
nand U1131 (N_1131,N_982,N_804);
nor U1132 (N_1132,N_906,N_891);
nand U1133 (N_1133,N_873,N_828);
or U1134 (N_1134,N_963,N_908);
and U1135 (N_1135,N_988,N_979);
nor U1136 (N_1136,N_949,N_966);
and U1137 (N_1137,N_801,N_823);
nand U1138 (N_1138,N_917,N_834);
and U1139 (N_1139,N_836,N_977);
nor U1140 (N_1140,N_948,N_928);
nor U1141 (N_1141,N_915,N_898);
nor U1142 (N_1142,N_941,N_968);
nor U1143 (N_1143,N_811,N_867);
or U1144 (N_1144,N_924,N_864);
or U1145 (N_1145,N_882,N_989);
and U1146 (N_1146,N_828,N_940);
nand U1147 (N_1147,N_916,N_861);
xor U1148 (N_1148,N_888,N_858);
and U1149 (N_1149,N_850,N_942);
nand U1150 (N_1150,N_942,N_857);
and U1151 (N_1151,N_819,N_967);
nand U1152 (N_1152,N_968,N_938);
nor U1153 (N_1153,N_831,N_847);
nor U1154 (N_1154,N_851,N_967);
and U1155 (N_1155,N_872,N_864);
or U1156 (N_1156,N_956,N_982);
nor U1157 (N_1157,N_805,N_988);
or U1158 (N_1158,N_944,N_871);
nand U1159 (N_1159,N_896,N_814);
nor U1160 (N_1160,N_887,N_805);
or U1161 (N_1161,N_984,N_990);
nor U1162 (N_1162,N_919,N_972);
and U1163 (N_1163,N_823,N_811);
nor U1164 (N_1164,N_800,N_991);
xnor U1165 (N_1165,N_935,N_918);
nor U1166 (N_1166,N_859,N_960);
nor U1167 (N_1167,N_830,N_838);
nor U1168 (N_1168,N_957,N_960);
nand U1169 (N_1169,N_906,N_882);
or U1170 (N_1170,N_853,N_926);
nor U1171 (N_1171,N_891,N_844);
and U1172 (N_1172,N_930,N_830);
nor U1173 (N_1173,N_865,N_923);
or U1174 (N_1174,N_945,N_950);
nand U1175 (N_1175,N_985,N_856);
nand U1176 (N_1176,N_918,N_984);
or U1177 (N_1177,N_975,N_988);
nor U1178 (N_1178,N_810,N_910);
nand U1179 (N_1179,N_944,N_884);
or U1180 (N_1180,N_884,N_869);
xor U1181 (N_1181,N_801,N_904);
nor U1182 (N_1182,N_837,N_817);
nand U1183 (N_1183,N_888,N_954);
nor U1184 (N_1184,N_875,N_844);
or U1185 (N_1185,N_876,N_921);
or U1186 (N_1186,N_931,N_819);
nor U1187 (N_1187,N_832,N_907);
nand U1188 (N_1188,N_884,N_865);
nand U1189 (N_1189,N_893,N_952);
and U1190 (N_1190,N_996,N_965);
and U1191 (N_1191,N_873,N_947);
nor U1192 (N_1192,N_934,N_893);
nand U1193 (N_1193,N_810,N_948);
or U1194 (N_1194,N_990,N_805);
nand U1195 (N_1195,N_954,N_897);
nor U1196 (N_1196,N_867,N_909);
nand U1197 (N_1197,N_846,N_851);
and U1198 (N_1198,N_955,N_933);
and U1199 (N_1199,N_959,N_937);
nand U1200 (N_1200,N_1017,N_1139);
nand U1201 (N_1201,N_1108,N_1042);
nor U1202 (N_1202,N_1171,N_1013);
nor U1203 (N_1203,N_1162,N_1047);
and U1204 (N_1204,N_1161,N_1164);
nor U1205 (N_1205,N_1031,N_1011);
nand U1206 (N_1206,N_1051,N_1127);
nor U1207 (N_1207,N_1155,N_1055);
nand U1208 (N_1208,N_1122,N_1094);
nand U1209 (N_1209,N_1098,N_1030);
nand U1210 (N_1210,N_1039,N_1109);
or U1211 (N_1211,N_1079,N_1145);
nor U1212 (N_1212,N_1008,N_1197);
and U1213 (N_1213,N_1115,N_1172);
and U1214 (N_1214,N_1028,N_1080);
nand U1215 (N_1215,N_1140,N_1173);
nand U1216 (N_1216,N_1018,N_1129);
nand U1217 (N_1217,N_1100,N_1043);
and U1218 (N_1218,N_1069,N_1001);
nor U1219 (N_1219,N_1167,N_1006);
xor U1220 (N_1220,N_1007,N_1072);
and U1221 (N_1221,N_1132,N_1163);
nor U1222 (N_1222,N_1104,N_1189);
nor U1223 (N_1223,N_1009,N_1074);
and U1224 (N_1224,N_1123,N_1199);
nand U1225 (N_1225,N_1023,N_1148);
nand U1226 (N_1226,N_1086,N_1093);
and U1227 (N_1227,N_1137,N_1185);
or U1228 (N_1228,N_1166,N_1087);
or U1229 (N_1229,N_1063,N_1078);
and U1230 (N_1230,N_1022,N_1095);
nor U1231 (N_1231,N_1113,N_1062);
nor U1232 (N_1232,N_1107,N_1136);
nor U1233 (N_1233,N_1082,N_1056);
nor U1234 (N_1234,N_1154,N_1182);
and U1235 (N_1235,N_1065,N_1010);
nand U1236 (N_1236,N_1125,N_1119);
and U1237 (N_1237,N_1046,N_1057);
nand U1238 (N_1238,N_1138,N_1091);
and U1239 (N_1239,N_1120,N_1053);
nand U1240 (N_1240,N_1160,N_1038);
nor U1241 (N_1241,N_1179,N_1012);
nor U1242 (N_1242,N_1124,N_1060);
and U1243 (N_1243,N_1196,N_1186);
nand U1244 (N_1244,N_1158,N_1076);
xor U1245 (N_1245,N_1090,N_1116);
nor U1246 (N_1246,N_1000,N_1066);
nand U1247 (N_1247,N_1143,N_1170);
and U1248 (N_1248,N_1024,N_1105);
nor U1249 (N_1249,N_1111,N_1044);
or U1250 (N_1250,N_1178,N_1102);
nand U1251 (N_1251,N_1058,N_1188);
nand U1252 (N_1252,N_1150,N_1067);
and U1253 (N_1253,N_1190,N_1005);
and U1254 (N_1254,N_1131,N_1121);
nand U1255 (N_1255,N_1177,N_1027);
and U1256 (N_1256,N_1133,N_1097);
or U1257 (N_1257,N_1004,N_1029);
and U1258 (N_1258,N_1151,N_1184);
nor U1259 (N_1259,N_1157,N_1075);
and U1260 (N_1260,N_1073,N_1002);
and U1261 (N_1261,N_1134,N_1141);
nor U1262 (N_1262,N_1103,N_1025);
nor U1263 (N_1263,N_1033,N_1019);
and U1264 (N_1264,N_1142,N_1165);
nor U1265 (N_1265,N_1037,N_1096);
and U1266 (N_1266,N_1176,N_1088);
or U1267 (N_1267,N_1020,N_1045);
or U1268 (N_1268,N_1036,N_1149);
xor U1269 (N_1269,N_1003,N_1193);
nor U1270 (N_1270,N_1135,N_1052);
nor U1271 (N_1271,N_1049,N_1180);
nand U1272 (N_1272,N_1153,N_1181);
nor U1273 (N_1273,N_1083,N_1175);
nor U1274 (N_1274,N_1112,N_1014);
or U1275 (N_1275,N_1128,N_1068);
and U1276 (N_1276,N_1050,N_1092);
or U1277 (N_1277,N_1198,N_1085);
nor U1278 (N_1278,N_1034,N_1117);
or U1279 (N_1279,N_1130,N_1021);
nor U1280 (N_1280,N_1152,N_1126);
xnor U1281 (N_1281,N_1183,N_1118);
and U1282 (N_1282,N_1081,N_1159);
and U1283 (N_1283,N_1101,N_1084);
nor U1284 (N_1284,N_1110,N_1144);
nor U1285 (N_1285,N_1015,N_1061);
nand U1286 (N_1286,N_1156,N_1048);
or U1287 (N_1287,N_1195,N_1070);
and U1288 (N_1288,N_1192,N_1026);
nand U1289 (N_1289,N_1099,N_1191);
and U1290 (N_1290,N_1089,N_1106);
nor U1291 (N_1291,N_1146,N_1041);
or U1292 (N_1292,N_1059,N_1114);
and U1293 (N_1293,N_1016,N_1169);
nand U1294 (N_1294,N_1032,N_1147);
nand U1295 (N_1295,N_1194,N_1054);
xnor U1296 (N_1296,N_1174,N_1035);
nor U1297 (N_1297,N_1040,N_1071);
and U1298 (N_1298,N_1077,N_1064);
nor U1299 (N_1299,N_1168,N_1187);
and U1300 (N_1300,N_1185,N_1164);
nand U1301 (N_1301,N_1058,N_1048);
or U1302 (N_1302,N_1199,N_1007);
or U1303 (N_1303,N_1117,N_1056);
or U1304 (N_1304,N_1103,N_1179);
and U1305 (N_1305,N_1084,N_1052);
or U1306 (N_1306,N_1041,N_1090);
nand U1307 (N_1307,N_1013,N_1144);
nor U1308 (N_1308,N_1172,N_1181);
and U1309 (N_1309,N_1153,N_1162);
nor U1310 (N_1310,N_1055,N_1168);
nor U1311 (N_1311,N_1033,N_1145);
nor U1312 (N_1312,N_1055,N_1156);
nor U1313 (N_1313,N_1070,N_1126);
nand U1314 (N_1314,N_1062,N_1064);
nand U1315 (N_1315,N_1187,N_1093);
nor U1316 (N_1316,N_1059,N_1189);
and U1317 (N_1317,N_1010,N_1060);
nor U1318 (N_1318,N_1009,N_1078);
nor U1319 (N_1319,N_1146,N_1121);
nand U1320 (N_1320,N_1199,N_1124);
and U1321 (N_1321,N_1026,N_1040);
or U1322 (N_1322,N_1016,N_1129);
nand U1323 (N_1323,N_1189,N_1024);
xnor U1324 (N_1324,N_1164,N_1033);
nor U1325 (N_1325,N_1176,N_1133);
or U1326 (N_1326,N_1105,N_1036);
and U1327 (N_1327,N_1176,N_1131);
nand U1328 (N_1328,N_1122,N_1118);
and U1329 (N_1329,N_1081,N_1082);
or U1330 (N_1330,N_1072,N_1052);
nor U1331 (N_1331,N_1112,N_1077);
and U1332 (N_1332,N_1175,N_1119);
nor U1333 (N_1333,N_1043,N_1192);
nor U1334 (N_1334,N_1046,N_1036);
nand U1335 (N_1335,N_1137,N_1125);
nor U1336 (N_1336,N_1183,N_1135);
nand U1337 (N_1337,N_1013,N_1177);
and U1338 (N_1338,N_1139,N_1005);
xnor U1339 (N_1339,N_1102,N_1081);
or U1340 (N_1340,N_1126,N_1114);
nor U1341 (N_1341,N_1129,N_1162);
nor U1342 (N_1342,N_1138,N_1068);
and U1343 (N_1343,N_1159,N_1071);
nor U1344 (N_1344,N_1037,N_1135);
or U1345 (N_1345,N_1196,N_1138);
and U1346 (N_1346,N_1115,N_1120);
or U1347 (N_1347,N_1130,N_1163);
nand U1348 (N_1348,N_1164,N_1078);
nand U1349 (N_1349,N_1128,N_1123);
or U1350 (N_1350,N_1028,N_1001);
or U1351 (N_1351,N_1199,N_1111);
or U1352 (N_1352,N_1042,N_1080);
nor U1353 (N_1353,N_1129,N_1098);
nand U1354 (N_1354,N_1112,N_1005);
xnor U1355 (N_1355,N_1032,N_1031);
and U1356 (N_1356,N_1144,N_1103);
nand U1357 (N_1357,N_1140,N_1123);
or U1358 (N_1358,N_1001,N_1095);
and U1359 (N_1359,N_1192,N_1080);
and U1360 (N_1360,N_1121,N_1088);
or U1361 (N_1361,N_1144,N_1071);
xnor U1362 (N_1362,N_1082,N_1010);
or U1363 (N_1363,N_1135,N_1153);
and U1364 (N_1364,N_1108,N_1139);
or U1365 (N_1365,N_1179,N_1168);
nor U1366 (N_1366,N_1156,N_1178);
nand U1367 (N_1367,N_1160,N_1177);
nand U1368 (N_1368,N_1042,N_1084);
and U1369 (N_1369,N_1122,N_1146);
nor U1370 (N_1370,N_1110,N_1196);
xnor U1371 (N_1371,N_1198,N_1007);
nor U1372 (N_1372,N_1136,N_1097);
nor U1373 (N_1373,N_1038,N_1165);
and U1374 (N_1374,N_1072,N_1129);
nor U1375 (N_1375,N_1062,N_1069);
and U1376 (N_1376,N_1161,N_1115);
nor U1377 (N_1377,N_1103,N_1155);
nand U1378 (N_1378,N_1196,N_1188);
nor U1379 (N_1379,N_1120,N_1082);
and U1380 (N_1380,N_1114,N_1108);
nor U1381 (N_1381,N_1169,N_1124);
or U1382 (N_1382,N_1125,N_1076);
nor U1383 (N_1383,N_1141,N_1174);
nand U1384 (N_1384,N_1152,N_1086);
or U1385 (N_1385,N_1086,N_1061);
nand U1386 (N_1386,N_1136,N_1004);
and U1387 (N_1387,N_1036,N_1057);
or U1388 (N_1388,N_1095,N_1182);
nand U1389 (N_1389,N_1003,N_1063);
or U1390 (N_1390,N_1199,N_1133);
nor U1391 (N_1391,N_1143,N_1028);
nand U1392 (N_1392,N_1048,N_1029);
or U1393 (N_1393,N_1018,N_1126);
nand U1394 (N_1394,N_1060,N_1190);
or U1395 (N_1395,N_1192,N_1033);
or U1396 (N_1396,N_1040,N_1198);
nor U1397 (N_1397,N_1159,N_1020);
and U1398 (N_1398,N_1025,N_1100);
and U1399 (N_1399,N_1127,N_1166);
or U1400 (N_1400,N_1395,N_1213);
or U1401 (N_1401,N_1299,N_1247);
nand U1402 (N_1402,N_1346,N_1349);
and U1403 (N_1403,N_1362,N_1365);
and U1404 (N_1404,N_1369,N_1323);
and U1405 (N_1405,N_1236,N_1356);
and U1406 (N_1406,N_1387,N_1277);
nor U1407 (N_1407,N_1237,N_1228);
or U1408 (N_1408,N_1378,N_1211);
xnor U1409 (N_1409,N_1389,N_1363);
nor U1410 (N_1410,N_1278,N_1344);
nor U1411 (N_1411,N_1215,N_1243);
or U1412 (N_1412,N_1245,N_1287);
nand U1413 (N_1413,N_1286,N_1251);
or U1414 (N_1414,N_1290,N_1386);
nor U1415 (N_1415,N_1264,N_1309);
or U1416 (N_1416,N_1273,N_1242);
nor U1417 (N_1417,N_1212,N_1210);
xor U1418 (N_1418,N_1391,N_1267);
nand U1419 (N_1419,N_1366,N_1229);
nor U1420 (N_1420,N_1218,N_1260);
nand U1421 (N_1421,N_1393,N_1246);
and U1422 (N_1422,N_1382,N_1216);
nand U1423 (N_1423,N_1300,N_1310);
or U1424 (N_1424,N_1308,N_1312);
nand U1425 (N_1425,N_1253,N_1303);
or U1426 (N_1426,N_1222,N_1291);
nor U1427 (N_1427,N_1330,N_1332);
and U1428 (N_1428,N_1374,N_1252);
nor U1429 (N_1429,N_1219,N_1351);
and U1430 (N_1430,N_1331,N_1345);
and U1431 (N_1431,N_1294,N_1232);
nand U1432 (N_1432,N_1347,N_1311);
or U1433 (N_1433,N_1274,N_1234);
and U1434 (N_1434,N_1240,N_1248);
and U1435 (N_1435,N_1367,N_1319);
and U1436 (N_1436,N_1329,N_1301);
or U1437 (N_1437,N_1372,N_1326);
or U1438 (N_1438,N_1279,N_1205);
nor U1439 (N_1439,N_1202,N_1307);
or U1440 (N_1440,N_1288,N_1271);
or U1441 (N_1441,N_1322,N_1257);
nand U1442 (N_1442,N_1226,N_1272);
nand U1443 (N_1443,N_1385,N_1204);
and U1444 (N_1444,N_1342,N_1263);
nand U1445 (N_1445,N_1354,N_1358);
nor U1446 (N_1446,N_1353,N_1266);
or U1447 (N_1447,N_1233,N_1209);
or U1448 (N_1448,N_1324,N_1390);
nand U1449 (N_1449,N_1275,N_1224);
or U1450 (N_1450,N_1328,N_1207);
nor U1451 (N_1451,N_1384,N_1268);
and U1452 (N_1452,N_1217,N_1350);
or U1453 (N_1453,N_1298,N_1348);
or U1454 (N_1454,N_1373,N_1225);
nand U1455 (N_1455,N_1368,N_1317);
or U1456 (N_1456,N_1297,N_1315);
nor U1457 (N_1457,N_1361,N_1285);
nand U1458 (N_1458,N_1270,N_1316);
or U1459 (N_1459,N_1220,N_1338);
nand U1460 (N_1460,N_1280,N_1321);
or U1461 (N_1461,N_1293,N_1206);
nand U1462 (N_1462,N_1254,N_1289);
or U1463 (N_1463,N_1364,N_1357);
and U1464 (N_1464,N_1325,N_1269);
nor U1465 (N_1465,N_1244,N_1335);
nand U1466 (N_1466,N_1398,N_1295);
or U1467 (N_1467,N_1370,N_1313);
and U1468 (N_1468,N_1360,N_1231);
and U1469 (N_1469,N_1339,N_1276);
nor U1470 (N_1470,N_1359,N_1337);
nand U1471 (N_1471,N_1304,N_1320);
nand U1472 (N_1472,N_1375,N_1397);
nand U1473 (N_1473,N_1340,N_1223);
and U1474 (N_1474,N_1230,N_1305);
nor U1475 (N_1475,N_1296,N_1221);
and U1476 (N_1476,N_1388,N_1292);
and U1477 (N_1477,N_1262,N_1343);
nand U1478 (N_1478,N_1333,N_1250);
nand U1479 (N_1479,N_1265,N_1258);
and U1480 (N_1480,N_1235,N_1399);
nor U1481 (N_1481,N_1283,N_1259);
nor U1482 (N_1482,N_1241,N_1256);
nor U1483 (N_1483,N_1396,N_1381);
nand U1484 (N_1484,N_1392,N_1318);
nand U1485 (N_1485,N_1282,N_1302);
nor U1486 (N_1486,N_1394,N_1239);
or U1487 (N_1487,N_1314,N_1261);
and U1488 (N_1488,N_1380,N_1355);
and U1489 (N_1489,N_1327,N_1341);
and U1490 (N_1490,N_1281,N_1371);
or U1491 (N_1491,N_1201,N_1249);
and U1492 (N_1492,N_1377,N_1208);
and U1493 (N_1493,N_1284,N_1334);
nand U1494 (N_1494,N_1306,N_1379);
nor U1495 (N_1495,N_1383,N_1200);
and U1496 (N_1496,N_1203,N_1376);
nand U1497 (N_1497,N_1352,N_1238);
and U1498 (N_1498,N_1227,N_1255);
nand U1499 (N_1499,N_1336,N_1214);
or U1500 (N_1500,N_1270,N_1259);
and U1501 (N_1501,N_1383,N_1393);
nor U1502 (N_1502,N_1318,N_1281);
nand U1503 (N_1503,N_1265,N_1274);
and U1504 (N_1504,N_1212,N_1236);
nor U1505 (N_1505,N_1366,N_1330);
and U1506 (N_1506,N_1292,N_1314);
and U1507 (N_1507,N_1392,N_1233);
xnor U1508 (N_1508,N_1236,N_1323);
and U1509 (N_1509,N_1218,N_1214);
or U1510 (N_1510,N_1334,N_1296);
nor U1511 (N_1511,N_1225,N_1340);
nand U1512 (N_1512,N_1207,N_1343);
or U1513 (N_1513,N_1313,N_1270);
or U1514 (N_1514,N_1212,N_1387);
nand U1515 (N_1515,N_1343,N_1220);
nor U1516 (N_1516,N_1285,N_1380);
nand U1517 (N_1517,N_1326,N_1267);
nand U1518 (N_1518,N_1237,N_1211);
or U1519 (N_1519,N_1266,N_1276);
xor U1520 (N_1520,N_1321,N_1233);
and U1521 (N_1521,N_1340,N_1302);
xnor U1522 (N_1522,N_1217,N_1336);
nand U1523 (N_1523,N_1229,N_1323);
or U1524 (N_1524,N_1275,N_1360);
nand U1525 (N_1525,N_1215,N_1277);
nor U1526 (N_1526,N_1376,N_1244);
nand U1527 (N_1527,N_1270,N_1307);
or U1528 (N_1528,N_1226,N_1387);
and U1529 (N_1529,N_1320,N_1352);
and U1530 (N_1530,N_1237,N_1372);
and U1531 (N_1531,N_1232,N_1288);
nor U1532 (N_1532,N_1237,N_1359);
nor U1533 (N_1533,N_1336,N_1250);
or U1534 (N_1534,N_1232,N_1279);
or U1535 (N_1535,N_1264,N_1311);
nand U1536 (N_1536,N_1227,N_1376);
nor U1537 (N_1537,N_1272,N_1294);
xor U1538 (N_1538,N_1371,N_1241);
nand U1539 (N_1539,N_1345,N_1395);
and U1540 (N_1540,N_1295,N_1247);
nand U1541 (N_1541,N_1310,N_1374);
or U1542 (N_1542,N_1338,N_1297);
or U1543 (N_1543,N_1364,N_1283);
or U1544 (N_1544,N_1230,N_1321);
nand U1545 (N_1545,N_1368,N_1259);
and U1546 (N_1546,N_1249,N_1362);
nor U1547 (N_1547,N_1234,N_1303);
nor U1548 (N_1548,N_1274,N_1295);
and U1549 (N_1549,N_1286,N_1283);
and U1550 (N_1550,N_1207,N_1221);
nor U1551 (N_1551,N_1251,N_1336);
or U1552 (N_1552,N_1363,N_1241);
or U1553 (N_1553,N_1316,N_1393);
or U1554 (N_1554,N_1307,N_1364);
and U1555 (N_1555,N_1362,N_1349);
and U1556 (N_1556,N_1346,N_1238);
nand U1557 (N_1557,N_1362,N_1286);
nor U1558 (N_1558,N_1277,N_1308);
or U1559 (N_1559,N_1282,N_1232);
xnor U1560 (N_1560,N_1250,N_1342);
nor U1561 (N_1561,N_1376,N_1272);
xnor U1562 (N_1562,N_1332,N_1364);
nor U1563 (N_1563,N_1319,N_1281);
and U1564 (N_1564,N_1337,N_1221);
and U1565 (N_1565,N_1360,N_1349);
nand U1566 (N_1566,N_1265,N_1350);
nor U1567 (N_1567,N_1229,N_1236);
nor U1568 (N_1568,N_1256,N_1331);
xnor U1569 (N_1569,N_1307,N_1387);
nor U1570 (N_1570,N_1268,N_1361);
nor U1571 (N_1571,N_1382,N_1278);
and U1572 (N_1572,N_1242,N_1214);
or U1573 (N_1573,N_1214,N_1384);
and U1574 (N_1574,N_1381,N_1218);
nand U1575 (N_1575,N_1313,N_1205);
nand U1576 (N_1576,N_1287,N_1242);
nand U1577 (N_1577,N_1354,N_1316);
and U1578 (N_1578,N_1371,N_1229);
nor U1579 (N_1579,N_1352,N_1294);
or U1580 (N_1580,N_1229,N_1277);
or U1581 (N_1581,N_1309,N_1396);
nor U1582 (N_1582,N_1237,N_1242);
and U1583 (N_1583,N_1358,N_1374);
nand U1584 (N_1584,N_1261,N_1342);
nor U1585 (N_1585,N_1386,N_1363);
nand U1586 (N_1586,N_1242,N_1352);
or U1587 (N_1587,N_1283,N_1353);
and U1588 (N_1588,N_1216,N_1201);
nor U1589 (N_1589,N_1328,N_1271);
xor U1590 (N_1590,N_1342,N_1270);
nand U1591 (N_1591,N_1221,N_1318);
and U1592 (N_1592,N_1289,N_1300);
or U1593 (N_1593,N_1278,N_1211);
or U1594 (N_1594,N_1310,N_1203);
nand U1595 (N_1595,N_1322,N_1294);
nand U1596 (N_1596,N_1224,N_1271);
or U1597 (N_1597,N_1236,N_1226);
nand U1598 (N_1598,N_1291,N_1250);
or U1599 (N_1599,N_1261,N_1396);
nand U1600 (N_1600,N_1591,N_1558);
nor U1601 (N_1601,N_1475,N_1574);
nor U1602 (N_1602,N_1585,N_1433);
and U1603 (N_1603,N_1445,N_1427);
nand U1604 (N_1604,N_1476,N_1536);
nand U1605 (N_1605,N_1509,N_1417);
xor U1606 (N_1606,N_1401,N_1527);
nand U1607 (N_1607,N_1500,N_1549);
or U1608 (N_1608,N_1537,N_1529);
nor U1609 (N_1609,N_1485,N_1424);
and U1610 (N_1610,N_1598,N_1520);
nand U1611 (N_1611,N_1579,N_1566);
and U1612 (N_1612,N_1588,N_1457);
or U1613 (N_1613,N_1434,N_1564);
nand U1614 (N_1614,N_1420,N_1575);
xnor U1615 (N_1615,N_1451,N_1590);
nand U1616 (N_1616,N_1543,N_1547);
nand U1617 (N_1617,N_1493,N_1593);
nor U1618 (N_1618,N_1405,N_1570);
nand U1619 (N_1619,N_1435,N_1453);
nand U1620 (N_1620,N_1511,N_1423);
nor U1621 (N_1621,N_1463,N_1545);
nor U1622 (N_1622,N_1583,N_1592);
and U1623 (N_1623,N_1525,N_1496);
nor U1624 (N_1624,N_1490,N_1473);
nand U1625 (N_1625,N_1440,N_1554);
nand U1626 (N_1626,N_1444,N_1548);
and U1627 (N_1627,N_1404,N_1594);
and U1628 (N_1628,N_1409,N_1430);
or U1629 (N_1629,N_1526,N_1540);
and U1630 (N_1630,N_1534,N_1448);
nor U1631 (N_1631,N_1582,N_1449);
and U1632 (N_1632,N_1516,N_1524);
or U1633 (N_1633,N_1481,N_1474);
nor U1634 (N_1634,N_1480,N_1429);
or U1635 (N_1635,N_1452,N_1454);
or U1636 (N_1636,N_1519,N_1572);
nor U1637 (N_1637,N_1568,N_1421);
or U1638 (N_1638,N_1542,N_1479);
or U1639 (N_1639,N_1502,N_1556);
or U1640 (N_1640,N_1415,N_1400);
or U1641 (N_1641,N_1486,N_1467);
or U1642 (N_1642,N_1447,N_1406);
nor U1643 (N_1643,N_1470,N_1532);
and U1644 (N_1644,N_1505,N_1407);
nor U1645 (N_1645,N_1541,N_1513);
or U1646 (N_1646,N_1498,N_1472);
and U1647 (N_1647,N_1555,N_1563);
nor U1648 (N_1648,N_1517,N_1597);
or U1649 (N_1649,N_1512,N_1422);
or U1650 (N_1650,N_1408,N_1497);
and U1651 (N_1651,N_1441,N_1521);
or U1652 (N_1652,N_1494,N_1403);
and U1653 (N_1653,N_1455,N_1514);
xnor U1654 (N_1654,N_1539,N_1478);
nand U1655 (N_1655,N_1468,N_1495);
nor U1656 (N_1656,N_1567,N_1425);
nand U1657 (N_1657,N_1442,N_1553);
nand U1658 (N_1658,N_1589,N_1487);
or U1659 (N_1659,N_1535,N_1544);
or U1660 (N_1660,N_1464,N_1414);
or U1661 (N_1661,N_1483,N_1416);
nand U1662 (N_1662,N_1492,N_1489);
nor U1663 (N_1663,N_1538,N_1462);
nor U1664 (N_1664,N_1561,N_1569);
nor U1665 (N_1665,N_1531,N_1507);
nor U1666 (N_1666,N_1431,N_1595);
and U1667 (N_1667,N_1508,N_1411);
nand U1668 (N_1668,N_1458,N_1584);
nand U1669 (N_1669,N_1410,N_1576);
nand U1670 (N_1670,N_1501,N_1402);
nor U1671 (N_1671,N_1565,N_1426);
nor U1672 (N_1672,N_1523,N_1438);
or U1673 (N_1673,N_1587,N_1586);
nor U1674 (N_1674,N_1412,N_1436);
nand U1675 (N_1675,N_1450,N_1581);
nor U1676 (N_1676,N_1506,N_1552);
and U1677 (N_1677,N_1499,N_1491);
nand U1678 (N_1678,N_1530,N_1466);
nor U1679 (N_1679,N_1459,N_1546);
and U1680 (N_1680,N_1557,N_1469);
and U1681 (N_1681,N_1419,N_1428);
or U1682 (N_1682,N_1456,N_1443);
nor U1683 (N_1683,N_1432,N_1518);
nor U1684 (N_1684,N_1533,N_1599);
or U1685 (N_1685,N_1580,N_1488);
and U1686 (N_1686,N_1504,N_1573);
nand U1687 (N_1687,N_1446,N_1515);
or U1688 (N_1688,N_1503,N_1577);
or U1689 (N_1689,N_1437,N_1439);
or U1690 (N_1690,N_1482,N_1461);
or U1691 (N_1691,N_1559,N_1528);
or U1692 (N_1692,N_1562,N_1484);
or U1693 (N_1693,N_1596,N_1578);
or U1694 (N_1694,N_1571,N_1413);
or U1695 (N_1695,N_1465,N_1551);
and U1696 (N_1696,N_1550,N_1560);
nand U1697 (N_1697,N_1418,N_1522);
and U1698 (N_1698,N_1477,N_1471);
or U1699 (N_1699,N_1460,N_1510);
and U1700 (N_1700,N_1563,N_1549);
xor U1701 (N_1701,N_1549,N_1447);
nand U1702 (N_1702,N_1570,N_1540);
or U1703 (N_1703,N_1525,N_1492);
nand U1704 (N_1704,N_1490,N_1595);
or U1705 (N_1705,N_1478,N_1565);
or U1706 (N_1706,N_1417,N_1562);
and U1707 (N_1707,N_1467,N_1543);
nand U1708 (N_1708,N_1499,N_1500);
nor U1709 (N_1709,N_1559,N_1490);
nand U1710 (N_1710,N_1438,N_1518);
nand U1711 (N_1711,N_1424,N_1562);
and U1712 (N_1712,N_1413,N_1548);
nand U1713 (N_1713,N_1513,N_1423);
nor U1714 (N_1714,N_1475,N_1497);
and U1715 (N_1715,N_1584,N_1530);
nor U1716 (N_1716,N_1514,N_1499);
or U1717 (N_1717,N_1414,N_1499);
or U1718 (N_1718,N_1439,N_1412);
and U1719 (N_1719,N_1423,N_1443);
nor U1720 (N_1720,N_1524,N_1491);
or U1721 (N_1721,N_1405,N_1564);
nand U1722 (N_1722,N_1513,N_1481);
or U1723 (N_1723,N_1468,N_1528);
nand U1724 (N_1724,N_1402,N_1464);
nor U1725 (N_1725,N_1560,N_1419);
nand U1726 (N_1726,N_1441,N_1589);
nor U1727 (N_1727,N_1471,N_1534);
nand U1728 (N_1728,N_1497,N_1569);
and U1729 (N_1729,N_1408,N_1487);
nor U1730 (N_1730,N_1447,N_1477);
nand U1731 (N_1731,N_1452,N_1515);
nor U1732 (N_1732,N_1484,N_1437);
or U1733 (N_1733,N_1400,N_1580);
or U1734 (N_1734,N_1525,N_1592);
and U1735 (N_1735,N_1554,N_1588);
nor U1736 (N_1736,N_1598,N_1490);
nand U1737 (N_1737,N_1501,N_1422);
or U1738 (N_1738,N_1402,N_1578);
nand U1739 (N_1739,N_1482,N_1455);
nor U1740 (N_1740,N_1510,N_1501);
nor U1741 (N_1741,N_1443,N_1451);
and U1742 (N_1742,N_1575,N_1464);
and U1743 (N_1743,N_1544,N_1572);
nor U1744 (N_1744,N_1567,N_1516);
and U1745 (N_1745,N_1473,N_1425);
or U1746 (N_1746,N_1451,N_1437);
nor U1747 (N_1747,N_1575,N_1467);
or U1748 (N_1748,N_1421,N_1486);
nand U1749 (N_1749,N_1533,N_1493);
nand U1750 (N_1750,N_1422,N_1576);
nor U1751 (N_1751,N_1425,N_1453);
nor U1752 (N_1752,N_1536,N_1540);
nand U1753 (N_1753,N_1480,N_1414);
and U1754 (N_1754,N_1489,N_1584);
or U1755 (N_1755,N_1414,N_1596);
and U1756 (N_1756,N_1451,N_1576);
nor U1757 (N_1757,N_1422,N_1464);
and U1758 (N_1758,N_1474,N_1468);
and U1759 (N_1759,N_1487,N_1426);
nand U1760 (N_1760,N_1584,N_1515);
and U1761 (N_1761,N_1482,N_1402);
and U1762 (N_1762,N_1506,N_1581);
and U1763 (N_1763,N_1560,N_1555);
and U1764 (N_1764,N_1494,N_1564);
nor U1765 (N_1765,N_1441,N_1536);
and U1766 (N_1766,N_1587,N_1452);
or U1767 (N_1767,N_1553,N_1482);
nor U1768 (N_1768,N_1549,N_1543);
or U1769 (N_1769,N_1406,N_1474);
or U1770 (N_1770,N_1428,N_1512);
nand U1771 (N_1771,N_1418,N_1415);
nand U1772 (N_1772,N_1432,N_1439);
nor U1773 (N_1773,N_1491,N_1408);
nor U1774 (N_1774,N_1528,N_1527);
and U1775 (N_1775,N_1433,N_1431);
or U1776 (N_1776,N_1529,N_1594);
nand U1777 (N_1777,N_1596,N_1446);
or U1778 (N_1778,N_1518,N_1408);
nand U1779 (N_1779,N_1514,N_1474);
or U1780 (N_1780,N_1484,N_1440);
nand U1781 (N_1781,N_1553,N_1588);
or U1782 (N_1782,N_1489,N_1408);
or U1783 (N_1783,N_1503,N_1476);
and U1784 (N_1784,N_1462,N_1571);
nand U1785 (N_1785,N_1572,N_1531);
and U1786 (N_1786,N_1431,N_1537);
and U1787 (N_1787,N_1466,N_1417);
and U1788 (N_1788,N_1574,N_1430);
nor U1789 (N_1789,N_1520,N_1416);
nor U1790 (N_1790,N_1403,N_1446);
or U1791 (N_1791,N_1415,N_1580);
xnor U1792 (N_1792,N_1577,N_1582);
nor U1793 (N_1793,N_1599,N_1455);
nand U1794 (N_1794,N_1535,N_1411);
nor U1795 (N_1795,N_1585,N_1422);
and U1796 (N_1796,N_1498,N_1453);
nor U1797 (N_1797,N_1447,N_1485);
and U1798 (N_1798,N_1405,N_1530);
nand U1799 (N_1799,N_1501,N_1436);
and U1800 (N_1800,N_1601,N_1716);
nor U1801 (N_1801,N_1723,N_1640);
or U1802 (N_1802,N_1791,N_1693);
nand U1803 (N_1803,N_1798,N_1797);
nand U1804 (N_1804,N_1764,N_1769);
or U1805 (N_1805,N_1712,N_1661);
and U1806 (N_1806,N_1653,N_1650);
nor U1807 (N_1807,N_1702,N_1708);
and U1808 (N_1808,N_1608,N_1612);
or U1809 (N_1809,N_1799,N_1795);
nor U1810 (N_1810,N_1753,N_1613);
or U1811 (N_1811,N_1666,N_1718);
or U1812 (N_1812,N_1629,N_1768);
or U1813 (N_1813,N_1647,N_1634);
and U1814 (N_1814,N_1743,N_1686);
and U1815 (N_1815,N_1742,N_1618);
nand U1816 (N_1816,N_1658,N_1733);
and U1817 (N_1817,N_1793,N_1725);
or U1818 (N_1818,N_1651,N_1739);
or U1819 (N_1819,N_1681,N_1737);
and U1820 (N_1820,N_1638,N_1731);
nand U1821 (N_1821,N_1636,N_1679);
and U1822 (N_1822,N_1747,N_1691);
nor U1823 (N_1823,N_1602,N_1694);
or U1824 (N_1824,N_1677,N_1687);
nand U1825 (N_1825,N_1690,N_1751);
nand U1826 (N_1826,N_1724,N_1709);
nand U1827 (N_1827,N_1748,N_1741);
or U1828 (N_1828,N_1643,N_1667);
nor U1829 (N_1829,N_1727,N_1683);
and U1830 (N_1830,N_1624,N_1635);
or U1831 (N_1831,N_1715,N_1639);
nand U1832 (N_1832,N_1784,N_1621);
and U1833 (N_1833,N_1755,N_1663);
or U1834 (N_1834,N_1730,N_1657);
and U1835 (N_1835,N_1785,N_1699);
nand U1836 (N_1836,N_1756,N_1628);
and U1837 (N_1837,N_1631,N_1622);
nand U1838 (N_1838,N_1705,N_1703);
or U1839 (N_1839,N_1692,N_1761);
or U1840 (N_1840,N_1777,N_1706);
nand U1841 (N_1841,N_1788,N_1668);
nand U1842 (N_1842,N_1776,N_1728);
and U1843 (N_1843,N_1675,N_1664);
nor U1844 (N_1844,N_1637,N_1645);
or U1845 (N_1845,N_1646,N_1732);
or U1846 (N_1846,N_1685,N_1611);
nor U1847 (N_1847,N_1656,N_1654);
and U1848 (N_1848,N_1700,N_1697);
nor U1849 (N_1849,N_1746,N_1772);
or U1850 (N_1850,N_1678,N_1696);
or U1851 (N_1851,N_1662,N_1794);
nand U1852 (N_1852,N_1680,N_1620);
and U1853 (N_1853,N_1649,N_1787);
nor U1854 (N_1854,N_1790,N_1779);
and U1855 (N_1855,N_1786,N_1606);
nand U1856 (N_1856,N_1676,N_1695);
and U1857 (N_1857,N_1641,N_1757);
nor U1858 (N_1858,N_1609,N_1762);
and U1859 (N_1859,N_1758,N_1783);
or U1860 (N_1860,N_1615,N_1669);
nand U1861 (N_1861,N_1735,N_1754);
nor U1862 (N_1862,N_1796,N_1774);
nor U1863 (N_1863,N_1689,N_1648);
and U1864 (N_1864,N_1672,N_1642);
nand U1865 (N_1865,N_1652,N_1660);
nor U1866 (N_1866,N_1770,N_1750);
nand U1867 (N_1867,N_1632,N_1633);
and U1868 (N_1868,N_1720,N_1603);
or U1869 (N_1869,N_1710,N_1734);
and U1870 (N_1870,N_1736,N_1607);
and U1871 (N_1871,N_1729,N_1665);
nand U1872 (N_1872,N_1738,N_1616);
nor U1873 (N_1873,N_1759,N_1673);
nor U1874 (N_1874,N_1684,N_1614);
nor U1875 (N_1875,N_1711,N_1604);
nor U1876 (N_1876,N_1659,N_1745);
and U1877 (N_1877,N_1780,N_1771);
or U1878 (N_1878,N_1655,N_1688);
nand U1879 (N_1879,N_1627,N_1671);
and U1880 (N_1880,N_1717,N_1752);
nand U1881 (N_1881,N_1701,N_1674);
xor U1882 (N_1882,N_1778,N_1781);
nand U1883 (N_1883,N_1792,N_1617);
nand U1884 (N_1884,N_1726,N_1744);
nor U1885 (N_1885,N_1714,N_1719);
nor U1886 (N_1886,N_1789,N_1707);
nor U1887 (N_1887,N_1749,N_1722);
or U1888 (N_1888,N_1630,N_1760);
nor U1889 (N_1889,N_1765,N_1625);
or U1890 (N_1890,N_1704,N_1766);
and U1891 (N_1891,N_1782,N_1767);
nor U1892 (N_1892,N_1682,N_1763);
nor U1893 (N_1893,N_1619,N_1626);
nand U1894 (N_1894,N_1721,N_1698);
and U1895 (N_1895,N_1740,N_1713);
nor U1896 (N_1896,N_1670,N_1775);
xor U1897 (N_1897,N_1610,N_1605);
and U1898 (N_1898,N_1773,N_1600);
nor U1899 (N_1899,N_1623,N_1644);
and U1900 (N_1900,N_1741,N_1618);
and U1901 (N_1901,N_1688,N_1784);
nand U1902 (N_1902,N_1794,N_1730);
and U1903 (N_1903,N_1774,N_1736);
nor U1904 (N_1904,N_1743,N_1632);
and U1905 (N_1905,N_1724,N_1644);
xor U1906 (N_1906,N_1764,N_1757);
nand U1907 (N_1907,N_1709,N_1720);
or U1908 (N_1908,N_1652,N_1621);
nand U1909 (N_1909,N_1739,N_1645);
nor U1910 (N_1910,N_1789,N_1791);
nand U1911 (N_1911,N_1750,N_1683);
and U1912 (N_1912,N_1605,N_1755);
or U1913 (N_1913,N_1664,N_1711);
or U1914 (N_1914,N_1680,N_1761);
nand U1915 (N_1915,N_1764,N_1784);
and U1916 (N_1916,N_1714,N_1765);
nand U1917 (N_1917,N_1735,N_1678);
nand U1918 (N_1918,N_1760,N_1715);
nand U1919 (N_1919,N_1611,N_1645);
nor U1920 (N_1920,N_1624,N_1799);
or U1921 (N_1921,N_1772,N_1663);
nand U1922 (N_1922,N_1777,N_1633);
and U1923 (N_1923,N_1636,N_1781);
nand U1924 (N_1924,N_1645,N_1765);
nand U1925 (N_1925,N_1703,N_1748);
nor U1926 (N_1926,N_1723,N_1771);
nand U1927 (N_1927,N_1798,N_1778);
nand U1928 (N_1928,N_1721,N_1705);
xor U1929 (N_1929,N_1607,N_1721);
or U1930 (N_1930,N_1785,N_1731);
and U1931 (N_1931,N_1766,N_1646);
or U1932 (N_1932,N_1641,N_1753);
and U1933 (N_1933,N_1695,N_1696);
nand U1934 (N_1934,N_1798,N_1630);
and U1935 (N_1935,N_1782,N_1681);
or U1936 (N_1936,N_1647,N_1749);
or U1937 (N_1937,N_1634,N_1669);
nand U1938 (N_1938,N_1678,N_1729);
nand U1939 (N_1939,N_1796,N_1792);
and U1940 (N_1940,N_1715,N_1651);
and U1941 (N_1941,N_1622,N_1662);
xnor U1942 (N_1942,N_1619,N_1760);
and U1943 (N_1943,N_1600,N_1659);
nor U1944 (N_1944,N_1782,N_1716);
nor U1945 (N_1945,N_1713,N_1651);
nand U1946 (N_1946,N_1614,N_1603);
nand U1947 (N_1947,N_1610,N_1701);
nor U1948 (N_1948,N_1698,N_1729);
or U1949 (N_1949,N_1772,N_1676);
and U1950 (N_1950,N_1603,N_1705);
or U1951 (N_1951,N_1650,N_1664);
or U1952 (N_1952,N_1699,N_1744);
or U1953 (N_1953,N_1609,N_1606);
nand U1954 (N_1954,N_1711,N_1723);
nor U1955 (N_1955,N_1653,N_1785);
or U1956 (N_1956,N_1783,N_1784);
nand U1957 (N_1957,N_1693,N_1729);
nor U1958 (N_1958,N_1631,N_1744);
nand U1959 (N_1959,N_1725,N_1605);
xnor U1960 (N_1960,N_1797,N_1648);
and U1961 (N_1961,N_1799,N_1676);
nand U1962 (N_1962,N_1699,N_1628);
nor U1963 (N_1963,N_1694,N_1615);
nor U1964 (N_1964,N_1752,N_1664);
nand U1965 (N_1965,N_1686,N_1766);
or U1966 (N_1966,N_1637,N_1708);
and U1967 (N_1967,N_1710,N_1685);
nor U1968 (N_1968,N_1755,N_1666);
or U1969 (N_1969,N_1757,N_1710);
nor U1970 (N_1970,N_1620,N_1763);
or U1971 (N_1971,N_1769,N_1693);
and U1972 (N_1972,N_1771,N_1642);
nor U1973 (N_1973,N_1676,N_1651);
nand U1974 (N_1974,N_1759,N_1687);
and U1975 (N_1975,N_1681,N_1711);
nand U1976 (N_1976,N_1689,N_1727);
and U1977 (N_1977,N_1726,N_1661);
or U1978 (N_1978,N_1672,N_1770);
and U1979 (N_1979,N_1664,N_1682);
and U1980 (N_1980,N_1621,N_1794);
nand U1981 (N_1981,N_1600,N_1717);
or U1982 (N_1982,N_1773,N_1632);
and U1983 (N_1983,N_1744,N_1785);
or U1984 (N_1984,N_1762,N_1765);
nor U1985 (N_1985,N_1642,N_1640);
nor U1986 (N_1986,N_1698,N_1746);
nor U1987 (N_1987,N_1785,N_1769);
nor U1988 (N_1988,N_1764,N_1688);
nor U1989 (N_1989,N_1701,N_1692);
or U1990 (N_1990,N_1651,N_1722);
nand U1991 (N_1991,N_1701,N_1739);
and U1992 (N_1992,N_1767,N_1737);
nand U1993 (N_1993,N_1706,N_1621);
nor U1994 (N_1994,N_1782,N_1694);
and U1995 (N_1995,N_1734,N_1661);
nor U1996 (N_1996,N_1722,N_1778);
nand U1997 (N_1997,N_1748,N_1763);
or U1998 (N_1998,N_1730,N_1718);
or U1999 (N_1999,N_1688,N_1711);
nor U2000 (N_2000,N_1845,N_1991);
nor U2001 (N_2001,N_1866,N_1958);
or U2002 (N_2002,N_1922,N_1835);
nand U2003 (N_2003,N_1888,N_1996);
or U2004 (N_2004,N_1880,N_1803);
and U2005 (N_2005,N_1965,N_1911);
or U2006 (N_2006,N_1993,N_1893);
and U2007 (N_2007,N_1907,N_1906);
and U2008 (N_2008,N_1817,N_1925);
and U2009 (N_2009,N_1995,N_1889);
nand U2010 (N_2010,N_1920,N_1836);
or U2011 (N_2011,N_1820,N_1834);
nor U2012 (N_2012,N_1840,N_1932);
nor U2013 (N_2013,N_1942,N_1884);
nand U2014 (N_2014,N_1927,N_1998);
and U2015 (N_2015,N_1939,N_1864);
nor U2016 (N_2016,N_1908,N_1838);
or U2017 (N_2017,N_1807,N_1854);
and U2018 (N_2018,N_1897,N_1941);
nand U2019 (N_2019,N_1881,N_1848);
or U2020 (N_2020,N_1891,N_1956);
or U2021 (N_2021,N_1940,N_1858);
or U2022 (N_2022,N_1978,N_1861);
nor U2023 (N_2023,N_1987,N_1806);
nor U2024 (N_2024,N_1930,N_1938);
nand U2025 (N_2025,N_1839,N_1819);
nand U2026 (N_2026,N_1808,N_1842);
and U2027 (N_2027,N_1865,N_1831);
nand U2028 (N_2028,N_1997,N_1871);
and U2029 (N_2029,N_1933,N_1830);
nor U2030 (N_2030,N_1989,N_1900);
nor U2031 (N_2031,N_1878,N_1915);
and U2032 (N_2032,N_1948,N_1802);
nand U2033 (N_2033,N_1928,N_1818);
nor U2034 (N_2034,N_1877,N_1868);
or U2035 (N_2035,N_1847,N_1981);
nand U2036 (N_2036,N_1971,N_1916);
nand U2037 (N_2037,N_1859,N_1934);
or U2038 (N_2038,N_1990,N_1999);
and U2039 (N_2039,N_1918,N_1936);
and U2040 (N_2040,N_1944,N_1849);
and U2041 (N_2041,N_1821,N_1811);
and U2042 (N_2042,N_1919,N_1954);
and U2043 (N_2043,N_1872,N_1892);
nand U2044 (N_2044,N_1822,N_1975);
or U2045 (N_2045,N_1825,N_1979);
xnor U2046 (N_2046,N_1853,N_1909);
nor U2047 (N_2047,N_1984,N_1846);
nand U2048 (N_2048,N_1823,N_1955);
nand U2049 (N_2049,N_1976,N_1982);
or U2050 (N_2050,N_1945,N_1994);
and U2051 (N_2051,N_1968,N_1953);
or U2052 (N_2052,N_1841,N_1829);
nand U2053 (N_2053,N_1901,N_1857);
and U2054 (N_2054,N_1950,N_1809);
nand U2055 (N_2055,N_1812,N_1905);
nor U2056 (N_2056,N_1910,N_1876);
nor U2057 (N_2057,N_1903,N_1816);
nand U2058 (N_2058,N_1894,N_1960);
and U2059 (N_2059,N_1924,N_1935);
nand U2060 (N_2060,N_1844,N_1959);
nand U2061 (N_2061,N_1988,N_1804);
and U2062 (N_2062,N_1862,N_1828);
nand U2063 (N_2063,N_1929,N_1837);
nand U2064 (N_2064,N_1923,N_1867);
and U2065 (N_2065,N_1921,N_1969);
or U2066 (N_2066,N_1813,N_1885);
nor U2067 (N_2067,N_1850,N_1937);
nor U2068 (N_2068,N_1967,N_1952);
nor U2069 (N_2069,N_1814,N_1869);
nand U2070 (N_2070,N_1824,N_1800);
nand U2071 (N_2071,N_1801,N_1805);
nand U2072 (N_2072,N_1832,N_1947);
nor U2073 (N_2073,N_1943,N_1826);
or U2074 (N_2074,N_1873,N_1972);
nand U2075 (N_2075,N_1896,N_1833);
nand U2076 (N_2076,N_1913,N_1875);
and U2077 (N_2077,N_1904,N_1856);
or U2078 (N_2078,N_1827,N_1946);
nor U2079 (N_2079,N_1986,N_1902);
or U2080 (N_2080,N_1912,N_1970);
and U2081 (N_2081,N_1964,N_1926);
or U2082 (N_2082,N_1957,N_1863);
nand U2083 (N_2083,N_1874,N_1882);
nor U2084 (N_2084,N_1961,N_1898);
nor U2085 (N_2085,N_1815,N_1931);
nor U2086 (N_2086,N_1886,N_1977);
or U2087 (N_2087,N_1879,N_1852);
or U2088 (N_2088,N_1895,N_1974);
nand U2089 (N_2089,N_1951,N_1992);
or U2090 (N_2090,N_1890,N_1883);
and U2091 (N_2091,N_1949,N_1810);
or U2092 (N_2092,N_1914,N_1851);
nand U2093 (N_2093,N_1843,N_1917);
and U2094 (N_2094,N_1899,N_1980);
or U2095 (N_2095,N_1966,N_1962);
nand U2096 (N_2096,N_1963,N_1973);
and U2097 (N_2097,N_1887,N_1855);
nand U2098 (N_2098,N_1983,N_1985);
nor U2099 (N_2099,N_1870,N_1860);
nor U2100 (N_2100,N_1830,N_1952);
and U2101 (N_2101,N_1986,N_1894);
nand U2102 (N_2102,N_1953,N_1983);
nand U2103 (N_2103,N_1956,N_1912);
nand U2104 (N_2104,N_1851,N_1854);
or U2105 (N_2105,N_1812,N_1945);
nor U2106 (N_2106,N_1815,N_1969);
and U2107 (N_2107,N_1972,N_1979);
or U2108 (N_2108,N_1814,N_1895);
or U2109 (N_2109,N_1828,N_1810);
and U2110 (N_2110,N_1982,N_1858);
nand U2111 (N_2111,N_1956,N_1887);
nand U2112 (N_2112,N_1937,N_1941);
or U2113 (N_2113,N_1933,N_1993);
nand U2114 (N_2114,N_1874,N_1880);
nand U2115 (N_2115,N_1964,N_1803);
nand U2116 (N_2116,N_1994,N_1926);
and U2117 (N_2117,N_1858,N_1948);
nor U2118 (N_2118,N_1909,N_1990);
or U2119 (N_2119,N_1964,N_1921);
and U2120 (N_2120,N_1833,N_1882);
nor U2121 (N_2121,N_1898,N_1945);
nand U2122 (N_2122,N_1861,N_1859);
nor U2123 (N_2123,N_1868,N_1841);
and U2124 (N_2124,N_1969,N_1877);
and U2125 (N_2125,N_1874,N_1998);
nor U2126 (N_2126,N_1992,N_1817);
nor U2127 (N_2127,N_1821,N_1932);
and U2128 (N_2128,N_1912,N_1961);
nand U2129 (N_2129,N_1829,N_1974);
and U2130 (N_2130,N_1905,N_1975);
nand U2131 (N_2131,N_1994,N_1904);
xnor U2132 (N_2132,N_1982,N_1964);
and U2133 (N_2133,N_1879,N_1806);
or U2134 (N_2134,N_1968,N_1806);
nand U2135 (N_2135,N_1804,N_1921);
and U2136 (N_2136,N_1803,N_1875);
nand U2137 (N_2137,N_1884,N_1899);
or U2138 (N_2138,N_1874,N_1961);
nand U2139 (N_2139,N_1949,N_1858);
and U2140 (N_2140,N_1988,N_1976);
and U2141 (N_2141,N_1883,N_1956);
nand U2142 (N_2142,N_1842,N_1911);
nand U2143 (N_2143,N_1951,N_1837);
nor U2144 (N_2144,N_1877,N_1944);
nor U2145 (N_2145,N_1915,N_1917);
or U2146 (N_2146,N_1874,N_1994);
nand U2147 (N_2147,N_1970,N_1965);
nand U2148 (N_2148,N_1838,N_1949);
or U2149 (N_2149,N_1847,N_1997);
nor U2150 (N_2150,N_1938,N_1848);
nor U2151 (N_2151,N_1835,N_1980);
or U2152 (N_2152,N_1917,N_1853);
and U2153 (N_2153,N_1897,N_1831);
and U2154 (N_2154,N_1952,N_1954);
nor U2155 (N_2155,N_1897,N_1866);
or U2156 (N_2156,N_1989,N_1821);
nand U2157 (N_2157,N_1800,N_1857);
nor U2158 (N_2158,N_1825,N_1896);
and U2159 (N_2159,N_1842,N_1891);
or U2160 (N_2160,N_1808,N_1945);
or U2161 (N_2161,N_1899,N_1922);
nand U2162 (N_2162,N_1864,N_1899);
nand U2163 (N_2163,N_1829,N_1925);
nand U2164 (N_2164,N_1904,N_1907);
or U2165 (N_2165,N_1866,N_1850);
or U2166 (N_2166,N_1980,N_1868);
nor U2167 (N_2167,N_1822,N_1840);
or U2168 (N_2168,N_1931,N_1857);
nor U2169 (N_2169,N_1873,N_1984);
nor U2170 (N_2170,N_1908,N_1804);
and U2171 (N_2171,N_1800,N_1981);
xnor U2172 (N_2172,N_1963,N_1965);
and U2173 (N_2173,N_1835,N_1940);
or U2174 (N_2174,N_1939,N_1849);
nor U2175 (N_2175,N_1984,N_1980);
or U2176 (N_2176,N_1867,N_1801);
and U2177 (N_2177,N_1997,N_1970);
or U2178 (N_2178,N_1858,N_1826);
or U2179 (N_2179,N_1972,N_1916);
nor U2180 (N_2180,N_1939,N_1968);
and U2181 (N_2181,N_1962,N_1827);
or U2182 (N_2182,N_1911,N_1981);
or U2183 (N_2183,N_1959,N_1833);
nand U2184 (N_2184,N_1984,N_1928);
nand U2185 (N_2185,N_1905,N_1963);
xor U2186 (N_2186,N_1933,N_1960);
nor U2187 (N_2187,N_1904,N_1932);
nand U2188 (N_2188,N_1918,N_1955);
or U2189 (N_2189,N_1991,N_1803);
or U2190 (N_2190,N_1915,N_1885);
nand U2191 (N_2191,N_1821,N_1976);
and U2192 (N_2192,N_1912,N_1847);
nor U2193 (N_2193,N_1863,N_1948);
nand U2194 (N_2194,N_1838,N_1973);
or U2195 (N_2195,N_1822,N_1823);
and U2196 (N_2196,N_1930,N_1913);
nor U2197 (N_2197,N_1817,N_1880);
or U2198 (N_2198,N_1992,N_1988);
nor U2199 (N_2199,N_1988,N_1862);
nor U2200 (N_2200,N_2054,N_2180);
and U2201 (N_2201,N_2135,N_2134);
xor U2202 (N_2202,N_2048,N_2116);
xnor U2203 (N_2203,N_2169,N_2042);
nor U2204 (N_2204,N_2035,N_2174);
or U2205 (N_2205,N_2052,N_2003);
nor U2206 (N_2206,N_2165,N_2000);
nand U2207 (N_2207,N_2031,N_2027);
and U2208 (N_2208,N_2160,N_2198);
and U2209 (N_2209,N_2190,N_2058);
or U2210 (N_2210,N_2140,N_2087);
and U2211 (N_2211,N_2127,N_2094);
nor U2212 (N_2212,N_2005,N_2168);
or U2213 (N_2213,N_2059,N_2008);
nor U2214 (N_2214,N_2050,N_2150);
xnor U2215 (N_2215,N_2046,N_2018);
nand U2216 (N_2216,N_2128,N_2184);
nor U2217 (N_2217,N_2117,N_2104);
nand U2218 (N_2218,N_2107,N_2191);
or U2219 (N_2219,N_2033,N_2110);
nor U2220 (N_2220,N_2171,N_2179);
or U2221 (N_2221,N_2068,N_2075);
nor U2222 (N_2222,N_2113,N_2026);
nand U2223 (N_2223,N_2044,N_2152);
nand U2224 (N_2224,N_2125,N_2072);
or U2225 (N_2225,N_2036,N_2069);
xnor U2226 (N_2226,N_2162,N_2067);
nor U2227 (N_2227,N_2154,N_2100);
and U2228 (N_2228,N_2095,N_2196);
or U2229 (N_2229,N_2158,N_2090);
and U2230 (N_2230,N_2017,N_2138);
nor U2231 (N_2231,N_2178,N_2193);
nor U2232 (N_2232,N_2010,N_2002);
and U2233 (N_2233,N_2009,N_2092);
nand U2234 (N_2234,N_2012,N_2151);
nor U2235 (N_2235,N_2022,N_2091);
nor U2236 (N_2236,N_2019,N_2115);
or U2237 (N_2237,N_2132,N_2028);
nor U2238 (N_2238,N_2175,N_2182);
and U2239 (N_2239,N_2041,N_2149);
nand U2240 (N_2240,N_2065,N_2124);
nor U2241 (N_2241,N_2172,N_2056);
or U2242 (N_2242,N_2030,N_2089);
xor U2243 (N_2243,N_2070,N_2083);
or U2244 (N_2244,N_2157,N_2006);
nor U2245 (N_2245,N_2133,N_2185);
nand U2246 (N_2246,N_2137,N_2040);
or U2247 (N_2247,N_2187,N_2093);
nand U2248 (N_2248,N_2163,N_2101);
nand U2249 (N_2249,N_2079,N_2118);
and U2250 (N_2250,N_2146,N_2007);
or U2251 (N_2251,N_2081,N_2103);
and U2252 (N_2252,N_2020,N_2139);
and U2253 (N_2253,N_2098,N_2176);
nand U2254 (N_2254,N_2064,N_2167);
or U2255 (N_2255,N_2161,N_2084);
nand U2256 (N_2256,N_2164,N_2086);
and U2257 (N_2257,N_2108,N_2129);
xor U2258 (N_2258,N_2077,N_2085);
nand U2259 (N_2259,N_2024,N_2194);
and U2260 (N_2260,N_2057,N_2120);
nand U2261 (N_2261,N_2177,N_2076);
and U2262 (N_2262,N_2004,N_2147);
or U2263 (N_2263,N_2114,N_2192);
nor U2264 (N_2264,N_2155,N_2080);
nor U2265 (N_2265,N_2156,N_2038);
or U2266 (N_2266,N_2032,N_2188);
and U2267 (N_2267,N_2142,N_2061);
nor U2268 (N_2268,N_2014,N_2088);
nand U2269 (N_2269,N_2049,N_2173);
nand U2270 (N_2270,N_2066,N_2097);
nand U2271 (N_2271,N_2063,N_2122);
xor U2272 (N_2272,N_2099,N_2023);
nand U2273 (N_2273,N_2109,N_2071);
nor U2274 (N_2274,N_2021,N_2170);
or U2275 (N_2275,N_2034,N_2148);
and U2276 (N_2276,N_2073,N_2145);
nand U2277 (N_2277,N_2186,N_2130);
and U2278 (N_2278,N_2053,N_2105);
and U2279 (N_2279,N_2078,N_2143);
or U2280 (N_2280,N_2153,N_2037);
or U2281 (N_2281,N_2136,N_2111);
or U2282 (N_2282,N_2060,N_2102);
nor U2283 (N_2283,N_2144,N_2123);
nand U2284 (N_2284,N_2011,N_2166);
and U2285 (N_2285,N_2001,N_2112);
or U2286 (N_2286,N_2141,N_2016);
nand U2287 (N_2287,N_2183,N_2199);
or U2288 (N_2288,N_2043,N_2045);
nor U2289 (N_2289,N_2082,N_2189);
nand U2290 (N_2290,N_2029,N_2121);
and U2291 (N_2291,N_2039,N_2126);
and U2292 (N_2292,N_2131,N_2195);
nand U2293 (N_2293,N_2051,N_2106);
and U2294 (N_2294,N_2096,N_2181);
or U2295 (N_2295,N_2159,N_2062);
nand U2296 (N_2296,N_2055,N_2074);
and U2297 (N_2297,N_2047,N_2025);
nor U2298 (N_2298,N_2015,N_2197);
nand U2299 (N_2299,N_2119,N_2013);
or U2300 (N_2300,N_2185,N_2159);
nor U2301 (N_2301,N_2165,N_2152);
and U2302 (N_2302,N_2131,N_2160);
or U2303 (N_2303,N_2091,N_2043);
and U2304 (N_2304,N_2030,N_2065);
and U2305 (N_2305,N_2150,N_2189);
nand U2306 (N_2306,N_2047,N_2066);
and U2307 (N_2307,N_2101,N_2064);
and U2308 (N_2308,N_2115,N_2053);
nor U2309 (N_2309,N_2065,N_2103);
and U2310 (N_2310,N_2000,N_2052);
or U2311 (N_2311,N_2036,N_2025);
and U2312 (N_2312,N_2049,N_2102);
nor U2313 (N_2313,N_2076,N_2121);
and U2314 (N_2314,N_2070,N_2119);
nor U2315 (N_2315,N_2032,N_2130);
or U2316 (N_2316,N_2081,N_2137);
nor U2317 (N_2317,N_2190,N_2192);
or U2318 (N_2318,N_2127,N_2013);
and U2319 (N_2319,N_2036,N_2191);
nor U2320 (N_2320,N_2021,N_2154);
nand U2321 (N_2321,N_2047,N_2166);
nand U2322 (N_2322,N_2158,N_2037);
nor U2323 (N_2323,N_2075,N_2053);
nand U2324 (N_2324,N_2177,N_2199);
nor U2325 (N_2325,N_2126,N_2178);
and U2326 (N_2326,N_2192,N_2184);
or U2327 (N_2327,N_2037,N_2000);
and U2328 (N_2328,N_2136,N_2188);
or U2329 (N_2329,N_2151,N_2022);
nand U2330 (N_2330,N_2014,N_2148);
nor U2331 (N_2331,N_2171,N_2074);
and U2332 (N_2332,N_2188,N_2054);
nand U2333 (N_2333,N_2176,N_2189);
nor U2334 (N_2334,N_2190,N_2174);
and U2335 (N_2335,N_2159,N_2059);
nand U2336 (N_2336,N_2112,N_2031);
xor U2337 (N_2337,N_2170,N_2178);
nand U2338 (N_2338,N_2035,N_2148);
or U2339 (N_2339,N_2055,N_2096);
nor U2340 (N_2340,N_2006,N_2101);
nand U2341 (N_2341,N_2198,N_2164);
and U2342 (N_2342,N_2161,N_2067);
and U2343 (N_2343,N_2187,N_2034);
nor U2344 (N_2344,N_2060,N_2163);
or U2345 (N_2345,N_2079,N_2081);
or U2346 (N_2346,N_2177,N_2038);
and U2347 (N_2347,N_2081,N_2030);
nand U2348 (N_2348,N_2005,N_2018);
or U2349 (N_2349,N_2056,N_2072);
or U2350 (N_2350,N_2172,N_2111);
and U2351 (N_2351,N_2156,N_2185);
or U2352 (N_2352,N_2136,N_2032);
nor U2353 (N_2353,N_2144,N_2104);
and U2354 (N_2354,N_2041,N_2110);
or U2355 (N_2355,N_2034,N_2082);
and U2356 (N_2356,N_2074,N_2176);
nor U2357 (N_2357,N_2130,N_2143);
nor U2358 (N_2358,N_2175,N_2057);
xnor U2359 (N_2359,N_2153,N_2145);
nor U2360 (N_2360,N_2062,N_2060);
and U2361 (N_2361,N_2127,N_2086);
nand U2362 (N_2362,N_2062,N_2061);
or U2363 (N_2363,N_2118,N_2170);
nor U2364 (N_2364,N_2060,N_2138);
nor U2365 (N_2365,N_2011,N_2195);
and U2366 (N_2366,N_2183,N_2171);
nand U2367 (N_2367,N_2029,N_2067);
nor U2368 (N_2368,N_2178,N_2106);
and U2369 (N_2369,N_2168,N_2160);
and U2370 (N_2370,N_2147,N_2186);
and U2371 (N_2371,N_2003,N_2065);
or U2372 (N_2372,N_2119,N_2114);
and U2373 (N_2373,N_2085,N_2036);
nand U2374 (N_2374,N_2183,N_2012);
nor U2375 (N_2375,N_2103,N_2011);
nor U2376 (N_2376,N_2142,N_2062);
nand U2377 (N_2377,N_2008,N_2198);
and U2378 (N_2378,N_2164,N_2170);
or U2379 (N_2379,N_2079,N_2111);
xnor U2380 (N_2380,N_2100,N_2034);
nand U2381 (N_2381,N_2020,N_2163);
nand U2382 (N_2382,N_2063,N_2199);
nor U2383 (N_2383,N_2188,N_2038);
and U2384 (N_2384,N_2008,N_2071);
and U2385 (N_2385,N_2096,N_2145);
and U2386 (N_2386,N_2045,N_2134);
and U2387 (N_2387,N_2012,N_2056);
nand U2388 (N_2388,N_2008,N_2021);
nor U2389 (N_2389,N_2016,N_2113);
nand U2390 (N_2390,N_2155,N_2183);
nand U2391 (N_2391,N_2058,N_2147);
nand U2392 (N_2392,N_2017,N_2196);
or U2393 (N_2393,N_2148,N_2115);
nand U2394 (N_2394,N_2007,N_2192);
and U2395 (N_2395,N_2185,N_2054);
and U2396 (N_2396,N_2113,N_2098);
or U2397 (N_2397,N_2158,N_2131);
nand U2398 (N_2398,N_2172,N_2101);
nand U2399 (N_2399,N_2007,N_2015);
or U2400 (N_2400,N_2206,N_2259);
nand U2401 (N_2401,N_2333,N_2260);
or U2402 (N_2402,N_2345,N_2284);
nor U2403 (N_2403,N_2384,N_2386);
nor U2404 (N_2404,N_2231,N_2373);
nand U2405 (N_2405,N_2318,N_2283);
or U2406 (N_2406,N_2200,N_2289);
nand U2407 (N_2407,N_2346,N_2272);
and U2408 (N_2408,N_2217,N_2304);
xnor U2409 (N_2409,N_2311,N_2293);
or U2410 (N_2410,N_2308,N_2353);
nor U2411 (N_2411,N_2341,N_2327);
nand U2412 (N_2412,N_2285,N_2392);
nand U2413 (N_2413,N_2256,N_2339);
nand U2414 (N_2414,N_2383,N_2253);
xor U2415 (N_2415,N_2312,N_2249);
or U2416 (N_2416,N_2296,N_2230);
and U2417 (N_2417,N_2270,N_2251);
or U2418 (N_2418,N_2224,N_2320);
and U2419 (N_2419,N_2239,N_2374);
or U2420 (N_2420,N_2324,N_2314);
or U2421 (N_2421,N_2279,N_2243);
nand U2422 (N_2422,N_2273,N_2381);
and U2423 (N_2423,N_2370,N_2330);
nor U2424 (N_2424,N_2378,N_2263);
or U2425 (N_2425,N_2335,N_2238);
or U2426 (N_2426,N_2218,N_2380);
nand U2427 (N_2427,N_2264,N_2375);
and U2428 (N_2428,N_2344,N_2219);
and U2429 (N_2429,N_2385,N_2241);
and U2430 (N_2430,N_2315,N_2306);
nor U2431 (N_2431,N_2332,N_2365);
or U2432 (N_2432,N_2229,N_2313);
nand U2433 (N_2433,N_2292,N_2240);
nor U2434 (N_2434,N_2236,N_2280);
or U2435 (N_2435,N_2287,N_2212);
or U2436 (N_2436,N_2286,N_2294);
and U2437 (N_2437,N_2393,N_2355);
nand U2438 (N_2438,N_2337,N_2237);
nor U2439 (N_2439,N_2310,N_2371);
and U2440 (N_2440,N_2201,N_2362);
nand U2441 (N_2441,N_2208,N_2268);
or U2442 (N_2442,N_2363,N_2359);
or U2443 (N_2443,N_2319,N_2343);
nor U2444 (N_2444,N_2220,N_2336);
xnor U2445 (N_2445,N_2399,N_2334);
or U2446 (N_2446,N_2338,N_2356);
nor U2447 (N_2447,N_2303,N_2203);
or U2448 (N_2448,N_2248,N_2369);
nor U2449 (N_2449,N_2396,N_2367);
nor U2450 (N_2450,N_2269,N_2357);
nor U2451 (N_2451,N_2209,N_2326);
nand U2452 (N_2452,N_2349,N_2271);
and U2453 (N_2453,N_2202,N_2305);
nand U2454 (N_2454,N_2290,N_2258);
nor U2455 (N_2455,N_2226,N_2348);
or U2456 (N_2456,N_2277,N_2216);
and U2457 (N_2457,N_2382,N_2210);
and U2458 (N_2458,N_2321,N_2276);
and U2459 (N_2459,N_2261,N_2309);
and U2460 (N_2460,N_2300,N_2204);
and U2461 (N_2461,N_2390,N_2213);
or U2462 (N_2462,N_2351,N_2211);
and U2463 (N_2463,N_2347,N_2398);
nor U2464 (N_2464,N_2257,N_2372);
and U2465 (N_2465,N_2267,N_2215);
nand U2466 (N_2466,N_2235,N_2297);
nor U2467 (N_2467,N_2228,N_2282);
nor U2468 (N_2468,N_2262,N_2266);
or U2469 (N_2469,N_2274,N_2288);
nand U2470 (N_2470,N_2205,N_2227);
xor U2471 (N_2471,N_2299,N_2342);
nor U2472 (N_2472,N_2395,N_2387);
and U2473 (N_2473,N_2222,N_2354);
nand U2474 (N_2474,N_2225,N_2207);
or U2475 (N_2475,N_2397,N_2246);
and U2476 (N_2476,N_2265,N_2302);
nand U2477 (N_2477,N_2223,N_2301);
nor U2478 (N_2478,N_2323,N_2278);
nand U2479 (N_2479,N_2316,N_2352);
nand U2480 (N_2480,N_2242,N_2340);
nor U2481 (N_2481,N_2214,N_2329);
nand U2482 (N_2482,N_2275,N_2368);
nor U2483 (N_2483,N_2325,N_2358);
xor U2484 (N_2484,N_2254,N_2244);
nand U2485 (N_2485,N_2291,N_2233);
or U2486 (N_2486,N_2247,N_2350);
or U2487 (N_2487,N_2317,N_2328);
and U2488 (N_2488,N_2307,N_2388);
and U2489 (N_2489,N_2281,N_2252);
xnor U2490 (N_2490,N_2361,N_2391);
or U2491 (N_2491,N_2379,N_2376);
nor U2492 (N_2492,N_2255,N_2221);
nand U2493 (N_2493,N_2364,N_2234);
nor U2494 (N_2494,N_2389,N_2366);
and U2495 (N_2495,N_2377,N_2232);
nand U2496 (N_2496,N_2295,N_2322);
and U2497 (N_2497,N_2360,N_2298);
nand U2498 (N_2498,N_2331,N_2394);
nor U2499 (N_2499,N_2245,N_2250);
and U2500 (N_2500,N_2296,N_2244);
or U2501 (N_2501,N_2389,N_2202);
and U2502 (N_2502,N_2340,N_2223);
xnor U2503 (N_2503,N_2257,N_2374);
or U2504 (N_2504,N_2360,N_2286);
or U2505 (N_2505,N_2227,N_2330);
or U2506 (N_2506,N_2314,N_2203);
nor U2507 (N_2507,N_2369,N_2222);
nor U2508 (N_2508,N_2201,N_2393);
or U2509 (N_2509,N_2326,N_2330);
nor U2510 (N_2510,N_2275,N_2388);
nor U2511 (N_2511,N_2205,N_2224);
nor U2512 (N_2512,N_2315,N_2288);
nand U2513 (N_2513,N_2324,N_2243);
or U2514 (N_2514,N_2204,N_2347);
or U2515 (N_2515,N_2243,N_2254);
xor U2516 (N_2516,N_2376,N_2383);
or U2517 (N_2517,N_2245,N_2361);
nand U2518 (N_2518,N_2372,N_2250);
or U2519 (N_2519,N_2216,N_2242);
and U2520 (N_2520,N_2275,N_2361);
nand U2521 (N_2521,N_2354,N_2313);
nand U2522 (N_2522,N_2306,N_2374);
nand U2523 (N_2523,N_2248,N_2233);
nand U2524 (N_2524,N_2267,N_2293);
nand U2525 (N_2525,N_2328,N_2331);
nor U2526 (N_2526,N_2285,N_2347);
nand U2527 (N_2527,N_2289,N_2318);
and U2528 (N_2528,N_2212,N_2350);
or U2529 (N_2529,N_2284,N_2336);
or U2530 (N_2530,N_2203,N_2246);
nor U2531 (N_2531,N_2209,N_2217);
nor U2532 (N_2532,N_2238,N_2266);
and U2533 (N_2533,N_2324,N_2248);
nand U2534 (N_2534,N_2269,N_2336);
and U2535 (N_2535,N_2330,N_2347);
and U2536 (N_2536,N_2225,N_2285);
nand U2537 (N_2537,N_2227,N_2392);
nor U2538 (N_2538,N_2298,N_2204);
nand U2539 (N_2539,N_2338,N_2379);
nand U2540 (N_2540,N_2399,N_2273);
and U2541 (N_2541,N_2227,N_2266);
or U2542 (N_2542,N_2269,N_2395);
nand U2543 (N_2543,N_2251,N_2266);
or U2544 (N_2544,N_2339,N_2292);
nor U2545 (N_2545,N_2358,N_2252);
nor U2546 (N_2546,N_2290,N_2341);
nor U2547 (N_2547,N_2266,N_2333);
and U2548 (N_2548,N_2302,N_2262);
and U2549 (N_2549,N_2374,N_2217);
nor U2550 (N_2550,N_2228,N_2218);
nor U2551 (N_2551,N_2331,N_2377);
or U2552 (N_2552,N_2364,N_2252);
or U2553 (N_2553,N_2212,N_2357);
or U2554 (N_2554,N_2250,N_2211);
nor U2555 (N_2555,N_2298,N_2296);
or U2556 (N_2556,N_2253,N_2334);
nor U2557 (N_2557,N_2233,N_2344);
and U2558 (N_2558,N_2386,N_2355);
or U2559 (N_2559,N_2370,N_2293);
and U2560 (N_2560,N_2318,N_2312);
and U2561 (N_2561,N_2290,N_2235);
or U2562 (N_2562,N_2345,N_2367);
and U2563 (N_2563,N_2379,N_2385);
nand U2564 (N_2564,N_2219,N_2209);
and U2565 (N_2565,N_2215,N_2394);
nor U2566 (N_2566,N_2348,N_2394);
or U2567 (N_2567,N_2292,N_2259);
nor U2568 (N_2568,N_2373,N_2321);
nor U2569 (N_2569,N_2268,N_2384);
and U2570 (N_2570,N_2227,N_2236);
nand U2571 (N_2571,N_2394,N_2351);
and U2572 (N_2572,N_2268,N_2383);
and U2573 (N_2573,N_2278,N_2336);
or U2574 (N_2574,N_2383,N_2365);
nand U2575 (N_2575,N_2250,N_2397);
nand U2576 (N_2576,N_2211,N_2393);
and U2577 (N_2577,N_2221,N_2216);
nor U2578 (N_2578,N_2210,N_2272);
and U2579 (N_2579,N_2377,N_2262);
nand U2580 (N_2580,N_2320,N_2352);
or U2581 (N_2581,N_2216,N_2265);
nand U2582 (N_2582,N_2353,N_2315);
nor U2583 (N_2583,N_2393,N_2311);
nor U2584 (N_2584,N_2392,N_2359);
or U2585 (N_2585,N_2270,N_2291);
and U2586 (N_2586,N_2243,N_2344);
nand U2587 (N_2587,N_2345,N_2226);
nor U2588 (N_2588,N_2226,N_2364);
or U2589 (N_2589,N_2287,N_2293);
and U2590 (N_2590,N_2343,N_2270);
and U2591 (N_2591,N_2321,N_2213);
or U2592 (N_2592,N_2292,N_2229);
or U2593 (N_2593,N_2225,N_2239);
or U2594 (N_2594,N_2375,N_2328);
nand U2595 (N_2595,N_2382,N_2350);
nand U2596 (N_2596,N_2357,N_2221);
and U2597 (N_2597,N_2355,N_2374);
nand U2598 (N_2598,N_2371,N_2386);
and U2599 (N_2599,N_2378,N_2228);
or U2600 (N_2600,N_2519,N_2430);
nor U2601 (N_2601,N_2481,N_2467);
nor U2602 (N_2602,N_2419,N_2508);
or U2603 (N_2603,N_2468,N_2535);
or U2604 (N_2604,N_2490,N_2546);
and U2605 (N_2605,N_2543,N_2536);
nor U2606 (N_2606,N_2584,N_2484);
or U2607 (N_2607,N_2588,N_2573);
nand U2608 (N_2608,N_2445,N_2453);
or U2609 (N_2609,N_2450,N_2500);
or U2610 (N_2610,N_2458,N_2593);
nand U2611 (N_2611,N_2568,N_2581);
nor U2612 (N_2612,N_2447,N_2437);
nor U2613 (N_2613,N_2489,N_2492);
and U2614 (N_2614,N_2542,N_2544);
nor U2615 (N_2615,N_2572,N_2531);
or U2616 (N_2616,N_2442,N_2582);
and U2617 (N_2617,N_2518,N_2425);
nor U2618 (N_2618,N_2553,N_2406);
nor U2619 (N_2619,N_2441,N_2505);
or U2620 (N_2620,N_2548,N_2448);
nand U2621 (N_2621,N_2552,N_2459);
nand U2622 (N_2622,N_2583,N_2504);
and U2623 (N_2623,N_2452,N_2549);
nor U2624 (N_2624,N_2525,N_2407);
nand U2625 (N_2625,N_2440,N_2408);
nor U2626 (N_2626,N_2513,N_2520);
and U2627 (N_2627,N_2416,N_2592);
nand U2628 (N_2628,N_2483,N_2558);
nor U2629 (N_2629,N_2559,N_2578);
nor U2630 (N_2630,N_2574,N_2455);
nand U2631 (N_2631,N_2598,N_2511);
nor U2632 (N_2632,N_2554,N_2521);
and U2633 (N_2633,N_2556,N_2576);
or U2634 (N_2634,N_2527,N_2497);
and U2635 (N_2635,N_2404,N_2538);
nand U2636 (N_2636,N_2461,N_2493);
and U2637 (N_2637,N_2462,N_2495);
or U2638 (N_2638,N_2514,N_2571);
nand U2639 (N_2639,N_2491,N_2402);
nand U2640 (N_2640,N_2526,N_2503);
or U2641 (N_2641,N_2512,N_2522);
nor U2642 (N_2642,N_2565,N_2411);
nor U2643 (N_2643,N_2537,N_2560);
or U2644 (N_2644,N_2569,N_2469);
nor U2645 (N_2645,N_2443,N_2541);
nor U2646 (N_2646,N_2475,N_2501);
xor U2647 (N_2647,N_2436,N_2479);
nand U2648 (N_2648,N_2524,N_2426);
or U2649 (N_2649,N_2597,N_2456);
nor U2650 (N_2650,N_2446,N_2562);
or U2651 (N_2651,N_2439,N_2463);
or U2652 (N_2652,N_2557,N_2400);
or U2653 (N_2653,N_2488,N_2540);
nand U2654 (N_2654,N_2473,N_2551);
nor U2655 (N_2655,N_2561,N_2580);
nand U2656 (N_2656,N_2486,N_2494);
and U2657 (N_2657,N_2516,N_2499);
nor U2658 (N_2658,N_2424,N_2529);
nor U2659 (N_2659,N_2451,N_2471);
or U2660 (N_2660,N_2547,N_2575);
nand U2661 (N_2661,N_2431,N_2550);
and U2662 (N_2662,N_2566,N_2434);
nand U2663 (N_2663,N_2496,N_2465);
nand U2664 (N_2664,N_2466,N_2413);
or U2665 (N_2665,N_2405,N_2534);
and U2666 (N_2666,N_2594,N_2401);
and U2667 (N_2667,N_2433,N_2596);
or U2668 (N_2668,N_2482,N_2435);
or U2669 (N_2669,N_2589,N_2570);
nand U2670 (N_2670,N_2586,N_2506);
nand U2671 (N_2671,N_2507,N_2528);
and U2672 (N_2672,N_2474,N_2478);
nor U2673 (N_2673,N_2533,N_2595);
nand U2674 (N_2674,N_2599,N_2444);
or U2675 (N_2675,N_2422,N_2421);
and U2676 (N_2676,N_2539,N_2567);
or U2677 (N_2677,N_2485,N_2454);
or U2678 (N_2678,N_2410,N_2487);
or U2679 (N_2679,N_2480,N_2412);
nor U2680 (N_2680,N_2470,N_2428);
and U2681 (N_2681,N_2517,N_2498);
nor U2682 (N_2682,N_2432,N_2476);
nand U2683 (N_2683,N_2457,N_2510);
nand U2684 (N_2684,N_2420,N_2429);
nor U2685 (N_2685,N_2403,N_2417);
nand U2686 (N_2686,N_2591,N_2423);
nor U2687 (N_2687,N_2438,N_2460);
nor U2688 (N_2688,N_2564,N_2502);
and U2689 (N_2689,N_2515,N_2590);
nor U2690 (N_2690,N_2472,N_2587);
or U2691 (N_2691,N_2449,N_2545);
nor U2692 (N_2692,N_2577,N_2555);
and U2693 (N_2693,N_2530,N_2427);
nor U2694 (N_2694,N_2585,N_2418);
or U2695 (N_2695,N_2579,N_2477);
nand U2696 (N_2696,N_2563,N_2509);
and U2697 (N_2697,N_2532,N_2415);
or U2698 (N_2698,N_2523,N_2464);
nand U2699 (N_2699,N_2414,N_2409);
nor U2700 (N_2700,N_2593,N_2545);
nor U2701 (N_2701,N_2465,N_2493);
and U2702 (N_2702,N_2596,N_2571);
and U2703 (N_2703,N_2496,N_2554);
xnor U2704 (N_2704,N_2439,N_2503);
and U2705 (N_2705,N_2405,N_2570);
nand U2706 (N_2706,N_2523,N_2412);
nor U2707 (N_2707,N_2516,N_2522);
and U2708 (N_2708,N_2474,N_2429);
nand U2709 (N_2709,N_2549,N_2513);
and U2710 (N_2710,N_2418,N_2443);
or U2711 (N_2711,N_2429,N_2406);
and U2712 (N_2712,N_2475,N_2436);
and U2713 (N_2713,N_2557,N_2467);
xnor U2714 (N_2714,N_2562,N_2421);
or U2715 (N_2715,N_2466,N_2492);
or U2716 (N_2716,N_2505,N_2595);
nor U2717 (N_2717,N_2510,N_2587);
or U2718 (N_2718,N_2540,N_2479);
and U2719 (N_2719,N_2454,N_2544);
nand U2720 (N_2720,N_2596,N_2512);
xor U2721 (N_2721,N_2409,N_2408);
and U2722 (N_2722,N_2517,N_2582);
nand U2723 (N_2723,N_2401,N_2544);
or U2724 (N_2724,N_2474,N_2444);
and U2725 (N_2725,N_2456,N_2516);
nand U2726 (N_2726,N_2468,N_2494);
and U2727 (N_2727,N_2503,N_2447);
and U2728 (N_2728,N_2423,N_2421);
and U2729 (N_2729,N_2512,N_2537);
and U2730 (N_2730,N_2477,N_2565);
nor U2731 (N_2731,N_2419,N_2480);
and U2732 (N_2732,N_2469,N_2578);
nor U2733 (N_2733,N_2419,N_2471);
or U2734 (N_2734,N_2472,N_2425);
nand U2735 (N_2735,N_2412,N_2513);
nand U2736 (N_2736,N_2557,N_2532);
or U2737 (N_2737,N_2551,N_2445);
nand U2738 (N_2738,N_2419,N_2429);
or U2739 (N_2739,N_2577,N_2469);
nor U2740 (N_2740,N_2579,N_2478);
nor U2741 (N_2741,N_2502,N_2542);
and U2742 (N_2742,N_2575,N_2425);
nand U2743 (N_2743,N_2464,N_2402);
nor U2744 (N_2744,N_2550,N_2508);
xnor U2745 (N_2745,N_2533,N_2492);
xnor U2746 (N_2746,N_2467,N_2544);
nand U2747 (N_2747,N_2458,N_2588);
nand U2748 (N_2748,N_2433,N_2517);
nand U2749 (N_2749,N_2582,N_2403);
nand U2750 (N_2750,N_2502,N_2416);
and U2751 (N_2751,N_2594,N_2490);
or U2752 (N_2752,N_2520,N_2581);
or U2753 (N_2753,N_2482,N_2461);
nor U2754 (N_2754,N_2489,N_2495);
nand U2755 (N_2755,N_2437,N_2467);
or U2756 (N_2756,N_2461,N_2442);
or U2757 (N_2757,N_2433,N_2406);
nor U2758 (N_2758,N_2592,N_2490);
and U2759 (N_2759,N_2495,N_2491);
nor U2760 (N_2760,N_2410,N_2574);
nor U2761 (N_2761,N_2575,N_2500);
xnor U2762 (N_2762,N_2534,N_2469);
nand U2763 (N_2763,N_2526,N_2554);
nor U2764 (N_2764,N_2433,N_2475);
and U2765 (N_2765,N_2424,N_2457);
nor U2766 (N_2766,N_2458,N_2414);
and U2767 (N_2767,N_2470,N_2542);
nand U2768 (N_2768,N_2506,N_2530);
nand U2769 (N_2769,N_2463,N_2517);
nor U2770 (N_2770,N_2567,N_2585);
and U2771 (N_2771,N_2518,N_2460);
and U2772 (N_2772,N_2425,N_2565);
nor U2773 (N_2773,N_2583,N_2467);
or U2774 (N_2774,N_2555,N_2554);
nor U2775 (N_2775,N_2528,N_2586);
nand U2776 (N_2776,N_2527,N_2433);
nand U2777 (N_2777,N_2579,N_2556);
nand U2778 (N_2778,N_2419,N_2555);
nand U2779 (N_2779,N_2438,N_2476);
nand U2780 (N_2780,N_2549,N_2472);
nor U2781 (N_2781,N_2412,N_2409);
or U2782 (N_2782,N_2540,N_2589);
nand U2783 (N_2783,N_2429,N_2518);
or U2784 (N_2784,N_2457,N_2522);
nor U2785 (N_2785,N_2501,N_2582);
and U2786 (N_2786,N_2584,N_2478);
or U2787 (N_2787,N_2564,N_2428);
and U2788 (N_2788,N_2404,N_2483);
nor U2789 (N_2789,N_2407,N_2475);
nor U2790 (N_2790,N_2598,N_2414);
nor U2791 (N_2791,N_2423,N_2496);
or U2792 (N_2792,N_2480,N_2478);
or U2793 (N_2793,N_2480,N_2587);
nand U2794 (N_2794,N_2400,N_2513);
nand U2795 (N_2795,N_2504,N_2557);
or U2796 (N_2796,N_2518,N_2411);
xnor U2797 (N_2797,N_2597,N_2409);
nor U2798 (N_2798,N_2513,N_2477);
and U2799 (N_2799,N_2514,N_2559);
and U2800 (N_2800,N_2642,N_2781);
nor U2801 (N_2801,N_2796,N_2668);
xnor U2802 (N_2802,N_2712,N_2605);
and U2803 (N_2803,N_2609,N_2624);
nand U2804 (N_2804,N_2688,N_2734);
nor U2805 (N_2805,N_2627,N_2662);
nor U2806 (N_2806,N_2720,N_2697);
or U2807 (N_2807,N_2726,N_2762);
or U2808 (N_2808,N_2665,N_2764);
or U2809 (N_2809,N_2717,N_2696);
nor U2810 (N_2810,N_2746,N_2659);
xnor U2811 (N_2811,N_2719,N_2692);
nand U2812 (N_2812,N_2767,N_2608);
nand U2813 (N_2813,N_2647,N_2669);
and U2814 (N_2814,N_2655,N_2775);
nand U2815 (N_2815,N_2693,N_2721);
or U2816 (N_2816,N_2760,N_2643);
nor U2817 (N_2817,N_2610,N_2792);
nor U2818 (N_2818,N_2616,N_2711);
nand U2819 (N_2819,N_2735,N_2741);
nand U2820 (N_2820,N_2667,N_2615);
and U2821 (N_2821,N_2634,N_2748);
and U2822 (N_2822,N_2695,N_2701);
nor U2823 (N_2823,N_2736,N_2744);
nor U2824 (N_2824,N_2705,N_2670);
nor U2825 (N_2825,N_2638,N_2739);
nand U2826 (N_2826,N_2745,N_2779);
and U2827 (N_2827,N_2679,N_2621);
nand U2828 (N_2828,N_2788,N_2786);
and U2829 (N_2829,N_2718,N_2689);
and U2830 (N_2830,N_2780,N_2639);
nand U2831 (N_2831,N_2755,N_2797);
nand U2832 (N_2832,N_2682,N_2602);
nand U2833 (N_2833,N_2672,N_2600);
or U2834 (N_2834,N_2683,N_2607);
or U2835 (N_2835,N_2675,N_2790);
and U2836 (N_2836,N_2687,N_2770);
or U2837 (N_2837,N_2614,N_2731);
or U2838 (N_2838,N_2623,N_2759);
and U2839 (N_2839,N_2691,N_2740);
and U2840 (N_2840,N_2631,N_2771);
nand U2841 (N_2841,N_2628,N_2650);
or U2842 (N_2842,N_2793,N_2657);
nor U2843 (N_2843,N_2632,N_2603);
and U2844 (N_2844,N_2730,N_2722);
xor U2845 (N_2845,N_2795,N_2799);
nand U2846 (N_2846,N_2749,N_2651);
or U2847 (N_2847,N_2728,N_2769);
or U2848 (N_2848,N_2787,N_2622);
nand U2849 (N_2849,N_2676,N_2648);
or U2850 (N_2850,N_2686,N_2646);
or U2851 (N_2851,N_2751,N_2625);
and U2852 (N_2852,N_2747,N_2737);
nor U2853 (N_2853,N_2654,N_2753);
nand U2854 (N_2854,N_2777,N_2708);
or U2855 (N_2855,N_2791,N_2611);
nor U2856 (N_2856,N_2633,N_2703);
nor U2857 (N_2857,N_2698,N_2773);
nor U2858 (N_2858,N_2617,N_2680);
nand U2859 (N_2859,N_2757,N_2626);
or U2860 (N_2860,N_2715,N_2727);
or U2861 (N_2861,N_2723,N_2699);
nand U2862 (N_2862,N_2778,N_2644);
nand U2863 (N_2863,N_2794,N_2684);
and U2864 (N_2864,N_2690,N_2613);
nor U2865 (N_2865,N_2635,N_2782);
and U2866 (N_2866,N_2758,N_2776);
nand U2867 (N_2867,N_2750,N_2700);
nor U2868 (N_2868,N_2707,N_2704);
or U2869 (N_2869,N_2702,N_2754);
nor U2870 (N_2870,N_2619,N_2729);
nand U2871 (N_2871,N_2636,N_2725);
and U2872 (N_2872,N_2706,N_2783);
and U2873 (N_2873,N_2716,N_2685);
nand U2874 (N_2874,N_2653,N_2601);
or U2875 (N_2875,N_2694,N_2671);
nand U2876 (N_2876,N_2630,N_2606);
nor U2877 (N_2877,N_2738,N_2714);
and U2878 (N_2878,N_2743,N_2629);
and U2879 (N_2879,N_2677,N_2798);
and U2880 (N_2880,N_2742,N_2656);
xnor U2881 (N_2881,N_2620,N_2724);
and U2882 (N_2882,N_2774,N_2763);
and U2883 (N_2883,N_2666,N_2612);
nor U2884 (N_2884,N_2664,N_2637);
or U2885 (N_2885,N_2649,N_2673);
and U2886 (N_2886,N_2645,N_2785);
nand U2887 (N_2887,N_2663,N_2765);
nand U2888 (N_2888,N_2784,N_2752);
nand U2889 (N_2889,N_2618,N_2660);
or U2890 (N_2890,N_2640,N_2709);
nor U2891 (N_2891,N_2674,N_2678);
or U2892 (N_2892,N_2768,N_2658);
or U2893 (N_2893,N_2661,N_2710);
and U2894 (N_2894,N_2652,N_2772);
nand U2895 (N_2895,N_2766,N_2681);
and U2896 (N_2896,N_2733,N_2713);
and U2897 (N_2897,N_2641,N_2761);
or U2898 (N_2898,N_2732,N_2789);
nor U2899 (N_2899,N_2604,N_2756);
or U2900 (N_2900,N_2674,N_2781);
nor U2901 (N_2901,N_2682,N_2692);
nand U2902 (N_2902,N_2695,N_2668);
nand U2903 (N_2903,N_2614,N_2777);
nor U2904 (N_2904,N_2751,N_2785);
nand U2905 (N_2905,N_2689,N_2741);
and U2906 (N_2906,N_2738,N_2793);
or U2907 (N_2907,N_2631,N_2708);
or U2908 (N_2908,N_2732,N_2700);
and U2909 (N_2909,N_2647,N_2730);
nor U2910 (N_2910,N_2651,N_2774);
and U2911 (N_2911,N_2796,N_2643);
xor U2912 (N_2912,N_2668,N_2627);
nor U2913 (N_2913,N_2673,N_2763);
nand U2914 (N_2914,N_2676,N_2737);
or U2915 (N_2915,N_2648,N_2691);
or U2916 (N_2916,N_2769,N_2754);
nand U2917 (N_2917,N_2600,N_2731);
or U2918 (N_2918,N_2619,N_2709);
nand U2919 (N_2919,N_2703,N_2718);
nand U2920 (N_2920,N_2713,N_2760);
or U2921 (N_2921,N_2640,N_2643);
nor U2922 (N_2922,N_2728,N_2708);
and U2923 (N_2923,N_2600,N_2742);
nand U2924 (N_2924,N_2694,N_2677);
nand U2925 (N_2925,N_2790,N_2633);
nor U2926 (N_2926,N_2747,N_2729);
and U2927 (N_2927,N_2784,N_2680);
or U2928 (N_2928,N_2709,N_2717);
and U2929 (N_2929,N_2792,N_2657);
and U2930 (N_2930,N_2681,N_2764);
nor U2931 (N_2931,N_2657,N_2781);
and U2932 (N_2932,N_2671,N_2747);
or U2933 (N_2933,N_2708,N_2797);
and U2934 (N_2934,N_2678,N_2685);
or U2935 (N_2935,N_2702,N_2796);
nor U2936 (N_2936,N_2668,N_2663);
or U2937 (N_2937,N_2778,N_2697);
nand U2938 (N_2938,N_2751,N_2793);
and U2939 (N_2939,N_2703,N_2762);
or U2940 (N_2940,N_2791,N_2683);
or U2941 (N_2941,N_2626,N_2717);
nor U2942 (N_2942,N_2671,N_2798);
nor U2943 (N_2943,N_2702,N_2704);
nor U2944 (N_2944,N_2735,N_2787);
and U2945 (N_2945,N_2644,N_2759);
nand U2946 (N_2946,N_2748,N_2668);
nand U2947 (N_2947,N_2742,N_2671);
and U2948 (N_2948,N_2797,N_2611);
and U2949 (N_2949,N_2764,N_2675);
and U2950 (N_2950,N_2616,N_2701);
or U2951 (N_2951,N_2726,N_2640);
nand U2952 (N_2952,N_2781,N_2662);
and U2953 (N_2953,N_2629,N_2707);
or U2954 (N_2954,N_2614,N_2630);
or U2955 (N_2955,N_2684,N_2781);
nor U2956 (N_2956,N_2661,N_2726);
and U2957 (N_2957,N_2666,N_2674);
and U2958 (N_2958,N_2695,N_2786);
nand U2959 (N_2959,N_2633,N_2662);
nor U2960 (N_2960,N_2633,N_2678);
and U2961 (N_2961,N_2679,N_2685);
or U2962 (N_2962,N_2765,N_2645);
nand U2963 (N_2963,N_2775,N_2656);
or U2964 (N_2964,N_2669,N_2606);
nor U2965 (N_2965,N_2617,N_2762);
nand U2966 (N_2966,N_2796,N_2762);
nand U2967 (N_2967,N_2750,N_2767);
nor U2968 (N_2968,N_2683,N_2728);
nor U2969 (N_2969,N_2736,N_2626);
nor U2970 (N_2970,N_2734,N_2719);
and U2971 (N_2971,N_2703,N_2604);
nand U2972 (N_2972,N_2680,N_2786);
and U2973 (N_2973,N_2768,N_2669);
nand U2974 (N_2974,N_2724,N_2767);
and U2975 (N_2975,N_2720,N_2609);
nand U2976 (N_2976,N_2644,N_2695);
nor U2977 (N_2977,N_2710,N_2677);
and U2978 (N_2978,N_2736,N_2749);
or U2979 (N_2979,N_2632,N_2711);
nand U2980 (N_2980,N_2785,N_2757);
nor U2981 (N_2981,N_2640,N_2790);
nor U2982 (N_2982,N_2618,N_2706);
or U2983 (N_2983,N_2636,N_2699);
or U2984 (N_2984,N_2686,N_2776);
nand U2985 (N_2985,N_2772,N_2754);
and U2986 (N_2986,N_2709,N_2753);
nor U2987 (N_2987,N_2665,N_2772);
nor U2988 (N_2988,N_2716,N_2632);
nor U2989 (N_2989,N_2653,N_2674);
and U2990 (N_2990,N_2657,N_2670);
or U2991 (N_2991,N_2645,N_2782);
and U2992 (N_2992,N_2779,N_2695);
or U2993 (N_2993,N_2775,N_2704);
nor U2994 (N_2994,N_2684,N_2770);
nor U2995 (N_2995,N_2740,N_2670);
or U2996 (N_2996,N_2667,N_2715);
and U2997 (N_2997,N_2797,N_2796);
and U2998 (N_2998,N_2620,N_2780);
or U2999 (N_2999,N_2743,N_2715);
nand UO_0 (O_0,N_2837,N_2917);
or UO_1 (O_1,N_2921,N_2892);
nand UO_2 (O_2,N_2934,N_2935);
or UO_3 (O_3,N_2931,N_2924);
and UO_4 (O_4,N_2802,N_2918);
nor UO_5 (O_5,N_2806,N_2888);
or UO_6 (O_6,N_2875,N_2862);
nand UO_7 (O_7,N_2803,N_2982);
nand UO_8 (O_8,N_2913,N_2833);
or UO_9 (O_9,N_2940,N_2811);
nand UO_10 (O_10,N_2828,N_2815);
and UO_11 (O_11,N_2844,N_2852);
or UO_12 (O_12,N_2867,N_2958);
nand UO_13 (O_13,N_2963,N_2971);
or UO_14 (O_14,N_2933,N_2952);
nand UO_15 (O_15,N_2826,N_2981);
or UO_16 (O_16,N_2987,N_2871);
nor UO_17 (O_17,N_2832,N_2807);
and UO_18 (O_18,N_2996,N_2907);
and UO_19 (O_19,N_2962,N_2980);
and UO_20 (O_20,N_2883,N_2973);
and UO_21 (O_21,N_2863,N_2894);
and UO_22 (O_22,N_2847,N_2884);
or UO_23 (O_23,N_2845,N_2860);
or UO_24 (O_24,N_2813,N_2912);
nand UO_25 (O_25,N_2881,N_2910);
and UO_26 (O_26,N_2843,N_2974);
nand UO_27 (O_27,N_2817,N_2842);
nand UO_28 (O_28,N_2870,N_2868);
and UO_29 (O_29,N_2998,N_2818);
or UO_30 (O_30,N_2930,N_2941);
and UO_31 (O_31,N_2967,N_2919);
or UO_32 (O_32,N_2887,N_2994);
or UO_33 (O_33,N_2923,N_2808);
nor UO_34 (O_34,N_2893,N_2915);
nand UO_35 (O_35,N_2976,N_2947);
nor UO_36 (O_36,N_2873,N_2819);
xnor UO_37 (O_37,N_2890,N_2951);
nor UO_38 (O_38,N_2966,N_2834);
or UO_39 (O_39,N_2926,N_2920);
nand UO_40 (O_40,N_2928,N_2820);
and UO_41 (O_41,N_2929,N_2932);
nand UO_42 (O_42,N_2911,N_2972);
nor UO_43 (O_43,N_2827,N_2897);
or UO_44 (O_44,N_2969,N_2825);
or UO_45 (O_45,N_2876,N_2960);
nand UO_46 (O_46,N_2851,N_2809);
nor UO_47 (O_47,N_2838,N_2992);
nand UO_48 (O_48,N_2841,N_2985);
and UO_49 (O_49,N_2950,N_2885);
nand UO_50 (O_50,N_2814,N_2872);
or UO_51 (O_51,N_2999,N_2936);
nand UO_52 (O_52,N_2943,N_2965);
nand UO_53 (O_53,N_2800,N_2908);
nor UO_54 (O_54,N_2961,N_2927);
nor UO_55 (O_55,N_2900,N_2849);
nor UO_56 (O_56,N_2954,N_2948);
nor UO_57 (O_57,N_2895,N_2836);
nor UO_58 (O_58,N_2901,N_2988);
or UO_59 (O_59,N_2970,N_2922);
nor UO_60 (O_60,N_2939,N_2821);
nand UO_61 (O_61,N_2977,N_2856);
or UO_62 (O_62,N_2964,N_2906);
or UO_63 (O_63,N_2801,N_2953);
nor UO_64 (O_64,N_2830,N_2916);
nor UO_65 (O_65,N_2882,N_2861);
xor UO_66 (O_66,N_2984,N_2831);
or UO_67 (O_67,N_2839,N_2903);
nand UO_68 (O_68,N_2978,N_2989);
nor UO_69 (O_69,N_2848,N_2983);
and UO_70 (O_70,N_2902,N_2829);
or UO_71 (O_71,N_2975,N_2986);
and UO_72 (O_72,N_2914,N_2835);
nand UO_73 (O_73,N_2938,N_2904);
nand UO_74 (O_74,N_2822,N_2846);
xnor UO_75 (O_75,N_2812,N_2959);
nor UO_76 (O_76,N_2855,N_2991);
nor UO_77 (O_77,N_2898,N_2993);
nor UO_78 (O_78,N_2816,N_2823);
nand UO_79 (O_79,N_2891,N_2854);
nand UO_80 (O_80,N_2879,N_2864);
nand UO_81 (O_81,N_2858,N_2886);
and UO_82 (O_82,N_2857,N_2909);
or UO_83 (O_83,N_2956,N_2942);
and UO_84 (O_84,N_2874,N_2804);
or UO_85 (O_85,N_2866,N_2949);
nor UO_86 (O_86,N_2896,N_2877);
and UO_87 (O_87,N_2995,N_2840);
nand UO_88 (O_88,N_2853,N_2869);
nor UO_89 (O_89,N_2944,N_2880);
or UO_90 (O_90,N_2824,N_2899);
and UO_91 (O_91,N_2946,N_2955);
and UO_92 (O_92,N_2878,N_2957);
nand UO_93 (O_93,N_2997,N_2937);
or UO_94 (O_94,N_2979,N_2945);
or UO_95 (O_95,N_2990,N_2810);
or UO_96 (O_96,N_2865,N_2905);
nor UO_97 (O_97,N_2925,N_2889);
or UO_98 (O_98,N_2859,N_2968);
and UO_99 (O_99,N_2805,N_2850);
or UO_100 (O_100,N_2867,N_2813);
or UO_101 (O_101,N_2976,N_2961);
and UO_102 (O_102,N_2858,N_2935);
or UO_103 (O_103,N_2860,N_2904);
nor UO_104 (O_104,N_2967,N_2978);
or UO_105 (O_105,N_2963,N_2807);
or UO_106 (O_106,N_2835,N_2805);
or UO_107 (O_107,N_2801,N_2885);
and UO_108 (O_108,N_2879,N_2810);
nand UO_109 (O_109,N_2803,N_2816);
nand UO_110 (O_110,N_2884,N_2859);
nand UO_111 (O_111,N_2814,N_2849);
nor UO_112 (O_112,N_2926,N_2916);
nor UO_113 (O_113,N_2966,N_2887);
or UO_114 (O_114,N_2966,N_2959);
nor UO_115 (O_115,N_2918,N_2922);
nor UO_116 (O_116,N_2988,N_2896);
nand UO_117 (O_117,N_2865,N_2923);
or UO_118 (O_118,N_2918,N_2841);
or UO_119 (O_119,N_2946,N_2884);
nand UO_120 (O_120,N_2870,N_2839);
nand UO_121 (O_121,N_2802,N_2819);
and UO_122 (O_122,N_2956,N_2982);
and UO_123 (O_123,N_2937,N_2855);
and UO_124 (O_124,N_2812,N_2832);
and UO_125 (O_125,N_2974,N_2925);
or UO_126 (O_126,N_2894,N_2887);
and UO_127 (O_127,N_2937,N_2947);
and UO_128 (O_128,N_2833,N_2981);
or UO_129 (O_129,N_2846,N_2841);
nor UO_130 (O_130,N_2903,N_2945);
nor UO_131 (O_131,N_2884,N_2977);
or UO_132 (O_132,N_2923,N_2912);
nor UO_133 (O_133,N_2971,N_2841);
nor UO_134 (O_134,N_2930,N_2831);
nand UO_135 (O_135,N_2874,N_2951);
and UO_136 (O_136,N_2930,N_2925);
and UO_137 (O_137,N_2839,N_2954);
or UO_138 (O_138,N_2874,N_2986);
nor UO_139 (O_139,N_2904,N_2834);
nor UO_140 (O_140,N_2835,N_2895);
and UO_141 (O_141,N_2985,N_2850);
or UO_142 (O_142,N_2863,N_2845);
nor UO_143 (O_143,N_2999,N_2981);
or UO_144 (O_144,N_2942,N_2915);
or UO_145 (O_145,N_2946,N_2853);
nor UO_146 (O_146,N_2942,N_2809);
and UO_147 (O_147,N_2993,N_2860);
or UO_148 (O_148,N_2913,N_2872);
and UO_149 (O_149,N_2862,N_2936);
or UO_150 (O_150,N_2962,N_2811);
nand UO_151 (O_151,N_2879,N_2933);
xnor UO_152 (O_152,N_2975,N_2997);
or UO_153 (O_153,N_2814,N_2808);
nor UO_154 (O_154,N_2833,N_2977);
nor UO_155 (O_155,N_2848,N_2803);
nand UO_156 (O_156,N_2981,N_2936);
and UO_157 (O_157,N_2980,N_2908);
and UO_158 (O_158,N_2860,N_2989);
and UO_159 (O_159,N_2896,N_2904);
and UO_160 (O_160,N_2986,N_2939);
nand UO_161 (O_161,N_2870,N_2983);
xor UO_162 (O_162,N_2868,N_2930);
and UO_163 (O_163,N_2962,N_2991);
nand UO_164 (O_164,N_2945,N_2918);
nor UO_165 (O_165,N_2848,N_2939);
or UO_166 (O_166,N_2931,N_2980);
nor UO_167 (O_167,N_2989,N_2853);
or UO_168 (O_168,N_2866,N_2881);
and UO_169 (O_169,N_2972,N_2905);
or UO_170 (O_170,N_2833,N_2890);
and UO_171 (O_171,N_2926,N_2964);
nor UO_172 (O_172,N_2904,N_2806);
nand UO_173 (O_173,N_2821,N_2827);
or UO_174 (O_174,N_2947,N_2936);
and UO_175 (O_175,N_2827,N_2815);
or UO_176 (O_176,N_2860,N_2926);
nor UO_177 (O_177,N_2811,N_2955);
nor UO_178 (O_178,N_2956,N_2874);
or UO_179 (O_179,N_2951,N_2835);
nor UO_180 (O_180,N_2986,N_2885);
or UO_181 (O_181,N_2980,N_2813);
or UO_182 (O_182,N_2941,N_2847);
xor UO_183 (O_183,N_2998,N_2962);
or UO_184 (O_184,N_2877,N_2942);
nand UO_185 (O_185,N_2803,N_2943);
and UO_186 (O_186,N_2972,N_2861);
and UO_187 (O_187,N_2842,N_2865);
xor UO_188 (O_188,N_2806,N_2970);
and UO_189 (O_189,N_2808,N_2813);
nor UO_190 (O_190,N_2847,N_2899);
nand UO_191 (O_191,N_2822,N_2944);
and UO_192 (O_192,N_2832,N_2872);
nand UO_193 (O_193,N_2808,N_2918);
and UO_194 (O_194,N_2962,N_2942);
nor UO_195 (O_195,N_2865,N_2965);
nand UO_196 (O_196,N_2841,N_2813);
and UO_197 (O_197,N_2926,N_2879);
and UO_198 (O_198,N_2887,N_2982);
nand UO_199 (O_199,N_2812,N_2826);
nor UO_200 (O_200,N_2812,N_2879);
nand UO_201 (O_201,N_2950,N_2900);
nand UO_202 (O_202,N_2896,N_2848);
and UO_203 (O_203,N_2932,N_2985);
or UO_204 (O_204,N_2998,N_2892);
nand UO_205 (O_205,N_2941,N_2873);
nand UO_206 (O_206,N_2880,N_2878);
and UO_207 (O_207,N_2848,N_2835);
nor UO_208 (O_208,N_2945,N_2957);
and UO_209 (O_209,N_2979,N_2838);
and UO_210 (O_210,N_2998,N_2873);
and UO_211 (O_211,N_2806,N_2871);
or UO_212 (O_212,N_2823,N_2930);
and UO_213 (O_213,N_2848,N_2915);
nor UO_214 (O_214,N_2825,N_2856);
and UO_215 (O_215,N_2948,N_2837);
nand UO_216 (O_216,N_2804,N_2810);
and UO_217 (O_217,N_2981,N_2870);
nor UO_218 (O_218,N_2834,N_2972);
nor UO_219 (O_219,N_2998,N_2943);
nand UO_220 (O_220,N_2845,N_2801);
and UO_221 (O_221,N_2808,N_2944);
nand UO_222 (O_222,N_2942,N_2997);
or UO_223 (O_223,N_2989,N_2918);
or UO_224 (O_224,N_2890,N_2801);
or UO_225 (O_225,N_2803,N_2915);
and UO_226 (O_226,N_2838,N_2822);
nor UO_227 (O_227,N_2926,N_2984);
nor UO_228 (O_228,N_2937,N_2945);
and UO_229 (O_229,N_2941,N_2883);
nand UO_230 (O_230,N_2976,N_2834);
and UO_231 (O_231,N_2922,N_2835);
nand UO_232 (O_232,N_2885,N_2844);
or UO_233 (O_233,N_2842,N_2931);
nand UO_234 (O_234,N_2826,N_2997);
and UO_235 (O_235,N_2804,N_2840);
and UO_236 (O_236,N_2822,N_2860);
nor UO_237 (O_237,N_2867,N_2851);
and UO_238 (O_238,N_2849,N_2847);
and UO_239 (O_239,N_2801,N_2852);
or UO_240 (O_240,N_2923,N_2881);
nor UO_241 (O_241,N_2867,N_2921);
and UO_242 (O_242,N_2949,N_2909);
nand UO_243 (O_243,N_2818,N_2856);
or UO_244 (O_244,N_2917,N_2987);
nor UO_245 (O_245,N_2930,N_2981);
or UO_246 (O_246,N_2881,N_2834);
nor UO_247 (O_247,N_2920,N_2977);
nor UO_248 (O_248,N_2894,N_2908);
and UO_249 (O_249,N_2909,N_2898);
nand UO_250 (O_250,N_2832,N_2860);
nand UO_251 (O_251,N_2893,N_2873);
and UO_252 (O_252,N_2878,N_2944);
or UO_253 (O_253,N_2946,N_2931);
or UO_254 (O_254,N_2989,N_2900);
nor UO_255 (O_255,N_2947,N_2852);
nand UO_256 (O_256,N_2908,N_2976);
nor UO_257 (O_257,N_2862,N_2823);
nand UO_258 (O_258,N_2926,N_2946);
and UO_259 (O_259,N_2956,N_2935);
and UO_260 (O_260,N_2963,N_2837);
nor UO_261 (O_261,N_2995,N_2845);
and UO_262 (O_262,N_2900,N_2850);
or UO_263 (O_263,N_2950,N_2813);
nor UO_264 (O_264,N_2826,N_2965);
or UO_265 (O_265,N_2807,N_2885);
and UO_266 (O_266,N_2996,N_2890);
nor UO_267 (O_267,N_2901,N_2816);
nor UO_268 (O_268,N_2933,N_2957);
nor UO_269 (O_269,N_2860,N_2983);
nor UO_270 (O_270,N_2912,N_2830);
nor UO_271 (O_271,N_2843,N_2834);
or UO_272 (O_272,N_2912,N_2874);
nor UO_273 (O_273,N_2861,N_2984);
or UO_274 (O_274,N_2818,N_2944);
nand UO_275 (O_275,N_2985,N_2951);
xor UO_276 (O_276,N_2999,N_2806);
and UO_277 (O_277,N_2864,N_2975);
and UO_278 (O_278,N_2824,N_2809);
and UO_279 (O_279,N_2892,N_2904);
nand UO_280 (O_280,N_2824,N_2946);
or UO_281 (O_281,N_2839,N_2999);
and UO_282 (O_282,N_2992,N_2896);
or UO_283 (O_283,N_2878,N_2925);
nor UO_284 (O_284,N_2884,N_2831);
and UO_285 (O_285,N_2852,N_2854);
nand UO_286 (O_286,N_2905,N_2990);
and UO_287 (O_287,N_2914,N_2843);
and UO_288 (O_288,N_2917,N_2850);
and UO_289 (O_289,N_2884,N_2895);
nand UO_290 (O_290,N_2864,N_2808);
and UO_291 (O_291,N_2919,N_2993);
nand UO_292 (O_292,N_2897,N_2914);
and UO_293 (O_293,N_2832,N_2813);
nand UO_294 (O_294,N_2926,N_2954);
nand UO_295 (O_295,N_2980,N_2945);
or UO_296 (O_296,N_2851,N_2995);
or UO_297 (O_297,N_2936,N_2903);
and UO_298 (O_298,N_2974,N_2966);
nand UO_299 (O_299,N_2827,N_2833);
nand UO_300 (O_300,N_2848,N_2830);
or UO_301 (O_301,N_2997,N_2864);
nand UO_302 (O_302,N_2828,N_2995);
nand UO_303 (O_303,N_2991,N_2848);
and UO_304 (O_304,N_2842,N_2906);
or UO_305 (O_305,N_2882,N_2879);
nand UO_306 (O_306,N_2866,N_2887);
nor UO_307 (O_307,N_2947,N_2921);
nand UO_308 (O_308,N_2907,N_2806);
nand UO_309 (O_309,N_2994,N_2822);
nor UO_310 (O_310,N_2914,N_2932);
and UO_311 (O_311,N_2881,N_2807);
or UO_312 (O_312,N_2876,N_2882);
and UO_313 (O_313,N_2936,N_2908);
or UO_314 (O_314,N_2837,N_2918);
or UO_315 (O_315,N_2955,N_2834);
or UO_316 (O_316,N_2925,N_2840);
and UO_317 (O_317,N_2917,N_2977);
nand UO_318 (O_318,N_2947,N_2970);
and UO_319 (O_319,N_2880,N_2840);
and UO_320 (O_320,N_2873,N_2803);
xnor UO_321 (O_321,N_2937,N_2826);
nand UO_322 (O_322,N_2929,N_2940);
nand UO_323 (O_323,N_2993,N_2937);
and UO_324 (O_324,N_2832,N_2926);
or UO_325 (O_325,N_2928,N_2875);
nor UO_326 (O_326,N_2866,N_2982);
or UO_327 (O_327,N_2800,N_2981);
xnor UO_328 (O_328,N_2907,N_2986);
and UO_329 (O_329,N_2944,N_2924);
nand UO_330 (O_330,N_2898,N_2896);
nand UO_331 (O_331,N_2899,N_2931);
nor UO_332 (O_332,N_2939,N_2866);
or UO_333 (O_333,N_2832,N_2909);
or UO_334 (O_334,N_2841,N_2970);
and UO_335 (O_335,N_2871,N_2912);
or UO_336 (O_336,N_2805,N_2959);
nor UO_337 (O_337,N_2896,N_2883);
or UO_338 (O_338,N_2923,N_2843);
nor UO_339 (O_339,N_2963,N_2809);
or UO_340 (O_340,N_2880,N_2946);
nor UO_341 (O_341,N_2985,N_2828);
or UO_342 (O_342,N_2836,N_2884);
nand UO_343 (O_343,N_2943,N_2919);
xor UO_344 (O_344,N_2850,N_2839);
and UO_345 (O_345,N_2962,N_2802);
and UO_346 (O_346,N_2939,N_2873);
and UO_347 (O_347,N_2885,N_2848);
and UO_348 (O_348,N_2868,N_2857);
or UO_349 (O_349,N_2909,N_2860);
nand UO_350 (O_350,N_2833,N_2920);
and UO_351 (O_351,N_2915,N_2996);
and UO_352 (O_352,N_2810,N_2815);
nand UO_353 (O_353,N_2942,N_2994);
or UO_354 (O_354,N_2970,N_2938);
or UO_355 (O_355,N_2873,N_2971);
and UO_356 (O_356,N_2992,N_2908);
and UO_357 (O_357,N_2978,N_2957);
nor UO_358 (O_358,N_2808,N_2995);
nor UO_359 (O_359,N_2906,N_2959);
or UO_360 (O_360,N_2882,N_2921);
and UO_361 (O_361,N_2964,N_2841);
nor UO_362 (O_362,N_2888,N_2876);
or UO_363 (O_363,N_2996,N_2809);
nor UO_364 (O_364,N_2909,N_2831);
nor UO_365 (O_365,N_2854,N_2853);
nand UO_366 (O_366,N_2916,N_2953);
nor UO_367 (O_367,N_2964,N_2806);
nor UO_368 (O_368,N_2831,N_2961);
and UO_369 (O_369,N_2836,N_2946);
nor UO_370 (O_370,N_2927,N_2803);
and UO_371 (O_371,N_2891,N_2974);
nand UO_372 (O_372,N_2801,N_2903);
nand UO_373 (O_373,N_2992,N_2811);
nor UO_374 (O_374,N_2987,N_2827);
nor UO_375 (O_375,N_2833,N_2880);
nor UO_376 (O_376,N_2912,N_2930);
or UO_377 (O_377,N_2850,N_2843);
or UO_378 (O_378,N_2937,N_2815);
or UO_379 (O_379,N_2977,N_2967);
xor UO_380 (O_380,N_2932,N_2964);
and UO_381 (O_381,N_2927,N_2982);
and UO_382 (O_382,N_2931,N_2861);
or UO_383 (O_383,N_2939,N_2841);
nand UO_384 (O_384,N_2912,N_2989);
and UO_385 (O_385,N_2832,N_2898);
nor UO_386 (O_386,N_2962,N_2848);
and UO_387 (O_387,N_2934,N_2881);
nor UO_388 (O_388,N_2890,N_2808);
or UO_389 (O_389,N_2975,N_2932);
or UO_390 (O_390,N_2835,N_2886);
nor UO_391 (O_391,N_2987,N_2865);
or UO_392 (O_392,N_2969,N_2907);
and UO_393 (O_393,N_2830,N_2875);
nor UO_394 (O_394,N_2956,N_2881);
or UO_395 (O_395,N_2905,N_2940);
or UO_396 (O_396,N_2951,N_2863);
and UO_397 (O_397,N_2833,N_2875);
nand UO_398 (O_398,N_2813,N_2821);
nor UO_399 (O_399,N_2820,N_2917);
nand UO_400 (O_400,N_2949,N_2961);
nor UO_401 (O_401,N_2989,N_2830);
and UO_402 (O_402,N_2849,N_2868);
nor UO_403 (O_403,N_2801,N_2861);
nor UO_404 (O_404,N_2966,N_2921);
or UO_405 (O_405,N_2886,N_2929);
nor UO_406 (O_406,N_2915,N_2824);
nand UO_407 (O_407,N_2954,N_2816);
nor UO_408 (O_408,N_2832,N_2983);
xor UO_409 (O_409,N_2817,N_2898);
and UO_410 (O_410,N_2832,N_2852);
or UO_411 (O_411,N_2941,N_2850);
and UO_412 (O_412,N_2828,N_2826);
or UO_413 (O_413,N_2998,N_2970);
or UO_414 (O_414,N_2906,N_2875);
nand UO_415 (O_415,N_2969,N_2873);
nand UO_416 (O_416,N_2986,N_2888);
nor UO_417 (O_417,N_2831,N_2927);
nand UO_418 (O_418,N_2883,N_2982);
nand UO_419 (O_419,N_2827,N_2928);
nor UO_420 (O_420,N_2816,N_2810);
or UO_421 (O_421,N_2920,N_2903);
nand UO_422 (O_422,N_2824,N_2813);
nand UO_423 (O_423,N_2884,N_2958);
or UO_424 (O_424,N_2983,N_2801);
nor UO_425 (O_425,N_2880,N_2998);
and UO_426 (O_426,N_2996,N_2917);
or UO_427 (O_427,N_2898,N_2889);
nor UO_428 (O_428,N_2953,N_2819);
or UO_429 (O_429,N_2981,N_2899);
nand UO_430 (O_430,N_2969,N_2860);
nor UO_431 (O_431,N_2965,N_2861);
nor UO_432 (O_432,N_2987,N_2975);
and UO_433 (O_433,N_2805,N_2884);
or UO_434 (O_434,N_2911,N_2985);
or UO_435 (O_435,N_2842,N_2845);
or UO_436 (O_436,N_2847,N_2805);
nor UO_437 (O_437,N_2908,N_2930);
nand UO_438 (O_438,N_2828,N_2926);
xnor UO_439 (O_439,N_2988,N_2925);
or UO_440 (O_440,N_2855,N_2934);
nor UO_441 (O_441,N_2846,N_2943);
and UO_442 (O_442,N_2964,N_2937);
nor UO_443 (O_443,N_2893,N_2919);
and UO_444 (O_444,N_2884,N_2985);
nand UO_445 (O_445,N_2899,N_2883);
nor UO_446 (O_446,N_2803,N_2936);
or UO_447 (O_447,N_2889,N_2807);
nor UO_448 (O_448,N_2920,N_2959);
or UO_449 (O_449,N_2848,N_2936);
and UO_450 (O_450,N_2844,N_2977);
or UO_451 (O_451,N_2918,N_2853);
nor UO_452 (O_452,N_2969,N_2904);
nand UO_453 (O_453,N_2846,N_2915);
xnor UO_454 (O_454,N_2863,N_2838);
or UO_455 (O_455,N_2877,N_2956);
and UO_456 (O_456,N_2847,N_2905);
xor UO_457 (O_457,N_2880,N_2951);
and UO_458 (O_458,N_2815,N_2903);
and UO_459 (O_459,N_2812,N_2962);
or UO_460 (O_460,N_2863,N_2857);
or UO_461 (O_461,N_2850,N_2913);
nand UO_462 (O_462,N_2849,N_2965);
and UO_463 (O_463,N_2846,N_2881);
nor UO_464 (O_464,N_2867,N_2825);
nand UO_465 (O_465,N_2806,N_2886);
or UO_466 (O_466,N_2812,N_2823);
and UO_467 (O_467,N_2811,N_2843);
or UO_468 (O_468,N_2803,N_2889);
nor UO_469 (O_469,N_2930,N_2994);
nand UO_470 (O_470,N_2890,N_2820);
or UO_471 (O_471,N_2972,N_2832);
or UO_472 (O_472,N_2869,N_2981);
and UO_473 (O_473,N_2920,N_2852);
or UO_474 (O_474,N_2981,N_2885);
or UO_475 (O_475,N_2983,N_2952);
or UO_476 (O_476,N_2913,N_2838);
nor UO_477 (O_477,N_2912,N_2945);
nor UO_478 (O_478,N_2887,N_2871);
and UO_479 (O_479,N_2966,N_2811);
or UO_480 (O_480,N_2874,N_2913);
or UO_481 (O_481,N_2810,N_2896);
nand UO_482 (O_482,N_2965,N_2997);
or UO_483 (O_483,N_2820,N_2838);
xnor UO_484 (O_484,N_2890,N_2829);
or UO_485 (O_485,N_2870,N_2985);
nor UO_486 (O_486,N_2986,N_2841);
and UO_487 (O_487,N_2896,N_2820);
and UO_488 (O_488,N_2912,N_2896);
and UO_489 (O_489,N_2898,N_2892);
and UO_490 (O_490,N_2808,N_2812);
nand UO_491 (O_491,N_2929,N_2830);
xnor UO_492 (O_492,N_2949,N_2979);
nor UO_493 (O_493,N_2931,N_2901);
nor UO_494 (O_494,N_2865,N_2870);
nor UO_495 (O_495,N_2995,N_2926);
and UO_496 (O_496,N_2975,N_2803);
or UO_497 (O_497,N_2827,N_2992);
nor UO_498 (O_498,N_2846,N_2910);
or UO_499 (O_499,N_2887,N_2909);
endmodule