module basic_500_3000_500_3_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_61,In_146);
or U1 (N_1,In_113,In_463);
nand U2 (N_2,In_465,In_181);
or U3 (N_3,In_459,In_250);
nand U4 (N_4,In_353,In_243);
nor U5 (N_5,In_97,In_110);
nand U6 (N_6,In_211,In_68);
or U7 (N_7,In_261,In_185);
nor U8 (N_8,In_258,In_270);
and U9 (N_9,In_107,In_182);
nor U10 (N_10,In_260,In_143);
nor U11 (N_11,In_288,In_118);
and U12 (N_12,In_10,In_434);
nand U13 (N_13,In_452,In_173);
nor U14 (N_14,In_318,In_282);
nor U15 (N_15,In_404,In_160);
nand U16 (N_16,In_251,In_338);
nand U17 (N_17,In_73,In_219);
and U18 (N_18,In_337,In_429);
or U19 (N_19,In_9,In_153);
and U20 (N_20,In_364,In_58);
and U21 (N_21,In_204,In_474);
and U22 (N_22,In_319,In_16);
nor U23 (N_23,In_191,In_433);
nand U24 (N_24,In_129,In_169);
and U25 (N_25,In_460,In_451);
and U26 (N_26,In_327,In_490);
or U27 (N_27,In_131,In_362);
nor U28 (N_28,In_90,In_303);
and U29 (N_29,In_194,In_215);
and U30 (N_30,In_158,In_218);
nor U31 (N_31,In_388,In_144);
xnor U32 (N_32,In_438,In_343);
or U33 (N_33,In_128,In_398);
and U34 (N_34,In_187,In_467);
nand U35 (N_35,In_223,In_171);
nand U36 (N_36,In_83,In_120);
or U37 (N_37,In_381,In_385);
nor U38 (N_38,In_109,In_217);
or U39 (N_39,In_313,In_414);
and U40 (N_40,In_279,In_172);
or U41 (N_41,In_448,In_96);
nor U42 (N_42,In_111,In_70);
nand U43 (N_43,In_253,In_292);
nor U44 (N_44,In_401,In_55);
or U45 (N_45,In_254,In_415);
and U46 (N_46,In_491,In_0);
nor U47 (N_47,In_295,In_445);
and U48 (N_48,In_413,In_287);
and U49 (N_49,In_165,In_209);
nand U50 (N_50,In_48,In_168);
or U51 (N_51,In_389,In_375);
or U52 (N_52,In_267,In_477);
or U53 (N_53,In_486,In_485);
or U54 (N_54,In_115,In_36);
nand U55 (N_55,In_335,In_314);
nand U56 (N_56,In_371,In_345);
and U57 (N_57,In_259,In_102);
xnor U58 (N_58,In_37,In_59);
nand U59 (N_59,In_476,In_472);
or U60 (N_60,In_84,In_482);
or U61 (N_61,In_346,In_101);
nor U62 (N_62,In_207,In_344);
nor U63 (N_63,In_391,In_141);
nor U64 (N_64,In_22,In_149);
nor U65 (N_65,In_498,In_402);
xor U66 (N_66,In_213,In_376);
nand U67 (N_67,In_71,In_435);
nand U68 (N_68,In_306,In_138);
nand U69 (N_69,In_290,In_4);
nand U70 (N_70,In_273,In_432);
and U71 (N_71,In_237,In_315);
nand U72 (N_72,In_228,In_98);
or U73 (N_73,In_400,In_423);
nand U74 (N_74,In_457,In_492);
or U75 (N_75,In_12,In_24);
nand U76 (N_76,In_412,In_494);
or U77 (N_77,In_82,In_293);
or U78 (N_78,In_323,In_167);
nand U79 (N_79,In_57,In_67);
nor U80 (N_80,In_196,In_484);
and U81 (N_81,In_252,In_363);
nand U82 (N_82,In_195,In_33);
nand U83 (N_83,In_152,In_39);
nor U84 (N_84,In_235,In_332);
nor U85 (N_85,In_136,In_179);
and U86 (N_86,In_430,In_373);
or U87 (N_87,In_454,In_284);
xnor U88 (N_88,In_123,In_407);
or U89 (N_89,In_473,In_134);
and U90 (N_90,In_75,In_54);
nor U91 (N_91,In_446,In_236);
nor U92 (N_92,In_437,In_458);
nand U93 (N_93,In_379,In_221);
nor U94 (N_94,In_377,In_92);
and U95 (N_95,In_367,In_289);
and U96 (N_96,In_63,In_17);
or U97 (N_97,In_480,In_390);
nor U98 (N_98,In_66,In_244);
or U99 (N_99,In_25,In_21);
nor U100 (N_100,In_449,In_330);
or U101 (N_101,In_190,In_317);
nand U102 (N_102,In_62,In_368);
or U103 (N_103,In_140,In_359);
and U104 (N_104,In_495,In_424);
nand U105 (N_105,In_88,In_114);
nor U106 (N_106,In_122,In_208);
nor U107 (N_107,In_395,In_304);
or U108 (N_108,In_333,In_370);
and U109 (N_109,In_198,In_18);
or U110 (N_110,In_307,In_358);
and U111 (N_111,In_443,In_422);
and U112 (N_112,In_233,In_15);
nor U113 (N_113,In_72,In_489);
or U114 (N_114,In_366,In_47);
and U115 (N_115,In_226,In_431);
nand U116 (N_116,In_135,In_214);
or U117 (N_117,In_311,In_40);
nand U118 (N_118,In_483,In_188);
or U119 (N_119,In_369,In_89);
or U120 (N_120,In_447,In_297);
and U121 (N_121,In_356,In_283);
xnor U122 (N_122,In_103,In_340);
and U123 (N_123,In_155,In_41);
and U124 (N_124,In_268,In_466);
nor U125 (N_125,In_121,In_248);
and U126 (N_126,In_201,In_163);
nand U127 (N_127,In_200,In_99);
and U128 (N_128,In_20,In_199);
nor U129 (N_129,In_456,In_230);
nor U130 (N_130,In_396,In_420);
and U131 (N_131,In_79,In_210);
nand U132 (N_132,In_291,In_28);
nand U133 (N_133,In_387,In_416);
and U134 (N_134,In_372,In_23);
nand U135 (N_135,In_32,In_126);
nor U136 (N_136,In_357,In_76);
nor U137 (N_137,In_46,In_132);
nor U138 (N_138,In_108,In_475);
xnor U139 (N_139,In_440,In_471);
and U140 (N_140,In_334,In_321);
nand U141 (N_141,In_499,In_159);
or U142 (N_142,In_100,In_418);
nor U143 (N_143,In_139,In_7);
or U144 (N_144,In_453,In_470);
and U145 (N_145,In_352,In_350);
nand U146 (N_146,In_374,In_257);
nor U147 (N_147,In_479,In_240);
and U148 (N_148,In_275,In_50);
or U149 (N_149,In_239,In_203);
nor U150 (N_150,In_478,In_394);
and U151 (N_151,In_469,In_263);
xor U152 (N_152,In_180,In_410);
nand U153 (N_153,In_220,In_405);
or U154 (N_154,In_234,In_104);
xor U155 (N_155,In_302,In_316);
or U156 (N_156,In_274,In_5);
nor U157 (N_157,In_427,In_74);
or U158 (N_158,In_80,In_52);
and U159 (N_159,In_308,In_409);
and U160 (N_160,In_51,In_331);
nand U161 (N_161,In_81,In_225);
or U162 (N_162,In_264,In_487);
and U163 (N_163,In_202,In_265);
and U164 (N_164,In_6,In_271);
or U165 (N_165,In_64,In_178);
xnor U166 (N_166,In_69,In_276);
nand U167 (N_167,In_497,In_266);
and U168 (N_168,In_269,In_241);
and U169 (N_169,In_309,In_148);
and U170 (N_170,In_162,In_324);
nand U171 (N_171,In_142,In_166);
or U172 (N_172,In_85,In_34);
xnor U173 (N_173,In_339,In_14);
nor U174 (N_174,In_382,In_384);
and U175 (N_175,In_300,In_13);
or U176 (N_176,In_326,In_247);
nor U177 (N_177,In_305,In_1);
or U178 (N_178,In_493,In_31);
nand U179 (N_179,In_496,In_176);
and U180 (N_180,In_53,In_329);
or U181 (N_181,In_42,In_127);
nand U182 (N_182,In_222,In_450);
nor U183 (N_183,In_193,In_238);
nor U184 (N_184,In_242,In_347);
nor U185 (N_185,In_245,In_2);
nor U186 (N_186,In_216,In_310);
nor U187 (N_187,In_137,In_403);
and U188 (N_188,In_78,In_19);
or U189 (N_189,In_278,In_86);
nand U190 (N_190,In_380,In_348);
nand U191 (N_191,In_154,In_355);
and U192 (N_192,In_299,In_232);
nand U193 (N_193,In_349,In_11);
or U194 (N_194,In_49,In_341);
and U195 (N_195,In_93,In_184);
or U196 (N_196,In_38,In_462);
nor U197 (N_197,In_189,In_481);
or U198 (N_198,In_45,In_336);
nor U199 (N_199,In_361,In_44);
nand U200 (N_200,In_43,In_322);
nor U201 (N_201,In_312,In_119);
and U202 (N_202,In_351,In_164);
nor U203 (N_203,In_262,In_112);
nand U204 (N_204,In_419,In_342);
nor U205 (N_205,In_325,In_227);
and U206 (N_206,In_212,In_392);
and U207 (N_207,In_436,In_393);
or U208 (N_208,In_426,In_170);
nand U209 (N_209,In_328,In_87);
nand U210 (N_210,In_125,In_124);
nand U211 (N_211,In_157,In_206);
nand U212 (N_212,In_183,In_105);
xor U213 (N_213,In_439,In_29);
and U214 (N_214,In_35,In_116);
or U215 (N_215,In_286,In_224);
xnor U216 (N_216,In_399,In_229);
or U217 (N_217,In_147,In_91);
or U218 (N_218,In_145,In_378);
nand U219 (N_219,In_417,In_175);
nand U220 (N_220,In_455,In_397);
nand U221 (N_221,In_360,In_280);
nand U222 (N_222,In_26,In_27);
nand U223 (N_223,In_272,In_186);
nor U224 (N_224,In_246,In_256);
or U225 (N_225,In_77,In_461);
nor U226 (N_226,In_161,In_386);
nor U227 (N_227,In_192,In_320);
nor U228 (N_228,In_8,In_277);
and U229 (N_229,In_408,In_285);
and U230 (N_230,In_177,In_464);
and U231 (N_231,In_205,In_174);
nor U232 (N_232,In_150,In_94);
or U233 (N_233,In_488,In_298);
and U234 (N_234,In_130,In_30);
nor U235 (N_235,In_249,In_95);
nor U236 (N_236,In_117,In_468);
nand U237 (N_237,In_151,In_133);
nand U238 (N_238,In_60,In_411);
nand U239 (N_239,In_106,In_406);
nor U240 (N_240,In_365,In_65);
or U241 (N_241,In_197,In_296);
nand U242 (N_242,In_421,In_231);
nor U243 (N_243,In_428,In_3);
or U244 (N_244,In_156,In_354);
nor U245 (N_245,In_281,In_294);
nor U246 (N_246,In_444,In_255);
or U247 (N_247,In_383,In_301);
nand U248 (N_248,In_425,In_56);
and U249 (N_249,In_442,In_441);
or U250 (N_250,In_114,In_170);
or U251 (N_251,In_69,In_402);
or U252 (N_252,In_11,In_20);
and U253 (N_253,In_336,In_448);
nand U254 (N_254,In_257,In_100);
or U255 (N_255,In_15,In_395);
nand U256 (N_256,In_385,In_322);
nor U257 (N_257,In_148,In_308);
nor U258 (N_258,In_185,In_367);
or U259 (N_259,In_195,In_21);
and U260 (N_260,In_397,In_350);
or U261 (N_261,In_402,In_337);
nor U262 (N_262,In_312,In_428);
nor U263 (N_263,In_443,In_332);
or U264 (N_264,In_381,In_438);
and U265 (N_265,In_254,In_46);
or U266 (N_266,In_395,In_121);
nor U267 (N_267,In_366,In_499);
and U268 (N_268,In_63,In_324);
or U269 (N_269,In_42,In_348);
nand U270 (N_270,In_157,In_364);
nor U271 (N_271,In_371,In_115);
or U272 (N_272,In_316,In_406);
nand U273 (N_273,In_10,In_57);
or U274 (N_274,In_149,In_464);
and U275 (N_275,In_385,In_319);
or U276 (N_276,In_156,In_75);
or U277 (N_277,In_317,In_397);
nand U278 (N_278,In_337,In_345);
and U279 (N_279,In_119,In_146);
or U280 (N_280,In_445,In_47);
and U281 (N_281,In_266,In_97);
nand U282 (N_282,In_83,In_254);
nand U283 (N_283,In_353,In_193);
or U284 (N_284,In_37,In_185);
or U285 (N_285,In_109,In_346);
or U286 (N_286,In_171,In_465);
or U287 (N_287,In_450,In_414);
or U288 (N_288,In_12,In_342);
and U289 (N_289,In_82,In_84);
or U290 (N_290,In_197,In_394);
nor U291 (N_291,In_427,In_441);
nand U292 (N_292,In_337,In_103);
nand U293 (N_293,In_278,In_433);
xor U294 (N_294,In_381,In_464);
nand U295 (N_295,In_270,In_319);
xor U296 (N_296,In_409,In_313);
and U297 (N_297,In_340,In_368);
nand U298 (N_298,In_67,In_491);
nand U299 (N_299,In_281,In_8);
nand U300 (N_300,In_237,In_287);
or U301 (N_301,In_250,In_388);
or U302 (N_302,In_309,In_308);
nand U303 (N_303,In_164,In_76);
nand U304 (N_304,In_271,In_170);
nand U305 (N_305,In_298,In_237);
and U306 (N_306,In_441,In_322);
and U307 (N_307,In_44,In_193);
nor U308 (N_308,In_305,In_347);
and U309 (N_309,In_2,In_484);
and U310 (N_310,In_268,In_62);
or U311 (N_311,In_362,In_196);
and U312 (N_312,In_123,In_252);
nand U313 (N_313,In_12,In_107);
and U314 (N_314,In_223,In_422);
or U315 (N_315,In_263,In_94);
and U316 (N_316,In_7,In_314);
or U317 (N_317,In_368,In_121);
or U318 (N_318,In_400,In_36);
nor U319 (N_319,In_101,In_452);
and U320 (N_320,In_13,In_259);
nand U321 (N_321,In_389,In_41);
nand U322 (N_322,In_204,In_98);
nand U323 (N_323,In_141,In_32);
and U324 (N_324,In_357,In_474);
nand U325 (N_325,In_111,In_414);
and U326 (N_326,In_82,In_202);
and U327 (N_327,In_312,In_222);
or U328 (N_328,In_453,In_242);
nor U329 (N_329,In_369,In_51);
xor U330 (N_330,In_270,In_162);
nor U331 (N_331,In_6,In_147);
and U332 (N_332,In_176,In_412);
and U333 (N_333,In_141,In_377);
and U334 (N_334,In_450,In_348);
nand U335 (N_335,In_99,In_98);
or U336 (N_336,In_33,In_181);
nor U337 (N_337,In_251,In_86);
or U338 (N_338,In_214,In_330);
or U339 (N_339,In_413,In_427);
nand U340 (N_340,In_192,In_244);
nor U341 (N_341,In_367,In_477);
and U342 (N_342,In_149,In_368);
nor U343 (N_343,In_465,In_90);
and U344 (N_344,In_172,In_299);
and U345 (N_345,In_268,In_19);
nor U346 (N_346,In_449,In_172);
nor U347 (N_347,In_319,In_405);
nand U348 (N_348,In_327,In_315);
and U349 (N_349,In_101,In_278);
or U350 (N_350,In_43,In_194);
nand U351 (N_351,In_273,In_35);
and U352 (N_352,In_245,In_290);
or U353 (N_353,In_155,In_434);
nand U354 (N_354,In_401,In_14);
and U355 (N_355,In_129,In_497);
or U356 (N_356,In_85,In_137);
nor U357 (N_357,In_139,In_307);
or U358 (N_358,In_436,In_97);
or U359 (N_359,In_191,In_288);
or U360 (N_360,In_380,In_385);
nor U361 (N_361,In_8,In_395);
and U362 (N_362,In_272,In_400);
or U363 (N_363,In_245,In_202);
nand U364 (N_364,In_490,In_93);
nor U365 (N_365,In_189,In_371);
or U366 (N_366,In_264,In_47);
nor U367 (N_367,In_204,In_403);
or U368 (N_368,In_277,In_491);
nand U369 (N_369,In_229,In_30);
and U370 (N_370,In_372,In_234);
nor U371 (N_371,In_98,In_153);
nand U372 (N_372,In_177,In_495);
and U373 (N_373,In_93,In_119);
nand U374 (N_374,In_218,In_477);
and U375 (N_375,In_331,In_314);
nor U376 (N_376,In_190,In_9);
nand U377 (N_377,In_260,In_120);
and U378 (N_378,In_344,In_250);
nand U379 (N_379,In_392,In_131);
or U380 (N_380,In_367,In_108);
or U381 (N_381,In_106,In_497);
or U382 (N_382,In_124,In_264);
nor U383 (N_383,In_123,In_1);
and U384 (N_384,In_488,In_404);
nand U385 (N_385,In_436,In_341);
and U386 (N_386,In_37,In_222);
nor U387 (N_387,In_154,In_144);
nor U388 (N_388,In_186,In_125);
and U389 (N_389,In_466,In_484);
or U390 (N_390,In_243,In_124);
or U391 (N_391,In_363,In_455);
and U392 (N_392,In_307,In_308);
nand U393 (N_393,In_265,In_61);
nor U394 (N_394,In_39,In_105);
xnor U395 (N_395,In_217,In_302);
nor U396 (N_396,In_71,In_144);
nor U397 (N_397,In_40,In_456);
and U398 (N_398,In_164,In_5);
or U399 (N_399,In_491,In_163);
or U400 (N_400,In_191,In_468);
nand U401 (N_401,In_421,In_319);
nand U402 (N_402,In_424,In_310);
nor U403 (N_403,In_259,In_164);
and U404 (N_404,In_51,In_57);
or U405 (N_405,In_376,In_130);
xnor U406 (N_406,In_26,In_122);
and U407 (N_407,In_203,In_260);
and U408 (N_408,In_20,In_170);
and U409 (N_409,In_272,In_190);
nor U410 (N_410,In_263,In_416);
nand U411 (N_411,In_422,In_464);
or U412 (N_412,In_2,In_464);
nor U413 (N_413,In_153,In_131);
nor U414 (N_414,In_212,In_342);
nor U415 (N_415,In_186,In_375);
nand U416 (N_416,In_33,In_305);
nor U417 (N_417,In_40,In_186);
or U418 (N_418,In_301,In_179);
and U419 (N_419,In_15,In_419);
or U420 (N_420,In_304,In_71);
nand U421 (N_421,In_455,In_40);
or U422 (N_422,In_15,In_140);
nor U423 (N_423,In_91,In_468);
nor U424 (N_424,In_350,In_282);
xor U425 (N_425,In_7,In_413);
xor U426 (N_426,In_128,In_166);
nand U427 (N_427,In_279,In_167);
nor U428 (N_428,In_129,In_364);
or U429 (N_429,In_45,In_153);
nor U430 (N_430,In_260,In_224);
nor U431 (N_431,In_409,In_296);
nand U432 (N_432,In_199,In_336);
or U433 (N_433,In_85,In_6);
and U434 (N_434,In_199,In_291);
nor U435 (N_435,In_316,In_226);
nand U436 (N_436,In_32,In_248);
and U437 (N_437,In_352,In_255);
or U438 (N_438,In_429,In_219);
nor U439 (N_439,In_370,In_156);
nand U440 (N_440,In_489,In_103);
nor U441 (N_441,In_255,In_224);
nor U442 (N_442,In_431,In_316);
nand U443 (N_443,In_398,In_247);
or U444 (N_444,In_25,In_55);
nand U445 (N_445,In_144,In_378);
and U446 (N_446,In_286,In_258);
and U447 (N_447,In_203,In_401);
and U448 (N_448,In_52,In_317);
nor U449 (N_449,In_280,In_187);
nor U450 (N_450,In_70,In_326);
and U451 (N_451,In_397,In_235);
nand U452 (N_452,In_439,In_305);
and U453 (N_453,In_131,In_202);
or U454 (N_454,In_293,In_2);
or U455 (N_455,In_303,In_413);
and U456 (N_456,In_395,In_228);
or U457 (N_457,In_429,In_476);
nand U458 (N_458,In_347,In_268);
nand U459 (N_459,In_251,In_168);
nand U460 (N_460,In_253,In_299);
and U461 (N_461,In_275,In_82);
nand U462 (N_462,In_257,In_256);
nand U463 (N_463,In_49,In_307);
and U464 (N_464,In_95,In_214);
and U465 (N_465,In_33,In_308);
nor U466 (N_466,In_324,In_72);
nor U467 (N_467,In_371,In_65);
or U468 (N_468,In_238,In_276);
nand U469 (N_469,In_458,In_134);
nor U470 (N_470,In_459,In_163);
or U471 (N_471,In_99,In_114);
xor U472 (N_472,In_239,In_159);
nand U473 (N_473,In_361,In_6);
nor U474 (N_474,In_139,In_155);
nand U475 (N_475,In_489,In_207);
nor U476 (N_476,In_62,In_453);
nand U477 (N_477,In_437,In_247);
and U478 (N_478,In_376,In_77);
nor U479 (N_479,In_402,In_265);
or U480 (N_480,In_253,In_473);
or U481 (N_481,In_465,In_249);
and U482 (N_482,In_172,In_454);
nor U483 (N_483,In_421,In_481);
nor U484 (N_484,In_182,In_127);
or U485 (N_485,In_272,In_354);
and U486 (N_486,In_375,In_363);
nor U487 (N_487,In_25,In_459);
and U488 (N_488,In_392,In_252);
nor U489 (N_489,In_126,In_228);
xnor U490 (N_490,In_489,In_25);
nor U491 (N_491,In_464,In_383);
and U492 (N_492,In_43,In_464);
and U493 (N_493,In_462,In_155);
nand U494 (N_494,In_71,In_410);
or U495 (N_495,In_300,In_25);
or U496 (N_496,In_45,In_460);
and U497 (N_497,In_115,In_187);
nor U498 (N_498,In_255,In_486);
and U499 (N_499,In_384,In_238);
nor U500 (N_500,In_474,In_306);
and U501 (N_501,In_210,In_266);
or U502 (N_502,In_4,In_42);
nor U503 (N_503,In_437,In_428);
or U504 (N_504,In_181,In_241);
nand U505 (N_505,In_67,In_202);
nand U506 (N_506,In_198,In_429);
and U507 (N_507,In_119,In_394);
or U508 (N_508,In_157,In_132);
nor U509 (N_509,In_254,In_178);
and U510 (N_510,In_460,In_241);
nand U511 (N_511,In_336,In_172);
xor U512 (N_512,In_197,In_101);
nor U513 (N_513,In_10,In_439);
or U514 (N_514,In_314,In_95);
nor U515 (N_515,In_241,In_313);
nand U516 (N_516,In_43,In_287);
nand U517 (N_517,In_53,In_416);
nand U518 (N_518,In_421,In_369);
nor U519 (N_519,In_116,In_472);
nand U520 (N_520,In_208,In_138);
and U521 (N_521,In_147,In_157);
and U522 (N_522,In_276,In_158);
and U523 (N_523,In_440,In_398);
nand U524 (N_524,In_414,In_2);
and U525 (N_525,In_110,In_90);
and U526 (N_526,In_146,In_459);
or U527 (N_527,In_159,In_394);
nor U528 (N_528,In_22,In_431);
nor U529 (N_529,In_120,In_199);
and U530 (N_530,In_351,In_419);
or U531 (N_531,In_341,In_256);
nand U532 (N_532,In_5,In_344);
xnor U533 (N_533,In_401,In_5);
and U534 (N_534,In_13,In_403);
nor U535 (N_535,In_156,In_0);
nor U536 (N_536,In_141,In_487);
nand U537 (N_537,In_415,In_158);
nand U538 (N_538,In_436,In_269);
or U539 (N_539,In_231,In_68);
or U540 (N_540,In_340,In_483);
or U541 (N_541,In_140,In_244);
nand U542 (N_542,In_233,In_116);
nand U543 (N_543,In_138,In_236);
or U544 (N_544,In_101,In_325);
nor U545 (N_545,In_177,In_24);
xnor U546 (N_546,In_297,In_355);
nand U547 (N_547,In_329,In_67);
or U548 (N_548,In_379,In_281);
nand U549 (N_549,In_5,In_177);
or U550 (N_550,In_110,In_277);
nand U551 (N_551,In_183,In_123);
nand U552 (N_552,In_111,In_35);
nor U553 (N_553,In_428,In_302);
or U554 (N_554,In_488,In_34);
and U555 (N_555,In_266,In_101);
nand U556 (N_556,In_499,In_373);
nand U557 (N_557,In_307,In_54);
or U558 (N_558,In_257,In_442);
nand U559 (N_559,In_183,In_448);
nor U560 (N_560,In_161,In_199);
and U561 (N_561,In_65,In_4);
and U562 (N_562,In_173,In_17);
or U563 (N_563,In_494,In_9);
and U564 (N_564,In_254,In_268);
or U565 (N_565,In_327,In_24);
nor U566 (N_566,In_369,In_318);
nor U567 (N_567,In_372,In_449);
or U568 (N_568,In_48,In_314);
and U569 (N_569,In_450,In_191);
nor U570 (N_570,In_306,In_139);
and U571 (N_571,In_434,In_36);
nand U572 (N_572,In_73,In_206);
nor U573 (N_573,In_460,In_439);
nand U574 (N_574,In_228,In_91);
or U575 (N_575,In_335,In_395);
nand U576 (N_576,In_104,In_312);
and U577 (N_577,In_499,In_80);
nand U578 (N_578,In_475,In_146);
nor U579 (N_579,In_441,In_161);
nor U580 (N_580,In_389,In_210);
or U581 (N_581,In_390,In_294);
or U582 (N_582,In_99,In_432);
nor U583 (N_583,In_371,In_366);
nor U584 (N_584,In_450,In_285);
nor U585 (N_585,In_127,In_213);
and U586 (N_586,In_382,In_80);
nand U587 (N_587,In_151,In_177);
and U588 (N_588,In_304,In_2);
nand U589 (N_589,In_340,In_199);
and U590 (N_590,In_346,In_171);
and U591 (N_591,In_370,In_112);
nor U592 (N_592,In_108,In_221);
nand U593 (N_593,In_95,In_225);
nor U594 (N_594,In_120,In_102);
and U595 (N_595,In_371,In_448);
and U596 (N_596,In_63,In_469);
or U597 (N_597,In_236,In_164);
and U598 (N_598,In_364,In_70);
or U599 (N_599,In_151,In_293);
and U600 (N_600,In_127,In_484);
xnor U601 (N_601,In_495,In_114);
and U602 (N_602,In_377,In_61);
nor U603 (N_603,In_104,In_48);
nor U604 (N_604,In_198,In_107);
and U605 (N_605,In_272,In_373);
nor U606 (N_606,In_392,In_436);
and U607 (N_607,In_328,In_320);
or U608 (N_608,In_436,In_443);
and U609 (N_609,In_412,In_228);
or U610 (N_610,In_67,In_364);
or U611 (N_611,In_141,In_281);
or U612 (N_612,In_211,In_311);
or U613 (N_613,In_434,In_80);
and U614 (N_614,In_393,In_235);
nand U615 (N_615,In_332,In_471);
nor U616 (N_616,In_236,In_469);
and U617 (N_617,In_494,In_373);
or U618 (N_618,In_362,In_350);
nor U619 (N_619,In_403,In_188);
nand U620 (N_620,In_306,In_88);
or U621 (N_621,In_51,In_459);
and U622 (N_622,In_244,In_178);
or U623 (N_623,In_34,In_474);
nor U624 (N_624,In_214,In_179);
and U625 (N_625,In_54,In_291);
nor U626 (N_626,In_292,In_313);
or U627 (N_627,In_315,In_336);
or U628 (N_628,In_166,In_97);
and U629 (N_629,In_278,In_157);
or U630 (N_630,In_190,In_80);
and U631 (N_631,In_118,In_443);
and U632 (N_632,In_454,In_295);
or U633 (N_633,In_68,In_220);
and U634 (N_634,In_354,In_125);
or U635 (N_635,In_396,In_272);
nor U636 (N_636,In_99,In_81);
and U637 (N_637,In_321,In_274);
nand U638 (N_638,In_337,In_370);
or U639 (N_639,In_378,In_457);
and U640 (N_640,In_156,In_58);
nand U641 (N_641,In_139,In_122);
nor U642 (N_642,In_39,In_370);
nor U643 (N_643,In_210,In_137);
or U644 (N_644,In_351,In_353);
nor U645 (N_645,In_81,In_375);
or U646 (N_646,In_368,In_32);
and U647 (N_647,In_360,In_336);
and U648 (N_648,In_16,In_27);
and U649 (N_649,In_436,In_27);
nand U650 (N_650,In_16,In_216);
and U651 (N_651,In_40,In_38);
or U652 (N_652,In_115,In_71);
nand U653 (N_653,In_65,In_207);
or U654 (N_654,In_187,In_73);
and U655 (N_655,In_66,In_228);
nor U656 (N_656,In_401,In_105);
nand U657 (N_657,In_121,In_332);
and U658 (N_658,In_37,In_62);
nand U659 (N_659,In_103,In_288);
and U660 (N_660,In_173,In_449);
nor U661 (N_661,In_205,In_366);
or U662 (N_662,In_464,In_467);
nand U663 (N_663,In_180,In_474);
xnor U664 (N_664,In_399,In_158);
and U665 (N_665,In_261,In_315);
and U666 (N_666,In_407,In_353);
nand U667 (N_667,In_479,In_454);
nand U668 (N_668,In_151,In_351);
nand U669 (N_669,In_29,In_224);
xor U670 (N_670,In_325,In_29);
nand U671 (N_671,In_446,In_215);
and U672 (N_672,In_274,In_121);
and U673 (N_673,In_239,In_287);
or U674 (N_674,In_174,In_422);
and U675 (N_675,In_318,In_46);
nor U676 (N_676,In_68,In_277);
and U677 (N_677,In_157,In_232);
nand U678 (N_678,In_294,In_429);
nor U679 (N_679,In_123,In_219);
nand U680 (N_680,In_175,In_127);
nor U681 (N_681,In_399,In_351);
and U682 (N_682,In_404,In_102);
and U683 (N_683,In_373,In_270);
or U684 (N_684,In_29,In_287);
nor U685 (N_685,In_345,In_481);
nand U686 (N_686,In_28,In_494);
and U687 (N_687,In_208,In_178);
and U688 (N_688,In_392,In_344);
nand U689 (N_689,In_153,In_305);
nor U690 (N_690,In_210,In_66);
and U691 (N_691,In_498,In_69);
nor U692 (N_692,In_474,In_325);
and U693 (N_693,In_429,In_335);
and U694 (N_694,In_348,In_38);
nor U695 (N_695,In_129,In_394);
and U696 (N_696,In_201,In_115);
or U697 (N_697,In_306,In_181);
nand U698 (N_698,In_437,In_116);
nor U699 (N_699,In_243,In_78);
or U700 (N_700,In_4,In_331);
and U701 (N_701,In_166,In_17);
and U702 (N_702,In_170,In_379);
nor U703 (N_703,In_310,In_26);
or U704 (N_704,In_354,In_186);
or U705 (N_705,In_399,In_276);
nor U706 (N_706,In_84,In_438);
nand U707 (N_707,In_139,In_262);
nor U708 (N_708,In_15,In_345);
nor U709 (N_709,In_388,In_67);
and U710 (N_710,In_265,In_326);
nand U711 (N_711,In_348,In_207);
or U712 (N_712,In_129,In_317);
nand U713 (N_713,In_137,In_294);
nand U714 (N_714,In_409,In_437);
nand U715 (N_715,In_197,In_270);
and U716 (N_716,In_416,In_484);
nand U717 (N_717,In_297,In_227);
nor U718 (N_718,In_443,In_322);
or U719 (N_719,In_350,In_60);
or U720 (N_720,In_121,In_379);
nor U721 (N_721,In_484,In_361);
and U722 (N_722,In_427,In_364);
nand U723 (N_723,In_78,In_418);
nand U724 (N_724,In_14,In_487);
or U725 (N_725,In_117,In_364);
nand U726 (N_726,In_406,In_245);
nand U727 (N_727,In_322,In_113);
nand U728 (N_728,In_337,In_460);
and U729 (N_729,In_148,In_304);
and U730 (N_730,In_462,In_316);
xor U731 (N_731,In_234,In_315);
nor U732 (N_732,In_429,In_439);
nor U733 (N_733,In_335,In_334);
nand U734 (N_734,In_85,In_19);
nor U735 (N_735,In_62,In_370);
or U736 (N_736,In_336,In_301);
nor U737 (N_737,In_276,In_271);
xor U738 (N_738,In_74,In_393);
xnor U739 (N_739,In_165,In_358);
and U740 (N_740,In_499,In_107);
and U741 (N_741,In_361,In_300);
and U742 (N_742,In_450,In_445);
and U743 (N_743,In_110,In_485);
or U744 (N_744,In_303,In_212);
and U745 (N_745,In_265,In_413);
nand U746 (N_746,In_35,In_414);
and U747 (N_747,In_461,In_6);
or U748 (N_748,In_90,In_21);
nor U749 (N_749,In_415,In_474);
and U750 (N_750,In_17,In_8);
and U751 (N_751,In_23,In_96);
or U752 (N_752,In_11,In_177);
or U753 (N_753,In_331,In_96);
and U754 (N_754,In_256,In_185);
and U755 (N_755,In_334,In_148);
nand U756 (N_756,In_181,In_175);
and U757 (N_757,In_115,In_372);
nand U758 (N_758,In_127,In_269);
nor U759 (N_759,In_491,In_14);
and U760 (N_760,In_453,In_1);
nor U761 (N_761,In_316,In_402);
and U762 (N_762,In_9,In_191);
and U763 (N_763,In_265,In_352);
or U764 (N_764,In_402,In_16);
nand U765 (N_765,In_177,In_153);
and U766 (N_766,In_116,In_238);
or U767 (N_767,In_62,In_257);
or U768 (N_768,In_26,In_433);
nand U769 (N_769,In_198,In_357);
nor U770 (N_770,In_62,In_352);
nand U771 (N_771,In_206,In_470);
and U772 (N_772,In_218,In_144);
nand U773 (N_773,In_423,In_63);
nand U774 (N_774,In_49,In_277);
nor U775 (N_775,In_226,In_495);
or U776 (N_776,In_247,In_432);
and U777 (N_777,In_2,In_309);
or U778 (N_778,In_348,In_137);
nor U779 (N_779,In_292,In_139);
nand U780 (N_780,In_69,In_270);
nor U781 (N_781,In_124,In_94);
and U782 (N_782,In_415,In_60);
nor U783 (N_783,In_320,In_421);
and U784 (N_784,In_292,In_61);
and U785 (N_785,In_172,In_244);
and U786 (N_786,In_392,In_102);
and U787 (N_787,In_198,In_287);
and U788 (N_788,In_59,In_19);
and U789 (N_789,In_235,In_270);
nand U790 (N_790,In_397,In_185);
nand U791 (N_791,In_408,In_199);
or U792 (N_792,In_405,In_15);
nand U793 (N_793,In_251,In_326);
or U794 (N_794,In_261,In_58);
nor U795 (N_795,In_69,In_499);
nand U796 (N_796,In_50,In_38);
and U797 (N_797,In_96,In_84);
and U798 (N_798,In_115,In_426);
or U799 (N_799,In_381,In_289);
nand U800 (N_800,In_138,In_2);
and U801 (N_801,In_48,In_396);
nor U802 (N_802,In_184,In_167);
or U803 (N_803,In_402,In_410);
and U804 (N_804,In_365,In_267);
nand U805 (N_805,In_19,In_410);
or U806 (N_806,In_279,In_421);
nor U807 (N_807,In_322,In_26);
nor U808 (N_808,In_236,In_407);
nand U809 (N_809,In_226,In_346);
and U810 (N_810,In_416,In_371);
or U811 (N_811,In_199,In_167);
or U812 (N_812,In_454,In_234);
nand U813 (N_813,In_322,In_334);
and U814 (N_814,In_389,In_343);
nand U815 (N_815,In_156,In_465);
nor U816 (N_816,In_428,In_65);
nand U817 (N_817,In_7,In_410);
and U818 (N_818,In_98,In_252);
nor U819 (N_819,In_33,In_134);
and U820 (N_820,In_411,In_215);
nand U821 (N_821,In_406,In_67);
nand U822 (N_822,In_181,In_270);
or U823 (N_823,In_411,In_369);
nor U824 (N_824,In_7,In_405);
and U825 (N_825,In_203,In_410);
nor U826 (N_826,In_142,In_66);
nor U827 (N_827,In_15,In_454);
and U828 (N_828,In_285,In_277);
and U829 (N_829,In_113,In_269);
and U830 (N_830,In_175,In_236);
or U831 (N_831,In_85,In_11);
and U832 (N_832,In_384,In_493);
nand U833 (N_833,In_53,In_83);
and U834 (N_834,In_110,In_397);
nand U835 (N_835,In_252,In_142);
nor U836 (N_836,In_448,In_292);
or U837 (N_837,In_164,In_387);
nor U838 (N_838,In_45,In_306);
nand U839 (N_839,In_334,In_199);
nand U840 (N_840,In_331,In_35);
or U841 (N_841,In_456,In_368);
and U842 (N_842,In_55,In_68);
xor U843 (N_843,In_319,In_133);
or U844 (N_844,In_408,In_365);
or U845 (N_845,In_245,In_369);
or U846 (N_846,In_59,In_395);
nor U847 (N_847,In_226,In_361);
nor U848 (N_848,In_342,In_106);
xor U849 (N_849,In_490,In_401);
or U850 (N_850,In_305,In_40);
and U851 (N_851,In_454,In_265);
nand U852 (N_852,In_141,In_237);
nor U853 (N_853,In_489,In_70);
nor U854 (N_854,In_197,In_116);
nor U855 (N_855,In_257,In_485);
xor U856 (N_856,In_25,In_233);
nand U857 (N_857,In_183,In_211);
or U858 (N_858,In_450,In_161);
xor U859 (N_859,In_363,In_347);
or U860 (N_860,In_26,In_181);
nor U861 (N_861,In_366,In_187);
and U862 (N_862,In_176,In_277);
and U863 (N_863,In_430,In_128);
and U864 (N_864,In_355,In_83);
and U865 (N_865,In_68,In_315);
and U866 (N_866,In_280,In_203);
xnor U867 (N_867,In_462,In_296);
and U868 (N_868,In_170,In_262);
nand U869 (N_869,In_284,In_32);
nand U870 (N_870,In_441,In_274);
or U871 (N_871,In_3,In_137);
nor U872 (N_872,In_94,In_494);
and U873 (N_873,In_484,In_265);
nor U874 (N_874,In_57,In_288);
xor U875 (N_875,In_456,In_444);
nand U876 (N_876,In_77,In_335);
nand U877 (N_877,In_60,In_402);
or U878 (N_878,In_208,In_492);
nand U879 (N_879,In_108,In_252);
or U880 (N_880,In_283,In_489);
and U881 (N_881,In_54,In_62);
nor U882 (N_882,In_352,In_103);
or U883 (N_883,In_24,In_283);
nand U884 (N_884,In_415,In_76);
nand U885 (N_885,In_394,In_267);
or U886 (N_886,In_179,In_209);
or U887 (N_887,In_320,In_317);
and U888 (N_888,In_390,In_142);
and U889 (N_889,In_7,In_53);
nand U890 (N_890,In_73,In_130);
and U891 (N_891,In_354,In_169);
and U892 (N_892,In_62,In_333);
and U893 (N_893,In_426,In_490);
nor U894 (N_894,In_363,In_422);
xor U895 (N_895,In_173,In_160);
and U896 (N_896,In_7,In_282);
nand U897 (N_897,In_332,In_183);
nor U898 (N_898,In_58,In_128);
or U899 (N_899,In_482,In_113);
nor U900 (N_900,In_145,In_485);
nor U901 (N_901,In_483,In_165);
nand U902 (N_902,In_383,In_355);
or U903 (N_903,In_67,In_294);
nand U904 (N_904,In_225,In_344);
or U905 (N_905,In_150,In_470);
nand U906 (N_906,In_100,In_373);
and U907 (N_907,In_71,In_182);
nand U908 (N_908,In_213,In_362);
and U909 (N_909,In_45,In_344);
nor U910 (N_910,In_381,In_104);
and U911 (N_911,In_233,In_23);
and U912 (N_912,In_431,In_349);
and U913 (N_913,In_319,In_397);
or U914 (N_914,In_201,In_478);
or U915 (N_915,In_490,In_231);
xnor U916 (N_916,In_200,In_250);
or U917 (N_917,In_466,In_169);
nor U918 (N_918,In_287,In_33);
nand U919 (N_919,In_346,In_282);
nor U920 (N_920,In_48,In_185);
and U921 (N_921,In_237,In_158);
and U922 (N_922,In_214,In_393);
nand U923 (N_923,In_419,In_181);
nand U924 (N_924,In_408,In_434);
and U925 (N_925,In_84,In_443);
or U926 (N_926,In_441,In_360);
or U927 (N_927,In_183,In_478);
nand U928 (N_928,In_329,In_495);
nor U929 (N_929,In_212,In_489);
or U930 (N_930,In_34,In_326);
nor U931 (N_931,In_455,In_435);
and U932 (N_932,In_144,In_402);
nand U933 (N_933,In_67,In_209);
nand U934 (N_934,In_423,In_32);
or U935 (N_935,In_46,In_390);
or U936 (N_936,In_8,In_241);
nor U937 (N_937,In_357,In_169);
nor U938 (N_938,In_452,In_106);
and U939 (N_939,In_175,In_102);
and U940 (N_940,In_159,In_285);
or U941 (N_941,In_345,In_347);
or U942 (N_942,In_54,In_156);
or U943 (N_943,In_257,In_117);
nand U944 (N_944,In_215,In_294);
nor U945 (N_945,In_432,In_23);
and U946 (N_946,In_469,In_305);
and U947 (N_947,In_157,In_489);
xor U948 (N_948,In_6,In_254);
or U949 (N_949,In_320,In_249);
and U950 (N_950,In_431,In_193);
nand U951 (N_951,In_302,In_378);
and U952 (N_952,In_145,In_143);
nor U953 (N_953,In_464,In_425);
nor U954 (N_954,In_391,In_271);
and U955 (N_955,In_13,In_400);
and U956 (N_956,In_275,In_62);
nand U957 (N_957,In_18,In_213);
or U958 (N_958,In_351,In_160);
xor U959 (N_959,In_319,In_131);
nand U960 (N_960,In_352,In_438);
or U961 (N_961,In_368,In_258);
and U962 (N_962,In_285,In_337);
and U963 (N_963,In_69,In_110);
or U964 (N_964,In_401,In_377);
nor U965 (N_965,In_209,In_81);
and U966 (N_966,In_348,In_286);
or U967 (N_967,In_53,In_209);
nand U968 (N_968,In_10,In_363);
nand U969 (N_969,In_132,In_285);
or U970 (N_970,In_301,In_78);
nor U971 (N_971,In_333,In_37);
nor U972 (N_972,In_327,In_298);
or U973 (N_973,In_67,In_445);
nand U974 (N_974,In_493,In_379);
and U975 (N_975,In_434,In_362);
nand U976 (N_976,In_406,In_495);
nor U977 (N_977,In_38,In_129);
nor U978 (N_978,In_391,In_337);
nand U979 (N_979,In_409,In_89);
nand U980 (N_980,In_185,In_8);
nand U981 (N_981,In_469,In_269);
and U982 (N_982,In_154,In_78);
and U983 (N_983,In_410,In_63);
or U984 (N_984,In_344,In_412);
nor U985 (N_985,In_210,In_96);
nor U986 (N_986,In_148,In_433);
and U987 (N_987,In_59,In_51);
or U988 (N_988,In_459,In_252);
nor U989 (N_989,In_1,In_179);
and U990 (N_990,In_67,In_371);
or U991 (N_991,In_428,In_106);
nand U992 (N_992,In_417,In_118);
or U993 (N_993,In_59,In_461);
and U994 (N_994,In_99,In_145);
or U995 (N_995,In_151,In_135);
nor U996 (N_996,In_458,In_122);
and U997 (N_997,In_445,In_433);
and U998 (N_998,In_180,In_342);
xor U999 (N_999,In_165,In_328);
nand U1000 (N_1000,N_741,N_202);
or U1001 (N_1001,N_31,N_439);
or U1002 (N_1002,N_615,N_375);
nand U1003 (N_1003,N_938,N_595);
nor U1004 (N_1004,N_292,N_896);
nand U1005 (N_1005,N_980,N_672);
or U1006 (N_1006,N_951,N_817);
nand U1007 (N_1007,N_689,N_102);
nor U1008 (N_1008,N_236,N_855);
and U1009 (N_1009,N_631,N_358);
nand U1010 (N_1010,N_321,N_420);
or U1011 (N_1011,N_942,N_688);
nand U1012 (N_1012,N_758,N_536);
or U1013 (N_1013,N_651,N_493);
and U1014 (N_1014,N_281,N_393);
or U1015 (N_1015,N_655,N_422);
nand U1016 (N_1016,N_490,N_796);
or U1017 (N_1017,N_242,N_440);
nand U1018 (N_1018,N_705,N_154);
or U1019 (N_1019,N_526,N_497);
nor U1020 (N_1020,N_240,N_710);
nor U1021 (N_1021,N_157,N_426);
nand U1022 (N_1022,N_712,N_891);
or U1023 (N_1023,N_153,N_419);
nor U1024 (N_1024,N_427,N_706);
nor U1025 (N_1025,N_748,N_642);
or U1026 (N_1026,N_830,N_747);
nor U1027 (N_1027,N_895,N_336);
nor U1028 (N_1028,N_786,N_926);
or U1029 (N_1029,N_750,N_108);
nor U1030 (N_1030,N_367,N_607);
or U1031 (N_1031,N_789,N_576);
nand U1032 (N_1032,N_871,N_775);
nor U1033 (N_1033,N_990,N_673);
and U1034 (N_1034,N_838,N_144);
nand U1035 (N_1035,N_67,N_351);
or U1036 (N_1036,N_355,N_88);
nor U1037 (N_1037,N_235,N_64);
nor U1038 (N_1038,N_380,N_40);
and U1039 (N_1039,N_641,N_908);
or U1040 (N_1040,N_658,N_620);
nand U1041 (N_1041,N_720,N_514);
nor U1042 (N_1042,N_289,N_820);
nand U1043 (N_1043,N_209,N_975);
nor U1044 (N_1044,N_774,N_32);
or U1045 (N_1045,N_145,N_928);
nand U1046 (N_1046,N_643,N_534);
or U1047 (N_1047,N_294,N_208);
or U1048 (N_1048,N_234,N_508);
nand U1049 (N_1049,N_738,N_33);
and U1050 (N_1050,N_918,N_396);
or U1051 (N_1051,N_905,N_379);
or U1052 (N_1052,N_699,N_737);
or U1053 (N_1053,N_589,N_191);
or U1054 (N_1054,N_310,N_695);
nor U1055 (N_1055,N_877,N_499);
nor U1056 (N_1056,N_487,N_99);
and U1057 (N_1057,N_256,N_834);
xnor U1058 (N_1058,N_482,N_697);
nor U1059 (N_1059,N_225,N_219);
nor U1060 (N_1060,N_403,N_561);
nand U1061 (N_1061,N_185,N_765);
xnor U1062 (N_1062,N_1,N_611);
or U1063 (N_1063,N_675,N_100);
nand U1064 (N_1064,N_696,N_46);
nand U1065 (N_1065,N_792,N_170);
or U1066 (N_1066,N_969,N_458);
nor U1067 (N_1067,N_199,N_733);
nor U1068 (N_1068,N_183,N_645);
and U1069 (N_1069,N_62,N_264);
and U1070 (N_1070,N_117,N_498);
nand U1071 (N_1071,N_684,N_198);
nor U1072 (N_1072,N_441,N_754);
and U1073 (N_1073,N_999,N_285);
or U1074 (N_1074,N_119,N_880);
or U1075 (N_1075,N_272,N_401);
or U1076 (N_1076,N_868,N_411);
nand U1077 (N_1077,N_172,N_38);
nor U1078 (N_1078,N_863,N_408);
and U1079 (N_1079,N_342,N_163);
and U1080 (N_1080,N_692,N_494);
nor U1081 (N_1081,N_448,N_939);
and U1082 (N_1082,N_110,N_557);
or U1083 (N_1083,N_174,N_715);
nand U1084 (N_1084,N_309,N_548);
and U1085 (N_1085,N_295,N_719);
or U1086 (N_1086,N_934,N_782);
or U1087 (N_1087,N_988,N_621);
and U1088 (N_1088,N_9,N_936);
nor U1089 (N_1089,N_146,N_878);
nand U1090 (N_1090,N_12,N_873);
and U1091 (N_1091,N_950,N_510);
nand U1092 (N_1092,N_237,N_231);
or U1093 (N_1093,N_843,N_276);
and U1094 (N_1094,N_676,N_43);
nand U1095 (N_1095,N_967,N_708);
and U1096 (N_1096,N_997,N_644);
nand U1097 (N_1097,N_280,N_86);
and U1098 (N_1098,N_524,N_727);
or U1099 (N_1099,N_192,N_619);
nor U1100 (N_1100,N_47,N_909);
or U1101 (N_1101,N_844,N_653);
nand U1102 (N_1102,N_160,N_654);
nand U1103 (N_1103,N_771,N_279);
nand U1104 (N_1104,N_543,N_109);
and U1105 (N_1105,N_34,N_17);
or U1106 (N_1106,N_244,N_884);
nand U1107 (N_1107,N_875,N_399);
xnor U1108 (N_1108,N_320,N_69);
or U1109 (N_1109,N_215,N_177);
nor U1110 (N_1110,N_204,N_666);
nand U1111 (N_1111,N_816,N_691);
nand U1112 (N_1112,N_565,N_2);
and U1113 (N_1113,N_386,N_663);
and U1114 (N_1114,N_932,N_155);
xnor U1115 (N_1115,N_677,N_790);
nand U1116 (N_1116,N_716,N_819);
nor U1117 (N_1117,N_943,N_468);
or U1118 (N_1118,N_729,N_753);
or U1119 (N_1119,N_679,N_520);
and U1120 (N_1120,N_196,N_89);
nor U1121 (N_1121,N_150,N_944);
nand U1122 (N_1122,N_70,N_869);
and U1123 (N_1123,N_555,N_913);
nor U1124 (N_1124,N_148,N_303);
or U1125 (N_1125,N_731,N_463);
nand U1126 (N_1126,N_897,N_904);
and U1127 (N_1127,N_372,N_232);
nor U1128 (N_1128,N_324,N_703);
or U1129 (N_1129,N_914,N_867);
nand U1130 (N_1130,N_718,N_63);
nand U1131 (N_1131,N_288,N_374);
nor U1132 (N_1132,N_349,N_728);
or U1133 (N_1133,N_559,N_362);
nand U1134 (N_1134,N_413,N_251);
or U1135 (N_1135,N_646,N_945);
or U1136 (N_1136,N_302,N_252);
xnor U1137 (N_1137,N_756,N_560);
or U1138 (N_1138,N_609,N_814);
nor U1139 (N_1139,N_888,N_533);
nand U1140 (N_1140,N_462,N_258);
xnor U1141 (N_1141,N_762,N_501);
and U1142 (N_1142,N_428,N_656);
or U1143 (N_1143,N_622,N_745);
nand U1144 (N_1144,N_120,N_392);
nor U1145 (N_1145,N_248,N_881);
nor U1146 (N_1146,N_902,N_356);
and U1147 (N_1147,N_261,N_734);
or U1148 (N_1148,N_637,N_469);
or U1149 (N_1149,N_767,N_348);
and U1150 (N_1150,N_485,N_958);
or U1151 (N_1151,N_424,N_903);
nand U1152 (N_1152,N_509,N_103);
and U1153 (N_1153,N_948,N_42);
nor U1154 (N_1154,N_532,N_801);
and U1155 (N_1155,N_805,N_492);
and U1156 (N_1156,N_769,N_152);
nand U1157 (N_1157,N_304,N_22);
or U1158 (N_1158,N_573,N_173);
and U1159 (N_1159,N_388,N_528);
nor U1160 (N_1160,N_13,N_981);
xor U1161 (N_1161,N_78,N_800);
or U1162 (N_1162,N_55,N_200);
and U1163 (N_1163,N_544,N_563);
nor U1164 (N_1164,N_373,N_466);
or U1165 (N_1165,N_478,N_243);
nand U1166 (N_1166,N_992,N_704);
xor U1167 (N_1167,N_553,N_887);
nor U1168 (N_1168,N_384,N_925);
nor U1169 (N_1169,N_118,N_898);
nor U1170 (N_1170,N_768,N_323);
nand U1171 (N_1171,N_591,N_278);
nand U1172 (N_1172,N_147,N_328);
or U1173 (N_1173,N_124,N_390);
and U1174 (N_1174,N_586,N_95);
nand U1175 (N_1175,N_125,N_452);
nor U1176 (N_1176,N_505,N_171);
or U1177 (N_1177,N_317,N_134);
nand U1178 (N_1178,N_851,N_450);
or U1179 (N_1179,N_29,N_343);
nand U1180 (N_1180,N_957,N_19);
nor U1181 (N_1181,N_389,N_860);
nor U1182 (N_1182,N_809,N_126);
nand U1183 (N_1183,N_203,N_847);
nand U1184 (N_1184,N_600,N_984);
and U1185 (N_1185,N_269,N_92);
nand U1186 (N_1186,N_812,N_841);
xnor U1187 (N_1187,N_977,N_305);
or U1188 (N_1188,N_636,N_395);
nand U1189 (N_1189,N_156,N_449);
nor U1190 (N_1190,N_971,N_588);
or U1191 (N_1191,N_111,N_791);
or U1192 (N_1192,N_26,N_484);
or U1193 (N_1193,N_723,N_453);
or U1194 (N_1194,N_630,N_569);
nor U1195 (N_1195,N_85,N_79);
and U1196 (N_1196,N_680,N_429);
nand U1197 (N_1197,N_854,N_283);
or U1198 (N_1198,N_810,N_24);
nor U1199 (N_1199,N_71,N_72);
and U1200 (N_1200,N_227,N_551);
nor U1201 (N_1201,N_836,N_973);
nor U1202 (N_1202,N_139,N_443);
or U1203 (N_1203,N_627,N_927);
nor U1204 (N_1204,N_430,N_730);
and U1205 (N_1205,N_333,N_832);
or U1206 (N_1206,N_787,N_23);
and U1207 (N_1207,N_341,N_955);
or U1208 (N_1208,N_385,N_923);
nand U1209 (N_1209,N_239,N_476);
or U1210 (N_1210,N_3,N_329);
xnor U1211 (N_1211,N_802,N_193);
nor U1212 (N_1212,N_477,N_907);
nor U1213 (N_1213,N_678,N_519);
or U1214 (N_1214,N_30,N_580);
nand U1215 (N_1215,N_364,N_725);
xor U1216 (N_1216,N_314,N_489);
and U1217 (N_1217,N_906,N_94);
or U1218 (N_1218,N_701,N_149);
and U1219 (N_1219,N_550,N_795);
nor U1220 (N_1220,N_217,N_601);
nor U1221 (N_1221,N_683,N_241);
and U1222 (N_1222,N_603,N_66);
nor U1223 (N_1223,N_178,N_371);
and U1224 (N_1224,N_82,N_604);
nor U1225 (N_1225,N_352,N_554);
nand U1226 (N_1226,N_978,N_121);
nand U1227 (N_1227,N_797,N_182);
and U1228 (N_1228,N_825,N_253);
or U1229 (N_1229,N_562,N_807);
or U1230 (N_1230,N_432,N_194);
or U1231 (N_1231,N_517,N_783);
and U1232 (N_1232,N_886,N_968);
nand U1233 (N_1233,N_518,N_598);
nor U1234 (N_1234,N_911,N_53);
xor U1235 (N_1235,N_872,N_436);
or U1236 (N_1236,N_97,N_665);
nand U1237 (N_1237,N_360,N_785);
nand U1238 (N_1238,N_639,N_531);
and U1239 (N_1239,N_540,N_625);
nor U1240 (N_1240,N_506,N_406);
nor U1241 (N_1241,N_274,N_77);
or U1242 (N_1242,N_267,N_180);
and U1243 (N_1243,N_931,N_27);
or U1244 (N_1244,N_381,N_457);
nor U1245 (N_1245,N_681,N_229);
nand U1246 (N_1246,N_254,N_87);
nor U1247 (N_1247,N_864,N_318);
nand U1248 (N_1248,N_726,N_579);
nor U1249 (N_1249,N_467,N_961);
or U1250 (N_1250,N_11,N_778);
and U1251 (N_1251,N_25,N_949);
nor U1252 (N_1252,N_83,N_35);
or U1253 (N_1253,N_45,N_915);
or U1254 (N_1254,N_410,N_512);
nor U1255 (N_1255,N_447,N_660);
nand U1256 (N_1256,N_599,N_165);
nor U1257 (N_1257,N_974,N_37);
nand U1258 (N_1258,N_255,N_52);
and U1259 (N_1259,N_885,N_772);
or U1260 (N_1260,N_434,N_0);
nor U1261 (N_1261,N_982,N_744);
nand U1262 (N_1262,N_166,N_585);
nand U1263 (N_1263,N_799,N_417);
or U1264 (N_1264,N_8,N_995);
nand U1265 (N_1265,N_670,N_921);
nand U1266 (N_1266,N_777,N_766);
or U1267 (N_1267,N_500,N_416);
nand U1268 (N_1268,N_14,N_284);
nor U1269 (N_1269,N_346,N_856);
or U1270 (N_1270,N_471,N_940);
nand U1271 (N_1271,N_142,N_287);
and U1272 (N_1272,N_488,N_865);
or U1273 (N_1273,N_634,N_788);
nor U1274 (N_1274,N_188,N_158);
and U1275 (N_1275,N_979,N_649);
and U1276 (N_1276,N_808,N_337);
and U1277 (N_1277,N_848,N_539);
or U1278 (N_1278,N_21,N_402);
and U1279 (N_1279,N_535,N_301);
nand U1280 (N_1280,N_291,N_542);
nor U1281 (N_1281,N_459,N_168);
nand U1282 (N_1282,N_404,N_347);
nand U1283 (N_1283,N_525,N_76);
nor U1284 (N_1284,N_567,N_889);
nand U1285 (N_1285,N_425,N_954);
and U1286 (N_1286,N_717,N_377);
and U1287 (N_1287,N_610,N_922);
or U1288 (N_1288,N_306,N_529);
nand U1289 (N_1289,N_376,N_818);
xor U1290 (N_1290,N_702,N_214);
or U1291 (N_1291,N_273,N_370);
and U1292 (N_1292,N_39,N_590);
nand U1293 (N_1293,N_41,N_138);
or U1294 (N_1294,N_275,N_763);
or U1295 (N_1295,N_319,N_835);
and U1296 (N_1296,N_104,N_455);
or U1297 (N_1297,N_826,N_44);
nor U1298 (N_1298,N_647,N_365);
nor U1299 (N_1299,N_749,N_136);
or U1300 (N_1300,N_823,N_472);
nand U1301 (N_1301,N_606,N_901);
or U1302 (N_1302,N_164,N_58);
nor U1303 (N_1303,N_614,N_549);
or U1304 (N_1304,N_986,N_594);
or U1305 (N_1305,N_249,N_547);
nand U1306 (N_1306,N_383,N_315);
nor U1307 (N_1307,N_828,N_616);
nand U1308 (N_1308,N_363,N_311);
or U1309 (N_1309,N_20,N_760);
and U1310 (N_1310,N_68,N_247);
nor U1311 (N_1311,N_238,N_857);
nand U1312 (N_1312,N_861,N_698);
or U1313 (N_1313,N_344,N_866);
nand U1314 (N_1314,N_369,N_228);
nand U1315 (N_1315,N_546,N_602);
nand U1316 (N_1316,N_740,N_205);
or U1317 (N_1317,N_206,N_690);
and U1318 (N_1318,N_815,N_659);
and U1319 (N_1319,N_596,N_127);
or U1320 (N_1320,N_211,N_822);
or U1321 (N_1321,N_299,N_475);
or U1322 (N_1322,N_359,N_521);
or U1323 (N_1323,N_956,N_640);
or U1324 (N_1324,N_582,N_638);
and U1325 (N_1325,N_798,N_724);
nor U1326 (N_1326,N_899,N_60);
and U1327 (N_1327,N_496,N_910);
or U1328 (N_1328,N_4,N_435);
or U1329 (N_1329,N_335,N_946);
nor U1330 (N_1330,N_538,N_963);
and U1331 (N_1331,N_972,N_858);
nand U1332 (N_1332,N_137,N_316);
or U1333 (N_1333,N_714,N_368);
nand U1334 (N_1334,N_423,N_779);
or U1335 (N_1335,N_587,N_57);
nor U1336 (N_1336,N_226,N_732);
nor U1337 (N_1337,N_98,N_132);
nor U1338 (N_1338,N_130,N_994);
nor U1339 (N_1339,N_378,N_507);
or U1340 (N_1340,N_633,N_128);
or U1341 (N_1341,N_682,N_743);
and U1342 (N_1342,N_742,N_755);
nor U1343 (N_1343,N_709,N_541);
and U1344 (N_1344,N_883,N_503);
or U1345 (N_1345,N_106,N_129);
or U1346 (N_1346,N_141,N_18);
and U1347 (N_1347,N_618,N_821);
nor U1348 (N_1348,N_220,N_387);
nor U1349 (N_1349,N_10,N_920);
or U1350 (N_1350,N_187,N_530);
or U1351 (N_1351,N_960,N_222);
nor U1352 (N_1352,N_407,N_876);
or U1353 (N_1353,N_652,N_929);
and U1354 (N_1354,N_916,N_933);
nor U1355 (N_1355,N_250,N_481);
or U1356 (N_1356,N_894,N_334);
and U1357 (N_1357,N_837,N_114);
xnor U1358 (N_1358,N_246,N_307);
or U1359 (N_1359,N_56,N_224);
nand U1360 (N_1360,N_846,N_605);
nor U1361 (N_1361,N_842,N_260);
or U1362 (N_1362,N_985,N_575);
nand U1363 (N_1363,N_523,N_81);
and U1364 (N_1364,N_735,N_265);
nor U1365 (N_1365,N_859,N_759);
nor U1366 (N_1366,N_806,N_218);
nor U1367 (N_1367,N_721,N_840);
nand U1368 (N_1368,N_568,N_711);
or U1369 (N_1369,N_179,N_919);
nor U1370 (N_1370,N_917,N_437);
nor U1371 (N_1371,N_572,N_752);
nand U1372 (N_1372,N_632,N_882);
or U1373 (N_1373,N_470,N_340);
nor U1374 (N_1374,N_181,N_444);
or U1375 (N_1375,N_593,N_257);
nor U1376 (N_1376,N_935,N_515);
and U1377 (N_1377,N_223,N_613);
and U1378 (N_1378,N_564,N_233);
or U1379 (N_1379,N_537,N_694);
or U1380 (N_1380,N_176,N_707);
nor U1381 (N_1381,N_297,N_286);
xnor U1382 (N_1382,N_577,N_73);
nand U1383 (N_1383,N_671,N_51);
and U1384 (N_1384,N_879,N_578);
nor U1385 (N_1385,N_930,N_433);
or U1386 (N_1386,N_668,N_201);
xor U1387 (N_1387,N_438,N_456);
or U1388 (N_1388,N_313,N_282);
or U1389 (N_1389,N_833,N_461);
and U1390 (N_1390,N_421,N_271);
nor U1391 (N_1391,N_687,N_405);
nor U1392 (N_1392,N_105,N_397);
nor U1393 (N_1393,N_845,N_451);
and U1394 (N_1394,N_780,N_839);
and U1395 (N_1395,N_391,N_811);
nor U1396 (N_1396,N_268,N_75);
and U1397 (N_1397,N_870,N_213);
nor U1398 (N_1398,N_570,N_983);
and U1399 (N_1399,N_93,N_502);
and U1400 (N_1400,N_366,N_685);
nor U1401 (N_1401,N_84,N_991);
nor U1402 (N_1402,N_331,N_480);
nand U1403 (N_1403,N_516,N_113);
or U1404 (N_1404,N_414,N_608);
nand U1405 (N_1405,N_28,N_300);
or U1406 (N_1406,N_976,N_167);
nand U1407 (N_1407,N_966,N_140);
nand U1408 (N_1408,N_626,N_850);
nand U1409 (N_1409,N_513,N_612);
nand U1410 (N_1410,N_61,N_184);
and U1411 (N_1411,N_736,N_998);
nor U1412 (N_1412,N_629,N_827);
and U1413 (N_1413,N_277,N_195);
nor U1414 (N_1414,N_327,N_353);
and U1415 (N_1415,N_545,N_454);
nor U1416 (N_1416,N_804,N_54);
nor U1417 (N_1417,N_965,N_59);
or U1418 (N_1418,N_824,N_853);
or U1419 (N_1419,N_831,N_5);
nor U1420 (N_1420,N_230,N_266);
nand U1421 (N_1421,N_382,N_207);
nor U1422 (N_1422,N_216,N_412);
nor U1423 (N_1423,N_761,N_332);
or U1424 (N_1424,N_65,N_662);
nor U1425 (N_1425,N_739,N_667);
nand U1426 (N_1426,N_354,N_162);
and U1427 (N_1427,N_409,N_900);
nand U1428 (N_1428,N_361,N_624);
and U1429 (N_1429,N_628,N_617);
nor U1430 (N_1430,N_80,N_583);
or U1431 (N_1431,N_350,N_263);
and U1432 (N_1432,N_491,N_339);
nor U1433 (N_1433,N_245,N_221);
nand U1434 (N_1434,N_357,N_293);
nor U1435 (N_1435,N_270,N_15);
nand U1436 (N_1436,N_296,N_924);
or U1437 (N_1437,N_345,N_597);
nand U1438 (N_1438,N_959,N_190);
nand U1439 (N_1439,N_326,N_581);
nand U1440 (N_1440,N_669,N_49);
nand U1441 (N_1441,N_486,N_479);
nand U1442 (N_1442,N_169,N_210);
nand U1443 (N_1443,N_657,N_592);
nor U1444 (N_1444,N_674,N_937);
or U1445 (N_1445,N_115,N_186);
nor U1446 (N_1446,N_50,N_308);
nor U1447 (N_1447,N_947,N_48);
or U1448 (N_1448,N_661,N_693);
and U1449 (N_1449,N_751,N_133);
or U1450 (N_1450,N_793,N_952);
nand U1451 (N_1451,N_571,N_445);
nor U1452 (N_1452,N_970,N_398);
nor U1453 (N_1453,N_849,N_552);
or U1454 (N_1454,N_135,N_189);
nor U1455 (N_1455,N_648,N_962);
nor U1456 (N_1456,N_298,N_941);
nor U1457 (N_1457,N_131,N_338);
or U1458 (N_1458,N_16,N_322);
or U1459 (N_1459,N_764,N_143);
nor U1460 (N_1460,N_74,N_803);
and U1461 (N_1461,N_773,N_862);
and U1462 (N_1462,N_330,N_465);
and U1463 (N_1463,N_107,N_558);
nor U1464 (N_1464,N_953,N_197);
or U1465 (N_1465,N_116,N_650);
or U1466 (N_1466,N_122,N_829);
nand U1467 (N_1467,N_784,N_874);
and U1468 (N_1468,N_852,N_996);
nand U1469 (N_1469,N_700,N_664);
and U1470 (N_1470,N_794,N_431);
nand U1471 (N_1471,N_101,N_912);
or U1472 (N_1472,N_556,N_713);
nor U1473 (N_1473,N_474,N_90);
nor U1474 (N_1474,N_394,N_91);
or U1475 (N_1475,N_722,N_159);
and U1476 (N_1476,N_446,N_175);
or U1477 (N_1477,N_987,N_770);
nor U1478 (N_1478,N_325,N_893);
and U1479 (N_1479,N_96,N_993);
nor U1480 (N_1480,N_460,N_890);
and U1481 (N_1481,N_6,N_312);
and U1482 (N_1482,N_746,N_473);
or U1483 (N_1483,N_964,N_686);
nand U1484 (N_1484,N_161,N_442);
nand U1485 (N_1485,N_7,N_757);
or U1486 (N_1486,N_415,N_259);
nand U1487 (N_1487,N_584,N_504);
nor U1488 (N_1488,N_511,N_112);
or U1489 (N_1489,N_262,N_123);
nor U1490 (N_1490,N_892,N_522);
nor U1491 (N_1491,N_574,N_781);
nor U1492 (N_1492,N_418,N_495);
nand U1493 (N_1493,N_623,N_776);
nor U1494 (N_1494,N_527,N_483);
nand U1495 (N_1495,N_464,N_566);
or U1496 (N_1496,N_212,N_36);
nor U1497 (N_1497,N_813,N_151);
nor U1498 (N_1498,N_400,N_989);
and U1499 (N_1499,N_635,N_290);
and U1500 (N_1500,N_10,N_448);
nor U1501 (N_1501,N_434,N_80);
and U1502 (N_1502,N_601,N_528);
or U1503 (N_1503,N_677,N_180);
nor U1504 (N_1504,N_522,N_112);
or U1505 (N_1505,N_320,N_335);
nand U1506 (N_1506,N_615,N_620);
nor U1507 (N_1507,N_160,N_668);
nor U1508 (N_1508,N_697,N_820);
or U1509 (N_1509,N_780,N_937);
or U1510 (N_1510,N_854,N_912);
nand U1511 (N_1511,N_438,N_419);
or U1512 (N_1512,N_415,N_8);
and U1513 (N_1513,N_257,N_458);
and U1514 (N_1514,N_14,N_665);
nand U1515 (N_1515,N_907,N_488);
or U1516 (N_1516,N_882,N_593);
nand U1517 (N_1517,N_595,N_631);
nand U1518 (N_1518,N_640,N_791);
or U1519 (N_1519,N_225,N_781);
or U1520 (N_1520,N_157,N_821);
or U1521 (N_1521,N_495,N_34);
and U1522 (N_1522,N_19,N_46);
nand U1523 (N_1523,N_15,N_368);
or U1524 (N_1524,N_92,N_857);
or U1525 (N_1525,N_222,N_529);
and U1526 (N_1526,N_851,N_536);
nor U1527 (N_1527,N_895,N_584);
nor U1528 (N_1528,N_858,N_482);
nor U1529 (N_1529,N_935,N_472);
or U1530 (N_1530,N_72,N_801);
nand U1531 (N_1531,N_414,N_82);
or U1532 (N_1532,N_500,N_51);
nor U1533 (N_1533,N_800,N_941);
and U1534 (N_1534,N_296,N_919);
and U1535 (N_1535,N_232,N_758);
nand U1536 (N_1536,N_877,N_102);
nor U1537 (N_1537,N_306,N_940);
and U1538 (N_1538,N_362,N_650);
nand U1539 (N_1539,N_406,N_576);
or U1540 (N_1540,N_210,N_460);
nand U1541 (N_1541,N_480,N_484);
nor U1542 (N_1542,N_595,N_223);
or U1543 (N_1543,N_192,N_352);
nand U1544 (N_1544,N_877,N_825);
and U1545 (N_1545,N_381,N_475);
nor U1546 (N_1546,N_627,N_621);
and U1547 (N_1547,N_375,N_656);
nand U1548 (N_1548,N_622,N_472);
nor U1549 (N_1549,N_101,N_753);
nor U1550 (N_1550,N_767,N_897);
nor U1551 (N_1551,N_382,N_232);
nor U1552 (N_1552,N_758,N_133);
nor U1553 (N_1553,N_472,N_909);
nand U1554 (N_1554,N_931,N_321);
and U1555 (N_1555,N_508,N_643);
and U1556 (N_1556,N_837,N_934);
or U1557 (N_1557,N_875,N_957);
and U1558 (N_1558,N_772,N_864);
or U1559 (N_1559,N_164,N_69);
nor U1560 (N_1560,N_299,N_714);
nor U1561 (N_1561,N_871,N_537);
nor U1562 (N_1562,N_876,N_448);
or U1563 (N_1563,N_479,N_104);
and U1564 (N_1564,N_489,N_494);
nor U1565 (N_1565,N_889,N_465);
or U1566 (N_1566,N_413,N_931);
nand U1567 (N_1567,N_522,N_435);
or U1568 (N_1568,N_739,N_330);
or U1569 (N_1569,N_60,N_87);
xor U1570 (N_1570,N_470,N_680);
xnor U1571 (N_1571,N_304,N_991);
and U1572 (N_1572,N_16,N_866);
nor U1573 (N_1573,N_182,N_668);
nand U1574 (N_1574,N_619,N_671);
xor U1575 (N_1575,N_966,N_70);
and U1576 (N_1576,N_991,N_676);
or U1577 (N_1577,N_578,N_737);
or U1578 (N_1578,N_628,N_399);
nor U1579 (N_1579,N_850,N_562);
nand U1580 (N_1580,N_134,N_657);
or U1581 (N_1581,N_66,N_659);
or U1582 (N_1582,N_605,N_766);
or U1583 (N_1583,N_792,N_798);
or U1584 (N_1584,N_808,N_999);
or U1585 (N_1585,N_241,N_505);
and U1586 (N_1586,N_498,N_799);
nor U1587 (N_1587,N_780,N_997);
or U1588 (N_1588,N_686,N_98);
and U1589 (N_1589,N_374,N_549);
and U1590 (N_1590,N_3,N_109);
xnor U1591 (N_1591,N_94,N_578);
nand U1592 (N_1592,N_531,N_987);
or U1593 (N_1593,N_155,N_851);
or U1594 (N_1594,N_47,N_552);
nor U1595 (N_1595,N_927,N_293);
nand U1596 (N_1596,N_521,N_198);
nand U1597 (N_1597,N_209,N_533);
nor U1598 (N_1598,N_141,N_936);
nor U1599 (N_1599,N_100,N_49);
or U1600 (N_1600,N_340,N_337);
and U1601 (N_1601,N_887,N_716);
and U1602 (N_1602,N_166,N_807);
nor U1603 (N_1603,N_120,N_911);
nand U1604 (N_1604,N_872,N_143);
xnor U1605 (N_1605,N_895,N_22);
or U1606 (N_1606,N_449,N_101);
or U1607 (N_1607,N_870,N_743);
nor U1608 (N_1608,N_515,N_606);
and U1609 (N_1609,N_432,N_370);
nand U1610 (N_1610,N_406,N_584);
nor U1611 (N_1611,N_320,N_814);
or U1612 (N_1612,N_581,N_221);
and U1613 (N_1613,N_420,N_349);
and U1614 (N_1614,N_545,N_381);
or U1615 (N_1615,N_432,N_504);
nor U1616 (N_1616,N_775,N_25);
and U1617 (N_1617,N_429,N_515);
nor U1618 (N_1618,N_658,N_200);
nand U1619 (N_1619,N_655,N_661);
and U1620 (N_1620,N_363,N_858);
nand U1621 (N_1621,N_4,N_459);
nand U1622 (N_1622,N_270,N_400);
or U1623 (N_1623,N_342,N_341);
nor U1624 (N_1624,N_21,N_23);
nor U1625 (N_1625,N_532,N_867);
or U1626 (N_1626,N_790,N_945);
and U1627 (N_1627,N_290,N_275);
nor U1628 (N_1628,N_104,N_958);
and U1629 (N_1629,N_652,N_193);
nand U1630 (N_1630,N_761,N_326);
or U1631 (N_1631,N_87,N_320);
and U1632 (N_1632,N_177,N_830);
nor U1633 (N_1633,N_889,N_753);
nand U1634 (N_1634,N_769,N_179);
nand U1635 (N_1635,N_582,N_776);
or U1636 (N_1636,N_385,N_420);
and U1637 (N_1637,N_182,N_278);
nor U1638 (N_1638,N_147,N_47);
nand U1639 (N_1639,N_64,N_161);
nand U1640 (N_1640,N_243,N_913);
or U1641 (N_1641,N_87,N_927);
and U1642 (N_1642,N_205,N_952);
nor U1643 (N_1643,N_443,N_25);
xor U1644 (N_1644,N_488,N_672);
and U1645 (N_1645,N_244,N_863);
nand U1646 (N_1646,N_492,N_422);
and U1647 (N_1647,N_375,N_696);
or U1648 (N_1648,N_637,N_47);
nand U1649 (N_1649,N_976,N_645);
and U1650 (N_1650,N_724,N_574);
and U1651 (N_1651,N_819,N_125);
and U1652 (N_1652,N_916,N_175);
and U1653 (N_1653,N_304,N_876);
or U1654 (N_1654,N_944,N_539);
nand U1655 (N_1655,N_918,N_496);
or U1656 (N_1656,N_294,N_289);
and U1657 (N_1657,N_898,N_643);
and U1658 (N_1658,N_91,N_557);
nor U1659 (N_1659,N_696,N_585);
and U1660 (N_1660,N_351,N_54);
xnor U1661 (N_1661,N_635,N_186);
nor U1662 (N_1662,N_214,N_18);
and U1663 (N_1663,N_59,N_107);
or U1664 (N_1664,N_83,N_930);
nor U1665 (N_1665,N_361,N_664);
nor U1666 (N_1666,N_563,N_266);
and U1667 (N_1667,N_218,N_430);
nand U1668 (N_1668,N_8,N_499);
and U1669 (N_1669,N_381,N_878);
or U1670 (N_1670,N_961,N_650);
nand U1671 (N_1671,N_524,N_648);
and U1672 (N_1672,N_151,N_436);
or U1673 (N_1673,N_903,N_946);
and U1674 (N_1674,N_168,N_432);
or U1675 (N_1675,N_288,N_394);
or U1676 (N_1676,N_601,N_914);
or U1677 (N_1677,N_709,N_883);
nor U1678 (N_1678,N_847,N_441);
nand U1679 (N_1679,N_364,N_665);
nand U1680 (N_1680,N_138,N_506);
and U1681 (N_1681,N_585,N_405);
nand U1682 (N_1682,N_250,N_526);
nand U1683 (N_1683,N_868,N_717);
and U1684 (N_1684,N_36,N_300);
and U1685 (N_1685,N_946,N_40);
nand U1686 (N_1686,N_747,N_78);
nand U1687 (N_1687,N_666,N_724);
or U1688 (N_1688,N_962,N_931);
and U1689 (N_1689,N_613,N_128);
and U1690 (N_1690,N_348,N_129);
and U1691 (N_1691,N_853,N_807);
nor U1692 (N_1692,N_672,N_891);
nand U1693 (N_1693,N_786,N_9);
and U1694 (N_1694,N_292,N_735);
or U1695 (N_1695,N_36,N_965);
and U1696 (N_1696,N_880,N_789);
nor U1697 (N_1697,N_570,N_184);
nor U1698 (N_1698,N_83,N_101);
nand U1699 (N_1699,N_546,N_533);
or U1700 (N_1700,N_479,N_294);
and U1701 (N_1701,N_261,N_686);
xor U1702 (N_1702,N_15,N_891);
and U1703 (N_1703,N_656,N_625);
and U1704 (N_1704,N_594,N_258);
or U1705 (N_1705,N_868,N_179);
nor U1706 (N_1706,N_661,N_901);
and U1707 (N_1707,N_846,N_635);
nor U1708 (N_1708,N_750,N_79);
nor U1709 (N_1709,N_58,N_857);
or U1710 (N_1710,N_458,N_577);
and U1711 (N_1711,N_752,N_608);
nor U1712 (N_1712,N_211,N_331);
or U1713 (N_1713,N_436,N_412);
nand U1714 (N_1714,N_49,N_292);
nand U1715 (N_1715,N_884,N_537);
nor U1716 (N_1716,N_119,N_601);
or U1717 (N_1717,N_450,N_687);
or U1718 (N_1718,N_70,N_850);
and U1719 (N_1719,N_149,N_40);
or U1720 (N_1720,N_128,N_847);
nor U1721 (N_1721,N_88,N_201);
and U1722 (N_1722,N_598,N_509);
or U1723 (N_1723,N_987,N_528);
nand U1724 (N_1724,N_99,N_763);
or U1725 (N_1725,N_631,N_484);
nand U1726 (N_1726,N_772,N_861);
nor U1727 (N_1727,N_908,N_214);
xnor U1728 (N_1728,N_252,N_375);
nor U1729 (N_1729,N_927,N_893);
nor U1730 (N_1730,N_996,N_125);
nor U1731 (N_1731,N_874,N_119);
and U1732 (N_1732,N_942,N_225);
nor U1733 (N_1733,N_297,N_537);
and U1734 (N_1734,N_843,N_641);
and U1735 (N_1735,N_255,N_442);
or U1736 (N_1736,N_58,N_890);
and U1737 (N_1737,N_954,N_161);
nand U1738 (N_1738,N_986,N_214);
nand U1739 (N_1739,N_463,N_24);
or U1740 (N_1740,N_757,N_176);
and U1741 (N_1741,N_983,N_366);
nand U1742 (N_1742,N_155,N_204);
xor U1743 (N_1743,N_386,N_815);
and U1744 (N_1744,N_32,N_856);
and U1745 (N_1745,N_848,N_893);
and U1746 (N_1746,N_33,N_52);
nand U1747 (N_1747,N_643,N_798);
nand U1748 (N_1748,N_619,N_121);
and U1749 (N_1749,N_258,N_616);
nand U1750 (N_1750,N_262,N_511);
nand U1751 (N_1751,N_138,N_883);
and U1752 (N_1752,N_165,N_854);
and U1753 (N_1753,N_361,N_548);
and U1754 (N_1754,N_577,N_190);
xor U1755 (N_1755,N_765,N_389);
and U1756 (N_1756,N_779,N_141);
or U1757 (N_1757,N_577,N_626);
and U1758 (N_1758,N_65,N_910);
nor U1759 (N_1759,N_968,N_326);
xnor U1760 (N_1760,N_131,N_467);
and U1761 (N_1761,N_349,N_168);
nand U1762 (N_1762,N_851,N_511);
or U1763 (N_1763,N_401,N_887);
nand U1764 (N_1764,N_584,N_633);
nor U1765 (N_1765,N_550,N_864);
nand U1766 (N_1766,N_410,N_735);
and U1767 (N_1767,N_737,N_747);
and U1768 (N_1768,N_600,N_303);
nand U1769 (N_1769,N_485,N_482);
nand U1770 (N_1770,N_76,N_622);
nand U1771 (N_1771,N_76,N_653);
nor U1772 (N_1772,N_216,N_971);
or U1773 (N_1773,N_282,N_908);
or U1774 (N_1774,N_651,N_755);
nor U1775 (N_1775,N_826,N_834);
nor U1776 (N_1776,N_102,N_905);
or U1777 (N_1777,N_785,N_736);
and U1778 (N_1778,N_493,N_881);
and U1779 (N_1779,N_727,N_884);
or U1780 (N_1780,N_576,N_743);
and U1781 (N_1781,N_775,N_201);
and U1782 (N_1782,N_672,N_731);
nor U1783 (N_1783,N_835,N_941);
nand U1784 (N_1784,N_461,N_390);
nor U1785 (N_1785,N_343,N_366);
nor U1786 (N_1786,N_489,N_533);
or U1787 (N_1787,N_40,N_654);
and U1788 (N_1788,N_26,N_432);
nor U1789 (N_1789,N_349,N_553);
and U1790 (N_1790,N_20,N_803);
or U1791 (N_1791,N_353,N_206);
nor U1792 (N_1792,N_348,N_220);
and U1793 (N_1793,N_701,N_254);
and U1794 (N_1794,N_243,N_99);
nand U1795 (N_1795,N_97,N_67);
or U1796 (N_1796,N_177,N_163);
nor U1797 (N_1797,N_424,N_678);
nor U1798 (N_1798,N_464,N_237);
or U1799 (N_1799,N_771,N_652);
or U1800 (N_1800,N_769,N_271);
and U1801 (N_1801,N_323,N_299);
nor U1802 (N_1802,N_141,N_533);
nand U1803 (N_1803,N_946,N_526);
nand U1804 (N_1804,N_996,N_179);
and U1805 (N_1805,N_551,N_257);
and U1806 (N_1806,N_958,N_395);
and U1807 (N_1807,N_146,N_221);
or U1808 (N_1808,N_642,N_997);
or U1809 (N_1809,N_790,N_704);
or U1810 (N_1810,N_729,N_495);
xor U1811 (N_1811,N_744,N_36);
xnor U1812 (N_1812,N_180,N_235);
and U1813 (N_1813,N_259,N_178);
nor U1814 (N_1814,N_1,N_562);
nand U1815 (N_1815,N_70,N_410);
nor U1816 (N_1816,N_205,N_354);
nand U1817 (N_1817,N_460,N_379);
or U1818 (N_1818,N_135,N_164);
nand U1819 (N_1819,N_492,N_141);
or U1820 (N_1820,N_646,N_252);
and U1821 (N_1821,N_489,N_313);
or U1822 (N_1822,N_35,N_620);
nor U1823 (N_1823,N_474,N_920);
and U1824 (N_1824,N_947,N_554);
or U1825 (N_1825,N_333,N_863);
nor U1826 (N_1826,N_169,N_369);
nand U1827 (N_1827,N_239,N_804);
nor U1828 (N_1828,N_629,N_870);
nand U1829 (N_1829,N_421,N_967);
nand U1830 (N_1830,N_459,N_25);
nand U1831 (N_1831,N_422,N_281);
or U1832 (N_1832,N_300,N_849);
nand U1833 (N_1833,N_352,N_537);
nor U1834 (N_1834,N_433,N_585);
and U1835 (N_1835,N_647,N_953);
or U1836 (N_1836,N_158,N_359);
nand U1837 (N_1837,N_544,N_161);
or U1838 (N_1838,N_956,N_564);
nor U1839 (N_1839,N_408,N_195);
nand U1840 (N_1840,N_112,N_920);
nor U1841 (N_1841,N_265,N_839);
nand U1842 (N_1842,N_387,N_424);
and U1843 (N_1843,N_575,N_126);
nor U1844 (N_1844,N_493,N_36);
or U1845 (N_1845,N_915,N_884);
or U1846 (N_1846,N_800,N_300);
or U1847 (N_1847,N_764,N_754);
or U1848 (N_1848,N_342,N_854);
or U1849 (N_1849,N_547,N_437);
or U1850 (N_1850,N_661,N_375);
or U1851 (N_1851,N_58,N_246);
nor U1852 (N_1852,N_580,N_524);
and U1853 (N_1853,N_471,N_264);
nand U1854 (N_1854,N_194,N_233);
and U1855 (N_1855,N_895,N_311);
nand U1856 (N_1856,N_800,N_239);
nand U1857 (N_1857,N_257,N_309);
nor U1858 (N_1858,N_924,N_590);
nand U1859 (N_1859,N_337,N_459);
nor U1860 (N_1860,N_265,N_58);
and U1861 (N_1861,N_628,N_536);
xor U1862 (N_1862,N_89,N_47);
nand U1863 (N_1863,N_852,N_65);
nor U1864 (N_1864,N_235,N_590);
nand U1865 (N_1865,N_96,N_450);
nor U1866 (N_1866,N_142,N_402);
xor U1867 (N_1867,N_442,N_968);
nand U1868 (N_1868,N_119,N_561);
nor U1869 (N_1869,N_743,N_868);
or U1870 (N_1870,N_663,N_897);
or U1871 (N_1871,N_100,N_951);
or U1872 (N_1872,N_496,N_218);
nand U1873 (N_1873,N_61,N_299);
nand U1874 (N_1874,N_307,N_369);
or U1875 (N_1875,N_131,N_984);
and U1876 (N_1876,N_607,N_182);
or U1877 (N_1877,N_597,N_94);
nand U1878 (N_1878,N_944,N_845);
nor U1879 (N_1879,N_750,N_690);
nor U1880 (N_1880,N_325,N_823);
nor U1881 (N_1881,N_393,N_54);
and U1882 (N_1882,N_706,N_605);
or U1883 (N_1883,N_258,N_254);
and U1884 (N_1884,N_691,N_426);
nor U1885 (N_1885,N_435,N_379);
or U1886 (N_1886,N_450,N_72);
nand U1887 (N_1887,N_224,N_289);
nor U1888 (N_1888,N_306,N_729);
and U1889 (N_1889,N_656,N_391);
and U1890 (N_1890,N_586,N_622);
nand U1891 (N_1891,N_998,N_787);
nand U1892 (N_1892,N_956,N_886);
nor U1893 (N_1893,N_262,N_291);
nand U1894 (N_1894,N_875,N_765);
nor U1895 (N_1895,N_357,N_444);
and U1896 (N_1896,N_996,N_43);
nor U1897 (N_1897,N_205,N_363);
nor U1898 (N_1898,N_261,N_645);
nor U1899 (N_1899,N_831,N_573);
nor U1900 (N_1900,N_383,N_287);
nor U1901 (N_1901,N_501,N_83);
nand U1902 (N_1902,N_547,N_285);
nor U1903 (N_1903,N_746,N_784);
or U1904 (N_1904,N_829,N_176);
or U1905 (N_1905,N_830,N_829);
nor U1906 (N_1906,N_825,N_56);
nand U1907 (N_1907,N_844,N_432);
nand U1908 (N_1908,N_859,N_192);
or U1909 (N_1909,N_71,N_968);
nand U1910 (N_1910,N_664,N_847);
and U1911 (N_1911,N_472,N_845);
nor U1912 (N_1912,N_927,N_453);
xnor U1913 (N_1913,N_999,N_102);
and U1914 (N_1914,N_370,N_179);
and U1915 (N_1915,N_287,N_43);
and U1916 (N_1916,N_447,N_408);
and U1917 (N_1917,N_673,N_932);
or U1918 (N_1918,N_844,N_715);
and U1919 (N_1919,N_25,N_227);
and U1920 (N_1920,N_805,N_65);
nand U1921 (N_1921,N_966,N_222);
nand U1922 (N_1922,N_397,N_534);
nor U1923 (N_1923,N_840,N_134);
or U1924 (N_1924,N_192,N_697);
and U1925 (N_1925,N_90,N_673);
nor U1926 (N_1926,N_477,N_603);
and U1927 (N_1927,N_572,N_366);
nor U1928 (N_1928,N_821,N_488);
or U1929 (N_1929,N_667,N_943);
and U1930 (N_1930,N_695,N_529);
or U1931 (N_1931,N_675,N_789);
nand U1932 (N_1932,N_332,N_359);
and U1933 (N_1933,N_264,N_812);
or U1934 (N_1934,N_945,N_129);
nor U1935 (N_1935,N_90,N_611);
and U1936 (N_1936,N_393,N_81);
or U1937 (N_1937,N_819,N_278);
nand U1938 (N_1938,N_174,N_151);
nor U1939 (N_1939,N_819,N_760);
or U1940 (N_1940,N_360,N_239);
and U1941 (N_1941,N_492,N_624);
nor U1942 (N_1942,N_757,N_604);
or U1943 (N_1943,N_867,N_205);
nor U1944 (N_1944,N_163,N_739);
nand U1945 (N_1945,N_370,N_630);
nor U1946 (N_1946,N_991,N_162);
and U1947 (N_1947,N_724,N_937);
nand U1948 (N_1948,N_102,N_531);
nand U1949 (N_1949,N_857,N_621);
and U1950 (N_1950,N_877,N_808);
nor U1951 (N_1951,N_153,N_608);
nor U1952 (N_1952,N_795,N_844);
nor U1953 (N_1953,N_137,N_613);
or U1954 (N_1954,N_638,N_483);
nor U1955 (N_1955,N_612,N_478);
xnor U1956 (N_1956,N_304,N_394);
or U1957 (N_1957,N_442,N_790);
nand U1958 (N_1958,N_657,N_14);
or U1959 (N_1959,N_202,N_581);
nand U1960 (N_1960,N_40,N_333);
or U1961 (N_1961,N_711,N_363);
nor U1962 (N_1962,N_202,N_679);
or U1963 (N_1963,N_307,N_393);
and U1964 (N_1964,N_810,N_405);
or U1965 (N_1965,N_435,N_705);
or U1966 (N_1966,N_260,N_46);
nand U1967 (N_1967,N_811,N_856);
and U1968 (N_1968,N_703,N_680);
or U1969 (N_1969,N_859,N_57);
nand U1970 (N_1970,N_998,N_144);
nand U1971 (N_1971,N_703,N_563);
nand U1972 (N_1972,N_387,N_340);
nand U1973 (N_1973,N_64,N_84);
or U1974 (N_1974,N_72,N_629);
nor U1975 (N_1975,N_371,N_455);
nor U1976 (N_1976,N_449,N_890);
and U1977 (N_1977,N_353,N_380);
nor U1978 (N_1978,N_499,N_236);
or U1979 (N_1979,N_910,N_25);
nor U1980 (N_1980,N_244,N_927);
and U1981 (N_1981,N_102,N_529);
nand U1982 (N_1982,N_608,N_764);
nand U1983 (N_1983,N_110,N_960);
and U1984 (N_1984,N_275,N_994);
nand U1985 (N_1985,N_353,N_167);
nand U1986 (N_1986,N_971,N_744);
nand U1987 (N_1987,N_425,N_473);
or U1988 (N_1988,N_745,N_110);
nand U1989 (N_1989,N_843,N_32);
and U1990 (N_1990,N_915,N_421);
nor U1991 (N_1991,N_467,N_224);
nand U1992 (N_1992,N_900,N_18);
xnor U1993 (N_1993,N_309,N_955);
xnor U1994 (N_1994,N_46,N_585);
and U1995 (N_1995,N_739,N_581);
and U1996 (N_1996,N_734,N_640);
nand U1997 (N_1997,N_257,N_160);
nor U1998 (N_1998,N_916,N_531);
nor U1999 (N_1999,N_425,N_616);
and U2000 (N_2000,N_1151,N_1262);
nand U2001 (N_2001,N_1423,N_1464);
and U2002 (N_2002,N_1128,N_1880);
nand U2003 (N_2003,N_1341,N_1312);
nand U2004 (N_2004,N_1411,N_1957);
or U2005 (N_2005,N_1360,N_1031);
nand U2006 (N_2006,N_1167,N_1217);
or U2007 (N_2007,N_1791,N_1119);
nand U2008 (N_2008,N_1886,N_1304);
or U2009 (N_2009,N_1123,N_1111);
nand U2010 (N_2010,N_1853,N_1436);
and U2011 (N_2011,N_1546,N_1776);
nand U2012 (N_2012,N_1327,N_1744);
or U2013 (N_2013,N_1460,N_1682);
nand U2014 (N_2014,N_1252,N_1442);
nor U2015 (N_2015,N_1389,N_1543);
xor U2016 (N_2016,N_1889,N_1752);
and U2017 (N_2017,N_1154,N_1909);
nand U2018 (N_2018,N_1887,N_1751);
nand U2019 (N_2019,N_1103,N_1396);
or U2020 (N_2020,N_1882,N_1748);
nor U2021 (N_2021,N_1308,N_1617);
nor U2022 (N_2022,N_1350,N_1141);
and U2023 (N_2023,N_1471,N_1246);
nor U2024 (N_2024,N_1796,N_1004);
nand U2025 (N_2025,N_1229,N_1047);
nor U2026 (N_2026,N_1306,N_1615);
nor U2027 (N_2027,N_1062,N_1156);
nor U2028 (N_2028,N_1370,N_1509);
nand U2029 (N_2029,N_1907,N_1122);
nand U2030 (N_2030,N_1575,N_1714);
and U2031 (N_2031,N_1646,N_1079);
or U2032 (N_2032,N_1879,N_1037);
nand U2033 (N_2033,N_1032,N_1679);
and U2034 (N_2034,N_1121,N_1535);
nor U2035 (N_2035,N_1651,N_1457);
and U2036 (N_2036,N_1588,N_1768);
and U2037 (N_2037,N_1799,N_1200);
and U2038 (N_2038,N_1949,N_1135);
nor U2039 (N_2039,N_1481,N_1434);
or U2040 (N_2040,N_1400,N_1338);
or U2041 (N_2041,N_1024,N_1598);
nor U2042 (N_2042,N_1560,N_1028);
and U2043 (N_2043,N_1921,N_1737);
and U2044 (N_2044,N_1764,N_1956);
nor U2045 (N_2045,N_1629,N_1142);
and U2046 (N_2046,N_1426,N_1541);
and U2047 (N_2047,N_1124,N_1280);
nand U2048 (N_2048,N_1727,N_1045);
or U2049 (N_2049,N_1057,N_1131);
and U2050 (N_2050,N_1666,N_1248);
and U2051 (N_2051,N_1740,N_1494);
and U2052 (N_2052,N_1511,N_1240);
nor U2053 (N_2053,N_1066,N_1641);
or U2054 (N_2054,N_1258,N_1050);
nand U2055 (N_2055,N_1186,N_1081);
nand U2056 (N_2056,N_1166,N_1561);
or U2057 (N_2057,N_1673,N_1149);
nor U2058 (N_2058,N_1709,N_1242);
or U2059 (N_2059,N_1499,N_1275);
and U2060 (N_2060,N_1928,N_1427);
xor U2061 (N_2061,N_1516,N_1273);
nand U2062 (N_2062,N_1798,N_1146);
nor U2063 (N_2063,N_1595,N_1540);
and U2064 (N_2064,N_1072,N_1284);
nand U2065 (N_2065,N_1997,N_1754);
and U2066 (N_2066,N_1580,N_1602);
and U2067 (N_2067,N_1319,N_1894);
or U2068 (N_2068,N_1194,N_1895);
nand U2069 (N_2069,N_1048,N_1683);
or U2070 (N_2070,N_1844,N_1552);
or U2071 (N_2071,N_1946,N_1728);
and U2072 (N_2072,N_1850,N_1948);
nand U2073 (N_2073,N_1725,N_1906);
and U2074 (N_2074,N_1136,N_1969);
nand U2075 (N_2075,N_1971,N_1388);
nand U2076 (N_2076,N_1323,N_1978);
and U2077 (N_2077,N_1896,N_1099);
nor U2078 (N_2078,N_1385,N_1571);
nor U2079 (N_2079,N_1624,N_1719);
nor U2080 (N_2080,N_1623,N_1745);
or U2081 (N_2081,N_1771,N_1954);
and U2082 (N_2082,N_1467,N_1923);
or U2083 (N_2083,N_1660,N_1721);
nand U2084 (N_2084,N_1581,N_1374);
nor U2085 (N_2085,N_1981,N_1170);
and U2086 (N_2086,N_1572,N_1036);
nand U2087 (N_2087,N_1030,N_1184);
xor U2088 (N_2088,N_1443,N_1428);
nand U2089 (N_2089,N_1658,N_1608);
nand U2090 (N_2090,N_1074,N_1147);
xnor U2091 (N_2091,N_1309,N_1840);
or U2092 (N_2092,N_1049,N_1318);
nor U2093 (N_2093,N_1778,N_1414);
nor U2094 (N_2094,N_1846,N_1484);
nor U2095 (N_2095,N_1455,N_1401);
nand U2096 (N_2096,N_1181,N_1349);
and U2097 (N_2097,N_1579,N_1652);
and U2098 (N_2098,N_1817,N_1266);
nand U2099 (N_2099,N_1253,N_1953);
and U2100 (N_2100,N_1902,N_1645);
nand U2101 (N_2101,N_1684,N_1854);
or U2102 (N_2102,N_1230,N_1508);
or U2103 (N_2103,N_1178,N_1755);
and U2104 (N_2104,N_1819,N_1209);
and U2105 (N_2105,N_1247,N_1218);
nand U2106 (N_2106,N_1769,N_1500);
or U2107 (N_2107,N_1664,N_1775);
and U2108 (N_2108,N_1991,N_1298);
nand U2109 (N_2109,N_1493,N_1314);
nand U2110 (N_2110,N_1576,N_1734);
nand U2111 (N_2111,N_1227,N_1591);
or U2112 (N_2112,N_1093,N_1279);
nor U2113 (N_2113,N_1449,N_1931);
or U2114 (N_2114,N_1251,N_1593);
nand U2115 (N_2115,N_1100,N_1597);
and U2116 (N_2116,N_1925,N_1980);
nand U2117 (N_2117,N_1067,N_1017);
or U2118 (N_2118,N_1342,N_1568);
nand U2119 (N_2119,N_1272,N_1694);
nor U2120 (N_2120,N_1935,N_1526);
or U2121 (N_2121,N_1618,N_1406);
xnor U2122 (N_2122,N_1559,N_1006);
and U2123 (N_2123,N_1000,N_1988);
nand U2124 (N_2124,N_1270,N_1678);
nor U2125 (N_2125,N_1225,N_1089);
nand U2126 (N_2126,N_1422,N_1452);
nor U2127 (N_2127,N_1235,N_1310);
nand U2128 (N_2128,N_1289,N_1205);
or U2129 (N_2129,N_1912,N_1107);
xnor U2130 (N_2130,N_1356,N_1334);
and U2131 (N_2131,N_1808,N_1655);
or U2132 (N_2132,N_1930,N_1013);
and U2133 (N_2133,N_1998,N_1905);
nand U2134 (N_2134,N_1269,N_1790);
nand U2135 (N_2135,N_1398,N_1491);
nor U2136 (N_2136,N_1291,N_1842);
nor U2137 (N_2137,N_1035,N_1650);
nand U2138 (N_2138,N_1403,N_1478);
nand U2139 (N_2139,N_1736,N_1685);
xnor U2140 (N_2140,N_1897,N_1346);
xor U2141 (N_2141,N_1361,N_1090);
and U2142 (N_2142,N_1920,N_1022);
or U2143 (N_2143,N_1976,N_1465);
nand U2144 (N_2144,N_1249,N_1340);
and U2145 (N_2145,N_1900,N_1566);
or U2146 (N_2146,N_1451,N_1355);
nand U2147 (N_2147,N_1809,N_1753);
nand U2148 (N_2148,N_1105,N_1102);
xor U2149 (N_2149,N_1375,N_1758);
nand U2150 (N_2150,N_1885,N_1545);
and U2151 (N_2151,N_1332,N_1760);
or U2152 (N_2152,N_1497,N_1005);
and U2153 (N_2153,N_1155,N_1109);
and U2154 (N_2154,N_1926,N_1250);
or U2155 (N_2155,N_1870,N_1807);
nand U2156 (N_2156,N_1795,N_1527);
and U2157 (N_2157,N_1642,N_1640);
and U2158 (N_2158,N_1762,N_1033);
or U2159 (N_2159,N_1717,N_1199);
or U2160 (N_2160,N_1787,N_1483);
or U2161 (N_2161,N_1667,N_1945);
and U2162 (N_2162,N_1805,N_1486);
and U2163 (N_2163,N_1430,N_1616);
or U2164 (N_2164,N_1958,N_1419);
and U2165 (N_2165,N_1607,N_1255);
or U2166 (N_2166,N_1773,N_1782);
or U2167 (N_2167,N_1772,N_1357);
and U2168 (N_2168,N_1082,N_1404);
and U2169 (N_2169,N_1635,N_1992);
or U2170 (N_2170,N_1139,N_1722);
and U2171 (N_2171,N_1127,N_1183);
nand U2172 (N_2172,N_1029,N_1365);
nor U2173 (N_2173,N_1814,N_1697);
and U2174 (N_2174,N_1282,N_1890);
and U2175 (N_2175,N_1120,N_1162);
nand U2176 (N_2176,N_1116,N_1631);
nor U2177 (N_2177,N_1838,N_1822);
and U2178 (N_2178,N_1061,N_1522);
nor U2179 (N_2179,N_1055,N_1399);
or U2180 (N_2180,N_1379,N_1784);
or U2181 (N_2181,N_1803,N_1381);
and U2182 (N_2182,N_1321,N_1779);
nor U2183 (N_2183,N_1816,N_1830);
or U2184 (N_2184,N_1704,N_1876);
or U2185 (N_2185,N_1437,N_1010);
nand U2186 (N_2186,N_1831,N_1354);
or U2187 (N_2187,N_1636,N_1690);
nor U2188 (N_2188,N_1197,N_1416);
or U2189 (N_2189,N_1176,N_1852);
and U2190 (N_2190,N_1910,N_1950);
nand U2191 (N_2191,N_1555,N_1833);
and U2192 (N_2192,N_1777,N_1695);
nor U2193 (N_2193,N_1573,N_1182);
nor U2194 (N_2194,N_1832,N_1532);
nand U2195 (N_2195,N_1390,N_1649);
nor U2196 (N_2196,N_1968,N_1875);
and U2197 (N_2197,N_1490,N_1175);
nor U2198 (N_2198,N_1421,N_1440);
nand U2199 (N_2199,N_1080,N_1007);
xnor U2200 (N_2200,N_1157,N_1610);
nand U2201 (N_2201,N_1513,N_1707);
or U2202 (N_2202,N_1330,N_1256);
or U2203 (N_2203,N_1731,N_1461);
and U2204 (N_2204,N_1908,N_1232);
xnor U2205 (N_2205,N_1418,N_1820);
and U2206 (N_2206,N_1628,N_1553);
nor U2207 (N_2207,N_1883,N_1094);
nand U2208 (N_2208,N_1002,N_1533);
xnor U2209 (N_2209,N_1244,N_1405);
or U2210 (N_2210,N_1936,N_1689);
and U2211 (N_2211,N_1158,N_1039);
and U2212 (N_2212,N_1963,N_1989);
nand U2213 (N_2213,N_1480,N_1322);
xor U2214 (N_2214,N_1397,N_1387);
nand U2215 (N_2215,N_1245,N_1632);
nor U2216 (N_2216,N_1821,N_1104);
or U2217 (N_2217,N_1520,N_1849);
and U2218 (N_2218,N_1380,N_1671);
or U2219 (N_2219,N_1215,N_1008);
or U2220 (N_2220,N_1172,N_1362);
or U2221 (N_2221,N_1085,N_1818);
nor U2222 (N_2222,N_1841,N_1300);
xor U2223 (N_2223,N_1425,N_1196);
nand U2224 (N_2224,N_1320,N_1564);
or U2225 (N_2225,N_1653,N_1877);
and U2226 (N_2226,N_1961,N_1868);
nor U2227 (N_2227,N_1274,N_1661);
nand U2228 (N_2228,N_1797,N_1363);
and U2229 (N_2229,N_1382,N_1899);
nor U2230 (N_2230,N_1892,N_1523);
and U2231 (N_2231,N_1058,N_1019);
nor U2232 (N_2232,N_1324,N_1095);
and U2233 (N_2233,N_1222,N_1625);
nor U2234 (N_2234,N_1757,N_1974);
or U2235 (N_2235,N_1829,N_1469);
nor U2236 (N_2236,N_1506,N_1474);
nor U2237 (N_2237,N_1743,N_1839);
or U2238 (N_2238,N_1530,N_1501);
or U2239 (N_2239,N_1496,N_1171);
or U2240 (N_2240,N_1582,N_1348);
and U2241 (N_2241,N_1152,N_1177);
nand U2242 (N_2242,N_1088,N_1410);
and U2243 (N_2243,N_1164,N_1488);
or U2244 (N_2244,N_1701,N_1601);
or U2245 (N_2245,N_1145,N_1932);
nand U2246 (N_2246,N_1479,N_1210);
nor U2247 (N_2247,N_1054,N_1051);
nor U2248 (N_2248,N_1525,N_1993);
nand U2249 (N_2249,N_1789,N_1687);
or U2250 (N_2250,N_1187,N_1703);
nand U2251 (N_2251,N_1518,N_1710);
and U2252 (N_2252,N_1943,N_1848);
or U2253 (N_2253,N_1369,N_1009);
or U2254 (N_2254,N_1583,N_1173);
and U2255 (N_2255,N_1016,N_1806);
nor U2256 (N_2256,N_1216,N_1444);
nor U2257 (N_2257,N_1189,N_1940);
or U2258 (N_2258,N_1115,N_1371);
nand U2259 (N_2259,N_1763,N_1871);
and U2260 (N_2260,N_1160,N_1878);
and U2261 (N_2261,N_1929,N_1294);
or U2262 (N_2262,N_1825,N_1512);
or U2263 (N_2263,N_1335,N_1718);
and U2264 (N_2264,N_1433,N_1148);
and U2265 (N_2265,N_1134,N_1015);
nor U2266 (N_2266,N_1391,N_1698);
nand U2267 (N_2267,N_1857,N_1383);
and U2268 (N_2268,N_1515,N_1605);
nand U2269 (N_2269,N_1505,N_1236);
or U2270 (N_2270,N_1872,N_1358);
nand U2271 (N_2271,N_1691,N_1578);
nor U2272 (N_2272,N_1053,N_1263);
nand U2273 (N_2273,N_1344,N_1407);
nand U2274 (N_2274,N_1287,N_1693);
nand U2275 (N_2275,N_1549,N_1804);
nand U2276 (N_2276,N_1786,N_1688);
or U2277 (N_2277,N_1634,N_1783);
nand U2278 (N_2278,N_1705,N_1092);
or U2279 (N_2279,N_1677,N_1656);
or U2280 (N_2280,N_1001,N_1059);
and U2281 (N_2281,N_1959,N_1860);
and U2282 (N_2282,N_1609,N_1027);
or U2283 (N_2283,N_1378,N_1137);
or U2284 (N_2284,N_1668,N_1307);
or U2285 (N_2285,N_1285,N_1219);
nand U2286 (N_2286,N_1223,N_1812);
nand U2287 (N_2287,N_1845,N_1101);
nor U2288 (N_2288,N_1238,N_1723);
nand U2289 (N_2289,N_1746,N_1241);
nor U2290 (N_2290,N_1475,N_1811);
or U2291 (N_2291,N_1408,N_1052);
nor U2292 (N_2292,N_1918,N_1524);
and U2293 (N_2293,N_1861,N_1952);
nor U2294 (N_2294,N_1973,N_1233);
nand U2295 (N_2295,N_1563,N_1977);
and U2296 (N_2296,N_1014,N_1916);
nand U2297 (N_2297,N_1586,N_1622);
or U2298 (N_2298,N_1585,N_1901);
nor U2299 (N_2299,N_1767,N_1303);
and U2300 (N_2300,N_1316,N_1828);
nand U2301 (N_2301,N_1738,N_1866);
and U2302 (N_2302,N_1662,N_1402);
nor U2303 (N_2303,N_1299,N_1392);
xnor U2304 (N_2304,N_1445,N_1198);
nor U2305 (N_2305,N_1364,N_1788);
nand U2306 (N_2306,N_1712,N_1025);
nand U2307 (N_2307,N_1489,N_1268);
and U2308 (N_2308,N_1510,N_1732);
nor U2309 (N_2309,N_1603,N_1700);
or U2310 (N_2310,N_1325,N_1960);
nor U2311 (N_2311,N_1587,N_1277);
nand U2312 (N_2312,N_1858,N_1888);
nor U2313 (N_2313,N_1647,N_1826);
or U2314 (N_2314,N_1112,N_1020);
or U2315 (N_2315,N_1458,N_1810);
and U2316 (N_2316,N_1078,N_1542);
nor U2317 (N_2317,N_1937,N_1212);
nand U2318 (N_2318,N_1669,N_1503);
and U2319 (N_2319,N_1359,N_1292);
and U2320 (N_2320,N_1794,N_1823);
and U2321 (N_2321,N_1118,N_1163);
xnor U2322 (N_2322,N_1999,N_1130);
or U2323 (N_2323,N_1420,N_1011);
and U2324 (N_2324,N_1729,N_1295);
nor U2325 (N_2325,N_1681,N_1781);
nand U2326 (N_2326,N_1686,N_1550);
nor U2327 (N_2327,N_1674,N_1132);
or U2328 (N_2328,N_1023,N_1915);
nand U2329 (N_2329,N_1529,N_1495);
and U2330 (N_2330,N_1676,N_1947);
or U2331 (N_2331,N_1528,N_1975);
or U2332 (N_2332,N_1620,N_1800);
or U2333 (N_2333,N_1613,N_1046);
nand U2334 (N_2334,N_1574,N_1409);
nand U2335 (N_2335,N_1126,N_1672);
or U2336 (N_2336,N_1502,N_1836);
and U2337 (N_2337,N_1627,N_1352);
and U2338 (N_2338,N_1942,N_1188);
or U2339 (N_2339,N_1429,N_1435);
or U2340 (N_2340,N_1290,N_1565);
nand U2341 (N_2341,N_1174,N_1113);
or U2342 (N_2342,N_1333,N_1534);
nor U2343 (N_2343,N_1326,N_1551);
nor U2344 (N_2344,N_1243,N_1264);
nor U2345 (N_2345,N_1477,N_1168);
or U2346 (N_2346,N_1539,N_1463);
and U2347 (N_2347,N_1995,N_1473);
nor U2348 (N_2348,N_1075,N_1278);
nor U2349 (N_2349,N_1125,N_1468);
nand U2350 (N_2350,N_1498,N_1675);
or U2351 (N_2351,N_1336,N_1133);
nor U2352 (N_2352,N_1231,N_1372);
or U2353 (N_2353,N_1296,N_1742);
and U2354 (N_2354,N_1611,N_1874);
and U2355 (N_2355,N_1547,N_1454);
nor U2356 (N_2356,N_1206,N_1544);
or U2357 (N_2357,N_1612,N_1366);
and U2358 (N_2358,N_1643,N_1076);
or U2359 (N_2359,N_1856,N_1485);
or U2360 (N_2360,N_1064,N_1161);
or U2361 (N_2361,N_1190,N_1234);
xor U2362 (N_2362,N_1070,N_1413);
or U2363 (N_2363,N_1276,N_1557);
or U2364 (N_2364,N_1815,N_1487);
and U2365 (N_2365,N_1305,N_1042);
nand U2366 (N_2366,N_1087,N_1110);
or U2367 (N_2367,N_1570,N_1599);
and U2368 (N_2368,N_1747,N_1670);
or U2369 (N_2369,N_1680,N_1985);
and U2370 (N_2370,N_1211,N_1548);
and U2371 (N_2371,N_1281,N_1898);
nor U2372 (N_2372,N_1117,N_1749);
and U2373 (N_2373,N_1556,N_1891);
or U2374 (N_2374,N_1893,N_1780);
and U2375 (N_2375,N_1692,N_1302);
nand U2376 (N_2376,N_1637,N_1741);
or U2377 (N_2377,N_1944,N_1267);
nor U2378 (N_2378,N_1699,N_1271);
or U2379 (N_2379,N_1084,N_1453);
nor U2380 (N_2380,N_1012,N_1884);
nand U2381 (N_2381,N_1470,N_1766);
or U2382 (N_2382,N_1328,N_1143);
or U2383 (N_2383,N_1432,N_1914);
and U2384 (N_2384,N_1792,N_1091);
nand U2385 (N_2385,N_1201,N_1716);
or U2386 (N_2386,N_1855,N_1619);
nand U2387 (N_2387,N_1043,N_1638);
nand U2388 (N_2388,N_1696,N_1204);
and U2389 (N_2389,N_1129,N_1260);
nand U2390 (N_2390,N_1447,N_1114);
and U2391 (N_2391,N_1873,N_1865);
and U2392 (N_2392,N_1606,N_1140);
nand U2393 (N_2393,N_1073,N_1034);
and U2394 (N_2394,N_1600,N_1904);
and U2395 (N_2395,N_1317,N_1180);
nand U2396 (N_2396,N_1862,N_1538);
and U2397 (N_2397,N_1824,N_1730);
and U2398 (N_2398,N_1195,N_1715);
and U2399 (N_2399,N_1519,N_1867);
or U2400 (N_2400,N_1972,N_1395);
and U2401 (N_2401,N_1859,N_1086);
and U2402 (N_2402,N_1733,N_1724);
and U2403 (N_2403,N_1964,N_1922);
nand U2404 (N_2404,N_1351,N_1759);
or U2405 (N_2405,N_1329,N_1739);
nor U2406 (N_2406,N_1951,N_1237);
nor U2407 (N_2407,N_1265,N_1827);
nand U2408 (N_2408,N_1663,N_1462);
and U2409 (N_2409,N_1517,N_1060);
nor U2410 (N_2410,N_1417,N_1630);
and U2411 (N_2411,N_1596,N_1626);
and U2412 (N_2412,N_1331,N_1415);
nand U2413 (N_2413,N_1315,N_1514);
or U2414 (N_2414,N_1106,N_1228);
and U2415 (N_2415,N_1644,N_1569);
or U2416 (N_2416,N_1590,N_1881);
nor U2417 (N_2417,N_1504,N_1970);
or U2418 (N_2418,N_1982,N_1621);
or U2419 (N_2419,N_1214,N_1917);
nor U2420 (N_2420,N_1239,N_1531);
or U2421 (N_2421,N_1720,N_1903);
and U2422 (N_2422,N_1735,N_1301);
or U2423 (N_2423,N_1311,N_1785);
or U2424 (N_2424,N_1208,N_1224);
nand U2425 (N_2425,N_1837,N_1144);
nor U2426 (N_2426,N_1774,N_1040);
nand U2427 (N_2427,N_1657,N_1802);
or U2428 (N_2428,N_1038,N_1343);
or U2429 (N_2429,N_1756,N_1869);
nand U2430 (N_2430,N_1192,N_1983);
nand U2431 (N_2431,N_1337,N_1288);
or U2432 (N_2432,N_1507,N_1955);
and U2433 (N_2433,N_1077,N_1063);
and U2434 (N_2434,N_1584,N_1367);
nor U2435 (N_2435,N_1967,N_1431);
and U2436 (N_2436,N_1558,N_1456);
or U2437 (N_2437,N_1376,N_1843);
and U2438 (N_2438,N_1313,N_1254);
or U2439 (N_2439,N_1185,N_1933);
or U2440 (N_2440,N_1990,N_1345);
nor U2441 (N_2441,N_1965,N_1577);
and U2442 (N_2442,N_1924,N_1614);
nand U2443 (N_2443,N_1412,N_1987);
nor U2444 (N_2444,N_1446,N_1283);
or U2445 (N_2445,N_1203,N_1220);
and U2446 (N_2446,N_1394,N_1919);
or U2447 (N_2447,N_1438,N_1353);
or U2448 (N_2448,N_1293,N_1018);
nand U2449 (N_2449,N_1659,N_1384);
and U2450 (N_2450,N_1979,N_1770);
or U2451 (N_2451,N_1927,N_1153);
and U2452 (N_2452,N_1633,N_1984);
or U2453 (N_2453,N_1521,N_1226);
and U2454 (N_2454,N_1138,N_1286);
and U2455 (N_2455,N_1068,N_1562);
nand U2456 (N_2456,N_1996,N_1257);
nor U2457 (N_2457,N_1847,N_1368);
nand U2458 (N_2458,N_1448,N_1207);
nor U2459 (N_2459,N_1261,N_1913);
nand U2460 (N_2460,N_1994,N_1834);
and U2461 (N_2461,N_1108,N_1386);
nor U2462 (N_2462,N_1179,N_1472);
or U2463 (N_2463,N_1726,N_1835);
nand U2464 (N_2464,N_1864,N_1750);
or U2465 (N_2465,N_1911,N_1041);
nand U2466 (N_2466,N_1459,N_1339);
nand U2467 (N_2467,N_1793,N_1986);
nand U2468 (N_2468,N_1056,N_1592);
and U2469 (N_2469,N_1259,N_1393);
or U2470 (N_2470,N_1567,N_1191);
nand U2471 (N_2471,N_1377,N_1941);
nand U2472 (N_2472,N_1639,N_1938);
and U2473 (N_2473,N_1813,N_1713);
nor U2474 (N_2474,N_1083,N_1851);
nand U2475 (N_2475,N_1065,N_1466);
nand U2476 (N_2476,N_1439,N_1193);
nand U2477 (N_2477,N_1554,N_1003);
nor U2478 (N_2478,N_1213,N_1648);
nor U2479 (N_2479,N_1476,N_1096);
and U2480 (N_2480,N_1711,N_1424);
nor U2481 (N_2481,N_1021,N_1536);
nor U2482 (N_2482,N_1202,N_1159);
nor U2483 (N_2483,N_1169,N_1604);
and U2484 (N_2484,N_1761,N_1966);
or U2485 (N_2485,N_1069,N_1537);
nand U2486 (N_2486,N_1589,N_1150);
and U2487 (N_2487,N_1934,N_1044);
and U2488 (N_2488,N_1702,N_1450);
nand U2489 (N_2489,N_1026,N_1665);
and U2490 (N_2490,N_1097,N_1441);
or U2491 (N_2491,N_1863,N_1765);
nand U2492 (N_2492,N_1098,N_1962);
or U2493 (N_2493,N_1347,N_1939);
nor U2494 (N_2494,N_1706,N_1165);
or U2495 (N_2495,N_1297,N_1482);
or U2496 (N_2496,N_1801,N_1373);
or U2497 (N_2497,N_1071,N_1594);
nand U2498 (N_2498,N_1221,N_1708);
or U2499 (N_2499,N_1492,N_1654);
nor U2500 (N_2500,N_1084,N_1722);
or U2501 (N_2501,N_1236,N_1341);
and U2502 (N_2502,N_1625,N_1096);
nor U2503 (N_2503,N_1651,N_1224);
and U2504 (N_2504,N_1845,N_1313);
or U2505 (N_2505,N_1034,N_1424);
nor U2506 (N_2506,N_1044,N_1005);
nor U2507 (N_2507,N_1159,N_1521);
and U2508 (N_2508,N_1684,N_1980);
nand U2509 (N_2509,N_1593,N_1015);
and U2510 (N_2510,N_1322,N_1469);
nor U2511 (N_2511,N_1041,N_1247);
or U2512 (N_2512,N_1439,N_1406);
or U2513 (N_2513,N_1005,N_1064);
nand U2514 (N_2514,N_1331,N_1323);
and U2515 (N_2515,N_1889,N_1240);
and U2516 (N_2516,N_1663,N_1030);
or U2517 (N_2517,N_1344,N_1503);
or U2518 (N_2518,N_1737,N_1907);
nor U2519 (N_2519,N_1532,N_1057);
or U2520 (N_2520,N_1407,N_1043);
nand U2521 (N_2521,N_1891,N_1764);
nor U2522 (N_2522,N_1721,N_1979);
nand U2523 (N_2523,N_1680,N_1112);
and U2524 (N_2524,N_1653,N_1394);
and U2525 (N_2525,N_1994,N_1000);
and U2526 (N_2526,N_1582,N_1346);
or U2527 (N_2527,N_1352,N_1695);
nand U2528 (N_2528,N_1543,N_1545);
or U2529 (N_2529,N_1030,N_1267);
nor U2530 (N_2530,N_1219,N_1932);
nand U2531 (N_2531,N_1910,N_1528);
nor U2532 (N_2532,N_1333,N_1099);
and U2533 (N_2533,N_1722,N_1217);
nand U2534 (N_2534,N_1877,N_1284);
or U2535 (N_2535,N_1160,N_1366);
nand U2536 (N_2536,N_1711,N_1940);
nor U2537 (N_2537,N_1915,N_1327);
nor U2538 (N_2538,N_1448,N_1568);
and U2539 (N_2539,N_1740,N_1547);
or U2540 (N_2540,N_1443,N_1179);
nor U2541 (N_2541,N_1273,N_1406);
nand U2542 (N_2542,N_1437,N_1951);
nand U2543 (N_2543,N_1717,N_1959);
and U2544 (N_2544,N_1876,N_1722);
xor U2545 (N_2545,N_1809,N_1220);
nor U2546 (N_2546,N_1103,N_1246);
nor U2547 (N_2547,N_1076,N_1149);
nand U2548 (N_2548,N_1408,N_1767);
and U2549 (N_2549,N_1936,N_1003);
nand U2550 (N_2550,N_1548,N_1426);
nor U2551 (N_2551,N_1913,N_1253);
nor U2552 (N_2552,N_1800,N_1185);
and U2553 (N_2553,N_1780,N_1006);
and U2554 (N_2554,N_1787,N_1464);
nand U2555 (N_2555,N_1401,N_1235);
or U2556 (N_2556,N_1702,N_1906);
nand U2557 (N_2557,N_1223,N_1719);
nand U2558 (N_2558,N_1481,N_1594);
nor U2559 (N_2559,N_1066,N_1044);
and U2560 (N_2560,N_1673,N_1677);
or U2561 (N_2561,N_1990,N_1447);
or U2562 (N_2562,N_1660,N_1419);
nand U2563 (N_2563,N_1800,N_1934);
nor U2564 (N_2564,N_1031,N_1162);
nor U2565 (N_2565,N_1307,N_1252);
or U2566 (N_2566,N_1952,N_1011);
nor U2567 (N_2567,N_1717,N_1251);
nor U2568 (N_2568,N_1478,N_1570);
nand U2569 (N_2569,N_1905,N_1016);
and U2570 (N_2570,N_1800,N_1932);
nand U2571 (N_2571,N_1703,N_1256);
or U2572 (N_2572,N_1434,N_1521);
nand U2573 (N_2573,N_1277,N_1519);
and U2574 (N_2574,N_1925,N_1392);
or U2575 (N_2575,N_1881,N_1789);
nor U2576 (N_2576,N_1908,N_1975);
nor U2577 (N_2577,N_1347,N_1493);
and U2578 (N_2578,N_1143,N_1310);
nor U2579 (N_2579,N_1229,N_1327);
or U2580 (N_2580,N_1880,N_1191);
and U2581 (N_2581,N_1078,N_1992);
nor U2582 (N_2582,N_1756,N_1946);
or U2583 (N_2583,N_1757,N_1018);
nor U2584 (N_2584,N_1479,N_1873);
nor U2585 (N_2585,N_1843,N_1812);
nand U2586 (N_2586,N_1590,N_1845);
or U2587 (N_2587,N_1225,N_1316);
nor U2588 (N_2588,N_1067,N_1771);
nand U2589 (N_2589,N_1266,N_1848);
and U2590 (N_2590,N_1630,N_1316);
and U2591 (N_2591,N_1853,N_1004);
nand U2592 (N_2592,N_1544,N_1845);
and U2593 (N_2593,N_1629,N_1965);
nand U2594 (N_2594,N_1495,N_1118);
nand U2595 (N_2595,N_1690,N_1831);
nor U2596 (N_2596,N_1529,N_1768);
or U2597 (N_2597,N_1406,N_1428);
and U2598 (N_2598,N_1802,N_1484);
nand U2599 (N_2599,N_1271,N_1089);
nand U2600 (N_2600,N_1084,N_1316);
or U2601 (N_2601,N_1568,N_1098);
nor U2602 (N_2602,N_1372,N_1630);
or U2603 (N_2603,N_1592,N_1091);
and U2604 (N_2604,N_1339,N_1440);
nand U2605 (N_2605,N_1358,N_1261);
nand U2606 (N_2606,N_1995,N_1706);
and U2607 (N_2607,N_1891,N_1875);
nand U2608 (N_2608,N_1945,N_1555);
nor U2609 (N_2609,N_1878,N_1115);
or U2610 (N_2610,N_1613,N_1488);
nor U2611 (N_2611,N_1833,N_1997);
nand U2612 (N_2612,N_1535,N_1010);
or U2613 (N_2613,N_1659,N_1479);
nor U2614 (N_2614,N_1162,N_1479);
and U2615 (N_2615,N_1935,N_1534);
or U2616 (N_2616,N_1569,N_1062);
and U2617 (N_2617,N_1033,N_1936);
xor U2618 (N_2618,N_1708,N_1790);
and U2619 (N_2619,N_1274,N_1122);
or U2620 (N_2620,N_1106,N_1643);
nand U2621 (N_2621,N_1558,N_1288);
and U2622 (N_2622,N_1687,N_1340);
and U2623 (N_2623,N_1071,N_1240);
or U2624 (N_2624,N_1441,N_1703);
nand U2625 (N_2625,N_1164,N_1754);
nand U2626 (N_2626,N_1087,N_1215);
and U2627 (N_2627,N_1347,N_1248);
or U2628 (N_2628,N_1164,N_1272);
nand U2629 (N_2629,N_1552,N_1157);
and U2630 (N_2630,N_1648,N_1912);
or U2631 (N_2631,N_1477,N_1764);
nor U2632 (N_2632,N_1646,N_1378);
and U2633 (N_2633,N_1631,N_1410);
and U2634 (N_2634,N_1313,N_1611);
nand U2635 (N_2635,N_1764,N_1090);
and U2636 (N_2636,N_1598,N_1131);
nor U2637 (N_2637,N_1452,N_1551);
and U2638 (N_2638,N_1274,N_1933);
nand U2639 (N_2639,N_1093,N_1469);
nand U2640 (N_2640,N_1099,N_1684);
nand U2641 (N_2641,N_1171,N_1656);
xor U2642 (N_2642,N_1069,N_1640);
or U2643 (N_2643,N_1598,N_1612);
and U2644 (N_2644,N_1324,N_1516);
or U2645 (N_2645,N_1791,N_1270);
nand U2646 (N_2646,N_1009,N_1990);
nor U2647 (N_2647,N_1248,N_1720);
nand U2648 (N_2648,N_1703,N_1346);
nor U2649 (N_2649,N_1915,N_1440);
nand U2650 (N_2650,N_1921,N_1248);
nor U2651 (N_2651,N_1111,N_1489);
and U2652 (N_2652,N_1231,N_1476);
or U2653 (N_2653,N_1720,N_1381);
or U2654 (N_2654,N_1377,N_1641);
and U2655 (N_2655,N_1601,N_1735);
and U2656 (N_2656,N_1529,N_1223);
nor U2657 (N_2657,N_1884,N_1317);
nor U2658 (N_2658,N_1611,N_1578);
xor U2659 (N_2659,N_1307,N_1367);
and U2660 (N_2660,N_1030,N_1328);
or U2661 (N_2661,N_1455,N_1192);
or U2662 (N_2662,N_1499,N_1916);
nor U2663 (N_2663,N_1321,N_1745);
nor U2664 (N_2664,N_1878,N_1723);
or U2665 (N_2665,N_1533,N_1906);
or U2666 (N_2666,N_1055,N_1848);
nand U2667 (N_2667,N_1505,N_1360);
or U2668 (N_2668,N_1873,N_1845);
nor U2669 (N_2669,N_1263,N_1537);
and U2670 (N_2670,N_1138,N_1572);
nand U2671 (N_2671,N_1022,N_1828);
or U2672 (N_2672,N_1834,N_1342);
nand U2673 (N_2673,N_1548,N_1300);
nor U2674 (N_2674,N_1934,N_1668);
or U2675 (N_2675,N_1045,N_1957);
nand U2676 (N_2676,N_1612,N_1114);
or U2677 (N_2677,N_1744,N_1698);
or U2678 (N_2678,N_1265,N_1821);
xnor U2679 (N_2679,N_1026,N_1421);
and U2680 (N_2680,N_1470,N_1558);
and U2681 (N_2681,N_1134,N_1455);
or U2682 (N_2682,N_1037,N_1753);
nand U2683 (N_2683,N_1829,N_1390);
or U2684 (N_2684,N_1420,N_1143);
nor U2685 (N_2685,N_1803,N_1618);
or U2686 (N_2686,N_1735,N_1351);
and U2687 (N_2687,N_1577,N_1431);
nor U2688 (N_2688,N_1107,N_1769);
and U2689 (N_2689,N_1907,N_1432);
nor U2690 (N_2690,N_1110,N_1633);
nand U2691 (N_2691,N_1742,N_1425);
nand U2692 (N_2692,N_1933,N_1700);
nor U2693 (N_2693,N_1255,N_1650);
nand U2694 (N_2694,N_1599,N_1687);
or U2695 (N_2695,N_1889,N_1244);
or U2696 (N_2696,N_1320,N_1532);
and U2697 (N_2697,N_1774,N_1783);
nand U2698 (N_2698,N_1361,N_1818);
and U2699 (N_2699,N_1148,N_1689);
and U2700 (N_2700,N_1400,N_1768);
and U2701 (N_2701,N_1740,N_1844);
nor U2702 (N_2702,N_1474,N_1146);
nor U2703 (N_2703,N_1227,N_1268);
nor U2704 (N_2704,N_1312,N_1250);
nor U2705 (N_2705,N_1366,N_1091);
and U2706 (N_2706,N_1700,N_1052);
nand U2707 (N_2707,N_1696,N_1932);
nand U2708 (N_2708,N_1450,N_1333);
and U2709 (N_2709,N_1424,N_1502);
and U2710 (N_2710,N_1046,N_1492);
and U2711 (N_2711,N_1505,N_1955);
or U2712 (N_2712,N_1343,N_1172);
and U2713 (N_2713,N_1346,N_1821);
or U2714 (N_2714,N_1987,N_1436);
or U2715 (N_2715,N_1483,N_1165);
or U2716 (N_2716,N_1103,N_1899);
nand U2717 (N_2717,N_1640,N_1044);
nor U2718 (N_2718,N_1435,N_1888);
nand U2719 (N_2719,N_1069,N_1908);
xnor U2720 (N_2720,N_1705,N_1005);
xor U2721 (N_2721,N_1869,N_1937);
nand U2722 (N_2722,N_1671,N_1651);
xor U2723 (N_2723,N_1166,N_1651);
and U2724 (N_2724,N_1357,N_1421);
nand U2725 (N_2725,N_1087,N_1810);
nand U2726 (N_2726,N_1269,N_1777);
nor U2727 (N_2727,N_1737,N_1905);
nor U2728 (N_2728,N_1408,N_1693);
or U2729 (N_2729,N_1393,N_1225);
and U2730 (N_2730,N_1245,N_1299);
and U2731 (N_2731,N_1109,N_1437);
nand U2732 (N_2732,N_1002,N_1638);
nand U2733 (N_2733,N_1392,N_1969);
nor U2734 (N_2734,N_1721,N_1671);
and U2735 (N_2735,N_1010,N_1478);
nand U2736 (N_2736,N_1192,N_1346);
nor U2737 (N_2737,N_1028,N_1724);
or U2738 (N_2738,N_1067,N_1251);
nor U2739 (N_2739,N_1677,N_1033);
nor U2740 (N_2740,N_1460,N_1371);
nand U2741 (N_2741,N_1471,N_1909);
and U2742 (N_2742,N_1411,N_1139);
and U2743 (N_2743,N_1100,N_1160);
nor U2744 (N_2744,N_1385,N_1930);
nand U2745 (N_2745,N_1937,N_1370);
or U2746 (N_2746,N_1783,N_1518);
and U2747 (N_2747,N_1272,N_1217);
nand U2748 (N_2748,N_1064,N_1728);
nor U2749 (N_2749,N_1708,N_1907);
and U2750 (N_2750,N_1517,N_1906);
nor U2751 (N_2751,N_1832,N_1096);
and U2752 (N_2752,N_1095,N_1752);
nor U2753 (N_2753,N_1873,N_1531);
nand U2754 (N_2754,N_1667,N_1495);
and U2755 (N_2755,N_1644,N_1829);
or U2756 (N_2756,N_1363,N_1494);
nor U2757 (N_2757,N_1242,N_1140);
nor U2758 (N_2758,N_1669,N_1364);
nand U2759 (N_2759,N_1179,N_1536);
or U2760 (N_2760,N_1742,N_1034);
and U2761 (N_2761,N_1838,N_1929);
nor U2762 (N_2762,N_1165,N_1225);
nor U2763 (N_2763,N_1249,N_1343);
nand U2764 (N_2764,N_1651,N_1433);
nand U2765 (N_2765,N_1578,N_1152);
or U2766 (N_2766,N_1448,N_1344);
nor U2767 (N_2767,N_1118,N_1141);
nand U2768 (N_2768,N_1152,N_1405);
and U2769 (N_2769,N_1610,N_1764);
nor U2770 (N_2770,N_1008,N_1831);
and U2771 (N_2771,N_1550,N_1356);
or U2772 (N_2772,N_1708,N_1836);
or U2773 (N_2773,N_1828,N_1166);
nor U2774 (N_2774,N_1727,N_1254);
and U2775 (N_2775,N_1724,N_1397);
and U2776 (N_2776,N_1315,N_1277);
or U2777 (N_2777,N_1798,N_1061);
nand U2778 (N_2778,N_1256,N_1997);
nor U2779 (N_2779,N_1771,N_1090);
nor U2780 (N_2780,N_1833,N_1862);
and U2781 (N_2781,N_1087,N_1497);
nor U2782 (N_2782,N_1970,N_1661);
and U2783 (N_2783,N_1640,N_1421);
and U2784 (N_2784,N_1211,N_1100);
nor U2785 (N_2785,N_1495,N_1474);
nor U2786 (N_2786,N_1905,N_1685);
or U2787 (N_2787,N_1842,N_1477);
nand U2788 (N_2788,N_1946,N_1848);
or U2789 (N_2789,N_1429,N_1374);
or U2790 (N_2790,N_1904,N_1804);
or U2791 (N_2791,N_1773,N_1702);
nand U2792 (N_2792,N_1090,N_1337);
nand U2793 (N_2793,N_1167,N_1679);
or U2794 (N_2794,N_1612,N_1313);
nor U2795 (N_2795,N_1843,N_1746);
and U2796 (N_2796,N_1037,N_1629);
or U2797 (N_2797,N_1557,N_1255);
xnor U2798 (N_2798,N_1338,N_1187);
nor U2799 (N_2799,N_1057,N_1178);
nand U2800 (N_2800,N_1133,N_1214);
and U2801 (N_2801,N_1262,N_1086);
or U2802 (N_2802,N_1914,N_1665);
nor U2803 (N_2803,N_1880,N_1494);
or U2804 (N_2804,N_1188,N_1872);
or U2805 (N_2805,N_1397,N_1865);
nand U2806 (N_2806,N_1264,N_1580);
and U2807 (N_2807,N_1401,N_1833);
or U2808 (N_2808,N_1271,N_1728);
nor U2809 (N_2809,N_1793,N_1864);
and U2810 (N_2810,N_1277,N_1479);
xnor U2811 (N_2811,N_1658,N_1950);
or U2812 (N_2812,N_1570,N_1774);
nand U2813 (N_2813,N_1381,N_1217);
and U2814 (N_2814,N_1946,N_1610);
and U2815 (N_2815,N_1338,N_1945);
nand U2816 (N_2816,N_1146,N_1996);
nand U2817 (N_2817,N_1836,N_1266);
and U2818 (N_2818,N_1574,N_1577);
nand U2819 (N_2819,N_1370,N_1652);
nor U2820 (N_2820,N_1841,N_1754);
or U2821 (N_2821,N_1559,N_1221);
and U2822 (N_2822,N_1716,N_1509);
nor U2823 (N_2823,N_1375,N_1811);
xor U2824 (N_2824,N_1905,N_1004);
nand U2825 (N_2825,N_1435,N_1562);
or U2826 (N_2826,N_1880,N_1552);
or U2827 (N_2827,N_1693,N_1975);
and U2828 (N_2828,N_1283,N_1543);
or U2829 (N_2829,N_1875,N_1825);
nand U2830 (N_2830,N_1330,N_1895);
nor U2831 (N_2831,N_1871,N_1736);
nand U2832 (N_2832,N_1158,N_1078);
and U2833 (N_2833,N_1341,N_1749);
and U2834 (N_2834,N_1207,N_1264);
nand U2835 (N_2835,N_1266,N_1183);
nor U2836 (N_2836,N_1752,N_1796);
nor U2837 (N_2837,N_1569,N_1652);
or U2838 (N_2838,N_1471,N_1760);
nor U2839 (N_2839,N_1016,N_1488);
nand U2840 (N_2840,N_1579,N_1946);
nor U2841 (N_2841,N_1232,N_1430);
nand U2842 (N_2842,N_1990,N_1510);
xor U2843 (N_2843,N_1155,N_1650);
or U2844 (N_2844,N_1394,N_1515);
xnor U2845 (N_2845,N_1858,N_1513);
and U2846 (N_2846,N_1892,N_1213);
and U2847 (N_2847,N_1404,N_1463);
and U2848 (N_2848,N_1301,N_1311);
and U2849 (N_2849,N_1726,N_1618);
nor U2850 (N_2850,N_1145,N_1083);
or U2851 (N_2851,N_1910,N_1091);
and U2852 (N_2852,N_1636,N_1427);
or U2853 (N_2853,N_1504,N_1000);
nand U2854 (N_2854,N_1053,N_1039);
nor U2855 (N_2855,N_1379,N_1144);
nor U2856 (N_2856,N_1578,N_1258);
nand U2857 (N_2857,N_1368,N_1601);
nor U2858 (N_2858,N_1900,N_1401);
or U2859 (N_2859,N_1729,N_1224);
nand U2860 (N_2860,N_1895,N_1472);
nor U2861 (N_2861,N_1894,N_1633);
nand U2862 (N_2862,N_1814,N_1873);
or U2863 (N_2863,N_1121,N_1920);
nor U2864 (N_2864,N_1125,N_1167);
and U2865 (N_2865,N_1244,N_1722);
and U2866 (N_2866,N_1778,N_1136);
nor U2867 (N_2867,N_1646,N_1366);
or U2868 (N_2868,N_1332,N_1181);
and U2869 (N_2869,N_1926,N_1024);
nor U2870 (N_2870,N_1151,N_1034);
and U2871 (N_2871,N_1191,N_1399);
or U2872 (N_2872,N_1374,N_1141);
nand U2873 (N_2873,N_1542,N_1344);
or U2874 (N_2874,N_1348,N_1544);
nor U2875 (N_2875,N_1786,N_1236);
nor U2876 (N_2876,N_1505,N_1743);
nor U2877 (N_2877,N_1109,N_1623);
nor U2878 (N_2878,N_1563,N_1551);
nor U2879 (N_2879,N_1889,N_1748);
or U2880 (N_2880,N_1803,N_1161);
and U2881 (N_2881,N_1653,N_1389);
and U2882 (N_2882,N_1701,N_1342);
and U2883 (N_2883,N_1817,N_1418);
or U2884 (N_2884,N_1918,N_1298);
nand U2885 (N_2885,N_1570,N_1568);
and U2886 (N_2886,N_1052,N_1171);
and U2887 (N_2887,N_1418,N_1645);
and U2888 (N_2888,N_1102,N_1740);
or U2889 (N_2889,N_1530,N_1959);
or U2890 (N_2890,N_1654,N_1406);
or U2891 (N_2891,N_1102,N_1618);
or U2892 (N_2892,N_1524,N_1764);
and U2893 (N_2893,N_1444,N_1253);
nor U2894 (N_2894,N_1301,N_1037);
or U2895 (N_2895,N_1212,N_1566);
or U2896 (N_2896,N_1139,N_1099);
and U2897 (N_2897,N_1855,N_1125);
and U2898 (N_2898,N_1431,N_1903);
and U2899 (N_2899,N_1402,N_1606);
nand U2900 (N_2900,N_1247,N_1252);
nor U2901 (N_2901,N_1737,N_1807);
or U2902 (N_2902,N_1482,N_1895);
and U2903 (N_2903,N_1473,N_1895);
or U2904 (N_2904,N_1576,N_1495);
nor U2905 (N_2905,N_1243,N_1808);
or U2906 (N_2906,N_1446,N_1247);
and U2907 (N_2907,N_1782,N_1097);
or U2908 (N_2908,N_1601,N_1398);
xnor U2909 (N_2909,N_1973,N_1726);
nor U2910 (N_2910,N_1519,N_1023);
or U2911 (N_2911,N_1408,N_1336);
and U2912 (N_2912,N_1573,N_1791);
or U2913 (N_2913,N_1238,N_1473);
or U2914 (N_2914,N_1922,N_1307);
nor U2915 (N_2915,N_1463,N_1519);
nor U2916 (N_2916,N_1959,N_1146);
or U2917 (N_2917,N_1792,N_1637);
or U2918 (N_2918,N_1723,N_1569);
and U2919 (N_2919,N_1118,N_1786);
or U2920 (N_2920,N_1895,N_1920);
or U2921 (N_2921,N_1151,N_1726);
nand U2922 (N_2922,N_1861,N_1671);
xor U2923 (N_2923,N_1662,N_1335);
nor U2924 (N_2924,N_1216,N_1020);
and U2925 (N_2925,N_1177,N_1312);
and U2926 (N_2926,N_1692,N_1372);
nand U2927 (N_2927,N_1915,N_1202);
and U2928 (N_2928,N_1565,N_1246);
nand U2929 (N_2929,N_1531,N_1216);
xor U2930 (N_2930,N_1621,N_1869);
or U2931 (N_2931,N_1971,N_1582);
or U2932 (N_2932,N_1682,N_1118);
and U2933 (N_2933,N_1224,N_1857);
nand U2934 (N_2934,N_1236,N_1105);
nand U2935 (N_2935,N_1129,N_1816);
nor U2936 (N_2936,N_1390,N_1566);
nor U2937 (N_2937,N_1402,N_1544);
or U2938 (N_2938,N_1571,N_1984);
nand U2939 (N_2939,N_1325,N_1229);
nor U2940 (N_2940,N_1056,N_1805);
nor U2941 (N_2941,N_1170,N_1495);
nor U2942 (N_2942,N_1996,N_1685);
and U2943 (N_2943,N_1649,N_1385);
and U2944 (N_2944,N_1498,N_1696);
xor U2945 (N_2945,N_1345,N_1880);
nor U2946 (N_2946,N_1819,N_1936);
nand U2947 (N_2947,N_1904,N_1909);
xor U2948 (N_2948,N_1158,N_1382);
and U2949 (N_2949,N_1882,N_1004);
xor U2950 (N_2950,N_1394,N_1661);
and U2951 (N_2951,N_1032,N_1750);
or U2952 (N_2952,N_1685,N_1760);
and U2953 (N_2953,N_1078,N_1074);
nor U2954 (N_2954,N_1518,N_1525);
and U2955 (N_2955,N_1962,N_1925);
and U2956 (N_2956,N_1152,N_1121);
nand U2957 (N_2957,N_1549,N_1168);
or U2958 (N_2958,N_1093,N_1730);
nor U2959 (N_2959,N_1385,N_1430);
nor U2960 (N_2960,N_1673,N_1053);
and U2961 (N_2961,N_1385,N_1738);
nand U2962 (N_2962,N_1912,N_1398);
nand U2963 (N_2963,N_1085,N_1426);
nor U2964 (N_2964,N_1020,N_1614);
nor U2965 (N_2965,N_1429,N_1746);
or U2966 (N_2966,N_1056,N_1268);
and U2967 (N_2967,N_1045,N_1424);
nor U2968 (N_2968,N_1189,N_1395);
nor U2969 (N_2969,N_1060,N_1791);
xnor U2970 (N_2970,N_1644,N_1082);
xor U2971 (N_2971,N_1159,N_1750);
nor U2972 (N_2972,N_1219,N_1446);
or U2973 (N_2973,N_1449,N_1149);
and U2974 (N_2974,N_1780,N_1498);
nor U2975 (N_2975,N_1523,N_1837);
nand U2976 (N_2976,N_1702,N_1633);
or U2977 (N_2977,N_1161,N_1689);
or U2978 (N_2978,N_1195,N_1184);
or U2979 (N_2979,N_1607,N_1114);
nand U2980 (N_2980,N_1333,N_1578);
or U2981 (N_2981,N_1949,N_1270);
nand U2982 (N_2982,N_1925,N_1261);
nor U2983 (N_2983,N_1305,N_1089);
and U2984 (N_2984,N_1267,N_1052);
or U2985 (N_2985,N_1906,N_1475);
nor U2986 (N_2986,N_1244,N_1411);
or U2987 (N_2987,N_1645,N_1959);
or U2988 (N_2988,N_1759,N_1725);
nand U2989 (N_2989,N_1157,N_1179);
and U2990 (N_2990,N_1031,N_1271);
and U2991 (N_2991,N_1492,N_1006);
or U2992 (N_2992,N_1212,N_1816);
and U2993 (N_2993,N_1344,N_1792);
or U2994 (N_2994,N_1760,N_1901);
or U2995 (N_2995,N_1205,N_1346);
xor U2996 (N_2996,N_1525,N_1074);
or U2997 (N_2997,N_1744,N_1939);
xor U2998 (N_2998,N_1352,N_1855);
or U2999 (N_2999,N_1756,N_1219);
nor UO_0 (O_0,N_2043,N_2029);
nor UO_1 (O_1,N_2066,N_2440);
nand UO_2 (O_2,N_2719,N_2847);
or UO_3 (O_3,N_2574,N_2340);
or UO_4 (O_4,N_2800,N_2081);
nor UO_5 (O_5,N_2497,N_2271);
nand UO_6 (O_6,N_2698,N_2456);
nand UO_7 (O_7,N_2225,N_2390);
nor UO_8 (O_8,N_2695,N_2069);
and UO_9 (O_9,N_2203,N_2825);
nor UO_10 (O_10,N_2108,N_2495);
or UO_11 (O_11,N_2168,N_2607);
nand UO_12 (O_12,N_2504,N_2701);
and UO_13 (O_13,N_2486,N_2033);
and UO_14 (O_14,N_2062,N_2822);
nand UO_15 (O_15,N_2065,N_2215);
nand UO_16 (O_16,N_2393,N_2539);
nand UO_17 (O_17,N_2529,N_2976);
nand UO_18 (O_18,N_2214,N_2133);
nor UO_19 (O_19,N_2363,N_2293);
and UO_20 (O_20,N_2230,N_2110);
nand UO_21 (O_21,N_2921,N_2312);
and UO_22 (O_22,N_2437,N_2920);
and UO_23 (O_23,N_2439,N_2139);
xor UO_24 (O_24,N_2585,N_2469);
nand UO_25 (O_25,N_2858,N_2808);
or UO_26 (O_26,N_2927,N_2697);
nor UO_27 (O_27,N_2406,N_2886);
nand UO_28 (O_28,N_2678,N_2008);
nor UO_29 (O_29,N_2127,N_2465);
and UO_30 (O_30,N_2028,N_2377);
and UO_31 (O_31,N_2019,N_2454);
and UO_32 (O_32,N_2334,N_2746);
and UO_33 (O_33,N_2654,N_2897);
and UO_34 (O_34,N_2975,N_2207);
nor UO_35 (O_35,N_2423,N_2167);
or UO_36 (O_36,N_2570,N_2755);
or UO_37 (O_37,N_2200,N_2226);
nand UO_38 (O_38,N_2795,N_2217);
nor UO_39 (O_39,N_2621,N_2474);
and UO_40 (O_40,N_2670,N_2748);
and UO_41 (O_41,N_2900,N_2205);
nor UO_42 (O_42,N_2606,N_2164);
or UO_43 (O_43,N_2949,N_2269);
and UO_44 (O_44,N_2517,N_2741);
nor UO_45 (O_45,N_2275,N_2890);
and UO_46 (O_46,N_2496,N_2535);
or UO_47 (O_47,N_2742,N_2191);
and UO_48 (O_48,N_2561,N_2418);
nand UO_49 (O_49,N_2716,N_2209);
and UO_50 (O_50,N_2778,N_2193);
nand UO_51 (O_51,N_2750,N_2893);
and UO_52 (O_52,N_2591,N_2389);
nor UO_53 (O_53,N_2986,N_2728);
xor UO_54 (O_54,N_2173,N_2202);
or UO_55 (O_55,N_2556,N_2219);
nor UO_56 (O_56,N_2938,N_2245);
nand UO_57 (O_57,N_2338,N_2336);
and UO_58 (O_58,N_2749,N_2330);
nand UO_59 (O_59,N_2305,N_2569);
and UO_60 (O_60,N_2930,N_2727);
and UO_61 (O_61,N_2672,N_2699);
and UO_62 (O_62,N_2025,N_2684);
or UO_63 (O_63,N_2589,N_2160);
nand UO_64 (O_64,N_2396,N_2934);
nand UO_65 (O_65,N_2853,N_2899);
nor UO_66 (O_66,N_2425,N_2368);
and UO_67 (O_67,N_2973,N_2652);
and UO_68 (O_68,N_2877,N_2827);
nor UO_69 (O_69,N_2985,N_2040);
nand UO_70 (O_70,N_2554,N_2462);
nand UO_71 (O_71,N_2012,N_2669);
or UO_72 (O_72,N_2067,N_2460);
or UO_73 (O_73,N_2981,N_2061);
and UO_74 (O_74,N_2763,N_2736);
and UO_75 (O_75,N_2918,N_2611);
or UO_76 (O_76,N_2919,N_2557);
nand UO_77 (O_77,N_2357,N_2280);
nor UO_78 (O_78,N_2403,N_2979);
nor UO_79 (O_79,N_2154,N_2449);
xnor UO_80 (O_80,N_2384,N_2265);
nand UO_81 (O_81,N_2325,N_2789);
and UO_82 (O_82,N_2461,N_2744);
and UO_83 (O_83,N_2580,N_2731);
or UO_84 (O_84,N_2596,N_2568);
and UO_85 (O_85,N_2941,N_2564);
or UO_86 (O_86,N_2706,N_2766);
or UO_87 (O_87,N_2958,N_2060);
or UO_88 (O_88,N_2785,N_2242);
and UO_89 (O_89,N_2448,N_2723);
nand UO_90 (O_90,N_2655,N_2031);
nor UO_91 (O_91,N_2828,N_2122);
nor UO_92 (O_92,N_2391,N_2013);
nand UO_93 (O_93,N_2965,N_2246);
nor UO_94 (O_94,N_2768,N_2422);
or UO_95 (O_95,N_2544,N_2240);
nor UO_96 (O_96,N_2453,N_2722);
and UO_97 (O_97,N_2832,N_2912);
and UO_98 (O_98,N_2306,N_2288);
or UO_99 (O_99,N_2296,N_2049);
or UO_100 (O_100,N_2547,N_2106);
nor UO_101 (O_101,N_2745,N_2186);
or UO_102 (O_102,N_2199,N_2213);
and UO_103 (O_103,N_2261,N_2378);
nor UO_104 (O_104,N_2364,N_2104);
xor UO_105 (O_105,N_2253,N_2468);
nor UO_106 (O_106,N_2907,N_2705);
and UO_107 (O_107,N_2720,N_2473);
nor UO_108 (O_108,N_2908,N_2955);
nor UO_109 (O_109,N_2775,N_2183);
or UO_110 (O_110,N_2159,N_2614);
and UO_111 (O_111,N_2002,N_2010);
nand UO_112 (O_112,N_2408,N_2479);
nor UO_113 (O_113,N_2414,N_2272);
nand UO_114 (O_114,N_2546,N_2201);
and UO_115 (O_115,N_2952,N_2349);
or UO_116 (O_116,N_2874,N_2058);
xnor UO_117 (O_117,N_2507,N_2519);
and UO_118 (O_118,N_2576,N_2289);
and UO_119 (O_119,N_2099,N_2683);
or UO_120 (O_120,N_2567,N_2345);
nand UO_121 (O_121,N_2928,N_2650);
and UO_122 (O_122,N_2362,N_2532);
or UO_123 (O_123,N_2274,N_2512);
or UO_124 (O_124,N_2365,N_2688);
or UO_125 (O_125,N_2888,N_2055);
or UO_126 (O_126,N_2170,N_2664);
nand UO_127 (O_127,N_2045,N_2590);
and UO_128 (O_128,N_2870,N_2150);
nand UO_129 (O_129,N_2627,N_2035);
or UO_130 (O_130,N_2392,N_2014);
and UO_131 (O_131,N_2846,N_2600);
or UO_132 (O_132,N_2320,N_2096);
and UO_133 (O_133,N_2476,N_2759);
and UO_134 (O_134,N_2830,N_2906);
and UO_135 (O_135,N_2936,N_2407);
or UO_136 (O_136,N_2374,N_2229);
or UO_137 (O_137,N_2884,N_2109);
and UO_138 (O_138,N_2948,N_2256);
or UO_139 (O_139,N_2451,N_2634);
nor UO_140 (O_140,N_2732,N_2550);
or UO_141 (O_141,N_2797,N_2356);
or UO_142 (O_142,N_2982,N_2583);
nor UO_143 (O_143,N_2447,N_2904);
and UO_144 (O_144,N_2779,N_2690);
or UO_145 (O_145,N_2794,N_2558);
nor UO_146 (O_146,N_2006,N_2347);
and UO_147 (O_147,N_2135,N_2780);
or UO_148 (O_148,N_2761,N_2582);
nand UO_149 (O_149,N_2604,N_2560);
and UO_150 (O_150,N_2679,N_2141);
and UO_151 (O_151,N_2433,N_2501);
nand UO_152 (O_152,N_2854,N_2087);
nand UO_153 (O_153,N_2233,N_2824);
and UO_154 (O_154,N_2594,N_2331);
and UO_155 (O_155,N_2381,N_2300);
nor UO_156 (O_156,N_2513,N_2971);
or UO_157 (O_157,N_2876,N_2277);
and UO_158 (O_158,N_2514,N_2605);
nor UO_159 (O_159,N_2799,N_2542);
nand UO_160 (O_160,N_2434,N_2939);
nor UO_161 (O_161,N_2562,N_2673);
and UO_162 (O_162,N_2659,N_2909);
nand UO_163 (O_163,N_2942,N_2538);
or UO_164 (O_164,N_2953,N_2868);
nor UO_165 (O_165,N_2711,N_2793);
nor UO_166 (O_166,N_2831,N_2735);
or UO_167 (O_167,N_2767,N_2691);
nor UO_168 (O_168,N_2675,N_2086);
nand UO_169 (O_169,N_2656,N_2136);
and UO_170 (O_170,N_2489,N_2103);
nand UO_171 (O_171,N_2641,N_2301);
or UO_172 (O_172,N_2525,N_2506);
or UO_173 (O_173,N_2865,N_2635);
nor UO_174 (O_174,N_2917,N_2487);
nor UO_175 (O_175,N_2329,N_2508);
or UO_176 (O_176,N_2577,N_2313);
nor UO_177 (O_177,N_2179,N_2764);
or UO_178 (O_178,N_2578,N_2208);
and UO_179 (O_179,N_2385,N_2250);
or UO_180 (O_180,N_2470,N_2176);
and UO_181 (O_181,N_2395,N_2812);
and UO_182 (O_182,N_2102,N_2530);
nor UO_183 (O_183,N_2171,N_2282);
and UO_184 (O_184,N_2236,N_2798);
nand UO_185 (O_185,N_2592,N_2639);
and UO_186 (O_186,N_2383,N_2297);
nand UO_187 (O_187,N_2784,N_2216);
or UO_188 (O_188,N_2581,N_2318);
or UO_189 (O_189,N_2411,N_2420);
nor UO_190 (O_190,N_2792,N_2911);
and UO_191 (O_191,N_2471,N_2760);
nand UO_192 (O_192,N_2980,N_2056);
and UO_193 (O_193,N_2555,N_2490);
nand UO_194 (O_194,N_2503,N_2991);
and UO_195 (O_195,N_2015,N_2630);
and UO_196 (O_196,N_2105,N_2817);
or UO_197 (O_197,N_2276,N_2048);
and UO_198 (O_198,N_2195,N_2042);
or UO_199 (O_199,N_2073,N_2116);
and UO_200 (O_200,N_2211,N_2839);
nor UO_201 (O_201,N_2153,N_2358);
nand UO_202 (O_202,N_2052,N_2409);
nand UO_203 (O_203,N_2316,N_2348);
and UO_204 (O_204,N_2412,N_2394);
nand UO_205 (O_205,N_2260,N_2126);
nand UO_206 (O_206,N_2146,N_2492);
and UO_207 (O_207,N_2415,N_2840);
nand UO_208 (O_208,N_2129,N_2163);
or UO_209 (O_209,N_2247,N_2889);
nor UO_210 (O_210,N_2252,N_2954);
or UO_211 (O_211,N_2835,N_2923);
nor UO_212 (O_212,N_2838,N_2047);
nor UO_213 (O_213,N_2397,N_2198);
and UO_214 (O_214,N_2937,N_2145);
nand UO_215 (O_215,N_2521,N_2815);
or UO_216 (O_216,N_2806,N_2227);
or UO_217 (O_217,N_2483,N_2180);
nand UO_218 (O_218,N_2914,N_2232);
or UO_219 (O_219,N_2323,N_2989);
nor UO_220 (O_220,N_2801,N_2730);
and UO_221 (O_221,N_2662,N_2873);
and UO_222 (O_222,N_2903,N_2834);
nor UO_223 (O_223,N_2974,N_2175);
or UO_224 (O_224,N_2050,N_2712);
and UO_225 (O_225,N_2729,N_2053);
nor UO_226 (O_226,N_2452,N_2431);
and UO_227 (O_227,N_2855,N_2617);
or UO_228 (O_228,N_2118,N_2072);
nor UO_229 (O_229,N_2960,N_2622);
nand UO_230 (O_230,N_2161,N_2291);
and UO_231 (O_231,N_2776,N_2113);
nand UO_232 (O_232,N_2543,N_2816);
nor UO_233 (O_233,N_2837,N_2399);
nor UO_234 (O_234,N_2077,N_2303);
nor UO_235 (O_235,N_2472,N_2457);
nor UO_236 (O_236,N_2147,N_2314);
or UO_237 (O_237,N_2355,N_2651);
nand UO_238 (O_238,N_2281,N_2572);
nand UO_239 (O_239,N_2726,N_2883);
and UO_240 (O_240,N_2427,N_2125);
nand UO_241 (O_241,N_2267,N_2114);
xor UO_242 (O_242,N_2747,N_2710);
and UO_243 (O_243,N_2255,N_2660);
and UO_244 (O_244,N_2970,N_2545);
nor UO_245 (O_245,N_2945,N_2803);
and UO_246 (O_246,N_2696,N_2478);
and UO_247 (O_247,N_2196,N_2894);
nor UO_248 (O_248,N_2511,N_2983);
nand UO_249 (O_249,N_2243,N_2769);
and UO_250 (O_250,N_2445,N_2814);
nor UO_251 (O_251,N_2804,N_2262);
nor UO_252 (O_252,N_2140,N_2857);
nor UO_253 (O_253,N_2095,N_2387);
or UO_254 (O_254,N_2924,N_2444);
or UO_255 (O_255,N_2925,N_2234);
or UO_256 (O_256,N_2823,N_2682);
nand UO_257 (O_257,N_2740,N_2608);
and UO_258 (O_258,N_2626,N_2707);
nor UO_259 (O_259,N_2629,N_2790);
or UO_260 (O_260,N_2661,N_2802);
nand UO_261 (O_261,N_2017,N_2926);
and UO_262 (O_262,N_2343,N_2184);
or UO_263 (O_263,N_2772,N_2488);
and UO_264 (O_264,N_2413,N_2177);
or UO_265 (O_265,N_2645,N_2382);
and UO_266 (O_266,N_2957,N_2197);
xor UO_267 (O_267,N_2480,N_2668);
nor UO_268 (O_268,N_2676,N_2999);
or UO_269 (O_269,N_2027,N_2148);
and UO_270 (O_270,N_2714,N_2475);
nand UO_271 (O_271,N_2637,N_2977);
nand UO_272 (O_272,N_2352,N_2872);
nor UO_273 (O_273,N_2571,N_2222);
nor UO_274 (O_274,N_2443,N_2950);
nor UO_275 (O_275,N_2204,N_2036);
or UO_276 (O_276,N_2088,N_2351);
or UO_277 (O_277,N_2692,N_2943);
or UO_278 (O_278,N_2713,N_2324);
nor UO_279 (O_279,N_2674,N_2625);
or UO_280 (O_280,N_2107,N_2494);
nand UO_281 (O_281,N_2644,N_2597);
and UO_282 (O_282,N_2956,N_2235);
nor UO_283 (O_283,N_2360,N_2375);
or UO_284 (O_284,N_2573,N_2717);
nor UO_285 (O_285,N_2285,N_2315);
and UO_286 (O_286,N_2063,N_2094);
or UO_287 (O_287,N_2026,N_2595);
nor UO_288 (O_288,N_2947,N_2988);
nand UO_289 (O_289,N_2231,N_2859);
nand UO_290 (O_290,N_2671,N_2738);
nor UO_291 (O_291,N_2498,N_2818);
nand UO_292 (O_292,N_2079,N_2820);
or UO_293 (O_293,N_2613,N_2638);
nand UO_294 (O_294,N_2327,N_2083);
nor UO_295 (O_295,N_2238,N_2528);
nand UO_296 (O_296,N_2221,N_2218);
nor UO_297 (O_297,N_2693,N_2155);
and UO_298 (O_298,N_2601,N_2781);
nor UO_299 (O_299,N_2533,N_2166);
and UO_300 (O_300,N_2700,N_2032);
and UO_301 (O_301,N_2867,N_2860);
nand UO_302 (O_302,N_2491,N_2584);
nor UO_303 (O_303,N_2875,N_2777);
and UO_304 (O_304,N_2034,N_2376);
and UO_305 (O_305,N_2257,N_2852);
or UO_306 (O_306,N_2003,N_2130);
or UO_307 (O_307,N_2144,N_2885);
nor UO_308 (O_308,N_2322,N_2881);
and UO_309 (O_309,N_2359,N_2092);
nand UO_310 (O_310,N_2754,N_2115);
or UO_311 (O_311,N_2553,N_2344);
nand UO_312 (O_312,N_2085,N_2984);
or UO_313 (O_313,N_2442,N_2786);
nand UO_314 (O_314,N_2510,N_2882);
nor UO_315 (O_315,N_2270,N_2878);
nor UO_316 (O_316,N_2829,N_2657);
or UO_317 (O_317,N_2551,N_2266);
or UO_318 (O_318,N_2430,N_2464);
nor UO_319 (O_319,N_2765,N_2987);
and UO_320 (O_320,N_2080,N_2286);
nand UO_321 (O_321,N_2251,N_2120);
and UO_322 (O_322,N_2350,N_2354);
and UO_323 (O_323,N_2123,N_2481);
or UO_324 (O_324,N_2646,N_2694);
nor UO_325 (O_325,N_2658,N_2178);
or UO_326 (O_326,N_2940,N_2076);
or UO_327 (O_327,N_2398,N_2739);
nor UO_328 (O_328,N_2887,N_2500);
or UO_329 (O_329,N_2810,N_2905);
nor UO_330 (O_330,N_2640,N_2421);
or UO_331 (O_331,N_2969,N_2902);
nand UO_332 (O_332,N_2826,N_2212);
and UO_333 (O_333,N_2933,N_2616);
or UO_334 (O_334,N_2993,N_2548);
or UO_335 (O_335,N_2680,N_2435);
or UO_336 (O_336,N_2400,N_2968);
nor UO_337 (O_337,N_2466,N_2192);
nand UO_338 (O_338,N_2609,N_2326);
nand UO_339 (O_339,N_2901,N_2278);
xor UO_340 (O_340,N_2997,N_2681);
or UO_341 (O_341,N_2788,N_2758);
or UO_342 (O_342,N_2011,N_2455);
nor UO_343 (O_343,N_2961,N_2405);
nor UO_344 (O_344,N_2292,N_2733);
nor UO_345 (O_345,N_2169,N_2084);
or UO_346 (O_346,N_2518,N_2963);
nand UO_347 (O_347,N_2485,N_2091);
nand UO_348 (O_348,N_2038,N_2866);
nand UO_349 (O_349,N_2703,N_2037);
or UO_350 (O_350,N_2811,N_2051);
or UO_351 (O_351,N_2307,N_2054);
and UO_352 (O_352,N_2515,N_2372);
or UO_353 (O_353,N_2715,N_2337);
nor UO_354 (O_354,N_2039,N_2782);
nor UO_355 (O_355,N_2241,N_2220);
or UO_356 (O_356,N_2524,N_2636);
xnor UO_357 (O_357,N_2725,N_2704);
nor UO_358 (O_358,N_2516,N_2962);
and UO_359 (O_359,N_2841,N_2845);
or UO_360 (O_360,N_2346,N_2990);
and UO_361 (O_361,N_2821,N_2332);
nor UO_362 (O_362,N_2353,N_2467);
or UO_363 (O_363,N_2724,N_2522);
nor UO_364 (O_364,N_2188,N_2311);
nor UO_365 (O_365,N_2935,N_2774);
and UO_366 (O_366,N_2157,N_2946);
nor UO_367 (O_367,N_2182,N_2268);
nand UO_368 (O_368,N_2996,N_2000);
and UO_369 (O_369,N_2005,N_2531);
nand UO_370 (O_370,N_2057,N_2290);
and UO_371 (O_371,N_2041,N_2566);
and UO_372 (O_372,N_2295,N_2895);
nand UO_373 (O_373,N_2787,N_2308);
nor UO_374 (O_374,N_2653,N_2438);
nor UO_375 (O_375,N_2709,N_2417);
and UO_376 (O_376,N_2602,N_2426);
or UO_377 (O_377,N_2059,N_2813);
nand UO_378 (O_378,N_2441,N_2138);
or UO_379 (O_379,N_2972,N_2022);
or UO_380 (O_380,N_2023,N_2624);
and UO_381 (O_381,N_2112,N_2922);
nand UO_382 (O_382,N_2064,N_2537);
or UO_383 (O_383,N_2223,N_2194);
or UO_384 (O_384,N_2879,N_2520);
nor UO_385 (O_385,N_2298,N_2910);
and UO_386 (O_386,N_2366,N_2482);
nand UO_387 (O_387,N_2552,N_2864);
or UO_388 (O_388,N_2689,N_2228);
nand UO_389 (O_389,N_2898,N_2666);
nor UO_390 (O_390,N_2317,N_2913);
and UO_391 (O_391,N_2001,N_2030);
or UO_392 (O_392,N_2967,N_2579);
or UO_393 (O_393,N_2143,N_2089);
nor UO_394 (O_394,N_2379,N_2007);
nand UO_395 (O_395,N_2565,N_2304);
or UO_396 (O_396,N_2998,N_2009);
and UO_397 (O_397,N_2299,N_2459);
nand UO_398 (O_398,N_2428,N_2410);
and UO_399 (O_399,N_2623,N_2279);
and UO_400 (O_400,N_2090,N_2302);
or UO_401 (O_401,N_2502,N_2540);
nand UO_402 (O_402,N_2162,N_2142);
nand UO_403 (O_403,N_2931,N_2563);
nand UO_404 (O_404,N_2667,N_2401);
and UO_405 (O_405,N_2446,N_2751);
nor UO_406 (O_406,N_2631,N_2335);
or UO_407 (O_407,N_2239,N_2371);
nand UO_408 (O_408,N_2734,N_2068);
and UO_409 (O_409,N_2493,N_2369);
and UO_410 (O_410,N_2074,N_2424);
and UO_411 (O_411,N_2499,N_2752);
or UO_412 (O_412,N_2137,N_2757);
nor UO_413 (O_413,N_2149,N_2992);
and UO_414 (O_414,N_2131,N_2458);
nor UO_415 (O_415,N_2342,N_2254);
or UO_416 (O_416,N_2809,N_2310);
and UO_417 (O_417,N_2783,N_2756);
or UO_418 (O_418,N_2134,N_2534);
nand UO_419 (O_419,N_2849,N_2586);
nand UO_420 (O_420,N_2477,N_2649);
nor UO_421 (O_421,N_2593,N_2258);
nor UO_422 (O_422,N_2093,N_2686);
nand UO_423 (O_423,N_2773,N_2844);
nand UO_424 (O_424,N_2848,N_2020);
nand UO_425 (O_425,N_2588,N_2891);
xor UO_426 (O_426,N_2615,N_2156);
nor UO_427 (O_427,N_2259,N_2319);
nor UO_428 (O_428,N_2484,N_2549);
nor UO_429 (O_429,N_2861,N_2187);
nor UO_430 (O_430,N_2172,N_2805);
and UO_431 (O_431,N_2018,N_2620);
nor UO_432 (O_432,N_2509,N_2836);
nor UO_433 (O_433,N_2328,N_2959);
nor UO_434 (O_434,N_2612,N_2665);
nand UO_435 (O_435,N_2599,N_2128);
or UO_436 (O_436,N_2158,N_2648);
nor UO_437 (O_437,N_2932,N_2915);
or UO_438 (O_438,N_2929,N_2819);
nor UO_439 (O_439,N_2995,N_2851);
nor UO_440 (O_440,N_2044,N_2070);
and UO_441 (O_441,N_2097,N_2856);
and UO_442 (O_442,N_2436,N_2450);
nand UO_443 (O_443,N_2463,N_2124);
and UO_444 (O_444,N_2370,N_2892);
nand UO_445 (O_445,N_2964,N_2016);
nand UO_446 (O_446,N_2951,N_2708);
nor UO_447 (O_447,N_2284,N_2633);
and UO_448 (O_448,N_2341,N_2121);
and UO_449 (O_449,N_2863,N_2966);
nand UO_450 (O_450,N_2046,N_2249);
and UO_451 (O_451,N_2807,N_2082);
and UO_452 (O_452,N_2432,N_2587);
or UO_453 (O_453,N_2685,N_2206);
xnor UO_454 (O_454,N_2174,N_2796);
nor UO_455 (O_455,N_2619,N_2185);
nand UO_456 (O_456,N_2264,N_2021);
nand UO_457 (O_457,N_2404,N_2618);
nor UO_458 (O_458,N_2833,N_2598);
or UO_459 (O_459,N_2843,N_2559);
and UO_460 (O_460,N_2119,N_2388);
nor UO_461 (O_461,N_2263,N_2224);
and UO_462 (O_462,N_2603,N_2632);
nand UO_463 (O_463,N_2075,N_2244);
xor UO_464 (O_464,N_2994,N_2541);
nor UO_465 (O_465,N_2287,N_2416);
nand UO_466 (O_466,N_2944,N_2189);
or UO_467 (O_467,N_2283,N_2737);
nor UO_468 (O_468,N_2101,N_2210);
nor UO_469 (O_469,N_2718,N_2643);
nand UO_470 (O_470,N_2294,N_2869);
or UO_471 (O_471,N_2321,N_2402);
or UO_472 (O_472,N_2373,N_2871);
nand UO_473 (O_473,N_2100,N_2791);
nor UO_474 (O_474,N_2527,N_2610);
and UO_475 (O_475,N_2762,N_2663);
and UO_476 (O_476,N_2111,N_2880);
nand UO_477 (O_477,N_2190,N_2628);
or UO_478 (O_478,N_2575,N_2677);
nor UO_479 (O_479,N_2850,N_2526);
nor UO_480 (O_480,N_2721,N_2024);
or UO_481 (O_481,N_2339,N_2181);
nor UO_482 (O_482,N_2523,N_2248);
nor UO_483 (O_483,N_2743,N_2132);
or UO_484 (O_484,N_2165,N_2896);
nor UO_485 (O_485,N_2333,N_2505);
and UO_486 (O_486,N_2361,N_2419);
nor UO_487 (O_487,N_2770,N_2386);
and UO_488 (O_488,N_2429,N_2152);
and UO_489 (O_489,N_2071,N_2004);
nand UO_490 (O_490,N_2978,N_2117);
or UO_491 (O_491,N_2771,N_2078);
nand UO_492 (O_492,N_2380,N_2151);
or UO_493 (O_493,N_2273,N_2702);
nand UO_494 (O_494,N_2536,N_2862);
or UO_495 (O_495,N_2842,N_2916);
xnor UO_496 (O_496,N_2367,N_2098);
and UO_497 (O_497,N_2237,N_2687);
nand UO_498 (O_498,N_2309,N_2642);
nand UO_499 (O_499,N_2753,N_2647);
endmodule