module basic_1000_10000_1500_50_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_242,In_964);
and U1 (N_1,In_42,In_335);
nor U2 (N_2,In_220,In_650);
nand U3 (N_3,In_171,In_752);
nor U4 (N_4,In_622,In_380);
and U5 (N_5,In_515,In_336);
and U6 (N_6,In_233,In_236);
or U7 (N_7,In_549,In_929);
or U8 (N_8,In_900,In_391);
nand U9 (N_9,In_795,In_701);
xnor U10 (N_10,In_405,In_50);
xor U11 (N_11,In_30,In_189);
nand U12 (N_12,In_247,In_545);
and U13 (N_13,In_522,In_858);
nand U14 (N_14,In_796,In_175);
nor U15 (N_15,In_847,In_610);
nor U16 (N_16,In_994,In_925);
nor U17 (N_17,In_750,In_412);
nor U18 (N_18,In_587,In_179);
nor U19 (N_19,In_376,In_834);
and U20 (N_20,In_79,In_846);
nand U21 (N_21,In_18,In_867);
or U22 (N_22,In_197,In_347);
nand U23 (N_23,In_161,In_895);
nor U24 (N_24,In_186,In_300);
and U25 (N_25,In_501,In_539);
nand U26 (N_26,In_629,In_862);
xnor U27 (N_27,In_209,In_26);
and U28 (N_28,In_960,In_893);
nor U29 (N_29,In_86,In_309);
or U30 (N_30,In_708,In_681);
nand U31 (N_31,In_368,In_976);
and U32 (N_32,In_147,In_955);
xor U33 (N_33,In_485,In_678);
nor U34 (N_34,In_855,In_593);
and U35 (N_35,In_136,In_879);
or U36 (N_36,In_956,In_34);
nor U37 (N_37,In_148,In_452);
nor U38 (N_38,In_384,In_657);
nand U39 (N_39,In_748,In_154);
nand U40 (N_40,In_824,In_513);
xnor U41 (N_41,In_205,In_794);
or U42 (N_42,In_224,In_397);
nand U43 (N_43,In_17,In_516);
and U44 (N_44,In_658,In_971);
nand U45 (N_45,In_385,In_98);
nand U46 (N_46,In_825,In_132);
nand U47 (N_47,In_281,In_108);
nor U48 (N_48,In_965,In_341);
nor U49 (N_49,In_201,In_835);
nor U50 (N_50,In_936,In_266);
nand U51 (N_51,In_655,In_686);
nor U52 (N_52,In_454,In_69);
and U53 (N_53,In_554,In_364);
xnor U54 (N_54,In_781,In_393);
or U55 (N_55,In_354,In_520);
or U56 (N_56,In_100,In_315);
xor U57 (N_57,In_165,In_723);
nor U58 (N_58,In_221,In_45);
or U59 (N_59,In_359,In_427);
and U60 (N_60,In_959,In_606);
or U61 (N_61,In_537,In_51);
xor U62 (N_62,In_719,In_143);
nor U63 (N_63,In_754,In_417);
nand U64 (N_64,In_730,In_637);
or U65 (N_65,In_429,In_386);
or U66 (N_66,In_901,In_41);
or U67 (N_67,In_909,In_786);
nand U68 (N_68,In_255,In_96);
and U69 (N_69,In_387,In_667);
xor U70 (N_70,In_902,In_728);
nand U71 (N_71,In_897,In_431);
nor U72 (N_72,In_478,In_511);
nand U73 (N_73,In_905,In_624);
nor U74 (N_74,In_910,In_532);
or U75 (N_75,In_396,In_72);
nand U76 (N_76,In_816,In_665);
or U77 (N_77,In_115,In_907);
nand U78 (N_78,In_456,In_920);
or U79 (N_79,In_12,In_872);
and U80 (N_80,In_293,In_107);
or U81 (N_81,In_371,In_819);
and U82 (N_82,In_267,In_174);
or U83 (N_83,In_196,In_297);
or U84 (N_84,In_878,In_704);
nand U85 (N_85,In_156,In_225);
xor U86 (N_86,In_780,In_131);
and U87 (N_87,In_285,In_235);
or U88 (N_88,In_164,In_152);
nand U89 (N_89,In_813,In_725);
nor U90 (N_90,In_601,In_477);
or U91 (N_91,In_807,In_635);
nor U92 (N_92,In_882,In_552);
nor U93 (N_93,In_425,In_614);
or U94 (N_94,In_198,In_159);
and U95 (N_95,In_973,In_519);
or U96 (N_96,In_767,In_863);
nand U97 (N_97,In_696,In_842);
and U98 (N_98,In_663,In_646);
nor U99 (N_99,In_258,In_617);
nor U100 (N_100,In_713,In_495);
or U101 (N_101,In_660,In_978);
nor U102 (N_102,In_38,In_669);
nand U103 (N_103,In_13,In_88);
or U104 (N_104,In_721,In_782);
or U105 (N_105,In_349,In_560);
nor U106 (N_106,In_49,In_351);
nor U107 (N_107,In_303,In_679);
or U108 (N_108,In_697,In_649);
and U109 (N_109,In_944,In_917);
or U110 (N_110,In_125,In_54);
nor U111 (N_111,In_765,In_6);
and U112 (N_112,In_590,In_366);
nand U113 (N_113,In_906,In_158);
nor U114 (N_114,In_742,In_567);
xor U115 (N_115,In_968,In_533);
and U116 (N_116,In_287,In_972);
nor U117 (N_117,In_231,In_426);
or U118 (N_118,In_966,In_317);
nor U119 (N_119,In_607,In_555);
and U120 (N_120,In_316,In_237);
nand U121 (N_121,In_591,In_67);
or U122 (N_122,In_430,In_980);
nor U123 (N_123,In_421,In_117);
and U124 (N_124,In_250,In_949);
or U125 (N_125,In_451,In_603);
and U126 (N_126,In_10,In_62);
nor U127 (N_127,In_135,In_428);
nor U128 (N_128,In_999,In_463);
nand U129 (N_129,In_302,In_940);
or U130 (N_130,In_140,In_975);
nor U131 (N_131,In_234,In_640);
nand U132 (N_132,In_656,In_358);
and U133 (N_133,In_784,In_155);
or U134 (N_134,In_829,In_307);
nand U135 (N_135,In_283,In_841);
nand U136 (N_136,In_203,In_691);
or U137 (N_137,In_311,In_71);
xnor U138 (N_138,In_129,In_547);
or U139 (N_139,In_103,In_321);
and U140 (N_140,In_613,In_791);
xnor U141 (N_141,In_184,In_828);
nand U142 (N_142,In_861,In_680);
nor U143 (N_143,In_373,In_296);
and U144 (N_144,In_566,In_832);
or U145 (N_145,In_180,In_333);
nand U146 (N_146,In_468,In_268);
and U147 (N_147,In_584,In_724);
or U148 (N_148,In_772,In_469);
or U149 (N_149,In_625,In_390);
nor U150 (N_150,In_888,In_729);
or U151 (N_151,In_139,In_749);
or U152 (N_152,In_173,In_743);
nor U153 (N_153,In_213,In_798);
nand U154 (N_154,In_239,In_407);
or U155 (N_155,In_602,In_588);
nand U156 (N_156,In_238,In_416);
nand U157 (N_157,In_151,In_859);
xnor U158 (N_158,In_693,In_204);
nand U159 (N_159,In_970,In_612);
xnor U160 (N_160,In_487,In_776);
nand U161 (N_161,In_571,In_361);
nand U162 (N_162,In_369,In_460);
nor U163 (N_163,In_223,In_36);
or U164 (N_164,In_831,In_924);
or U165 (N_165,In_314,In_434);
and U166 (N_166,In_318,In_80);
xnor U167 (N_167,In_40,In_853);
and U168 (N_168,In_214,In_432);
nand U169 (N_169,In_413,In_137);
nand U170 (N_170,In_123,In_181);
nor U171 (N_171,In_77,In_792);
or U172 (N_172,In_66,In_114);
and U173 (N_173,In_483,In_465);
or U174 (N_174,In_676,In_443);
nand U175 (N_175,In_875,In_930);
nand U176 (N_176,In_53,In_838);
nor U177 (N_177,In_672,In_46);
or U178 (N_178,In_176,In_95);
and U179 (N_179,In_264,In_563);
or U180 (N_180,In_251,In_133);
xnor U181 (N_181,In_20,In_542);
or U182 (N_182,In_177,In_865);
or U183 (N_183,In_219,In_328);
and U184 (N_184,In_746,In_496);
nand U185 (N_185,In_439,In_894);
or U186 (N_186,In_726,In_438);
xnor U187 (N_187,In_664,In_382);
or U188 (N_188,In_569,In_762);
and U189 (N_189,In_883,In_575);
nand U190 (N_190,In_28,In_561);
or U191 (N_191,In_922,In_172);
xnor U192 (N_192,In_923,In_104);
nand U193 (N_193,In_365,In_357);
or U194 (N_194,In_524,In_339);
nor U195 (N_195,In_868,In_144);
nand U196 (N_196,In_609,In_422);
or U197 (N_197,In_941,In_689);
and U198 (N_198,In_475,In_709);
and U199 (N_199,In_306,In_653);
nand U200 (N_200,In_279,N_34);
nand U201 (N_201,In_23,In_111);
or U202 (N_202,In_619,In_134);
nand U203 (N_203,In_948,In_937);
or U204 (N_204,N_130,In_806);
and U205 (N_205,In_128,N_102);
or U206 (N_206,In_168,In_869);
or U207 (N_207,In_755,N_115);
nor U208 (N_208,In_24,In_630);
and U209 (N_209,In_331,In_277);
and U210 (N_210,In_820,N_55);
nand U211 (N_211,In_898,In_11);
nor U212 (N_212,In_3,N_98);
nand U213 (N_213,In_886,In_102);
or U214 (N_214,N_88,In_259);
and U215 (N_215,N_155,N_120);
or U216 (N_216,In_774,In_810);
nand U217 (N_217,In_984,In_903);
and U218 (N_218,In_170,In_580);
or U219 (N_219,N_175,In_805);
or U220 (N_220,In_313,In_594);
and U221 (N_221,N_17,In_821);
nor U222 (N_222,In_195,N_62);
or U223 (N_223,In_256,In_716);
nor U224 (N_224,In_482,In_65);
and U225 (N_225,N_190,In_839);
and U226 (N_226,N_144,In_811);
nor U227 (N_227,In_378,In_288);
and U228 (N_228,In_210,In_352);
nor U229 (N_229,In_344,In_671);
xnor U230 (N_230,In_733,In_15);
or U231 (N_231,In_446,In_301);
xnor U232 (N_232,In_493,N_199);
nand U233 (N_233,In_827,N_111);
or U234 (N_234,In_727,In_866);
and U235 (N_235,In_536,N_91);
nand U236 (N_236,N_1,In_435);
and U237 (N_237,N_26,N_140);
and U238 (N_238,In_249,In_411);
nor U239 (N_239,In_127,In_260);
nor U240 (N_240,N_21,In_803);
and U241 (N_241,In_324,N_126);
nand U242 (N_242,N_27,In_535);
and U243 (N_243,In_589,In_476);
nor U244 (N_244,In_974,In_626);
nand U245 (N_245,In_299,In_325);
or U246 (N_246,In_70,N_152);
nand U247 (N_247,In_444,In_799);
xor U248 (N_248,N_57,N_142);
nor U249 (N_249,N_70,In_169);
nor U250 (N_250,In_632,In_962);
xor U251 (N_251,In_720,In_83);
nand U252 (N_252,In_912,In_119);
nand U253 (N_253,In_712,In_891);
and U254 (N_254,In_271,In_753);
or U255 (N_255,In_740,In_698);
nor U256 (N_256,N_41,In_388);
and U257 (N_257,N_122,In_802);
nand U258 (N_258,In_950,In_138);
nor U259 (N_259,In_541,In_94);
nor U260 (N_260,N_149,N_53);
nand U261 (N_261,N_75,In_330);
or U262 (N_262,In_568,In_166);
and U263 (N_263,In_84,In_130);
xor U264 (N_264,In_215,In_768);
and U265 (N_265,In_346,N_89);
nor U266 (N_266,N_176,In_56);
nor U267 (N_267,N_92,In_928);
and U268 (N_268,In_526,In_202);
and U269 (N_269,In_793,In_73);
xnor U270 (N_270,In_101,In_448);
nand U271 (N_271,In_738,N_153);
and U272 (N_272,In_192,In_852);
and U273 (N_273,In_836,N_136);
or U274 (N_274,In_737,N_5);
nor U275 (N_275,In_471,N_133);
nor U276 (N_276,In_916,In_497);
or U277 (N_277,N_112,N_181);
and U278 (N_278,In_599,N_81);
nor U279 (N_279,N_83,In_914);
nor U280 (N_280,In_340,In_415);
nor U281 (N_281,In_817,In_885);
xor U282 (N_282,N_78,In_27);
or U283 (N_283,In_890,In_703);
nand U284 (N_284,N_196,In_503);
xor U285 (N_285,N_97,In_921);
or U286 (N_286,N_170,In_932);
and U287 (N_287,In_22,In_450);
nor U288 (N_288,In_360,N_116);
nand U289 (N_289,N_195,In_78);
nor U290 (N_290,N_174,N_45);
and U291 (N_291,In_744,In_605);
nand U292 (N_292,In_194,In_269);
and U293 (N_293,N_117,In_441);
and U294 (N_294,In_783,In_685);
nand U295 (N_295,N_84,N_86);
or U296 (N_296,In_342,In_75);
and U297 (N_297,In_892,In_453);
xnor U298 (N_298,In_800,In_870);
or U299 (N_299,In_860,In_559);
xor U300 (N_300,N_138,In_608);
nand U301 (N_301,In_332,In_739);
nor U302 (N_302,In_375,In_377);
xor U303 (N_303,In_759,N_159);
nand U304 (N_304,In_583,In_634);
and U305 (N_305,In_777,In_467);
or U306 (N_306,In_464,N_186);
nand U307 (N_307,In_934,In_120);
nor U308 (N_308,In_178,In_280);
and U309 (N_309,In_229,In_801);
nor U310 (N_310,In_254,N_118);
nand U311 (N_311,In_546,In_570);
nor U312 (N_312,N_99,N_163);
nand U313 (N_313,In_145,In_498);
nand U314 (N_314,In_286,In_993);
nor U315 (N_315,In_291,In_500);
nand U316 (N_316,In_642,In_988);
or U317 (N_317,In_523,N_18);
or U318 (N_318,In_402,N_69);
or U319 (N_319,In_410,In_815);
or U320 (N_320,In_48,In_760);
nor U321 (N_321,In_187,N_108);
and U322 (N_322,In_284,In_531);
and U323 (N_323,In_323,In_769);
xor U324 (N_324,In_82,N_182);
and U325 (N_325,In_981,In_673);
or U326 (N_326,N_36,In_688);
nor U327 (N_327,N_54,In_37);
or U328 (N_328,In_241,N_39);
and U329 (N_329,N_147,N_6);
nor U330 (N_330,N_106,In_581);
nor U331 (N_331,In_39,In_926);
nand U332 (N_332,In_735,N_67);
nand U333 (N_333,In_779,In_756);
nand U334 (N_334,In_850,In_418);
nand U335 (N_335,In_864,In_113);
or U336 (N_336,In_245,In_206);
and U337 (N_337,In_350,In_908);
and U338 (N_338,In_492,In_833);
nor U339 (N_339,In_992,In_983);
or U340 (N_340,N_38,In_913);
and U341 (N_341,In_0,In_97);
nand U342 (N_342,In_99,In_690);
or U343 (N_343,In_272,N_37);
nand U344 (N_344,In_751,In_506);
nand U345 (N_345,N_134,N_31);
and U346 (N_346,In_362,In_871);
or U347 (N_347,In_666,In_991);
nor U348 (N_348,N_124,In_822);
nand U349 (N_349,In_639,In_732);
nand U350 (N_350,N_119,In_52);
and U351 (N_351,In_700,In_212);
xnor U352 (N_352,In_491,In_572);
or U353 (N_353,In_674,N_85);
nor U354 (N_354,In_731,In_499);
nand U355 (N_355,In_844,In_440);
xor U356 (N_356,In_32,N_168);
nand U357 (N_357,In_345,In_633);
and U358 (N_358,N_59,In_207);
nand U359 (N_359,In_507,In_761);
nor U360 (N_360,In_409,N_79);
xnor U361 (N_361,In_63,In_851);
or U362 (N_362,N_135,In_353);
xor U363 (N_363,N_184,In_564);
and U364 (N_364,In_76,In_785);
nand U365 (N_365,In_2,In_967);
nand U366 (N_366,In_618,In_677);
and U367 (N_367,In_33,N_46);
xnor U368 (N_368,N_65,In_338);
nand U369 (N_369,In_643,In_433);
xnor U370 (N_370,N_127,In_320);
or U371 (N_371,In_586,In_694);
nand U372 (N_372,N_194,In_363);
xnor U373 (N_373,In_8,N_185);
nand U374 (N_374,In_521,N_48);
nand U375 (N_375,In_931,In_400);
and U376 (N_376,In_232,In_124);
or U377 (N_377,In_979,N_107);
or U378 (N_378,In_947,In_474);
and U379 (N_379,N_110,N_191);
nand U380 (N_380,In_420,In_876);
xnor U381 (N_381,N_2,In_556);
nor U382 (N_382,N_11,In_797);
or U383 (N_383,In_595,In_216);
nor U384 (N_384,N_183,In_278);
and U385 (N_385,In_74,In_647);
xor U386 (N_386,In_843,In_35);
nor U387 (N_387,In_406,In_969);
and U388 (N_388,In_459,In_510);
or U389 (N_389,In_322,In_557);
nand U390 (N_390,In_436,N_50);
nand U391 (N_391,In_585,In_757);
or U392 (N_392,In_734,In_211);
or U393 (N_393,In_227,In_675);
and U394 (N_394,In_551,In_848);
or U395 (N_395,In_163,N_137);
or U396 (N_396,In_329,N_188);
nor U397 (N_397,N_40,In_228);
nand U398 (N_398,In_529,In_379);
or U399 (N_399,N_77,In_505);
nand U400 (N_400,In_651,N_197);
nand U401 (N_401,In_473,N_209);
and U402 (N_402,N_266,In_57);
nand U403 (N_403,N_379,In_14);
and U404 (N_404,N_154,In_190);
nand U405 (N_405,In_193,N_282);
nor U406 (N_406,N_359,N_222);
nor U407 (N_407,In_543,In_995);
and U408 (N_408,In_918,N_43);
nand U409 (N_409,In_706,In_200);
or U410 (N_410,In_403,In_60);
and U411 (N_411,N_229,In_604);
nand U412 (N_412,In_312,N_319);
xnor U413 (N_413,N_391,In_919);
or U414 (N_414,In_684,N_241);
or U415 (N_415,N_93,In_683);
nand U416 (N_416,In_356,N_272);
nand U417 (N_417,N_369,In_383);
nor U418 (N_418,In_118,N_165);
nand U419 (N_419,N_132,N_227);
nand U420 (N_420,In_621,In_659);
nor U421 (N_421,In_771,In_488);
nand U422 (N_422,In_945,N_269);
or U423 (N_423,N_384,N_28);
nor U424 (N_424,In_857,N_245);
or U425 (N_425,In_787,In_248);
and U426 (N_426,N_24,N_247);
nand U427 (N_427,In_788,In_85);
nand U428 (N_428,In_81,N_56);
nor U429 (N_429,In_109,In_58);
or U430 (N_430,N_216,N_210);
nor U431 (N_431,N_273,In_442);
nand U432 (N_432,In_270,N_389);
or U433 (N_433,In_222,N_123);
nor U434 (N_434,N_313,In_183);
nand U435 (N_435,N_299,N_283);
nor U436 (N_436,In_600,N_20);
and U437 (N_437,N_16,N_7);
nor U438 (N_438,N_10,N_330);
or U439 (N_439,In_16,In_9);
nor U440 (N_440,In_31,N_347);
nand U441 (N_441,In_544,In_823);
and U442 (N_442,In_89,N_214);
xor U443 (N_443,In_304,N_345);
or U444 (N_444,In_447,N_254);
nor U445 (N_445,N_87,N_255);
or U446 (N_446,N_315,In_789);
nor U447 (N_447,In_598,N_145);
or U448 (N_448,N_173,N_44);
or U449 (N_449,N_179,In_933);
nand U450 (N_450,In_208,N_52);
nor U451 (N_451,In_479,N_326);
and U452 (N_452,N_259,In_951);
and U453 (N_453,In_562,N_230);
nand U454 (N_454,In_636,N_354);
or U455 (N_455,In_308,In_935);
nor U456 (N_456,N_198,In_226);
nand U457 (N_457,In_401,N_338);
nand U458 (N_458,N_382,N_146);
nand U459 (N_459,N_355,In_722);
or U460 (N_460,In_576,In_990);
xnor U461 (N_461,In_424,N_340);
xnor U462 (N_462,In_404,N_22);
or U463 (N_463,N_335,N_246);
nand U464 (N_464,N_162,N_208);
nor U465 (N_465,N_318,In_707);
nor U466 (N_466,In_687,N_339);
nand U467 (N_467,In_1,In_484);
or U468 (N_468,N_169,N_257);
and U469 (N_469,N_393,N_337);
and U470 (N_470,N_29,In_292);
and U471 (N_471,In_141,In_389);
nand U472 (N_472,N_302,N_160);
nor U473 (N_473,N_213,N_212);
nand U474 (N_474,In_381,In_274);
nand U475 (N_475,In_408,N_156);
nand U476 (N_476,N_343,In_305);
nor U477 (N_477,In_942,In_4);
nor U478 (N_478,In_628,In_641);
or U479 (N_479,N_218,N_248);
nand U480 (N_480,N_289,N_151);
xor U481 (N_481,In_550,N_223);
nor U482 (N_482,In_939,In_43);
nand U483 (N_483,N_13,In_877);
or U484 (N_484,In_142,In_504);
nand U485 (N_485,N_268,In_958);
nor U486 (N_486,N_320,N_220);
xnor U487 (N_487,In_263,N_297);
or U488 (N_488,In_162,In_961);
nor U489 (N_489,N_281,N_178);
nor U490 (N_490,N_94,In_809);
or U491 (N_491,N_15,In_25);
or U492 (N_492,In_326,N_244);
nor U493 (N_493,In_957,N_287);
or U494 (N_494,N_399,In_597);
xnor U495 (N_495,N_357,N_296);
nand U496 (N_496,N_392,N_23);
nand U497 (N_497,N_274,N_217);
nand U498 (N_498,N_306,N_301);
or U499 (N_499,In_188,N_262);
or U500 (N_500,In_873,N_192);
and U501 (N_501,In_611,N_30);
or U502 (N_502,In_741,N_291);
xnor U503 (N_503,N_189,In_199);
or U504 (N_504,In_889,In_514);
and U505 (N_505,N_71,N_279);
nor U506 (N_506,In_348,In_764);
xor U507 (N_507,In_182,In_718);
and U508 (N_508,In_808,N_237);
nor U509 (N_509,N_322,N_386);
xor U510 (N_510,N_51,In_59);
and U511 (N_511,In_538,In_682);
nor U512 (N_512,N_323,In_19);
nor U513 (N_513,In_87,In_692);
nand U514 (N_514,N_284,In_5);
nor U515 (N_515,In_92,N_200);
and U516 (N_516,In_573,N_60);
nand U517 (N_517,N_187,In_93);
nor U518 (N_518,In_518,In_508);
and U519 (N_519,In_273,In_414);
xor U520 (N_520,In_310,N_61);
or U521 (N_521,N_35,In_620);
nand U522 (N_522,N_157,In_711);
nor U523 (N_523,In_915,In_419);
nand U524 (N_524,N_303,N_387);
or U525 (N_525,N_225,N_314);
xnor U526 (N_526,N_271,N_397);
xnor U527 (N_527,In_7,N_113);
or U528 (N_528,In_631,N_381);
or U529 (N_529,In_710,In_998);
and U530 (N_530,In_481,In_509);
or U531 (N_531,N_277,N_288);
nand U532 (N_532,In_217,In_294);
nand U533 (N_533,N_234,N_377);
or U534 (N_534,In_399,N_215);
xnor U535 (N_535,N_105,In_64);
nand U536 (N_536,N_295,In_982);
and U537 (N_537,N_261,In_953);
nand U538 (N_538,N_321,In_160);
or U539 (N_539,N_104,In_480);
nand U540 (N_540,In_55,N_224);
nor U541 (N_541,N_285,In_887);
xnor U542 (N_542,N_150,In_29);
and U543 (N_543,N_292,N_311);
nand U544 (N_544,In_527,N_211);
nor U545 (N_545,In_616,N_240);
and U546 (N_546,In_105,In_985);
or U547 (N_547,N_180,In_627);
and U548 (N_548,In_489,N_239);
nor U549 (N_549,In_874,N_206);
xnor U550 (N_550,In_327,In_374);
nand U551 (N_551,In_804,N_202);
nand U552 (N_552,In_392,In_295);
and U553 (N_553,N_344,In_840);
nor U554 (N_554,In_997,In_398);
nor U555 (N_555,N_324,N_264);
nor U556 (N_556,N_366,In_705);
or U557 (N_557,In_261,In_775);
or U558 (N_558,In_826,In_778);
xnor U559 (N_559,In_90,N_385);
or U560 (N_560,In_638,N_374);
or U561 (N_561,N_109,In_343);
xnor U562 (N_562,N_252,N_331);
nand U563 (N_563,In_517,N_63);
nor U564 (N_564,N_114,N_103);
and U565 (N_565,N_380,N_263);
xnor U566 (N_566,N_376,N_243);
nor U567 (N_567,In_191,N_346);
nand U568 (N_568,N_90,N_0);
nand U569 (N_569,In_230,N_249);
nor U570 (N_570,In_943,N_367);
and U571 (N_571,In_121,N_364);
and U572 (N_572,In_996,N_19);
or U573 (N_573,In_150,N_96);
nand U574 (N_574,In_699,N_143);
or U575 (N_575,N_350,N_342);
nor U576 (N_576,N_276,N_305);
or U577 (N_577,In_582,In_494);
and U578 (N_578,In_856,In_21);
and U579 (N_579,N_228,In_437);
and U580 (N_580,N_32,In_702);
or U581 (N_581,N_4,In_763);
or U582 (N_582,In_337,In_167);
and U583 (N_583,N_9,In_246);
nor U584 (N_584,In_91,In_257);
nor U585 (N_585,N_394,N_207);
nand U586 (N_586,N_14,In_252);
nand U587 (N_587,In_845,N_365);
nand U588 (N_588,N_253,In_854);
nand U589 (N_589,In_458,In_548);
nor U590 (N_590,N_251,N_336);
or U591 (N_591,N_327,In_880);
nand U592 (N_592,N_290,In_911);
and U593 (N_593,N_328,N_298);
nand U594 (N_594,In_445,In_540);
or U595 (N_595,N_221,N_370);
nand U596 (N_596,In_989,In_490);
or U597 (N_597,In_334,N_353);
or U598 (N_598,In_987,N_82);
and U599 (N_599,N_356,In_355);
or U600 (N_600,In_112,N_445);
or U601 (N_601,N_569,N_522);
and U602 (N_602,N_68,N_172);
nand U603 (N_603,N_73,N_493);
nor U604 (N_604,N_158,In_394);
nand U605 (N_605,N_470,N_538);
or U606 (N_606,In_986,N_576);
and U607 (N_607,N_437,N_129);
xnor U608 (N_608,N_378,N_586);
nand U609 (N_609,In_282,In_276);
and U610 (N_610,N_525,N_532);
or U611 (N_611,N_461,N_405);
xor U612 (N_612,N_574,N_242);
and U613 (N_613,N_520,N_372);
nor U614 (N_614,N_448,N_238);
and U615 (N_615,N_420,N_487);
and U616 (N_616,N_164,N_599);
nand U617 (N_617,N_581,N_415);
nand U618 (N_618,In_455,N_100);
xor U619 (N_619,In_185,N_352);
and U620 (N_620,N_8,N_515);
nor U621 (N_621,N_422,N_275);
or U622 (N_622,N_554,N_250);
nor U623 (N_623,In_814,In_615);
nand U624 (N_624,N_465,N_585);
nand U625 (N_625,N_469,N_462);
nor U626 (N_626,In_963,N_390);
or U627 (N_627,N_517,N_267);
and U628 (N_628,N_425,N_543);
or U629 (N_629,N_80,N_358);
or U630 (N_630,N_451,N_76);
and U631 (N_631,In_662,N_499);
nor U632 (N_632,N_598,In_670);
or U633 (N_633,N_429,In_512);
nand U634 (N_634,In_654,N_478);
nand U635 (N_635,N_235,In_736);
nor U636 (N_636,N_395,In_977);
or U637 (N_637,N_233,In_44);
or U638 (N_638,N_505,In_747);
or U639 (N_639,In_157,N_546);
nor U640 (N_640,N_513,N_526);
and U641 (N_641,N_480,N_547);
or U642 (N_642,N_236,N_558);
and U643 (N_643,N_500,In_462);
nor U644 (N_644,N_286,In_899);
xor U645 (N_645,In_574,N_590);
nand U646 (N_646,N_527,N_430);
nand U647 (N_647,N_64,N_441);
nand U648 (N_648,N_432,N_424);
nor U649 (N_649,N_433,N_593);
and U650 (N_650,N_572,N_258);
and U651 (N_651,N_417,N_597);
or U652 (N_652,N_431,In_466);
and U653 (N_653,N_495,N_413);
or U654 (N_654,N_219,N_460);
and U655 (N_655,N_360,N_396);
nand U656 (N_656,In_290,N_583);
xnor U657 (N_657,N_440,In_837);
and U658 (N_658,In_644,In_370);
nor U659 (N_659,N_447,N_491);
and U660 (N_660,N_204,In_122);
nand U661 (N_661,In_812,In_884);
and U662 (N_662,In_146,In_652);
nand U663 (N_663,N_471,In_745);
or U664 (N_664,In_623,N_294);
nor U665 (N_665,N_66,In_714);
and U666 (N_666,N_479,In_153);
nand U667 (N_667,N_439,N_456);
nand U668 (N_668,N_457,N_524);
and U669 (N_669,In_952,N_125);
nor U670 (N_670,In_367,N_121);
and U671 (N_671,N_412,N_473);
nand U672 (N_672,N_485,N_72);
or U673 (N_673,N_551,N_595);
and U674 (N_674,N_231,In_790);
nor U675 (N_675,In_946,N_193);
nand U676 (N_676,N_349,N_587);
nand U677 (N_677,In_502,N_427);
xnor U678 (N_678,N_428,N_332);
and U679 (N_679,N_573,N_363);
xnor U680 (N_680,N_549,N_452);
or U681 (N_681,In_116,N_12);
or U682 (N_682,In_298,N_278);
or U683 (N_683,N_453,N_270);
nor U684 (N_684,In_461,In_579);
or U685 (N_685,N_203,In_265);
nand U686 (N_686,N_423,In_661);
and U687 (N_687,In_954,N_406);
and U688 (N_688,N_421,N_438);
or U689 (N_689,N_444,N_171);
nor U690 (N_690,N_541,N_476);
and U691 (N_691,N_404,N_463);
and U692 (N_692,N_566,In_648);
nor U693 (N_693,N_362,In_849);
nor U694 (N_694,N_410,N_443);
or U695 (N_695,In_578,N_166);
nor U696 (N_696,N_531,In_253);
xnor U697 (N_697,N_398,N_466);
nor U698 (N_698,In_449,In_47);
nor U699 (N_699,N_161,In_262);
and U700 (N_700,N_486,In_457);
xor U701 (N_701,In_472,N_455);
or U702 (N_702,N_101,N_474);
and U703 (N_703,N_502,N_512);
nor U704 (N_704,In_553,N_33);
and U705 (N_705,In_61,N_435);
nand U706 (N_706,N_307,N_594);
xnor U707 (N_707,In_695,N_260);
and U708 (N_708,In_818,N_131);
and U709 (N_709,N_436,N_167);
nor U710 (N_710,N_459,N_563);
or U711 (N_711,N_506,N_42);
nand U712 (N_712,N_300,N_401);
or U713 (N_713,In_596,N_361);
and U714 (N_714,N_310,N_511);
and U715 (N_715,N_567,N_559);
nand U716 (N_716,N_494,N_434);
nand U717 (N_717,N_582,N_141);
or U718 (N_718,In_717,In_106);
or U719 (N_719,N_498,N_148);
or U720 (N_720,In_830,N_552);
or U721 (N_721,N_312,N_539);
xor U722 (N_722,N_484,N_467);
nand U723 (N_723,N_536,N_596);
nor U724 (N_724,N_368,In_773);
and U725 (N_725,In_525,N_458);
and U726 (N_726,In_668,N_523);
and U727 (N_727,N_373,In_244);
xor U728 (N_728,N_293,N_577);
nand U729 (N_729,N_490,N_177);
nand U730 (N_730,N_521,N_309);
and U731 (N_731,N_333,N_589);
and U732 (N_732,N_308,N_557);
nand U733 (N_733,N_492,N_426);
and U734 (N_734,N_496,N_508);
nor U735 (N_735,N_442,In_528);
nor U736 (N_736,N_483,N_58);
nand U737 (N_737,In_126,N_529);
nand U738 (N_738,N_555,N_482);
nand U739 (N_739,N_501,N_416);
nand U740 (N_740,In_218,N_450);
and U741 (N_741,N_419,N_516);
nor U742 (N_742,In_530,N_418);
or U743 (N_743,N_304,N_568);
nand U744 (N_744,N_226,N_560);
nor U745 (N_745,N_265,In_645);
or U746 (N_746,N_280,N_348);
or U747 (N_747,N_316,N_139);
nor U748 (N_748,N_475,N_407);
and U749 (N_749,N_561,N_556);
nand U750 (N_750,N_472,N_530);
or U751 (N_751,N_548,N_383);
nor U752 (N_752,N_497,N_400);
nor U753 (N_753,N_550,N_388);
or U754 (N_754,N_571,In_486);
nand U755 (N_755,In_715,N_519);
nor U756 (N_756,N_553,N_95);
xnor U757 (N_757,N_503,N_3);
nand U758 (N_758,In_275,N_518);
or U759 (N_759,N_446,N_351);
nand U760 (N_760,In_592,N_481);
nand U761 (N_761,N_584,N_545);
nand U762 (N_762,N_489,In_395);
and U763 (N_763,N_564,In_881);
or U764 (N_764,N_580,N_540);
or U765 (N_765,In_758,N_371);
nor U766 (N_766,N_454,N_317);
or U767 (N_767,N_409,N_528);
nor U768 (N_768,N_579,N_449);
nand U769 (N_769,N_468,In_904);
xnor U770 (N_770,N_535,N_488);
nand U771 (N_771,N_588,In_149);
nand U772 (N_772,N_575,N_341);
or U773 (N_773,N_534,N_570);
or U774 (N_774,In_896,N_375);
or U775 (N_775,N_477,In_927);
nor U776 (N_776,In_319,In_68);
and U777 (N_777,N_411,N_542);
and U778 (N_778,In_558,N_562);
nand U779 (N_779,N_256,N_49);
and U780 (N_780,N_504,N_25);
nor U781 (N_781,N_408,N_74);
nand U782 (N_782,N_507,N_402);
nor U783 (N_783,In_577,N_464);
and U784 (N_784,N_403,N_591);
and U785 (N_785,N_544,N_578);
or U786 (N_786,In_470,N_514);
nand U787 (N_787,N_509,In_243);
nand U788 (N_788,In_938,N_232);
and U789 (N_789,In_770,In_110);
or U790 (N_790,In_766,N_334);
and U791 (N_791,N_201,In_240);
and U792 (N_792,N_533,In_423);
or U793 (N_793,N_414,N_325);
and U794 (N_794,N_592,In_565);
or U795 (N_795,N_47,In_289);
xor U796 (N_796,N_537,N_205);
nor U797 (N_797,In_534,N_329);
xnor U798 (N_798,N_128,N_510);
nand U799 (N_799,N_565,In_372);
nor U800 (N_800,N_688,N_629);
or U801 (N_801,N_611,N_753);
nor U802 (N_802,N_699,N_706);
or U803 (N_803,N_681,N_683);
nor U804 (N_804,N_632,N_695);
nor U805 (N_805,N_672,N_797);
nor U806 (N_806,N_731,N_679);
nand U807 (N_807,N_690,N_618);
or U808 (N_808,N_612,N_643);
and U809 (N_809,N_741,N_658);
or U810 (N_810,N_662,N_669);
nor U811 (N_811,N_746,N_694);
nor U812 (N_812,N_736,N_635);
nor U813 (N_813,N_607,N_602);
and U814 (N_814,N_640,N_685);
or U815 (N_815,N_762,N_682);
xnor U816 (N_816,N_704,N_772);
nor U817 (N_817,N_677,N_754);
nor U818 (N_818,N_768,N_633);
nand U819 (N_819,N_788,N_614);
nor U820 (N_820,N_723,N_654);
xnor U821 (N_821,N_705,N_744);
nor U822 (N_822,N_742,N_789);
or U823 (N_823,N_661,N_714);
nand U824 (N_824,N_752,N_710);
nand U825 (N_825,N_657,N_739);
or U826 (N_826,N_738,N_622);
nor U827 (N_827,N_783,N_769);
or U828 (N_828,N_606,N_724);
nand U829 (N_829,N_634,N_794);
or U830 (N_830,N_638,N_605);
nor U831 (N_831,N_758,N_743);
or U832 (N_832,N_718,N_603);
xor U833 (N_833,N_767,N_787);
nor U834 (N_834,N_627,N_616);
nor U835 (N_835,N_621,N_792);
nor U836 (N_836,N_798,N_747);
nand U837 (N_837,N_760,N_697);
nor U838 (N_838,N_755,N_732);
and U839 (N_839,N_692,N_790);
nand U840 (N_840,N_701,N_795);
or U841 (N_841,N_650,N_676);
or U842 (N_842,N_785,N_703);
nand U843 (N_843,N_784,N_648);
or U844 (N_844,N_719,N_680);
nor U845 (N_845,N_759,N_749);
nand U846 (N_846,N_781,N_615);
and U847 (N_847,N_745,N_619);
nand U848 (N_848,N_660,N_637);
nand U849 (N_849,N_691,N_735);
xor U850 (N_850,N_601,N_678);
nand U851 (N_851,N_709,N_748);
nand U852 (N_852,N_720,N_791);
and U853 (N_853,N_675,N_777);
nand U854 (N_854,N_712,N_771);
and U855 (N_855,N_740,N_670);
nand U856 (N_856,N_655,N_793);
and U857 (N_857,N_668,N_666);
nor U858 (N_858,N_716,N_763);
xnor U859 (N_859,N_689,N_631);
nor U860 (N_860,N_715,N_673);
nand U861 (N_861,N_778,N_707);
and U862 (N_862,N_725,N_761);
and U863 (N_863,N_617,N_737);
and U864 (N_864,N_729,N_713);
nand U865 (N_865,N_757,N_649);
and U866 (N_866,N_647,N_604);
xnor U867 (N_867,N_652,N_799);
nand U868 (N_868,N_733,N_646);
or U869 (N_869,N_645,N_727);
xor U870 (N_870,N_651,N_628);
nor U871 (N_871,N_779,N_696);
nor U872 (N_872,N_613,N_730);
nor U873 (N_873,N_653,N_711);
or U874 (N_874,N_667,N_734);
nor U875 (N_875,N_756,N_600);
nor U876 (N_876,N_774,N_620);
nor U877 (N_877,N_770,N_722);
nand U878 (N_878,N_610,N_636);
nor U879 (N_879,N_693,N_674);
or U880 (N_880,N_644,N_624);
and U881 (N_881,N_642,N_765);
nand U882 (N_882,N_702,N_626);
nand U883 (N_883,N_623,N_728);
or U884 (N_884,N_721,N_750);
nand U885 (N_885,N_609,N_641);
or U886 (N_886,N_684,N_665);
and U887 (N_887,N_708,N_687);
or U888 (N_888,N_782,N_700);
xnor U889 (N_889,N_608,N_764);
nand U890 (N_890,N_775,N_656);
nor U891 (N_891,N_786,N_671);
nand U892 (N_892,N_766,N_659);
nand U893 (N_893,N_686,N_751);
or U894 (N_894,N_773,N_780);
nand U895 (N_895,N_698,N_664);
nand U896 (N_896,N_726,N_625);
or U897 (N_897,N_796,N_630);
nand U898 (N_898,N_663,N_639);
or U899 (N_899,N_776,N_717);
nand U900 (N_900,N_766,N_785);
or U901 (N_901,N_698,N_633);
or U902 (N_902,N_777,N_788);
nor U903 (N_903,N_789,N_733);
or U904 (N_904,N_760,N_607);
nand U905 (N_905,N_793,N_799);
nand U906 (N_906,N_707,N_680);
and U907 (N_907,N_615,N_792);
or U908 (N_908,N_771,N_794);
nor U909 (N_909,N_796,N_751);
or U910 (N_910,N_664,N_791);
nor U911 (N_911,N_676,N_738);
or U912 (N_912,N_780,N_610);
and U913 (N_913,N_792,N_761);
nor U914 (N_914,N_750,N_636);
and U915 (N_915,N_618,N_673);
or U916 (N_916,N_738,N_624);
or U917 (N_917,N_658,N_738);
nand U918 (N_918,N_751,N_649);
xor U919 (N_919,N_724,N_744);
nand U920 (N_920,N_751,N_643);
xnor U921 (N_921,N_764,N_781);
and U922 (N_922,N_693,N_606);
or U923 (N_923,N_612,N_720);
nand U924 (N_924,N_657,N_772);
nand U925 (N_925,N_774,N_646);
nand U926 (N_926,N_726,N_747);
nor U927 (N_927,N_619,N_687);
or U928 (N_928,N_779,N_796);
and U929 (N_929,N_612,N_629);
nor U930 (N_930,N_750,N_743);
and U931 (N_931,N_727,N_610);
nand U932 (N_932,N_624,N_630);
or U933 (N_933,N_746,N_712);
xor U934 (N_934,N_738,N_604);
and U935 (N_935,N_677,N_799);
nand U936 (N_936,N_718,N_671);
and U937 (N_937,N_663,N_779);
nand U938 (N_938,N_707,N_672);
nand U939 (N_939,N_635,N_772);
nor U940 (N_940,N_745,N_776);
and U941 (N_941,N_772,N_600);
and U942 (N_942,N_706,N_638);
and U943 (N_943,N_676,N_698);
nor U944 (N_944,N_772,N_617);
or U945 (N_945,N_644,N_664);
or U946 (N_946,N_724,N_774);
or U947 (N_947,N_686,N_684);
or U948 (N_948,N_611,N_659);
nand U949 (N_949,N_749,N_692);
nor U950 (N_950,N_684,N_751);
xnor U951 (N_951,N_623,N_742);
nor U952 (N_952,N_611,N_689);
and U953 (N_953,N_633,N_702);
xor U954 (N_954,N_651,N_726);
nor U955 (N_955,N_658,N_606);
nand U956 (N_956,N_760,N_666);
or U957 (N_957,N_776,N_719);
and U958 (N_958,N_789,N_787);
nand U959 (N_959,N_678,N_609);
or U960 (N_960,N_795,N_749);
and U961 (N_961,N_693,N_735);
and U962 (N_962,N_680,N_764);
or U963 (N_963,N_757,N_612);
nand U964 (N_964,N_664,N_753);
and U965 (N_965,N_780,N_729);
nand U966 (N_966,N_631,N_695);
nor U967 (N_967,N_773,N_752);
and U968 (N_968,N_612,N_754);
or U969 (N_969,N_745,N_644);
or U970 (N_970,N_764,N_753);
and U971 (N_971,N_603,N_707);
nor U972 (N_972,N_753,N_698);
or U973 (N_973,N_631,N_753);
nor U974 (N_974,N_789,N_628);
and U975 (N_975,N_642,N_654);
or U976 (N_976,N_781,N_772);
nor U977 (N_977,N_772,N_770);
and U978 (N_978,N_639,N_786);
nand U979 (N_979,N_795,N_620);
xor U980 (N_980,N_793,N_620);
and U981 (N_981,N_652,N_720);
nor U982 (N_982,N_704,N_690);
or U983 (N_983,N_693,N_720);
and U984 (N_984,N_659,N_705);
or U985 (N_985,N_634,N_758);
nor U986 (N_986,N_667,N_626);
and U987 (N_987,N_696,N_706);
and U988 (N_988,N_670,N_696);
xnor U989 (N_989,N_626,N_623);
or U990 (N_990,N_757,N_711);
and U991 (N_991,N_725,N_704);
nor U992 (N_992,N_661,N_609);
or U993 (N_993,N_762,N_680);
xnor U994 (N_994,N_781,N_774);
or U995 (N_995,N_621,N_628);
or U996 (N_996,N_717,N_755);
nand U997 (N_997,N_705,N_751);
xnor U998 (N_998,N_648,N_681);
and U999 (N_999,N_605,N_670);
or U1000 (N_1000,N_971,N_826);
nor U1001 (N_1001,N_885,N_848);
and U1002 (N_1002,N_858,N_898);
or U1003 (N_1003,N_820,N_925);
and U1004 (N_1004,N_903,N_956);
nand U1005 (N_1005,N_837,N_976);
or U1006 (N_1006,N_849,N_984);
and U1007 (N_1007,N_827,N_910);
and U1008 (N_1008,N_933,N_936);
nor U1009 (N_1009,N_899,N_831);
nor U1010 (N_1010,N_913,N_891);
xor U1011 (N_1011,N_901,N_962);
or U1012 (N_1012,N_834,N_996);
and U1013 (N_1013,N_875,N_959);
and U1014 (N_1014,N_836,N_992);
nor U1015 (N_1015,N_816,N_921);
xnor U1016 (N_1016,N_987,N_886);
and U1017 (N_1017,N_947,N_884);
nand U1018 (N_1018,N_985,N_894);
nor U1019 (N_1019,N_988,N_832);
nand U1020 (N_1020,N_995,N_920);
or U1021 (N_1021,N_852,N_945);
and U1022 (N_1022,N_845,N_978);
nand U1023 (N_1023,N_991,N_912);
or U1024 (N_1024,N_919,N_879);
and U1025 (N_1025,N_941,N_895);
nand U1026 (N_1026,N_954,N_949);
nand U1027 (N_1027,N_844,N_865);
nor U1028 (N_1028,N_951,N_969);
or U1029 (N_1029,N_887,N_839);
nor U1030 (N_1030,N_923,N_904);
and U1031 (N_1031,N_840,N_808);
or U1032 (N_1032,N_915,N_909);
or U1033 (N_1033,N_952,N_880);
nand U1034 (N_1034,N_935,N_868);
nor U1035 (N_1035,N_950,N_893);
nand U1036 (N_1036,N_997,N_859);
or U1037 (N_1037,N_938,N_857);
nor U1038 (N_1038,N_823,N_841);
nand U1039 (N_1039,N_866,N_994);
and U1040 (N_1040,N_967,N_943);
xnor U1041 (N_1041,N_811,N_964);
or U1042 (N_1042,N_932,N_908);
nor U1043 (N_1043,N_902,N_800);
nand U1044 (N_1044,N_927,N_854);
nor U1045 (N_1045,N_860,N_888);
nor U1046 (N_1046,N_804,N_822);
nand U1047 (N_1047,N_813,N_977);
and U1048 (N_1048,N_917,N_983);
nand U1049 (N_1049,N_892,N_851);
xnor U1050 (N_1050,N_944,N_924);
xnor U1051 (N_1051,N_821,N_825);
and U1052 (N_1052,N_957,N_855);
nand U1053 (N_1053,N_807,N_883);
and U1054 (N_1054,N_981,N_905);
nor U1055 (N_1055,N_877,N_801);
nand U1056 (N_1056,N_942,N_802);
nand U1057 (N_1057,N_930,N_937);
xor U1058 (N_1058,N_968,N_872);
xor U1059 (N_1059,N_934,N_989);
nand U1060 (N_1060,N_843,N_970);
nand U1061 (N_1061,N_830,N_846);
nand U1062 (N_1062,N_805,N_907);
and U1063 (N_1063,N_931,N_874);
nor U1064 (N_1064,N_958,N_817);
or U1065 (N_1065,N_815,N_955);
and U1066 (N_1066,N_914,N_916);
nand U1067 (N_1067,N_828,N_850);
or U1068 (N_1068,N_960,N_838);
and U1069 (N_1069,N_812,N_890);
xor U1070 (N_1070,N_922,N_806);
and U1071 (N_1071,N_829,N_900);
and U1072 (N_1072,N_870,N_990);
xor U1073 (N_1073,N_966,N_972);
nor U1074 (N_1074,N_819,N_999);
and U1075 (N_1075,N_869,N_835);
xor U1076 (N_1076,N_864,N_876);
and U1077 (N_1077,N_998,N_939);
and U1078 (N_1078,N_881,N_906);
nand U1079 (N_1079,N_929,N_963);
or U1080 (N_1080,N_982,N_861);
or U1081 (N_1081,N_975,N_979);
nand U1082 (N_1082,N_833,N_842);
and U1083 (N_1083,N_948,N_856);
nand U1084 (N_1084,N_911,N_862);
nor U1085 (N_1085,N_889,N_873);
or U1086 (N_1086,N_803,N_878);
nand U1087 (N_1087,N_973,N_897);
xnor U1088 (N_1088,N_814,N_993);
xor U1089 (N_1089,N_961,N_810);
nand U1090 (N_1090,N_863,N_928);
nand U1091 (N_1091,N_824,N_946);
nand U1092 (N_1092,N_871,N_974);
or U1093 (N_1093,N_986,N_896);
xnor U1094 (N_1094,N_940,N_853);
or U1095 (N_1095,N_965,N_867);
and U1096 (N_1096,N_847,N_918);
nor U1097 (N_1097,N_953,N_926);
and U1098 (N_1098,N_882,N_980);
or U1099 (N_1099,N_818,N_809);
nand U1100 (N_1100,N_900,N_920);
and U1101 (N_1101,N_866,N_903);
or U1102 (N_1102,N_981,N_889);
nand U1103 (N_1103,N_919,N_923);
or U1104 (N_1104,N_958,N_952);
nand U1105 (N_1105,N_991,N_860);
and U1106 (N_1106,N_904,N_847);
nand U1107 (N_1107,N_958,N_883);
nor U1108 (N_1108,N_884,N_971);
xor U1109 (N_1109,N_866,N_882);
and U1110 (N_1110,N_903,N_825);
nor U1111 (N_1111,N_834,N_911);
nand U1112 (N_1112,N_876,N_857);
nor U1113 (N_1113,N_880,N_858);
nand U1114 (N_1114,N_875,N_921);
or U1115 (N_1115,N_856,N_812);
nand U1116 (N_1116,N_963,N_961);
and U1117 (N_1117,N_822,N_936);
or U1118 (N_1118,N_942,N_800);
nor U1119 (N_1119,N_817,N_996);
nor U1120 (N_1120,N_869,N_935);
xor U1121 (N_1121,N_844,N_963);
nor U1122 (N_1122,N_858,N_804);
nand U1123 (N_1123,N_820,N_997);
xor U1124 (N_1124,N_994,N_992);
and U1125 (N_1125,N_928,N_986);
or U1126 (N_1126,N_966,N_953);
and U1127 (N_1127,N_955,N_910);
and U1128 (N_1128,N_819,N_885);
and U1129 (N_1129,N_993,N_855);
and U1130 (N_1130,N_906,N_993);
xnor U1131 (N_1131,N_876,N_964);
nand U1132 (N_1132,N_921,N_969);
nand U1133 (N_1133,N_995,N_817);
and U1134 (N_1134,N_887,N_824);
nand U1135 (N_1135,N_845,N_976);
or U1136 (N_1136,N_951,N_828);
and U1137 (N_1137,N_987,N_838);
and U1138 (N_1138,N_899,N_930);
nand U1139 (N_1139,N_904,N_931);
nand U1140 (N_1140,N_934,N_880);
nor U1141 (N_1141,N_966,N_861);
nand U1142 (N_1142,N_868,N_931);
or U1143 (N_1143,N_844,N_979);
and U1144 (N_1144,N_948,N_803);
and U1145 (N_1145,N_898,N_907);
and U1146 (N_1146,N_925,N_995);
and U1147 (N_1147,N_828,N_970);
nand U1148 (N_1148,N_856,N_912);
and U1149 (N_1149,N_840,N_908);
nor U1150 (N_1150,N_854,N_839);
or U1151 (N_1151,N_803,N_890);
nand U1152 (N_1152,N_854,N_902);
nor U1153 (N_1153,N_891,N_903);
nor U1154 (N_1154,N_814,N_922);
and U1155 (N_1155,N_966,N_896);
nand U1156 (N_1156,N_804,N_845);
xor U1157 (N_1157,N_833,N_809);
and U1158 (N_1158,N_971,N_876);
and U1159 (N_1159,N_951,N_820);
or U1160 (N_1160,N_820,N_838);
nor U1161 (N_1161,N_830,N_849);
xor U1162 (N_1162,N_969,N_893);
and U1163 (N_1163,N_821,N_813);
and U1164 (N_1164,N_880,N_956);
nor U1165 (N_1165,N_913,N_976);
and U1166 (N_1166,N_880,N_885);
or U1167 (N_1167,N_886,N_855);
nand U1168 (N_1168,N_815,N_883);
nor U1169 (N_1169,N_964,N_842);
and U1170 (N_1170,N_933,N_919);
nor U1171 (N_1171,N_990,N_841);
and U1172 (N_1172,N_818,N_825);
nor U1173 (N_1173,N_879,N_906);
and U1174 (N_1174,N_813,N_906);
or U1175 (N_1175,N_937,N_894);
nor U1176 (N_1176,N_861,N_900);
and U1177 (N_1177,N_940,N_972);
and U1178 (N_1178,N_971,N_877);
and U1179 (N_1179,N_812,N_953);
nor U1180 (N_1180,N_897,N_867);
or U1181 (N_1181,N_976,N_973);
nand U1182 (N_1182,N_935,N_949);
nor U1183 (N_1183,N_990,N_838);
and U1184 (N_1184,N_814,N_837);
or U1185 (N_1185,N_854,N_938);
and U1186 (N_1186,N_854,N_910);
nand U1187 (N_1187,N_974,N_973);
and U1188 (N_1188,N_944,N_915);
nand U1189 (N_1189,N_897,N_938);
xor U1190 (N_1190,N_800,N_890);
nor U1191 (N_1191,N_936,N_810);
nor U1192 (N_1192,N_999,N_984);
or U1193 (N_1193,N_852,N_919);
and U1194 (N_1194,N_873,N_923);
or U1195 (N_1195,N_953,N_894);
nand U1196 (N_1196,N_800,N_925);
nor U1197 (N_1197,N_982,N_862);
and U1198 (N_1198,N_951,N_940);
xor U1199 (N_1199,N_848,N_947);
and U1200 (N_1200,N_1067,N_1132);
or U1201 (N_1201,N_1052,N_1019);
and U1202 (N_1202,N_1042,N_1073);
nand U1203 (N_1203,N_1030,N_1010);
nand U1204 (N_1204,N_1155,N_1154);
nor U1205 (N_1205,N_1021,N_1151);
or U1206 (N_1206,N_1059,N_1036);
nor U1207 (N_1207,N_1029,N_1153);
and U1208 (N_1208,N_1011,N_1003);
nand U1209 (N_1209,N_1148,N_1039);
or U1210 (N_1210,N_1183,N_1034);
and U1211 (N_1211,N_1186,N_1123);
and U1212 (N_1212,N_1165,N_1041);
and U1213 (N_1213,N_1138,N_1009);
nor U1214 (N_1214,N_1134,N_1054);
and U1215 (N_1215,N_1127,N_1187);
or U1216 (N_1216,N_1157,N_1178);
or U1217 (N_1217,N_1121,N_1177);
or U1218 (N_1218,N_1096,N_1063);
xnor U1219 (N_1219,N_1159,N_1184);
and U1220 (N_1220,N_1000,N_1026);
or U1221 (N_1221,N_1158,N_1008);
and U1222 (N_1222,N_1197,N_1195);
and U1223 (N_1223,N_1180,N_1025);
nand U1224 (N_1224,N_1128,N_1112);
and U1225 (N_1225,N_1002,N_1005);
or U1226 (N_1226,N_1049,N_1056);
and U1227 (N_1227,N_1001,N_1190);
xor U1228 (N_1228,N_1028,N_1131);
nand U1229 (N_1229,N_1044,N_1004);
or U1230 (N_1230,N_1174,N_1020);
xnor U1231 (N_1231,N_1164,N_1137);
or U1232 (N_1232,N_1014,N_1037);
nor U1233 (N_1233,N_1161,N_1104);
or U1234 (N_1234,N_1198,N_1140);
or U1235 (N_1235,N_1007,N_1182);
nor U1236 (N_1236,N_1080,N_1070);
or U1237 (N_1237,N_1167,N_1109);
xnor U1238 (N_1238,N_1160,N_1101);
nor U1239 (N_1239,N_1102,N_1013);
nor U1240 (N_1240,N_1051,N_1126);
nor U1241 (N_1241,N_1156,N_1094);
nor U1242 (N_1242,N_1193,N_1032);
nand U1243 (N_1243,N_1108,N_1199);
or U1244 (N_1244,N_1168,N_1081);
nor U1245 (N_1245,N_1117,N_1045);
and U1246 (N_1246,N_1082,N_1103);
and U1247 (N_1247,N_1083,N_1194);
or U1248 (N_1248,N_1120,N_1087);
nand U1249 (N_1249,N_1053,N_1139);
or U1250 (N_1250,N_1068,N_1040);
nor U1251 (N_1251,N_1192,N_1012);
xor U1252 (N_1252,N_1097,N_1050);
and U1253 (N_1253,N_1114,N_1122);
nor U1254 (N_1254,N_1033,N_1110);
nand U1255 (N_1255,N_1107,N_1118);
nor U1256 (N_1256,N_1043,N_1149);
or U1257 (N_1257,N_1055,N_1006);
and U1258 (N_1258,N_1060,N_1115);
nand U1259 (N_1259,N_1035,N_1062);
nor U1260 (N_1260,N_1058,N_1099);
xor U1261 (N_1261,N_1088,N_1038);
and U1262 (N_1262,N_1146,N_1173);
nor U1263 (N_1263,N_1077,N_1119);
nand U1264 (N_1264,N_1022,N_1085);
nor U1265 (N_1265,N_1057,N_1172);
and U1266 (N_1266,N_1130,N_1106);
nor U1267 (N_1267,N_1191,N_1144);
nor U1268 (N_1268,N_1145,N_1024);
or U1269 (N_1269,N_1046,N_1162);
nand U1270 (N_1270,N_1179,N_1092);
and U1271 (N_1271,N_1015,N_1072);
nand U1272 (N_1272,N_1074,N_1089);
nand U1273 (N_1273,N_1018,N_1091);
nor U1274 (N_1274,N_1176,N_1129);
or U1275 (N_1275,N_1076,N_1185);
nor U1276 (N_1276,N_1031,N_1133);
nand U1277 (N_1277,N_1066,N_1152);
or U1278 (N_1278,N_1111,N_1065);
nor U1279 (N_1279,N_1023,N_1163);
nor U1280 (N_1280,N_1116,N_1095);
or U1281 (N_1281,N_1086,N_1135);
and U1282 (N_1282,N_1071,N_1027);
nand U1283 (N_1283,N_1017,N_1189);
or U1284 (N_1284,N_1175,N_1143);
nand U1285 (N_1285,N_1125,N_1064);
or U1286 (N_1286,N_1113,N_1169);
and U1287 (N_1287,N_1150,N_1048);
nor U1288 (N_1288,N_1196,N_1141);
xor U1289 (N_1289,N_1100,N_1090);
nor U1290 (N_1290,N_1016,N_1188);
nand U1291 (N_1291,N_1181,N_1069);
xor U1292 (N_1292,N_1075,N_1078);
nor U1293 (N_1293,N_1142,N_1105);
nor U1294 (N_1294,N_1147,N_1061);
and U1295 (N_1295,N_1136,N_1047);
nor U1296 (N_1296,N_1093,N_1170);
and U1297 (N_1297,N_1084,N_1124);
nor U1298 (N_1298,N_1098,N_1079);
nand U1299 (N_1299,N_1171,N_1166);
xnor U1300 (N_1300,N_1081,N_1084);
xnor U1301 (N_1301,N_1030,N_1027);
nand U1302 (N_1302,N_1035,N_1036);
nor U1303 (N_1303,N_1012,N_1036);
or U1304 (N_1304,N_1131,N_1132);
or U1305 (N_1305,N_1175,N_1150);
or U1306 (N_1306,N_1108,N_1197);
and U1307 (N_1307,N_1198,N_1000);
nor U1308 (N_1308,N_1068,N_1015);
nand U1309 (N_1309,N_1032,N_1030);
nor U1310 (N_1310,N_1029,N_1034);
nand U1311 (N_1311,N_1054,N_1172);
or U1312 (N_1312,N_1190,N_1097);
or U1313 (N_1313,N_1082,N_1097);
nor U1314 (N_1314,N_1047,N_1089);
and U1315 (N_1315,N_1126,N_1017);
or U1316 (N_1316,N_1089,N_1030);
and U1317 (N_1317,N_1174,N_1024);
nor U1318 (N_1318,N_1167,N_1013);
or U1319 (N_1319,N_1092,N_1094);
nor U1320 (N_1320,N_1146,N_1044);
or U1321 (N_1321,N_1130,N_1076);
and U1322 (N_1322,N_1016,N_1084);
nand U1323 (N_1323,N_1106,N_1043);
nor U1324 (N_1324,N_1140,N_1040);
xnor U1325 (N_1325,N_1186,N_1070);
and U1326 (N_1326,N_1174,N_1064);
and U1327 (N_1327,N_1009,N_1159);
nor U1328 (N_1328,N_1141,N_1082);
nand U1329 (N_1329,N_1139,N_1061);
nor U1330 (N_1330,N_1108,N_1044);
nand U1331 (N_1331,N_1019,N_1167);
and U1332 (N_1332,N_1056,N_1079);
nand U1333 (N_1333,N_1135,N_1134);
nor U1334 (N_1334,N_1051,N_1145);
or U1335 (N_1335,N_1056,N_1083);
nor U1336 (N_1336,N_1017,N_1123);
nand U1337 (N_1337,N_1181,N_1129);
nand U1338 (N_1338,N_1050,N_1156);
nand U1339 (N_1339,N_1140,N_1102);
nand U1340 (N_1340,N_1168,N_1051);
and U1341 (N_1341,N_1125,N_1111);
nor U1342 (N_1342,N_1071,N_1001);
and U1343 (N_1343,N_1131,N_1179);
and U1344 (N_1344,N_1022,N_1139);
nand U1345 (N_1345,N_1057,N_1038);
or U1346 (N_1346,N_1144,N_1091);
nor U1347 (N_1347,N_1177,N_1012);
nor U1348 (N_1348,N_1147,N_1138);
and U1349 (N_1349,N_1128,N_1016);
or U1350 (N_1350,N_1122,N_1116);
and U1351 (N_1351,N_1126,N_1043);
nor U1352 (N_1352,N_1168,N_1014);
nand U1353 (N_1353,N_1155,N_1005);
nor U1354 (N_1354,N_1074,N_1022);
xnor U1355 (N_1355,N_1005,N_1041);
or U1356 (N_1356,N_1064,N_1040);
nor U1357 (N_1357,N_1033,N_1003);
or U1358 (N_1358,N_1168,N_1045);
nor U1359 (N_1359,N_1106,N_1173);
nor U1360 (N_1360,N_1137,N_1065);
and U1361 (N_1361,N_1029,N_1126);
nand U1362 (N_1362,N_1132,N_1081);
nand U1363 (N_1363,N_1079,N_1077);
and U1364 (N_1364,N_1035,N_1086);
and U1365 (N_1365,N_1118,N_1187);
and U1366 (N_1366,N_1194,N_1097);
nand U1367 (N_1367,N_1006,N_1029);
and U1368 (N_1368,N_1149,N_1112);
nand U1369 (N_1369,N_1181,N_1051);
and U1370 (N_1370,N_1008,N_1027);
nand U1371 (N_1371,N_1156,N_1140);
nand U1372 (N_1372,N_1145,N_1018);
nor U1373 (N_1373,N_1107,N_1135);
nand U1374 (N_1374,N_1053,N_1095);
nor U1375 (N_1375,N_1013,N_1070);
and U1376 (N_1376,N_1058,N_1160);
and U1377 (N_1377,N_1071,N_1149);
nand U1378 (N_1378,N_1050,N_1145);
or U1379 (N_1379,N_1015,N_1190);
nand U1380 (N_1380,N_1152,N_1120);
nor U1381 (N_1381,N_1087,N_1165);
or U1382 (N_1382,N_1080,N_1092);
nand U1383 (N_1383,N_1111,N_1177);
nand U1384 (N_1384,N_1171,N_1108);
nand U1385 (N_1385,N_1122,N_1038);
nand U1386 (N_1386,N_1136,N_1137);
nand U1387 (N_1387,N_1130,N_1160);
and U1388 (N_1388,N_1165,N_1099);
xnor U1389 (N_1389,N_1057,N_1176);
nor U1390 (N_1390,N_1193,N_1033);
nand U1391 (N_1391,N_1170,N_1140);
nand U1392 (N_1392,N_1052,N_1196);
nand U1393 (N_1393,N_1074,N_1030);
and U1394 (N_1394,N_1030,N_1107);
nor U1395 (N_1395,N_1167,N_1056);
or U1396 (N_1396,N_1150,N_1061);
nand U1397 (N_1397,N_1159,N_1127);
nor U1398 (N_1398,N_1109,N_1160);
xnor U1399 (N_1399,N_1120,N_1197);
nand U1400 (N_1400,N_1364,N_1329);
xnor U1401 (N_1401,N_1297,N_1384);
or U1402 (N_1402,N_1207,N_1245);
nor U1403 (N_1403,N_1261,N_1208);
and U1404 (N_1404,N_1291,N_1358);
nand U1405 (N_1405,N_1222,N_1340);
nor U1406 (N_1406,N_1242,N_1317);
and U1407 (N_1407,N_1273,N_1354);
or U1408 (N_1408,N_1314,N_1200);
or U1409 (N_1409,N_1378,N_1356);
nand U1410 (N_1410,N_1295,N_1370);
or U1411 (N_1411,N_1375,N_1269);
or U1412 (N_1412,N_1232,N_1316);
and U1413 (N_1413,N_1301,N_1395);
and U1414 (N_1414,N_1216,N_1205);
nand U1415 (N_1415,N_1266,N_1237);
nor U1416 (N_1416,N_1276,N_1377);
and U1417 (N_1417,N_1366,N_1257);
nand U1418 (N_1418,N_1248,N_1286);
and U1419 (N_1419,N_1213,N_1240);
nand U1420 (N_1420,N_1307,N_1253);
or U1421 (N_1421,N_1322,N_1380);
xnor U1422 (N_1422,N_1239,N_1325);
and U1423 (N_1423,N_1290,N_1318);
nand U1424 (N_1424,N_1323,N_1230);
nor U1425 (N_1425,N_1294,N_1350);
nand U1426 (N_1426,N_1399,N_1382);
or U1427 (N_1427,N_1376,N_1274);
nand U1428 (N_1428,N_1303,N_1236);
nor U1429 (N_1429,N_1394,N_1386);
nand U1430 (N_1430,N_1233,N_1228);
and U1431 (N_1431,N_1214,N_1202);
xor U1432 (N_1432,N_1343,N_1328);
nor U1433 (N_1433,N_1357,N_1255);
and U1434 (N_1434,N_1206,N_1372);
and U1435 (N_1435,N_1281,N_1288);
or U1436 (N_1436,N_1299,N_1246);
nand U1437 (N_1437,N_1298,N_1262);
and U1438 (N_1438,N_1341,N_1334);
and U1439 (N_1439,N_1263,N_1231);
nor U1440 (N_1440,N_1308,N_1385);
nand U1441 (N_1441,N_1272,N_1387);
nor U1442 (N_1442,N_1243,N_1339);
nand U1443 (N_1443,N_1300,N_1238);
nor U1444 (N_1444,N_1211,N_1275);
xnor U1445 (N_1445,N_1218,N_1355);
nor U1446 (N_1446,N_1363,N_1285);
nor U1447 (N_1447,N_1241,N_1333);
and U1448 (N_1448,N_1212,N_1360);
nor U1449 (N_1449,N_1381,N_1344);
and U1450 (N_1450,N_1305,N_1292);
nor U1451 (N_1451,N_1264,N_1215);
nand U1452 (N_1452,N_1210,N_1310);
nand U1453 (N_1453,N_1302,N_1280);
and U1454 (N_1454,N_1225,N_1311);
and U1455 (N_1455,N_1226,N_1304);
and U1456 (N_1456,N_1352,N_1379);
nor U1457 (N_1457,N_1369,N_1235);
nor U1458 (N_1458,N_1279,N_1327);
or U1459 (N_1459,N_1244,N_1217);
and U1460 (N_1460,N_1390,N_1251);
nand U1461 (N_1461,N_1320,N_1258);
and U1462 (N_1462,N_1271,N_1249);
or U1463 (N_1463,N_1338,N_1287);
xor U1464 (N_1464,N_1368,N_1351);
or U1465 (N_1465,N_1267,N_1362);
and U1466 (N_1466,N_1284,N_1342);
nand U1467 (N_1467,N_1234,N_1367);
nor U1468 (N_1468,N_1306,N_1309);
or U1469 (N_1469,N_1221,N_1278);
and U1470 (N_1470,N_1256,N_1247);
nor U1471 (N_1471,N_1346,N_1289);
and U1472 (N_1472,N_1321,N_1373);
nand U1473 (N_1473,N_1389,N_1396);
nor U1474 (N_1474,N_1393,N_1283);
nand U1475 (N_1475,N_1365,N_1348);
nor U1476 (N_1476,N_1204,N_1293);
nand U1477 (N_1477,N_1224,N_1220);
nor U1478 (N_1478,N_1331,N_1252);
or U1479 (N_1479,N_1250,N_1259);
nand U1480 (N_1480,N_1270,N_1223);
nor U1481 (N_1481,N_1347,N_1337);
and U1482 (N_1482,N_1229,N_1326);
or U1483 (N_1483,N_1383,N_1361);
or U1484 (N_1484,N_1349,N_1209);
xnor U1485 (N_1485,N_1203,N_1397);
and U1486 (N_1486,N_1315,N_1201);
and U1487 (N_1487,N_1260,N_1359);
nand U1488 (N_1488,N_1296,N_1312);
nor U1489 (N_1489,N_1374,N_1388);
nand U1490 (N_1490,N_1391,N_1227);
and U1491 (N_1491,N_1392,N_1265);
xor U1492 (N_1492,N_1282,N_1336);
or U1493 (N_1493,N_1313,N_1371);
nor U1494 (N_1494,N_1398,N_1268);
or U1495 (N_1495,N_1277,N_1219);
xor U1496 (N_1496,N_1335,N_1330);
and U1497 (N_1497,N_1332,N_1353);
or U1498 (N_1498,N_1324,N_1319);
nand U1499 (N_1499,N_1254,N_1345);
nor U1500 (N_1500,N_1237,N_1240);
nand U1501 (N_1501,N_1360,N_1251);
nor U1502 (N_1502,N_1356,N_1352);
nor U1503 (N_1503,N_1375,N_1382);
and U1504 (N_1504,N_1250,N_1397);
or U1505 (N_1505,N_1243,N_1202);
nor U1506 (N_1506,N_1206,N_1355);
nand U1507 (N_1507,N_1322,N_1246);
nor U1508 (N_1508,N_1397,N_1239);
and U1509 (N_1509,N_1241,N_1240);
and U1510 (N_1510,N_1228,N_1341);
and U1511 (N_1511,N_1222,N_1285);
xnor U1512 (N_1512,N_1220,N_1348);
and U1513 (N_1513,N_1262,N_1367);
and U1514 (N_1514,N_1252,N_1317);
and U1515 (N_1515,N_1332,N_1386);
nand U1516 (N_1516,N_1362,N_1349);
nand U1517 (N_1517,N_1288,N_1360);
nand U1518 (N_1518,N_1210,N_1224);
nor U1519 (N_1519,N_1389,N_1315);
xnor U1520 (N_1520,N_1390,N_1399);
nand U1521 (N_1521,N_1245,N_1251);
xnor U1522 (N_1522,N_1323,N_1318);
nand U1523 (N_1523,N_1218,N_1260);
nor U1524 (N_1524,N_1362,N_1384);
nand U1525 (N_1525,N_1233,N_1317);
and U1526 (N_1526,N_1375,N_1300);
or U1527 (N_1527,N_1282,N_1321);
and U1528 (N_1528,N_1398,N_1369);
nor U1529 (N_1529,N_1373,N_1236);
xor U1530 (N_1530,N_1220,N_1331);
nor U1531 (N_1531,N_1211,N_1248);
or U1532 (N_1532,N_1248,N_1355);
nor U1533 (N_1533,N_1243,N_1387);
nand U1534 (N_1534,N_1397,N_1343);
xnor U1535 (N_1535,N_1291,N_1349);
xor U1536 (N_1536,N_1274,N_1318);
xnor U1537 (N_1537,N_1326,N_1379);
or U1538 (N_1538,N_1305,N_1229);
and U1539 (N_1539,N_1237,N_1244);
or U1540 (N_1540,N_1283,N_1239);
nand U1541 (N_1541,N_1221,N_1363);
xnor U1542 (N_1542,N_1232,N_1396);
xnor U1543 (N_1543,N_1348,N_1223);
or U1544 (N_1544,N_1231,N_1309);
nor U1545 (N_1545,N_1380,N_1225);
nand U1546 (N_1546,N_1395,N_1268);
nand U1547 (N_1547,N_1282,N_1250);
and U1548 (N_1548,N_1253,N_1278);
or U1549 (N_1549,N_1358,N_1386);
and U1550 (N_1550,N_1285,N_1309);
xnor U1551 (N_1551,N_1281,N_1270);
and U1552 (N_1552,N_1233,N_1288);
or U1553 (N_1553,N_1394,N_1235);
nor U1554 (N_1554,N_1240,N_1312);
nand U1555 (N_1555,N_1241,N_1304);
and U1556 (N_1556,N_1365,N_1219);
or U1557 (N_1557,N_1385,N_1332);
nor U1558 (N_1558,N_1226,N_1252);
or U1559 (N_1559,N_1230,N_1394);
nor U1560 (N_1560,N_1253,N_1323);
nand U1561 (N_1561,N_1279,N_1237);
or U1562 (N_1562,N_1388,N_1262);
and U1563 (N_1563,N_1233,N_1245);
nor U1564 (N_1564,N_1205,N_1233);
nand U1565 (N_1565,N_1262,N_1324);
or U1566 (N_1566,N_1341,N_1266);
and U1567 (N_1567,N_1306,N_1280);
xor U1568 (N_1568,N_1209,N_1278);
nand U1569 (N_1569,N_1264,N_1341);
nand U1570 (N_1570,N_1377,N_1226);
nor U1571 (N_1571,N_1396,N_1293);
or U1572 (N_1572,N_1208,N_1210);
or U1573 (N_1573,N_1389,N_1387);
nor U1574 (N_1574,N_1313,N_1238);
xor U1575 (N_1575,N_1331,N_1308);
nand U1576 (N_1576,N_1300,N_1203);
and U1577 (N_1577,N_1398,N_1263);
xor U1578 (N_1578,N_1357,N_1301);
and U1579 (N_1579,N_1212,N_1340);
xor U1580 (N_1580,N_1362,N_1248);
nor U1581 (N_1581,N_1254,N_1212);
nand U1582 (N_1582,N_1329,N_1208);
nand U1583 (N_1583,N_1381,N_1296);
xor U1584 (N_1584,N_1214,N_1300);
nand U1585 (N_1585,N_1266,N_1258);
nand U1586 (N_1586,N_1272,N_1304);
nand U1587 (N_1587,N_1202,N_1369);
and U1588 (N_1588,N_1306,N_1241);
nand U1589 (N_1589,N_1219,N_1221);
or U1590 (N_1590,N_1398,N_1241);
nand U1591 (N_1591,N_1253,N_1304);
nand U1592 (N_1592,N_1383,N_1208);
and U1593 (N_1593,N_1289,N_1396);
or U1594 (N_1594,N_1202,N_1353);
nor U1595 (N_1595,N_1275,N_1373);
nor U1596 (N_1596,N_1306,N_1277);
nor U1597 (N_1597,N_1260,N_1284);
or U1598 (N_1598,N_1269,N_1360);
and U1599 (N_1599,N_1269,N_1313);
nand U1600 (N_1600,N_1529,N_1456);
nand U1601 (N_1601,N_1448,N_1592);
nor U1602 (N_1602,N_1468,N_1508);
nand U1603 (N_1603,N_1413,N_1541);
xor U1604 (N_1604,N_1569,N_1572);
nand U1605 (N_1605,N_1543,N_1493);
nor U1606 (N_1606,N_1513,N_1531);
or U1607 (N_1607,N_1522,N_1482);
nor U1608 (N_1608,N_1471,N_1480);
and U1609 (N_1609,N_1527,N_1442);
and U1610 (N_1610,N_1537,N_1488);
xor U1611 (N_1611,N_1492,N_1417);
nand U1612 (N_1612,N_1574,N_1596);
and U1613 (N_1613,N_1577,N_1426);
nand U1614 (N_1614,N_1521,N_1547);
and U1615 (N_1615,N_1447,N_1431);
nor U1616 (N_1616,N_1584,N_1459);
nand U1617 (N_1617,N_1504,N_1416);
or U1618 (N_1618,N_1441,N_1528);
or U1619 (N_1619,N_1515,N_1418);
or U1620 (N_1620,N_1490,N_1420);
nand U1621 (N_1621,N_1552,N_1463);
xor U1622 (N_1622,N_1562,N_1495);
or U1623 (N_1623,N_1429,N_1462);
or U1624 (N_1624,N_1449,N_1533);
or U1625 (N_1625,N_1491,N_1581);
nand U1626 (N_1626,N_1517,N_1410);
or U1627 (N_1627,N_1496,N_1599);
nor U1628 (N_1628,N_1408,N_1545);
nor U1629 (N_1629,N_1489,N_1444);
nand U1630 (N_1630,N_1433,N_1419);
nor U1631 (N_1631,N_1503,N_1475);
or U1632 (N_1632,N_1576,N_1403);
nor U1633 (N_1633,N_1587,N_1523);
nor U1634 (N_1634,N_1405,N_1483);
nand U1635 (N_1635,N_1556,N_1579);
xor U1636 (N_1636,N_1402,N_1555);
and U1637 (N_1637,N_1437,N_1564);
and U1638 (N_1638,N_1506,N_1518);
nor U1639 (N_1639,N_1477,N_1565);
or U1640 (N_1640,N_1434,N_1571);
nor U1641 (N_1641,N_1414,N_1512);
and U1642 (N_1642,N_1500,N_1466);
nor U1643 (N_1643,N_1582,N_1575);
or U1644 (N_1644,N_1485,N_1542);
and U1645 (N_1645,N_1567,N_1461);
nand U1646 (N_1646,N_1597,N_1554);
nand U1647 (N_1647,N_1526,N_1425);
nand U1648 (N_1648,N_1532,N_1510);
nand U1649 (N_1649,N_1481,N_1427);
nor U1650 (N_1650,N_1558,N_1538);
or U1651 (N_1651,N_1559,N_1585);
nand U1652 (N_1652,N_1573,N_1422);
nor U1653 (N_1653,N_1458,N_1453);
nor U1654 (N_1654,N_1401,N_1476);
and U1655 (N_1655,N_1446,N_1516);
nor U1656 (N_1656,N_1535,N_1469);
nor U1657 (N_1657,N_1568,N_1406);
and U1658 (N_1658,N_1566,N_1474);
and U1659 (N_1659,N_1594,N_1544);
or U1660 (N_1660,N_1472,N_1409);
nand U1661 (N_1661,N_1487,N_1494);
or U1662 (N_1662,N_1451,N_1470);
and U1663 (N_1663,N_1539,N_1583);
nor U1664 (N_1664,N_1550,N_1435);
nor U1665 (N_1665,N_1589,N_1548);
nand U1666 (N_1666,N_1530,N_1588);
nor U1667 (N_1667,N_1452,N_1524);
and U1668 (N_1668,N_1455,N_1478);
nor U1669 (N_1669,N_1505,N_1553);
or U1670 (N_1670,N_1436,N_1595);
or U1671 (N_1671,N_1473,N_1563);
xnor U1672 (N_1672,N_1497,N_1560);
or U1673 (N_1673,N_1432,N_1525);
and U1674 (N_1674,N_1590,N_1519);
nand U1675 (N_1675,N_1514,N_1499);
nor U1676 (N_1676,N_1467,N_1593);
and U1677 (N_1677,N_1501,N_1421);
nor U1678 (N_1678,N_1443,N_1520);
xnor U1679 (N_1679,N_1540,N_1546);
nor U1680 (N_1680,N_1407,N_1536);
nor U1681 (N_1681,N_1465,N_1507);
and U1682 (N_1682,N_1428,N_1598);
nand U1683 (N_1683,N_1534,N_1509);
nand U1684 (N_1684,N_1423,N_1586);
and U1685 (N_1685,N_1498,N_1440);
or U1686 (N_1686,N_1486,N_1549);
or U1687 (N_1687,N_1511,N_1561);
nand U1688 (N_1688,N_1454,N_1412);
and U1689 (N_1689,N_1484,N_1457);
nor U1690 (N_1690,N_1591,N_1570);
nor U1691 (N_1691,N_1578,N_1400);
or U1692 (N_1692,N_1464,N_1460);
and U1693 (N_1693,N_1404,N_1424);
xnor U1694 (N_1694,N_1450,N_1439);
xnor U1695 (N_1695,N_1551,N_1438);
and U1696 (N_1696,N_1580,N_1502);
nor U1697 (N_1697,N_1445,N_1415);
xor U1698 (N_1698,N_1411,N_1479);
nor U1699 (N_1699,N_1557,N_1430);
xnor U1700 (N_1700,N_1442,N_1440);
nor U1701 (N_1701,N_1514,N_1564);
nand U1702 (N_1702,N_1446,N_1545);
nor U1703 (N_1703,N_1465,N_1555);
nand U1704 (N_1704,N_1530,N_1446);
nand U1705 (N_1705,N_1413,N_1563);
nor U1706 (N_1706,N_1434,N_1426);
or U1707 (N_1707,N_1561,N_1543);
and U1708 (N_1708,N_1490,N_1574);
nand U1709 (N_1709,N_1513,N_1432);
nand U1710 (N_1710,N_1597,N_1549);
xor U1711 (N_1711,N_1569,N_1534);
and U1712 (N_1712,N_1544,N_1548);
and U1713 (N_1713,N_1492,N_1533);
and U1714 (N_1714,N_1557,N_1594);
nand U1715 (N_1715,N_1492,N_1443);
nor U1716 (N_1716,N_1523,N_1479);
nor U1717 (N_1717,N_1552,N_1561);
or U1718 (N_1718,N_1445,N_1560);
nand U1719 (N_1719,N_1419,N_1507);
xor U1720 (N_1720,N_1413,N_1500);
or U1721 (N_1721,N_1404,N_1489);
xor U1722 (N_1722,N_1544,N_1434);
or U1723 (N_1723,N_1459,N_1512);
or U1724 (N_1724,N_1530,N_1538);
or U1725 (N_1725,N_1546,N_1499);
or U1726 (N_1726,N_1401,N_1502);
and U1727 (N_1727,N_1533,N_1454);
or U1728 (N_1728,N_1473,N_1576);
nand U1729 (N_1729,N_1503,N_1481);
and U1730 (N_1730,N_1530,N_1569);
nand U1731 (N_1731,N_1552,N_1590);
nor U1732 (N_1732,N_1585,N_1504);
nand U1733 (N_1733,N_1556,N_1411);
nand U1734 (N_1734,N_1449,N_1493);
and U1735 (N_1735,N_1496,N_1426);
nor U1736 (N_1736,N_1566,N_1454);
nand U1737 (N_1737,N_1567,N_1482);
nor U1738 (N_1738,N_1455,N_1475);
or U1739 (N_1739,N_1511,N_1529);
and U1740 (N_1740,N_1439,N_1443);
and U1741 (N_1741,N_1489,N_1599);
or U1742 (N_1742,N_1564,N_1555);
nand U1743 (N_1743,N_1420,N_1407);
nor U1744 (N_1744,N_1551,N_1492);
nand U1745 (N_1745,N_1539,N_1575);
nand U1746 (N_1746,N_1505,N_1587);
nor U1747 (N_1747,N_1512,N_1570);
nor U1748 (N_1748,N_1525,N_1576);
or U1749 (N_1749,N_1592,N_1456);
nor U1750 (N_1750,N_1490,N_1408);
or U1751 (N_1751,N_1548,N_1422);
or U1752 (N_1752,N_1415,N_1403);
or U1753 (N_1753,N_1577,N_1419);
nand U1754 (N_1754,N_1512,N_1407);
nand U1755 (N_1755,N_1506,N_1583);
nor U1756 (N_1756,N_1556,N_1472);
nand U1757 (N_1757,N_1567,N_1402);
or U1758 (N_1758,N_1595,N_1531);
or U1759 (N_1759,N_1432,N_1550);
nand U1760 (N_1760,N_1492,N_1461);
nand U1761 (N_1761,N_1557,N_1515);
and U1762 (N_1762,N_1581,N_1521);
and U1763 (N_1763,N_1503,N_1484);
nand U1764 (N_1764,N_1584,N_1418);
or U1765 (N_1765,N_1535,N_1549);
or U1766 (N_1766,N_1517,N_1405);
or U1767 (N_1767,N_1431,N_1499);
and U1768 (N_1768,N_1419,N_1576);
and U1769 (N_1769,N_1490,N_1597);
or U1770 (N_1770,N_1529,N_1531);
nor U1771 (N_1771,N_1464,N_1575);
nor U1772 (N_1772,N_1418,N_1511);
and U1773 (N_1773,N_1444,N_1469);
or U1774 (N_1774,N_1417,N_1504);
or U1775 (N_1775,N_1437,N_1450);
nor U1776 (N_1776,N_1543,N_1564);
xor U1777 (N_1777,N_1503,N_1412);
nor U1778 (N_1778,N_1532,N_1431);
xnor U1779 (N_1779,N_1491,N_1577);
and U1780 (N_1780,N_1534,N_1590);
nand U1781 (N_1781,N_1519,N_1463);
or U1782 (N_1782,N_1518,N_1562);
and U1783 (N_1783,N_1548,N_1431);
xnor U1784 (N_1784,N_1445,N_1587);
xor U1785 (N_1785,N_1534,N_1403);
nor U1786 (N_1786,N_1583,N_1571);
or U1787 (N_1787,N_1535,N_1486);
nand U1788 (N_1788,N_1506,N_1588);
or U1789 (N_1789,N_1473,N_1407);
or U1790 (N_1790,N_1574,N_1434);
nor U1791 (N_1791,N_1449,N_1485);
nor U1792 (N_1792,N_1535,N_1424);
nand U1793 (N_1793,N_1436,N_1432);
nand U1794 (N_1794,N_1413,N_1493);
nor U1795 (N_1795,N_1508,N_1409);
nor U1796 (N_1796,N_1570,N_1533);
or U1797 (N_1797,N_1597,N_1548);
or U1798 (N_1798,N_1588,N_1462);
nor U1799 (N_1799,N_1596,N_1582);
nand U1800 (N_1800,N_1724,N_1604);
nor U1801 (N_1801,N_1776,N_1644);
or U1802 (N_1802,N_1679,N_1799);
nor U1803 (N_1803,N_1703,N_1698);
xnor U1804 (N_1804,N_1757,N_1655);
or U1805 (N_1805,N_1700,N_1663);
nor U1806 (N_1806,N_1603,N_1717);
nor U1807 (N_1807,N_1742,N_1768);
nand U1808 (N_1808,N_1601,N_1719);
nand U1809 (N_1809,N_1647,N_1634);
and U1810 (N_1810,N_1760,N_1783);
or U1811 (N_1811,N_1710,N_1685);
nand U1812 (N_1812,N_1635,N_1779);
and U1813 (N_1813,N_1752,N_1649);
and U1814 (N_1814,N_1730,N_1781);
and U1815 (N_1815,N_1751,N_1739);
xnor U1816 (N_1816,N_1636,N_1676);
and U1817 (N_1817,N_1640,N_1766);
or U1818 (N_1818,N_1639,N_1792);
nor U1819 (N_1819,N_1729,N_1771);
and U1820 (N_1820,N_1615,N_1780);
xnor U1821 (N_1821,N_1697,N_1622);
and U1822 (N_1822,N_1756,N_1787);
nand U1823 (N_1823,N_1723,N_1687);
nand U1824 (N_1824,N_1797,N_1628);
or U1825 (N_1825,N_1788,N_1732);
or U1826 (N_1826,N_1795,N_1782);
or U1827 (N_1827,N_1664,N_1632);
nor U1828 (N_1828,N_1642,N_1621);
or U1829 (N_1829,N_1674,N_1606);
and U1830 (N_1830,N_1608,N_1683);
nand U1831 (N_1831,N_1708,N_1706);
nand U1832 (N_1832,N_1662,N_1716);
xor U1833 (N_1833,N_1772,N_1747);
or U1834 (N_1834,N_1633,N_1619);
nor U1835 (N_1835,N_1623,N_1793);
or U1836 (N_1836,N_1738,N_1680);
xnor U1837 (N_1837,N_1785,N_1670);
nand U1838 (N_1838,N_1722,N_1629);
and U1839 (N_1839,N_1727,N_1753);
and U1840 (N_1840,N_1651,N_1614);
or U1841 (N_1841,N_1611,N_1652);
nor U1842 (N_1842,N_1654,N_1607);
or U1843 (N_1843,N_1746,N_1713);
nand U1844 (N_1844,N_1759,N_1627);
xor U1845 (N_1845,N_1744,N_1733);
nor U1846 (N_1846,N_1696,N_1602);
xor U1847 (N_1847,N_1682,N_1789);
nand U1848 (N_1848,N_1638,N_1725);
nand U1849 (N_1849,N_1677,N_1758);
and U1850 (N_1850,N_1686,N_1688);
xnor U1851 (N_1851,N_1726,N_1743);
nand U1852 (N_1852,N_1650,N_1714);
xnor U1853 (N_1853,N_1728,N_1731);
nand U1854 (N_1854,N_1645,N_1736);
nor U1855 (N_1855,N_1796,N_1624);
and U1856 (N_1856,N_1612,N_1798);
nand U1857 (N_1857,N_1720,N_1734);
or U1858 (N_1858,N_1765,N_1770);
nor U1859 (N_1859,N_1620,N_1681);
and U1860 (N_1860,N_1660,N_1721);
and U1861 (N_1861,N_1745,N_1653);
nor U1862 (N_1862,N_1661,N_1630);
xnor U1863 (N_1863,N_1672,N_1626);
xor U1864 (N_1864,N_1666,N_1673);
or U1865 (N_1865,N_1605,N_1637);
nand U1866 (N_1866,N_1616,N_1618);
nand U1867 (N_1867,N_1718,N_1689);
and U1868 (N_1868,N_1643,N_1699);
or U1869 (N_1869,N_1773,N_1600);
xor U1870 (N_1870,N_1669,N_1707);
nor U1871 (N_1871,N_1786,N_1657);
or U1872 (N_1872,N_1684,N_1778);
nand U1873 (N_1873,N_1748,N_1695);
or U1874 (N_1874,N_1763,N_1694);
or U1875 (N_1875,N_1755,N_1737);
xor U1876 (N_1876,N_1646,N_1774);
nor U1877 (N_1877,N_1794,N_1690);
nand U1878 (N_1878,N_1784,N_1692);
nand U1879 (N_1879,N_1702,N_1775);
nor U1880 (N_1880,N_1658,N_1659);
or U1881 (N_1881,N_1675,N_1648);
nand U1882 (N_1882,N_1631,N_1705);
nor U1883 (N_1883,N_1656,N_1667);
nand U1884 (N_1884,N_1791,N_1712);
nand U1885 (N_1885,N_1691,N_1764);
xor U1886 (N_1886,N_1641,N_1617);
nand U1887 (N_1887,N_1678,N_1767);
and U1888 (N_1888,N_1693,N_1715);
xnor U1889 (N_1889,N_1741,N_1671);
xnor U1890 (N_1890,N_1665,N_1761);
nand U1891 (N_1891,N_1610,N_1749);
or U1892 (N_1892,N_1735,N_1709);
or U1893 (N_1893,N_1625,N_1754);
and U1894 (N_1894,N_1790,N_1609);
and U1895 (N_1895,N_1668,N_1777);
nand U1896 (N_1896,N_1750,N_1769);
and U1897 (N_1897,N_1740,N_1704);
or U1898 (N_1898,N_1701,N_1613);
nand U1899 (N_1899,N_1711,N_1762);
xor U1900 (N_1900,N_1733,N_1687);
nand U1901 (N_1901,N_1689,N_1608);
or U1902 (N_1902,N_1792,N_1628);
and U1903 (N_1903,N_1631,N_1703);
nand U1904 (N_1904,N_1722,N_1755);
and U1905 (N_1905,N_1707,N_1776);
or U1906 (N_1906,N_1724,N_1743);
or U1907 (N_1907,N_1728,N_1750);
nand U1908 (N_1908,N_1792,N_1624);
xor U1909 (N_1909,N_1714,N_1657);
and U1910 (N_1910,N_1614,N_1662);
nand U1911 (N_1911,N_1621,N_1747);
nand U1912 (N_1912,N_1613,N_1621);
or U1913 (N_1913,N_1795,N_1696);
or U1914 (N_1914,N_1695,N_1684);
and U1915 (N_1915,N_1636,N_1692);
nor U1916 (N_1916,N_1767,N_1649);
and U1917 (N_1917,N_1609,N_1796);
or U1918 (N_1918,N_1773,N_1624);
nor U1919 (N_1919,N_1751,N_1695);
xor U1920 (N_1920,N_1723,N_1752);
and U1921 (N_1921,N_1776,N_1712);
nor U1922 (N_1922,N_1697,N_1761);
xor U1923 (N_1923,N_1770,N_1766);
and U1924 (N_1924,N_1747,N_1762);
nor U1925 (N_1925,N_1612,N_1734);
nand U1926 (N_1926,N_1624,N_1672);
or U1927 (N_1927,N_1789,N_1633);
and U1928 (N_1928,N_1606,N_1718);
or U1929 (N_1929,N_1729,N_1615);
nor U1930 (N_1930,N_1799,N_1797);
nor U1931 (N_1931,N_1683,N_1750);
or U1932 (N_1932,N_1601,N_1777);
or U1933 (N_1933,N_1690,N_1753);
nor U1934 (N_1934,N_1759,N_1771);
or U1935 (N_1935,N_1750,N_1753);
nand U1936 (N_1936,N_1601,N_1788);
and U1937 (N_1937,N_1668,N_1667);
and U1938 (N_1938,N_1680,N_1626);
and U1939 (N_1939,N_1672,N_1710);
nand U1940 (N_1940,N_1730,N_1665);
nand U1941 (N_1941,N_1652,N_1657);
or U1942 (N_1942,N_1716,N_1626);
nor U1943 (N_1943,N_1643,N_1654);
and U1944 (N_1944,N_1610,N_1658);
or U1945 (N_1945,N_1662,N_1668);
nor U1946 (N_1946,N_1677,N_1711);
or U1947 (N_1947,N_1686,N_1624);
and U1948 (N_1948,N_1726,N_1757);
nand U1949 (N_1949,N_1687,N_1601);
or U1950 (N_1950,N_1786,N_1735);
nor U1951 (N_1951,N_1781,N_1745);
nand U1952 (N_1952,N_1603,N_1669);
nand U1953 (N_1953,N_1772,N_1665);
and U1954 (N_1954,N_1650,N_1790);
nor U1955 (N_1955,N_1763,N_1703);
nor U1956 (N_1956,N_1608,N_1775);
nand U1957 (N_1957,N_1662,N_1760);
nor U1958 (N_1958,N_1667,N_1770);
or U1959 (N_1959,N_1634,N_1759);
nand U1960 (N_1960,N_1620,N_1689);
and U1961 (N_1961,N_1684,N_1645);
and U1962 (N_1962,N_1608,N_1609);
and U1963 (N_1963,N_1606,N_1603);
nand U1964 (N_1964,N_1613,N_1691);
nor U1965 (N_1965,N_1607,N_1600);
or U1966 (N_1966,N_1656,N_1736);
and U1967 (N_1967,N_1637,N_1788);
nand U1968 (N_1968,N_1789,N_1631);
or U1969 (N_1969,N_1733,N_1748);
xor U1970 (N_1970,N_1666,N_1665);
nand U1971 (N_1971,N_1615,N_1635);
and U1972 (N_1972,N_1700,N_1677);
nand U1973 (N_1973,N_1790,N_1701);
xnor U1974 (N_1974,N_1797,N_1605);
or U1975 (N_1975,N_1672,N_1601);
nor U1976 (N_1976,N_1738,N_1759);
or U1977 (N_1977,N_1727,N_1663);
xor U1978 (N_1978,N_1737,N_1653);
and U1979 (N_1979,N_1716,N_1624);
or U1980 (N_1980,N_1628,N_1696);
xor U1981 (N_1981,N_1742,N_1711);
xnor U1982 (N_1982,N_1627,N_1628);
nand U1983 (N_1983,N_1696,N_1750);
nor U1984 (N_1984,N_1734,N_1663);
nor U1985 (N_1985,N_1654,N_1624);
nor U1986 (N_1986,N_1600,N_1690);
or U1987 (N_1987,N_1758,N_1772);
and U1988 (N_1988,N_1761,N_1636);
xnor U1989 (N_1989,N_1669,N_1622);
and U1990 (N_1990,N_1673,N_1729);
xor U1991 (N_1991,N_1775,N_1705);
xor U1992 (N_1992,N_1720,N_1646);
nor U1993 (N_1993,N_1645,N_1602);
or U1994 (N_1994,N_1664,N_1602);
and U1995 (N_1995,N_1629,N_1668);
xnor U1996 (N_1996,N_1653,N_1601);
nand U1997 (N_1997,N_1784,N_1731);
or U1998 (N_1998,N_1699,N_1725);
or U1999 (N_1999,N_1672,N_1641);
nand U2000 (N_2000,N_1899,N_1897);
nor U2001 (N_2001,N_1964,N_1985);
nor U2002 (N_2002,N_1821,N_1843);
nand U2003 (N_2003,N_1888,N_1959);
or U2004 (N_2004,N_1979,N_1890);
and U2005 (N_2005,N_1997,N_1858);
xor U2006 (N_2006,N_1823,N_1913);
nand U2007 (N_2007,N_1983,N_1884);
nand U2008 (N_2008,N_1999,N_1931);
and U2009 (N_2009,N_1977,N_1834);
nand U2010 (N_2010,N_1819,N_1947);
nand U2011 (N_2011,N_1911,N_1809);
and U2012 (N_2012,N_1831,N_1830);
nand U2013 (N_2013,N_1989,N_1838);
nand U2014 (N_2014,N_1863,N_1956);
or U2015 (N_2015,N_1871,N_1867);
nor U2016 (N_2016,N_1820,N_1854);
or U2017 (N_2017,N_1986,N_1844);
and U2018 (N_2018,N_1875,N_1877);
and U2019 (N_2019,N_1827,N_1816);
or U2020 (N_2020,N_1857,N_1924);
nor U2021 (N_2021,N_1958,N_1992);
and U2022 (N_2022,N_1932,N_1852);
nand U2023 (N_2023,N_1876,N_1918);
xor U2024 (N_2024,N_1869,N_1960);
nor U2025 (N_2025,N_1800,N_1904);
nand U2026 (N_2026,N_1967,N_1900);
nand U2027 (N_2027,N_1920,N_1984);
xor U2028 (N_2028,N_1982,N_1970);
nand U2029 (N_2029,N_1923,N_1865);
nor U2030 (N_2030,N_1998,N_1901);
or U2031 (N_2031,N_1889,N_1872);
and U2032 (N_2032,N_1829,N_1939);
nand U2033 (N_2033,N_1946,N_1929);
xnor U2034 (N_2034,N_1938,N_1811);
nor U2035 (N_2035,N_1935,N_1808);
nand U2036 (N_2036,N_1914,N_1933);
and U2037 (N_2037,N_1953,N_1822);
nor U2038 (N_2038,N_1955,N_1882);
nand U2039 (N_2039,N_1801,N_1883);
or U2040 (N_2040,N_1978,N_1824);
nor U2041 (N_2041,N_1954,N_1804);
or U2042 (N_2042,N_1928,N_1893);
nand U2043 (N_2043,N_1862,N_1995);
and U2044 (N_2044,N_1826,N_1942);
and U2045 (N_2045,N_1891,N_1870);
and U2046 (N_2046,N_1910,N_1895);
or U2047 (N_2047,N_1813,N_1806);
and U2048 (N_2048,N_1969,N_1845);
or U2049 (N_2049,N_1856,N_1837);
nand U2050 (N_2050,N_1803,N_1952);
or U2051 (N_2051,N_1907,N_1990);
nand U2052 (N_2052,N_1915,N_1850);
or U2053 (N_2053,N_1925,N_1868);
and U2054 (N_2054,N_1817,N_1896);
and U2055 (N_2055,N_1963,N_1934);
nor U2056 (N_2056,N_1842,N_1941);
and U2057 (N_2057,N_1859,N_1885);
xnor U2058 (N_2058,N_1951,N_1987);
and U2059 (N_2059,N_1917,N_1840);
nor U2060 (N_2060,N_1905,N_1881);
xnor U2061 (N_2061,N_1825,N_1849);
and U2062 (N_2062,N_1957,N_1873);
nand U2063 (N_2063,N_1846,N_1880);
nand U2064 (N_2064,N_1972,N_1861);
nand U2065 (N_2065,N_1878,N_1912);
nand U2066 (N_2066,N_1903,N_1994);
nand U2067 (N_2067,N_1835,N_1805);
or U2068 (N_2068,N_1906,N_1927);
nor U2069 (N_2069,N_1949,N_1996);
nor U2070 (N_2070,N_1810,N_1828);
nor U2071 (N_2071,N_1836,N_1973);
nand U2072 (N_2072,N_1866,N_1909);
and U2073 (N_2073,N_1833,N_1965);
nor U2074 (N_2074,N_1926,N_1894);
nand U2075 (N_2075,N_1945,N_1980);
nor U2076 (N_2076,N_1937,N_1874);
nand U2077 (N_2077,N_1892,N_1807);
or U2078 (N_2078,N_1860,N_1887);
and U2079 (N_2079,N_1848,N_1993);
nand U2080 (N_2080,N_1902,N_1847);
nand U2081 (N_2081,N_1940,N_1864);
nand U2082 (N_2082,N_1812,N_1841);
nor U2083 (N_2083,N_1919,N_1802);
or U2084 (N_2084,N_1961,N_1948);
and U2085 (N_2085,N_1922,N_1975);
nor U2086 (N_2086,N_1886,N_1930);
and U2087 (N_2087,N_1832,N_1851);
xor U2088 (N_2088,N_1981,N_1879);
and U2089 (N_2089,N_1943,N_1971);
nand U2090 (N_2090,N_1916,N_1815);
and U2091 (N_2091,N_1908,N_1962);
nor U2092 (N_2092,N_1991,N_1936);
nand U2093 (N_2093,N_1898,N_1818);
xor U2094 (N_2094,N_1855,N_1988);
xnor U2095 (N_2095,N_1814,N_1950);
xnor U2096 (N_2096,N_1839,N_1921);
nand U2097 (N_2097,N_1944,N_1974);
nor U2098 (N_2098,N_1968,N_1853);
and U2099 (N_2099,N_1966,N_1976);
and U2100 (N_2100,N_1965,N_1810);
or U2101 (N_2101,N_1880,N_1886);
or U2102 (N_2102,N_1934,N_1940);
and U2103 (N_2103,N_1867,N_1920);
or U2104 (N_2104,N_1836,N_1952);
xnor U2105 (N_2105,N_1873,N_1827);
nand U2106 (N_2106,N_1925,N_1954);
nand U2107 (N_2107,N_1890,N_1868);
or U2108 (N_2108,N_1937,N_1970);
or U2109 (N_2109,N_1847,N_1906);
and U2110 (N_2110,N_1834,N_1830);
and U2111 (N_2111,N_1871,N_1924);
or U2112 (N_2112,N_1812,N_1923);
nor U2113 (N_2113,N_1934,N_1982);
nand U2114 (N_2114,N_1856,N_1977);
and U2115 (N_2115,N_1848,N_1832);
and U2116 (N_2116,N_1959,N_1891);
nor U2117 (N_2117,N_1983,N_1972);
or U2118 (N_2118,N_1868,N_1865);
and U2119 (N_2119,N_1948,N_1875);
xor U2120 (N_2120,N_1955,N_1964);
or U2121 (N_2121,N_1900,N_1979);
nand U2122 (N_2122,N_1871,N_1851);
nor U2123 (N_2123,N_1860,N_1921);
or U2124 (N_2124,N_1870,N_1985);
nand U2125 (N_2125,N_1833,N_1857);
nor U2126 (N_2126,N_1912,N_1806);
nor U2127 (N_2127,N_1960,N_1915);
nor U2128 (N_2128,N_1972,N_1813);
nand U2129 (N_2129,N_1923,N_1881);
and U2130 (N_2130,N_1890,N_1975);
nand U2131 (N_2131,N_1815,N_1926);
or U2132 (N_2132,N_1864,N_1952);
and U2133 (N_2133,N_1913,N_1825);
nand U2134 (N_2134,N_1952,N_1943);
nor U2135 (N_2135,N_1877,N_1822);
nor U2136 (N_2136,N_1962,N_1926);
nor U2137 (N_2137,N_1850,N_1810);
and U2138 (N_2138,N_1809,N_1979);
and U2139 (N_2139,N_1916,N_1942);
xnor U2140 (N_2140,N_1904,N_1943);
or U2141 (N_2141,N_1993,N_1876);
nand U2142 (N_2142,N_1997,N_1857);
or U2143 (N_2143,N_1901,N_1824);
and U2144 (N_2144,N_1829,N_1911);
and U2145 (N_2145,N_1925,N_1989);
nor U2146 (N_2146,N_1857,N_1832);
and U2147 (N_2147,N_1869,N_1985);
or U2148 (N_2148,N_1966,N_1937);
and U2149 (N_2149,N_1848,N_1809);
xor U2150 (N_2150,N_1847,N_1983);
nor U2151 (N_2151,N_1912,N_1981);
or U2152 (N_2152,N_1944,N_1940);
and U2153 (N_2153,N_1822,N_1908);
nor U2154 (N_2154,N_1972,N_1842);
or U2155 (N_2155,N_1901,N_1839);
nor U2156 (N_2156,N_1987,N_1917);
and U2157 (N_2157,N_1997,N_1961);
nor U2158 (N_2158,N_1901,N_1858);
xnor U2159 (N_2159,N_1823,N_1966);
nor U2160 (N_2160,N_1908,N_1970);
or U2161 (N_2161,N_1974,N_1947);
nand U2162 (N_2162,N_1932,N_1995);
and U2163 (N_2163,N_1954,N_1864);
nand U2164 (N_2164,N_1851,N_1986);
or U2165 (N_2165,N_1804,N_1845);
nor U2166 (N_2166,N_1994,N_1950);
and U2167 (N_2167,N_1932,N_1918);
or U2168 (N_2168,N_1935,N_1890);
nand U2169 (N_2169,N_1895,N_1848);
nor U2170 (N_2170,N_1912,N_1938);
nor U2171 (N_2171,N_1865,N_1850);
nor U2172 (N_2172,N_1863,N_1803);
and U2173 (N_2173,N_1900,N_1877);
nor U2174 (N_2174,N_1935,N_1989);
and U2175 (N_2175,N_1879,N_1976);
and U2176 (N_2176,N_1928,N_1901);
and U2177 (N_2177,N_1883,N_1928);
and U2178 (N_2178,N_1912,N_1950);
and U2179 (N_2179,N_1935,N_1934);
nand U2180 (N_2180,N_1896,N_1925);
and U2181 (N_2181,N_1965,N_1877);
xor U2182 (N_2182,N_1884,N_1845);
xnor U2183 (N_2183,N_1912,N_1989);
nor U2184 (N_2184,N_1911,N_1962);
and U2185 (N_2185,N_1880,N_1904);
nor U2186 (N_2186,N_1862,N_1878);
nor U2187 (N_2187,N_1895,N_1887);
or U2188 (N_2188,N_1863,N_1815);
nor U2189 (N_2189,N_1941,N_1860);
and U2190 (N_2190,N_1865,N_1826);
nand U2191 (N_2191,N_1946,N_1836);
and U2192 (N_2192,N_1806,N_1929);
or U2193 (N_2193,N_1849,N_1996);
or U2194 (N_2194,N_1840,N_1801);
or U2195 (N_2195,N_1875,N_1980);
and U2196 (N_2196,N_1914,N_1985);
and U2197 (N_2197,N_1835,N_1894);
or U2198 (N_2198,N_1904,N_1976);
nor U2199 (N_2199,N_1988,N_1878);
nor U2200 (N_2200,N_2008,N_2030);
nand U2201 (N_2201,N_2049,N_2115);
nor U2202 (N_2202,N_2058,N_2134);
nor U2203 (N_2203,N_2188,N_2136);
nand U2204 (N_2204,N_2164,N_2198);
or U2205 (N_2205,N_2040,N_2138);
and U2206 (N_2206,N_2137,N_2003);
nor U2207 (N_2207,N_2035,N_2123);
xnor U2208 (N_2208,N_2166,N_2154);
or U2209 (N_2209,N_2048,N_2026);
nand U2210 (N_2210,N_2055,N_2036);
nor U2211 (N_2211,N_2087,N_2183);
and U2212 (N_2212,N_2075,N_2015);
or U2213 (N_2213,N_2106,N_2014);
nand U2214 (N_2214,N_2100,N_2090);
and U2215 (N_2215,N_2047,N_2020);
nor U2216 (N_2216,N_2065,N_2152);
and U2217 (N_2217,N_2129,N_2174);
and U2218 (N_2218,N_2162,N_2175);
nor U2219 (N_2219,N_2051,N_2000);
nor U2220 (N_2220,N_2170,N_2176);
and U2221 (N_2221,N_2028,N_2172);
nor U2222 (N_2222,N_2144,N_2022);
nand U2223 (N_2223,N_2073,N_2041);
and U2224 (N_2224,N_2156,N_2013);
and U2225 (N_2225,N_2007,N_2159);
nand U2226 (N_2226,N_2187,N_2112);
nand U2227 (N_2227,N_2093,N_2179);
nor U2228 (N_2228,N_2023,N_2119);
nand U2229 (N_2229,N_2109,N_2042);
and U2230 (N_2230,N_2088,N_2155);
xor U2231 (N_2231,N_2016,N_2089);
nand U2232 (N_2232,N_2105,N_2113);
xor U2233 (N_2233,N_2095,N_2169);
and U2234 (N_2234,N_2128,N_2104);
nand U2235 (N_2235,N_2146,N_2149);
nor U2236 (N_2236,N_2139,N_2182);
and U2237 (N_2237,N_2173,N_2191);
nor U2238 (N_2238,N_2045,N_2120);
nand U2239 (N_2239,N_2143,N_2083);
nor U2240 (N_2240,N_2130,N_2084);
or U2241 (N_2241,N_2181,N_2163);
nor U2242 (N_2242,N_2079,N_2150);
nand U2243 (N_2243,N_2186,N_2027);
and U2244 (N_2244,N_2068,N_2012);
nor U2245 (N_2245,N_2161,N_2011);
nand U2246 (N_2246,N_2001,N_2018);
and U2247 (N_2247,N_2124,N_2133);
xor U2248 (N_2248,N_2009,N_2140);
nor U2249 (N_2249,N_2178,N_2078);
or U2250 (N_2250,N_2094,N_2033);
or U2251 (N_2251,N_2092,N_2039);
and U2252 (N_2252,N_2168,N_2102);
nand U2253 (N_2253,N_2190,N_2167);
or U2254 (N_2254,N_2010,N_2158);
and U2255 (N_2255,N_2085,N_2153);
or U2256 (N_2256,N_2029,N_2116);
nand U2257 (N_2257,N_2070,N_2147);
nor U2258 (N_2258,N_2103,N_2184);
or U2259 (N_2259,N_2086,N_2050);
nor U2260 (N_2260,N_2122,N_2031);
nand U2261 (N_2261,N_2072,N_2132);
nor U2262 (N_2262,N_2197,N_2141);
and U2263 (N_2263,N_2193,N_2034);
nand U2264 (N_2264,N_2037,N_2151);
nand U2265 (N_2265,N_2192,N_2056);
nor U2266 (N_2266,N_2077,N_2101);
and U2267 (N_2267,N_2004,N_2189);
or U2268 (N_2268,N_2062,N_2064);
nand U2269 (N_2269,N_2098,N_2021);
nor U2270 (N_2270,N_2121,N_2135);
or U2271 (N_2271,N_2160,N_2024);
or U2272 (N_2272,N_2125,N_2131);
xor U2273 (N_2273,N_2043,N_2061);
nand U2274 (N_2274,N_2006,N_2196);
and U2275 (N_2275,N_2057,N_2082);
or U2276 (N_2276,N_2180,N_2091);
or U2277 (N_2277,N_2096,N_2145);
nand U2278 (N_2278,N_2046,N_2017);
nor U2279 (N_2279,N_2142,N_2019);
and U2280 (N_2280,N_2165,N_2108);
and U2281 (N_2281,N_2118,N_2071);
and U2282 (N_2282,N_2059,N_2076);
and U2283 (N_2283,N_2052,N_2063);
or U2284 (N_2284,N_2157,N_2097);
nor U2285 (N_2285,N_2107,N_2032);
or U2286 (N_2286,N_2044,N_2195);
nor U2287 (N_2287,N_2053,N_2081);
or U2288 (N_2288,N_2074,N_2002);
or U2289 (N_2289,N_2038,N_2117);
and U2290 (N_2290,N_2080,N_2194);
nor U2291 (N_2291,N_2025,N_2067);
nand U2292 (N_2292,N_2069,N_2199);
and U2293 (N_2293,N_2005,N_2114);
nand U2294 (N_2294,N_2054,N_2066);
nand U2295 (N_2295,N_2110,N_2148);
nor U2296 (N_2296,N_2111,N_2171);
nand U2297 (N_2297,N_2126,N_2060);
or U2298 (N_2298,N_2127,N_2185);
nand U2299 (N_2299,N_2177,N_2099);
nor U2300 (N_2300,N_2126,N_2089);
or U2301 (N_2301,N_2075,N_2188);
and U2302 (N_2302,N_2045,N_2101);
nor U2303 (N_2303,N_2068,N_2141);
and U2304 (N_2304,N_2152,N_2113);
nor U2305 (N_2305,N_2121,N_2189);
and U2306 (N_2306,N_2030,N_2163);
and U2307 (N_2307,N_2117,N_2160);
and U2308 (N_2308,N_2007,N_2078);
nand U2309 (N_2309,N_2176,N_2093);
nor U2310 (N_2310,N_2111,N_2146);
xor U2311 (N_2311,N_2103,N_2019);
xor U2312 (N_2312,N_2122,N_2195);
nor U2313 (N_2313,N_2066,N_2028);
nor U2314 (N_2314,N_2081,N_2069);
nand U2315 (N_2315,N_2117,N_2178);
and U2316 (N_2316,N_2130,N_2051);
nand U2317 (N_2317,N_2130,N_2007);
and U2318 (N_2318,N_2025,N_2102);
or U2319 (N_2319,N_2168,N_2178);
nor U2320 (N_2320,N_2127,N_2026);
or U2321 (N_2321,N_2045,N_2141);
nor U2322 (N_2322,N_2011,N_2159);
nor U2323 (N_2323,N_2004,N_2088);
or U2324 (N_2324,N_2056,N_2014);
or U2325 (N_2325,N_2019,N_2156);
and U2326 (N_2326,N_2020,N_2022);
xor U2327 (N_2327,N_2190,N_2032);
and U2328 (N_2328,N_2189,N_2147);
and U2329 (N_2329,N_2184,N_2119);
nand U2330 (N_2330,N_2166,N_2010);
or U2331 (N_2331,N_2170,N_2085);
nand U2332 (N_2332,N_2084,N_2127);
or U2333 (N_2333,N_2068,N_2078);
nand U2334 (N_2334,N_2151,N_2093);
nand U2335 (N_2335,N_2052,N_2121);
or U2336 (N_2336,N_2076,N_2108);
nand U2337 (N_2337,N_2121,N_2199);
and U2338 (N_2338,N_2110,N_2169);
or U2339 (N_2339,N_2069,N_2119);
nor U2340 (N_2340,N_2020,N_2026);
nor U2341 (N_2341,N_2192,N_2163);
nand U2342 (N_2342,N_2156,N_2122);
nand U2343 (N_2343,N_2018,N_2144);
and U2344 (N_2344,N_2041,N_2001);
nor U2345 (N_2345,N_2117,N_2150);
xnor U2346 (N_2346,N_2192,N_2059);
nand U2347 (N_2347,N_2165,N_2192);
and U2348 (N_2348,N_2180,N_2190);
nor U2349 (N_2349,N_2020,N_2096);
xnor U2350 (N_2350,N_2164,N_2185);
nor U2351 (N_2351,N_2135,N_2157);
nand U2352 (N_2352,N_2187,N_2133);
nor U2353 (N_2353,N_2090,N_2143);
nand U2354 (N_2354,N_2067,N_2183);
nor U2355 (N_2355,N_2127,N_2199);
or U2356 (N_2356,N_2131,N_2041);
nand U2357 (N_2357,N_2098,N_2135);
nand U2358 (N_2358,N_2188,N_2000);
and U2359 (N_2359,N_2189,N_2024);
xnor U2360 (N_2360,N_2123,N_2157);
nor U2361 (N_2361,N_2147,N_2063);
xor U2362 (N_2362,N_2142,N_2056);
xnor U2363 (N_2363,N_2042,N_2110);
nor U2364 (N_2364,N_2013,N_2169);
and U2365 (N_2365,N_2029,N_2000);
and U2366 (N_2366,N_2000,N_2032);
xnor U2367 (N_2367,N_2123,N_2050);
nand U2368 (N_2368,N_2082,N_2052);
or U2369 (N_2369,N_2049,N_2123);
or U2370 (N_2370,N_2071,N_2104);
nand U2371 (N_2371,N_2109,N_2058);
and U2372 (N_2372,N_2070,N_2058);
xor U2373 (N_2373,N_2124,N_2040);
nand U2374 (N_2374,N_2183,N_2009);
or U2375 (N_2375,N_2165,N_2154);
nor U2376 (N_2376,N_2051,N_2170);
nor U2377 (N_2377,N_2198,N_2076);
and U2378 (N_2378,N_2162,N_2159);
nand U2379 (N_2379,N_2182,N_2055);
nand U2380 (N_2380,N_2069,N_2077);
nor U2381 (N_2381,N_2103,N_2067);
xor U2382 (N_2382,N_2133,N_2128);
nand U2383 (N_2383,N_2038,N_2188);
nand U2384 (N_2384,N_2181,N_2043);
xor U2385 (N_2385,N_2135,N_2134);
or U2386 (N_2386,N_2132,N_2029);
and U2387 (N_2387,N_2132,N_2109);
nor U2388 (N_2388,N_2138,N_2038);
xor U2389 (N_2389,N_2197,N_2034);
and U2390 (N_2390,N_2192,N_2186);
and U2391 (N_2391,N_2048,N_2049);
nor U2392 (N_2392,N_2186,N_2197);
and U2393 (N_2393,N_2134,N_2094);
nor U2394 (N_2394,N_2058,N_2042);
nor U2395 (N_2395,N_2133,N_2007);
and U2396 (N_2396,N_2136,N_2079);
and U2397 (N_2397,N_2105,N_2172);
or U2398 (N_2398,N_2118,N_2095);
nor U2399 (N_2399,N_2056,N_2044);
xor U2400 (N_2400,N_2273,N_2245);
or U2401 (N_2401,N_2352,N_2247);
nor U2402 (N_2402,N_2292,N_2279);
nand U2403 (N_2403,N_2232,N_2394);
nand U2404 (N_2404,N_2288,N_2264);
nor U2405 (N_2405,N_2240,N_2252);
nor U2406 (N_2406,N_2384,N_2363);
nor U2407 (N_2407,N_2333,N_2297);
and U2408 (N_2408,N_2319,N_2393);
nor U2409 (N_2409,N_2275,N_2258);
or U2410 (N_2410,N_2312,N_2294);
nand U2411 (N_2411,N_2299,N_2260);
or U2412 (N_2412,N_2224,N_2242);
and U2413 (N_2413,N_2385,N_2296);
or U2414 (N_2414,N_2381,N_2308);
nor U2415 (N_2415,N_2383,N_2391);
or U2416 (N_2416,N_2227,N_2338);
and U2417 (N_2417,N_2217,N_2213);
and U2418 (N_2418,N_2397,N_2379);
nand U2419 (N_2419,N_2238,N_2348);
and U2420 (N_2420,N_2358,N_2257);
xnor U2421 (N_2421,N_2298,N_2289);
nand U2422 (N_2422,N_2216,N_2321);
nand U2423 (N_2423,N_2337,N_2351);
or U2424 (N_2424,N_2377,N_2225);
and U2425 (N_2425,N_2203,N_2277);
nor U2426 (N_2426,N_2331,N_2369);
and U2427 (N_2427,N_2340,N_2345);
xnor U2428 (N_2428,N_2235,N_2282);
nand U2429 (N_2429,N_2211,N_2218);
or U2430 (N_2430,N_2353,N_2220);
nor U2431 (N_2431,N_2243,N_2311);
nor U2432 (N_2432,N_2278,N_2214);
nand U2433 (N_2433,N_2293,N_2269);
xnor U2434 (N_2434,N_2259,N_2303);
and U2435 (N_2435,N_2274,N_2263);
and U2436 (N_2436,N_2389,N_2283);
or U2437 (N_2437,N_2329,N_2230);
nand U2438 (N_2438,N_2241,N_2309);
and U2439 (N_2439,N_2368,N_2370);
nor U2440 (N_2440,N_2207,N_2209);
nor U2441 (N_2441,N_2271,N_2254);
xnor U2442 (N_2442,N_2356,N_2205);
or U2443 (N_2443,N_2307,N_2326);
or U2444 (N_2444,N_2251,N_2380);
nor U2445 (N_2445,N_2323,N_2372);
nand U2446 (N_2446,N_2202,N_2320);
or U2447 (N_2447,N_2272,N_2302);
nand U2448 (N_2448,N_2233,N_2374);
or U2449 (N_2449,N_2346,N_2316);
nand U2450 (N_2450,N_2362,N_2342);
nor U2451 (N_2451,N_2206,N_2276);
xnor U2452 (N_2452,N_2317,N_2215);
xnor U2453 (N_2453,N_2244,N_2250);
and U2454 (N_2454,N_2341,N_2328);
and U2455 (N_2455,N_2366,N_2344);
nor U2456 (N_2456,N_2304,N_2210);
nand U2457 (N_2457,N_2390,N_2228);
or U2458 (N_2458,N_2246,N_2367);
or U2459 (N_2459,N_2253,N_2359);
and U2460 (N_2460,N_2334,N_2347);
or U2461 (N_2461,N_2315,N_2221);
or U2462 (N_2462,N_2229,N_2350);
nand U2463 (N_2463,N_2286,N_2261);
nand U2464 (N_2464,N_2285,N_2236);
nor U2465 (N_2465,N_2310,N_2332);
nand U2466 (N_2466,N_2318,N_2399);
xnor U2467 (N_2467,N_2270,N_2314);
nand U2468 (N_2468,N_2212,N_2290);
nor U2469 (N_2469,N_2256,N_2313);
nor U2470 (N_2470,N_2339,N_2291);
xnor U2471 (N_2471,N_2208,N_2200);
nor U2472 (N_2472,N_2231,N_2357);
and U2473 (N_2473,N_2300,N_2262);
nor U2474 (N_2474,N_2284,N_2239);
nor U2475 (N_2475,N_2325,N_2219);
xnor U2476 (N_2476,N_2223,N_2201);
nand U2477 (N_2477,N_2398,N_2226);
or U2478 (N_2478,N_2361,N_2255);
xor U2479 (N_2479,N_2249,N_2281);
nand U2480 (N_2480,N_2355,N_2267);
and U2481 (N_2481,N_2301,N_2360);
or U2482 (N_2482,N_2378,N_2382);
or U2483 (N_2483,N_2222,N_2327);
and U2484 (N_2484,N_2396,N_2266);
nor U2485 (N_2485,N_2386,N_2324);
nand U2486 (N_2486,N_2204,N_2354);
or U2487 (N_2487,N_2237,N_2306);
or U2488 (N_2488,N_2280,N_2388);
nand U2489 (N_2489,N_2395,N_2373);
and U2490 (N_2490,N_2248,N_2265);
xor U2491 (N_2491,N_2387,N_2322);
and U2492 (N_2492,N_2371,N_2295);
nor U2493 (N_2493,N_2392,N_2268);
nand U2494 (N_2494,N_2335,N_2343);
or U2495 (N_2495,N_2305,N_2364);
and U2496 (N_2496,N_2336,N_2349);
nand U2497 (N_2497,N_2365,N_2375);
and U2498 (N_2498,N_2376,N_2234);
or U2499 (N_2499,N_2330,N_2287);
nand U2500 (N_2500,N_2256,N_2263);
xnor U2501 (N_2501,N_2393,N_2398);
xnor U2502 (N_2502,N_2398,N_2209);
and U2503 (N_2503,N_2200,N_2210);
xor U2504 (N_2504,N_2352,N_2378);
or U2505 (N_2505,N_2215,N_2309);
xor U2506 (N_2506,N_2215,N_2224);
or U2507 (N_2507,N_2268,N_2366);
xnor U2508 (N_2508,N_2231,N_2254);
nand U2509 (N_2509,N_2338,N_2262);
xnor U2510 (N_2510,N_2356,N_2354);
and U2511 (N_2511,N_2259,N_2261);
nor U2512 (N_2512,N_2337,N_2367);
xnor U2513 (N_2513,N_2272,N_2390);
nand U2514 (N_2514,N_2349,N_2296);
nor U2515 (N_2515,N_2348,N_2343);
nor U2516 (N_2516,N_2334,N_2212);
and U2517 (N_2517,N_2260,N_2361);
nand U2518 (N_2518,N_2344,N_2393);
or U2519 (N_2519,N_2384,N_2299);
nand U2520 (N_2520,N_2256,N_2288);
and U2521 (N_2521,N_2349,N_2253);
nor U2522 (N_2522,N_2336,N_2318);
and U2523 (N_2523,N_2326,N_2342);
nand U2524 (N_2524,N_2275,N_2221);
nor U2525 (N_2525,N_2386,N_2399);
nor U2526 (N_2526,N_2349,N_2208);
or U2527 (N_2527,N_2351,N_2330);
nand U2528 (N_2528,N_2289,N_2264);
xnor U2529 (N_2529,N_2263,N_2251);
xnor U2530 (N_2530,N_2381,N_2208);
or U2531 (N_2531,N_2314,N_2219);
and U2532 (N_2532,N_2363,N_2245);
and U2533 (N_2533,N_2308,N_2341);
nand U2534 (N_2534,N_2312,N_2246);
nand U2535 (N_2535,N_2280,N_2290);
nand U2536 (N_2536,N_2303,N_2287);
xor U2537 (N_2537,N_2385,N_2321);
nor U2538 (N_2538,N_2317,N_2298);
or U2539 (N_2539,N_2354,N_2289);
xor U2540 (N_2540,N_2359,N_2265);
nand U2541 (N_2541,N_2238,N_2373);
nand U2542 (N_2542,N_2302,N_2374);
nor U2543 (N_2543,N_2275,N_2316);
or U2544 (N_2544,N_2229,N_2381);
nor U2545 (N_2545,N_2219,N_2383);
nand U2546 (N_2546,N_2367,N_2208);
nand U2547 (N_2547,N_2256,N_2225);
nor U2548 (N_2548,N_2275,N_2280);
or U2549 (N_2549,N_2228,N_2331);
nor U2550 (N_2550,N_2224,N_2252);
or U2551 (N_2551,N_2206,N_2251);
nand U2552 (N_2552,N_2337,N_2399);
or U2553 (N_2553,N_2332,N_2205);
nor U2554 (N_2554,N_2217,N_2291);
or U2555 (N_2555,N_2396,N_2363);
and U2556 (N_2556,N_2225,N_2217);
nand U2557 (N_2557,N_2340,N_2207);
xnor U2558 (N_2558,N_2268,N_2341);
or U2559 (N_2559,N_2381,N_2385);
nor U2560 (N_2560,N_2230,N_2377);
nor U2561 (N_2561,N_2204,N_2324);
or U2562 (N_2562,N_2296,N_2204);
or U2563 (N_2563,N_2303,N_2227);
and U2564 (N_2564,N_2344,N_2376);
or U2565 (N_2565,N_2368,N_2394);
nor U2566 (N_2566,N_2223,N_2232);
nor U2567 (N_2567,N_2237,N_2228);
or U2568 (N_2568,N_2280,N_2282);
or U2569 (N_2569,N_2315,N_2334);
nand U2570 (N_2570,N_2237,N_2236);
nand U2571 (N_2571,N_2264,N_2307);
nor U2572 (N_2572,N_2376,N_2359);
nor U2573 (N_2573,N_2218,N_2246);
nor U2574 (N_2574,N_2387,N_2240);
or U2575 (N_2575,N_2244,N_2337);
nor U2576 (N_2576,N_2227,N_2378);
and U2577 (N_2577,N_2313,N_2355);
or U2578 (N_2578,N_2332,N_2299);
or U2579 (N_2579,N_2226,N_2242);
nand U2580 (N_2580,N_2357,N_2305);
nand U2581 (N_2581,N_2386,N_2218);
or U2582 (N_2582,N_2332,N_2295);
or U2583 (N_2583,N_2278,N_2395);
and U2584 (N_2584,N_2355,N_2218);
or U2585 (N_2585,N_2369,N_2353);
and U2586 (N_2586,N_2235,N_2391);
nor U2587 (N_2587,N_2375,N_2226);
and U2588 (N_2588,N_2277,N_2208);
or U2589 (N_2589,N_2366,N_2220);
nor U2590 (N_2590,N_2277,N_2252);
and U2591 (N_2591,N_2387,N_2262);
nand U2592 (N_2592,N_2210,N_2353);
nand U2593 (N_2593,N_2303,N_2256);
nand U2594 (N_2594,N_2319,N_2238);
nor U2595 (N_2595,N_2240,N_2293);
nor U2596 (N_2596,N_2220,N_2330);
or U2597 (N_2597,N_2251,N_2365);
nand U2598 (N_2598,N_2322,N_2382);
and U2599 (N_2599,N_2285,N_2362);
and U2600 (N_2600,N_2483,N_2414);
xor U2601 (N_2601,N_2441,N_2401);
xnor U2602 (N_2602,N_2436,N_2474);
or U2603 (N_2603,N_2548,N_2428);
xnor U2604 (N_2604,N_2422,N_2449);
and U2605 (N_2605,N_2546,N_2582);
nand U2606 (N_2606,N_2453,N_2400);
nor U2607 (N_2607,N_2542,N_2520);
nand U2608 (N_2608,N_2413,N_2557);
nor U2609 (N_2609,N_2438,N_2465);
xnor U2610 (N_2610,N_2549,N_2540);
nor U2611 (N_2611,N_2530,N_2518);
or U2612 (N_2612,N_2470,N_2408);
nand U2613 (N_2613,N_2425,N_2497);
nor U2614 (N_2614,N_2507,N_2416);
xor U2615 (N_2615,N_2552,N_2502);
and U2616 (N_2616,N_2519,N_2473);
and U2617 (N_2617,N_2471,N_2469);
nor U2618 (N_2618,N_2431,N_2543);
nor U2619 (N_2619,N_2529,N_2409);
and U2620 (N_2620,N_2435,N_2440);
or U2621 (N_2621,N_2587,N_2584);
nor U2622 (N_2622,N_2464,N_2411);
nor U2623 (N_2623,N_2484,N_2446);
and U2624 (N_2624,N_2573,N_2420);
and U2625 (N_2625,N_2568,N_2515);
and U2626 (N_2626,N_2439,N_2569);
xnor U2627 (N_2627,N_2472,N_2514);
or U2628 (N_2628,N_2496,N_2426);
nor U2629 (N_2629,N_2545,N_2579);
nor U2630 (N_2630,N_2551,N_2555);
nor U2631 (N_2631,N_2479,N_2506);
and U2632 (N_2632,N_2585,N_2434);
nand U2633 (N_2633,N_2563,N_2537);
nand U2634 (N_2634,N_2457,N_2522);
nand U2635 (N_2635,N_2583,N_2580);
and U2636 (N_2636,N_2547,N_2432);
or U2637 (N_2637,N_2565,N_2419);
nor U2638 (N_2638,N_2480,N_2450);
and U2639 (N_2639,N_2593,N_2445);
or U2640 (N_2640,N_2444,N_2533);
nand U2641 (N_2641,N_2576,N_2499);
nand U2642 (N_2642,N_2427,N_2481);
and U2643 (N_2643,N_2487,N_2406);
nor U2644 (N_2644,N_2458,N_2577);
and U2645 (N_2645,N_2451,N_2417);
or U2646 (N_2646,N_2594,N_2571);
nor U2647 (N_2647,N_2508,N_2477);
nor U2648 (N_2648,N_2410,N_2491);
nor U2649 (N_2649,N_2558,N_2505);
or U2650 (N_2650,N_2561,N_2556);
nor U2651 (N_2651,N_2592,N_2448);
nand U2652 (N_2652,N_2504,N_2463);
and U2653 (N_2653,N_2534,N_2415);
nor U2654 (N_2654,N_2482,N_2589);
nor U2655 (N_2655,N_2509,N_2452);
nand U2656 (N_2656,N_2586,N_2575);
nor U2657 (N_2657,N_2488,N_2468);
nor U2658 (N_2658,N_2424,N_2437);
nand U2659 (N_2659,N_2403,N_2532);
and U2660 (N_2660,N_2566,N_2429);
nand U2661 (N_2661,N_2466,N_2503);
nor U2662 (N_2662,N_2538,N_2500);
and U2663 (N_2663,N_2524,N_2486);
nand U2664 (N_2664,N_2531,N_2559);
nor U2665 (N_2665,N_2536,N_2567);
nor U2666 (N_2666,N_2513,N_2490);
or U2667 (N_2667,N_2418,N_2516);
nor U2668 (N_2668,N_2478,N_2599);
nor U2669 (N_2669,N_2517,N_2544);
and U2670 (N_2670,N_2562,N_2535);
nand U2671 (N_2671,N_2595,N_2447);
and U2672 (N_2672,N_2404,N_2527);
nand U2673 (N_2673,N_2495,N_2525);
nand U2674 (N_2674,N_2476,N_2412);
nor U2675 (N_2675,N_2421,N_2407);
nand U2676 (N_2676,N_2493,N_2402);
nand U2677 (N_2677,N_2581,N_2405);
xnor U2678 (N_2678,N_2523,N_2485);
nand U2679 (N_2679,N_2462,N_2494);
nand U2680 (N_2680,N_2430,N_2455);
nor U2681 (N_2681,N_2489,N_2591);
and U2682 (N_2682,N_2578,N_2572);
and U2683 (N_2683,N_2554,N_2596);
and U2684 (N_2684,N_2498,N_2443);
nand U2685 (N_2685,N_2521,N_2512);
and U2686 (N_2686,N_2433,N_2528);
nor U2687 (N_2687,N_2461,N_2539);
nand U2688 (N_2688,N_2442,N_2570);
or U2689 (N_2689,N_2564,N_2526);
nand U2690 (N_2690,N_2598,N_2574);
nand U2691 (N_2691,N_2560,N_2511);
and U2692 (N_2692,N_2501,N_2423);
nor U2693 (N_2693,N_2460,N_2454);
and U2694 (N_2694,N_2475,N_2467);
nand U2695 (N_2695,N_2588,N_2541);
and U2696 (N_2696,N_2550,N_2456);
nor U2697 (N_2697,N_2597,N_2459);
nor U2698 (N_2698,N_2492,N_2590);
nand U2699 (N_2699,N_2553,N_2510);
or U2700 (N_2700,N_2599,N_2428);
nand U2701 (N_2701,N_2541,N_2522);
or U2702 (N_2702,N_2475,N_2447);
nor U2703 (N_2703,N_2425,N_2554);
nor U2704 (N_2704,N_2472,N_2569);
or U2705 (N_2705,N_2409,N_2559);
nor U2706 (N_2706,N_2420,N_2597);
nor U2707 (N_2707,N_2417,N_2478);
xnor U2708 (N_2708,N_2446,N_2536);
xnor U2709 (N_2709,N_2526,N_2420);
xor U2710 (N_2710,N_2538,N_2527);
nor U2711 (N_2711,N_2559,N_2404);
xnor U2712 (N_2712,N_2541,N_2447);
or U2713 (N_2713,N_2579,N_2524);
nand U2714 (N_2714,N_2477,N_2500);
or U2715 (N_2715,N_2465,N_2480);
or U2716 (N_2716,N_2557,N_2409);
or U2717 (N_2717,N_2406,N_2497);
nand U2718 (N_2718,N_2575,N_2478);
nor U2719 (N_2719,N_2556,N_2432);
or U2720 (N_2720,N_2583,N_2414);
and U2721 (N_2721,N_2541,N_2436);
nand U2722 (N_2722,N_2462,N_2543);
or U2723 (N_2723,N_2550,N_2580);
nor U2724 (N_2724,N_2444,N_2436);
or U2725 (N_2725,N_2557,N_2554);
and U2726 (N_2726,N_2549,N_2515);
or U2727 (N_2727,N_2435,N_2472);
or U2728 (N_2728,N_2487,N_2426);
and U2729 (N_2729,N_2492,N_2403);
xnor U2730 (N_2730,N_2545,N_2416);
xnor U2731 (N_2731,N_2497,N_2507);
xor U2732 (N_2732,N_2519,N_2444);
nor U2733 (N_2733,N_2521,N_2590);
nor U2734 (N_2734,N_2562,N_2419);
xor U2735 (N_2735,N_2543,N_2495);
nor U2736 (N_2736,N_2445,N_2503);
xor U2737 (N_2737,N_2591,N_2534);
or U2738 (N_2738,N_2431,N_2467);
or U2739 (N_2739,N_2504,N_2488);
and U2740 (N_2740,N_2431,N_2583);
and U2741 (N_2741,N_2548,N_2577);
or U2742 (N_2742,N_2477,N_2545);
nand U2743 (N_2743,N_2544,N_2558);
and U2744 (N_2744,N_2441,N_2413);
or U2745 (N_2745,N_2537,N_2492);
and U2746 (N_2746,N_2443,N_2430);
and U2747 (N_2747,N_2418,N_2508);
and U2748 (N_2748,N_2456,N_2521);
and U2749 (N_2749,N_2524,N_2569);
nor U2750 (N_2750,N_2448,N_2430);
and U2751 (N_2751,N_2584,N_2506);
nor U2752 (N_2752,N_2589,N_2407);
or U2753 (N_2753,N_2472,N_2545);
or U2754 (N_2754,N_2407,N_2543);
nand U2755 (N_2755,N_2462,N_2402);
and U2756 (N_2756,N_2427,N_2417);
or U2757 (N_2757,N_2578,N_2573);
nor U2758 (N_2758,N_2484,N_2482);
and U2759 (N_2759,N_2480,N_2429);
and U2760 (N_2760,N_2409,N_2598);
nand U2761 (N_2761,N_2524,N_2592);
nand U2762 (N_2762,N_2428,N_2521);
or U2763 (N_2763,N_2472,N_2542);
or U2764 (N_2764,N_2472,N_2457);
nor U2765 (N_2765,N_2426,N_2400);
xor U2766 (N_2766,N_2466,N_2474);
or U2767 (N_2767,N_2523,N_2505);
nor U2768 (N_2768,N_2448,N_2485);
nor U2769 (N_2769,N_2455,N_2463);
or U2770 (N_2770,N_2562,N_2472);
nor U2771 (N_2771,N_2578,N_2550);
nor U2772 (N_2772,N_2440,N_2593);
nand U2773 (N_2773,N_2470,N_2461);
or U2774 (N_2774,N_2409,N_2405);
or U2775 (N_2775,N_2423,N_2499);
or U2776 (N_2776,N_2583,N_2401);
or U2777 (N_2777,N_2454,N_2499);
and U2778 (N_2778,N_2465,N_2470);
nand U2779 (N_2779,N_2517,N_2531);
nor U2780 (N_2780,N_2558,N_2589);
xor U2781 (N_2781,N_2492,N_2478);
or U2782 (N_2782,N_2403,N_2432);
and U2783 (N_2783,N_2534,N_2562);
or U2784 (N_2784,N_2429,N_2575);
xnor U2785 (N_2785,N_2564,N_2587);
or U2786 (N_2786,N_2413,N_2454);
nand U2787 (N_2787,N_2579,N_2448);
or U2788 (N_2788,N_2510,N_2494);
xor U2789 (N_2789,N_2498,N_2584);
and U2790 (N_2790,N_2503,N_2590);
or U2791 (N_2791,N_2438,N_2569);
or U2792 (N_2792,N_2584,N_2495);
nor U2793 (N_2793,N_2556,N_2510);
or U2794 (N_2794,N_2533,N_2500);
nor U2795 (N_2795,N_2501,N_2470);
nor U2796 (N_2796,N_2471,N_2542);
xnor U2797 (N_2797,N_2436,N_2489);
and U2798 (N_2798,N_2578,N_2592);
and U2799 (N_2799,N_2500,N_2455);
xnor U2800 (N_2800,N_2758,N_2662);
xor U2801 (N_2801,N_2722,N_2693);
and U2802 (N_2802,N_2659,N_2733);
and U2803 (N_2803,N_2633,N_2764);
or U2804 (N_2804,N_2717,N_2670);
xor U2805 (N_2805,N_2695,N_2635);
and U2806 (N_2806,N_2634,N_2753);
xnor U2807 (N_2807,N_2624,N_2643);
nand U2808 (N_2808,N_2611,N_2734);
and U2809 (N_2809,N_2649,N_2678);
or U2810 (N_2810,N_2770,N_2762);
nor U2811 (N_2811,N_2781,N_2682);
and U2812 (N_2812,N_2653,N_2701);
or U2813 (N_2813,N_2656,N_2631);
nand U2814 (N_2814,N_2752,N_2616);
xor U2815 (N_2815,N_2772,N_2789);
or U2816 (N_2816,N_2606,N_2680);
nand U2817 (N_2817,N_2795,N_2687);
and U2818 (N_2818,N_2736,N_2663);
nor U2819 (N_2819,N_2709,N_2674);
or U2820 (N_2820,N_2614,N_2726);
nor U2821 (N_2821,N_2760,N_2676);
nand U2822 (N_2822,N_2765,N_2748);
or U2823 (N_2823,N_2655,N_2694);
nand U2824 (N_2824,N_2700,N_2637);
or U2825 (N_2825,N_2714,N_2690);
xnor U2826 (N_2826,N_2615,N_2608);
nor U2827 (N_2827,N_2605,N_2792);
nand U2828 (N_2828,N_2688,N_2739);
nand U2829 (N_2829,N_2667,N_2636);
or U2830 (N_2830,N_2738,N_2671);
or U2831 (N_2831,N_2706,N_2645);
nand U2832 (N_2832,N_2679,N_2602);
or U2833 (N_2833,N_2707,N_2669);
or U2834 (N_2834,N_2672,N_2740);
nand U2835 (N_2835,N_2697,N_2625);
and U2836 (N_2836,N_2704,N_2683);
and U2837 (N_2837,N_2673,N_2767);
nor U2838 (N_2838,N_2775,N_2730);
nor U2839 (N_2839,N_2743,N_2612);
or U2840 (N_2840,N_2621,N_2689);
and U2841 (N_2841,N_2696,N_2731);
and U2842 (N_2842,N_2619,N_2749);
nor U2843 (N_2843,N_2661,N_2677);
nand U2844 (N_2844,N_2725,N_2604);
xnor U2845 (N_2845,N_2627,N_2600);
or U2846 (N_2846,N_2703,N_2620);
and U2847 (N_2847,N_2640,N_2675);
nor U2848 (N_2848,N_2724,N_2638);
nor U2849 (N_2849,N_2757,N_2771);
nor U2850 (N_2850,N_2729,N_2745);
nand U2851 (N_2851,N_2681,N_2668);
nor U2852 (N_2852,N_2756,N_2723);
nor U2853 (N_2853,N_2735,N_2618);
and U2854 (N_2854,N_2647,N_2708);
nand U2855 (N_2855,N_2776,N_2773);
nand U2856 (N_2856,N_2794,N_2732);
nor U2857 (N_2857,N_2641,N_2780);
and U2858 (N_2858,N_2737,N_2657);
or U2859 (N_2859,N_2711,N_2744);
xor U2860 (N_2860,N_2742,N_2755);
nand U2861 (N_2861,N_2665,N_2710);
nand U2862 (N_2862,N_2763,N_2769);
and U2863 (N_2863,N_2651,N_2774);
nor U2864 (N_2864,N_2713,N_2629);
nor U2865 (N_2865,N_2628,N_2796);
and U2866 (N_2866,N_2626,N_2718);
nand U2867 (N_2867,N_2652,N_2685);
or U2868 (N_2868,N_2728,N_2658);
nor U2869 (N_2869,N_2632,N_2650);
and U2870 (N_2870,N_2784,N_2759);
or U2871 (N_2871,N_2721,N_2746);
xor U2872 (N_2872,N_2747,N_2610);
nor U2873 (N_2873,N_2798,N_2720);
nor U2874 (N_2874,N_2654,N_2754);
or U2875 (N_2875,N_2768,N_2786);
nand U2876 (N_2876,N_2719,N_2686);
nor U2877 (N_2877,N_2785,N_2639);
nand U2878 (N_2878,N_2666,N_2727);
or U2879 (N_2879,N_2630,N_2761);
or U2880 (N_2880,N_2705,N_2788);
nor U2881 (N_2881,N_2623,N_2692);
or U2882 (N_2882,N_2751,N_2698);
nor U2883 (N_2883,N_2793,N_2715);
nand U2884 (N_2884,N_2648,N_2787);
nor U2885 (N_2885,N_2609,N_2684);
or U2886 (N_2886,N_2642,N_2782);
nor U2887 (N_2887,N_2699,N_2601);
xnor U2888 (N_2888,N_2777,N_2617);
nor U2889 (N_2889,N_2741,N_2778);
and U2890 (N_2890,N_2791,N_2660);
or U2891 (N_2891,N_2644,N_2766);
nor U2892 (N_2892,N_2750,N_2607);
or U2893 (N_2893,N_2799,N_2613);
or U2894 (N_2894,N_2691,N_2622);
and U2895 (N_2895,N_2779,N_2646);
nand U2896 (N_2896,N_2797,N_2790);
or U2897 (N_2897,N_2702,N_2664);
nand U2898 (N_2898,N_2712,N_2603);
and U2899 (N_2899,N_2783,N_2716);
and U2900 (N_2900,N_2740,N_2645);
xor U2901 (N_2901,N_2691,N_2791);
nand U2902 (N_2902,N_2631,N_2753);
nand U2903 (N_2903,N_2699,N_2736);
nor U2904 (N_2904,N_2709,N_2761);
nor U2905 (N_2905,N_2668,N_2674);
nor U2906 (N_2906,N_2739,N_2620);
or U2907 (N_2907,N_2751,N_2770);
or U2908 (N_2908,N_2784,N_2799);
and U2909 (N_2909,N_2675,N_2776);
nand U2910 (N_2910,N_2674,N_2630);
nor U2911 (N_2911,N_2640,N_2747);
nand U2912 (N_2912,N_2729,N_2670);
nand U2913 (N_2913,N_2776,N_2625);
nand U2914 (N_2914,N_2702,N_2619);
xor U2915 (N_2915,N_2728,N_2741);
and U2916 (N_2916,N_2690,N_2646);
nor U2917 (N_2917,N_2726,N_2664);
and U2918 (N_2918,N_2770,N_2760);
and U2919 (N_2919,N_2754,N_2756);
nor U2920 (N_2920,N_2609,N_2686);
xnor U2921 (N_2921,N_2676,N_2700);
nand U2922 (N_2922,N_2671,N_2767);
nor U2923 (N_2923,N_2724,N_2646);
and U2924 (N_2924,N_2602,N_2731);
nand U2925 (N_2925,N_2675,N_2656);
and U2926 (N_2926,N_2654,N_2651);
or U2927 (N_2927,N_2636,N_2732);
or U2928 (N_2928,N_2610,N_2654);
or U2929 (N_2929,N_2672,N_2749);
nand U2930 (N_2930,N_2698,N_2690);
nor U2931 (N_2931,N_2638,N_2673);
or U2932 (N_2932,N_2767,N_2781);
and U2933 (N_2933,N_2711,N_2777);
or U2934 (N_2934,N_2714,N_2796);
and U2935 (N_2935,N_2694,N_2717);
and U2936 (N_2936,N_2705,N_2645);
and U2937 (N_2937,N_2644,N_2671);
nand U2938 (N_2938,N_2628,N_2635);
and U2939 (N_2939,N_2704,N_2715);
and U2940 (N_2940,N_2682,N_2630);
and U2941 (N_2941,N_2640,N_2650);
nor U2942 (N_2942,N_2670,N_2740);
nor U2943 (N_2943,N_2767,N_2736);
xor U2944 (N_2944,N_2654,N_2717);
and U2945 (N_2945,N_2636,N_2615);
nor U2946 (N_2946,N_2685,N_2785);
and U2947 (N_2947,N_2777,N_2610);
nand U2948 (N_2948,N_2682,N_2754);
or U2949 (N_2949,N_2616,N_2759);
nor U2950 (N_2950,N_2678,N_2603);
nand U2951 (N_2951,N_2746,N_2674);
and U2952 (N_2952,N_2658,N_2746);
and U2953 (N_2953,N_2727,N_2661);
nand U2954 (N_2954,N_2687,N_2682);
xor U2955 (N_2955,N_2719,N_2706);
nand U2956 (N_2956,N_2791,N_2681);
nand U2957 (N_2957,N_2745,N_2728);
nor U2958 (N_2958,N_2625,N_2742);
and U2959 (N_2959,N_2747,N_2647);
nor U2960 (N_2960,N_2678,N_2783);
nand U2961 (N_2961,N_2627,N_2781);
nor U2962 (N_2962,N_2724,N_2671);
nor U2963 (N_2963,N_2750,N_2673);
and U2964 (N_2964,N_2607,N_2743);
xor U2965 (N_2965,N_2710,N_2655);
and U2966 (N_2966,N_2618,N_2725);
or U2967 (N_2967,N_2690,N_2668);
nand U2968 (N_2968,N_2714,N_2657);
nor U2969 (N_2969,N_2768,N_2602);
and U2970 (N_2970,N_2637,N_2738);
or U2971 (N_2971,N_2799,N_2682);
nand U2972 (N_2972,N_2726,N_2777);
nor U2973 (N_2973,N_2733,N_2637);
or U2974 (N_2974,N_2769,N_2745);
xor U2975 (N_2975,N_2670,N_2644);
and U2976 (N_2976,N_2704,N_2649);
nor U2977 (N_2977,N_2638,N_2642);
nand U2978 (N_2978,N_2765,N_2650);
or U2979 (N_2979,N_2657,N_2705);
or U2980 (N_2980,N_2790,N_2686);
nor U2981 (N_2981,N_2654,N_2608);
and U2982 (N_2982,N_2747,N_2769);
or U2983 (N_2983,N_2717,N_2737);
nand U2984 (N_2984,N_2698,N_2713);
and U2985 (N_2985,N_2785,N_2753);
nor U2986 (N_2986,N_2717,N_2691);
and U2987 (N_2987,N_2749,N_2700);
nor U2988 (N_2988,N_2633,N_2783);
and U2989 (N_2989,N_2622,N_2627);
nor U2990 (N_2990,N_2660,N_2790);
or U2991 (N_2991,N_2738,N_2717);
nor U2992 (N_2992,N_2741,N_2615);
nor U2993 (N_2993,N_2606,N_2676);
nand U2994 (N_2994,N_2735,N_2663);
nand U2995 (N_2995,N_2764,N_2695);
or U2996 (N_2996,N_2722,N_2708);
nor U2997 (N_2997,N_2713,N_2686);
or U2998 (N_2998,N_2766,N_2742);
and U2999 (N_2999,N_2621,N_2704);
and U3000 (N_3000,N_2858,N_2982);
nand U3001 (N_3001,N_2821,N_2867);
or U3002 (N_3002,N_2979,N_2899);
and U3003 (N_3003,N_2803,N_2960);
nor U3004 (N_3004,N_2835,N_2871);
or U3005 (N_3005,N_2817,N_2865);
nor U3006 (N_3006,N_2988,N_2903);
xnor U3007 (N_3007,N_2869,N_2838);
or U3008 (N_3008,N_2964,N_2857);
nor U3009 (N_3009,N_2890,N_2894);
or U3010 (N_3010,N_2965,N_2834);
or U3011 (N_3011,N_2991,N_2856);
and U3012 (N_3012,N_2936,N_2874);
xnor U3013 (N_3013,N_2848,N_2962);
nand U3014 (N_3014,N_2901,N_2978);
nor U3015 (N_3015,N_2843,N_2918);
nand U3016 (N_3016,N_2981,N_2908);
xnor U3017 (N_3017,N_2854,N_2833);
xnor U3018 (N_3018,N_2912,N_2888);
or U3019 (N_3019,N_2829,N_2887);
nor U3020 (N_3020,N_2975,N_2992);
nand U3021 (N_3021,N_2997,N_2845);
nand U3022 (N_3022,N_2976,N_2818);
nand U3023 (N_3023,N_2961,N_2813);
and U3024 (N_3024,N_2830,N_2985);
nor U3025 (N_3025,N_2973,N_2996);
or U3026 (N_3026,N_2836,N_2823);
nor U3027 (N_3027,N_2900,N_2902);
nor U3028 (N_3028,N_2863,N_2841);
and U3029 (N_3029,N_2827,N_2941);
and U3030 (N_3030,N_2950,N_2926);
nand U3031 (N_3031,N_2876,N_2947);
and U3032 (N_3032,N_2882,N_2907);
or U3033 (N_3033,N_2989,N_2939);
and U3034 (N_3034,N_2970,N_2972);
xor U3035 (N_3035,N_2878,N_2967);
or U3036 (N_3036,N_2873,N_2940);
and U3037 (N_3037,N_2971,N_2849);
or U3038 (N_3038,N_2969,N_2955);
and U3039 (N_3039,N_2993,N_2855);
or U3040 (N_3040,N_2910,N_2828);
nor U3041 (N_3041,N_2801,N_2884);
or U3042 (N_3042,N_2898,N_2889);
and U3043 (N_3043,N_2806,N_2850);
xnor U3044 (N_3044,N_2933,N_2897);
and U3045 (N_3045,N_2915,N_2824);
nor U3046 (N_3046,N_2914,N_2994);
and U3047 (N_3047,N_2942,N_2859);
or U3048 (N_3048,N_2956,N_2814);
nand U3049 (N_3049,N_2820,N_2802);
and U3050 (N_3050,N_2983,N_2919);
nor U3051 (N_3051,N_2846,N_2911);
and U3052 (N_3052,N_2864,N_2847);
and U3053 (N_3053,N_2966,N_2822);
nand U3054 (N_3054,N_2987,N_2990);
or U3055 (N_3055,N_2935,N_2922);
nor U3056 (N_3056,N_2812,N_2826);
or U3057 (N_3057,N_2881,N_2963);
nand U3058 (N_3058,N_2905,N_2807);
nor U3059 (N_3059,N_2825,N_2862);
and U3060 (N_3060,N_2938,N_2808);
and U3061 (N_3061,N_2923,N_2877);
and U3062 (N_3062,N_2949,N_2954);
and U3063 (N_3063,N_2952,N_2944);
nand U3064 (N_3064,N_2892,N_2931);
and U3065 (N_3065,N_2895,N_2872);
xnor U3066 (N_3066,N_2932,N_2831);
xnor U3067 (N_3067,N_2948,N_2909);
or U3068 (N_3068,N_2860,N_2883);
and U3069 (N_3069,N_2800,N_2880);
or U3070 (N_3070,N_2832,N_2861);
and U3071 (N_3071,N_2946,N_2925);
and U3072 (N_3072,N_2842,N_2930);
or U3073 (N_3073,N_2998,N_2809);
and U3074 (N_3074,N_2886,N_2968);
or U3075 (N_3075,N_2891,N_2851);
and U3076 (N_3076,N_2805,N_2943);
and U3077 (N_3077,N_2945,N_2837);
nor U3078 (N_3078,N_2896,N_2819);
nor U3079 (N_3079,N_2866,N_2906);
or U3080 (N_3080,N_2974,N_2951);
nand U3081 (N_3081,N_2924,N_2893);
xnor U3082 (N_3082,N_2959,N_2999);
xnor U3083 (N_3083,N_2839,N_2852);
nor U3084 (N_3084,N_2885,N_2816);
or U3085 (N_3085,N_2958,N_2840);
or U3086 (N_3086,N_2875,N_2957);
nand U3087 (N_3087,N_2937,N_2904);
or U3088 (N_3088,N_2916,N_2804);
xor U3089 (N_3089,N_2980,N_2917);
xor U3090 (N_3090,N_2815,N_2853);
and U3091 (N_3091,N_2929,N_2986);
nand U3092 (N_3092,N_2920,N_2927);
or U3093 (N_3093,N_2953,N_2934);
nand U3094 (N_3094,N_2977,N_2870);
xnor U3095 (N_3095,N_2995,N_2913);
nand U3096 (N_3096,N_2868,N_2921);
and U3097 (N_3097,N_2984,N_2879);
or U3098 (N_3098,N_2844,N_2928);
and U3099 (N_3099,N_2811,N_2810);
and U3100 (N_3100,N_2985,N_2837);
and U3101 (N_3101,N_2943,N_2963);
and U3102 (N_3102,N_2982,N_2847);
or U3103 (N_3103,N_2942,N_2845);
nand U3104 (N_3104,N_2939,N_2964);
xnor U3105 (N_3105,N_2984,N_2918);
and U3106 (N_3106,N_2889,N_2974);
nor U3107 (N_3107,N_2957,N_2991);
nor U3108 (N_3108,N_2986,N_2827);
and U3109 (N_3109,N_2855,N_2915);
nor U3110 (N_3110,N_2962,N_2946);
nand U3111 (N_3111,N_2864,N_2804);
nor U3112 (N_3112,N_2922,N_2881);
nand U3113 (N_3113,N_2954,N_2881);
and U3114 (N_3114,N_2819,N_2818);
nor U3115 (N_3115,N_2868,N_2913);
and U3116 (N_3116,N_2906,N_2891);
nor U3117 (N_3117,N_2839,N_2973);
xnor U3118 (N_3118,N_2859,N_2827);
xnor U3119 (N_3119,N_2887,N_2922);
and U3120 (N_3120,N_2989,N_2913);
and U3121 (N_3121,N_2887,N_2999);
nor U3122 (N_3122,N_2971,N_2941);
nand U3123 (N_3123,N_2922,N_2940);
and U3124 (N_3124,N_2845,N_2861);
nand U3125 (N_3125,N_2898,N_2904);
and U3126 (N_3126,N_2926,N_2861);
nand U3127 (N_3127,N_2907,N_2889);
or U3128 (N_3128,N_2908,N_2891);
nor U3129 (N_3129,N_2876,N_2839);
nor U3130 (N_3130,N_2855,N_2999);
nor U3131 (N_3131,N_2937,N_2851);
nand U3132 (N_3132,N_2952,N_2862);
nor U3133 (N_3133,N_2882,N_2944);
nand U3134 (N_3134,N_2810,N_2973);
nor U3135 (N_3135,N_2994,N_2960);
xnor U3136 (N_3136,N_2839,N_2832);
nand U3137 (N_3137,N_2869,N_2999);
nor U3138 (N_3138,N_2892,N_2927);
or U3139 (N_3139,N_2952,N_2814);
nor U3140 (N_3140,N_2818,N_2901);
or U3141 (N_3141,N_2960,N_2868);
or U3142 (N_3142,N_2858,N_2846);
and U3143 (N_3143,N_2983,N_2950);
nand U3144 (N_3144,N_2928,N_2986);
nor U3145 (N_3145,N_2899,N_2822);
and U3146 (N_3146,N_2893,N_2956);
xnor U3147 (N_3147,N_2957,N_2931);
nor U3148 (N_3148,N_2911,N_2973);
xnor U3149 (N_3149,N_2957,N_2919);
nor U3150 (N_3150,N_2816,N_2937);
nand U3151 (N_3151,N_2858,N_2945);
and U3152 (N_3152,N_2922,N_2977);
nand U3153 (N_3153,N_2934,N_2833);
or U3154 (N_3154,N_2993,N_2863);
or U3155 (N_3155,N_2911,N_2951);
nor U3156 (N_3156,N_2893,N_2823);
and U3157 (N_3157,N_2920,N_2885);
nand U3158 (N_3158,N_2948,N_2912);
and U3159 (N_3159,N_2917,N_2860);
and U3160 (N_3160,N_2998,N_2847);
nand U3161 (N_3161,N_2832,N_2879);
nand U3162 (N_3162,N_2982,N_2869);
xor U3163 (N_3163,N_2972,N_2906);
nand U3164 (N_3164,N_2823,N_2946);
or U3165 (N_3165,N_2908,N_2804);
nand U3166 (N_3166,N_2953,N_2978);
and U3167 (N_3167,N_2889,N_2875);
or U3168 (N_3168,N_2957,N_2819);
or U3169 (N_3169,N_2902,N_2871);
and U3170 (N_3170,N_2900,N_2921);
and U3171 (N_3171,N_2853,N_2842);
nand U3172 (N_3172,N_2957,N_2900);
and U3173 (N_3173,N_2834,N_2814);
nand U3174 (N_3174,N_2829,N_2940);
or U3175 (N_3175,N_2979,N_2824);
and U3176 (N_3176,N_2904,N_2951);
or U3177 (N_3177,N_2926,N_2969);
nor U3178 (N_3178,N_2898,N_2942);
nor U3179 (N_3179,N_2920,N_2800);
xor U3180 (N_3180,N_2843,N_2926);
nand U3181 (N_3181,N_2895,N_2834);
or U3182 (N_3182,N_2807,N_2987);
nor U3183 (N_3183,N_2968,N_2805);
nor U3184 (N_3184,N_2850,N_2924);
nor U3185 (N_3185,N_2952,N_2926);
nand U3186 (N_3186,N_2928,N_2840);
nand U3187 (N_3187,N_2841,N_2800);
and U3188 (N_3188,N_2840,N_2993);
nor U3189 (N_3189,N_2884,N_2964);
nor U3190 (N_3190,N_2858,N_2864);
or U3191 (N_3191,N_2902,N_2808);
or U3192 (N_3192,N_2848,N_2911);
or U3193 (N_3193,N_2946,N_2945);
nor U3194 (N_3194,N_2828,N_2852);
and U3195 (N_3195,N_2950,N_2801);
xnor U3196 (N_3196,N_2853,N_2814);
and U3197 (N_3197,N_2836,N_2890);
or U3198 (N_3198,N_2966,N_2961);
nand U3199 (N_3199,N_2942,N_2862);
and U3200 (N_3200,N_3169,N_3150);
nand U3201 (N_3201,N_3052,N_3151);
or U3202 (N_3202,N_3030,N_3176);
nor U3203 (N_3203,N_3121,N_3028);
and U3204 (N_3204,N_3119,N_3088);
and U3205 (N_3205,N_3006,N_3011);
nand U3206 (N_3206,N_3120,N_3100);
and U3207 (N_3207,N_3079,N_3132);
and U3208 (N_3208,N_3089,N_3177);
and U3209 (N_3209,N_3145,N_3170);
or U3210 (N_3210,N_3020,N_3140);
nand U3211 (N_3211,N_3154,N_3174);
or U3212 (N_3212,N_3005,N_3083);
nand U3213 (N_3213,N_3070,N_3199);
xor U3214 (N_3214,N_3043,N_3185);
and U3215 (N_3215,N_3036,N_3061);
and U3216 (N_3216,N_3153,N_3110);
nor U3217 (N_3217,N_3179,N_3002);
and U3218 (N_3218,N_3197,N_3192);
nand U3219 (N_3219,N_3040,N_3095);
xor U3220 (N_3220,N_3064,N_3082);
or U3221 (N_3221,N_3125,N_3035);
nor U3222 (N_3222,N_3022,N_3039);
nand U3223 (N_3223,N_3105,N_3168);
nor U3224 (N_3224,N_3129,N_3034);
or U3225 (N_3225,N_3045,N_3114);
and U3226 (N_3226,N_3060,N_3056);
and U3227 (N_3227,N_3108,N_3144);
nand U3228 (N_3228,N_3147,N_3055);
xnor U3229 (N_3229,N_3081,N_3159);
nor U3230 (N_3230,N_3023,N_3024);
nor U3231 (N_3231,N_3071,N_3063);
xor U3232 (N_3232,N_3075,N_3085);
nand U3233 (N_3233,N_3026,N_3093);
nor U3234 (N_3234,N_3065,N_3086);
and U3235 (N_3235,N_3103,N_3098);
xnor U3236 (N_3236,N_3037,N_3092);
or U3237 (N_3237,N_3193,N_3091);
nand U3238 (N_3238,N_3090,N_3021);
and U3239 (N_3239,N_3104,N_3107);
or U3240 (N_3240,N_3112,N_3138);
xnor U3241 (N_3241,N_3115,N_3068);
xor U3242 (N_3242,N_3001,N_3111);
nand U3243 (N_3243,N_3102,N_3164);
and U3244 (N_3244,N_3166,N_3027);
xnor U3245 (N_3245,N_3155,N_3141);
xor U3246 (N_3246,N_3073,N_3015);
nand U3247 (N_3247,N_3069,N_3135);
and U3248 (N_3248,N_3188,N_3072);
and U3249 (N_3249,N_3186,N_3101);
or U3250 (N_3250,N_3167,N_3087);
and U3251 (N_3251,N_3181,N_3018);
nor U3252 (N_3252,N_3084,N_3156);
and U3253 (N_3253,N_3127,N_3117);
and U3254 (N_3254,N_3049,N_3126);
or U3255 (N_3255,N_3007,N_3157);
nor U3256 (N_3256,N_3050,N_3152);
nand U3257 (N_3257,N_3076,N_3031);
and U3258 (N_3258,N_3122,N_3017);
nor U3259 (N_3259,N_3053,N_3118);
and U3260 (N_3260,N_3146,N_3190);
and U3261 (N_3261,N_3080,N_3148);
nor U3262 (N_3262,N_3171,N_3124);
xnor U3263 (N_3263,N_3062,N_3183);
or U3264 (N_3264,N_3025,N_3175);
or U3265 (N_3265,N_3046,N_3184);
and U3266 (N_3266,N_3099,N_3149);
and U3267 (N_3267,N_3038,N_3191);
nor U3268 (N_3268,N_3010,N_3019);
nand U3269 (N_3269,N_3160,N_3042);
and U3270 (N_3270,N_3123,N_3033);
nand U3271 (N_3271,N_3077,N_3012);
xnor U3272 (N_3272,N_3016,N_3074);
nor U3273 (N_3273,N_3047,N_3158);
nand U3274 (N_3274,N_3182,N_3109);
xor U3275 (N_3275,N_3009,N_3032);
nand U3276 (N_3276,N_3162,N_3136);
nand U3277 (N_3277,N_3173,N_3097);
nor U3278 (N_3278,N_3134,N_3059);
nand U3279 (N_3279,N_3094,N_3044);
and U3280 (N_3280,N_3195,N_3066);
nand U3281 (N_3281,N_3058,N_3004);
or U3282 (N_3282,N_3051,N_3165);
nor U3283 (N_3283,N_3013,N_3196);
or U3284 (N_3284,N_3048,N_3130);
and U3285 (N_3285,N_3133,N_3172);
xnor U3286 (N_3286,N_3198,N_3189);
nor U3287 (N_3287,N_3161,N_3113);
and U3288 (N_3288,N_3128,N_3096);
nand U3289 (N_3289,N_3078,N_3180);
nand U3290 (N_3290,N_3057,N_3163);
nor U3291 (N_3291,N_3143,N_3194);
xnor U3292 (N_3292,N_3116,N_3187);
xor U3293 (N_3293,N_3178,N_3137);
or U3294 (N_3294,N_3000,N_3014);
nand U3295 (N_3295,N_3131,N_3139);
or U3296 (N_3296,N_3106,N_3041);
nor U3297 (N_3297,N_3054,N_3029);
nand U3298 (N_3298,N_3003,N_3067);
nor U3299 (N_3299,N_3142,N_3008);
and U3300 (N_3300,N_3151,N_3037);
nand U3301 (N_3301,N_3036,N_3157);
nor U3302 (N_3302,N_3077,N_3041);
and U3303 (N_3303,N_3045,N_3122);
nor U3304 (N_3304,N_3092,N_3086);
nand U3305 (N_3305,N_3074,N_3080);
or U3306 (N_3306,N_3144,N_3015);
xor U3307 (N_3307,N_3092,N_3169);
xor U3308 (N_3308,N_3026,N_3125);
nor U3309 (N_3309,N_3038,N_3124);
and U3310 (N_3310,N_3138,N_3027);
nor U3311 (N_3311,N_3021,N_3141);
and U3312 (N_3312,N_3101,N_3116);
nand U3313 (N_3313,N_3037,N_3181);
xnor U3314 (N_3314,N_3186,N_3100);
nor U3315 (N_3315,N_3165,N_3138);
or U3316 (N_3316,N_3021,N_3028);
or U3317 (N_3317,N_3044,N_3147);
nand U3318 (N_3318,N_3117,N_3071);
or U3319 (N_3319,N_3181,N_3020);
or U3320 (N_3320,N_3017,N_3185);
nand U3321 (N_3321,N_3016,N_3009);
nor U3322 (N_3322,N_3015,N_3027);
or U3323 (N_3323,N_3113,N_3003);
and U3324 (N_3324,N_3164,N_3107);
xnor U3325 (N_3325,N_3071,N_3180);
nand U3326 (N_3326,N_3064,N_3147);
xor U3327 (N_3327,N_3151,N_3064);
or U3328 (N_3328,N_3189,N_3169);
or U3329 (N_3329,N_3135,N_3043);
nand U3330 (N_3330,N_3117,N_3101);
nand U3331 (N_3331,N_3073,N_3064);
or U3332 (N_3332,N_3063,N_3123);
nand U3333 (N_3333,N_3122,N_3066);
nand U3334 (N_3334,N_3091,N_3130);
xnor U3335 (N_3335,N_3038,N_3128);
nand U3336 (N_3336,N_3009,N_3161);
and U3337 (N_3337,N_3094,N_3098);
nand U3338 (N_3338,N_3018,N_3082);
nand U3339 (N_3339,N_3174,N_3004);
nor U3340 (N_3340,N_3195,N_3002);
nor U3341 (N_3341,N_3154,N_3082);
nand U3342 (N_3342,N_3191,N_3142);
and U3343 (N_3343,N_3023,N_3013);
and U3344 (N_3344,N_3056,N_3084);
nand U3345 (N_3345,N_3065,N_3133);
nor U3346 (N_3346,N_3126,N_3112);
nand U3347 (N_3347,N_3138,N_3172);
nand U3348 (N_3348,N_3069,N_3190);
and U3349 (N_3349,N_3164,N_3148);
nand U3350 (N_3350,N_3058,N_3109);
nor U3351 (N_3351,N_3149,N_3068);
nor U3352 (N_3352,N_3194,N_3150);
or U3353 (N_3353,N_3123,N_3189);
nor U3354 (N_3354,N_3070,N_3075);
or U3355 (N_3355,N_3117,N_3105);
nor U3356 (N_3356,N_3162,N_3147);
or U3357 (N_3357,N_3048,N_3114);
nand U3358 (N_3358,N_3048,N_3034);
xnor U3359 (N_3359,N_3099,N_3161);
and U3360 (N_3360,N_3056,N_3006);
nand U3361 (N_3361,N_3197,N_3013);
nor U3362 (N_3362,N_3052,N_3032);
nor U3363 (N_3363,N_3077,N_3169);
nor U3364 (N_3364,N_3146,N_3107);
or U3365 (N_3365,N_3055,N_3109);
and U3366 (N_3366,N_3128,N_3041);
or U3367 (N_3367,N_3015,N_3189);
nand U3368 (N_3368,N_3117,N_3150);
and U3369 (N_3369,N_3127,N_3168);
nor U3370 (N_3370,N_3198,N_3089);
or U3371 (N_3371,N_3119,N_3145);
nor U3372 (N_3372,N_3026,N_3051);
nor U3373 (N_3373,N_3009,N_3138);
nand U3374 (N_3374,N_3190,N_3135);
xor U3375 (N_3375,N_3044,N_3067);
nor U3376 (N_3376,N_3134,N_3157);
or U3377 (N_3377,N_3081,N_3036);
nor U3378 (N_3378,N_3034,N_3049);
nand U3379 (N_3379,N_3066,N_3157);
or U3380 (N_3380,N_3082,N_3053);
and U3381 (N_3381,N_3030,N_3173);
nor U3382 (N_3382,N_3084,N_3151);
or U3383 (N_3383,N_3015,N_3180);
nor U3384 (N_3384,N_3109,N_3038);
and U3385 (N_3385,N_3022,N_3152);
nand U3386 (N_3386,N_3141,N_3177);
and U3387 (N_3387,N_3057,N_3052);
xnor U3388 (N_3388,N_3097,N_3089);
or U3389 (N_3389,N_3109,N_3168);
nand U3390 (N_3390,N_3146,N_3139);
and U3391 (N_3391,N_3071,N_3038);
nor U3392 (N_3392,N_3182,N_3030);
and U3393 (N_3393,N_3062,N_3052);
and U3394 (N_3394,N_3046,N_3062);
and U3395 (N_3395,N_3010,N_3071);
nand U3396 (N_3396,N_3155,N_3130);
or U3397 (N_3397,N_3129,N_3061);
or U3398 (N_3398,N_3004,N_3104);
nor U3399 (N_3399,N_3018,N_3102);
nand U3400 (N_3400,N_3276,N_3352);
nor U3401 (N_3401,N_3220,N_3268);
or U3402 (N_3402,N_3308,N_3343);
xor U3403 (N_3403,N_3226,N_3325);
xnor U3404 (N_3404,N_3238,N_3231);
and U3405 (N_3405,N_3374,N_3318);
or U3406 (N_3406,N_3299,N_3326);
and U3407 (N_3407,N_3236,N_3223);
nand U3408 (N_3408,N_3234,N_3337);
or U3409 (N_3409,N_3336,N_3255);
nor U3410 (N_3410,N_3302,N_3319);
and U3411 (N_3411,N_3244,N_3321);
nand U3412 (N_3412,N_3246,N_3263);
nor U3413 (N_3413,N_3216,N_3388);
nand U3414 (N_3414,N_3367,N_3225);
nor U3415 (N_3415,N_3399,N_3386);
or U3416 (N_3416,N_3202,N_3218);
or U3417 (N_3417,N_3331,N_3311);
and U3418 (N_3418,N_3254,N_3342);
or U3419 (N_3419,N_3382,N_3359);
xnor U3420 (N_3420,N_3240,N_3250);
nand U3421 (N_3421,N_3357,N_3376);
xnor U3422 (N_3422,N_3368,N_3329);
and U3423 (N_3423,N_3341,N_3340);
nand U3424 (N_3424,N_3345,N_3366);
or U3425 (N_3425,N_3380,N_3251);
nand U3426 (N_3426,N_3237,N_3282);
and U3427 (N_3427,N_3292,N_3389);
or U3428 (N_3428,N_3229,N_3230);
nand U3429 (N_3429,N_3204,N_3361);
nor U3430 (N_3430,N_3375,N_3260);
and U3431 (N_3431,N_3287,N_3372);
xnor U3432 (N_3432,N_3256,N_3378);
or U3433 (N_3433,N_3258,N_3264);
nor U3434 (N_3434,N_3232,N_3332);
nor U3435 (N_3435,N_3233,N_3398);
nor U3436 (N_3436,N_3315,N_3205);
nor U3437 (N_3437,N_3291,N_3309);
nor U3438 (N_3438,N_3297,N_3228);
and U3439 (N_3439,N_3206,N_3383);
or U3440 (N_3440,N_3358,N_3209);
and U3441 (N_3441,N_3212,N_3384);
and U3442 (N_3442,N_3377,N_3252);
xor U3443 (N_3443,N_3300,N_3215);
nor U3444 (N_3444,N_3243,N_3353);
nand U3445 (N_3445,N_3270,N_3265);
nor U3446 (N_3446,N_3211,N_3271);
nand U3447 (N_3447,N_3281,N_3219);
and U3448 (N_3448,N_3327,N_3248);
or U3449 (N_3449,N_3347,N_3253);
nand U3450 (N_3450,N_3285,N_3245);
or U3451 (N_3451,N_3391,N_3339);
xor U3452 (N_3452,N_3390,N_3235);
and U3453 (N_3453,N_3279,N_3272);
nor U3454 (N_3454,N_3289,N_3266);
or U3455 (N_3455,N_3294,N_3333);
nand U3456 (N_3456,N_3280,N_3392);
or U3457 (N_3457,N_3262,N_3314);
or U3458 (N_3458,N_3210,N_3394);
nor U3459 (N_3459,N_3356,N_3334);
or U3460 (N_3460,N_3365,N_3381);
and U3461 (N_3461,N_3305,N_3387);
and U3462 (N_3462,N_3295,N_3323);
nand U3463 (N_3463,N_3267,N_3364);
nand U3464 (N_3464,N_3274,N_3301);
nor U3465 (N_3465,N_3203,N_3363);
nor U3466 (N_3466,N_3330,N_3393);
nand U3467 (N_3467,N_3328,N_3249);
nand U3468 (N_3468,N_3369,N_3239);
and U3469 (N_3469,N_3395,N_3261);
xnor U3470 (N_3470,N_3227,N_3348);
nor U3471 (N_3471,N_3354,N_3370);
or U3472 (N_3472,N_3290,N_3257);
or U3473 (N_3473,N_3278,N_3360);
nor U3474 (N_3474,N_3385,N_3217);
nand U3475 (N_3475,N_3277,N_3346);
nor U3476 (N_3476,N_3201,N_3284);
nand U3477 (N_3477,N_3306,N_3371);
xor U3478 (N_3478,N_3335,N_3303);
xnor U3479 (N_3479,N_3313,N_3247);
xor U3480 (N_3480,N_3222,N_3338);
or U3481 (N_3481,N_3379,N_3273);
nor U3482 (N_3482,N_3310,N_3259);
nand U3483 (N_3483,N_3269,N_3349);
and U3484 (N_3484,N_3324,N_3397);
or U3485 (N_3485,N_3317,N_3224);
or U3486 (N_3486,N_3242,N_3208);
or U3487 (N_3487,N_3275,N_3214);
nor U3488 (N_3488,N_3344,N_3312);
and U3489 (N_3489,N_3316,N_3283);
or U3490 (N_3490,N_3207,N_3288);
nor U3491 (N_3491,N_3221,N_3307);
nand U3492 (N_3492,N_3241,N_3355);
and U3493 (N_3493,N_3213,N_3322);
nor U3494 (N_3494,N_3298,N_3304);
or U3495 (N_3495,N_3320,N_3351);
xnor U3496 (N_3496,N_3362,N_3350);
and U3497 (N_3497,N_3296,N_3286);
and U3498 (N_3498,N_3293,N_3396);
nor U3499 (N_3499,N_3200,N_3373);
and U3500 (N_3500,N_3322,N_3299);
and U3501 (N_3501,N_3322,N_3269);
and U3502 (N_3502,N_3378,N_3382);
nand U3503 (N_3503,N_3273,N_3240);
and U3504 (N_3504,N_3391,N_3242);
nand U3505 (N_3505,N_3315,N_3387);
or U3506 (N_3506,N_3250,N_3317);
nor U3507 (N_3507,N_3265,N_3259);
nor U3508 (N_3508,N_3284,N_3245);
nand U3509 (N_3509,N_3381,N_3391);
and U3510 (N_3510,N_3336,N_3387);
xor U3511 (N_3511,N_3208,N_3265);
nor U3512 (N_3512,N_3357,N_3244);
nand U3513 (N_3513,N_3258,N_3313);
nor U3514 (N_3514,N_3335,N_3381);
nand U3515 (N_3515,N_3227,N_3341);
xnor U3516 (N_3516,N_3367,N_3350);
and U3517 (N_3517,N_3259,N_3353);
or U3518 (N_3518,N_3378,N_3331);
or U3519 (N_3519,N_3338,N_3242);
or U3520 (N_3520,N_3297,N_3242);
and U3521 (N_3521,N_3249,N_3365);
and U3522 (N_3522,N_3235,N_3218);
and U3523 (N_3523,N_3367,N_3265);
or U3524 (N_3524,N_3218,N_3312);
or U3525 (N_3525,N_3393,N_3267);
or U3526 (N_3526,N_3247,N_3218);
nand U3527 (N_3527,N_3238,N_3351);
nor U3528 (N_3528,N_3336,N_3298);
and U3529 (N_3529,N_3342,N_3245);
nor U3530 (N_3530,N_3297,N_3304);
or U3531 (N_3531,N_3323,N_3373);
nor U3532 (N_3532,N_3270,N_3295);
nor U3533 (N_3533,N_3358,N_3397);
xnor U3534 (N_3534,N_3390,N_3394);
or U3535 (N_3535,N_3358,N_3382);
nand U3536 (N_3536,N_3284,N_3337);
xor U3537 (N_3537,N_3370,N_3216);
nor U3538 (N_3538,N_3211,N_3391);
or U3539 (N_3539,N_3222,N_3231);
and U3540 (N_3540,N_3204,N_3375);
nor U3541 (N_3541,N_3245,N_3253);
nor U3542 (N_3542,N_3254,N_3296);
or U3543 (N_3543,N_3342,N_3383);
or U3544 (N_3544,N_3358,N_3295);
xnor U3545 (N_3545,N_3231,N_3316);
or U3546 (N_3546,N_3270,N_3245);
nor U3547 (N_3547,N_3207,N_3276);
xnor U3548 (N_3548,N_3271,N_3257);
nor U3549 (N_3549,N_3368,N_3226);
and U3550 (N_3550,N_3300,N_3253);
xnor U3551 (N_3551,N_3307,N_3251);
and U3552 (N_3552,N_3200,N_3287);
and U3553 (N_3553,N_3248,N_3396);
or U3554 (N_3554,N_3295,N_3296);
xor U3555 (N_3555,N_3377,N_3283);
and U3556 (N_3556,N_3204,N_3312);
xor U3557 (N_3557,N_3367,N_3381);
nand U3558 (N_3558,N_3362,N_3388);
nor U3559 (N_3559,N_3360,N_3265);
nand U3560 (N_3560,N_3259,N_3201);
and U3561 (N_3561,N_3283,N_3350);
xor U3562 (N_3562,N_3283,N_3312);
xnor U3563 (N_3563,N_3257,N_3267);
or U3564 (N_3564,N_3348,N_3281);
nor U3565 (N_3565,N_3201,N_3234);
nand U3566 (N_3566,N_3263,N_3315);
and U3567 (N_3567,N_3284,N_3397);
or U3568 (N_3568,N_3223,N_3283);
nor U3569 (N_3569,N_3370,N_3237);
xnor U3570 (N_3570,N_3301,N_3360);
nor U3571 (N_3571,N_3261,N_3241);
nand U3572 (N_3572,N_3364,N_3210);
nand U3573 (N_3573,N_3278,N_3296);
and U3574 (N_3574,N_3393,N_3238);
and U3575 (N_3575,N_3360,N_3226);
nand U3576 (N_3576,N_3318,N_3366);
and U3577 (N_3577,N_3256,N_3279);
xor U3578 (N_3578,N_3294,N_3285);
nor U3579 (N_3579,N_3289,N_3334);
and U3580 (N_3580,N_3373,N_3305);
or U3581 (N_3581,N_3337,N_3332);
nand U3582 (N_3582,N_3273,N_3299);
or U3583 (N_3583,N_3235,N_3377);
or U3584 (N_3584,N_3293,N_3216);
nor U3585 (N_3585,N_3366,N_3375);
nor U3586 (N_3586,N_3318,N_3365);
and U3587 (N_3587,N_3325,N_3242);
xnor U3588 (N_3588,N_3208,N_3271);
or U3589 (N_3589,N_3337,N_3349);
and U3590 (N_3590,N_3261,N_3249);
and U3591 (N_3591,N_3390,N_3346);
nand U3592 (N_3592,N_3246,N_3266);
nor U3593 (N_3593,N_3281,N_3360);
and U3594 (N_3594,N_3373,N_3304);
nor U3595 (N_3595,N_3208,N_3277);
and U3596 (N_3596,N_3263,N_3257);
and U3597 (N_3597,N_3386,N_3303);
or U3598 (N_3598,N_3253,N_3381);
and U3599 (N_3599,N_3380,N_3235);
nand U3600 (N_3600,N_3501,N_3560);
nand U3601 (N_3601,N_3452,N_3514);
nor U3602 (N_3602,N_3496,N_3500);
and U3603 (N_3603,N_3423,N_3440);
or U3604 (N_3604,N_3550,N_3528);
xnor U3605 (N_3605,N_3539,N_3531);
nand U3606 (N_3606,N_3524,N_3599);
nor U3607 (N_3607,N_3545,N_3438);
or U3608 (N_3608,N_3458,N_3510);
nor U3609 (N_3609,N_3597,N_3480);
and U3610 (N_3610,N_3418,N_3554);
and U3611 (N_3611,N_3584,N_3596);
xnor U3612 (N_3612,N_3559,N_3478);
nand U3613 (N_3613,N_3561,N_3569);
or U3614 (N_3614,N_3400,N_3414);
nand U3615 (N_3615,N_3491,N_3562);
or U3616 (N_3616,N_3497,N_3534);
nor U3617 (N_3617,N_3588,N_3567);
xnor U3618 (N_3618,N_3499,N_3434);
or U3619 (N_3619,N_3557,N_3503);
and U3620 (N_3620,N_3530,N_3426);
nand U3621 (N_3621,N_3512,N_3495);
and U3622 (N_3622,N_3592,N_3445);
and U3623 (N_3623,N_3527,N_3536);
and U3624 (N_3624,N_3424,N_3506);
nand U3625 (N_3625,N_3430,N_3579);
nand U3626 (N_3626,N_3403,N_3543);
nor U3627 (N_3627,N_3407,N_3436);
and U3628 (N_3628,N_3410,N_3476);
or U3629 (N_3629,N_3577,N_3455);
nand U3630 (N_3630,N_3448,N_3515);
nand U3631 (N_3631,N_3553,N_3401);
nand U3632 (N_3632,N_3583,N_3493);
or U3633 (N_3633,N_3537,N_3513);
nand U3634 (N_3634,N_3429,N_3412);
and U3635 (N_3635,N_3463,N_3516);
nor U3636 (N_3636,N_3484,N_3415);
xnor U3637 (N_3637,N_3489,N_3581);
nand U3638 (N_3638,N_3441,N_3535);
xor U3639 (N_3639,N_3416,N_3533);
and U3640 (N_3640,N_3428,N_3435);
nor U3641 (N_3641,N_3548,N_3544);
nand U3642 (N_3642,N_3425,N_3482);
nand U3643 (N_3643,N_3477,N_3467);
or U3644 (N_3644,N_3479,N_3454);
and U3645 (N_3645,N_3413,N_3520);
or U3646 (N_3646,N_3421,N_3558);
nor U3647 (N_3647,N_3572,N_3508);
nor U3648 (N_3648,N_3521,N_3585);
nor U3649 (N_3649,N_3565,N_3573);
xnor U3650 (N_3650,N_3465,N_3555);
nor U3651 (N_3651,N_3541,N_3402);
or U3652 (N_3652,N_3546,N_3447);
xor U3653 (N_3653,N_3486,N_3459);
nand U3654 (N_3654,N_3576,N_3466);
or U3655 (N_3655,N_3422,N_3474);
nand U3656 (N_3656,N_3504,N_3431);
xor U3657 (N_3657,N_3411,N_3589);
and U3658 (N_3658,N_3551,N_3575);
or U3659 (N_3659,N_3487,N_3442);
xnor U3660 (N_3660,N_3409,N_3517);
and U3661 (N_3661,N_3502,N_3494);
xnor U3662 (N_3662,N_3450,N_3519);
or U3663 (N_3663,N_3590,N_3507);
or U3664 (N_3664,N_3488,N_3439);
or U3665 (N_3665,N_3571,N_3468);
and U3666 (N_3666,N_3570,N_3598);
and U3667 (N_3667,N_3523,N_3563);
nand U3668 (N_3668,N_3462,N_3580);
and U3669 (N_3669,N_3549,N_3595);
nand U3670 (N_3670,N_3451,N_3540);
or U3671 (N_3671,N_3470,N_3505);
nor U3672 (N_3672,N_3475,N_3481);
nand U3673 (N_3673,N_3511,N_3464);
xor U3674 (N_3674,N_3587,N_3568);
nor U3675 (N_3675,N_3483,N_3556);
nor U3676 (N_3676,N_3469,N_3538);
nand U3677 (N_3677,N_3498,N_3574);
nand U3678 (N_3678,N_3453,N_3582);
and U3679 (N_3679,N_3564,N_3525);
and U3680 (N_3680,N_3408,N_3485);
xor U3681 (N_3681,N_3419,N_3594);
nor U3682 (N_3682,N_3444,N_3417);
nor U3683 (N_3683,N_3472,N_3446);
nor U3684 (N_3684,N_3593,N_3492);
xor U3685 (N_3685,N_3433,N_3552);
and U3686 (N_3686,N_3443,N_3404);
or U3687 (N_3687,N_3456,N_3586);
nor U3688 (N_3688,N_3566,N_3471);
xnor U3689 (N_3689,N_3526,N_3532);
or U3690 (N_3690,N_3542,N_3522);
nor U3691 (N_3691,N_3473,N_3405);
or U3692 (N_3692,N_3406,N_3490);
nor U3693 (N_3693,N_3437,N_3457);
nor U3694 (N_3694,N_3432,N_3509);
or U3695 (N_3695,N_3427,N_3461);
nor U3696 (N_3696,N_3460,N_3518);
nor U3697 (N_3697,N_3529,N_3547);
xor U3698 (N_3698,N_3578,N_3591);
nand U3699 (N_3699,N_3449,N_3420);
nand U3700 (N_3700,N_3490,N_3493);
or U3701 (N_3701,N_3588,N_3571);
nor U3702 (N_3702,N_3446,N_3432);
or U3703 (N_3703,N_3445,N_3451);
nand U3704 (N_3704,N_3413,N_3458);
or U3705 (N_3705,N_3555,N_3529);
or U3706 (N_3706,N_3487,N_3587);
and U3707 (N_3707,N_3456,N_3544);
nor U3708 (N_3708,N_3491,N_3456);
nor U3709 (N_3709,N_3488,N_3454);
or U3710 (N_3710,N_3563,N_3412);
nand U3711 (N_3711,N_3406,N_3563);
and U3712 (N_3712,N_3588,N_3515);
nor U3713 (N_3713,N_3439,N_3466);
nor U3714 (N_3714,N_3498,N_3533);
nand U3715 (N_3715,N_3478,N_3505);
nand U3716 (N_3716,N_3540,N_3526);
or U3717 (N_3717,N_3433,N_3435);
nand U3718 (N_3718,N_3436,N_3475);
or U3719 (N_3719,N_3551,N_3590);
and U3720 (N_3720,N_3490,N_3538);
and U3721 (N_3721,N_3475,N_3522);
nor U3722 (N_3722,N_3447,N_3540);
and U3723 (N_3723,N_3581,N_3547);
or U3724 (N_3724,N_3453,N_3412);
nand U3725 (N_3725,N_3533,N_3521);
and U3726 (N_3726,N_3558,N_3466);
nor U3727 (N_3727,N_3549,N_3568);
nor U3728 (N_3728,N_3428,N_3530);
nor U3729 (N_3729,N_3419,N_3488);
nand U3730 (N_3730,N_3521,N_3477);
nor U3731 (N_3731,N_3468,N_3406);
nor U3732 (N_3732,N_3502,N_3454);
and U3733 (N_3733,N_3480,N_3554);
xnor U3734 (N_3734,N_3574,N_3561);
and U3735 (N_3735,N_3445,N_3519);
or U3736 (N_3736,N_3557,N_3440);
nand U3737 (N_3737,N_3443,N_3493);
or U3738 (N_3738,N_3556,N_3548);
xor U3739 (N_3739,N_3566,N_3567);
nand U3740 (N_3740,N_3435,N_3578);
or U3741 (N_3741,N_3440,N_3593);
nand U3742 (N_3742,N_3400,N_3443);
nand U3743 (N_3743,N_3523,N_3446);
or U3744 (N_3744,N_3575,N_3507);
and U3745 (N_3745,N_3594,N_3456);
or U3746 (N_3746,N_3464,N_3528);
nand U3747 (N_3747,N_3489,N_3550);
nand U3748 (N_3748,N_3422,N_3465);
nor U3749 (N_3749,N_3566,N_3515);
nor U3750 (N_3750,N_3470,N_3484);
nor U3751 (N_3751,N_3480,N_3506);
nand U3752 (N_3752,N_3551,N_3410);
xor U3753 (N_3753,N_3533,N_3497);
nand U3754 (N_3754,N_3549,N_3452);
nor U3755 (N_3755,N_3408,N_3554);
nand U3756 (N_3756,N_3423,N_3448);
nor U3757 (N_3757,N_3588,N_3439);
nor U3758 (N_3758,N_3408,N_3409);
nand U3759 (N_3759,N_3480,N_3451);
nor U3760 (N_3760,N_3578,N_3469);
nand U3761 (N_3761,N_3430,N_3554);
and U3762 (N_3762,N_3455,N_3431);
xor U3763 (N_3763,N_3561,N_3461);
or U3764 (N_3764,N_3596,N_3576);
and U3765 (N_3765,N_3484,N_3586);
and U3766 (N_3766,N_3524,N_3474);
or U3767 (N_3767,N_3418,N_3473);
or U3768 (N_3768,N_3449,N_3476);
nor U3769 (N_3769,N_3484,N_3536);
nor U3770 (N_3770,N_3557,N_3530);
nor U3771 (N_3771,N_3487,N_3556);
xnor U3772 (N_3772,N_3476,N_3599);
and U3773 (N_3773,N_3550,N_3543);
nand U3774 (N_3774,N_3435,N_3415);
and U3775 (N_3775,N_3461,N_3543);
and U3776 (N_3776,N_3588,N_3473);
nand U3777 (N_3777,N_3530,N_3412);
nand U3778 (N_3778,N_3533,N_3437);
or U3779 (N_3779,N_3591,N_3513);
xor U3780 (N_3780,N_3457,N_3413);
and U3781 (N_3781,N_3512,N_3544);
and U3782 (N_3782,N_3423,N_3583);
nand U3783 (N_3783,N_3562,N_3520);
nand U3784 (N_3784,N_3587,N_3405);
nor U3785 (N_3785,N_3499,N_3489);
nor U3786 (N_3786,N_3434,N_3451);
or U3787 (N_3787,N_3591,N_3401);
or U3788 (N_3788,N_3515,N_3461);
and U3789 (N_3789,N_3460,N_3430);
or U3790 (N_3790,N_3408,N_3439);
nor U3791 (N_3791,N_3433,N_3476);
and U3792 (N_3792,N_3431,N_3465);
nand U3793 (N_3793,N_3501,N_3555);
xnor U3794 (N_3794,N_3522,N_3548);
nor U3795 (N_3795,N_3567,N_3427);
and U3796 (N_3796,N_3568,N_3525);
nand U3797 (N_3797,N_3458,N_3557);
nor U3798 (N_3798,N_3434,N_3559);
nand U3799 (N_3799,N_3474,N_3461);
and U3800 (N_3800,N_3620,N_3632);
and U3801 (N_3801,N_3722,N_3721);
or U3802 (N_3802,N_3602,N_3629);
and U3803 (N_3803,N_3683,N_3713);
or U3804 (N_3804,N_3709,N_3610);
xnor U3805 (N_3805,N_3616,N_3724);
or U3806 (N_3806,N_3799,N_3678);
nand U3807 (N_3807,N_3670,N_3730);
or U3808 (N_3808,N_3635,N_3698);
and U3809 (N_3809,N_3703,N_3797);
nand U3810 (N_3810,N_3707,N_3735);
nor U3811 (N_3811,N_3691,N_3753);
nand U3812 (N_3812,N_3764,N_3762);
and U3813 (N_3813,N_3796,N_3771);
and U3814 (N_3814,N_3720,N_3666);
or U3815 (N_3815,N_3712,N_3785);
or U3816 (N_3816,N_3630,N_3768);
or U3817 (N_3817,N_3687,N_3706);
or U3818 (N_3818,N_3729,N_3790);
and U3819 (N_3819,N_3695,N_3614);
nand U3820 (N_3820,N_3773,N_3739);
xnor U3821 (N_3821,N_3612,N_3637);
nor U3822 (N_3822,N_3663,N_3767);
nor U3823 (N_3823,N_3743,N_3606);
nor U3824 (N_3824,N_3631,N_3717);
and U3825 (N_3825,N_3676,N_3646);
or U3826 (N_3826,N_3634,N_3798);
nor U3827 (N_3827,N_3696,N_3608);
nor U3828 (N_3828,N_3781,N_3626);
nand U3829 (N_3829,N_3752,N_3662);
nor U3830 (N_3830,N_3622,N_3701);
nand U3831 (N_3831,N_3652,N_3638);
and U3832 (N_3832,N_3688,N_3628);
nand U3833 (N_3833,N_3784,N_3783);
xnor U3834 (N_3834,N_3750,N_3601);
nand U3835 (N_3835,N_3760,N_3731);
nand U3836 (N_3836,N_3761,N_3742);
nand U3837 (N_3837,N_3748,N_3705);
nand U3838 (N_3838,N_3774,N_3672);
nor U3839 (N_3839,N_3759,N_3625);
or U3840 (N_3840,N_3741,N_3776);
nand U3841 (N_3841,N_3780,N_3793);
and U3842 (N_3842,N_3736,N_3653);
nand U3843 (N_3843,N_3747,N_3642);
or U3844 (N_3844,N_3636,N_3765);
nor U3845 (N_3845,N_3746,N_3795);
nor U3846 (N_3846,N_3681,N_3770);
nor U3847 (N_3847,N_3618,N_3684);
and U3848 (N_3848,N_3650,N_3699);
or U3849 (N_3849,N_3639,N_3613);
or U3850 (N_3850,N_3654,N_3737);
nor U3851 (N_3851,N_3690,N_3692);
nor U3852 (N_3852,N_3782,N_3775);
nand U3853 (N_3853,N_3671,N_3623);
nor U3854 (N_3854,N_3603,N_3751);
and U3855 (N_3855,N_3607,N_3674);
nor U3856 (N_3856,N_3749,N_3621);
nor U3857 (N_3857,N_3660,N_3697);
and U3858 (N_3858,N_3725,N_3609);
and U3859 (N_3859,N_3604,N_3728);
nor U3860 (N_3860,N_3791,N_3641);
nor U3861 (N_3861,N_3656,N_3754);
nand U3862 (N_3862,N_3716,N_3617);
nor U3863 (N_3863,N_3633,N_3605);
nor U3864 (N_3864,N_3682,N_3792);
or U3865 (N_3865,N_3675,N_3704);
or U3866 (N_3866,N_3667,N_3711);
nor U3867 (N_3867,N_3645,N_3644);
and U3868 (N_3868,N_3755,N_3665);
xor U3869 (N_3869,N_3772,N_3763);
nor U3870 (N_3870,N_3734,N_3611);
nor U3871 (N_3871,N_3640,N_3723);
nor U3872 (N_3872,N_3740,N_3651);
nor U3873 (N_3873,N_3715,N_3700);
nand U3874 (N_3874,N_3655,N_3680);
nand U3875 (N_3875,N_3669,N_3788);
nor U3876 (N_3876,N_3756,N_3710);
nand U3877 (N_3877,N_3619,N_3794);
or U3878 (N_3878,N_3769,N_3789);
nand U3879 (N_3879,N_3673,N_3757);
xnor U3880 (N_3880,N_3738,N_3693);
xor U3881 (N_3881,N_3664,N_3732);
nand U3882 (N_3882,N_3657,N_3659);
nor U3883 (N_3883,N_3727,N_3702);
and U3884 (N_3884,N_3714,N_3745);
nor U3885 (N_3885,N_3719,N_3766);
nand U3886 (N_3886,N_3694,N_3758);
and U3887 (N_3887,N_3679,N_3726);
or U3888 (N_3888,N_3744,N_3643);
nand U3889 (N_3889,N_3786,N_3778);
nor U3890 (N_3890,N_3647,N_3648);
nor U3891 (N_3891,N_3600,N_3718);
and U3892 (N_3892,N_3686,N_3689);
nor U3893 (N_3893,N_3615,N_3661);
nand U3894 (N_3894,N_3787,N_3777);
nor U3895 (N_3895,N_3649,N_3779);
nand U3896 (N_3896,N_3733,N_3708);
nor U3897 (N_3897,N_3658,N_3627);
and U3898 (N_3898,N_3685,N_3677);
nor U3899 (N_3899,N_3668,N_3624);
and U3900 (N_3900,N_3624,N_3738);
or U3901 (N_3901,N_3629,N_3760);
and U3902 (N_3902,N_3783,N_3750);
nor U3903 (N_3903,N_3736,N_3665);
nand U3904 (N_3904,N_3764,N_3652);
nor U3905 (N_3905,N_3685,N_3704);
and U3906 (N_3906,N_3713,N_3740);
or U3907 (N_3907,N_3640,N_3792);
or U3908 (N_3908,N_3621,N_3626);
nand U3909 (N_3909,N_3698,N_3606);
or U3910 (N_3910,N_3774,N_3652);
nand U3911 (N_3911,N_3704,N_3650);
or U3912 (N_3912,N_3779,N_3692);
or U3913 (N_3913,N_3675,N_3650);
or U3914 (N_3914,N_3693,N_3755);
xor U3915 (N_3915,N_3777,N_3757);
and U3916 (N_3916,N_3750,N_3660);
nand U3917 (N_3917,N_3643,N_3787);
or U3918 (N_3918,N_3612,N_3777);
nand U3919 (N_3919,N_3617,N_3623);
xnor U3920 (N_3920,N_3652,N_3673);
xor U3921 (N_3921,N_3620,N_3781);
or U3922 (N_3922,N_3675,N_3620);
nor U3923 (N_3923,N_3758,N_3794);
nor U3924 (N_3924,N_3626,N_3686);
nand U3925 (N_3925,N_3690,N_3733);
or U3926 (N_3926,N_3634,N_3621);
nor U3927 (N_3927,N_3606,N_3715);
nor U3928 (N_3928,N_3637,N_3692);
nand U3929 (N_3929,N_3786,N_3781);
nor U3930 (N_3930,N_3615,N_3679);
xor U3931 (N_3931,N_3616,N_3652);
or U3932 (N_3932,N_3761,N_3753);
or U3933 (N_3933,N_3732,N_3740);
and U3934 (N_3934,N_3610,N_3691);
and U3935 (N_3935,N_3670,N_3766);
or U3936 (N_3936,N_3706,N_3695);
nor U3937 (N_3937,N_3654,N_3784);
nor U3938 (N_3938,N_3770,N_3707);
or U3939 (N_3939,N_3792,N_3650);
and U3940 (N_3940,N_3765,N_3656);
and U3941 (N_3941,N_3633,N_3692);
nand U3942 (N_3942,N_3610,N_3761);
and U3943 (N_3943,N_3724,N_3683);
or U3944 (N_3944,N_3683,N_3617);
or U3945 (N_3945,N_3779,N_3699);
xnor U3946 (N_3946,N_3613,N_3754);
nand U3947 (N_3947,N_3765,N_3727);
or U3948 (N_3948,N_3611,N_3601);
and U3949 (N_3949,N_3631,N_3642);
nand U3950 (N_3950,N_3746,N_3771);
or U3951 (N_3951,N_3661,N_3646);
or U3952 (N_3952,N_3678,N_3613);
nor U3953 (N_3953,N_3753,N_3732);
nand U3954 (N_3954,N_3690,N_3728);
nand U3955 (N_3955,N_3754,N_3715);
xnor U3956 (N_3956,N_3685,N_3752);
nor U3957 (N_3957,N_3779,N_3654);
nor U3958 (N_3958,N_3779,N_3682);
or U3959 (N_3959,N_3799,N_3784);
nor U3960 (N_3960,N_3701,N_3660);
nor U3961 (N_3961,N_3655,N_3747);
and U3962 (N_3962,N_3784,N_3747);
nand U3963 (N_3963,N_3691,N_3646);
nor U3964 (N_3964,N_3728,N_3738);
nor U3965 (N_3965,N_3669,N_3680);
or U3966 (N_3966,N_3704,N_3601);
nand U3967 (N_3967,N_3794,N_3674);
and U3968 (N_3968,N_3645,N_3655);
nand U3969 (N_3969,N_3782,N_3681);
and U3970 (N_3970,N_3639,N_3793);
or U3971 (N_3971,N_3670,N_3754);
and U3972 (N_3972,N_3770,N_3640);
and U3973 (N_3973,N_3787,N_3666);
nand U3974 (N_3974,N_3734,N_3604);
and U3975 (N_3975,N_3691,N_3763);
and U3976 (N_3976,N_3602,N_3744);
nand U3977 (N_3977,N_3776,N_3723);
xor U3978 (N_3978,N_3704,N_3677);
or U3979 (N_3979,N_3771,N_3763);
nor U3980 (N_3980,N_3723,N_3609);
nor U3981 (N_3981,N_3709,N_3658);
xnor U3982 (N_3982,N_3795,N_3619);
and U3983 (N_3983,N_3697,N_3606);
or U3984 (N_3984,N_3778,N_3725);
nor U3985 (N_3985,N_3628,N_3686);
xor U3986 (N_3986,N_3634,N_3732);
or U3987 (N_3987,N_3712,N_3656);
nand U3988 (N_3988,N_3677,N_3748);
and U3989 (N_3989,N_3644,N_3660);
nand U3990 (N_3990,N_3650,N_3765);
nor U3991 (N_3991,N_3625,N_3738);
nor U3992 (N_3992,N_3765,N_3678);
nor U3993 (N_3993,N_3677,N_3778);
nor U3994 (N_3994,N_3727,N_3782);
xnor U3995 (N_3995,N_3726,N_3664);
nand U3996 (N_3996,N_3663,N_3655);
nand U3997 (N_3997,N_3625,N_3652);
nand U3998 (N_3998,N_3790,N_3781);
or U3999 (N_3999,N_3676,N_3714);
and U4000 (N_4000,N_3872,N_3887);
or U4001 (N_4001,N_3981,N_3905);
or U4002 (N_4002,N_3923,N_3853);
and U4003 (N_4003,N_3941,N_3976);
or U4004 (N_4004,N_3915,N_3866);
or U4005 (N_4005,N_3818,N_3878);
or U4006 (N_4006,N_3901,N_3879);
xor U4007 (N_4007,N_3978,N_3885);
nor U4008 (N_4008,N_3954,N_3994);
or U4009 (N_4009,N_3820,N_3826);
nand U4010 (N_4010,N_3964,N_3987);
and U4011 (N_4011,N_3971,N_3873);
or U4012 (N_4012,N_3880,N_3902);
or U4013 (N_4013,N_3936,N_3877);
nand U4014 (N_4014,N_3908,N_3824);
or U4015 (N_4015,N_3990,N_3926);
or U4016 (N_4016,N_3995,N_3910);
xnor U4017 (N_4017,N_3808,N_3802);
or U4018 (N_4018,N_3865,N_3825);
and U4019 (N_4019,N_3958,N_3858);
nor U4020 (N_4020,N_3860,N_3803);
nand U4021 (N_4021,N_3851,N_3983);
nor U4022 (N_4022,N_3848,N_3919);
nand U4023 (N_4023,N_3817,N_3822);
nand U4024 (N_4024,N_3998,N_3918);
nand U4025 (N_4025,N_3973,N_3811);
or U4026 (N_4026,N_3881,N_3831);
or U4027 (N_4027,N_3934,N_3969);
nor U4028 (N_4028,N_3986,N_3884);
xnor U4029 (N_4029,N_3943,N_3830);
or U4030 (N_4030,N_3862,N_3835);
or U4031 (N_4031,N_3871,N_3847);
nand U4032 (N_4032,N_3948,N_3875);
and U4033 (N_4033,N_3869,N_3975);
xnor U4034 (N_4034,N_3963,N_3819);
nor U4035 (N_4035,N_3967,N_3816);
and U4036 (N_4036,N_3886,N_3834);
nand U4037 (N_4037,N_3906,N_3841);
nor U4038 (N_4038,N_3989,N_3916);
nand U4039 (N_4039,N_3924,N_3947);
nand U4040 (N_4040,N_3845,N_3843);
and U4041 (N_4041,N_3974,N_3951);
xnor U4042 (N_4042,N_3933,N_3913);
nand U4043 (N_4043,N_3961,N_3813);
or U4044 (N_4044,N_3985,N_3827);
or U4045 (N_4045,N_3839,N_3999);
or U4046 (N_4046,N_3970,N_3997);
and U4047 (N_4047,N_3828,N_3868);
nand U4048 (N_4048,N_3836,N_3863);
and U4049 (N_4049,N_3829,N_3917);
and U4050 (N_4050,N_3892,N_3896);
and U4051 (N_4051,N_3833,N_3844);
nand U4052 (N_4052,N_3800,N_3946);
nor U4053 (N_4053,N_3903,N_3883);
nor U4054 (N_4054,N_3939,N_3991);
nor U4055 (N_4055,N_3935,N_3938);
xor U4056 (N_4056,N_3805,N_3952);
nand U4057 (N_4057,N_3979,N_3955);
and U4058 (N_4058,N_3942,N_3864);
nand U4059 (N_4059,N_3912,N_3837);
or U4060 (N_4060,N_3909,N_3992);
nand U4061 (N_4061,N_3932,N_3899);
nand U4062 (N_4062,N_3804,N_3890);
or U4063 (N_4063,N_3874,N_3925);
and U4064 (N_4064,N_3855,N_3815);
or U4065 (N_4065,N_3928,N_3982);
and U4066 (N_4066,N_3950,N_3888);
and U4067 (N_4067,N_3870,N_3895);
nor U4068 (N_4068,N_3840,N_3857);
xnor U4069 (N_4069,N_3859,N_3809);
xnor U4070 (N_4070,N_3968,N_3957);
and U4071 (N_4071,N_3977,N_3920);
xnor U4072 (N_4072,N_3842,N_3944);
nor U4073 (N_4073,N_3984,N_3993);
xnor U4074 (N_4074,N_3852,N_3861);
nand U4075 (N_4075,N_3931,N_3980);
nor U4076 (N_4076,N_3965,N_3945);
and U4077 (N_4077,N_3907,N_3900);
and U4078 (N_4078,N_3807,N_3856);
nor U4079 (N_4079,N_3810,N_3893);
or U4080 (N_4080,N_3882,N_3854);
nand U4081 (N_4081,N_3949,N_3801);
or U4082 (N_4082,N_3867,N_3914);
xnor U4083 (N_4083,N_3904,N_3806);
or U4084 (N_4084,N_3849,N_3897);
nand U4085 (N_4085,N_3927,N_3930);
or U4086 (N_4086,N_3814,N_3988);
nand U4087 (N_4087,N_3960,N_3921);
xor U4088 (N_4088,N_3876,N_3953);
or U4089 (N_4089,N_3821,N_3846);
nand U4090 (N_4090,N_3972,N_3823);
nor U4091 (N_4091,N_3937,N_3911);
or U4092 (N_4092,N_3838,N_3959);
or U4093 (N_4093,N_3962,N_3894);
or U4094 (N_4094,N_3812,N_3966);
xnor U4095 (N_4095,N_3850,N_3891);
nand U4096 (N_4096,N_3889,N_3996);
xnor U4097 (N_4097,N_3832,N_3922);
nand U4098 (N_4098,N_3940,N_3956);
xor U4099 (N_4099,N_3898,N_3929);
nand U4100 (N_4100,N_3887,N_3936);
nor U4101 (N_4101,N_3893,N_3975);
or U4102 (N_4102,N_3916,N_3819);
nand U4103 (N_4103,N_3852,N_3850);
nor U4104 (N_4104,N_3999,N_3851);
nor U4105 (N_4105,N_3824,N_3917);
or U4106 (N_4106,N_3833,N_3880);
nor U4107 (N_4107,N_3809,N_3893);
xnor U4108 (N_4108,N_3959,N_3953);
or U4109 (N_4109,N_3988,N_3940);
nand U4110 (N_4110,N_3976,N_3892);
nand U4111 (N_4111,N_3976,N_3820);
and U4112 (N_4112,N_3978,N_3950);
nor U4113 (N_4113,N_3973,N_3936);
or U4114 (N_4114,N_3988,N_3949);
or U4115 (N_4115,N_3972,N_3915);
xor U4116 (N_4116,N_3918,N_3908);
or U4117 (N_4117,N_3851,N_3923);
and U4118 (N_4118,N_3831,N_3970);
nand U4119 (N_4119,N_3868,N_3968);
or U4120 (N_4120,N_3998,N_3955);
nand U4121 (N_4121,N_3892,N_3855);
and U4122 (N_4122,N_3845,N_3884);
nor U4123 (N_4123,N_3825,N_3852);
nand U4124 (N_4124,N_3897,N_3978);
xor U4125 (N_4125,N_3915,N_3894);
or U4126 (N_4126,N_3925,N_3885);
and U4127 (N_4127,N_3855,N_3809);
nand U4128 (N_4128,N_3931,N_3807);
or U4129 (N_4129,N_3829,N_3888);
or U4130 (N_4130,N_3857,N_3831);
and U4131 (N_4131,N_3806,N_3830);
or U4132 (N_4132,N_3957,N_3901);
nor U4133 (N_4133,N_3885,N_3979);
nand U4134 (N_4134,N_3973,N_3827);
nor U4135 (N_4135,N_3825,N_3898);
nor U4136 (N_4136,N_3848,N_3856);
and U4137 (N_4137,N_3925,N_3805);
nand U4138 (N_4138,N_3833,N_3871);
nand U4139 (N_4139,N_3951,N_3932);
nand U4140 (N_4140,N_3959,N_3801);
nor U4141 (N_4141,N_3869,N_3987);
nand U4142 (N_4142,N_3888,N_3902);
or U4143 (N_4143,N_3868,N_3928);
nand U4144 (N_4144,N_3934,N_3968);
nor U4145 (N_4145,N_3886,N_3977);
or U4146 (N_4146,N_3998,N_3950);
nand U4147 (N_4147,N_3991,N_3863);
or U4148 (N_4148,N_3894,N_3911);
xor U4149 (N_4149,N_3972,N_3981);
nor U4150 (N_4150,N_3846,N_3926);
or U4151 (N_4151,N_3881,N_3991);
or U4152 (N_4152,N_3882,N_3972);
and U4153 (N_4153,N_3816,N_3997);
nand U4154 (N_4154,N_3840,N_3994);
nand U4155 (N_4155,N_3929,N_3955);
or U4156 (N_4156,N_3805,N_3908);
xnor U4157 (N_4157,N_3985,N_3823);
or U4158 (N_4158,N_3815,N_3832);
and U4159 (N_4159,N_3864,N_3899);
and U4160 (N_4160,N_3847,N_3825);
nor U4161 (N_4161,N_3864,N_3841);
nand U4162 (N_4162,N_3899,N_3838);
and U4163 (N_4163,N_3863,N_3984);
nand U4164 (N_4164,N_3990,N_3867);
nand U4165 (N_4165,N_3864,N_3928);
or U4166 (N_4166,N_3963,N_3885);
nand U4167 (N_4167,N_3868,N_3884);
nand U4168 (N_4168,N_3897,N_3985);
nor U4169 (N_4169,N_3859,N_3861);
or U4170 (N_4170,N_3901,N_3841);
and U4171 (N_4171,N_3999,N_3874);
or U4172 (N_4172,N_3851,N_3809);
or U4173 (N_4173,N_3953,N_3951);
or U4174 (N_4174,N_3871,N_3928);
nand U4175 (N_4175,N_3821,N_3975);
xnor U4176 (N_4176,N_3869,N_3983);
or U4177 (N_4177,N_3897,N_3934);
or U4178 (N_4178,N_3841,N_3824);
or U4179 (N_4179,N_3870,N_3953);
and U4180 (N_4180,N_3932,N_3937);
nor U4181 (N_4181,N_3809,N_3962);
or U4182 (N_4182,N_3903,N_3999);
or U4183 (N_4183,N_3887,N_3923);
nand U4184 (N_4184,N_3936,N_3830);
nand U4185 (N_4185,N_3999,N_3988);
nor U4186 (N_4186,N_3807,N_3949);
nor U4187 (N_4187,N_3956,N_3866);
or U4188 (N_4188,N_3964,N_3914);
or U4189 (N_4189,N_3945,N_3817);
and U4190 (N_4190,N_3983,N_3921);
or U4191 (N_4191,N_3938,N_3851);
or U4192 (N_4192,N_3882,N_3804);
or U4193 (N_4193,N_3918,N_3836);
or U4194 (N_4194,N_3882,N_3927);
nand U4195 (N_4195,N_3974,N_3897);
nand U4196 (N_4196,N_3802,N_3908);
or U4197 (N_4197,N_3905,N_3886);
xor U4198 (N_4198,N_3847,N_3968);
and U4199 (N_4199,N_3846,N_3844);
and U4200 (N_4200,N_4153,N_4038);
or U4201 (N_4201,N_4198,N_4003);
xor U4202 (N_4202,N_4194,N_4135);
nand U4203 (N_4203,N_4181,N_4188);
or U4204 (N_4204,N_4175,N_4160);
nand U4205 (N_4205,N_4088,N_4069);
nor U4206 (N_4206,N_4056,N_4016);
nor U4207 (N_4207,N_4070,N_4063);
and U4208 (N_4208,N_4112,N_4171);
or U4209 (N_4209,N_4074,N_4140);
or U4210 (N_4210,N_4180,N_4080);
or U4211 (N_4211,N_4119,N_4129);
or U4212 (N_4212,N_4136,N_4048);
or U4213 (N_4213,N_4001,N_4137);
or U4214 (N_4214,N_4092,N_4067);
and U4215 (N_4215,N_4057,N_4085);
nor U4216 (N_4216,N_4115,N_4009);
xor U4217 (N_4217,N_4053,N_4169);
nor U4218 (N_4218,N_4018,N_4103);
nor U4219 (N_4219,N_4022,N_4060);
xnor U4220 (N_4220,N_4150,N_4086);
and U4221 (N_4221,N_4064,N_4146);
nor U4222 (N_4222,N_4131,N_4004);
and U4223 (N_4223,N_4174,N_4000);
xor U4224 (N_4224,N_4095,N_4141);
xnor U4225 (N_4225,N_4111,N_4072);
and U4226 (N_4226,N_4079,N_4168);
or U4227 (N_4227,N_4091,N_4030);
and U4228 (N_4228,N_4139,N_4149);
and U4229 (N_4229,N_4005,N_4076);
nand U4230 (N_4230,N_4190,N_4010);
xor U4231 (N_4231,N_4024,N_4020);
nor U4232 (N_4232,N_4002,N_4100);
or U4233 (N_4233,N_4037,N_4156);
and U4234 (N_4234,N_4148,N_4101);
or U4235 (N_4235,N_4179,N_4107);
and U4236 (N_4236,N_4033,N_4071);
or U4237 (N_4237,N_4138,N_4089);
nand U4238 (N_4238,N_4128,N_4196);
nand U4239 (N_4239,N_4161,N_4118);
and U4240 (N_4240,N_4051,N_4078);
or U4241 (N_4241,N_4054,N_4124);
or U4242 (N_4242,N_4110,N_4102);
nand U4243 (N_4243,N_4015,N_4090);
nor U4244 (N_4244,N_4039,N_4096);
nand U4245 (N_4245,N_4127,N_4026);
and U4246 (N_4246,N_4025,N_4104);
nand U4247 (N_4247,N_4049,N_4028);
or U4248 (N_4248,N_4029,N_4176);
and U4249 (N_4249,N_4084,N_4155);
nor U4250 (N_4250,N_4183,N_4162);
nand U4251 (N_4251,N_4130,N_4159);
and U4252 (N_4252,N_4152,N_4185);
and U4253 (N_4253,N_4012,N_4065);
and U4254 (N_4254,N_4113,N_4094);
xor U4255 (N_4255,N_4031,N_4133);
nand U4256 (N_4256,N_4173,N_4027);
nand U4257 (N_4257,N_4062,N_4117);
nor U4258 (N_4258,N_4134,N_4041);
nor U4259 (N_4259,N_4109,N_4077);
and U4260 (N_4260,N_4036,N_4093);
and U4261 (N_4261,N_4158,N_4034);
nor U4262 (N_4262,N_4166,N_4098);
or U4263 (N_4263,N_4035,N_4178);
and U4264 (N_4264,N_4019,N_4099);
and U4265 (N_4265,N_4132,N_4055);
nand U4266 (N_4266,N_4042,N_4187);
or U4267 (N_4267,N_4114,N_4043);
nor U4268 (N_4268,N_4106,N_4145);
or U4269 (N_4269,N_4105,N_4083);
nor U4270 (N_4270,N_4052,N_4047);
nor U4271 (N_4271,N_4108,N_4165);
nor U4272 (N_4272,N_4182,N_4046);
nor U4273 (N_4273,N_4157,N_4144);
xor U4274 (N_4274,N_4032,N_4170);
and U4275 (N_4275,N_4040,N_4058);
nor U4276 (N_4276,N_4142,N_4021);
nand U4277 (N_4277,N_4151,N_4050);
nor U4278 (N_4278,N_4081,N_4044);
nand U4279 (N_4279,N_4121,N_4184);
and U4280 (N_4280,N_4097,N_4172);
xor U4281 (N_4281,N_4116,N_4006);
or U4282 (N_4282,N_4191,N_4143);
nor U4283 (N_4283,N_4073,N_4122);
or U4284 (N_4284,N_4186,N_4199);
nor U4285 (N_4285,N_4177,N_4167);
or U4286 (N_4286,N_4075,N_4087);
nand U4287 (N_4287,N_4147,N_4013);
and U4288 (N_4288,N_4014,N_4007);
and U4289 (N_4289,N_4008,N_4068);
or U4290 (N_4290,N_4082,N_4017);
and U4291 (N_4291,N_4163,N_4061);
nand U4292 (N_4292,N_4197,N_4154);
and U4293 (N_4293,N_4045,N_4125);
and U4294 (N_4294,N_4195,N_4123);
nor U4295 (N_4295,N_4059,N_4189);
and U4296 (N_4296,N_4164,N_4023);
nor U4297 (N_4297,N_4126,N_4011);
nand U4298 (N_4298,N_4066,N_4193);
nand U4299 (N_4299,N_4120,N_4192);
and U4300 (N_4300,N_4011,N_4148);
xnor U4301 (N_4301,N_4029,N_4191);
nand U4302 (N_4302,N_4110,N_4116);
xnor U4303 (N_4303,N_4032,N_4033);
and U4304 (N_4304,N_4135,N_4021);
nand U4305 (N_4305,N_4028,N_4169);
and U4306 (N_4306,N_4193,N_4018);
nor U4307 (N_4307,N_4021,N_4011);
or U4308 (N_4308,N_4088,N_4175);
or U4309 (N_4309,N_4042,N_4115);
nor U4310 (N_4310,N_4040,N_4105);
nor U4311 (N_4311,N_4185,N_4079);
and U4312 (N_4312,N_4132,N_4115);
nor U4313 (N_4313,N_4115,N_4054);
nor U4314 (N_4314,N_4049,N_4165);
nand U4315 (N_4315,N_4196,N_4134);
nor U4316 (N_4316,N_4093,N_4129);
nand U4317 (N_4317,N_4111,N_4125);
nand U4318 (N_4318,N_4062,N_4005);
or U4319 (N_4319,N_4074,N_4061);
xnor U4320 (N_4320,N_4167,N_4178);
and U4321 (N_4321,N_4062,N_4151);
nor U4322 (N_4322,N_4005,N_4157);
nand U4323 (N_4323,N_4127,N_4045);
and U4324 (N_4324,N_4105,N_4086);
xnor U4325 (N_4325,N_4153,N_4095);
nand U4326 (N_4326,N_4114,N_4040);
or U4327 (N_4327,N_4139,N_4187);
xnor U4328 (N_4328,N_4054,N_4057);
xor U4329 (N_4329,N_4157,N_4079);
xnor U4330 (N_4330,N_4042,N_4166);
and U4331 (N_4331,N_4053,N_4066);
or U4332 (N_4332,N_4118,N_4100);
or U4333 (N_4333,N_4178,N_4097);
nand U4334 (N_4334,N_4060,N_4096);
and U4335 (N_4335,N_4022,N_4167);
nor U4336 (N_4336,N_4003,N_4171);
and U4337 (N_4337,N_4128,N_4008);
or U4338 (N_4338,N_4119,N_4147);
and U4339 (N_4339,N_4027,N_4174);
nand U4340 (N_4340,N_4166,N_4012);
or U4341 (N_4341,N_4169,N_4186);
and U4342 (N_4342,N_4006,N_4078);
and U4343 (N_4343,N_4032,N_4085);
and U4344 (N_4344,N_4196,N_4141);
xor U4345 (N_4345,N_4169,N_4087);
or U4346 (N_4346,N_4025,N_4042);
nand U4347 (N_4347,N_4014,N_4096);
and U4348 (N_4348,N_4134,N_4056);
and U4349 (N_4349,N_4191,N_4178);
and U4350 (N_4350,N_4060,N_4068);
nor U4351 (N_4351,N_4113,N_4118);
xor U4352 (N_4352,N_4163,N_4028);
nor U4353 (N_4353,N_4068,N_4065);
nor U4354 (N_4354,N_4032,N_4095);
and U4355 (N_4355,N_4004,N_4167);
and U4356 (N_4356,N_4174,N_4091);
nand U4357 (N_4357,N_4131,N_4125);
or U4358 (N_4358,N_4001,N_4173);
nand U4359 (N_4359,N_4120,N_4154);
or U4360 (N_4360,N_4110,N_4038);
or U4361 (N_4361,N_4157,N_4042);
nor U4362 (N_4362,N_4173,N_4094);
xnor U4363 (N_4363,N_4160,N_4120);
nor U4364 (N_4364,N_4104,N_4191);
nor U4365 (N_4365,N_4026,N_4042);
or U4366 (N_4366,N_4003,N_4023);
or U4367 (N_4367,N_4142,N_4151);
and U4368 (N_4368,N_4059,N_4061);
nand U4369 (N_4369,N_4042,N_4050);
nand U4370 (N_4370,N_4181,N_4016);
nand U4371 (N_4371,N_4169,N_4009);
xnor U4372 (N_4372,N_4059,N_4120);
and U4373 (N_4373,N_4070,N_4137);
and U4374 (N_4374,N_4103,N_4157);
and U4375 (N_4375,N_4121,N_4002);
nor U4376 (N_4376,N_4099,N_4129);
or U4377 (N_4377,N_4048,N_4081);
nand U4378 (N_4378,N_4116,N_4090);
or U4379 (N_4379,N_4099,N_4181);
nor U4380 (N_4380,N_4046,N_4074);
or U4381 (N_4381,N_4072,N_4171);
nand U4382 (N_4382,N_4152,N_4140);
nor U4383 (N_4383,N_4158,N_4009);
nor U4384 (N_4384,N_4151,N_4057);
nand U4385 (N_4385,N_4145,N_4115);
nand U4386 (N_4386,N_4014,N_4114);
and U4387 (N_4387,N_4055,N_4128);
or U4388 (N_4388,N_4026,N_4180);
or U4389 (N_4389,N_4076,N_4017);
or U4390 (N_4390,N_4144,N_4039);
nand U4391 (N_4391,N_4172,N_4148);
nor U4392 (N_4392,N_4077,N_4091);
and U4393 (N_4393,N_4021,N_4152);
and U4394 (N_4394,N_4165,N_4025);
nor U4395 (N_4395,N_4123,N_4071);
or U4396 (N_4396,N_4032,N_4011);
nand U4397 (N_4397,N_4144,N_4117);
and U4398 (N_4398,N_4125,N_4102);
or U4399 (N_4399,N_4114,N_4166);
and U4400 (N_4400,N_4342,N_4336);
or U4401 (N_4401,N_4317,N_4314);
xnor U4402 (N_4402,N_4221,N_4270);
and U4403 (N_4403,N_4209,N_4361);
xor U4404 (N_4404,N_4331,N_4379);
and U4405 (N_4405,N_4367,N_4309);
and U4406 (N_4406,N_4234,N_4204);
nand U4407 (N_4407,N_4318,N_4358);
nor U4408 (N_4408,N_4246,N_4321);
or U4409 (N_4409,N_4232,N_4214);
nand U4410 (N_4410,N_4371,N_4264);
nand U4411 (N_4411,N_4368,N_4304);
nand U4412 (N_4412,N_4299,N_4308);
nand U4413 (N_4413,N_4260,N_4266);
and U4414 (N_4414,N_4273,N_4354);
and U4415 (N_4415,N_4230,N_4384);
nand U4416 (N_4416,N_4202,N_4286);
and U4417 (N_4417,N_4282,N_4377);
or U4418 (N_4418,N_4236,N_4280);
nand U4419 (N_4419,N_4330,N_4243);
or U4420 (N_4420,N_4364,N_4393);
nand U4421 (N_4421,N_4210,N_4378);
xor U4422 (N_4422,N_4238,N_4211);
nor U4423 (N_4423,N_4303,N_4240);
nand U4424 (N_4424,N_4271,N_4278);
nand U4425 (N_4425,N_4255,N_4279);
xor U4426 (N_4426,N_4227,N_4207);
or U4427 (N_4427,N_4373,N_4229);
nor U4428 (N_4428,N_4360,N_4383);
xnor U4429 (N_4429,N_4281,N_4294);
or U4430 (N_4430,N_4370,N_4355);
or U4431 (N_4431,N_4224,N_4313);
nor U4432 (N_4432,N_4352,N_4348);
nor U4433 (N_4433,N_4253,N_4349);
xnor U4434 (N_4434,N_4268,N_4375);
or U4435 (N_4435,N_4293,N_4263);
and U4436 (N_4436,N_4385,N_4212);
nand U4437 (N_4437,N_4285,N_4335);
nand U4438 (N_4438,N_4257,N_4269);
nor U4439 (N_4439,N_4256,N_4362);
nor U4440 (N_4440,N_4247,N_4341);
nand U4441 (N_4441,N_4295,N_4311);
and U4442 (N_4442,N_4220,N_4276);
nor U4443 (N_4443,N_4326,N_4283);
and U4444 (N_4444,N_4296,N_4325);
xnor U4445 (N_4445,N_4334,N_4218);
xnor U4446 (N_4446,N_4327,N_4213);
nand U4447 (N_4447,N_4252,N_4267);
nor U4448 (N_4448,N_4366,N_4392);
xor U4449 (N_4449,N_4201,N_4292);
nand U4450 (N_4450,N_4231,N_4237);
xnor U4451 (N_4451,N_4217,N_4215);
nor U4452 (N_4452,N_4245,N_4225);
nand U4453 (N_4453,N_4332,N_4391);
and U4454 (N_4454,N_4346,N_4275);
and U4455 (N_4455,N_4388,N_4259);
and U4456 (N_4456,N_4301,N_4387);
and U4457 (N_4457,N_4249,N_4380);
nor U4458 (N_4458,N_4251,N_4297);
nor U4459 (N_4459,N_4395,N_4343);
xor U4460 (N_4460,N_4351,N_4329);
nor U4461 (N_4461,N_4200,N_4356);
or U4462 (N_4462,N_4262,N_4381);
nand U4463 (N_4463,N_4310,N_4265);
nor U4464 (N_4464,N_4382,N_4248);
nor U4465 (N_4465,N_4250,N_4219);
and U4466 (N_4466,N_4222,N_4372);
nand U4467 (N_4467,N_4376,N_4386);
nand U4468 (N_4468,N_4261,N_4398);
or U4469 (N_4469,N_4307,N_4345);
nor U4470 (N_4470,N_4289,N_4272);
or U4471 (N_4471,N_4233,N_4205);
nor U4472 (N_4472,N_4337,N_4396);
nand U4473 (N_4473,N_4223,N_4340);
and U4474 (N_4474,N_4369,N_4365);
nor U4475 (N_4475,N_4390,N_4288);
nor U4476 (N_4476,N_4274,N_4322);
nand U4477 (N_4477,N_4298,N_4235);
or U4478 (N_4478,N_4357,N_4239);
and U4479 (N_4479,N_4312,N_4258);
and U4480 (N_4480,N_4284,N_4320);
xnor U4481 (N_4481,N_4359,N_4350);
or U4482 (N_4482,N_4305,N_4300);
xor U4483 (N_4483,N_4287,N_4344);
nor U4484 (N_4484,N_4302,N_4324);
nor U4485 (N_4485,N_4339,N_4397);
and U4486 (N_4486,N_4363,N_4228);
nand U4487 (N_4487,N_4290,N_4306);
xor U4488 (N_4488,N_4277,N_4208);
nand U4489 (N_4489,N_4328,N_4241);
nor U4490 (N_4490,N_4353,N_4389);
and U4491 (N_4491,N_4333,N_4291);
nor U4492 (N_4492,N_4394,N_4226);
or U4493 (N_4493,N_4206,N_4203);
nor U4494 (N_4494,N_4319,N_4315);
nor U4495 (N_4495,N_4254,N_4216);
nand U4496 (N_4496,N_4244,N_4399);
or U4497 (N_4497,N_4338,N_4242);
and U4498 (N_4498,N_4347,N_4316);
or U4499 (N_4499,N_4323,N_4374);
and U4500 (N_4500,N_4219,N_4274);
and U4501 (N_4501,N_4228,N_4247);
and U4502 (N_4502,N_4240,N_4236);
or U4503 (N_4503,N_4254,N_4363);
nor U4504 (N_4504,N_4266,N_4258);
or U4505 (N_4505,N_4302,N_4391);
nor U4506 (N_4506,N_4354,N_4275);
nand U4507 (N_4507,N_4396,N_4283);
xor U4508 (N_4508,N_4289,N_4227);
and U4509 (N_4509,N_4370,N_4379);
and U4510 (N_4510,N_4239,N_4320);
or U4511 (N_4511,N_4229,N_4359);
or U4512 (N_4512,N_4362,N_4357);
or U4513 (N_4513,N_4375,N_4249);
nand U4514 (N_4514,N_4213,N_4320);
xor U4515 (N_4515,N_4380,N_4344);
nor U4516 (N_4516,N_4207,N_4274);
nor U4517 (N_4517,N_4235,N_4398);
or U4518 (N_4518,N_4314,N_4338);
nor U4519 (N_4519,N_4233,N_4379);
and U4520 (N_4520,N_4204,N_4388);
nand U4521 (N_4521,N_4317,N_4321);
and U4522 (N_4522,N_4397,N_4253);
or U4523 (N_4523,N_4305,N_4378);
and U4524 (N_4524,N_4375,N_4349);
nor U4525 (N_4525,N_4376,N_4341);
and U4526 (N_4526,N_4256,N_4235);
and U4527 (N_4527,N_4223,N_4241);
or U4528 (N_4528,N_4216,N_4219);
nand U4529 (N_4529,N_4348,N_4329);
or U4530 (N_4530,N_4356,N_4304);
nand U4531 (N_4531,N_4338,N_4277);
nand U4532 (N_4532,N_4279,N_4354);
or U4533 (N_4533,N_4235,N_4269);
and U4534 (N_4534,N_4204,N_4380);
and U4535 (N_4535,N_4208,N_4396);
nand U4536 (N_4536,N_4367,N_4315);
xnor U4537 (N_4537,N_4328,N_4396);
nand U4538 (N_4538,N_4321,N_4397);
nor U4539 (N_4539,N_4370,N_4325);
nand U4540 (N_4540,N_4301,N_4275);
nand U4541 (N_4541,N_4342,N_4323);
and U4542 (N_4542,N_4376,N_4379);
and U4543 (N_4543,N_4398,N_4384);
xor U4544 (N_4544,N_4377,N_4206);
nor U4545 (N_4545,N_4234,N_4322);
nor U4546 (N_4546,N_4328,N_4283);
nand U4547 (N_4547,N_4386,N_4277);
xnor U4548 (N_4548,N_4258,N_4203);
nand U4549 (N_4549,N_4243,N_4360);
or U4550 (N_4550,N_4259,N_4284);
nor U4551 (N_4551,N_4238,N_4272);
nor U4552 (N_4552,N_4207,N_4203);
or U4553 (N_4553,N_4206,N_4325);
nand U4554 (N_4554,N_4232,N_4305);
xnor U4555 (N_4555,N_4289,N_4352);
or U4556 (N_4556,N_4282,N_4311);
xnor U4557 (N_4557,N_4259,N_4209);
nor U4558 (N_4558,N_4343,N_4289);
nand U4559 (N_4559,N_4243,N_4204);
or U4560 (N_4560,N_4361,N_4383);
or U4561 (N_4561,N_4382,N_4211);
nor U4562 (N_4562,N_4201,N_4210);
or U4563 (N_4563,N_4305,N_4329);
or U4564 (N_4564,N_4317,N_4223);
xor U4565 (N_4565,N_4373,N_4393);
or U4566 (N_4566,N_4274,N_4349);
or U4567 (N_4567,N_4306,N_4326);
nand U4568 (N_4568,N_4338,N_4226);
xnor U4569 (N_4569,N_4288,N_4370);
or U4570 (N_4570,N_4236,N_4296);
nand U4571 (N_4571,N_4213,N_4205);
nand U4572 (N_4572,N_4218,N_4350);
nand U4573 (N_4573,N_4329,N_4325);
nor U4574 (N_4574,N_4219,N_4207);
and U4575 (N_4575,N_4256,N_4233);
nor U4576 (N_4576,N_4331,N_4346);
or U4577 (N_4577,N_4271,N_4276);
xnor U4578 (N_4578,N_4274,N_4214);
nor U4579 (N_4579,N_4280,N_4210);
nor U4580 (N_4580,N_4231,N_4215);
xnor U4581 (N_4581,N_4309,N_4254);
nand U4582 (N_4582,N_4291,N_4378);
or U4583 (N_4583,N_4327,N_4210);
and U4584 (N_4584,N_4282,N_4234);
nand U4585 (N_4585,N_4388,N_4345);
or U4586 (N_4586,N_4224,N_4254);
or U4587 (N_4587,N_4305,N_4335);
nand U4588 (N_4588,N_4380,N_4339);
and U4589 (N_4589,N_4259,N_4327);
and U4590 (N_4590,N_4367,N_4222);
and U4591 (N_4591,N_4351,N_4259);
or U4592 (N_4592,N_4212,N_4381);
or U4593 (N_4593,N_4296,N_4350);
and U4594 (N_4594,N_4295,N_4276);
or U4595 (N_4595,N_4326,N_4222);
and U4596 (N_4596,N_4369,N_4377);
nor U4597 (N_4597,N_4281,N_4259);
nor U4598 (N_4598,N_4287,N_4211);
and U4599 (N_4599,N_4216,N_4208);
or U4600 (N_4600,N_4407,N_4594);
nand U4601 (N_4601,N_4494,N_4546);
xnor U4602 (N_4602,N_4482,N_4503);
or U4603 (N_4603,N_4458,N_4457);
nand U4604 (N_4604,N_4590,N_4505);
nand U4605 (N_4605,N_4549,N_4571);
nor U4606 (N_4606,N_4514,N_4422);
or U4607 (N_4607,N_4557,N_4472);
nor U4608 (N_4608,N_4499,N_4525);
or U4609 (N_4609,N_4544,N_4403);
nand U4610 (N_4610,N_4412,N_4461);
or U4611 (N_4611,N_4535,N_4460);
nor U4612 (N_4612,N_4483,N_4405);
and U4613 (N_4613,N_4596,N_4523);
nand U4614 (N_4614,N_4443,N_4400);
nor U4615 (N_4615,N_4495,N_4589);
nand U4616 (N_4616,N_4498,N_4513);
or U4617 (N_4617,N_4552,N_4473);
or U4618 (N_4618,N_4551,N_4532);
or U4619 (N_4619,N_4444,N_4423);
or U4620 (N_4620,N_4517,N_4441);
nor U4621 (N_4621,N_4559,N_4575);
and U4622 (N_4622,N_4468,N_4593);
or U4623 (N_4623,N_4521,N_4566);
xnor U4624 (N_4624,N_4480,N_4475);
nor U4625 (N_4625,N_4582,N_4402);
xnor U4626 (N_4626,N_4538,N_4406);
nand U4627 (N_4627,N_4516,N_4476);
nor U4628 (N_4628,N_4564,N_4448);
or U4629 (N_4629,N_4567,N_4466);
or U4630 (N_4630,N_4536,N_4592);
nor U4631 (N_4631,N_4562,N_4428);
or U4632 (N_4632,N_4479,N_4464);
and U4633 (N_4633,N_4452,N_4417);
xor U4634 (N_4634,N_4580,N_4599);
and U4635 (N_4635,N_4573,N_4435);
or U4636 (N_4636,N_4539,N_4509);
or U4637 (N_4637,N_4433,N_4486);
and U4638 (N_4638,N_4547,N_4508);
or U4639 (N_4639,N_4426,N_4478);
nand U4640 (N_4640,N_4543,N_4447);
and U4641 (N_4641,N_4431,N_4568);
nand U4642 (N_4642,N_4404,N_4492);
nor U4643 (N_4643,N_4463,N_4484);
xnor U4644 (N_4644,N_4556,N_4462);
nand U4645 (N_4645,N_4455,N_4507);
nor U4646 (N_4646,N_4453,N_4579);
nand U4647 (N_4647,N_4519,N_4491);
nand U4648 (N_4648,N_4572,N_4489);
nor U4649 (N_4649,N_4563,N_4548);
nand U4650 (N_4650,N_4511,N_4595);
nor U4651 (N_4651,N_4555,N_4429);
and U4652 (N_4652,N_4526,N_4597);
nand U4653 (N_4653,N_4474,N_4533);
or U4654 (N_4654,N_4554,N_4530);
nor U4655 (N_4655,N_4527,N_4424);
or U4656 (N_4656,N_4588,N_4454);
nor U4657 (N_4657,N_4477,N_4410);
or U4658 (N_4658,N_4459,N_4471);
nand U4659 (N_4659,N_4541,N_4550);
nand U4660 (N_4660,N_4416,N_4467);
or U4661 (N_4661,N_4570,N_4581);
or U4662 (N_4662,N_4577,N_4419);
or U4663 (N_4663,N_4487,N_4500);
nand U4664 (N_4664,N_4502,N_4438);
and U4665 (N_4665,N_4470,N_4427);
and U4666 (N_4666,N_4411,N_4430);
or U4667 (N_4667,N_4560,N_4565);
nor U4668 (N_4668,N_4481,N_4506);
nand U4669 (N_4669,N_4488,N_4520);
nor U4670 (N_4670,N_4576,N_4425);
nand U4671 (N_4671,N_4583,N_4445);
or U4672 (N_4672,N_4465,N_4409);
nor U4673 (N_4673,N_4542,N_4584);
nor U4674 (N_4674,N_4469,N_4432);
or U4675 (N_4675,N_4531,N_4558);
nand U4676 (N_4676,N_4518,N_4450);
and U4677 (N_4677,N_4540,N_4586);
or U4678 (N_4678,N_4436,N_4537);
nand U4679 (N_4679,N_4497,N_4534);
or U4680 (N_4680,N_4493,N_4449);
xnor U4681 (N_4681,N_4529,N_4578);
xnor U4682 (N_4682,N_4442,N_4598);
and U4683 (N_4683,N_4420,N_4415);
nand U4684 (N_4684,N_4408,N_4587);
and U4685 (N_4685,N_4413,N_4451);
or U4686 (N_4686,N_4434,N_4439);
nand U4687 (N_4687,N_4485,N_4522);
nor U4688 (N_4688,N_4591,N_4561);
nor U4689 (N_4689,N_4524,N_4515);
and U4690 (N_4690,N_4553,N_4545);
and U4691 (N_4691,N_4414,N_4585);
and U4692 (N_4692,N_4446,N_4574);
nor U4693 (N_4693,N_4418,N_4456);
xor U4694 (N_4694,N_4440,N_4512);
nand U4695 (N_4695,N_4510,N_4421);
nand U4696 (N_4696,N_4501,N_4437);
or U4697 (N_4697,N_4569,N_4528);
nand U4698 (N_4698,N_4504,N_4401);
nand U4699 (N_4699,N_4490,N_4496);
nor U4700 (N_4700,N_4453,N_4498);
or U4701 (N_4701,N_4400,N_4552);
nand U4702 (N_4702,N_4494,N_4410);
or U4703 (N_4703,N_4579,N_4472);
and U4704 (N_4704,N_4533,N_4428);
and U4705 (N_4705,N_4566,N_4450);
or U4706 (N_4706,N_4569,N_4436);
and U4707 (N_4707,N_4575,N_4538);
nand U4708 (N_4708,N_4548,N_4572);
and U4709 (N_4709,N_4453,N_4531);
and U4710 (N_4710,N_4483,N_4495);
xor U4711 (N_4711,N_4589,N_4559);
nor U4712 (N_4712,N_4434,N_4411);
and U4713 (N_4713,N_4540,N_4556);
nand U4714 (N_4714,N_4528,N_4487);
nand U4715 (N_4715,N_4439,N_4454);
nand U4716 (N_4716,N_4494,N_4416);
nor U4717 (N_4717,N_4541,N_4504);
xnor U4718 (N_4718,N_4401,N_4435);
or U4719 (N_4719,N_4462,N_4591);
nand U4720 (N_4720,N_4455,N_4543);
nand U4721 (N_4721,N_4443,N_4577);
nor U4722 (N_4722,N_4460,N_4434);
and U4723 (N_4723,N_4465,N_4492);
nor U4724 (N_4724,N_4530,N_4574);
nor U4725 (N_4725,N_4468,N_4560);
xnor U4726 (N_4726,N_4515,N_4442);
or U4727 (N_4727,N_4486,N_4541);
nand U4728 (N_4728,N_4557,N_4599);
nor U4729 (N_4729,N_4506,N_4443);
or U4730 (N_4730,N_4466,N_4408);
and U4731 (N_4731,N_4582,N_4430);
and U4732 (N_4732,N_4535,N_4592);
nand U4733 (N_4733,N_4526,N_4513);
xnor U4734 (N_4734,N_4514,N_4411);
and U4735 (N_4735,N_4550,N_4508);
or U4736 (N_4736,N_4477,N_4454);
or U4737 (N_4737,N_4424,N_4503);
nand U4738 (N_4738,N_4409,N_4509);
and U4739 (N_4739,N_4475,N_4543);
nand U4740 (N_4740,N_4462,N_4584);
xnor U4741 (N_4741,N_4470,N_4414);
nor U4742 (N_4742,N_4441,N_4529);
or U4743 (N_4743,N_4430,N_4458);
nor U4744 (N_4744,N_4507,N_4480);
nor U4745 (N_4745,N_4426,N_4403);
nand U4746 (N_4746,N_4558,N_4590);
nor U4747 (N_4747,N_4466,N_4450);
nand U4748 (N_4748,N_4410,N_4483);
or U4749 (N_4749,N_4400,N_4546);
and U4750 (N_4750,N_4468,N_4503);
and U4751 (N_4751,N_4575,N_4567);
nor U4752 (N_4752,N_4478,N_4544);
or U4753 (N_4753,N_4558,N_4475);
or U4754 (N_4754,N_4531,N_4469);
or U4755 (N_4755,N_4492,N_4535);
nand U4756 (N_4756,N_4567,N_4598);
nor U4757 (N_4757,N_4437,N_4523);
or U4758 (N_4758,N_4512,N_4496);
nor U4759 (N_4759,N_4466,N_4418);
nand U4760 (N_4760,N_4586,N_4416);
and U4761 (N_4761,N_4419,N_4584);
and U4762 (N_4762,N_4584,N_4441);
or U4763 (N_4763,N_4595,N_4478);
nand U4764 (N_4764,N_4468,N_4426);
nand U4765 (N_4765,N_4471,N_4402);
nand U4766 (N_4766,N_4493,N_4457);
and U4767 (N_4767,N_4529,N_4404);
xor U4768 (N_4768,N_4425,N_4417);
and U4769 (N_4769,N_4403,N_4512);
nand U4770 (N_4770,N_4545,N_4589);
nand U4771 (N_4771,N_4549,N_4459);
nand U4772 (N_4772,N_4439,N_4458);
or U4773 (N_4773,N_4586,N_4566);
nand U4774 (N_4774,N_4598,N_4564);
nand U4775 (N_4775,N_4420,N_4574);
nor U4776 (N_4776,N_4447,N_4435);
nand U4777 (N_4777,N_4548,N_4488);
or U4778 (N_4778,N_4517,N_4526);
nor U4779 (N_4779,N_4584,N_4595);
nor U4780 (N_4780,N_4520,N_4430);
nor U4781 (N_4781,N_4433,N_4530);
and U4782 (N_4782,N_4466,N_4597);
nand U4783 (N_4783,N_4437,N_4511);
or U4784 (N_4784,N_4500,N_4559);
nand U4785 (N_4785,N_4543,N_4480);
or U4786 (N_4786,N_4507,N_4531);
xnor U4787 (N_4787,N_4503,N_4580);
nor U4788 (N_4788,N_4553,N_4475);
nor U4789 (N_4789,N_4527,N_4469);
nor U4790 (N_4790,N_4599,N_4594);
nor U4791 (N_4791,N_4555,N_4511);
or U4792 (N_4792,N_4580,N_4437);
nand U4793 (N_4793,N_4488,N_4446);
and U4794 (N_4794,N_4518,N_4527);
nand U4795 (N_4795,N_4466,N_4479);
nor U4796 (N_4796,N_4509,N_4432);
and U4797 (N_4797,N_4433,N_4594);
nor U4798 (N_4798,N_4452,N_4538);
xnor U4799 (N_4799,N_4567,N_4430);
and U4800 (N_4800,N_4656,N_4784);
nand U4801 (N_4801,N_4693,N_4663);
nor U4802 (N_4802,N_4670,N_4654);
and U4803 (N_4803,N_4721,N_4671);
or U4804 (N_4804,N_4692,N_4638);
nor U4805 (N_4805,N_4660,N_4715);
nor U4806 (N_4806,N_4706,N_4792);
or U4807 (N_4807,N_4610,N_4606);
nand U4808 (N_4808,N_4644,N_4748);
or U4809 (N_4809,N_4636,N_4783);
nand U4810 (N_4810,N_4680,N_4623);
and U4811 (N_4811,N_4752,N_4666);
nor U4812 (N_4812,N_4705,N_4684);
nand U4813 (N_4813,N_4642,N_4697);
or U4814 (N_4814,N_4796,N_4719);
nor U4815 (N_4815,N_4790,N_4678);
or U4816 (N_4816,N_4708,N_4793);
nor U4817 (N_4817,N_4758,N_4755);
or U4818 (N_4818,N_4676,N_4789);
nor U4819 (N_4819,N_4608,N_4648);
or U4820 (N_4820,N_4627,N_4720);
or U4821 (N_4821,N_4780,N_4767);
nor U4822 (N_4822,N_4762,N_4728);
xor U4823 (N_4823,N_4735,N_4731);
nand U4824 (N_4824,N_4640,N_4659);
and U4825 (N_4825,N_4766,N_4723);
or U4826 (N_4826,N_4774,N_4739);
or U4827 (N_4827,N_4702,N_4617);
and U4828 (N_4828,N_4629,N_4730);
or U4829 (N_4829,N_4717,N_4622);
nand U4830 (N_4830,N_4737,N_4611);
and U4831 (N_4831,N_4729,N_4794);
and U4832 (N_4832,N_4782,N_4797);
and U4833 (N_4833,N_4616,N_4649);
xnor U4834 (N_4834,N_4677,N_4734);
and U4835 (N_4835,N_4637,N_4685);
or U4836 (N_4836,N_4612,N_4750);
and U4837 (N_4837,N_4768,N_4679);
nand U4838 (N_4838,N_4691,N_4603);
nor U4839 (N_4839,N_4736,N_4672);
or U4840 (N_4840,N_4615,N_4652);
nand U4841 (N_4841,N_4760,N_4632);
xnor U4842 (N_4842,N_4740,N_4700);
or U4843 (N_4843,N_4624,N_4669);
nor U4844 (N_4844,N_4694,N_4744);
or U4845 (N_4845,N_4620,N_4714);
nand U4846 (N_4846,N_4698,N_4711);
or U4847 (N_4847,N_4618,N_4635);
nor U4848 (N_4848,N_4732,N_4749);
and U4849 (N_4849,N_4746,N_4709);
or U4850 (N_4850,N_4772,N_4621);
nand U4851 (N_4851,N_4764,N_4619);
nand U4852 (N_4852,N_4742,N_4687);
and U4853 (N_4853,N_4724,N_4609);
nand U4854 (N_4854,N_4759,N_4614);
or U4855 (N_4855,N_4773,N_4605);
xor U4856 (N_4856,N_4795,N_4765);
and U4857 (N_4857,N_4668,N_4645);
or U4858 (N_4858,N_4798,N_4696);
nand U4859 (N_4859,N_4761,N_4630);
xnor U4860 (N_4860,N_4776,N_4665);
or U4861 (N_4861,N_4655,N_4602);
and U4862 (N_4862,N_4770,N_4754);
nor U4863 (N_4863,N_4653,N_4788);
nor U4864 (N_4864,N_4707,N_4778);
and U4865 (N_4865,N_4777,N_4681);
and U4866 (N_4866,N_4771,N_4787);
xor U4867 (N_4867,N_4633,N_4704);
xnor U4868 (N_4868,N_4718,N_4799);
nand U4869 (N_4869,N_4791,N_4607);
nor U4870 (N_4870,N_4674,N_4639);
xor U4871 (N_4871,N_4662,N_4786);
or U4872 (N_4872,N_4745,N_4647);
nor U4873 (N_4873,N_4625,N_4601);
or U4874 (N_4874,N_4689,N_4743);
and U4875 (N_4875,N_4600,N_4710);
or U4876 (N_4876,N_4650,N_4667);
or U4877 (N_4877,N_4695,N_4683);
nand U4878 (N_4878,N_4713,N_4741);
xnor U4879 (N_4879,N_4775,N_4733);
nand U4880 (N_4880,N_4634,N_4781);
or U4881 (N_4881,N_4628,N_4701);
and U4882 (N_4882,N_4726,N_4722);
and U4883 (N_4883,N_4613,N_4769);
nand U4884 (N_4884,N_4626,N_4712);
xnor U4885 (N_4885,N_4688,N_4753);
or U4886 (N_4886,N_4747,N_4725);
and U4887 (N_4887,N_4716,N_4738);
and U4888 (N_4888,N_4673,N_4646);
nand U4889 (N_4889,N_4785,N_4682);
nand U4890 (N_4890,N_4703,N_4658);
or U4891 (N_4891,N_4657,N_4641);
and U4892 (N_4892,N_4631,N_4690);
or U4893 (N_4893,N_4699,N_4757);
nand U4894 (N_4894,N_4675,N_4664);
nor U4895 (N_4895,N_4779,N_4686);
nor U4896 (N_4896,N_4727,N_4751);
or U4897 (N_4897,N_4661,N_4756);
nand U4898 (N_4898,N_4643,N_4763);
and U4899 (N_4899,N_4651,N_4604);
and U4900 (N_4900,N_4714,N_4786);
and U4901 (N_4901,N_4636,N_4748);
nor U4902 (N_4902,N_4734,N_4657);
or U4903 (N_4903,N_4705,N_4766);
nand U4904 (N_4904,N_4607,N_4737);
or U4905 (N_4905,N_4747,N_4627);
nor U4906 (N_4906,N_4657,N_4619);
nand U4907 (N_4907,N_4792,N_4781);
and U4908 (N_4908,N_4726,N_4601);
nor U4909 (N_4909,N_4624,N_4675);
and U4910 (N_4910,N_4797,N_4764);
nor U4911 (N_4911,N_4709,N_4616);
and U4912 (N_4912,N_4786,N_4620);
nand U4913 (N_4913,N_4735,N_4696);
nand U4914 (N_4914,N_4746,N_4660);
and U4915 (N_4915,N_4794,N_4759);
nand U4916 (N_4916,N_4714,N_4631);
and U4917 (N_4917,N_4770,N_4682);
or U4918 (N_4918,N_4724,N_4715);
or U4919 (N_4919,N_4605,N_4758);
nand U4920 (N_4920,N_4775,N_4631);
and U4921 (N_4921,N_4606,N_4786);
nand U4922 (N_4922,N_4651,N_4770);
nor U4923 (N_4923,N_4751,N_4760);
or U4924 (N_4924,N_4720,N_4709);
nor U4925 (N_4925,N_4616,N_4739);
nand U4926 (N_4926,N_4737,N_4629);
and U4927 (N_4927,N_4674,N_4726);
nand U4928 (N_4928,N_4716,N_4731);
xnor U4929 (N_4929,N_4612,N_4774);
nor U4930 (N_4930,N_4736,N_4746);
nor U4931 (N_4931,N_4759,N_4608);
or U4932 (N_4932,N_4789,N_4619);
nor U4933 (N_4933,N_4708,N_4765);
nand U4934 (N_4934,N_4604,N_4734);
or U4935 (N_4935,N_4634,N_4730);
nand U4936 (N_4936,N_4605,N_4696);
and U4937 (N_4937,N_4798,N_4703);
nor U4938 (N_4938,N_4753,N_4786);
or U4939 (N_4939,N_4738,N_4635);
or U4940 (N_4940,N_4779,N_4618);
xnor U4941 (N_4941,N_4780,N_4792);
nand U4942 (N_4942,N_4753,N_4694);
or U4943 (N_4943,N_4675,N_4788);
nand U4944 (N_4944,N_4769,N_4659);
nand U4945 (N_4945,N_4742,N_4780);
and U4946 (N_4946,N_4734,N_4730);
or U4947 (N_4947,N_4772,N_4724);
nor U4948 (N_4948,N_4624,N_4720);
nand U4949 (N_4949,N_4647,N_4747);
nor U4950 (N_4950,N_4758,N_4721);
or U4951 (N_4951,N_4688,N_4774);
or U4952 (N_4952,N_4745,N_4620);
or U4953 (N_4953,N_4728,N_4791);
nand U4954 (N_4954,N_4733,N_4618);
and U4955 (N_4955,N_4700,N_4769);
or U4956 (N_4956,N_4720,N_4649);
or U4957 (N_4957,N_4681,N_4612);
nand U4958 (N_4958,N_4714,N_4690);
or U4959 (N_4959,N_4715,N_4696);
nand U4960 (N_4960,N_4692,N_4683);
nand U4961 (N_4961,N_4661,N_4770);
and U4962 (N_4962,N_4720,N_4770);
nor U4963 (N_4963,N_4730,N_4684);
nor U4964 (N_4964,N_4793,N_4778);
nand U4965 (N_4965,N_4657,N_4659);
and U4966 (N_4966,N_4727,N_4604);
xor U4967 (N_4967,N_4779,N_4769);
nand U4968 (N_4968,N_4758,N_4772);
nor U4969 (N_4969,N_4774,N_4694);
nand U4970 (N_4970,N_4610,N_4604);
nand U4971 (N_4971,N_4645,N_4768);
nand U4972 (N_4972,N_4684,N_4628);
nor U4973 (N_4973,N_4757,N_4659);
nor U4974 (N_4974,N_4709,N_4656);
xor U4975 (N_4975,N_4760,N_4675);
and U4976 (N_4976,N_4628,N_4788);
or U4977 (N_4977,N_4767,N_4728);
nand U4978 (N_4978,N_4658,N_4655);
and U4979 (N_4979,N_4628,N_4764);
or U4980 (N_4980,N_4626,N_4795);
and U4981 (N_4981,N_4613,N_4751);
nor U4982 (N_4982,N_4642,N_4799);
nand U4983 (N_4983,N_4703,N_4742);
xor U4984 (N_4984,N_4703,N_4752);
nand U4985 (N_4985,N_4664,N_4618);
nor U4986 (N_4986,N_4748,N_4784);
nor U4987 (N_4987,N_4769,N_4797);
xnor U4988 (N_4988,N_4606,N_4602);
or U4989 (N_4989,N_4785,N_4763);
or U4990 (N_4990,N_4701,N_4757);
or U4991 (N_4991,N_4674,N_4622);
nand U4992 (N_4992,N_4636,N_4714);
nand U4993 (N_4993,N_4771,N_4790);
nor U4994 (N_4994,N_4600,N_4647);
or U4995 (N_4995,N_4628,N_4668);
xnor U4996 (N_4996,N_4740,N_4634);
nand U4997 (N_4997,N_4766,N_4720);
or U4998 (N_4998,N_4780,N_4620);
or U4999 (N_4999,N_4690,N_4757);
and U5000 (N_5000,N_4859,N_4829);
and U5001 (N_5001,N_4836,N_4920);
or U5002 (N_5002,N_4833,N_4997);
or U5003 (N_5003,N_4953,N_4895);
nor U5004 (N_5004,N_4897,N_4924);
or U5005 (N_5005,N_4929,N_4881);
and U5006 (N_5006,N_4839,N_4978);
and U5007 (N_5007,N_4800,N_4838);
nor U5008 (N_5008,N_4828,N_4840);
nand U5009 (N_5009,N_4898,N_4979);
xnor U5010 (N_5010,N_4983,N_4863);
and U5011 (N_5011,N_4891,N_4821);
or U5012 (N_5012,N_4921,N_4827);
or U5013 (N_5013,N_4817,N_4893);
nand U5014 (N_5014,N_4906,N_4845);
nor U5015 (N_5015,N_4857,N_4855);
and U5016 (N_5016,N_4832,N_4938);
nor U5017 (N_5017,N_4972,N_4974);
nor U5018 (N_5018,N_4948,N_4903);
nand U5019 (N_5019,N_4804,N_4909);
xnor U5020 (N_5020,N_4888,N_4882);
and U5021 (N_5021,N_4914,N_4816);
and U5022 (N_5022,N_4968,N_4989);
and U5023 (N_5023,N_4981,N_4900);
nand U5024 (N_5024,N_4835,N_4995);
and U5025 (N_5025,N_4885,N_4904);
xnor U5026 (N_5026,N_4991,N_4907);
nand U5027 (N_5027,N_4826,N_4831);
or U5028 (N_5028,N_4962,N_4860);
and U5029 (N_5029,N_4858,N_4886);
nand U5030 (N_5030,N_4999,N_4889);
xnor U5031 (N_5031,N_4971,N_4915);
or U5032 (N_5032,N_4849,N_4823);
nand U5033 (N_5033,N_4892,N_4949);
xnor U5034 (N_5034,N_4925,N_4946);
and U5035 (N_5035,N_4861,N_4806);
nor U5036 (N_5036,N_4877,N_4865);
and U5037 (N_5037,N_4996,N_4864);
nor U5038 (N_5038,N_4967,N_4852);
nand U5039 (N_5039,N_4935,N_4950);
xnor U5040 (N_5040,N_4896,N_4808);
or U5041 (N_5041,N_4937,N_4847);
nor U5042 (N_5042,N_4809,N_4975);
or U5043 (N_5043,N_4956,N_4875);
nand U5044 (N_5044,N_4976,N_4854);
nand U5045 (N_5045,N_4912,N_4876);
or U5046 (N_5046,N_4952,N_4959);
nor U5047 (N_5047,N_4931,N_4830);
and U5048 (N_5048,N_4887,N_4998);
or U5049 (N_5049,N_4868,N_4862);
or U5050 (N_5050,N_4992,N_4943);
nand U5051 (N_5051,N_4807,N_4902);
nand U5052 (N_5052,N_4843,N_4936);
nor U5053 (N_5053,N_4918,N_4965);
or U5054 (N_5054,N_4872,N_4966);
nor U5055 (N_5055,N_4884,N_4805);
nand U5056 (N_5056,N_4987,N_4815);
or U5057 (N_5057,N_4947,N_4874);
and U5058 (N_5058,N_4811,N_4880);
and U5059 (N_5059,N_4867,N_4986);
nor U5060 (N_5060,N_4802,N_4942);
xnor U5061 (N_5061,N_4890,N_4837);
xnor U5062 (N_5062,N_4980,N_4970);
nand U5063 (N_5063,N_4848,N_4818);
xnor U5064 (N_5064,N_4955,N_4926);
or U5065 (N_5065,N_4982,N_4944);
nor U5066 (N_5066,N_4814,N_4825);
or U5067 (N_5067,N_4911,N_4941);
or U5068 (N_5068,N_4870,N_4810);
nor U5069 (N_5069,N_4913,N_4850);
or U5070 (N_5070,N_4939,N_4977);
xor U5071 (N_5071,N_4993,N_4969);
xor U5072 (N_5072,N_4908,N_4973);
xnor U5073 (N_5073,N_4985,N_4994);
nand U5074 (N_5074,N_4873,N_4813);
nor U5075 (N_5075,N_4899,N_4841);
nor U5076 (N_5076,N_4803,N_4923);
or U5077 (N_5077,N_4960,N_4834);
and U5078 (N_5078,N_4901,N_4961);
or U5079 (N_5079,N_4894,N_4984);
nand U5080 (N_5080,N_4842,N_4940);
and U5081 (N_5081,N_4846,N_4928);
or U5082 (N_5082,N_4917,N_4958);
xor U5083 (N_5083,N_4963,N_4934);
nand U5084 (N_5084,N_4822,N_4919);
nor U5085 (N_5085,N_4932,N_4945);
and U5086 (N_5086,N_4954,N_4905);
and U5087 (N_5087,N_4820,N_4883);
nor U5088 (N_5088,N_4819,N_4930);
and U5089 (N_5089,N_4824,N_4878);
and U5090 (N_5090,N_4853,N_4988);
or U5091 (N_5091,N_4951,N_4851);
or U5092 (N_5092,N_4844,N_4964);
nor U5093 (N_5093,N_4916,N_4910);
nor U5094 (N_5094,N_4869,N_4871);
nand U5095 (N_5095,N_4866,N_4933);
or U5096 (N_5096,N_4812,N_4879);
and U5097 (N_5097,N_4957,N_4990);
or U5098 (N_5098,N_4801,N_4927);
xor U5099 (N_5099,N_4922,N_4856);
and U5100 (N_5100,N_4970,N_4924);
or U5101 (N_5101,N_4856,N_4813);
xnor U5102 (N_5102,N_4851,N_4990);
and U5103 (N_5103,N_4890,N_4917);
and U5104 (N_5104,N_4893,N_4836);
nand U5105 (N_5105,N_4938,N_4838);
and U5106 (N_5106,N_4893,N_4966);
nand U5107 (N_5107,N_4929,N_4931);
nand U5108 (N_5108,N_4931,N_4961);
nor U5109 (N_5109,N_4805,N_4964);
nand U5110 (N_5110,N_4872,N_4851);
nand U5111 (N_5111,N_4952,N_4838);
nand U5112 (N_5112,N_4887,N_4840);
and U5113 (N_5113,N_4932,N_4967);
or U5114 (N_5114,N_4994,N_4843);
or U5115 (N_5115,N_4811,N_4992);
or U5116 (N_5116,N_4875,N_4857);
nor U5117 (N_5117,N_4818,N_4847);
xnor U5118 (N_5118,N_4855,N_4959);
and U5119 (N_5119,N_4963,N_4898);
nand U5120 (N_5120,N_4988,N_4852);
nor U5121 (N_5121,N_4996,N_4857);
and U5122 (N_5122,N_4976,N_4902);
nand U5123 (N_5123,N_4998,N_4864);
nand U5124 (N_5124,N_4827,N_4857);
nand U5125 (N_5125,N_4826,N_4850);
nand U5126 (N_5126,N_4950,N_4933);
or U5127 (N_5127,N_4990,N_4945);
and U5128 (N_5128,N_4813,N_4913);
nand U5129 (N_5129,N_4822,N_4869);
nor U5130 (N_5130,N_4998,N_4858);
nand U5131 (N_5131,N_4974,N_4981);
nor U5132 (N_5132,N_4964,N_4801);
nor U5133 (N_5133,N_4840,N_4869);
nand U5134 (N_5134,N_4832,N_4928);
or U5135 (N_5135,N_4906,N_4946);
nor U5136 (N_5136,N_4837,N_4957);
xor U5137 (N_5137,N_4971,N_4859);
or U5138 (N_5138,N_4849,N_4865);
and U5139 (N_5139,N_4997,N_4868);
nand U5140 (N_5140,N_4934,N_4942);
or U5141 (N_5141,N_4912,N_4961);
or U5142 (N_5142,N_4966,N_4923);
nor U5143 (N_5143,N_4921,N_4948);
nand U5144 (N_5144,N_4971,N_4959);
or U5145 (N_5145,N_4903,N_4997);
or U5146 (N_5146,N_4856,N_4901);
or U5147 (N_5147,N_4870,N_4984);
or U5148 (N_5148,N_4847,N_4855);
nor U5149 (N_5149,N_4819,N_4868);
nor U5150 (N_5150,N_4970,N_4899);
or U5151 (N_5151,N_4900,N_4817);
or U5152 (N_5152,N_4833,N_4973);
nor U5153 (N_5153,N_4997,N_4995);
and U5154 (N_5154,N_4812,N_4894);
nor U5155 (N_5155,N_4881,N_4837);
nand U5156 (N_5156,N_4867,N_4824);
and U5157 (N_5157,N_4824,N_4856);
or U5158 (N_5158,N_4928,N_4854);
and U5159 (N_5159,N_4816,N_4902);
nand U5160 (N_5160,N_4991,N_4968);
or U5161 (N_5161,N_4871,N_4929);
xnor U5162 (N_5162,N_4895,N_4866);
nand U5163 (N_5163,N_4867,N_4844);
or U5164 (N_5164,N_4813,N_4854);
and U5165 (N_5165,N_4891,N_4826);
nor U5166 (N_5166,N_4833,N_4827);
nor U5167 (N_5167,N_4830,N_4885);
and U5168 (N_5168,N_4919,N_4991);
xor U5169 (N_5169,N_4858,N_4991);
and U5170 (N_5170,N_4916,N_4979);
or U5171 (N_5171,N_4849,N_4890);
and U5172 (N_5172,N_4955,N_4908);
and U5173 (N_5173,N_4936,N_4902);
nor U5174 (N_5174,N_4978,N_4991);
or U5175 (N_5175,N_4850,N_4874);
or U5176 (N_5176,N_4872,N_4913);
or U5177 (N_5177,N_4986,N_4970);
and U5178 (N_5178,N_4897,N_4909);
and U5179 (N_5179,N_4963,N_4981);
xnor U5180 (N_5180,N_4817,N_4883);
xor U5181 (N_5181,N_4956,N_4998);
or U5182 (N_5182,N_4917,N_4870);
nand U5183 (N_5183,N_4981,N_4935);
and U5184 (N_5184,N_4821,N_4978);
nor U5185 (N_5185,N_4833,N_4852);
nor U5186 (N_5186,N_4927,N_4861);
nor U5187 (N_5187,N_4952,N_4873);
and U5188 (N_5188,N_4825,N_4847);
xor U5189 (N_5189,N_4875,N_4940);
nand U5190 (N_5190,N_4836,N_4906);
and U5191 (N_5191,N_4857,N_4989);
or U5192 (N_5192,N_4859,N_4977);
nand U5193 (N_5193,N_4820,N_4857);
nor U5194 (N_5194,N_4844,N_4941);
or U5195 (N_5195,N_4827,N_4849);
nand U5196 (N_5196,N_4822,N_4890);
nand U5197 (N_5197,N_4842,N_4921);
xnor U5198 (N_5198,N_4810,N_4808);
nor U5199 (N_5199,N_4944,N_4906);
nand U5200 (N_5200,N_5057,N_5087);
nor U5201 (N_5201,N_5167,N_5073);
and U5202 (N_5202,N_5126,N_5110);
nand U5203 (N_5203,N_5068,N_5078);
nand U5204 (N_5204,N_5076,N_5179);
or U5205 (N_5205,N_5180,N_5048);
nand U5206 (N_5206,N_5178,N_5099);
and U5207 (N_5207,N_5189,N_5187);
and U5208 (N_5208,N_5085,N_5197);
or U5209 (N_5209,N_5101,N_5047);
xnor U5210 (N_5210,N_5164,N_5031);
or U5211 (N_5211,N_5064,N_5091);
or U5212 (N_5212,N_5058,N_5062);
or U5213 (N_5213,N_5007,N_5116);
or U5214 (N_5214,N_5089,N_5098);
nor U5215 (N_5215,N_5102,N_5004);
and U5216 (N_5216,N_5111,N_5185);
nand U5217 (N_5217,N_5000,N_5186);
nand U5218 (N_5218,N_5115,N_5174);
nor U5219 (N_5219,N_5013,N_5108);
nor U5220 (N_5220,N_5077,N_5083);
nor U5221 (N_5221,N_5049,N_5139);
and U5222 (N_5222,N_5029,N_5191);
nor U5223 (N_5223,N_5154,N_5135);
nand U5224 (N_5224,N_5039,N_5005);
nand U5225 (N_5225,N_5021,N_5069);
nor U5226 (N_5226,N_5086,N_5024);
xor U5227 (N_5227,N_5141,N_5173);
nand U5228 (N_5228,N_5168,N_5018);
nand U5229 (N_5229,N_5149,N_5159);
or U5230 (N_5230,N_5063,N_5095);
or U5231 (N_5231,N_5026,N_5080);
and U5232 (N_5232,N_5146,N_5056);
or U5233 (N_5233,N_5041,N_5150);
nand U5234 (N_5234,N_5096,N_5106);
and U5235 (N_5235,N_5120,N_5156);
and U5236 (N_5236,N_5194,N_5015);
and U5237 (N_5237,N_5019,N_5025);
and U5238 (N_5238,N_5052,N_5012);
and U5239 (N_5239,N_5022,N_5045);
or U5240 (N_5240,N_5044,N_5046);
or U5241 (N_5241,N_5118,N_5145);
and U5242 (N_5242,N_5157,N_5059);
and U5243 (N_5243,N_5142,N_5132);
xnor U5244 (N_5244,N_5001,N_5067);
nor U5245 (N_5245,N_5065,N_5014);
nor U5246 (N_5246,N_5009,N_5107);
or U5247 (N_5247,N_5136,N_5158);
nand U5248 (N_5248,N_5100,N_5032);
nor U5249 (N_5249,N_5081,N_5036);
nand U5250 (N_5250,N_5193,N_5094);
nand U5251 (N_5251,N_5105,N_5104);
nand U5252 (N_5252,N_5103,N_5020);
nand U5253 (N_5253,N_5175,N_5079);
xnor U5254 (N_5254,N_5050,N_5190);
and U5255 (N_5255,N_5117,N_5030);
xor U5256 (N_5256,N_5184,N_5182);
nand U5257 (N_5257,N_5196,N_5043);
nor U5258 (N_5258,N_5016,N_5053);
nor U5259 (N_5259,N_5163,N_5148);
and U5260 (N_5260,N_5131,N_5133);
and U5261 (N_5261,N_5124,N_5055);
and U5262 (N_5262,N_5084,N_5040);
nand U5263 (N_5263,N_5090,N_5119);
or U5264 (N_5264,N_5181,N_5171);
xor U5265 (N_5265,N_5075,N_5147);
and U5266 (N_5266,N_5008,N_5088);
or U5267 (N_5267,N_5054,N_5137);
xnor U5268 (N_5268,N_5097,N_5114);
or U5269 (N_5269,N_5144,N_5122);
nand U5270 (N_5270,N_5134,N_5129);
xnor U5271 (N_5271,N_5035,N_5176);
or U5272 (N_5272,N_5130,N_5123);
nor U5273 (N_5273,N_5006,N_5121);
nand U5274 (N_5274,N_5003,N_5172);
or U5275 (N_5275,N_5010,N_5198);
xnor U5276 (N_5276,N_5112,N_5093);
and U5277 (N_5277,N_5143,N_5042);
nor U5278 (N_5278,N_5152,N_5127);
and U5279 (N_5279,N_5162,N_5017);
or U5280 (N_5280,N_5165,N_5074);
nand U5281 (N_5281,N_5188,N_5061);
nor U5282 (N_5282,N_5169,N_5151);
and U5283 (N_5283,N_5070,N_5192);
xnor U5284 (N_5284,N_5140,N_5060);
xnor U5285 (N_5285,N_5155,N_5027);
or U5286 (N_5286,N_5011,N_5161);
xor U5287 (N_5287,N_5034,N_5183);
xnor U5288 (N_5288,N_5128,N_5160);
nand U5289 (N_5289,N_5125,N_5023);
and U5290 (N_5290,N_5199,N_5028);
or U5291 (N_5291,N_5082,N_5072);
nor U5292 (N_5292,N_5109,N_5038);
nor U5293 (N_5293,N_5166,N_5113);
xnor U5294 (N_5294,N_5037,N_5066);
or U5295 (N_5295,N_5051,N_5195);
or U5296 (N_5296,N_5153,N_5092);
or U5297 (N_5297,N_5138,N_5170);
nor U5298 (N_5298,N_5071,N_5177);
nor U5299 (N_5299,N_5002,N_5033);
and U5300 (N_5300,N_5177,N_5087);
and U5301 (N_5301,N_5185,N_5131);
nand U5302 (N_5302,N_5004,N_5075);
or U5303 (N_5303,N_5058,N_5007);
nor U5304 (N_5304,N_5121,N_5104);
xor U5305 (N_5305,N_5021,N_5067);
or U5306 (N_5306,N_5135,N_5095);
nand U5307 (N_5307,N_5099,N_5069);
nor U5308 (N_5308,N_5008,N_5109);
nand U5309 (N_5309,N_5056,N_5061);
xor U5310 (N_5310,N_5012,N_5140);
and U5311 (N_5311,N_5166,N_5158);
or U5312 (N_5312,N_5057,N_5193);
nor U5313 (N_5313,N_5199,N_5184);
nor U5314 (N_5314,N_5014,N_5085);
nand U5315 (N_5315,N_5068,N_5122);
nand U5316 (N_5316,N_5171,N_5082);
nor U5317 (N_5317,N_5149,N_5111);
nand U5318 (N_5318,N_5124,N_5135);
nor U5319 (N_5319,N_5112,N_5012);
xnor U5320 (N_5320,N_5014,N_5182);
nor U5321 (N_5321,N_5014,N_5064);
nor U5322 (N_5322,N_5080,N_5040);
xor U5323 (N_5323,N_5006,N_5074);
nor U5324 (N_5324,N_5003,N_5101);
or U5325 (N_5325,N_5027,N_5173);
nand U5326 (N_5326,N_5013,N_5133);
nor U5327 (N_5327,N_5125,N_5129);
nor U5328 (N_5328,N_5064,N_5126);
nor U5329 (N_5329,N_5039,N_5127);
or U5330 (N_5330,N_5071,N_5111);
nor U5331 (N_5331,N_5018,N_5010);
nand U5332 (N_5332,N_5032,N_5166);
and U5333 (N_5333,N_5069,N_5001);
nand U5334 (N_5334,N_5188,N_5004);
and U5335 (N_5335,N_5081,N_5026);
nor U5336 (N_5336,N_5137,N_5040);
xor U5337 (N_5337,N_5141,N_5111);
and U5338 (N_5338,N_5100,N_5081);
or U5339 (N_5339,N_5044,N_5196);
or U5340 (N_5340,N_5105,N_5040);
and U5341 (N_5341,N_5108,N_5165);
nand U5342 (N_5342,N_5113,N_5163);
xor U5343 (N_5343,N_5098,N_5109);
nor U5344 (N_5344,N_5177,N_5080);
nor U5345 (N_5345,N_5053,N_5095);
xor U5346 (N_5346,N_5057,N_5052);
nor U5347 (N_5347,N_5023,N_5028);
nor U5348 (N_5348,N_5071,N_5042);
nand U5349 (N_5349,N_5172,N_5178);
nor U5350 (N_5350,N_5017,N_5174);
or U5351 (N_5351,N_5075,N_5196);
nor U5352 (N_5352,N_5192,N_5123);
and U5353 (N_5353,N_5004,N_5115);
and U5354 (N_5354,N_5176,N_5106);
or U5355 (N_5355,N_5187,N_5182);
nor U5356 (N_5356,N_5020,N_5128);
nand U5357 (N_5357,N_5130,N_5006);
nand U5358 (N_5358,N_5124,N_5005);
or U5359 (N_5359,N_5010,N_5058);
or U5360 (N_5360,N_5170,N_5021);
or U5361 (N_5361,N_5027,N_5154);
or U5362 (N_5362,N_5141,N_5013);
and U5363 (N_5363,N_5086,N_5017);
nand U5364 (N_5364,N_5191,N_5084);
nand U5365 (N_5365,N_5096,N_5152);
and U5366 (N_5366,N_5162,N_5075);
and U5367 (N_5367,N_5173,N_5117);
or U5368 (N_5368,N_5155,N_5072);
and U5369 (N_5369,N_5167,N_5034);
or U5370 (N_5370,N_5009,N_5072);
nor U5371 (N_5371,N_5149,N_5166);
nor U5372 (N_5372,N_5122,N_5049);
nand U5373 (N_5373,N_5084,N_5043);
and U5374 (N_5374,N_5034,N_5069);
and U5375 (N_5375,N_5187,N_5115);
and U5376 (N_5376,N_5068,N_5022);
nor U5377 (N_5377,N_5130,N_5190);
nor U5378 (N_5378,N_5197,N_5163);
or U5379 (N_5379,N_5091,N_5175);
and U5380 (N_5380,N_5106,N_5019);
and U5381 (N_5381,N_5104,N_5160);
or U5382 (N_5382,N_5194,N_5126);
or U5383 (N_5383,N_5188,N_5003);
or U5384 (N_5384,N_5088,N_5154);
nand U5385 (N_5385,N_5004,N_5153);
nand U5386 (N_5386,N_5173,N_5120);
and U5387 (N_5387,N_5190,N_5177);
and U5388 (N_5388,N_5099,N_5090);
nor U5389 (N_5389,N_5162,N_5168);
or U5390 (N_5390,N_5033,N_5069);
nand U5391 (N_5391,N_5111,N_5115);
and U5392 (N_5392,N_5024,N_5054);
nand U5393 (N_5393,N_5021,N_5026);
and U5394 (N_5394,N_5134,N_5067);
and U5395 (N_5395,N_5050,N_5137);
xnor U5396 (N_5396,N_5082,N_5056);
and U5397 (N_5397,N_5135,N_5110);
and U5398 (N_5398,N_5152,N_5141);
or U5399 (N_5399,N_5095,N_5103);
or U5400 (N_5400,N_5319,N_5230);
nor U5401 (N_5401,N_5292,N_5275);
nand U5402 (N_5402,N_5360,N_5308);
nand U5403 (N_5403,N_5260,N_5239);
and U5404 (N_5404,N_5256,N_5333);
and U5405 (N_5405,N_5370,N_5313);
or U5406 (N_5406,N_5394,N_5281);
or U5407 (N_5407,N_5271,N_5200);
nand U5408 (N_5408,N_5215,N_5395);
nand U5409 (N_5409,N_5302,N_5216);
nand U5410 (N_5410,N_5280,N_5342);
nor U5411 (N_5411,N_5225,N_5357);
or U5412 (N_5412,N_5262,N_5205);
nand U5413 (N_5413,N_5315,N_5380);
nand U5414 (N_5414,N_5329,N_5284);
or U5415 (N_5415,N_5353,N_5392);
and U5416 (N_5416,N_5373,N_5364);
or U5417 (N_5417,N_5252,N_5237);
nand U5418 (N_5418,N_5270,N_5391);
nand U5419 (N_5419,N_5258,N_5274);
or U5420 (N_5420,N_5249,N_5204);
or U5421 (N_5421,N_5365,N_5310);
nand U5422 (N_5422,N_5322,N_5299);
nor U5423 (N_5423,N_5378,N_5396);
nor U5424 (N_5424,N_5320,N_5351);
and U5425 (N_5425,N_5289,N_5301);
xnor U5426 (N_5426,N_5255,N_5387);
or U5427 (N_5427,N_5377,N_5375);
or U5428 (N_5428,N_5263,N_5221);
nor U5429 (N_5429,N_5226,N_5334);
xnor U5430 (N_5430,N_5296,N_5264);
nand U5431 (N_5431,N_5210,N_5367);
nor U5432 (N_5432,N_5203,N_5276);
or U5433 (N_5433,N_5350,N_5343);
nor U5434 (N_5434,N_5248,N_5337);
nand U5435 (N_5435,N_5345,N_5362);
or U5436 (N_5436,N_5311,N_5304);
nor U5437 (N_5437,N_5206,N_5366);
nand U5438 (N_5438,N_5385,N_5207);
nand U5439 (N_5439,N_5356,N_5389);
and U5440 (N_5440,N_5219,N_5303);
nand U5441 (N_5441,N_5243,N_5352);
nand U5442 (N_5442,N_5228,N_5214);
and U5443 (N_5443,N_5209,N_5268);
or U5444 (N_5444,N_5327,N_5306);
nand U5445 (N_5445,N_5349,N_5233);
nand U5446 (N_5446,N_5305,N_5359);
nand U5447 (N_5447,N_5282,N_5363);
and U5448 (N_5448,N_5323,N_5287);
nand U5449 (N_5449,N_5384,N_5261);
and U5450 (N_5450,N_5348,N_5266);
nand U5451 (N_5451,N_5201,N_5232);
and U5452 (N_5452,N_5321,N_5312);
and U5453 (N_5453,N_5398,N_5393);
nand U5454 (N_5454,N_5202,N_5355);
nor U5455 (N_5455,N_5347,N_5265);
and U5456 (N_5456,N_5257,N_5240);
or U5457 (N_5457,N_5212,N_5376);
and U5458 (N_5458,N_5235,N_5211);
xnor U5459 (N_5459,N_5244,N_5332);
nand U5460 (N_5460,N_5316,N_5241);
and U5461 (N_5461,N_5390,N_5330);
nand U5462 (N_5462,N_5379,N_5217);
xor U5463 (N_5463,N_5277,N_5336);
nor U5464 (N_5464,N_5234,N_5317);
nand U5465 (N_5465,N_5383,N_5227);
and U5466 (N_5466,N_5223,N_5229);
nand U5467 (N_5467,N_5288,N_5245);
nor U5468 (N_5468,N_5208,N_5369);
nand U5469 (N_5469,N_5259,N_5285);
nor U5470 (N_5470,N_5279,N_5326);
and U5471 (N_5471,N_5374,N_5382);
nand U5472 (N_5472,N_5290,N_5269);
and U5473 (N_5473,N_5251,N_5338);
xor U5474 (N_5474,N_5246,N_5340);
xnor U5475 (N_5475,N_5309,N_5335);
nand U5476 (N_5476,N_5253,N_5236);
nor U5477 (N_5477,N_5222,N_5298);
nand U5478 (N_5478,N_5224,N_5283);
xor U5479 (N_5479,N_5297,N_5361);
nand U5480 (N_5480,N_5368,N_5254);
or U5481 (N_5481,N_5346,N_5354);
nor U5482 (N_5482,N_5328,N_5386);
and U5483 (N_5483,N_5293,N_5358);
or U5484 (N_5484,N_5218,N_5286);
or U5485 (N_5485,N_5294,N_5381);
or U5486 (N_5486,N_5307,N_5278);
nand U5487 (N_5487,N_5291,N_5267);
and U5488 (N_5488,N_5250,N_5238);
xor U5489 (N_5489,N_5331,N_5231);
nor U5490 (N_5490,N_5339,N_5388);
and U5491 (N_5491,N_5371,N_5399);
nor U5492 (N_5492,N_5220,N_5344);
nor U5493 (N_5493,N_5314,N_5213);
nand U5494 (N_5494,N_5300,N_5272);
nand U5495 (N_5495,N_5397,N_5318);
and U5496 (N_5496,N_5295,N_5372);
or U5497 (N_5497,N_5325,N_5247);
or U5498 (N_5498,N_5341,N_5324);
nand U5499 (N_5499,N_5273,N_5242);
or U5500 (N_5500,N_5359,N_5399);
nor U5501 (N_5501,N_5235,N_5363);
nor U5502 (N_5502,N_5268,N_5337);
and U5503 (N_5503,N_5226,N_5295);
and U5504 (N_5504,N_5356,N_5232);
nor U5505 (N_5505,N_5251,N_5345);
nand U5506 (N_5506,N_5330,N_5398);
nand U5507 (N_5507,N_5323,N_5237);
and U5508 (N_5508,N_5284,N_5328);
nand U5509 (N_5509,N_5310,N_5213);
or U5510 (N_5510,N_5343,N_5373);
or U5511 (N_5511,N_5338,N_5302);
or U5512 (N_5512,N_5332,N_5279);
and U5513 (N_5513,N_5317,N_5332);
xor U5514 (N_5514,N_5244,N_5297);
or U5515 (N_5515,N_5306,N_5224);
nor U5516 (N_5516,N_5348,N_5295);
nand U5517 (N_5517,N_5341,N_5289);
nand U5518 (N_5518,N_5360,N_5246);
and U5519 (N_5519,N_5240,N_5238);
or U5520 (N_5520,N_5275,N_5333);
or U5521 (N_5521,N_5281,N_5302);
or U5522 (N_5522,N_5387,N_5299);
nor U5523 (N_5523,N_5398,N_5252);
nor U5524 (N_5524,N_5332,N_5395);
nor U5525 (N_5525,N_5240,N_5227);
or U5526 (N_5526,N_5366,N_5239);
or U5527 (N_5527,N_5305,N_5337);
nor U5528 (N_5528,N_5315,N_5220);
nor U5529 (N_5529,N_5267,N_5233);
xor U5530 (N_5530,N_5271,N_5388);
nor U5531 (N_5531,N_5350,N_5214);
nor U5532 (N_5532,N_5299,N_5392);
or U5533 (N_5533,N_5366,N_5270);
nor U5534 (N_5534,N_5393,N_5214);
or U5535 (N_5535,N_5298,N_5257);
nor U5536 (N_5536,N_5276,N_5388);
and U5537 (N_5537,N_5345,N_5356);
nor U5538 (N_5538,N_5278,N_5271);
nand U5539 (N_5539,N_5275,N_5318);
xor U5540 (N_5540,N_5297,N_5299);
nand U5541 (N_5541,N_5279,N_5384);
or U5542 (N_5542,N_5237,N_5368);
nand U5543 (N_5543,N_5391,N_5339);
and U5544 (N_5544,N_5252,N_5395);
nand U5545 (N_5545,N_5261,N_5274);
nor U5546 (N_5546,N_5335,N_5200);
xor U5547 (N_5547,N_5267,N_5343);
or U5548 (N_5548,N_5349,N_5229);
xnor U5549 (N_5549,N_5343,N_5317);
and U5550 (N_5550,N_5366,N_5308);
nand U5551 (N_5551,N_5240,N_5273);
nand U5552 (N_5552,N_5330,N_5238);
and U5553 (N_5553,N_5379,N_5352);
and U5554 (N_5554,N_5204,N_5340);
and U5555 (N_5555,N_5221,N_5335);
xor U5556 (N_5556,N_5323,N_5341);
nand U5557 (N_5557,N_5315,N_5346);
nor U5558 (N_5558,N_5371,N_5260);
or U5559 (N_5559,N_5232,N_5273);
or U5560 (N_5560,N_5291,N_5349);
or U5561 (N_5561,N_5229,N_5248);
and U5562 (N_5562,N_5287,N_5317);
or U5563 (N_5563,N_5294,N_5217);
and U5564 (N_5564,N_5357,N_5262);
and U5565 (N_5565,N_5213,N_5267);
nor U5566 (N_5566,N_5233,N_5324);
xor U5567 (N_5567,N_5311,N_5309);
and U5568 (N_5568,N_5346,N_5202);
and U5569 (N_5569,N_5287,N_5340);
or U5570 (N_5570,N_5257,N_5317);
nand U5571 (N_5571,N_5392,N_5301);
or U5572 (N_5572,N_5340,N_5276);
nor U5573 (N_5573,N_5331,N_5368);
nand U5574 (N_5574,N_5344,N_5213);
and U5575 (N_5575,N_5278,N_5378);
xnor U5576 (N_5576,N_5328,N_5334);
or U5577 (N_5577,N_5229,N_5247);
nor U5578 (N_5578,N_5275,N_5315);
nor U5579 (N_5579,N_5365,N_5320);
nor U5580 (N_5580,N_5219,N_5245);
or U5581 (N_5581,N_5246,N_5366);
or U5582 (N_5582,N_5251,N_5296);
nor U5583 (N_5583,N_5396,N_5363);
or U5584 (N_5584,N_5211,N_5273);
nor U5585 (N_5585,N_5229,N_5285);
nand U5586 (N_5586,N_5219,N_5226);
and U5587 (N_5587,N_5315,N_5334);
or U5588 (N_5588,N_5287,N_5212);
nor U5589 (N_5589,N_5327,N_5271);
and U5590 (N_5590,N_5234,N_5328);
nor U5591 (N_5591,N_5274,N_5260);
nor U5592 (N_5592,N_5381,N_5237);
xnor U5593 (N_5593,N_5209,N_5321);
or U5594 (N_5594,N_5341,N_5388);
nand U5595 (N_5595,N_5201,N_5217);
nor U5596 (N_5596,N_5365,N_5319);
and U5597 (N_5597,N_5375,N_5245);
nand U5598 (N_5598,N_5273,N_5205);
nand U5599 (N_5599,N_5303,N_5245);
nor U5600 (N_5600,N_5553,N_5499);
xor U5601 (N_5601,N_5425,N_5593);
and U5602 (N_5602,N_5554,N_5573);
or U5603 (N_5603,N_5580,N_5509);
and U5604 (N_5604,N_5511,N_5482);
nor U5605 (N_5605,N_5403,N_5417);
nor U5606 (N_5606,N_5419,N_5485);
or U5607 (N_5607,N_5585,N_5451);
nor U5608 (N_5608,N_5592,N_5457);
and U5609 (N_5609,N_5504,N_5527);
and U5610 (N_5610,N_5575,N_5543);
and U5611 (N_5611,N_5443,N_5507);
xor U5612 (N_5612,N_5413,N_5455);
xnor U5613 (N_5613,N_5587,N_5448);
nand U5614 (N_5614,N_5586,N_5437);
or U5615 (N_5615,N_5537,N_5547);
or U5616 (N_5616,N_5441,N_5463);
nand U5617 (N_5617,N_5564,N_5572);
nand U5618 (N_5618,N_5472,N_5541);
and U5619 (N_5619,N_5576,N_5544);
xnor U5620 (N_5620,N_5439,N_5461);
nand U5621 (N_5621,N_5508,N_5502);
or U5622 (N_5622,N_5578,N_5510);
nor U5623 (N_5623,N_5589,N_5440);
xnor U5624 (N_5624,N_5583,N_5428);
and U5625 (N_5625,N_5435,N_5549);
and U5626 (N_5626,N_5567,N_5471);
and U5627 (N_5627,N_5584,N_5429);
nor U5628 (N_5628,N_5422,N_5582);
or U5629 (N_5629,N_5453,N_5473);
nor U5630 (N_5630,N_5409,N_5464);
nand U5631 (N_5631,N_5469,N_5591);
nor U5632 (N_5632,N_5563,N_5513);
or U5633 (N_5633,N_5515,N_5460);
nor U5634 (N_5634,N_5481,N_5491);
nor U5635 (N_5635,N_5478,N_5528);
nor U5636 (N_5636,N_5494,N_5495);
nor U5637 (N_5637,N_5526,N_5447);
nor U5638 (N_5638,N_5488,N_5438);
nand U5639 (N_5639,N_5444,N_5529);
and U5640 (N_5640,N_5411,N_5432);
and U5641 (N_5641,N_5574,N_5466);
xnor U5642 (N_5642,N_5407,N_5487);
nor U5643 (N_5643,N_5459,N_5493);
nor U5644 (N_5644,N_5594,N_5420);
xnor U5645 (N_5645,N_5512,N_5421);
nor U5646 (N_5646,N_5501,N_5599);
and U5647 (N_5647,N_5490,N_5570);
nand U5648 (N_5648,N_5545,N_5500);
nor U5649 (N_5649,N_5579,N_5531);
or U5650 (N_5650,N_5568,N_5416);
nand U5651 (N_5651,N_5533,N_5524);
nand U5652 (N_5652,N_5497,N_5449);
nand U5653 (N_5653,N_5534,N_5402);
or U5654 (N_5654,N_5536,N_5598);
and U5655 (N_5655,N_5503,N_5535);
or U5656 (N_5656,N_5548,N_5517);
nor U5657 (N_5657,N_5551,N_5514);
nor U5658 (N_5658,N_5454,N_5446);
xor U5659 (N_5659,N_5569,N_5577);
nor U5660 (N_5660,N_5418,N_5516);
and U5661 (N_5661,N_5566,N_5562);
nor U5662 (N_5662,N_5597,N_5525);
and U5663 (N_5663,N_5571,N_5559);
nand U5664 (N_5664,N_5410,N_5476);
xnor U5665 (N_5665,N_5550,N_5458);
and U5666 (N_5666,N_5445,N_5484);
nor U5667 (N_5667,N_5467,N_5404);
nor U5668 (N_5668,N_5530,N_5452);
nand U5669 (N_5669,N_5412,N_5492);
and U5670 (N_5670,N_5468,N_5431);
xnor U5671 (N_5671,N_5498,N_5496);
and U5672 (N_5672,N_5540,N_5520);
or U5673 (N_5673,N_5479,N_5427);
nand U5674 (N_5674,N_5474,N_5522);
and U5675 (N_5675,N_5434,N_5521);
or U5676 (N_5676,N_5433,N_5539);
nor U5677 (N_5677,N_5442,N_5561);
xnor U5678 (N_5678,N_5552,N_5546);
and U5679 (N_5679,N_5462,N_5558);
nor U5680 (N_5680,N_5465,N_5406);
and U5681 (N_5681,N_5555,N_5557);
xnor U5682 (N_5682,N_5408,N_5523);
xor U5683 (N_5683,N_5532,N_5414);
xnor U5684 (N_5684,N_5519,N_5542);
and U5685 (N_5685,N_5565,N_5486);
nand U5686 (N_5686,N_5430,N_5506);
nor U5687 (N_5687,N_5475,N_5518);
nor U5688 (N_5688,N_5596,N_5400);
xor U5689 (N_5689,N_5560,N_5556);
or U5690 (N_5690,N_5450,N_5436);
or U5691 (N_5691,N_5456,N_5426);
and U5692 (N_5692,N_5538,N_5581);
and U5693 (N_5693,N_5595,N_5424);
nor U5694 (N_5694,N_5480,N_5470);
xor U5695 (N_5695,N_5477,N_5483);
nand U5696 (N_5696,N_5415,N_5401);
xnor U5697 (N_5697,N_5423,N_5505);
nand U5698 (N_5698,N_5590,N_5588);
and U5699 (N_5699,N_5489,N_5405);
nor U5700 (N_5700,N_5557,N_5416);
or U5701 (N_5701,N_5553,N_5504);
and U5702 (N_5702,N_5579,N_5416);
and U5703 (N_5703,N_5435,N_5532);
nor U5704 (N_5704,N_5582,N_5431);
or U5705 (N_5705,N_5489,N_5420);
nand U5706 (N_5706,N_5529,N_5472);
nor U5707 (N_5707,N_5454,N_5457);
or U5708 (N_5708,N_5572,N_5520);
and U5709 (N_5709,N_5443,N_5450);
and U5710 (N_5710,N_5555,N_5564);
xor U5711 (N_5711,N_5483,N_5402);
nor U5712 (N_5712,N_5571,N_5409);
or U5713 (N_5713,N_5430,N_5579);
nor U5714 (N_5714,N_5515,N_5558);
nor U5715 (N_5715,N_5513,N_5573);
nand U5716 (N_5716,N_5410,N_5479);
and U5717 (N_5717,N_5407,N_5494);
and U5718 (N_5718,N_5556,N_5432);
nand U5719 (N_5719,N_5498,N_5539);
nor U5720 (N_5720,N_5538,N_5447);
nand U5721 (N_5721,N_5582,N_5475);
nor U5722 (N_5722,N_5406,N_5476);
xnor U5723 (N_5723,N_5588,N_5580);
or U5724 (N_5724,N_5547,N_5594);
xor U5725 (N_5725,N_5549,N_5505);
or U5726 (N_5726,N_5523,N_5576);
nor U5727 (N_5727,N_5558,N_5586);
and U5728 (N_5728,N_5491,N_5476);
nor U5729 (N_5729,N_5456,N_5507);
xnor U5730 (N_5730,N_5526,N_5430);
nand U5731 (N_5731,N_5530,N_5512);
nor U5732 (N_5732,N_5589,N_5419);
nor U5733 (N_5733,N_5420,N_5555);
or U5734 (N_5734,N_5550,N_5553);
nand U5735 (N_5735,N_5401,N_5516);
xnor U5736 (N_5736,N_5513,N_5429);
xnor U5737 (N_5737,N_5491,N_5587);
or U5738 (N_5738,N_5417,N_5535);
nor U5739 (N_5739,N_5458,N_5488);
or U5740 (N_5740,N_5504,N_5510);
and U5741 (N_5741,N_5412,N_5529);
nand U5742 (N_5742,N_5529,N_5409);
nand U5743 (N_5743,N_5592,N_5577);
or U5744 (N_5744,N_5545,N_5421);
nor U5745 (N_5745,N_5517,N_5542);
nand U5746 (N_5746,N_5455,N_5545);
and U5747 (N_5747,N_5539,N_5439);
nor U5748 (N_5748,N_5491,N_5487);
nand U5749 (N_5749,N_5575,N_5456);
or U5750 (N_5750,N_5500,N_5556);
nand U5751 (N_5751,N_5456,N_5522);
and U5752 (N_5752,N_5457,N_5422);
nor U5753 (N_5753,N_5520,N_5522);
or U5754 (N_5754,N_5519,N_5413);
or U5755 (N_5755,N_5572,N_5547);
xnor U5756 (N_5756,N_5564,N_5561);
or U5757 (N_5757,N_5590,N_5416);
nand U5758 (N_5758,N_5592,N_5522);
nor U5759 (N_5759,N_5462,N_5518);
nor U5760 (N_5760,N_5525,N_5453);
or U5761 (N_5761,N_5461,N_5422);
nor U5762 (N_5762,N_5544,N_5552);
nand U5763 (N_5763,N_5483,N_5478);
or U5764 (N_5764,N_5433,N_5459);
or U5765 (N_5765,N_5571,N_5557);
or U5766 (N_5766,N_5462,N_5493);
or U5767 (N_5767,N_5532,N_5596);
and U5768 (N_5768,N_5461,N_5591);
xnor U5769 (N_5769,N_5521,N_5535);
xnor U5770 (N_5770,N_5538,N_5481);
nand U5771 (N_5771,N_5512,N_5407);
or U5772 (N_5772,N_5530,N_5565);
nor U5773 (N_5773,N_5411,N_5419);
or U5774 (N_5774,N_5452,N_5524);
nor U5775 (N_5775,N_5508,N_5466);
or U5776 (N_5776,N_5586,N_5515);
and U5777 (N_5777,N_5522,N_5572);
xor U5778 (N_5778,N_5452,N_5545);
xor U5779 (N_5779,N_5425,N_5456);
and U5780 (N_5780,N_5547,N_5552);
or U5781 (N_5781,N_5415,N_5597);
nand U5782 (N_5782,N_5539,N_5592);
or U5783 (N_5783,N_5544,N_5538);
nand U5784 (N_5784,N_5575,N_5401);
nor U5785 (N_5785,N_5458,N_5554);
or U5786 (N_5786,N_5579,N_5406);
or U5787 (N_5787,N_5497,N_5585);
nor U5788 (N_5788,N_5465,N_5501);
nand U5789 (N_5789,N_5580,N_5455);
nand U5790 (N_5790,N_5575,N_5595);
nor U5791 (N_5791,N_5486,N_5583);
nor U5792 (N_5792,N_5404,N_5537);
nor U5793 (N_5793,N_5400,N_5521);
xnor U5794 (N_5794,N_5571,N_5593);
nand U5795 (N_5795,N_5424,N_5563);
nor U5796 (N_5796,N_5445,N_5566);
or U5797 (N_5797,N_5451,N_5540);
and U5798 (N_5798,N_5524,N_5428);
and U5799 (N_5799,N_5439,N_5598);
xnor U5800 (N_5800,N_5636,N_5745);
nor U5801 (N_5801,N_5784,N_5642);
nand U5802 (N_5802,N_5600,N_5798);
or U5803 (N_5803,N_5631,N_5726);
nor U5804 (N_5804,N_5678,N_5752);
and U5805 (N_5805,N_5766,N_5786);
nand U5806 (N_5806,N_5604,N_5630);
nor U5807 (N_5807,N_5747,N_5684);
or U5808 (N_5808,N_5666,N_5613);
or U5809 (N_5809,N_5754,N_5669);
or U5810 (N_5810,N_5612,N_5789);
and U5811 (N_5811,N_5740,N_5717);
nand U5812 (N_5812,N_5788,N_5693);
nand U5813 (N_5813,N_5782,N_5775);
nor U5814 (N_5814,N_5688,N_5616);
and U5815 (N_5815,N_5773,N_5731);
nand U5816 (N_5816,N_5709,N_5750);
or U5817 (N_5817,N_5771,N_5695);
nor U5818 (N_5818,N_5626,N_5647);
or U5819 (N_5819,N_5755,N_5792);
or U5820 (N_5820,N_5710,N_5664);
and U5821 (N_5821,N_5627,N_5632);
nand U5822 (N_5822,N_5760,N_5690);
nand U5823 (N_5823,N_5624,N_5718);
or U5824 (N_5824,N_5661,N_5743);
xor U5825 (N_5825,N_5772,N_5790);
nor U5826 (N_5826,N_5674,N_5637);
and U5827 (N_5827,N_5656,N_5737);
or U5828 (N_5828,N_5719,N_5796);
nand U5829 (N_5829,N_5757,N_5645);
or U5830 (N_5830,N_5708,N_5702);
or U5831 (N_5831,N_5759,N_5667);
nor U5832 (N_5832,N_5668,N_5623);
or U5833 (N_5833,N_5749,N_5651);
nand U5834 (N_5834,N_5653,N_5783);
and U5835 (N_5835,N_5714,N_5671);
and U5836 (N_5836,N_5694,N_5751);
nor U5837 (N_5837,N_5780,N_5795);
or U5838 (N_5838,N_5625,N_5761);
or U5839 (N_5839,N_5662,N_5748);
nand U5840 (N_5840,N_5744,N_5776);
nor U5841 (N_5841,N_5727,N_5781);
and U5842 (N_5842,N_5793,N_5629);
nand U5843 (N_5843,N_5706,N_5730);
or U5844 (N_5844,N_5712,N_5652);
nor U5845 (N_5845,N_5621,N_5701);
and U5846 (N_5846,N_5725,N_5777);
and U5847 (N_5847,N_5670,N_5638);
or U5848 (N_5848,N_5665,N_5654);
and U5849 (N_5849,N_5763,N_5724);
and U5850 (N_5850,N_5635,N_5742);
and U5851 (N_5851,N_5650,N_5680);
or U5852 (N_5852,N_5799,N_5633);
and U5853 (N_5853,N_5681,N_5686);
nor U5854 (N_5854,N_5648,N_5735);
nor U5855 (N_5855,N_5617,N_5704);
and U5856 (N_5856,N_5663,N_5779);
xnor U5857 (N_5857,N_5672,N_5729);
or U5858 (N_5858,N_5608,N_5736);
and U5859 (N_5859,N_5762,N_5689);
and U5860 (N_5860,N_5699,N_5649);
nor U5861 (N_5861,N_5640,N_5646);
nor U5862 (N_5862,N_5739,N_5728);
nand U5863 (N_5863,N_5687,N_5696);
or U5864 (N_5864,N_5764,N_5676);
and U5865 (N_5865,N_5733,N_5715);
nand U5866 (N_5866,N_5673,N_5615);
and U5867 (N_5867,N_5614,N_5643);
nor U5868 (N_5868,N_5794,N_5606);
nand U5869 (N_5869,N_5660,N_5628);
xor U5870 (N_5870,N_5607,N_5787);
and U5871 (N_5871,N_5720,N_5698);
and U5872 (N_5872,N_5738,N_5723);
and U5873 (N_5873,N_5703,N_5716);
or U5874 (N_5874,N_5655,N_5721);
or U5875 (N_5875,N_5770,N_5697);
xor U5876 (N_5876,N_5765,N_5679);
xnor U5877 (N_5877,N_5611,N_5618);
nand U5878 (N_5878,N_5746,N_5641);
and U5879 (N_5879,N_5700,N_5610);
and U5880 (N_5880,N_5603,N_5644);
nor U5881 (N_5881,N_5683,N_5797);
nand U5882 (N_5882,N_5774,N_5734);
or U5883 (N_5883,N_5601,N_5741);
xnor U5884 (N_5884,N_5685,N_5657);
xor U5885 (N_5885,N_5692,N_5620);
or U5886 (N_5886,N_5659,N_5619);
and U5887 (N_5887,N_5622,N_5707);
and U5888 (N_5888,N_5758,N_5682);
nor U5889 (N_5889,N_5677,N_5711);
xor U5890 (N_5890,N_5767,N_5691);
xor U5891 (N_5891,N_5768,N_5753);
xnor U5892 (N_5892,N_5639,N_5722);
xnor U5893 (N_5893,N_5791,N_5634);
xnor U5894 (N_5894,N_5732,N_5609);
nand U5895 (N_5895,N_5602,N_5785);
xnor U5896 (N_5896,N_5658,N_5756);
or U5897 (N_5897,N_5605,N_5778);
and U5898 (N_5898,N_5675,N_5705);
xnor U5899 (N_5899,N_5713,N_5769);
and U5900 (N_5900,N_5780,N_5652);
or U5901 (N_5901,N_5723,N_5700);
or U5902 (N_5902,N_5609,N_5649);
nor U5903 (N_5903,N_5682,N_5799);
xor U5904 (N_5904,N_5708,N_5690);
and U5905 (N_5905,N_5774,N_5716);
nor U5906 (N_5906,N_5760,N_5769);
and U5907 (N_5907,N_5717,N_5730);
or U5908 (N_5908,N_5613,N_5660);
nor U5909 (N_5909,N_5781,N_5676);
or U5910 (N_5910,N_5775,N_5627);
nor U5911 (N_5911,N_5658,N_5785);
or U5912 (N_5912,N_5686,N_5778);
and U5913 (N_5913,N_5636,N_5761);
nand U5914 (N_5914,N_5750,N_5668);
nor U5915 (N_5915,N_5638,N_5702);
and U5916 (N_5916,N_5790,N_5765);
and U5917 (N_5917,N_5731,N_5799);
and U5918 (N_5918,N_5722,N_5760);
nor U5919 (N_5919,N_5651,N_5767);
nand U5920 (N_5920,N_5680,N_5701);
and U5921 (N_5921,N_5617,N_5655);
nand U5922 (N_5922,N_5630,N_5647);
xnor U5923 (N_5923,N_5721,N_5645);
or U5924 (N_5924,N_5721,N_5751);
and U5925 (N_5925,N_5776,N_5658);
or U5926 (N_5926,N_5654,N_5660);
or U5927 (N_5927,N_5667,N_5710);
and U5928 (N_5928,N_5739,N_5699);
nand U5929 (N_5929,N_5755,N_5782);
and U5930 (N_5930,N_5786,N_5661);
or U5931 (N_5931,N_5680,N_5741);
nor U5932 (N_5932,N_5634,N_5665);
nor U5933 (N_5933,N_5628,N_5751);
nand U5934 (N_5934,N_5634,N_5643);
nor U5935 (N_5935,N_5656,N_5752);
nor U5936 (N_5936,N_5679,N_5767);
nand U5937 (N_5937,N_5643,N_5765);
nor U5938 (N_5938,N_5721,N_5730);
xor U5939 (N_5939,N_5705,N_5715);
nand U5940 (N_5940,N_5744,N_5759);
xor U5941 (N_5941,N_5762,N_5799);
nand U5942 (N_5942,N_5740,N_5753);
nor U5943 (N_5943,N_5738,N_5616);
nor U5944 (N_5944,N_5695,N_5705);
and U5945 (N_5945,N_5775,N_5734);
xor U5946 (N_5946,N_5749,N_5605);
nor U5947 (N_5947,N_5655,N_5630);
xor U5948 (N_5948,N_5734,N_5688);
and U5949 (N_5949,N_5672,N_5630);
nand U5950 (N_5950,N_5717,N_5792);
nor U5951 (N_5951,N_5752,N_5749);
nor U5952 (N_5952,N_5623,N_5643);
or U5953 (N_5953,N_5668,N_5764);
nor U5954 (N_5954,N_5611,N_5792);
or U5955 (N_5955,N_5669,N_5667);
nand U5956 (N_5956,N_5600,N_5637);
and U5957 (N_5957,N_5690,N_5667);
or U5958 (N_5958,N_5697,N_5677);
and U5959 (N_5959,N_5744,N_5664);
and U5960 (N_5960,N_5762,N_5715);
xor U5961 (N_5961,N_5636,N_5746);
nor U5962 (N_5962,N_5727,N_5662);
nor U5963 (N_5963,N_5662,N_5608);
or U5964 (N_5964,N_5795,N_5660);
nor U5965 (N_5965,N_5629,N_5755);
or U5966 (N_5966,N_5682,N_5670);
and U5967 (N_5967,N_5678,N_5767);
and U5968 (N_5968,N_5692,N_5727);
nand U5969 (N_5969,N_5699,N_5758);
or U5970 (N_5970,N_5770,N_5702);
nand U5971 (N_5971,N_5639,N_5706);
or U5972 (N_5972,N_5641,N_5661);
or U5973 (N_5973,N_5713,N_5784);
nand U5974 (N_5974,N_5643,N_5616);
and U5975 (N_5975,N_5696,N_5633);
and U5976 (N_5976,N_5653,N_5649);
or U5977 (N_5977,N_5643,N_5747);
or U5978 (N_5978,N_5798,N_5629);
nor U5979 (N_5979,N_5633,N_5644);
or U5980 (N_5980,N_5736,N_5704);
nor U5981 (N_5981,N_5634,N_5629);
nor U5982 (N_5982,N_5727,N_5645);
and U5983 (N_5983,N_5601,N_5659);
nor U5984 (N_5984,N_5735,N_5664);
or U5985 (N_5985,N_5784,N_5755);
nand U5986 (N_5986,N_5631,N_5683);
or U5987 (N_5987,N_5742,N_5691);
nand U5988 (N_5988,N_5765,N_5763);
and U5989 (N_5989,N_5781,N_5600);
nand U5990 (N_5990,N_5618,N_5788);
nor U5991 (N_5991,N_5607,N_5758);
nor U5992 (N_5992,N_5796,N_5740);
and U5993 (N_5993,N_5689,N_5674);
nand U5994 (N_5994,N_5657,N_5727);
xor U5995 (N_5995,N_5678,N_5792);
xnor U5996 (N_5996,N_5655,N_5790);
xnor U5997 (N_5997,N_5733,N_5722);
or U5998 (N_5998,N_5647,N_5617);
or U5999 (N_5999,N_5782,N_5677);
and U6000 (N_6000,N_5816,N_5930);
nor U6001 (N_6001,N_5815,N_5952);
and U6002 (N_6002,N_5908,N_5905);
or U6003 (N_6003,N_5804,N_5928);
nand U6004 (N_6004,N_5951,N_5909);
or U6005 (N_6005,N_5808,N_5817);
nor U6006 (N_6006,N_5846,N_5894);
or U6007 (N_6007,N_5826,N_5964);
nand U6008 (N_6008,N_5861,N_5911);
nand U6009 (N_6009,N_5988,N_5802);
or U6010 (N_6010,N_5809,N_5903);
nor U6011 (N_6011,N_5874,N_5993);
xor U6012 (N_6012,N_5906,N_5933);
nor U6013 (N_6013,N_5866,N_5959);
nand U6014 (N_6014,N_5849,N_5892);
nor U6015 (N_6015,N_5879,N_5873);
and U6016 (N_6016,N_5961,N_5968);
nor U6017 (N_6017,N_5989,N_5818);
nor U6018 (N_6018,N_5848,N_5870);
xnor U6019 (N_6019,N_5991,N_5912);
and U6020 (N_6020,N_5992,N_5965);
xor U6021 (N_6021,N_5953,N_5925);
nor U6022 (N_6022,N_5958,N_5985);
and U6023 (N_6023,N_5916,N_5915);
nand U6024 (N_6024,N_5857,N_5843);
nand U6025 (N_6025,N_5881,N_5967);
or U6026 (N_6026,N_5910,N_5820);
nand U6027 (N_6027,N_5853,N_5929);
nor U6028 (N_6028,N_5976,N_5895);
or U6029 (N_6029,N_5875,N_5982);
xor U6030 (N_6030,N_5824,N_5842);
and U6031 (N_6031,N_5946,N_5887);
nor U6032 (N_6032,N_5821,N_5878);
nor U6033 (N_6033,N_5896,N_5858);
nand U6034 (N_6034,N_5863,N_5805);
nand U6035 (N_6035,N_5960,N_5859);
nand U6036 (N_6036,N_5987,N_5891);
and U6037 (N_6037,N_5830,N_5939);
nand U6038 (N_6038,N_5814,N_5867);
and U6039 (N_6039,N_5871,N_5913);
nand U6040 (N_6040,N_5917,N_5862);
and U6041 (N_6041,N_5810,N_5970);
nand U6042 (N_6042,N_5819,N_5851);
nor U6043 (N_6043,N_5944,N_5996);
or U6044 (N_6044,N_5995,N_5825);
nor U6045 (N_6045,N_5812,N_5977);
nor U6046 (N_6046,N_5948,N_5919);
or U6047 (N_6047,N_5837,N_5983);
nand U6048 (N_6048,N_5974,N_5957);
or U6049 (N_6049,N_5827,N_5907);
nor U6050 (N_6050,N_5803,N_5942);
nand U6051 (N_6051,N_5998,N_5923);
nand U6052 (N_6052,N_5860,N_5823);
nand U6053 (N_6053,N_5981,N_5836);
and U6054 (N_6054,N_5924,N_5828);
or U6055 (N_6055,N_5990,N_5832);
xnor U6056 (N_6056,N_5971,N_5885);
nand U6057 (N_6057,N_5954,N_5829);
or U6058 (N_6058,N_5893,N_5943);
and U6059 (N_6059,N_5868,N_5966);
and U6060 (N_6060,N_5940,N_5854);
nand U6061 (N_6061,N_5834,N_5955);
xnor U6062 (N_6062,N_5801,N_5922);
or U6063 (N_6063,N_5931,N_5950);
nor U6064 (N_6064,N_5947,N_5980);
or U6065 (N_6065,N_5888,N_5838);
and U6066 (N_6066,N_5877,N_5972);
nand U6067 (N_6067,N_5890,N_5844);
nand U6068 (N_6068,N_5926,N_5835);
and U6069 (N_6069,N_5855,N_5932);
and U6070 (N_6070,N_5872,N_5880);
and U6071 (N_6071,N_5833,N_5822);
nand U6072 (N_6072,N_5999,N_5869);
nand U6073 (N_6073,N_5921,N_5806);
and U6074 (N_6074,N_5986,N_5864);
xor U6075 (N_6075,N_5899,N_5898);
or U6076 (N_6076,N_5962,N_5938);
nor U6077 (N_6077,N_5984,N_5963);
nand U6078 (N_6078,N_5889,N_5945);
and U6079 (N_6079,N_5902,N_5969);
and U6080 (N_6080,N_5845,N_5839);
nand U6081 (N_6081,N_5800,N_5927);
or U6082 (N_6082,N_5841,N_5949);
xnor U6083 (N_6083,N_5876,N_5997);
nand U6084 (N_6084,N_5904,N_5883);
nor U6085 (N_6085,N_5918,N_5900);
nand U6086 (N_6086,N_5941,N_5937);
nand U6087 (N_6087,N_5934,N_5807);
nor U6088 (N_6088,N_5882,N_5840);
nand U6089 (N_6089,N_5956,N_5847);
nand U6090 (N_6090,N_5901,N_5831);
nand U6091 (N_6091,N_5813,N_5975);
and U6092 (N_6092,N_5886,N_5914);
nor U6093 (N_6093,N_5884,N_5994);
nor U6094 (N_6094,N_5897,N_5852);
nor U6095 (N_6095,N_5865,N_5973);
and U6096 (N_6096,N_5979,N_5936);
and U6097 (N_6097,N_5856,N_5978);
or U6098 (N_6098,N_5850,N_5935);
nand U6099 (N_6099,N_5920,N_5811);
or U6100 (N_6100,N_5917,N_5824);
or U6101 (N_6101,N_5926,N_5947);
and U6102 (N_6102,N_5982,N_5965);
and U6103 (N_6103,N_5934,N_5891);
and U6104 (N_6104,N_5912,N_5891);
nand U6105 (N_6105,N_5828,N_5876);
or U6106 (N_6106,N_5951,N_5859);
xnor U6107 (N_6107,N_5896,N_5847);
and U6108 (N_6108,N_5848,N_5971);
nand U6109 (N_6109,N_5964,N_5881);
nand U6110 (N_6110,N_5837,N_5844);
xor U6111 (N_6111,N_5806,N_5888);
nand U6112 (N_6112,N_5898,N_5842);
nor U6113 (N_6113,N_5971,N_5941);
nor U6114 (N_6114,N_5954,N_5824);
xnor U6115 (N_6115,N_5858,N_5829);
nand U6116 (N_6116,N_5866,N_5858);
and U6117 (N_6117,N_5808,N_5903);
nor U6118 (N_6118,N_5916,N_5836);
nand U6119 (N_6119,N_5866,N_5889);
nor U6120 (N_6120,N_5835,N_5915);
and U6121 (N_6121,N_5979,N_5861);
nand U6122 (N_6122,N_5947,N_5822);
and U6123 (N_6123,N_5973,N_5817);
or U6124 (N_6124,N_5818,N_5879);
and U6125 (N_6125,N_5967,N_5884);
nand U6126 (N_6126,N_5830,N_5930);
and U6127 (N_6127,N_5900,N_5922);
nor U6128 (N_6128,N_5848,N_5864);
nor U6129 (N_6129,N_5814,N_5885);
nor U6130 (N_6130,N_5823,N_5954);
and U6131 (N_6131,N_5937,N_5804);
and U6132 (N_6132,N_5906,N_5819);
or U6133 (N_6133,N_5990,N_5858);
nor U6134 (N_6134,N_5902,N_5918);
nor U6135 (N_6135,N_5831,N_5862);
or U6136 (N_6136,N_5927,N_5818);
nand U6137 (N_6137,N_5816,N_5828);
nor U6138 (N_6138,N_5898,N_5993);
or U6139 (N_6139,N_5914,N_5822);
or U6140 (N_6140,N_5820,N_5835);
or U6141 (N_6141,N_5849,N_5863);
and U6142 (N_6142,N_5837,N_5897);
or U6143 (N_6143,N_5804,N_5958);
nand U6144 (N_6144,N_5981,N_5932);
nand U6145 (N_6145,N_5884,N_5872);
nand U6146 (N_6146,N_5874,N_5840);
xnor U6147 (N_6147,N_5883,N_5818);
or U6148 (N_6148,N_5848,N_5984);
nor U6149 (N_6149,N_5963,N_5852);
and U6150 (N_6150,N_5824,N_5946);
xor U6151 (N_6151,N_5879,N_5976);
or U6152 (N_6152,N_5925,N_5932);
or U6153 (N_6153,N_5825,N_5989);
and U6154 (N_6154,N_5965,N_5953);
nand U6155 (N_6155,N_5870,N_5913);
and U6156 (N_6156,N_5900,N_5804);
nand U6157 (N_6157,N_5974,N_5818);
nor U6158 (N_6158,N_5831,N_5947);
nor U6159 (N_6159,N_5810,N_5876);
and U6160 (N_6160,N_5988,N_5986);
xnor U6161 (N_6161,N_5959,N_5989);
nor U6162 (N_6162,N_5817,N_5981);
xor U6163 (N_6163,N_5879,N_5866);
and U6164 (N_6164,N_5841,N_5816);
nand U6165 (N_6165,N_5995,N_5880);
and U6166 (N_6166,N_5970,N_5891);
or U6167 (N_6167,N_5951,N_5954);
nor U6168 (N_6168,N_5953,N_5890);
nand U6169 (N_6169,N_5905,N_5911);
xnor U6170 (N_6170,N_5826,N_5948);
and U6171 (N_6171,N_5974,N_5894);
or U6172 (N_6172,N_5942,N_5845);
nor U6173 (N_6173,N_5862,N_5850);
nor U6174 (N_6174,N_5979,N_5872);
nand U6175 (N_6175,N_5934,N_5816);
nand U6176 (N_6176,N_5868,N_5912);
nor U6177 (N_6177,N_5914,N_5936);
nor U6178 (N_6178,N_5827,N_5891);
nand U6179 (N_6179,N_5882,N_5846);
nand U6180 (N_6180,N_5959,N_5852);
or U6181 (N_6181,N_5893,N_5876);
and U6182 (N_6182,N_5892,N_5995);
nand U6183 (N_6183,N_5818,N_5874);
nor U6184 (N_6184,N_5804,N_5944);
nor U6185 (N_6185,N_5954,N_5985);
and U6186 (N_6186,N_5962,N_5807);
nand U6187 (N_6187,N_5885,N_5956);
or U6188 (N_6188,N_5950,N_5957);
and U6189 (N_6189,N_5808,N_5837);
nand U6190 (N_6190,N_5845,N_5861);
and U6191 (N_6191,N_5939,N_5849);
and U6192 (N_6192,N_5999,N_5827);
or U6193 (N_6193,N_5861,N_5901);
nor U6194 (N_6194,N_5856,N_5890);
or U6195 (N_6195,N_5860,N_5848);
xnor U6196 (N_6196,N_5939,N_5953);
or U6197 (N_6197,N_5816,N_5802);
nor U6198 (N_6198,N_5960,N_5803);
nor U6199 (N_6199,N_5998,N_5842);
and U6200 (N_6200,N_6127,N_6073);
nor U6201 (N_6201,N_6126,N_6132);
and U6202 (N_6202,N_6065,N_6137);
and U6203 (N_6203,N_6168,N_6020);
or U6204 (N_6204,N_6183,N_6199);
and U6205 (N_6205,N_6170,N_6110);
nor U6206 (N_6206,N_6023,N_6189);
nand U6207 (N_6207,N_6148,N_6094);
and U6208 (N_6208,N_6061,N_6048);
and U6209 (N_6209,N_6049,N_6143);
nor U6210 (N_6210,N_6090,N_6017);
and U6211 (N_6211,N_6008,N_6042);
nand U6212 (N_6212,N_6043,N_6003);
or U6213 (N_6213,N_6119,N_6033);
and U6214 (N_6214,N_6060,N_6192);
nor U6215 (N_6215,N_6153,N_6057);
or U6216 (N_6216,N_6150,N_6001);
nor U6217 (N_6217,N_6159,N_6149);
or U6218 (N_6218,N_6103,N_6051);
nor U6219 (N_6219,N_6147,N_6145);
or U6220 (N_6220,N_6022,N_6196);
nand U6221 (N_6221,N_6015,N_6026);
nand U6222 (N_6222,N_6117,N_6111);
or U6223 (N_6223,N_6059,N_6040);
nand U6224 (N_6224,N_6044,N_6013);
and U6225 (N_6225,N_6105,N_6114);
and U6226 (N_6226,N_6160,N_6169);
nor U6227 (N_6227,N_6056,N_6151);
and U6228 (N_6228,N_6144,N_6004);
nor U6229 (N_6229,N_6181,N_6108);
nor U6230 (N_6230,N_6064,N_6021);
and U6231 (N_6231,N_6188,N_6198);
and U6232 (N_6232,N_6138,N_6010);
nor U6233 (N_6233,N_6122,N_6082);
nor U6234 (N_6234,N_6070,N_6172);
nand U6235 (N_6235,N_6089,N_6068);
or U6236 (N_6236,N_6141,N_6165);
and U6237 (N_6237,N_6027,N_6152);
and U6238 (N_6238,N_6102,N_6037);
nor U6239 (N_6239,N_6133,N_6113);
nor U6240 (N_6240,N_6092,N_6054);
and U6241 (N_6241,N_6041,N_6036);
nor U6242 (N_6242,N_6128,N_6045);
or U6243 (N_6243,N_6055,N_6086);
or U6244 (N_6244,N_6072,N_6158);
nor U6245 (N_6245,N_6140,N_6193);
nor U6246 (N_6246,N_6115,N_6136);
or U6247 (N_6247,N_6075,N_6077);
xnor U6248 (N_6248,N_6069,N_6079);
and U6249 (N_6249,N_6104,N_6163);
nor U6250 (N_6250,N_6080,N_6050);
xor U6251 (N_6251,N_6078,N_6093);
xor U6252 (N_6252,N_6155,N_6175);
nand U6253 (N_6253,N_6171,N_6112);
nor U6254 (N_6254,N_6174,N_6028);
or U6255 (N_6255,N_6146,N_6074);
or U6256 (N_6256,N_6179,N_6118);
nand U6257 (N_6257,N_6030,N_6062);
nor U6258 (N_6258,N_6129,N_6035);
nor U6259 (N_6259,N_6025,N_6139);
or U6260 (N_6260,N_6047,N_6095);
or U6261 (N_6261,N_6098,N_6124);
nor U6262 (N_6262,N_6012,N_6076);
and U6263 (N_6263,N_6161,N_6000);
nor U6264 (N_6264,N_6187,N_6018);
nand U6265 (N_6265,N_6106,N_6011);
nor U6266 (N_6266,N_6002,N_6088);
and U6267 (N_6267,N_6007,N_6116);
or U6268 (N_6268,N_6123,N_6038);
or U6269 (N_6269,N_6186,N_6178);
and U6270 (N_6270,N_6087,N_6195);
or U6271 (N_6271,N_6034,N_6190);
and U6272 (N_6272,N_6180,N_6063);
nor U6273 (N_6273,N_6101,N_6052);
and U6274 (N_6274,N_6135,N_6100);
and U6275 (N_6275,N_6173,N_6016);
and U6276 (N_6276,N_6009,N_6058);
xnor U6277 (N_6277,N_6125,N_6019);
nor U6278 (N_6278,N_6131,N_6085);
and U6279 (N_6279,N_6014,N_6024);
nor U6280 (N_6280,N_6164,N_6005);
and U6281 (N_6281,N_6066,N_6029);
nor U6282 (N_6282,N_6091,N_6185);
or U6283 (N_6283,N_6177,N_6032);
nor U6284 (N_6284,N_6191,N_6154);
nor U6285 (N_6285,N_6067,N_6046);
nor U6286 (N_6286,N_6197,N_6157);
nand U6287 (N_6287,N_6142,N_6071);
and U6288 (N_6288,N_6167,N_6053);
nor U6289 (N_6289,N_6006,N_6194);
or U6290 (N_6290,N_6081,N_6097);
nor U6291 (N_6291,N_6162,N_6083);
xnor U6292 (N_6292,N_6134,N_6107);
and U6293 (N_6293,N_6182,N_6184);
xor U6294 (N_6294,N_6099,N_6130);
and U6295 (N_6295,N_6109,N_6176);
nor U6296 (N_6296,N_6120,N_6121);
and U6297 (N_6297,N_6156,N_6031);
or U6298 (N_6298,N_6084,N_6166);
xnor U6299 (N_6299,N_6039,N_6096);
and U6300 (N_6300,N_6144,N_6089);
and U6301 (N_6301,N_6065,N_6011);
or U6302 (N_6302,N_6004,N_6136);
and U6303 (N_6303,N_6070,N_6184);
nor U6304 (N_6304,N_6059,N_6131);
and U6305 (N_6305,N_6174,N_6055);
or U6306 (N_6306,N_6074,N_6116);
nor U6307 (N_6307,N_6175,N_6160);
or U6308 (N_6308,N_6011,N_6003);
and U6309 (N_6309,N_6010,N_6032);
and U6310 (N_6310,N_6000,N_6068);
nor U6311 (N_6311,N_6076,N_6007);
or U6312 (N_6312,N_6061,N_6185);
or U6313 (N_6313,N_6055,N_6175);
xor U6314 (N_6314,N_6097,N_6175);
xor U6315 (N_6315,N_6119,N_6176);
xnor U6316 (N_6316,N_6159,N_6084);
or U6317 (N_6317,N_6042,N_6092);
or U6318 (N_6318,N_6096,N_6130);
or U6319 (N_6319,N_6198,N_6030);
or U6320 (N_6320,N_6108,N_6193);
nor U6321 (N_6321,N_6171,N_6065);
nor U6322 (N_6322,N_6059,N_6096);
nand U6323 (N_6323,N_6098,N_6197);
nor U6324 (N_6324,N_6085,N_6142);
nor U6325 (N_6325,N_6057,N_6180);
nand U6326 (N_6326,N_6046,N_6123);
xor U6327 (N_6327,N_6117,N_6114);
xor U6328 (N_6328,N_6122,N_6187);
or U6329 (N_6329,N_6052,N_6137);
nand U6330 (N_6330,N_6091,N_6142);
or U6331 (N_6331,N_6174,N_6156);
nand U6332 (N_6332,N_6178,N_6062);
nor U6333 (N_6333,N_6181,N_6059);
or U6334 (N_6334,N_6023,N_6013);
nand U6335 (N_6335,N_6018,N_6194);
or U6336 (N_6336,N_6015,N_6088);
nor U6337 (N_6337,N_6166,N_6140);
or U6338 (N_6338,N_6132,N_6161);
xor U6339 (N_6339,N_6123,N_6047);
or U6340 (N_6340,N_6049,N_6128);
nor U6341 (N_6341,N_6059,N_6028);
nand U6342 (N_6342,N_6014,N_6005);
and U6343 (N_6343,N_6132,N_6198);
or U6344 (N_6344,N_6090,N_6113);
nor U6345 (N_6345,N_6097,N_6079);
xor U6346 (N_6346,N_6152,N_6068);
xnor U6347 (N_6347,N_6151,N_6000);
nand U6348 (N_6348,N_6125,N_6169);
xor U6349 (N_6349,N_6132,N_6007);
or U6350 (N_6350,N_6108,N_6188);
and U6351 (N_6351,N_6196,N_6061);
nand U6352 (N_6352,N_6050,N_6059);
nor U6353 (N_6353,N_6124,N_6025);
nor U6354 (N_6354,N_6187,N_6111);
and U6355 (N_6355,N_6080,N_6041);
or U6356 (N_6356,N_6148,N_6001);
xnor U6357 (N_6357,N_6035,N_6070);
or U6358 (N_6358,N_6156,N_6082);
nand U6359 (N_6359,N_6176,N_6083);
and U6360 (N_6360,N_6173,N_6181);
or U6361 (N_6361,N_6025,N_6027);
and U6362 (N_6362,N_6184,N_6118);
nor U6363 (N_6363,N_6124,N_6190);
nor U6364 (N_6364,N_6030,N_6038);
or U6365 (N_6365,N_6101,N_6035);
or U6366 (N_6366,N_6113,N_6054);
nor U6367 (N_6367,N_6041,N_6092);
and U6368 (N_6368,N_6111,N_6002);
nand U6369 (N_6369,N_6143,N_6031);
and U6370 (N_6370,N_6079,N_6103);
nand U6371 (N_6371,N_6022,N_6074);
xnor U6372 (N_6372,N_6043,N_6137);
nor U6373 (N_6373,N_6180,N_6106);
and U6374 (N_6374,N_6047,N_6017);
nor U6375 (N_6375,N_6116,N_6153);
nor U6376 (N_6376,N_6091,N_6098);
nand U6377 (N_6377,N_6152,N_6084);
xnor U6378 (N_6378,N_6044,N_6143);
nand U6379 (N_6379,N_6060,N_6035);
nand U6380 (N_6380,N_6050,N_6145);
nand U6381 (N_6381,N_6091,N_6178);
nor U6382 (N_6382,N_6169,N_6008);
nand U6383 (N_6383,N_6152,N_6077);
or U6384 (N_6384,N_6165,N_6128);
or U6385 (N_6385,N_6070,N_6155);
nor U6386 (N_6386,N_6030,N_6013);
and U6387 (N_6387,N_6094,N_6081);
nand U6388 (N_6388,N_6058,N_6071);
or U6389 (N_6389,N_6020,N_6076);
nand U6390 (N_6390,N_6124,N_6099);
nor U6391 (N_6391,N_6144,N_6112);
nand U6392 (N_6392,N_6112,N_6001);
xor U6393 (N_6393,N_6108,N_6060);
or U6394 (N_6394,N_6132,N_6101);
xor U6395 (N_6395,N_6149,N_6000);
and U6396 (N_6396,N_6006,N_6168);
nand U6397 (N_6397,N_6114,N_6188);
nand U6398 (N_6398,N_6108,N_6187);
and U6399 (N_6399,N_6129,N_6043);
nor U6400 (N_6400,N_6325,N_6332);
nor U6401 (N_6401,N_6383,N_6225);
or U6402 (N_6402,N_6276,N_6220);
or U6403 (N_6403,N_6208,N_6352);
and U6404 (N_6404,N_6290,N_6340);
xnor U6405 (N_6405,N_6275,N_6313);
xnor U6406 (N_6406,N_6282,N_6273);
nand U6407 (N_6407,N_6337,N_6360);
or U6408 (N_6408,N_6397,N_6288);
nand U6409 (N_6409,N_6326,N_6380);
or U6410 (N_6410,N_6212,N_6267);
nor U6411 (N_6411,N_6368,N_6201);
nor U6412 (N_6412,N_6219,N_6270);
nand U6413 (N_6413,N_6324,N_6364);
nor U6414 (N_6414,N_6293,N_6398);
nor U6415 (N_6415,N_6204,N_6287);
nor U6416 (N_6416,N_6256,N_6388);
nor U6417 (N_6417,N_6218,N_6215);
nand U6418 (N_6418,N_6314,N_6392);
or U6419 (N_6419,N_6378,N_6280);
or U6420 (N_6420,N_6214,N_6323);
and U6421 (N_6421,N_6330,N_6242);
and U6422 (N_6422,N_6381,N_6263);
nand U6423 (N_6423,N_6316,N_6306);
xor U6424 (N_6424,N_6370,N_6376);
nand U6425 (N_6425,N_6319,N_6346);
nand U6426 (N_6426,N_6229,N_6351);
and U6427 (N_6427,N_6265,N_6385);
nand U6428 (N_6428,N_6207,N_6240);
nand U6429 (N_6429,N_6343,N_6284);
nand U6430 (N_6430,N_6396,N_6234);
xor U6431 (N_6431,N_6205,N_6244);
nand U6432 (N_6432,N_6353,N_6252);
nand U6433 (N_6433,N_6236,N_6375);
or U6434 (N_6434,N_6302,N_6344);
or U6435 (N_6435,N_6298,N_6355);
or U6436 (N_6436,N_6329,N_6259);
nor U6437 (N_6437,N_6257,N_6338);
nand U6438 (N_6438,N_6292,N_6301);
or U6439 (N_6439,N_6248,N_6277);
xor U6440 (N_6440,N_6315,N_6361);
or U6441 (N_6441,N_6210,N_6300);
or U6442 (N_6442,N_6309,N_6349);
nand U6443 (N_6443,N_6320,N_6283);
nor U6444 (N_6444,N_6202,N_6232);
and U6445 (N_6445,N_6241,N_6262);
nand U6446 (N_6446,N_6391,N_6373);
or U6447 (N_6447,N_6399,N_6255);
or U6448 (N_6448,N_6253,N_6243);
nand U6449 (N_6449,N_6379,N_6278);
nor U6450 (N_6450,N_6228,N_6251);
xor U6451 (N_6451,N_6365,N_6356);
nand U6452 (N_6452,N_6374,N_6217);
or U6453 (N_6453,N_6341,N_6328);
and U6454 (N_6454,N_6239,N_6310);
and U6455 (N_6455,N_6258,N_6390);
and U6456 (N_6456,N_6261,N_6289);
nand U6457 (N_6457,N_6203,N_6221);
and U6458 (N_6458,N_6345,N_6359);
or U6459 (N_6459,N_6393,N_6387);
and U6460 (N_6460,N_6372,N_6342);
xor U6461 (N_6461,N_6333,N_6311);
nor U6462 (N_6462,N_6224,N_6335);
nand U6463 (N_6463,N_6297,N_6213);
nor U6464 (N_6464,N_6303,N_6296);
xor U6465 (N_6465,N_6233,N_6264);
or U6466 (N_6466,N_6331,N_6336);
nand U6467 (N_6467,N_6366,N_6238);
xor U6468 (N_6468,N_6295,N_6395);
nor U6469 (N_6469,N_6235,N_6305);
nor U6470 (N_6470,N_6227,N_6371);
or U6471 (N_6471,N_6386,N_6294);
or U6472 (N_6472,N_6307,N_6222);
or U6473 (N_6473,N_6272,N_6249);
or U6474 (N_6474,N_6285,N_6206);
nand U6475 (N_6475,N_6317,N_6377);
or U6476 (N_6476,N_6268,N_6304);
and U6477 (N_6477,N_6291,N_6274);
nor U6478 (N_6478,N_6237,N_6281);
or U6479 (N_6479,N_6394,N_6231);
nor U6480 (N_6480,N_6357,N_6247);
or U6481 (N_6481,N_6347,N_6216);
nand U6482 (N_6482,N_6354,N_6250);
nor U6483 (N_6483,N_6350,N_6384);
or U6484 (N_6484,N_6382,N_6322);
and U6485 (N_6485,N_6269,N_6266);
nor U6486 (N_6486,N_6348,N_6245);
and U6487 (N_6487,N_6339,N_6363);
xnor U6488 (N_6488,N_6254,N_6369);
xor U6489 (N_6489,N_6334,N_6367);
or U6490 (N_6490,N_6286,N_6246);
and U6491 (N_6491,N_6200,N_6271);
nor U6492 (N_6492,N_6312,N_6358);
xor U6493 (N_6493,N_6279,N_6299);
nand U6494 (N_6494,N_6260,N_6308);
and U6495 (N_6495,N_6230,N_6223);
nor U6496 (N_6496,N_6327,N_6209);
nand U6497 (N_6497,N_6318,N_6211);
and U6498 (N_6498,N_6226,N_6321);
and U6499 (N_6499,N_6362,N_6389);
and U6500 (N_6500,N_6240,N_6282);
nor U6501 (N_6501,N_6318,N_6377);
and U6502 (N_6502,N_6325,N_6224);
xor U6503 (N_6503,N_6302,N_6329);
or U6504 (N_6504,N_6292,N_6237);
nor U6505 (N_6505,N_6202,N_6380);
and U6506 (N_6506,N_6378,N_6202);
or U6507 (N_6507,N_6246,N_6269);
nand U6508 (N_6508,N_6366,N_6347);
nand U6509 (N_6509,N_6310,N_6357);
nor U6510 (N_6510,N_6321,N_6280);
and U6511 (N_6511,N_6259,N_6268);
nand U6512 (N_6512,N_6372,N_6258);
nor U6513 (N_6513,N_6350,N_6267);
and U6514 (N_6514,N_6207,N_6276);
or U6515 (N_6515,N_6362,N_6349);
nand U6516 (N_6516,N_6238,N_6379);
or U6517 (N_6517,N_6372,N_6268);
and U6518 (N_6518,N_6292,N_6206);
nand U6519 (N_6519,N_6208,N_6211);
and U6520 (N_6520,N_6243,N_6236);
nand U6521 (N_6521,N_6292,N_6288);
nor U6522 (N_6522,N_6334,N_6371);
xnor U6523 (N_6523,N_6339,N_6217);
or U6524 (N_6524,N_6243,N_6371);
and U6525 (N_6525,N_6394,N_6268);
nand U6526 (N_6526,N_6344,N_6298);
nand U6527 (N_6527,N_6372,N_6262);
and U6528 (N_6528,N_6322,N_6303);
and U6529 (N_6529,N_6346,N_6347);
nand U6530 (N_6530,N_6304,N_6266);
or U6531 (N_6531,N_6353,N_6354);
nor U6532 (N_6532,N_6390,N_6346);
nor U6533 (N_6533,N_6324,N_6367);
or U6534 (N_6534,N_6356,N_6245);
nor U6535 (N_6535,N_6329,N_6220);
nand U6536 (N_6536,N_6370,N_6365);
xor U6537 (N_6537,N_6388,N_6285);
xnor U6538 (N_6538,N_6380,N_6354);
nand U6539 (N_6539,N_6223,N_6321);
nor U6540 (N_6540,N_6326,N_6320);
and U6541 (N_6541,N_6212,N_6214);
nor U6542 (N_6542,N_6272,N_6375);
and U6543 (N_6543,N_6337,N_6376);
nand U6544 (N_6544,N_6382,N_6391);
or U6545 (N_6545,N_6265,N_6270);
nor U6546 (N_6546,N_6306,N_6278);
xnor U6547 (N_6547,N_6204,N_6320);
or U6548 (N_6548,N_6345,N_6250);
nand U6549 (N_6549,N_6287,N_6341);
nor U6550 (N_6550,N_6325,N_6395);
and U6551 (N_6551,N_6219,N_6290);
nor U6552 (N_6552,N_6396,N_6281);
or U6553 (N_6553,N_6301,N_6277);
or U6554 (N_6554,N_6350,N_6250);
or U6555 (N_6555,N_6344,N_6268);
and U6556 (N_6556,N_6348,N_6397);
nor U6557 (N_6557,N_6251,N_6327);
and U6558 (N_6558,N_6392,N_6284);
and U6559 (N_6559,N_6395,N_6357);
nand U6560 (N_6560,N_6386,N_6311);
and U6561 (N_6561,N_6366,N_6352);
and U6562 (N_6562,N_6232,N_6305);
xor U6563 (N_6563,N_6263,N_6321);
nand U6564 (N_6564,N_6384,N_6269);
nor U6565 (N_6565,N_6220,N_6362);
xnor U6566 (N_6566,N_6241,N_6339);
nand U6567 (N_6567,N_6335,N_6396);
nor U6568 (N_6568,N_6284,N_6298);
and U6569 (N_6569,N_6243,N_6224);
nand U6570 (N_6570,N_6210,N_6335);
nand U6571 (N_6571,N_6278,N_6397);
or U6572 (N_6572,N_6360,N_6234);
and U6573 (N_6573,N_6208,N_6387);
and U6574 (N_6574,N_6270,N_6230);
or U6575 (N_6575,N_6336,N_6232);
nand U6576 (N_6576,N_6219,N_6386);
or U6577 (N_6577,N_6316,N_6347);
or U6578 (N_6578,N_6273,N_6301);
or U6579 (N_6579,N_6249,N_6208);
nor U6580 (N_6580,N_6212,N_6336);
nand U6581 (N_6581,N_6347,N_6279);
nor U6582 (N_6582,N_6334,N_6369);
and U6583 (N_6583,N_6263,N_6359);
nor U6584 (N_6584,N_6221,N_6316);
nor U6585 (N_6585,N_6396,N_6359);
and U6586 (N_6586,N_6248,N_6313);
nand U6587 (N_6587,N_6386,N_6245);
or U6588 (N_6588,N_6269,N_6335);
and U6589 (N_6589,N_6368,N_6299);
nand U6590 (N_6590,N_6256,N_6284);
or U6591 (N_6591,N_6230,N_6287);
and U6592 (N_6592,N_6350,N_6225);
and U6593 (N_6593,N_6386,N_6334);
xor U6594 (N_6594,N_6317,N_6209);
nand U6595 (N_6595,N_6282,N_6275);
or U6596 (N_6596,N_6373,N_6220);
or U6597 (N_6597,N_6228,N_6312);
or U6598 (N_6598,N_6358,N_6275);
nand U6599 (N_6599,N_6295,N_6250);
nand U6600 (N_6600,N_6533,N_6525);
nand U6601 (N_6601,N_6414,N_6582);
and U6602 (N_6602,N_6500,N_6412);
or U6603 (N_6603,N_6438,N_6418);
nand U6604 (N_6604,N_6545,N_6492);
xor U6605 (N_6605,N_6439,N_6405);
nand U6606 (N_6606,N_6576,N_6477);
or U6607 (N_6607,N_6513,N_6583);
xor U6608 (N_6608,N_6512,N_6495);
and U6609 (N_6609,N_6486,N_6558);
or U6610 (N_6610,N_6510,N_6487);
or U6611 (N_6611,N_6449,N_6496);
and U6612 (N_6612,N_6432,N_6413);
nor U6613 (N_6613,N_6591,N_6419);
or U6614 (N_6614,N_6471,N_6503);
nand U6615 (N_6615,N_6567,N_6410);
nor U6616 (N_6616,N_6524,N_6521);
nor U6617 (N_6617,N_6548,N_6593);
nor U6618 (N_6618,N_6520,N_6584);
and U6619 (N_6619,N_6430,N_6522);
or U6620 (N_6620,N_6435,N_6482);
xnor U6621 (N_6621,N_6571,N_6407);
and U6622 (N_6622,N_6490,N_6401);
xnor U6623 (N_6623,N_6494,N_6462);
xor U6624 (N_6624,N_6529,N_6526);
nand U6625 (N_6625,N_6466,N_6577);
or U6626 (N_6626,N_6587,N_6504);
nor U6627 (N_6627,N_6458,N_6416);
or U6628 (N_6628,N_6427,N_6484);
and U6629 (N_6629,N_6590,N_6426);
nand U6630 (N_6630,N_6552,N_6415);
or U6631 (N_6631,N_6489,N_6443);
or U6632 (N_6632,N_6554,N_6553);
or U6633 (N_6633,N_6528,N_6517);
nand U6634 (N_6634,N_6408,N_6542);
nand U6635 (N_6635,N_6476,N_6537);
nor U6636 (N_6636,N_6468,N_6403);
nand U6637 (N_6637,N_6441,N_6561);
or U6638 (N_6638,N_6595,N_6469);
nand U6639 (N_6639,N_6580,N_6498);
xor U6640 (N_6640,N_6433,N_6404);
nor U6641 (N_6641,N_6511,N_6546);
and U6642 (N_6642,N_6472,N_6515);
nor U6643 (N_6643,N_6444,N_6569);
xor U6644 (N_6644,N_6594,N_6488);
and U6645 (N_6645,N_6452,N_6539);
nor U6646 (N_6646,N_6454,N_6457);
nor U6647 (N_6647,N_6464,N_6564);
xor U6648 (N_6648,N_6420,N_6448);
or U6649 (N_6649,N_6507,N_6586);
nor U6650 (N_6650,N_6424,N_6423);
nand U6651 (N_6651,N_6455,N_6480);
nand U6652 (N_6652,N_6575,N_6598);
nand U6653 (N_6653,N_6599,N_6499);
nand U6654 (N_6654,N_6400,N_6442);
xnor U6655 (N_6655,N_6453,N_6565);
nor U6656 (N_6656,N_6579,N_6562);
and U6657 (N_6657,N_6570,N_6436);
nor U6658 (N_6658,N_6541,N_6550);
and U6659 (N_6659,N_6514,N_6578);
nand U6660 (N_6660,N_6437,N_6516);
or U6661 (N_6661,N_6497,N_6532);
or U6662 (N_6662,N_6589,N_6588);
xnor U6663 (N_6663,N_6465,N_6535);
or U6664 (N_6664,N_6456,N_6483);
nand U6665 (N_6665,N_6451,N_6573);
nand U6666 (N_6666,N_6447,N_6509);
nor U6667 (N_6667,N_6460,N_6481);
nor U6668 (N_6668,N_6543,N_6425);
and U6669 (N_6669,N_6474,N_6402);
xnor U6670 (N_6670,N_6461,N_6429);
nor U6671 (N_6671,N_6563,N_6502);
and U6672 (N_6672,N_6479,N_6417);
and U6673 (N_6673,N_6549,N_6534);
and U6674 (N_6674,N_6556,N_6572);
nand U6675 (N_6675,N_6446,N_6478);
and U6676 (N_6676,N_6566,N_6523);
or U6677 (N_6677,N_6463,N_6544);
xor U6678 (N_6678,N_6559,N_6538);
or U6679 (N_6679,N_6597,N_6519);
xor U6680 (N_6680,N_6585,N_6581);
nand U6681 (N_6681,N_6527,N_6536);
nor U6682 (N_6682,N_6470,N_6518);
and U6683 (N_6683,N_6434,N_6568);
nand U6684 (N_6684,N_6411,N_6445);
nand U6685 (N_6685,N_6557,N_6592);
and U6686 (N_6686,N_6505,N_6547);
and U6687 (N_6687,N_6473,N_6551);
nand U6688 (N_6688,N_6467,N_6493);
nand U6689 (N_6689,N_6574,N_6450);
or U6690 (N_6690,N_6540,N_6530);
and U6691 (N_6691,N_6431,N_6501);
nand U6692 (N_6692,N_6459,N_6406);
nand U6693 (N_6693,N_6409,N_6421);
nor U6694 (N_6694,N_6531,N_6440);
and U6695 (N_6695,N_6422,N_6485);
xnor U6696 (N_6696,N_6560,N_6491);
or U6697 (N_6697,N_6555,N_6506);
or U6698 (N_6698,N_6475,N_6508);
nand U6699 (N_6699,N_6428,N_6596);
or U6700 (N_6700,N_6441,N_6419);
and U6701 (N_6701,N_6453,N_6475);
xnor U6702 (N_6702,N_6512,N_6577);
or U6703 (N_6703,N_6413,N_6596);
or U6704 (N_6704,N_6403,N_6431);
nand U6705 (N_6705,N_6464,N_6578);
nor U6706 (N_6706,N_6562,N_6480);
or U6707 (N_6707,N_6547,N_6561);
nor U6708 (N_6708,N_6404,N_6466);
nor U6709 (N_6709,N_6421,N_6405);
or U6710 (N_6710,N_6495,N_6532);
nor U6711 (N_6711,N_6430,N_6566);
or U6712 (N_6712,N_6460,N_6594);
xnor U6713 (N_6713,N_6588,N_6561);
nor U6714 (N_6714,N_6536,N_6517);
nand U6715 (N_6715,N_6584,N_6500);
nor U6716 (N_6716,N_6450,N_6581);
nand U6717 (N_6717,N_6402,N_6575);
and U6718 (N_6718,N_6453,N_6519);
nor U6719 (N_6719,N_6534,N_6489);
nand U6720 (N_6720,N_6564,N_6417);
or U6721 (N_6721,N_6461,N_6416);
xnor U6722 (N_6722,N_6525,N_6462);
or U6723 (N_6723,N_6541,N_6571);
xnor U6724 (N_6724,N_6545,N_6557);
nor U6725 (N_6725,N_6419,N_6533);
or U6726 (N_6726,N_6503,N_6502);
xnor U6727 (N_6727,N_6422,N_6520);
and U6728 (N_6728,N_6570,N_6434);
or U6729 (N_6729,N_6407,N_6587);
xnor U6730 (N_6730,N_6453,N_6512);
nand U6731 (N_6731,N_6483,N_6435);
nand U6732 (N_6732,N_6544,N_6592);
or U6733 (N_6733,N_6541,N_6537);
and U6734 (N_6734,N_6490,N_6461);
nand U6735 (N_6735,N_6529,N_6528);
nor U6736 (N_6736,N_6587,N_6569);
nand U6737 (N_6737,N_6441,N_6411);
or U6738 (N_6738,N_6491,N_6540);
nor U6739 (N_6739,N_6455,N_6430);
and U6740 (N_6740,N_6411,N_6491);
nor U6741 (N_6741,N_6539,N_6547);
nand U6742 (N_6742,N_6597,N_6465);
and U6743 (N_6743,N_6473,N_6469);
nor U6744 (N_6744,N_6551,N_6442);
nand U6745 (N_6745,N_6474,N_6459);
and U6746 (N_6746,N_6557,N_6585);
nor U6747 (N_6747,N_6490,N_6550);
nor U6748 (N_6748,N_6456,N_6402);
or U6749 (N_6749,N_6477,N_6471);
nand U6750 (N_6750,N_6578,N_6525);
and U6751 (N_6751,N_6439,N_6544);
nor U6752 (N_6752,N_6438,N_6532);
nand U6753 (N_6753,N_6569,N_6409);
nand U6754 (N_6754,N_6460,N_6470);
nand U6755 (N_6755,N_6532,N_6595);
nand U6756 (N_6756,N_6449,N_6591);
nand U6757 (N_6757,N_6450,N_6421);
or U6758 (N_6758,N_6422,N_6539);
nand U6759 (N_6759,N_6546,N_6570);
and U6760 (N_6760,N_6486,N_6488);
nor U6761 (N_6761,N_6570,N_6497);
nor U6762 (N_6762,N_6489,N_6481);
and U6763 (N_6763,N_6529,N_6480);
and U6764 (N_6764,N_6464,N_6570);
nor U6765 (N_6765,N_6492,N_6469);
and U6766 (N_6766,N_6431,N_6523);
nor U6767 (N_6767,N_6543,N_6592);
or U6768 (N_6768,N_6593,N_6481);
nand U6769 (N_6769,N_6533,N_6516);
nand U6770 (N_6770,N_6449,N_6436);
and U6771 (N_6771,N_6421,N_6539);
nor U6772 (N_6772,N_6464,N_6518);
and U6773 (N_6773,N_6545,N_6498);
and U6774 (N_6774,N_6400,N_6494);
and U6775 (N_6775,N_6583,N_6541);
nor U6776 (N_6776,N_6599,N_6461);
or U6777 (N_6777,N_6566,N_6512);
nor U6778 (N_6778,N_6547,N_6599);
or U6779 (N_6779,N_6534,N_6533);
and U6780 (N_6780,N_6535,N_6534);
and U6781 (N_6781,N_6505,N_6451);
nand U6782 (N_6782,N_6512,N_6501);
nor U6783 (N_6783,N_6539,N_6526);
and U6784 (N_6784,N_6410,N_6425);
xnor U6785 (N_6785,N_6516,N_6519);
nand U6786 (N_6786,N_6536,N_6589);
nand U6787 (N_6787,N_6417,N_6430);
nand U6788 (N_6788,N_6519,N_6407);
and U6789 (N_6789,N_6468,N_6507);
or U6790 (N_6790,N_6421,N_6565);
xor U6791 (N_6791,N_6555,N_6586);
or U6792 (N_6792,N_6511,N_6479);
and U6793 (N_6793,N_6474,N_6403);
xor U6794 (N_6794,N_6486,N_6400);
nor U6795 (N_6795,N_6568,N_6513);
xnor U6796 (N_6796,N_6566,N_6508);
nor U6797 (N_6797,N_6509,N_6541);
or U6798 (N_6798,N_6595,N_6527);
nand U6799 (N_6799,N_6412,N_6442);
or U6800 (N_6800,N_6786,N_6760);
or U6801 (N_6801,N_6702,N_6726);
nor U6802 (N_6802,N_6699,N_6703);
nor U6803 (N_6803,N_6776,N_6664);
nand U6804 (N_6804,N_6701,N_6693);
and U6805 (N_6805,N_6720,N_6649);
nor U6806 (N_6806,N_6688,N_6736);
xor U6807 (N_6807,N_6755,N_6759);
or U6808 (N_6808,N_6705,N_6644);
nand U6809 (N_6809,N_6606,N_6739);
and U6810 (N_6810,N_6653,N_6793);
and U6811 (N_6811,N_6682,N_6781);
and U6812 (N_6812,N_6747,N_6799);
or U6813 (N_6813,N_6618,N_6667);
nor U6814 (N_6814,N_6640,N_6729);
or U6815 (N_6815,N_6731,N_6609);
and U6816 (N_6816,N_6651,N_6741);
or U6817 (N_6817,N_6629,N_6764);
nand U6818 (N_6818,N_6724,N_6718);
nand U6819 (N_6819,N_6662,N_6633);
and U6820 (N_6820,N_6673,N_6770);
nand U6821 (N_6821,N_6738,N_6614);
and U6822 (N_6822,N_6771,N_6628);
nand U6823 (N_6823,N_6757,N_6773);
xnor U6824 (N_6824,N_6671,N_6756);
xor U6825 (N_6825,N_6743,N_6732);
nor U6826 (N_6826,N_6632,N_6767);
nor U6827 (N_6827,N_6657,N_6694);
xnor U6828 (N_6828,N_6650,N_6774);
nor U6829 (N_6829,N_6666,N_6615);
nor U6830 (N_6830,N_6636,N_6707);
or U6831 (N_6831,N_6772,N_6677);
and U6832 (N_6832,N_6656,N_6645);
and U6833 (N_6833,N_6601,N_6734);
and U6834 (N_6834,N_6605,N_6691);
or U6835 (N_6835,N_6658,N_6680);
or U6836 (N_6836,N_6692,N_6621);
and U6837 (N_6837,N_6622,N_6695);
or U6838 (N_6838,N_6643,N_6740);
nand U6839 (N_6839,N_6775,N_6672);
nor U6840 (N_6840,N_6730,N_6678);
nand U6841 (N_6841,N_6674,N_6608);
and U6842 (N_6842,N_6762,N_6652);
and U6843 (N_6843,N_6654,N_6696);
xor U6844 (N_6844,N_6780,N_6768);
and U6845 (N_6845,N_6709,N_6721);
xnor U6846 (N_6846,N_6687,N_6635);
nand U6847 (N_6847,N_6711,N_6625);
and U6848 (N_6848,N_6665,N_6675);
nand U6849 (N_6849,N_6727,N_6681);
and U6850 (N_6850,N_6697,N_6765);
or U6851 (N_6851,N_6600,N_6716);
and U6852 (N_6852,N_6642,N_6790);
or U6853 (N_6853,N_6639,N_6602);
and U6854 (N_6854,N_6616,N_6728);
and U6855 (N_6855,N_6604,N_6660);
nand U6856 (N_6856,N_6670,N_6723);
nand U6857 (N_6857,N_6637,N_6783);
or U6858 (N_6858,N_6782,N_6648);
or U6859 (N_6859,N_6769,N_6712);
nand U6860 (N_6860,N_6749,N_6742);
nand U6861 (N_6861,N_6626,N_6631);
xor U6862 (N_6862,N_6714,N_6686);
and U6863 (N_6863,N_6638,N_6634);
and U6864 (N_6864,N_6794,N_6763);
nor U6865 (N_6865,N_6704,N_6778);
nand U6866 (N_6866,N_6722,N_6684);
or U6867 (N_6867,N_6777,N_6607);
and U6868 (N_6868,N_6766,N_6737);
xnor U6869 (N_6869,N_6754,N_6717);
nand U6870 (N_6870,N_6708,N_6685);
nand U6871 (N_6871,N_6706,N_6624);
xnor U6872 (N_6872,N_6745,N_6611);
nand U6873 (N_6873,N_6795,N_6746);
nand U6874 (N_6874,N_6779,N_6627);
and U6875 (N_6875,N_6751,N_6784);
nand U6876 (N_6876,N_6752,N_6715);
nand U6877 (N_6877,N_6676,N_6619);
nand U6878 (N_6878,N_6797,N_6787);
nand U6879 (N_6879,N_6620,N_6744);
nor U6880 (N_6880,N_6612,N_6710);
nand U6881 (N_6881,N_6646,N_6735);
nand U6882 (N_6882,N_6719,N_6700);
and U6883 (N_6883,N_6750,N_6798);
nand U6884 (N_6884,N_6789,N_6796);
or U6885 (N_6885,N_6690,N_6661);
or U6886 (N_6886,N_6630,N_6617);
nor U6887 (N_6887,N_6659,N_6623);
nor U6888 (N_6888,N_6610,N_6679);
nor U6889 (N_6889,N_6788,N_6733);
and U6890 (N_6890,N_6613,N_6663);
nand U6891 (N_6891,N_6683,N_6669);
or U6892 (N_6892,N_6725,N_6647);
and U6893 (N_6893,N_6758,N_6785);
and U6894 (N_6894,N_6761,N_6603);
nand U6895 (N_6895,N_6753,N_6689);
nand U6896 (N_6896,N_6748,N_6641);
nor U6897 (N_6897,N_6791,N_6698);
and U6898 (N_6898,N_6655,N_6713);
nor U6899 (N_6899,N_6792,N_6668);
nor U6900 (N_6900,N_6642,N_6721);
nor U6901 (N_6901,N_6702,N_6648);
nor U6902 (N_6902,N_6786,N_6706);
nand U6903 (N_6903,N_6651,N_6716);
xnor U6904 (N_6904,N_6777,N_6688);
or U6905 (N_6905,N_6674,N_6667);
nand U6906 (N_6906,N_6704,N_6696);
and U6907 (N_6907,N_6600,N_6756);
or U6908 (N_6908,N_6759,N_6788);
nand U6909 (N_6909,N_6744,N_6720);
or U6910 (N_6910,N_6778,N_6663);
and U6911 (N_6911,N_6625,N_6720);
nor U6912 (N_6912,N_6765,N_6657);
nor U6913 (N_6913,N_6674,N_6653);
nand U6914 (N_6914,N_6676,N_6775);
or U6915 (N_6915,N_6755,N_6695);
and U6916 (N_6916,N_6706,N_6628);
nand U6917 (N_6917,N_6668,N_6635);
nor U6918 (N_6918,N_6606,N_6641);
and U6919 (N_6919,N_6777,N_6708);
or U6920 (N_6920,N_6757,N_6767);
nand U6921 (N_6921,N_6768,N_6755);
nand U6922 (N_6922,N_6739,N_6722);
or U6923 (N_6923,N_6713,N_6715);
and U6924 (N_6924,N_6697,N_6751);
nor U6925 (N_6925,N_6740,N_6629);
and U6926 (N_6926,N_6641,N_6698);
xor U6927 (N_6927,N_6784,N_6629);
or U6928 (N_6928,N_6684,N_6699);
nor U6929 (N_6929,N_6681,N_6601);
nor U6930 (N_6930,N_6756,N_6759);
xnor U6931 (N_6931,N_6653,N_6663);
nand U6932 (N_6932,N_6621,N_6737);
and U6933 (N_6933,N_6761,N_6782);
nor U6934 (N_6934,N_6606,N_6609);
nand U6935 (N_6935,N_6758,N_6702);
nand U6936 (N_6936,N_6728,N_6628);
nand U6937 (N_6937,N_6744,N_6636);
nor U6938 (N_6938,N_6687,N_6601);
and U6939 (N_6939,N_6752,N_6695);
nand U6940 (N_6940,N_6680,N_6603);
or U6941 (N_6941,N_6630,N_6650);
nand U6942 (N_6942,N_6604,N_6739);
nand U6943 (N_6943,N_6771,N_6635);
nand U6944 (N_6944,N_6791,N_6762);
nand U6945 (N_6945,N_6794,N_6680);
or U6946 (N_6946,N_6667,N_6728);
or U6947 (N_6947,N_6780,N_6608);
nand U6948 (N_6948,N_6664,N_6795);
and U6949 (N_6949,N_6742,N_6676);
xor U6950 (N_6950,N_6637,N_6606);
nand U6951 (N_6951,N_6608,N_6782);
or U6952 (N_6952,N_6765,N_6769);
nor U6953 (N_6953,N_6705,N_6680);
nand U6954 (N_6954,N_6697,N_6717);
and U6955 (N_6955,N_6645,N_6704);
nand U6956 (N_6956,N_6656,N_6778);
or U6957 (N_6957,N_6769,N_6777);
nand U6958 (N_6958,N_6743,N_6736);
nor U6959 (N_6959,N_6729,N_6743);
nand U6960 (N_6960,N_6711,N_6602);
nand U6961 (N_6961,N_6689,N_6719);
or U6962 (N_6962,N_6736,N_6675);
and U6963 (N_6963,N_6635,N_6716);
nor U6964 (N_6964,N_6638,N_6689);
nor U6965 (N_6965,N_6638,N_6707);
or U6966 (N_6966,N_6694,N_6697);
nand U6967 (N_6967,N_6664,N_6658);
or U6968 (N_6968,N_6633,N_6701);
nor U6969 (N_6969,N_6640,N_6652);
nor U6970 (N_6970,N_6699,N_6674);
nor U6971 (N_6971,N_6629,N_6772);
or U6972 (N_6972,N_6749,N_6662);
or U6973 (N_6973,N_6664,N_6637);
nand U6974 (N_6974,N_6644,N_6786);
nor U6975 (N_6975,N_6766,N_6681);
and U6976 (N_6976,N_6765,N_6720);
nand U6977 (N_6977,N_6721,N_6682);
or U6978 (N_6978,N_6659,N_6656);
nor U6979 (N_6979,N_6776,N_6683);
xor U6980 (N_6980,N_6760,N_6607);
or U6981 (N_6981,N_6742,N_6750);
and U6982 (N_6982,N_6608,N_6611);
nor U6983 (N_6983,N_6633,N_6660);
and U6984 (N_6984,N_6736,N_6601);
nand U6985 (N_6985,N_6750,N_6706);
nor U6986 (N_6986,N_6743,N_6675);
xor U6987 (N_6987,N_6779,N_6604);
xnor U6988 (N_6988,N_6659,N_6742);
nor U6989 (N_6989,N_6760,N_6761);
nor U6990 (N_6990,N_6678,N_6796);
nor U6991 (N_6991,N_6709,N_6668);
or U6992 (N_6992,N_6672,N_6708);
or U6993 (N_6993,N_6748,N_6620);
nor U6994 (N_6994,N_6763,N_6753);
nand U6995 (N_6995,N_6663,N_6743);
nor U6996 (N_6996,N_6666,N_6701);
nor U6997 (N_6997,N_6733,N_6752);
nor U6998 (N_6998,N_6741,N_6739);
or U6999 (N_6999,N_6665,N_6796);
nand U7000 (N_7000,N_6923,N_6881);
or U7001 (N_7001,N_6838,N_6896);
nor U7002 (N_7002,N_6824,N_6976);
or U7003 (N_7003,N_6915,N_6959);
xnor U7004 (N_7004,N_6984,N_6948);
xnor U7005 (N_7005,N_6912,N_6825);
nand U7006 (N_7006,N_6835,N_6810);
and U7007 (N_7007,N_6857,N_6911);
or U7008 (N_7008,N_6945,N_6919);
or U7009 (N_7009,N_6934,N_6932);
and U7010 (N_7010,N_6986,N_6843);
and U7011 (N_7011,N_6830,N_6883);
nor U7012 (N_7012,N_6929,N_6814);
or U7013 (N_7013,N_6858,N_6819);
and U7014 (N_7014,N_6813,N_6808);
and U7015 (N_7015,N_6886,N_6855);
nand U7016 (N_7016,N_6856,N_6894);
and U7017 (N_7017,N_6925,N_6867);
or U7018 (N_7018,N_6955,N_6837);
and U7019 (N_7019,N_6963,N_6887);
and U7020 (N_7020,N_6836,N_6816);
and U7021 (N_7021,N_6906,N_6820);
nand U7022 (N_7022,N_6943,N_6924);
nand U7023 (N_7023,N_6869,N_6998);
or U7024 (N_7024,N_6965,N_6922);
and U7025 (N_7025,N_6958,N_6988);
and U7026 (N_7026,N_6833,N_6954);
nand U7027 (N_7027,N_6875,N_6827);
or U7028 (N_7028,N_6975,N_6996);
nor U7029 (N_7029,N_6822,N_6933);
nor U7030 (N_7030,N_6844,N_6981);
nand U7031 (N_7031,N_6993,N_6885);
nand U7032 (N_7032,N_6862,N_6940);
nand U7033 (N_7033,N_6846,N_6851);
nand U7034 (N_7034,N_6980,N_6864);
xnor U7035 (N_7035,N_6860,N_6917);
or U7036 (N_7036,N_6870,N_6942);
or U7037 (N_7037,N_6977,N_6889);
xor U7038 (N_7038,N_6845,N_6903);
and U7039 (N_7039,N_6898,N_6831);
nand U7040 (N_7040,N_6890,N_6805);
and U7041 (N_7041,N_6931,N_6939);
nand U7042 (N_7042,N_6809,N_6928);
or U7043 (N_7043,N_6839,N_6953);
nor U7044 (N_7044,N_6910,N_6868);
nor U7045 (N_7045,N_6944,N_6826);
nand U7046 (N_7046,N_6907,N_6918);
and U7047 (N_7047,N_6821,N_6967);
nor U7048 (N_7048,N_6994,N_6876);
nand U7049 (N_7049,N_6987,N_6946);
nor U7050 (N_7050,N_6803,N_6848);
or U7051 (N_7051,N_6908,N_6916);
nand U7052 (N_7052,N_6937,N_6941);
and U7053 (N_7053,N_6828,N_6990);
nor U7054 (N_7054,N_6841,N_6812);
nand U7055 (N_7055,N_6802,N_6853);
or U7056 (N_7056,N_6927,N_6961);
nand U7057 (N_7057,N_6806,N_6930);
nor U7058 (N_7058,N_6871,N_6859);
and U7059 (N_7059,N_6829,N_6909);
nand U7060 (N_7060,N_6818,N_6950);
or U7061 (N_7061,N_6807,N_6952);
nor U7062 (N_7062,N_6879,N_6893);
and U7063 (N_7063,N_6823,N_6817);
or U7064 (N_7064,N_6949,N_6888);
or U7065 (N_7065,N_6991,N_6983);
nand U7066 (N_7066,N_6902,N_6951);
nor U7067 (N_7067,N_6849,N_6882);
nor U7068 (N_7068,N_6936,N_6880);
nor U7069 (N_7069,N_6995,N_6966);
nand U7070 (N_7070,N_6920,N_6974);
or U7071 (N_7071,N_6884,N_6962);
or U7072 (N_7072,N_6852,N_6904);
or U7073 (N_7073,N_6989,N_6947);
or U7074 (N_7074,N_6815,N_6847);
or U7075 (N_7075,N_6938,N_6874);
or U7076 (N_7076,N_6850,N_6968);
and U7077 (N_7077,N_6842,N_6897);
nand U7078 (N_7078,N_6804,N_6982);
xor U7079 (N_7079,N_6899,N_6800);
or U7080 (N_7080,N_6905,N_6891);
nor U7081 (N_7081,N_6834,N_6866);
and U7082 (N_7082,N_6811,N_6957);
xnor U7083 (N_7083,N_6872,N_6865);
nand U7084 (N_7084,N_6970,N_6972);
xor U7085 (N_7085,N_6985,N_6901);
nor U7086 (N_7086,N_6956,N_6863);
xor U7087 (N_7087,N_6877,N_6921);
nor U7088 (N_7088,N_6900,N_6895);
nand U7089 (N_7089,N_6854,N_6801);
nand U7090 (N_7090,N_6935,N_6999);
nor U7091 (N_7091,N_6861,N_6873);
or U7092 (N_7092,N_6979,N_6969);
and U7093 (N_7093,N_6914,N_6913);
nor U7094 (N_7094,N_6978,N_6892);
nor U7095 (N_7095,N_6926,N_6973);
or U7096 (N_7096,N_6992,N_6964);
nor U7097 (N_7097,N_6971,N_6997);
nand U7098 (N_7098,N_6832,N_6960);
xnor U7099 (N_7099,N_6840,N_6878);
nor U7100 (N_7100,N_6979,N_6829);
nor U7101 (N_7101,N_6918,N_6931);
or U7102 (N_7102,N_6867,N_6944);
nor U7103 (N_7103,N_6934,N_6994);
or U7104 (N_7104,N_6940,N_6835);
nor U7105 (N_7105,N_6931,N_6902);
and U7106 (N_7106,N_6899,N_6840);
nand U7107 (N_7107,N_6809,N_6810);
nand U7108 (N_7108,N_6843,N_6974);
nand U7109 (N_7109,N_6967,N_6918);
nor U7110 (N_7110,N_6857,N_6847);
nand U7111 (N_7111,N_6971,N_6946);
or U7112 (N_7112,N_6912,N_6922);
or U7113 (N_7113,N_6875,N_6921);
and U7114 (N_7114,N_6982,N_6908);
nand U7115 (N_7115,N_6914,N_6988);
nor U7116 (N_7116,N_6898,N_6918);
or U7117 (N_7117,N_6825,N_6940);
or U7118 (N_7118,N_6887,N_6946);
nand U7119 (N_7119,N_6885,N_6944);
nand U7120 (N_7120,N_6837,N_6941);
or U7121 (N_7121,N_6829,N_6848);
and U7122 (N_7122,N_6834,N_6868);
and U7123 (N_7123,N_6838,N_6940);
and U7124 (N_7124,N_6968,N_6911);
nor U7125 (N_7125,N_6895,N_6924);
nor U7126 (N_7126,N_6891,N_6851);
nand U7127 (N_7127,N_6822,N_6904);
xnor U7128 (N_7128,N_6896,N_6977);
nand U7129 (N_7129,N_6871,N_6989);
nor U7130 (N_7130,N_6931,N_6893);
and U7131 (N_7131,N_6872,N_6837);
nand U7132 (N_7132,N_6964,N_6894);
nand U7133 (N_7133,N_6815,N_6820);
xnor U7134 (N_7134,N_6842,N_6989);
nor U7135 (N_7135,N_6933,N_6894);
nand U7136 (N_7136,N_6866,N_6915);
nor U7137 (N_7137,N_6969,N_6941);
nand U7138 (N_7138,N_6881,N_6855);
or U7139 (N_7139,N_6936,N_6822);
or U7140 (N_7140,N_6873,N_6835);
nor U7141 (N_7141,N_6878,N_6958);
or U7142 (N_7142,N_6858,N_6947);
and U7143 (N_7143,N_6809,N_6891);
or U7144 (N_7144,N_6853,N_6900);
nand U7145 (N_7145,N_6905,N_6831);
or U7146 (N_7146,N_6992,N_6937);
nand U7147 (N_7147,N_6967,N_6800);
and U7148 (N_7148,N_6876,N_6953);
nand U7149 (N_7149,N_6936,N_6924);
nor U7150 (N_7150,N_6987,N_6805);
nor U7151 (N_7151,N_6824,N_6974);
and U7152 (N_7152,N_6963,N_6898);
nor U7153 (N_7153,N_6800,N_6900);
nand U7154 (N_7154,N_6971,N_6834);
and U7155 (N_7155,N_6908,N_6800);
and U7156 (N_7156,N_6994,N_6959);
and U7157 (N_7157,N_6912,N_6849);
or U7158 (N_7158,N_6956,N_6856);
and U7159 (N_7159,N_6957,N_6986);
xor U7160 (N_7160,N_6951,N_6868);
nor U7161 (N_7161,N_6877,N_6937);
or U7162 (N_7162,N_6824,N_6955);
or U7163 (N_7163,N_6904,N_6851);
and U7164 (N_7164,N_6842,N_6819);
and U7165 (N_7165,N_6920,N_6881);
xnor U7166 (N_7166,N_6879,N_6949);
xor U7167 (N_7167,N_6873,N_6952);
nand U7168 (N_7168,N_6997,N_6830);
or U7169 (N_7169,N_6898,N_6844);
and U7170 (N_7170,N_6988,N_6821);
or U7171 (N_7171,N_6839,N_6851);
nand U7172 (N_7172,N_6853,N_6959);
and U7173 (N_7173,N_6979,N_6935);
xnor U7174 (N_7174,N_6911,N_6905);
nand U7175 (N_7175,N_6846,N_6886);
and U7176 (N_7176,N_6982,N_6931);
nor U7177 (N_7177,N_6956,N_6995);
xor U7178 (N_7178,N_6914,N_6998);
nor U7179 (N_7179,N_6952,N_6975);
and U7180 (N_7180,N_6824,N_6985);
or U7181 (N_7181,N_6963,N_6939);
nand U7182 (N_7182,N_6872,N_6952);
and U7183 (N_7183,N_6906,N_6887);
nor U7184 (N_7184,N_6962,N_6829);
or U7185 (N_7185,N_6967,N_6923);
and U7186 (N_7186,N_6956,N_6991);
xor U7187 (N_7187,N_6802,N_6985);
nand U7188 (N_7188,N_6814,N_6910);
nor U7189 (N_7189,N_6959,N_6991);
nand U7190 (N_7190,N_6854,N_6996);
nor U7191 (N_7191,N_6930,N_6861);
or U7192 (N_7192,N_6828,N_6912);
nor U7193 (N_7193,N_6880,N_6883);
nor U7194 (N_7194,N_6811,N_6807);
and U7195 (N_7195,N_6953,N_6821);
nand U7196 (N_7196,N_6977,N_6902);
xnor U7197 (N_7197,N_6810,N_6845);
or U7198 (N_7198,N_6923,N_6837);
xor U7199 (N_7199,N_6924,N_6904);
nor U7200 (N_7200,N_7043,N_7035);
or U7201 (N_7201,N_7193,N_7109);
nor U7202 (N_7202,N_7128,N_7118);
nand U7203 (N_7203,N_7195,N_7047);
nand U7204 (N_7204,N_7105,N_7186);
or U7205 (N_7205,N_7031,N_7100);
and U7206 (N_7206,N_7165,N_7001);
xor U7207 (N_7207,N_7170,N_7082);
nor U7208 (N_7208,N_7180,N_7168);
and U7209 (N_7209,N_7067,N_7086);
or U7210 (N_7210,N_7009,N_7179);
nor U7211 (N_7211,N_7192,N_7199);
nor U7212 (N_7212,N_7171,N_7185);
nand U7213 (N_7213,N_7169,N_7056);
and U7214 (N_7214,N_7046,N_7142);
nor U7215 (N_7215,N_7116,N_7120);
nand U7216 (N_7216,N_7164,N_7194);
and U7217 (N_7217,N_7074,N_7093);
nor U7218 (N_7218,N_7097,N_7041);
and U7219 (N_7219,N_7136,N_7045);
and U7220 (N_7220,N_7071,N_7076);
and U7221 (N_7221,N_7022,N_7190);
and U7222 (N_7222,N_7036,N_7068);
or U7223 (N_7223,N_7040,N_7049);
or U7224 (N_7224,N_7063,N_7054);
and U7225 (N_7225,N_7052,N_7042);
or U7226 (N_7226,N_7184,N_7182);
nor U7227 (N_7227,N_7038,N_7122);
nand U7228 (N_7228,N_7079,N_7134);
nand U7229 (N_7229,N_7030,N_7197);
nor U7230 (N_7230,N_7150,N_7015);
and U7231 (N_7231,N_7191,N_7154);
xor U7232 (N_7232,N_7181,N_7152);
nor U7233 (N_7233,N_7085,N_7080);
and U7234 (N_7234,N_7138,N_7053);
nand U7235 (N_7235,N_7060,N_7000);
or U7236 (N_7236,N_7126,N_7070);
or U7237 (N_7237,N_7127,N_7177);
or U7238 (N_7238,N_7010,N_7011);
xnor U7239 (N_7239,N_7081,N_7024);
or U7240 (N_7240,N_7119,N_7123);
nor U7241 (N_7241,N_7151,N_7161);
nand U7242 (N_7242,N_7131,N_7007);
nor U7243 (N_7243,N_7026,N_7187);
nor U7244 (N_7244,N_7029,N_7106);
nor U7245 (N_7245,N_7178,N_7196);
or U7246 (N_7246,N_7146,N_7003);
and U7247 (N_7247,N_7064,N_7088);
xnor U7248 (N_7248,N_7176,N_7017);
nor U7249 (N_7249,N_7174,N_7143);
or U7250 (N_7250,N_7034,N_7175);
or U7251 (N_7251,N_7103,N_7008);
xor U7252 (N_7252,N_7051,N_7173);
nand U7253 (N_7253,N_7005,N_7061);
xor U7254 (N_7254,N_7065,N_7188);
and U7255 (N_7255,N_7050,N_7075);
nor U7256 (N_7256,N_7133,N_7004);
nor U7257 (N_7257,N_7167,N_7083);
xnor U7258 (N_7258,N_7139,N_7018);
nand U7259 (N_7259,N_7077,N_7025);
nor U7260 (N_7260,N_7058,N_7140);
and U7261 (N_7261,N_7013,N_7019);
nand U7262 (N_7262,N_7002,N_7091);
nand U7263 (N_7263,N_7166,N_7145);
nand U7264 (N_7264,N_7147,N_7027);
and U7265 (N_7265,N_7048,N_7033);
or U7266 (N_7266,N_7084,N_7144);
and U7267 (N_7267,N_7012,N_7117);
nor U7268 (N_7268,N_7078,N_7098);
nor U7269 (N_7269,N_7072,N_7066);
nand U7270 (N_7270,N_7155,N_7156);
or U7271 (N_7271,N_7102,N_7153);
nand U7272 (N_7272,N_7062,N_7044);
nand U7273 (N_7273,N_7069,N_7157);
and U7274 (N_7274,N_7130,N_7039);
nand U7275 (N_7275,N_7087,N_7028);
nand U7276 (N_7276,N_7014,N_7089);
nor U7277 (N_7277,N_7104,N_7137);
nand U7278 (N_7278,N_7073,N_7095);
nor U7279 (N_7279,N_7162,N_7032);
nor U7280 (N_7280,N_7108,N_7158);
nand U7281 (N_7281,N_7124,N_7135);
nand U7282 (N_7282,N_7037,N_7059);
nor U7283 (N_7283,N_7163,N_7183);
and U7284 (N_7284,N_7114,N_7148);
and U7285 (N_7285,N_7094,N_7113);
and U7286 (N_7286,N_7112,N_7121);
nor U7287 (N_7287,N_7016,N_7129);
and U7288 (N_7288,N_7189,N_7159);
and U7289 (N_7289,N_7132,N_7107);
nor U7290 (N_7290,N_7149,N_7006);
nor U7291 (N_7291,N_7110,N_7090);
nand U7292 (N_7292,N_7096,N_7020);
and U7293 (N_7293,N_7092,N_7115);
nand U7294 (N_7294,N_7172,N_7111);
xor U7295 (N_7295,N_7055,N_7101);
and U7296 (N_7296,N_7021,N_7057);
and U7297 (N_7297,N_7160,N_7023);
or U7298 (N_7298,N_7141,N_7099);
nor U7299 (N_7299,N_7198,N_7125);
xnor U7300 (N_7300,N_7113,N_7030);
nor U7301 (N_7301,N_7154,N_7075);
nor U7302 (N_7302,N_7122,N_7132);
nand U7303 (N_7303,N_7107,N_7044);
nor U7304 (N_7304,N_7184,N_7000);
nand U7305 (N_7305,N_7059,N_7119);
and U7306 (N_7306,N_7099,N_7162);
and U7307 (N_7307,N_7140,N_7093);
nand U7308 (N_7308,N_7066,N_7019);
xor U7309 (N_7309,N_7132,N_7100);
and U7310 (N_7310,N_7083,N_7041);
and U7311 (N_7311,N_7011,N_7001);
or U7312 (N_7312,N_7196,N_7148);
nor U7313 (N_7313,N_7021,N_7074);
nor U7314 (N_7314,N_7100,N_7098);
nand U7315 (N_7315,N_7006,N_7017);
and U7316 (N_7316,N_7185,N_7112);
and U7317 (N_7317,N_7135,N_7060);
or U7318 (N_7318,N_7037,N_7190);
or U7319 (N_7319,N_7005,N_7043);
and U7320 (N_7320,N_7126,N_7061);
and U7321 (N_7321,N_7137,N_7036);
and U7322 (N_7322,N_7098,N_7075);
and U7323 (N_7323,N_7148,N_7087);
nand U7324 (N_7324,N_7139,N_7014);
nand U7325 (N_7325,N_7185,N_7113);
and U7326 (N_7326,N_7097,N_7095);
nor U7327 (N_7327,N_7143,N_7121);
nand U7328 (N_7328,N_7182,N_7007);
or U7329 (N_7329,N_7187,N_7142);
and U7330 (N_7330,N_7122,N_7090);
xor U7331 (N_7331,N_7114,N_7034);
nand U7332 (N_7332,N_7087,N_7076);
nor U7333 (N_7333,N_7165,N_7109);
and U7334 (N_7334,N_7072,N_7193);
or U7335 (N_7335,N_7007,N_7141);
nand U7336 (N_7336,N_7011,N_7000);
nand U7337 (N_7337,N_7140,N_7114);
and U7338 (N_7338,N_7056,N_7011);
or U7339 (N_7339,N_7014,N_7078);
and U7340 (N_7340,N_7162,N_7186);
xnor U7341 (N_7341,N_7191,N_7029);
and U7342 (N_7342,N_7116,N_7036);
nor U7343 (N_7343,N_7171,N_7108);
nor U7344 (N_7344,N_7095,N_7063);
nor U7345 (N_7345,N_7185,N_7089);
nand U7346 (N_7346,N_7112,N_7198);
nor U7347 (N_7347,N_7132,N_7182);
and U7348 (N_7348,N_7004,N_7096);
nand U7349 (N_7349,N_7069,N_7058);
xnor U7350 (N_7350,N_7135,N_7092);
nand U7351 (N_7351,N_7131,N_7125);
nor U7352 (N_7352,N_7183,N_7035);
or U7353 (N_7353,N_7029,N_7149);
xnor U7354 (N_7354,N_7023,N_7192);
nand U7355 (N_7355,N_7013,N_7192);
or U7356 (N_7356,N_7065,N_7035);
nand U7357 (N_7357,N_7114,N_7195);
and U7358 (N_7358,N_7061,N_7130);
nand U7359 (N_7359,N_7143,N_7193);
nor U7360 (N_7360,N_7137,N_7017);
nor U7361 (N_7361,N_7047,N_7032);
nand U7362 (N_7362,N_7097,N_7152);
nor U7363 (N_7363,N_7097,N_7139);
and U7364 (N_7364,N_7008,N_7042);
or U7365 (N_7365,N_7039,N_7167);
nand U7366 (N_7366,N_7155,N_7137);
or U7367 (N_7367,N_7181,N_7179);
and U7368 (N_7368,N_7075,N_7028);
and U7369 (N_7369,N_7011,N_7082);
nor U7370 (N_7370,N_7097,N_7054);
nand U7371 (N_7371,N_7128,N_7022);
and U7372 (N_7372,N_7186,N_7074);
nor U7373 (N_7373,N_7159,N_7135);
and U7374 (N_7374,N_7155,N_7039);
nor U7375 (N_7375,N_7087,N_7061);
or U7376 (N_7376,N_7028,N_7055);
and U7377 (N_7377,N_7010,N_7005);
or U7378 (N_7378,N_7138,N_7147);
xnor U7379 (N_7379,N_7117,N_7070);
xnor U7380 (N_7380,N_7087,N_7151);
xor U7381 (N_7381,N_7104,N_7154);
or U7382 (N_7382,N_7178,N_7012);
and U7383 (N_7383,N_7020,N_7192);
and U7384 (N_7384,N_7042,N_7088);
or U7385 (N_7385,N_7199,N_7097);
or U7386 (N_7386,N_7093,N_7032);
and U7387 (N_7387,N_7080,N_7170);
or U7388 (N_7388,N_7120,N_7024);
xor U7389 (N_7389,N_7001,N_7035);
or U7390 (N_7390,N_7038,N_7138);
nor U7391 (N_7391,N_7142,N_7117);
and U7392 (N_7392,N_7057,N_7020);
nor U7393 (N_7393,N_7066,N_7183);
nand U7394 (N_7394,N_7002,N_7079);
xnor U7395 (N_7395,N_7152,N_7040);
or U7396 (N_7396,N_7156,N_7172);
nand U7397 (N_7397,N_7011,N_7089);
nor U7398 (N_7398,N_7139,N_7123);
or U7399 (N_7399,N_7159,N_7037);
nor U7400 (N_7400,N_7305,N_7276);
nor U7401 (N_7401,N_7274,N_7245);
and U7402 (N_7402,N_7353,N_7323);
nor U7403 (N_7403,N_7375,N_7285);
nor U7404 (N_7404,N_7265,N_7352);
nand U7405 (N_7405,N_7271,N_7381);
and U7406 (N_7406,N_7289,N_7288);
nor U7407 (N_7407,N_7244,N_7368);
and U7408 (N_7408,N_7234,N_7361);
nand U7409 (N_7409,N_7248,N_7383);
and U7410 (N_7410,N_7241,N_7255);
and U7411 (N_7411,N_7397,N_7219);
nor U7412 (N_7412,N_7238,N_7229);
nor U7413 (N_7413,N_7284,N_7396);
or U7414 (N_7414,N_7232,N_7363);
or U7415 (N_7415,N_7299,N_7348);
nor U7416 (N_7416,N_7332,N_7318);
nor U7417 (N_7417,N_7279,N_7200);
and U7418 (N_7418,N_7385,N_7326);
or U7419 (N_7419,N_7358,N_7384);
and U7420 (N_7420,N_7317,N_7399);
and U7421 (N_7421,N_7391,N_7224);
and U7422 (N_7422,N_7217,N_7294);
nand U7423 (N_7423,N_7307,N_7344);
and U7424 (N_7424,N_7388,N_7321);
and U7425 (N_7425,N_7333,N_7273);
and U7426 (N_7426,N_7339,N_7372);
nor U7427 (N_7427,N_7367,N_7283);
nand U7428 (N_7428,N_7356,N_7242);
and U7429 (N_7429,N_7312,N_7338);
and U7430 (N_7430,N_7309,N_7330);
or U7431 (N_7431,N_7233,N_7205);
and U7432 (N_7432,N_7331,N_7300);
xnor U7433 (N_7433,N_7237,N_7291);
nor U7434 (N_7434,N_7239,N_7351);
xor U7435 (N_7435,N_7313,N_7393);
and U7436 (N_7436,N_7267,N_7389);
nand U7437 (N_7437,N_7208,N_7382);
or U7438 (N_7438,N_7262,N_7207);
and U7439 (N_7439,N_7350,N_7204);
or U7440 (N_7440,N_7357,N_7322);
or U7441 (N_7441,N_7297,N_7249);
or U7442 (N_7442,N_7336,N_7302);
and U7443 (N_7443,N_7310,N_7226);
and U7444 (N_7444,N_7280,N_7227);
and U7445 (N_7445,N_7345,N_7213);
nand U7446 (N_7446,N_7268,N_7210);
nand U7447 (N_7447,N_7216,N_7370);
nand U7448 (N_7448,N_7214,N_7369);
and U7449 (N_7449,N_7236,N_7371);
and U7450 (N_7450,N_7247,N_7264);
and U7451 (N_7451,N_7304,N_7290);
nor U7452 (N_7452,N_7266,N_7292);
nor U7453 (N_7453,N_7203,N_7228);
nor U7454 (N_7454,N_7215,N_7329);
nor U7455 (N_7455,N_7254,N_7364);
nor U7456 (N_7456,N_7298,N_7324);
nor U7457 (N_7457,N_7281,N_7235);
or U7458 (N_7458,N_7306,N_7287);
and U7459 (N_7459,N_7296,N_7340);
or U7460 (N_7460,N_7349,N_7392);
or U7461 (N_7461,N_7209,N_7377);
nor U7462 (N_7462,N_7301,N_7202);
nor U7463 (N_7463,N_7355,N_7359);
nand U7464 (N_7464,N_7251,N_7286);
nand U7465 (N_7465,N_7257,N_7293);
nand U7466 (N_7466,N_7374,N_7394);
xnor U7467 (N_7467,N_7246,N_7218);
and U7468 (N_7468,N_7354,N_7320);
nor U7469 (N_7469,N_7315,N_7337);
or U7470 (N_7470,N_7259,N_7201);
nand U7471 (N_7471,N_7252,N_7362);
nor U7472 (N_7472,N_7282,N_7230);
nand U7473 (N_7473,N_7316,N_7319);
or U7474 (N_7474,N_7387,N_7328);
or U7475 (N_7475,N_7256,N_7211);
nor U7476 (N_7476,N_7272,N_7221);
or U7477 (N_7477,N_7376,N_7366);
nor U7478 (N_7478,N_7334,N_7303);
nand U7479 (N_7479,N_7258,N_7222);
and U7480 (N_7480,N_7390,N_7261);
nor U7481 (N_7481,N_7223,N_7263);
or U7482 (N_7482,N_7325,N_7269);
or U7483 (N_7483,N_7379,N_7335);
or U7484 (N_7484,N_7342,N_7277);
nand U7485 (N_7485,N_7378,N_7278);
or U7486 (N_7486,N_7212,N_7295);
nand U7487 (N_7487,N_7341,N_7243);
and U7488 (N_7488,N_7206,N_7395);
and U7489 (N_7489,N_7253,N_7220);
nand U7490 (N_7490,N_7347,N_7386);
and U7491 (N_7491,N_7231,N_7365);
nor U7492 (N_7492,N_7398,N_7260);
or U7493 (N_7493,N_7225,N_7360);
nor U7494 (N_7494,N_7327,N_7314);
nor U7495 (N_7495,N_7270,N_7373);
or U7496 (N_7496,N_7311,N_7308);
and U7497 (N_7497,N_7346,N_7275);
nor U7498 (N_7498,N_7250,N_7380);
or U7499 (N_7499,N_7240,N_7343);
xor U7500 (N_7500,N_7364,N_7380);
nor U7501 (N_7501,N_7288,N_7247);
nor U7502 (N_7502,N_7200,N_7314);
or U7503 (N_7503,N_7294,N_7302);
nor U7504 (N_7504,N_7382,N_7202);
or U7505 (N_7505,N_7304,N_7258);
nand U7506 (N_7506,N_7322,N_7392);
and U7507 (N_7507,N_7305,N_7345);
nand U7508 (N_7508,N_7298,N_7343);
nor U7509 (N_7509,N_7391,N_7346);
and U7510 (N_7510,N_7294,N_7224);
or U7511 (N_7511,N_7248,N_7317);
nand U7512 (N_7512,N_7202,N_7390);
nor U7513 (N_7513,N_7367,N_7254);
nand U7514 (N_7514,N_7373,N_7242);
nand U7515 (N_7515,N_7320,N_7349);
and U7516 (N_7516,N_7331,N_7377);
nand U7517 (N_7517,N_7272,N_7260);
xnor U7518 (N_7518,N_7342,N_7240);
or U7519 (N_7519,N_7341,N_7266);
or U7520 (N_7520,N_7262,N_7215);
nor U7521 (N_7521,N_7252,N_7388);
or U7522 (N_7522,N_7344,N_7328);
and U7523 (N_7523,N_7337,N_7256);
nand U7524 (N_7524,N_7306,N_7332);
nor U7525 (N_7525,N_7328,N_7295);
or U7526 (N_7526,N_7205,N_7332);
nor U7527 (N_7527,N_7369,N_7295);
or U7528 (N_7528,N_7307,N_7350);
nor U7529 (N_7529,N_7207,N_7257);
or U7530 (N_7530,N_7282,N_7258);
and U7531 (N_7531,N_7370,N_7371);
or U7532 (N_7532,N_7365,N_7271);
nor U7533 (N_7533,N_7321,N_7375);
or U7534 (N_7534,N_7310,N_7368);
nand U7535 (N_7535,N_7253,N_7202);
and U7536 (N_7536,N_7204,N_7245);
or U7537 (N_7537,N_7273,N_7222);
and U7538 (N_7538,N_7200,N_7357);
or U7539 (N_7539,N_7332,N_7322);
nand U7540 (N_7540,N_7297,N_7281);
nor U7541 (N_7541,N_7352,N_7270);
nand U7542 (N_7542,N_7325,N_7387);
or U7543 (N_7543,N_7267,N_7329);
nand U7544 (N_7544,N_7377,N_7295);
or U7545 (N_7545,N_7260,N_7251);
nand U7546 (N_7546,N_7200,N_7374);
or U7547 (N_7547,N_7292,N_7201);
or U7548 (N_7548,N_7307,N_7326);
or U7549 (N_7549,N_7344,N_7382);
nor U7550 (N_7550,N_7279,N_7385);
and U7551 (N_7551,N_7306,N_7220);
or U7552 (N_7552,N_7293,N_7376);
or U7553 (N_7553,N_7275,N_7234);
nor U7554 (N_7554,N_7222,N_7387);
nand U7555 (N_7555,N_7327,N_7345);
or U7556 (N_7556,N_7237,N_7295);
and U7557 (N_7557,N_7269,N_7263);
nor U7558 (N_7558,N_7253,N_7306);
or U7559 (N_7559,N_7286,N_7370);
xor U7560 (N_7560,N_7220,N_7344);
nand U7561 (N_7561,N_7290,N_7255);
nand U7562 (N_7562,N_7247,N_7244);
nand U7563 (N_7563,N_7272,N_7376);
nand U7564 (N_7564,N_7333,N_7308);
or U7565 (N_7565,N_7348,N_7362);
nand U7566 (N_7566,N_7338,N_7371);
and U7567 (N_7567,N_7347,N_7288);
or U7568 (N_7568,N_7280,N_7208);
nand U7569 (N_7569,N_7269,N_7306);
nand U7570 (N_7570,N_7344,N_7265);
nor U7571 (N_7571,N_7252,N_7396);
or U7572 (N_7572,N_7283,N_7265);
nand U7573 (N_7573,N_7355,N_7361);
nor U7574 (N_7574,N_7321,N_7259);
or U7575 (N_7575,N_7258,N_7329);
nand U7576 (N_7576,N_7293,N_7299);
xor U7577 (N_7577,N_7258,N_7390);
nand U7578 (N_7578,N_7290,N_7318);
and U7579 (N_7579,N_7270,N_7320);
nor U7580 (N_7580,N_7238,N_7370);
nand U7581 (N_7581,N_7395,N_7385);
nor U7582 (N_7582,N_7364,N_7289);
and U7583 (N_7583,N_7254,N_7260);
nor U7584 (N_7584,N_7375,N_7359);
and U7585 (N_7585,N_7269,N_7232);
and U7586 (N_7586,N_7287,N_7383);
xnor U7587 (N_7587,N_7334,N_7371);
and U7588 (N_7588,N_7323,N_7282);
nor U7589 (N_7589,N_7206,N_7356);
and U7590 (N_7590,N_7311,N_7338);
xor U7591 (N_7591,N_7276,N_7248);
nor U7592 (N_7592,N_7281,N_7363);
nand U7593 (N_7593,N_7363,N_7263);
and U7594 (N_7594,N_7352,N_7375);
and U7595 (N_7595,N_7385,N_7334);
xor U7596 (N_7596,N_7388,N_7265);
or U7597 (N_7597,N_7322,N_7372);
and U7598 (N_7598,N_7304,N_7278);
or U7599 (N_7599,N_7243,N_7214);
nor U7600 (N_7600,N_7452,N_7417);
nor U7601 (N_7601,N_7491,N_7431);
and U7602 (N_7602,N_7406,N_7411);
xor U7603 (N_7603,N_7530,N_7418);
nand U7604 (N_7604,N_7472,N_7589);
nor U7605 (N_7605,N_7427,N_7544);
nor U7606 (N_7606,N_7576,N_7451);
nor U7607 (N_7607,N_7499,N_7410);
nor U7608 (N_7608,N_7578,N_7446);
or U7609 (N_7609,N_7554,N_7400);
nand U7610 (N_7610,N_7414,N_7560);
or U7611 (N_7611,N_7433,N_7456);
nor U7612 (N_7612,N_7517,N_7422);
and U7613 (N_7613,N_7445,N_7520);
nor U7614 (N_7614,N_7466,N_7421);
nand U7615 (N_7615,N_7425,N_7535);
nor U7616 (N_7616,N_7519,N_7592);
xnor U7617 (N_7617,N_7436,N_7481);
nand U7618 (N_7618,N_7573,N_7563);
xor U7619 (N_7619,N_7542,N_7586);
nand U7620 (N_7620,N_7454,N_7462);
and U7621 (N_7621,N_7553,N_7523);
nor U7622 (N_7622,N_7558,N_7477);
xor U7623 (N_7623,N_7416,N_7412);
or U7624 (N_7624,N_7478,N_7450);
nor U7625 (N_7625,N_7470,N_7532);
nand U7626 (N_7626,N_7401,N_7480);
and U7627 (N_7627,N_7583,N_7531);
or U7628 (N_7628,N_7504,N_7484);
or U7629 (N_7629,N_7522,N_7571);
nor U7630 (N_7630,N_7419,N_7404);
nor U7631 (N_7631,N_7430,N_7424);
and U7632 (N_7632,N_7496,N_7533);
or U7633 (N_7633,N_7493,N_7527);
or U7634 (N_7634,N_7489,N_7521);
nor U7635 (N_7635,N_7525,N_7540);
nand U7636 (N_7636,N_7529,N_7460);
nor U7637 (N_7637,N_7465,N_7565);
or U7638 (N_7638,N_7428,N_7468);
or U7639 (N_7639,N_7413,N_7584);
or U7640 (N_7640,N_7596,N_7434);
or U7641 (N_7641,N_7572,N_7511);
or U7642 (N_7642,N_7500,N_7463);
or U7643 (N_7643,N_7409,N_7442);
or U7644 (N_7644,N_7551,N_7464);
nand U7645 (N_7645,N_7420,N_7506);
xnor U7646 (N_7646,N_7547,N_7469);
nand U7647 (N_7647,N_7582,N_7495);
nand U7648 (N_7648,N_7486,N_7588);
nor U7649 (N_7649,N_7497,N_7549);
and U7650 (N_7650,N_7515,N_7444);
or U7651 (N_7651,N_7552,N_7440);
or U7652 (N_7652,N_7429,N_7524);
nor U7653 (N_7653,N_7514,N_7590);
nor U7654 (N_7654,N_7453,N_7402);
and U7655 (N_7655,N_7562,N_7426);
or U7656 (N_7656,N_7455,N_7479);
or U7657 (N_7657,N_7593,N_7577);
and U7658 (N_7658,N_7567,N_7503);
and U7659 (N_7659,N_7541,N_7403);
nor U7660 (N_7660,N_7585,N_7534);
and U7661 (N_7661,N_7490,N_7518);
and U7662 (N_7662,N_7494,N_7483);
or U7663 (N_7663,N_7556,N_7509);
nand U7664 (N_7664,N_7580,N_7437);
or U7665 (N_7665,N_7512,N_7568);
xnor U7666 (N_7666,N_7447,N_7536);
nor U7667 (N_7667,N_7435,N_7594);
or U7668 (N_7668,N_7538,N_7459);
xnor U7669 (N_7669,N_7505,N_7581);
or U7670 (N_7670,N_7569,N_7439);
xor U7671 (N_7671,N_7566,N_7432);
and U7672 (N_7672,N_7526,N_7548);
nor U7673 (N_7673,N_7510,N_7407);
or U7674 (N_7674,N_7579,N_7543);
and U7675 (N_7675,N_7570,N_7476);
xnor U7676 (N_7676,N_7492,N_7598);
nand U7677 (N_7677,N_7539,N_7513);
nand U7678 (N_7678,N_7471,N_7443);
or U7679 (N_7679,N_7415,N_7423);
nand U7680 (N_7680,N_7474,N_7561);
nor U7681 (N_7681,N_7595,N_7597);
xnor U7682 (N_7682,N_7537,N_7559);
and U7683 (N_7683,N_7485,N_7575);
nor U7684 (N_7684,N_7449,N_7557);
and U7685 (N_7685,N_7488,N_7508);
and U7686 (N_7686,N_7564,N_7528);
and U7687 (N_7687,N_7507,N_7587);
nor U7688 (N_7688,N_7555,N_7457);
nor U7689 (N_7689,N_7501,N_7405);
xnor U7690 (N_7690,N_7448,N_7498);
and U7691 (N_7691,N_7574,N_7467);
or U7692 (N_7692,N_7458,N_7482);
nor U7693 (N_7693,N_7473,N_7408);
and U7694 (N_7694,N_7502,N_7475);
nor U7695 (N_7695,N_7591,N_7441);
nor U7696 (N_7696,N_7461,N_7516);
nor U7697 (N_7697,N_7550,N_7438);
nor U7698 (N_7698,N_7545,N_7487);
or U7699 (N_7699,N_7599,N_7546);
or U7700 (N_7700,N_7402,N_7529);
nor U7701 (N_7701,N_7440,N_7595);
nor U7702 (N_7702,N_7444,N_7544);
nor U7703 (N_7703,N_7492,N_7544);
and U7704 (N_7704,N_7567,N_7437);
and U7705 (N_7705,N_7522,N_7433);
and U7706 (N_7706,N_7459,N_7490);
nand U7707 (N_7707,N_7509,N_7521);
xor U7708 (N_7708,N_7449,N_7561);
nand U7709 (N_7709,N_7418,N_7493);
and U7710 (N_7710,N_7527,N_7453);
and U7711 (N_7711,N_7434,N_7565);
xor U7712 (N_7712,N_7421,N_7519);
or U7713 (N_7713,N_7483,N_7486);
nand U7714 (N_7714,N_7419,N_7534);
and U7715 (N_7715,N_7423,N_7545);
or U7716 (N_7716,N_7534,N_7434);
nor U7717 (N_7717,N_7561,N_7542);
or U7718 (N_7718,N_7434,N_7535);
nand U7719 (N_7719,N_7483,N_7487);
or U7720 (N_7720,N_7569,N_7405);
nor U7721 (N_7721,N_7492,N_7417);
nor U7722 (N_7722,N_7551,N_7514);
nor U7723 (N_7723,N_7514,N_7548);
xor U7724 (N_7724,N_7442,N_7572);
or U7725 (N_7725,N_7462,N_7544);
nor U7726 (N_7726,N_7493,N_7503);
and U7727 (N_7727,N_7481,N_7521);
nor U7728 (N_7728,N_7554,N_7446);
or U7729 (N_7729,N_7523,N_7486);
nand U7730 (N_7730,N_7432,N_7550);
and U7731 (N_7731,N_7428,N_7536);
or U7732 (N_7732,N_7450,N_7452);
or U7733 (N_7733,N_7590,N_7567);
or U7734 (N_7734,N_7478,N_7582);
nand U7735 (N_7735,N_7489,N_7556);
xnor U7736 (N_7736,N_7558,N_7456);
or U7737 (N_7737,N_7449,N_7545);
or U7738 (N_7738,N_7478,N_7579);
and U7739 (N_7739,N_7436,N_7430);
or U7740 (N_7740,N_7446,N_7510);
nor U7741 (N_7741,N_7509,N_7512);
xor U7742 (N_7742,N_7436,N_7416);
or U7743 (N_7743,N_7448,N_7433);
and U7744 (N_7744,N_7458,N_7512);
nor U7745 (N_7745,N_7457,N_7585);
xnor U7746 (N_7746,N_7421,N_7443);
and U7747 (N_7747,N_7463,N_7587);
nor U7748 (N_7748,N_7576,N_7592);
nand U7749 (N_7749,N_7413,N_7470);
or U7750 (N_7750,N_7414,N_7554);
or U7751 (N_7751,N_7584,N_7432);
or U7752 (N_7752,N_7565,N_7559);
nor U7753 (N_7753,N_7462,N_7450);
xor U7754 (N_7754,N_7402,N_7507);
nand U7755 (N_7755,N_7439,N_7436);
or U7756 (N_7756,N_7464,N_7402);
and U7757 (N_7757,N_7445,N_7459);
and U7758 (N_7758,N_7445,N_7406);
or U7759 (N_7759,N_7553,N_7425);
nor U7760 (N_7760,N_7515,N_7534);
and U7761 (N_7761,N_7496,N_7514);
and U7762 (N_7762,N_7524,N_7513);
or U7763 (N_7763,N_7483,N_7404);
or U7764 (N_7764,N_7582,N_7450);
or U7765 (N_7765,N_7590,N_7509);
nand U7766 (N_7766,N_7410,N_7405);
nand U7767 (N_7767,N_7450,N_7451);
nand U7768 (N_7768,N_7452,N_7583);
xnor U7769 (N_7769,N_7531,N_7410);
and U7770 (N_7770,N_7552,N_7507);
or U7771 (N_7771,N_7476,N_7443);
or U7772 (N_7772,N_7565,N_7501);
nor U7773 (N_7773,N_7475,N_7575);
xnor U7774 (N_7774,N_7578,N_7463);
nand U7775 (N_7775,N_7482,N_7574);
and U7776 (N_7776,N_7512,N_7429);
nand U7777 (N_7777,N_7462,N_7482);
and U7778 (N_7778,N_7483,N_7477);
or U7779 (N_7779,N_7425,N_7492);
xnor U7780 (N_7780,N_7515,N_7483);
or U7781 (N_7781,N_7490,N_7592);
or U7782 (N_7782,N_7562,N_7542);
nor U7783 (N_7783,N_7455,N_7450);
or U7784 (N_7784,N_7556,N_7498);
nor U7785 (N_7785,N_7487,N_7574);
nor U7786 (N_7786,N_7466,N_7468);
and U7787 (N_7787,N_7575,N_7599);
and U7788 (N_7788,N_7491,N_7560);
nor U7789 (N_7789,N_7402,N_7553);
xor U7790 (N_7790,N_7440,N_7467);
nor U7791 (N_7791,N_7520,N_7461);
and U7792 (N_7792,N_7448,N_7559);
xor U7793 (N_7793,N_7549,N_7595);
and U7794 (N_7794,N_7587,N_7479);
xnor U7795 (N_7795,N_7441,N_7404);
or U7796 (N_7796,N_7524,N_7517);
nor U7797 (N_7797,N_7429,N_7411);
xnor U7798 (N_7798,N_7442,N_7447);
nand U7799 (N_7799,N_7546,N_7436);
nor U7800 (N_7800,N_7787,N_7602);
and U7801 (N_7801,N_7664,N_7781);
or U7802 (N_7802,N_7732,N_7667);
nor U7803 (N_7803,N_7624,N_7691);
nand U7804 (N_7804,N_7701,N_7611);
and U7805 (N_7805,N_7789,N_7690);
nor U7806 (N_7806,N_7673,N_7730);
nor U7807 (N_7807,N_7772,N_7604);
nor U7808 (N_7808,N_7608,N_7776);
or U7809 (N_7809,N_7709,N_7767);
nor U7810 (N_7810,N_7766,N_7731);
or U7811 (N_7811,N_7606,N_7754);
or U7812 (N_7812,N_7721,N_7738);
nor U7813 (N_7813,N_7600,N_7728);
nand U7814 (N_7814,N_7746,N_7764);
and U7815 (N_7815,N_7720,N_7677);
nand U7816 (N_7816,N_7739,N_7693);
nor U7817 (N_7817,N_7678,N_7637);
or U7818 (N_7818,N_7626,N_7745);
nor U7819 (N_7819,N_7650,N_7785);
nor U7820 (N_7820,N_7669,N_7618);
nor U7821 (N_7821,N_7685,N_7699);
and U7822 (N_7822,N_7651,N_7694);
and U7823 (N_7823,N_7758,N_7793);
xnor U7824 (N_7824,N_7647,N_7706);
or U7825 (N_7825,N_7768,N_7703);
and U7826 (N_7826,N_7770,N_7665);
nor U7827 (N_7827,N_7695,N_7794);
nor U7828 (N_7828,N_7753,N_7773);
xor U7829 (N_7829,N_7654,N_7620);
and U7830 (N_7830,N_7632,N_7716);
nor U7831 (N_7831,N_7700,N_7751);
and U7832 (N_7832,N_7779,N_7780);
or U7833 (N_7833,N_7771,N_7712);
nand U7834 (N_7834,N_7639,N_7658);
and U7835 (N_7835,N_7653,N_7672);
xor U7836 (N_7836,N_7718,N_7666);
and U7837 (N_7837,N_7715,N_7765);
nor U7838 (N_7838,N_7757,N_7601);
nand U7839 (N_7839,N_7617,N_7725);
or U7840 (N_7840,N_7630,N_7625);
and U7841 (N_7841,N_7675,N_7670);
nand U7842 (N_7842,N_7643,N_7762);
nand U7843 (N_7843,N_7777,N_7747);
nand U7844 (N_7844,N_7641,N_7613);
nand U7845 (N_7845,N_7697,N_7682);
nor U7846 (N_7846,N_7760,N_7644);
nor U7847 (N_7847,N_7656,N_7707);
or U7848 (N_7848,N_7657,N_7610);
nand U7849 (N_7849,N_7796,N_7623);
or U7850 (N_7850,N_7742,N_7688);
and U7851 (N_7851,N_7714,N_7756);
and U7852 (N_7852,N_7784,N_7717);
nand U7853 (N_7853,N_7755,N_7638);
xnor U7854 (N_7854,N_7722,N_7680);
nor U7855 (N_7855,N_7659,N_7681);
nand U7856 (N_7856,N_7790,N_7686);
nand U7857 (N_7857,N_7615,N_7634);
nor U7858 (N_7858,N_7652,N_7735);
nor U7859 (N_7859,N_7698,N_7621);
or U7860 (N_7860,N_7786,N_7734);
nand U7861 (N_7861,N_7729,N_7640);
and U7862 (N_7862,N_7727,N_7740);
or U7863 (N_7863,N_7628,N_7798);
nor U7864 (N_7864,N_7689,N_7795);
and U7865 (N_7865,N_7614,N_7710);
nor U7866 (N_7866,N_7679,N_7629);
nor U7867 (N_7867,N_7791,N_7605);
nor U7868 (N_7868,N_7645,N_7642);
nand U7869 (N_7869,N_7799,N_7743);
nand U7870 (N_7870,N_7661,N_7708);
nand U7871 (N_7871,N_7683,N_7671);
nand U7872 (N_7872,N_7633,N_7763);
or U7873 (N_7873,N_7692,N_7687);
nand U7874 (N_7874,N_7646,N_7631);
or U7875 (N_7875,N_7724,N_7748);
nor U7876 (N_7876,N_7744,N_7775);
and U7877 (N_7877,N_7736,N_7603);
and U7878 (N_7878,N_7696,N_7711);
nor U7879 (N_7879,N_7663,N_7733);
nor U7880 (N_7880,N_7719,N_7741);
nand U7881 (N_7881,N_7797,N_7778);
and U7882 (N_7882,N_7660,N_7627);
nor U7883 (N_7883,N_7702,N_7609);
and U7884 (N_7884,N_7668,N_7761);
or U7885 (N_7885,N_7749,N_7713);
nand U7886 (N_7886,N_7792,N_7649);
nor U7887 (N_7887,N_7636,N_7684);
xor U7888 (N_7888,N_7655,N_7674);
nor U7889 (N_7889,N_7750,N_7676);
or U7890 (N_7890,N_7704,N_7616);
xnor U7891 (N_7891,N_7635,N_7622);
nor U7892 (N_7892,N_7774,N_7752);
or U7893 (N_7893,N_7726,N_7737);
nand U7894 (N_7894,N_7662,N_7723);
or U7895 (N_7895,N_7705,N_7759);
and U7896 (N_7896,N_7788,N_7612);
nor U7897 (N_7897,N_7769,N_7783);
and U7898 (N_7898,N_7648,N_7782);
and U7899 (N_7899,N_7619,N_7607);
or U7900 (N_7900,N_7695,N_7635);
or U7901 (N_7901,N_7752,N_7646);
nor U7902 (N_7902,N_7796,N_7682);
nand U7903 (N_7903,N_7730,N_7769);
and U7904 (N_7904,N_7603,N_7778);
or U7905 (N_7905,N_7622,N_7709);
nand U7906 (N_7906,N_7785,N_7606);
and U7907 (N_7907,N_7656,N_7765);
nand U7908 (N_7908,N_7715,N_7758);
nor U7909 (N_7909,N_7709,N_7720);
or U7910 (N_7910,N_7789,N_7787);
xor U7911 (N_7911,N_7611,N_7673);
nand U7912 (N_7912,N_7790,N_7701);
and U7913 (N_7913,N_7662,N_7627);
and U7914 (N_7914,N_7620,N_7662);
nor U7915 (N_7915,N_7689,N_7693);
nand U7916 (N_7916,N_7698,N_7775);
or U7917 (N_7917,N_7621,N_7616);
xor U7918 (N_7918,N_7676,N_7695);
nor U7919 (N_7919,N_7783,N_7618);
or U7920 (N_7920,N_7745,N_7732);
and U7921 (N_7921,N_7707,N_7640);
and U7922 (N_7922,N_7784,N_7655);
nand U7923 (N_7923,N_7702,N_7733);
or U7924 (N_7924,N_7699,N_7630);
xor U7925 (N_7925,N_7743,N_7740);
nand U7926 (N_7926,N_7722,N_7792);
nand U7927 (N_7927,N_7712,N_7703);
and U7928 (N_7928,N_7661,N_7742);
nor U7929 (N_7929,N_7652,N_7786);
and U7930 (N_7930,N_7793,N_7640);
xnor U7931 (N_7931,N_7630,N_7682);
and U7932 (N_7932,N_7782,N_7758);
nand U7933 (N_7933,N_7771,N_7766);
or U7934 (N_7934,N_7779,N_7797);
and U7935 (N_7935,N_7663,N_7727);
nor U7936 (N_7936,N_7612,N_7713);
or U7937 (N_7937,N_7624,N_7653);
and U7938 (N_7938,N_7760,N_7757);
or U7939 (N_7939,N_7797,N_7718);
nand U7940 (N_7940,N_7785,N_7712);
and U7941 (N_7941,N_7688,N_7629);
or U7942 (N_7942,N_7764,N_7662);
xor U7943 (N_7943,N_7753,N_7690);
nor U7944 (N_7944,N_7749,N_7651);
nor U7945 (N_7945,N_7724,N_7675);
nor U7946 (N_7946,N_7750,N_7633);
or U7947 (N_7947,N_7735,N_7612);
nand U7948 (N_7948,N_7768,N_7790);
xor U7949 (N_7949,N_7753,N_7611);
and U7950 (N_7950,N_7733,N_7790);
nand U7951 (N_7951,N_7684,N_7673);
nand U7952 (N_7952,N_7634,N_7797);
and U7953 (N_7953,N_7624,N_7644);
nand U7954 (N_7954,N_7708,N_7681);
nor U7955 (N_7955,N_7746,N_7688);
or U7956 (N_7956,N_7643,N_7657);
and U7957 (N_7957,N_7637,N_7777);
nor U7958 (N_7958,N_7625,N_7688);
nand U7959 (N_7959,N_7611,N_7724);
and U7960 (N_7960,N_7652,N_7634);
and U7961 (N_7961,N_7763,N_7667);
and U7962 (N_7962,N_7768,N_7780);
or U7963 (N_7963,N_7744,N_7735);
nand U7964 (N_7964,N_7611,N_7684);
nand U7965 (N_7965,N_7757,N_7784);
nor U7966 (N_7966,N_7651,N_7633);
nor U7967 (N_7967,N_7667,N_7605);
nand U7968 (N_7968,N_7744,N_7696);
or U7969 (N_7969,N_7650,N_7606);
nor U7970 (N_7970,N_7734,N_7610);
or U7971 (N_7971,N_7799,N_7648);
nor U7972 (N_7972,N_7779,N_7766);
xnor U7973 (N_7973,N_7615,N_7778);
xor U7974 (N_7974,N_7692,N_7738);
and U7975 (N_7975,N_7715,N_7635);
nor U7976 (N_7976,N_7682,N_7675);
nand U7977 (N_7977,N_7743,N_7715);
nor U7978 (N_7978,N_7717,N_7795);
nand U7979 (N_7979,N_7702,N_7634);
and U7980 (N_7980,N_7742,N_7676);
nor U7981 (N_7981,N_7618,N_7635);
and U7982 (N_7982,N_7696,N_7731);
and U7983 (N_7983,N_7644,N_7790);
or U7984 (N_7984,N_7753,N_7677);
xnor U7985 (N_7985,N_7607,N_7643);
and U7986 (N_7986,N_7788,N_7638);
and U7987 (N_7987,N_7638,N_7674);
or U7988 (N_7988,N_7631,N_7774);
or U7989 (N_7989,N_7777,N_7631);
nand U7990 (N_7990,N_7789,N_7688);
and U7991 (N_7991,N_7743,N_7770);
or U7992 (N_7992,N_7655,N_7708);
or U7993 (N_7993,N_7709,N_7659);
and U7994 (N_7994,N_7771,N_7718);
or U7995 (N_7995,N_7644,N_7712);
xnor U7996 (N_7996,N_7753,N_7602);
nor U7997 (N_7997,N_7647,N_7624);
nand U7998 (N_7998,N_7664,N_7603);
nand U7999 (N_7999,N_7633,N_7798);
nand U8000 (N_8000,N_7818,N_7865);
or U8001 (N_8001,N_7894,N_7832);
or U8002 (N_8002,N_7995,N_7926);
nand U8003 (N_8003,N_7891,N_7807);
or U8004 (N_8004,N_7964,N_7895);
nand U8005 (N_8005,N_7944,N_7848);
or U8006 (N_8006,N_7902,N_7933);
xnor U8007 (N_8007,N_7830,N_7973);
or U8008 (N_8008,N_7863,N_7859);
or U8009 (N_8009,N_7884,N_7831);
nand U8010 (N_8010,N_7864,N_7805);
nand U8011 (N_8011,N_7890,N_7941);
and U8012 (N_8012,N_7880,N_7892);
xor U8013 (N_8013,N_7938,N_7956);
or U8014 (N_8014,N_7827,N_7881);
nor U8015 (N_8015,N_7949,N_7867);
nand U8016 (N_8016,N_7850,N_7812);
xnor U8017 (N_8017,N_7950,N_7903);
or U8018 (N_8018,N_7911,N_7920);
nand U8019 (N_8019,N_7924,N_7959);
or U8020 (N_8020,N_7983,N_7861);
nand U8021 (N_8021,N_7978,N_7958);
nand U8022 (N_8022,N_7855,N_7815);
and U8023 (N_8023,N_7904,N_7997);
xor U8024 (N_8024,N_7838,N_7811);
and U8025 (N_8025,N_7803,N_7993);
nor U8026 (N_8026,N_7819,N_7946);
and U8027 (N_8027,N_7875,N_7960);
or U8028 (N_8028,N_7988,N_7921);
or U8029 (N_8029,N_7951,N_7856);
nand U8030 (N_8030,N_7847,N_7925);
nor U8031 (N_8031,N_7908,N_7947);
and U8032 (N_8032,N_7915,N_7910);
nand U8033 (N_8033,N_7874,N_7998);
or U8034 (N_8034,N_7808,N_7854);
nand U8035 (N_8035,N_7954,N_7940);
nand U8036 (N_8036,N_7916,N_7866);
or U8037 (N_8037,N_7844,N_7957);
or U8038 (N_8038,N_7918,N_7852);
or U8039 (N_8039,N_7984,N_7900);
nor U8040 (N_8040,N_7928,N_7932);
and U8041 (N_8041,N_7839,N_7842);
nor U8042 (N_8042,N_7857,N_7840);
or U8043 (N_8043,N_7929,N_7825);
or U8044 (N_8044,N_7979,N_7975);
nor U8045 (N_8045,N_7945,N_7965);
or U8046 (N_8046,N_7885,N_7898);
nand U8047 (N_8047,N_7943,N_7980);
and U8048 (N_8048,N_7886,N_7888);
nand U8049 (N_8049,N_7906,N_7942);
nand U8050 (N_8050,N_7824,N_7999);
and U8051 (N_8051,N_7834,N_7966);
nand U8052 (N_8052,N_7877,N_7953);
nor U8053 (N_8053,N_7948,N_7802);
xnor U8054 (N_8054,N_7851,N_7813);
or U8055 (N_8055,N_7937,N_7869);
and U8056 (N_8056,N_7853,N_7934);
nor U8057 (N_8057,N_7878,N_7905);
and U8058 (N_8058,N_7821,N_7955);
and U8059 (N_8059,N_7873,N_7914);
and U8060 (N_8060,N_7841,N_7835);
and U8061 (N_8061,N_7990,N_7846);
or U8062 (N_8062,N_7879,N_7801);
or U8063 (N_8063,N_7809,N_7935);
nor U8064 (N_8064,N_7913,N_7836);
nand U8065 (N_8065,N_7893,N_7816);
nor U8066 (N_8066,N_7822,N_7992);
or U8067 (N_8067,N_7837,N_7976);
nor U8068 (N_8068,N_7870,N_7981);
nor U8069 (N_8069,N_7994,N_7989);
xnor U8070 (N_8070,N_7917,N_7826);
and U8071 (N_8071,N_7883,N_7860);
nand U8072 (N_8072,N_7868,N_7972);
or U8073 (N_8073,N_7899,N_7974);
xnor U8074 (N_8074,N_7909,N_7887);
nor U8075 (N_8075,N_7996,N_7829);
or U8076 (N_8076,N_7897,N_7817);
or U8077 (N_8077,N_7896,N_7833);
nand U8078 (N_8078,N_7963,N_7889);
or U8079 (N_8079,N_7971,N_7814);
nor U8080 (N_8080,N_7862,N_7986);
and U8081 (N_8081,N_7843,N_7968);
nand U8082 (N_8082,N_7845,N_7923);
nand U8083 (N_8083,N_7849,N_7823);
nor U8084 (N_8084,N_7912,N_7882);
nor U8085 (N_8085,N_7806,N_7871);
nand U8086 (N_8086,N_7901,N_7828);
xnor U8087 (N_8087,N_7985,N_7876);
nor U8088 (N_8088,N_7991,N_7820);
nor U8089 (N_8089,N_7982,N_7922);
nand U8090 (N_8090,N_7939,N_7967);
nand U8091 (N_8091,N_7907,N_7961);
or U8092 (N_8092,N_7931,N_7936);
or U8093 (N_8093,N_7800,N_7969);
nand U8094 (N_8094,N_7927,N_7952);
nand U8095 (N_8095,N_7962,N_7919);
xnor U8096 (N_8096,N_7930,N_7872);
and U8097 (N_8097,N_7804,N_7858);
or U8098 (N_8098,N_7987,N_7810);
nand U8099 (N_8099,N_7970,N_7977);
or U8100 (N_8100,N_7893,N_7815);
nor U8101 (N_8101,N_7920,N_7955);
or U8102 (N_8102,N_7943,N_7869);
nand U8103 (N_8103,N_7932,N_7852);
nand U8104 (N_8104,N_7800,N_7995);
and U8105 (N_8105,N_7848,N_7904);
nand U8106 (N_8106,N_7888,N_7909);
xnor U8107 (N_8107,N_7818,N_7868);
or U8108 (N_8108,N_7844,N_7899);
nand U8109 (N_8109,N_7995,N_7826);
nand U8110 (N_8110,N_7998,N_7917);
xor U8111 (N_8111,N_7938,N_7824);
or U8112 (N_8112,N_7824,N_7964);
xnor U8113 (N_8113,N_7985,N_7809);
xnor U8114 (N_8114,N_7937,N_7959);
nand U8115 (N_8115,N_7857,N_7872);
nor U8116 (N_8116,N_7950,N_7820);
or U8117 (N_8117,N_7980,N_7948);
or U8118 (N_8118,N_7990,N_7940);
nand U8119 (N_8119,N_7804,N_7924);
nor U8120 (N_8120,N_7910,N_7858);
nand U8121 (N_8121,N_7967,N_7925);
or U8122 (N_8122,N_7944,N_7953);
nand U8123 (N_8123,N_7953,N_7924);
or U8124 (N_8124,N_7895,N_7924);
nand U8125 (N_8125,N_7832,N_7984);
xor U8126 (N_8126,N_7958,N_7833);
or U8127 (N_8127,N_7830,N_7853);
nand U8128 (N_8128,N_7827,N_7820);
nand U8129 (N_8129,N_7813,N_7966);
and U8130 (N_8130,N_7947,N_7910);
xor U8131 (N_8131,N_7843,N_7895);
nor U8132 (N_8132,N_7872,N_7982);
nand U8133 (N_8133,N_7986,N_7884);
nand U8134 (N_8134,N_7834,N_7921);
nand U8135 (N_8135,N_7963,N_7960);
nand U8136 (N_8136,N_7852,N_7964);
or U8137 (N_8137,N_7882,N_7921);
or U8138 (N_8138,N_7867,N_7806);
nor U8139 (N_8139,N_7967,N_7942);
nor U8140 (N_8140,N_7829,N_7945);
or U8141 (N_8141,N_7815,N_7868);
and U8142 (N_8142,N_7952,N_7800);
nor U8143 (N_8143,N_7817,N_7914);
nor U8144 (N_8144,N_7855,N_7964);
nand U8145 (N_8145,N_7889,N_7863);
and U8146 (N_8146,N_7965,N_7857);
or U8147 (N_8147,N_7975,N_7862);
nand U8148 (N_8148,N_7837,N_7957);
and U8149 (N_8149,N_7970,N_7814);
or U8150 (N_8150,N_7844,N_7984);
nand U8151 (N_8151,N_7814,N_7883);
nand U8152 (N_8152,N_7973,N_7863);
nand U8153 (N_8153,N_7906,N_7866);
and U8154 (N_8154,N_7842,N_7949);
nor U8155 (N_8155,N_7975,N_7838);
or U8156 (N_8156,N_7897,N_7919);
nor U8157 (N_8157,N_7833,N_7910);
xor U8158 (N_8158,N_7966,N_7953);
and U8159 (N_8159,N_7967,N_7983);
nor U8160 (N_8160,N_7890,N_7852);
nand U8161 (N_8161,N_7997,N_7939);
nor U8162 (N_8162,N_7980,N_7825);
and U8163 (N_8163,N_7896,N_7882);
or U8164 (N_8164,N_7922,N_7948);
and U8165 (N_8165,N_7827,N_7911);
nor U8166 (N_8166,N_7833,N_7952);
nand U8167 (N_8167,N_7894,N_7833);
xnor U8168 (N_8168,N_7976,N_7995);
nand U8169 (N_8169,N_7880,N_7918);
and U8170 (N_8170,N_7860,N_7865);
or U8171 (N_8171,N_7917,N_7972);
or U8172 (N_8172,N_7813,N_7847);
or U8173 (N_8173,N_7902,N_7971);
nor U8174 (N_8174,N_7995,N_7932);
or U8175 (N_8175,N_7973,N_7901);
xnor U8176 (N_8176,N_7855,N_7985);
and U8177 (N_8177,N_7888,N_7934);
or U8178 (N_8178,N_7874,N_7917);
or U8179 (N_8179,N_7811,N_7945);
nor U8180 (N_8180,N_7805,N_7824);
nor U8181 (N_8181,N_7809,N_7965);
nor U8182 (N_8182,N_7852,N_7870);
nand U8183 (N_8183,N_7952,N_7823);
xnor U8184 (N_8184,N_7996,N_7814);
nand U8185 (N_8185,N_7859,N_7988);
nor U8186 (N_8186,N_7985,N_7922);
and U8187 (N_8187,N_7838,N_7994);
nand U8188 (N_8188,N_7932,N_7870);
nor U8189 (N_8189,N_7910,N_7872);
nor U8190 (N_8190,N_7968,N_7922);
nand U8191 (N_8191,N_7955,N_7811);
or U8192 (N_8192,N_7979,N_7971);
or U8193 (N_8193,N_7825,N_7802);
or U8194 (N_8194,N_7900,N_7877);
or U8195 (N_8195,N_7995,N_7985);
and U8196 (N_8196,N_7807,N_7878);
or U8197 (N_8197,N_7907,N_7813);
nor U8198 (N_8198,N_7963,N_7809);
or U8199 (N_8199,N_7853,N_7813);
nor U8200 (N_8200,N_8074,N_8174);
nand U8201 (N_8201,N_8124,N_8046);
and U8202 (N_8202,N_8172,N_8035);
nand U8203 (N_8203,N_8187,N_8064);
or U8204 (N_8204,N_8019,N_8031);
nor U8205 (N_8205,N_8013,N_8041);
xnor U8206 (N_8206,N_8146,N_8003);
or U8207 (N_8207,N_8106,N_8156);
nor U8208 (N_8208,N_8092,N_8020);
nor U8209 (N_8209,N_8083,N_8097);
nand U8210 (N_8210,N_8079,N_8138);
or U8211 (N_8211,N_8080,N_8163);
or U8212 (N_8212,N_8112,N_8129);
and U8213 (N_8213,N_8175,N_8144);
and U8214 (N_8214,N_8023,N_8052);
and U8215 (N_8215,N_8186,N_8049);
nand U8216 (N_8216,N_8054,N_8040);
nand U8217 (N_8217,N_8090,N_8152);
nor U8218 (N_8218,N_8057,N_8076);
and U8219 (N_8219,N_8061,N_8102);
nand U8220 (N_8220,N_8139,N_8073);
and U8221 (N_8221,N_8117,N_8179);
nand U8222 (N_8222,N_8075,N_8119);
or U8223 (N_8223,N_8095,N_8167);
nor U8224 (N_8224,N_8012,N_8149);
or U8225 (N_8225,N_8063,N_8157);
or U8226 (N_8226,N_8050,N_8042);
nor U8227 (N_8227,N_8008,N_8010);
or U8228 (N_8228,N_8181,N_8105);
xor U8229 (N_8229,N_8184,N_8123);
or U8230 (N_8230,N_8059,N_8065);
xor U8231 (N_8231,N_8161,N_8016);
nor U8232 (N_8232,N_8150,N_8033);
or U8233 (N_8233,N_8196,N_8032);
and U8234 (N_8234,N_8062,N_8026);
nand U8235 (N_8235,N_8170,N_8017);
nor U8236 (N_8236,N_8081,N_8027);
nand U8237 (N_8237,N_8142,N_8143);
xor U8238 (N_8238,N_8193,N_8151);
and U8239 (N_8239,N_8141,N_8171);
nand U8240 (N_8240,N_8189,N_8067);
or U8241 (N_8241,N_8185,N_8096);
nor U8242 (N_8242,N_8120,N_8114);
nor U8243 (N_8243,N_8045,N_8018);
nand U8244 (N_8244,N_8029,N_8188);
and U8245 (N_8245,N_8145,N_8110);
nor U8246 (N_8246,N_8078,N_8028);
nor U8247 (N_8247,N_8055,N_8194);
and U8248 (N_8248,N_8037,N_8053);
and U8249 (N_8249,N_8159,N_8177);
and U8250 (N_8250,N_8158,N_8118);
and U8251 (N_8251,N_8101,N_8108);
and U8252 (N_8252,N_8051,N_8166);
and U8253 (N_8253,N_8169,N_8126);
nand U8254 (N_8254,N_8056,N_8190);
nor U8255 (N_8255,N_8134,N_8071);
nand U8256 (N_8256,N_8001,N_8128);
xor U8257 (N_8257,N_8094,N_8098);
nor U8258 (N_8258,N_8005,N_8111);
or U8259 (N_8259,N_8164,N_8022);
nand U8260 (N_8260,N_8021,N_8088);
nor U8261 (N_8261,N_8084,N_8038);
and U8262 (N_8262,N_8182,N_8116);
nor U8263 (N_8263,N_8007,N_8011);
and U8264 (N_8264,N_8072,N_8132);
nand U8265 (N_8265,N_8107,N_8048);
xor U8266 (N_8266,N_8133,N_8103);
or U8267 (N_8267,N_8004,N_8197);
nand U8268 (N_8268,N_8127,N_8085);
or U8269 (N_8269,N_8180,N_8137);
nand U8270 (N_8270,N_8115,N_8069);
or U8271 (N_8271,N_8178,N_8140);
or U8272 (N_8272,N_8099,N_8070);
nand U8273 (N_8273,N_8192,N_8100);
nand U8274 (N_8274,N_8025,N_8113);
or U8275 (N_8275,N_8086,N_8043);
xor U8276 (N_8276,N_8136,N_8036);
and U8277 (N_8277,N_8068,N_8131);
nand U8278 (N_8278,N_8148,N_8199);
nor U8279 (N_8279,N_8039,N_8047);
nor U8280 (N_8280,N_8044,N_8000);
or U8281 (N_8281,N_8058,N_8060);
xnor U8282 (N_8282,N_8066,N_8198);
nand U8283 (N_8283,N_8147,N_8122);
xnor U8284 (N_8284,N_8087,N_8162);
xnor U8285 (N_8285,N_8173,N_8121);
and U8286 (N_8286,N_8002,N_8160);
nor U8287 (N_8287,N_8014,N_8091);
nor U8288 (N_8288,N_8195,N_8176);
nand U8289 (N_8289,N_8155,N_8104);
xnor U8290 (N_8290,N_8089,N_8015);
and U8291 (N_8291,N_8006,N_8034);
nor U8292 (N_8292,N_8082,N_8191);
nor U8293 (N_8293,N_8153,N_8093);
and U8294 (N_8294,N_8135,N_8165);
nand U8295 (N_8295,N_8077,N_8168);
or U8296 (N_8296,N_8125,N_8030);
and U8297 (N_8297,N_8109,N_8024);
and U8298 (N_8298,N_8183,N_8154);
nor U8299 (N_8299,N_8130,N_8009);
xnor U8300 (N_8300,N_8102,N_8041);
nand U8301 (N_8301,N_8186,N_8098);
xor U8302 (N_8302,N_8185,N_8131);
or U8303 (N_8303,N_8022,N_8077);
nor U8304 (N_8304,N_8182,N_8181);
and U8305 (N_8305,N_8159,N_8065);
nor U8306 (N_8306,N_8038,N_8106);
nor U8307 (N_8307,N_8068,N_8023);
or U8308 (N_8308,N_8033,N_8103);
or U8309 (N_8309,N_8039,N_8060);
and U8310 (N_8310,N_8005,N_8109);
nand U8311 (N_8311,N_8069,N_8131);
nor U8312 (N_8312,N_8077,N_8162);
or U8313 (N_8313,N_8054,N_8006);
and U8314 (N_8314,N_8138,N_8188);
and U8315 (N_8315,N_8155,N_8068);
nor U8316 (N_8316,N_8092,N_8138);
xor U8317 (N_8317,N_8052,N_8177);
nand U8318 (N_8318,N_8053,N_8108);
nand U8319 (N_8319,N_8094,N_8121);
nand U8320 (N_8320,N_8134,N_8180);
nor U8321 (N_8321,N_8071,N_8181);
and U8322 (N_8322,N_8147,N_8028);
and U8323 (N_8323,N_8117,N_8173);
xor U8324 (N_8324,N_8066,N_8082);
or U8325 (N_8325,N_8013,N_8144);
and U8326 (N_8326,N_8019,N_8093);
nand U8327 (N_8327,N_8183,N_8057);
nor U8328 (N_8328,N_8154,N_8137);
xor U8329 (N_8329,N_8052,N_8151);
and U8330 (N_8330,N_8072,N_8008);
nand U8331 (N_8331,N_8114,N_8101);
nor U8332 (N_8332,N_8094,N_8048);
or U8333 (N_8333,N_8120,N_8106);
or U8334 (N_8334,N_8154,N_8091);
or U8335 (N_8335,N_8008,N_8061);
or U8336 (N_8336,N_8138,N_8052);
nand U8337 (N_8337,N_8115,N_8170);
or U8338 (N_8338,N_8188,N_8017);
and U8339 (N_8339,N_8155,N_8149);
nor U8340 (N_8340,N_8091,N_8022);
nand U8341 (N_8341,N_8091,N_8096);
or U8342 (N_8342,N_8095,N_8064);
or U8343 (N_8343,N_8160,N_8017);
and U8344 (N_8344,N_8044,N_8077);
or U8345 (N_8345,N_8052,N_8115);
nand U8346 (N_8346,N_8065,N_8110);
nor U8347 (N_8347,N_8194,N_8146);
nand U8348 (N_8348,N_8099,N_8183);
and U8349 (N_8349,N_8021,N_8067);
nor U8350 (N_8350,N_8000,N_8009);
or U8351 (N_8351,N_8198,N_8177);
or U8352 (N_8352,N_8045,N_8014);
or U8353 (N_8353,N_8142,N_8059);
and U8354 (N_8354,N_8157,N_8132);
nor U8355 (N_8355,N_8033,N_8170);
xor U8356 (N_8356,N_8077,N_8172);
or U8357 (N_8357,N_8045,N_8124);
nor U8358 (N_8358,N_8190,N_8146);
and U8359 (N_8359,N_8106,N_8036);
or U8360 (N_8360,N_8053,N_8173);
nand U8361 (N_8361,N_8105,N_8052);
nand U8362 (N_8362,N_8198,N_8155);
xor U8363 (N_8363,N_8196,N_8004);
nand U8364 (N_8364,N_8003,N_8170);
nand U8365 (N_8365,N_8041,N_8167);
and U8366 (N_8366,N_8081,N_8133);
nand U8367 (N_8367,N_8123,N_8079);
nand U8368 (N_8368,N_8153,N_8000);
nand U8369 (N_8369,N_8094,N_8066);
nor U8370 (N_8370,N_8089,N_8072);
xor U8371 (N_8371,N_8137,N_8129);
and U8372 (N_8372,N_8036,N_8160);
xnor U8373 (N_8373,N_8131,N_8045);
or U8374 (N_8374,N_8024,N_8128);
or U8375 (N_8375,N_8049,N_8198);
nor U8376 (N_8376,N_8000,N_8131);
and U8377 (N_8377,N_8026,N_8036);
and U8378 (N_8378,N_8143,N_8135);
and U8379 (N_8379,N_8084,N_8184);
nand U8380 (N_8380,N_8113,N_8145);
or U8381 (N_8381,N_8044,N_8160);
xor U8382 (N_8382,N_8161,N_8084);
nor U8383 (N_8383,N_8104,N_8028);
nor U8384 (N_8384,N_8074,N_8053);
nand U8385 (N_8385,N_8195,N_8189);
or U8386 (N_8386,N_8053,N_8150);
or U8387 (N_8387,N_8185,N_8172);
and U8388 (N_8388,N_8129,N_8157);
or U8389 (N_8389,N_8125,N_8011);
nor U8390 (N_8390,N_8038,N_8183);
or U8391 (N_8391,N_8173,N_8146);
xnor U8392 (N_8392,N_8180,N_8192);
or U8393 (N_8393,N_8185,N_8165);
and U8394 (N_8394,N_8153,N_8086);
and U8395 (N_8395,N_8075,N_8097);
or U8396 (N_8396,N_8153,N_8188);
nand U8397 (N_8397,N_8064,N_8081);
or U8398 (N_8398,N_8042,N_8095);
nand U8399 (N_8399,N_8156,N_8089);
nand U8400 (N_8400,N_8391,N_8212);
and U8401 (N_8401,N_8359,N_8250);
or U8402 (N_8402,N_8397,N_8375);
and U8403 (N_8403,N_8301,N_8219);
and U8404 (N_8404,N_8333,N_8394);
or U8405 (N_8405,N_8268,N_8277);
xnor U8406 (N_8406,N_8314,N_8207);
or U8407 (N_8407,N_8365,N_8396);
nand U8408 (N_8408,N_8327,N_8354);
xor U8409 (N_8409,N_8384,N_8349);
nand U8410 (N_8410,N_8217,N_8390);
xnor U8411 (N_8411,N_8246,N_8267);
nand U8412 (N_8412,N_8319,N_8290);
or U8413 (N_8413,N_8317,N_8280);
nand U8414 (N_8414,N_8329,N_8278);
nor U8415 (N_8415,N_8363,N_8369);
or U8416 (N_8416,N_8200,N_8379);
nand U8417 (N_8417,N_8241,N_8325);
or U8418 (N_8418,N_8370,N_8323);
nand U8419 (N_8419,N_8218,N_8353);
or U8420 (N_8420,N_8374,N_8331);
and U8421 (N_8421,N_8239,N_8203);
nor U8422 (N_8422,N_8324,N_8227);
and U8423 (N_8423,N_8381,N_8285);
and U8424 (N_8424,N_8233,N_8294);
and U8425 (N_8425,N_8265,N_8308);
nand U8426 (N_8426,N_8259,N_8266);
or U8427 (N_8427,N_8262,N_8240);
or U8428 (N_8428,N_8297,N_8235);
and U8429 (N_8429,N_8350,N_8242);
xnor U8430 (N_8430,N_8213,N_8335);
nor U8431 (N_8431,N_8348,N_8284);
or U8432 (N_8432,N_8292,N_8253);
nand U8433 (N_8433,N_8315,N_8274);
nor U8434 (N_8434,N_8307,N_8286);
and U8435 (N_8435,N_8205,N_8392);
nor U8436 (N_8436,N_8269,N_8321);
and U8437 (N_8437,N_8251,N_8377);
nor U8438 (N_8438,N_8313,N_8204);
or U8439 (N_8439,N_8380,N_8234);
or U8440 (N_8440,N_8326,N_8320);
and U8441 (N_8441,N_8249,N_8340);
nand U8442 (N_8442,N_8300,N_8322);
nand U8443 (N_8443,N_8398,N_8282);
or U8444 (N_8444,N_8245,N_8298);
xnor U8445 (N_8445,N_8368,N_8273);
nor U8446 (N_8446,N_8352,N_8395);
xnor U8447 (N_8447,N_8337,N_8376);
nor U8448 (N_8448,N_8338,N_8372);
nor U8449 (N_8449,N_8254,N_8371);
nand U8450 (N_8450,N_8385,N_8237);
and U8451 (N_8451,N_8276,N_8316);
and U8452 (N_8452,N_8393,N_8201);
or U8453 (N_8453,N_8305,N_8302);
nand U8454 (N_8454,N_8270,N_8378);
nand U8455 (N_8455,N_8351,N_8382);
xor U8456 (N_8456,N_8360,N_8347);
nand U8457 (N_8457,N_8231,N_8255);
and U8458 (N_8458,N_8358,N_8264);
nor U8459 (N_8459,N_8343,N_8342);
and U8460 (N_8460,N_8364,N_8222);
nor U8461 (N_8461,N_8328,N_8256);
xor U8462 (N_8462,N_8296,N_8383);
nor U8463 (N_8463,N_8216,N_8248);
nand U8464 (N_8464,N_8260,N_8209);
nand U8465 (N_8465,N_8388,N_8334);
or U8466 (N_8466,N_8202,N_8210);
or U8467 (N_8467,N_8220,N_8309);
nand U8468 (N_8468,N_8225,N_8362);
nor U8469 (N_8469,N_8211,N_8226);
nor U8470 (N_8470,N_8275,N_8312);
nor U8471 (N_8471,N_8229,N_8230);
nand U8472 (N_8472,N_8330,N_8306);
nand U8473 (N_8473,N_8357,N_8224);
nand U8474 (N_8474,N_8214,N_8208);
or U8475 (N_8475,N_8223,N_8244);
and U8476 (N_8476,N_8287,N_8339);
nor U8477 (N_8477,N_8346,N_8261);
and U8478 (N_8478,N_8272,N_8243);
nor U8479 (N_8479,N_8345,N_8271);
nor U8480 (N_8480,N_8238,N_8361);
or U8481 (N_8481,N_8336,N_8311);
nor U8482 (N_8482,N_8299,N_8252);
nor U8483 (N_8483,N_8257,N_8215);
nand U8484 (N_8484,N_8366,N_8304);
and U8485 (N_8485,N_8386,N_8247);
nor U8486 (N_8486,N_8356,N_8373);
nor U8487 (N_8487,N_8263,N_8279);
and U8488 (N_8488,N_8367,N_8399);
nor U8489 (N_8489,N_8387,N_8295);
nand U8490 (N_8490,N_8236,N_8310);
nand U8491 (N_8491,N_8281,N_8389);
nand U8492 (N_8492,N_8344,N_8288);
nor U8493 (N_8493,N_8318,N_8289);
nand U8494 (N_8494,N_8221,N_8303);
and U8495 (N_8495,N_8293,N_8291);
nand U8496 (N_8496,N_8206,N_8228);
nor U8497 (N_8497,N_8232,N_8283);
and U8498 (N_8498,N_8355,N_8341);
nand U8499 (N_8499,N_8258,N_8332);
and U8500 (N_8500,N_8279,N_8242);
nor U8501 (N_8501,N_8210,N_8231);
or U8502 (N_8502,N_8374,N_8260);
nand U8503 (N_8503,N_8277,N_8243);
or U8504 (N_8504,N_8304,N_8364);
or U8505 (N_8505,N_8228,N_8300);
nand U8506 (N_8506,N_8328,N_8266);
xnor U8507 (N_8507,N_8360,N_8242);
nor U8508 (N_8508,N_8328,N_8216);
nor U8509 (N_8509,N_8246,N_8221);
nand U8510 (N_8510,N_8205,N_8389);
and U8511 (N_8511,N_8201,N_8382);
nand U8512 (N_8512,N_8353,N_8336);
nor U8513 (N_8513,N_8288,N_8244);
nor U8514 (N_8514,N_8211,N_8314);
nor U8515 (N_8515,N_8356,N_8311);
nor U8516 (N_8516,N_8336,N_8335);
or U8517 (N_8517,N_8329,N_8289);
and U8518 (N_8518,N_8234,N_8356);
nand U8519 (N_8519,N_8370,N_8254);
nor U8520 (N_8520,N_8348,N_8279);
or U8521 (N_8521,N_8383,N_8362);
nor U8522 (N_8522,N_8303,N_8203);
nor U8523 (N_8523,N_8281,N_8352);
nor U8524 (N_8524,N_8285,N_8209);
and U8525 (N_8525,N_8244,N_8200);
nand U8526 (N_8526,N_8380,N_8214);
or U8527 (N_8527,N_8232,N_8326);
nor U8528 (N_8528,N_8237,N_8330);
and U8529 (N_8529,N_8331,N_8252);
or U8530 (N_8530,N_8374,N_8248);
or U8531 (N_8531,N_8244,N_8260);
or U8532 (N_8532,N_8380,N_8359);
and U8533 (N_8533,N_8381,N_8320);
and U8534 (N_8534,N_8235,N_8309);
nor U8535 (N_8535,N_8298,N_8348);
or U8536 (N_8536,N_8299,N_8215);
nand U8537 (N_8537,N_8382,N_8328);
nand U8538 (N_8538,N_8353,N_8288);
nand U8539 (N_8539,N_8241,N_8308);
or U8540 (N_8540,N_8389,N_8312);
nor U8541 (N_8541,N_8279,N_8221);
and U8542 (N_8542,N_8272,N_8394);
or U8543 (N_8543,N_8272,N_8369);
nor U8544 (N_8544,N_8331,N_8302);
nor U8545 (N_8545,N_8363,N_8255);
or U8546 (N_8546,N_8229,N_8253);
or U8547 (N_8547,N_8393,N_8298);
nor U8548 (N_8548,N_8362,N_8315);
nor U8549 (N_8549,N_8238,N_8365);
nor U8550 (N_8550,N_8277,N_8354);
nand U8551 (N_8551,N_8308,N_8314);
nand U8552 (N_8552,N_8287,N_8286);
nand U8553 (N_8553,N_8379,N_8261);
or U8554 (N_8554,N_8358,N_8316);
nor U8555 (N_8555,N_8393,N_8232);
nand U8556 (N_8556,N_8214,N_8396);
nand U8557 (N_8557,N_8387,N_8241);
xnor U8558 (N_8558,N_8281,N_8203);
nor U8559 (N_8559,N_8322,N_8287);
or U8560 (N_8560,N_8334,N_8224);
nor U8561 (N_8561,N_8248,N_8317);
and U8562 (N_8562,N_8309,N_8252);
nor U8563 (N_8563,N_8202,N_8235);
or U8564 (N_8564,N_8221,N_8201);
nor U8565 (N_8565,N_8356,N_8346);
xor U8566 (N_8566,N_8380,N_8242);
and U8567 (N_8567,N_8313,N_8394);
nor U8568 (N_8568,N_8398,N_8285);
nor U8569 (N_8569,N_8206,N_8275);
and U8570 (N_8570,N_8296,N_8319);
and U8571 (N_8571,N_8386,N_8366);
and U8572 (N_8572,N_8308,N_8303);
or U8573 (N_8573,N_8272,N_8290);
xnor U8574 (N_8574,N_8247,N_8239);
or U8575 (N_8575,N_8399,N_8305);
nor U8576 (N_8576,N_8217,N_8235);
nor U8577 (N_8577,N_8396,N_8358);
and U8578 (N_8578,N_8242,N_8371);
or U8579 (N_8579,N_8269,N_8246);
nor U8580 (N_8580,N_8222,N_8397);
xnor U8581 (N_8581,N_8370,N_8257);
nand U8582 (N_8582,N_8283,N_8200);
nand U8583 (N_8583,N_8327,N_8278);
and U8584 (N_8584,N_8341,N_8245);
or U8585 (N_8585,N_8316,N_8328);
nand U8586 (N_8586,N_8334,N_8311);
and U8587 (N_8587,N_8285,N_8279);
nor U8588 (N_8588,N_8256,N_8369);
xor U8589 (N_8589,N_8292,N_8335);
and U8590 (N_8590,N_8203,N_8290);
or U8591 (N_8591,N_8312,N_8373);
and U8592 (N_8592,N_8315,N_8343);
nand U8593 (N_8593,N_8200,N_8337);
and U8594 (N_8594,N_8393,N_8274);
nor U8595 (N_8595,N_8281,N_8347);
or U8596 (N_8596,N_8261,N_8270);
nor U8597 (N_8597,N_8250,N_8383);
or U8598 (N_8598,N_8398,N_8393);
nor U8599 (N_8599,N_8290,N_8229);
or U8600 (N_8600,N_8442,N_8573);
or U8601 (N_8601,N_8464,N_8452);
nand U8602 (N_8602,N_8517,N_8437);
nand U8603 (N_8603,N_8548,N_8420);
nor U8604 (N_8604,N_8447,N_8559);
and U8605 (N_8605,N_8500,N_8551);
nand U8606 (N_8606,N_8408,N_8443);
and U8607 (N_8607,N_8504,N_8554);
or U8608 (N_8608,N_8496,N_8401);
nand U8609 (N_8609,N_8450,N_8468);
and U8610 (N_8610,N_8595,N_8516);
nand U8611 (N_8611,N_8511,N_8484);
or U8612 (N_8612,N_8530,N_8421);
xor U8613 (N_8613,N_8415,N_8451);
nor U8614 (N_8614,N_8473,N_8485);
nor U8615 (N_8615,N_8429,N_8585);
and U8616 (N_8616,N_8491,N_8534);
or U8617 (N_8617,N_8509,N_8456);
or U8618 (N_8618,N_8409,N_8580);
xor U8619 (N_8619,N_8579,N_8584);
or U8620 (N_8620,N_8567,N_8432);
nor U8621 (N_8621,N_8527,N_8413);
nor U8622 (N_8622,N_8545,N_8556);
nand U8623 (N_8623,N_8419,N_8476);
or U8624 (N_8624,N_8402,N_8553);
and U8625 (N_8625,N_8482,N_8519);
and U8626 (N_8626,N_8588,N_8591);
nand U8627 (N_8627,N_8596,N_8459);
nor U8628 (N_8628,N_8577,N_8515);
or U8629 (N_8629,N_8542,N_8525);
or U8630 (N_8630,N_8520,N_8430);
xor U8631 (N_8631,N_8465,N_8466);
nand U8632 (N_8632,N_8490,N_8564);
and U8633 (N_8633,N_8457,N_8543);
and U8634 (N_8634,N_8470,N_8411);
or U8635 (N_8635,N_8449,N_8558);
nor U8636 (N_8636,N_8535,N_8441);
nor U8637 (N_8637,N_8507,N_8460);
or U8638 (N_8638,N_8404,N_8480);
or U8639 (N_8639,N_8494,N_8495);
and U8640 (N_8640,N_8546,N_8557);
nor U8641 (N_8641,N_8592,N_8533);
nor U8642 (N_8642,N_8555,N_8562);
nand U8643 (N_8643,N_8438,N_8563);
or U8644 (N_8644,N_8524,N_8424);
and U8645 (N_8645,N_8586,N_8568);
nand U8646 (N_8646,N_8467,N_8581);
nand U8647 (N_8647,N_8561,N_8400);
nand U8648 (N_8648,N_8486,N_8483);
xor U8649 (N_8649,N_8514,N_8532);
xnor U8650 (N_8650,N_8529,N_8418);
nand U8651 (N_8651,N_8547,N_8425);
or U8652 (N_8652,N_8422,N_8566);
or U8653 (N_8653,N_8410,N_8497);
and U8654 (N_8654,N_8599,N_8427);
xnor U8655 (N_8655,N_8598,N_8501);
and U8656 (N_8656,N_8407,N_8479);
nand U8657 (N_8657,N_8541,N_8576);
nand U8658 (N_8658,N_8458,N_8474);
and U8659 (N_8659,N_8569,N_8508);
and U8660 (N_8660,N_8471,N_8570);
or U8661 (N_8661,N_8445,N_8505);
and U8662 (N_8662,N_8489,N_8523);
nand U8663 (N_8663,N_8550,N_8440);
nor U8664 (N_8664,N_8502,N_8406);
or U8665 (N_8665,N_8454,N_8518);
xor U8666 (N_8666,N_8540,N_8423);
or U8667 (N_8667,N_8434,N_8469);
or U8668 (N_8668,N_8499,N_8510);
nand U8669 (N_8669,N_8582,N_8405);
or U8670 (N_8670,N_8487,N_8426);
and U8671 (N_8671,N_8575,N_8506);
nand U8672 (N_8672,N_8433,N_8572);
xor U8673 (N_8673,N_8403,N_8528);
xor U8674 (N_8674,N_8536,N_8417);
nand U8675 (N_8675,N_8436,N_8521);
or U8676 (N_8676,N_8560,N_8571);
or U8677 (N_8677,N_8565,N_8538);
xor U8678 (N_8678,N_8414,N_8578);
nor U8679 (N_8679,N_8594,N_8488);
and U8680 (N_8680,N_8444,N_8475);
nor U8681 (N_8681,N_8503,N_8492);
nand U8682 (N_8682,N_8537,N_8512);
and U8683 (N_8683,N_8498,N_8412);
nand U8684 (N_8684,N_8461,N_8428);
nor U8685 (N_8685,N_8526,N_8455);
and U8686 (N_8686,N_8446,N_8590);
xor U8687 (N_8687,N_8463,N_8593);
or U8688 (N_8688,N_8544,N_8574);
nor U8689 (N_8689,N_8462,N_8589);
and U8690 (N_8690,N_8453,N_8435);
or U8691 (N_8691,N_8448,N_8513);
nor U8692 (N_8692,N_8552,N_8416);
nand U8693 (N_8693,N_8478,N_8472);
nor U8694 (N_8694,N_8549,N_8539);
nand U8695 (N_8695,N_8531,N_8597);
and U8696 (N_8696,N_8522,N_8481);
or U8697 (N_8697,N_8439,N_8493);
and U8698 (N_8698,N_8431,N_8583);
nor U8699 (N_8699,N_8587,N_8477);
and U8700 (N_8700,N_8548,N_8589);
or U8701 (N_8701,N_8570,N_8583);
and U8702 (N_8702,N_8571,N_8426);
or U8703 (N_8703,N_8481,N_8425);
and U8704 (N_8704,N_8503,N_8481);
nor U8705 (N_8705,N_8564,N_8474);
and U8706 (N_8706,N_8480,N_8477);
xor U8707 (N_8707,N_8538,N_8462);
nor U8708 (N_8708,N_8591,N_8476);
and U8709 (N_8709,N_8454,N_8588);
nor U8710 (N_8710,N_8548,N_8519);
nor U8711 (N_8711,N_8507,N_8541);
nor U8712 (N_8712,N_8558,N_8459);
and U8713 (N_8713,N_8487,N_8445);
nor U8714 (N_8714,N_8448,N_8507);
nor U8715 (N_8715,N_8493,N_8581);
or U8716 (N_8716,N_8488,N_8477);
xor U8717 (N_8717,N_8552,N_8520);
and U8718 (N_8718,N_8441,N_8570);
nand U8719 (N_8719,N_8559,N_8431);
nand U8720 (N_8720,N_8560,N_8534);
nor U8721 (N_8721,N_8508,N_8475);
nor U8722 (N_8722,N_8452,N_8477);
or U8723 (N_8723,N_8457,N_8527);
xnor U8724 (N_8724,N_8549,N_8407);
or U8725 (N_8725,N_8555,N_8514);
xor U8726 (N_8726,N_8565,N_8469);
nand U8727 (N_8727,N_8492,N_8493);
nor U8728 (N_8728,N_8492,N_8462);
or U8729 (N_8729,N_8529,N_8515);
or U8730 (N_8730,N_8540,N_8562);
or U8731 (N_8731,N_8551,N_8593);
nor U8732 (N_8732,N_8409,N_8584);
and U8733 (N_8733,N_8443,N_8406);
and U8734 (N_8734,N_8518,N_8557);
nor U8735 (N_8735,N_8477,N_8538);
and U8736 (N_8736,N_8455,N_8483);
xor U8737 (N_8737,N_8581,N_8585);
nor U8738 (N_8738,N_8558,N_8551);
and U8739 (N_8739,N_8535,N_8446);
nor U8740 (N_8740,N_8433,N_8582);
or U8741 (N_8741,N_8469,N_8526);
nand U8742 (N_8742,N_8569,N_8533);
nor U8743 (N_8743,N_8408,N_8555);
and U8744 (N_8744,N_8524,N_8460);
and U8745 (N_8745,N_8468,N_8437);
xor U8746 (N_8746,N_8463,N_8582);
or U8747 (N_8747,N_8477,N_8546);
or U8748 (N_8748,N_8538,N_8490);
and U8749 (N_8749,N_8464,N_8522);
nor U8750 (N_8750,N_8591,N_8533);
or U8751 (N_8751,N_8567,N_8540);
xor U8752 (N_8752,N_8592,N_8418);
xor U8753 (N_8753,N_8411,N_8465);
or U8754 (N_8754,N_8402,N_8514);
nand U8755 (N_8755,N_8547,N_8542);
xnor U8756 (N_8756,N_8572,N_8574);
or U8757 (N_8757,N_8583,N_8512);
nor U8758 (N_8758,N_8443,N_8487);
and U8759 (N_8759,N_8446,N_8506);
or U8760 (N_8760,N_8433,N_8496);
and U8761 (N_8761,N_8525,N_8552);
nand U8762 (N_8762,N_8545,N_8550);
xnor U8763 (N_8763,N_8530,N_8563);
and U8764 (N_8764,N_8404,N_8497);
nand U8765 (N_8765,N_8448,N_8487);
nand U8766 (N_8766,N_8434,N_8526);
nor U8767 (N_8767,N_8498,N_8546);
nor U8768 (N_8768,N_8560,N_8406);
nand U8769 (N_8769,N_8455,N_8406);
and U8770 (N_8770,N_8429,N_8581);
and U8771 (N_8771,N_8469,N_8463);
or U8772 (N_8772,N_8512,N_8599);
nor U8773 (N_8773,N_8489,N_8495);
xnor U8774 (N_8774,N_8458,N_8408);
and U8775 (N_8775,N_8444,N_8427);
or U8776 (N_8776,N_8564,N_8594);
and U8777 (N_8777,N_8449,N_8411);
and U8778 (N_8778,N_8598,N_8507);
and U8779 (N_8779,N_8555,N_8406);
xnor U8780 (N_8780,N_8566,N_8496);
and U8781 (N_8781,N_8532,N_8546);
nor U8782 (N_8782,N_8587,N_8573);
nor U8783 (N_8783,N_8407,N_8512);
nand U8784 (N_8784,N_8583,N_8589);
and U8785 (N_8785,N_8421,N_8566);
nor U8786 (N_8786,N_8517,N_8516);
or U8787 (N_8787,N_8545,N_8458);
nand U8788 (N_8788,N_8589,N_8576);
and U8789 (N_8789,N_8594,N_8472);
nor U8790 (N_8790,N_8436,N_8460);
nor U8791 (N_8791,N_8420,N_8514);
nand U8792 (N_8792,N_8440,N_8546);
nand U8793 (N_8793,N_8428,N_8434);
and U8794 (N_8794,N_8534,N_8580);
or U8795 (N_8795,N_8552,N_8495);
nor U8796 (N_8796,N_8457,N_8576);
and U8797 (N_8797,N_8570,N_8557);
nand U8798 (N_8798,N_8577,N_8492);
xnor U8799 (N_8799,N_8529,N_8487);
nand U8800 (N_8800,N_8702,N_8772);
nor U8801 (N_8801,N_8770,N_8791);
nor U8802 (N_8802,N_8757,N_8676);
nor U8803 (N_8803,N_8799,N_8747);
and U8804 (N_8804,N_8653,N_8729);
or U8805 (N_8805,N_8739,N_8719);
or U8806 (N_8806,N_8704,N_8617);
or U8807 (N_8807,N_8635,N_8624);
and U8808 (N_8808,N_8661,N_8644);
nor U8809 (N_8809,N_8604,N_8793);
xnor U8810 (N_8810,N_8742,N_8693);
nor U8811 (N_8811,N_8795,N_8728);
or U8812 (N_8812,N_8792,N_8633);
or U8813 (N_8813,N_8701,N_8606);
and U8814 (N_8814,N_8616,N_8680);
nand U8815 (N_8815,N_8735,N_8683);
nor U8816 (N_8816,N_8748,N_8674);
or U8817 (N_8817,N_8749,N_8798);
or U8818 (N_8818,N_8695,N_8634);
nor U8819 (N_8819,N_8744,N_8767);
nor U8820 (N_8820,N_8672,N_8670);
and U8821 (N_8821,N_8629,N_8755);
nand U8822 (N_8822,N_8774,N_8658);
xor U8823 (N_8823,N_8756,N_8776);
nand U8824 (N_8824,N_8696,N_8602);
and U8825 (N_8825,N_8738,N_8609);
xor U8826 (N_8826,N_8732,N_8611);
and U8827 (N_8827,N_8766,N_8679);
xor U8828 (N_8828,N_8675,N_8768);
and U8829 (N_8829,N_8769,N_8773);
and U8830 (N_8830,N_8708,N_8651);
or U8831 (N_8831,N_8694,N_8669);
or U8832 (N_8832,N_8685,N_8631);
or U8833 (N_8833,N_8671,N_8745);
or U8834 (N_8834,N_8765,N_8614);
nor U8835 (N_8835,N_8613,N_8686);
nand U8836 (N_8836,N_8640,N_8706);
or U8837 (N_8837,N_8794,N_8657);
and U8838 (N_8838,N_8688,N_8715);
or U8839 (N_8839,N_8648,N_8625);
or U8840 (N_8840,N_8783,N_8668);
or U8841 (N_8841,N_8660,N_8750);
or U8842 (N_8842,N_8605,N_8779);
xor U8843 (N_8843,N_8678,N_8758);
xnor U8844 (N_8844,N_8726,N_8682);
or U8845 (N_8845,N_8796,N_8628);
and U8846 (N_8846,N_8626,N_8786);
nand U8847 (N_8847,N_8612,N_8788);
and U8848 (N_8848,N_8664,N_8673);
xnor U8849 (N_8849,N_8607,N_8622);
nand U8850 (N_8850,N_8785,N_8636);
nor U8851 (N_8851,N_8730,N_8659);
or U8852 (N_8852,N_8643,N_8781);
or U8853 (N_8853,N_8698,N_8615);
and U8854 (N_8854,N_8761,N_8649);
nand U8855 (N_8855,N_8717,N_8647);
and U8856 (N_8856,N_8752,N_8632);
nor U8857 (N_8857,N_8790,N_8754);
and U8858 (N_8858,N_8619,N_8618);
or U8859 (N_8859,N_8677,N_8684);
xor U8860 (N_8860,N_8700,N_8652);
nor U8861 (N_8861,N_8763,N_8665);
or U8862 (N_8862,N_8610,N_8630);
nor U8863 (N_8863,N_8703,N_8601);
or U8864 (N_8864,N_8603,N_8760);
and U8865 (N_8865,N_8713,N_8620);
and U8866 (N_8866,N_8650,N_8627);
nor U8867 (N_8867,N_8656,N_8787);
nor U8868 (N_8868,N_8782,N_8751);
and U8869 (N_8869,N_8645,N_8731);
and U8870 (N_8870,N_8716,N_8641);
xor U8871 (N_8871,N_8778,N_8721);
nor U8872 (N_8872,N_8734,N_8723);
or U8873 (N_8873,N_8762,N_8777);
nor U8874 (N_8874,N_8789,N_8663);
nand U8875 (N_8875,N_8689,N_8720);
and U8876 (N_8876,N_8727,N_8699);
nand U8877 (N_8877,N_8662,N_8737);
or U8878 (N_8878,N_8714,N_8771);
nor U8879 (N_8879,N_8759,N_8608);
nand U8880 (N_8880,N_8638,N_8600);
nand U8881 (N_8881,N_8621,N_8764);
nor U8882 (N_8882,N_8705,N_8753);
or U8883 (N_8883,N_8639,N_8692);
or U8884 (N_8884,N_8707,N_8784);
and U8885 (N_8885,N_8718,N_8775);
xnor U8886 (N_8886,N_8623,N_8697);
and U8887 (N_8887,N_8710,N_8797);
or U8888 (N_8888,N_8666,N_8681);
and U8889 (N_8889,N_8654,N_8711);
and U8890 (N_8890,N_8687,N_8637);
and U8891 (N_8891,N_8667,N_8724);
and U8892 (N_8892,N_8780,N_8709);
nor U8893 (N_8893,N_8712,N_8722);
xor U8894 (N_8894,N_8736,N_8642);
nor U8895 (N_8895,N_8725,N_8741);
and U8896 (N_8896,N_8733,N_8655);
xnor U8897 (N_8897,N_8690,N_8691);
nor U8898 (N_8898,N_8740,N_8646);
or U8899 (N_8899,N_8743,N_8746);
nand U8900 (N_8900,N_8720,N_8724);
nor U8901 (N_8901,N_8642,N_8743);
and U8902 (N_8902,N_8783,N_8772);
nor U8903 (N_8903,N_8723,N_8642);
or U8904 (N_8904,N_8712,N_8603);
nor U8905 (N_8905,N_8685,N_8707);
nand U8906 (N_8906,N_8618,N_8749);
nand U8907 (N_8907,N_8603,N_8784);
nor U8908 (N_8908,N_8791,N_8789);
nand U8909 (N_8909,N_8653,N_8681);
and U8910 (N_8910,N_8602,N_8742);
nand U8911 (N_8911,N_8778,N_8685);
nor U8912 (N_8912,N_8613,N_8608);
or U8913 (N_8913,N_8709,N_8679);
and U8914 (N_8914,N_8620,N_8678);
xnor U8915 (N_8915,N_8673,N_8757);
or U8916 (N_8916,N_8709,N_8767);
or U8917 (N_8917,N_8697,N_8728);
nand U8918 (N_8918,N_8608,N_8611);
or U8919 (N_8919,N_8726,N_8751);
nand U8920 (N_8920,N_8707,N_8642);
and U8921 (N_8921,N_8653,N_8614);
or U8922 (N_8922,N_8791,N_8761);
nor U8923 (N_8923,N_8799,N_8665);
nor U8924 (N_8924,N_8630,N_8686);
nor U8925 (N_8925,N_8600,N_8623);
nor U8926 (N_8926,N_8691,N_8701);
or U8927 (N_8927,N_8699,N_8600);
or U8928 (N_8928,N_8753,N_8653);
or U8929 (N_8929,N_8621,N_8704);
and U8930 (N_8930,N_8622,N_8678);
nand U8931 (N_8931,N_8744,N_8699);
and U8932 (N_8932,N_8795,N_8689);
nand U8933 (N_8933,N_8789,N_8621);
and U8934 (N_8934,N_8706,N_8686);
xnor U8935 (N_8935,N_8787,N_8796);
and U8936 (N_8936,N_8716,N_8614);
nor U8937 (N_8937,N_8617,N_8609);
nand U8938 (N_8938,N_8643,N_8779);
nor U8939 (N_8939,N_8727,N_8652);
and U8940 (N_8940,N_8711,N_8758);
xnor U8941 (N_8941,N_8653,N_8762);
nand U8942 (N_8942,N_8744,N_8736);
or U8943 (N_8943,N_8614,N_8777);
nand U8944 (N_8944,N_8759,N_8771);
and U8945 (N_8945,N_8678,N_8697);
nor U8946 (N_8946,N_8609,N_8602);
or U8947 (N_8947,N_8674,N_8670);
nand U8948 (N_8948,N_8602,N_8654);
and U8949 (N_8949,N_8735,N_8760);
and U8950 (N_8950,N_8788,N_8757);
nand U8951 (N_8951,N_8635,N_8630);
nor U8952 (N_8952,N_8743,N_8798);
xnor U8953 (N_8953,N_8715,N_8651);
nor U8954 (N_8954,N_8699,N_8718);
or U8955 (N_8955,N_8604,N_8716);
xnor U8956 (N_8956,N_8650,N_8790);
nor U8957 (N_8957,N_8780,N_8657);
nand U8958 (N_8958,N_8769,N_8657);
and U8959 (N_8959,N_8712,N_8615);
nor U8960 (N_8960,N_8785,N_8798);
nor U8961 (N_8961,N_8706,N_8617);
nor U8962 (N_8962,N_8695,N_8652);
nor U8963 (N_8963,N_8758,N_8796);
and U8964 (N_8964,N_8675,N_8773);
nor U8965 (N_8965,N_8682,N_8654);
nand U8966 (N_8966,N_8724,N_8616);
or U8967 (N_8967,N_8780,N_8675);
nand U8968 (N_8968,N_8623,N_8740);
nor U8969 (N_8969,N_8794,N_8687);
and U8970 (N_8970,N_8628,N_8667);
nor U8971 (N_8971,N_8659,N_8612);
nor U8972 (N_8972,N_8767,N_8647);
nand U8973 (N_8973,N_8650,N_8718);
or U8974 (N_8974,N_8697,N_8730);
and U8975 (N_8975,N_8621,N_8651);
and U8976 (N_8976,N_8744,N_8757);
nand U8977 (N_8977,N_8771,N_8760);
or U8978 (N_8978,N_8634,N_8644);
and U8979 (N_8979,N_8609,N_8676);
nand U8980 (N_8980,N_8662,N_8638);
nor U8981 (N_8981,N_8680,N_8706);
xnor U8982 (N_8982,N_8778,N_8711);
or U8983 (N_8983,N_8705,N_8642);
nor U8984 (N_8984,N_8732,N_8786);
nor U8985 (N_8985,N_8718,N_8671);
or U8986 (N_8986,N_8791,N_8683);
nand U8987 (N_8987,N_8740,N_8695);
and U8988 (N_8988,N_8604,N_8636);
nand U8989 (N_8989,N_8767,N_8612);
xor U8990 (N_8990,N_8703,N_8621);
xor U8991 (N_8991,N_8684,N_8671);
and U8992 (N_8992,N_8652,N_8707);
and U8993 (N_8993,N_8789,N_8665);
xnor U8994 (N_8994,N_8699,N_8717);
nor U8995 (N_8995,N_8654,N_8783);
and U8996 (N_8996,N_8684,N_8617);
and U8997 (N_8997,N_8797,N_8708);
nand U8998 (N_8998,N_8766,N_8676);
nand U8999 (N_8999,N_8721,N_8674);
nand U9000 (N_9000,N_8878,N_8806);
or U9001 (N_9001,N_8949,N_8983);
nand U9002 (N_9002,N_8800,N_8824);
or U9003 (N_9003,N_8977,N_8877);
and U9004 (N_9004,N_8873,N_8860);
nand U9005 (N_9005,N_8823,N_8930);
nand U9006 (N_9006,N_8929,N_8844);
or U9007 (N_9007,N_8887,N_8923);
or U9008 (N_9008,N_8845,N_8898);
nor U9009 (N_9009,N_8954,N_8828);
nand U9010 (N_9010,N_8960,N_8852);
and U9011 (N_9011,N_8999,N_8849);
nand U9012 (N_9012,N_8984,N_8918);
xor U9013 (N_9013,N_8833,N_8911);
nor U9014 (N_9014,N_8904,N_8856);
or U9015 (N_9015,N_8869,N_8858);
nand U9016 (N_9016,N_8836,N_8815);
or U9017 (N_9017,N_8958,N_8926);
nand U9018 (N_9018,N_8952,N_8972);
nand U9019 (N_9019,N_8995,N_8908);
nand U9020 (N_9020,N_8969,N_8892);
nand U9021 (N_9021,N_8853,N_8808);
or U9022 (N_9022,N_8834,N_8978);
nor U9023 (N_9023,N_8913,N_8990);
nand U9024 (N_9024,N_8835,N_8997);
and U9025 (N_9025,N_8927,N_8925);
and U9026 (N_9026,N_8967,N_8979);
xor U9027 (N_9027,N_8981,N_8850);
or U9028 (N_9028,N_8883,N_8946);
nand U9029 (N_9029,N_8945,N_8943);
or U9030 (N_9030,N_8826,N_8841);
or U9031 (N_9031,N_8859,N_8813);
nand U9032 (N_9032,N_8955,N_8980);
nand U9033 (N_9033,N_8821,N_8964);
or U9034 (N_9034,N_8837,N_8961);
xnor U9035 (N_9035,N_8819,N_8915);
xnor U9036 (N_9036,N_8963,N_8919);
or U9037 (N_9037,N_8912,N_8890);
nand U9038 (N_9038,N_8991,N_8801);
nand U9039 (N_9039,N_8920,N_8865);
or U9040 (N_9040,N_8965,N_8968);
or U9041 (N_9041,N_8811,N_8966);
or U9042 (N_9042,N_8917,N_8947);
and U9043 (N_9043,N_8818,N_8914);
and U9044 (N_9044,N_8922,N_8891);
nor U9045 (N_9045,N_8839,N_8827);
nor U9046 (N_9046,N_8897,N_8816);
nor U9047 (N_9047,N_8899,N_8886);
and U9048 (N_9048,N_8987,N_8875);
nor U9049 (N_9049,N_8907,N_8996);
nand U9050 (N_9050,N_8910,N_8989);
and U9051 (N_9051,N_8994,N_8934);
or U9052 (N_9052,N_8831,N_8896);
and U9053 (N_9053,N_8894,N_8956);
and U9054 (N_9054,N_8804,N_8951);
or U9055 (N_9055,N_8959,N_8931);
xor U9056 (N_9056,N_8851,N_8893);
or U9057 (N_9057,N_8957,N_8884);
and U9058 (N_9058,N_8879,N_8941);
or U9059 (N_9059,N_8832,N_8944);
nand U9060 (N_9060,N_8900,N_8822);
xnor U9061 (N_9061,N_8810,N_8942);
nor U9062 (N_9062,N_8974,N_8872);
nor U9063 (N_9063,N_8971,N_8939);
xnor U9064 (N_9064,N_8857,N_8985);
xor U9065 (N_9065,N_8848,N_8976);
or U9066 (N_9066,N_8829,N_8906);
nor U9067 (N_9067,N_8820,N_8905);
xnor U9068 (N_9068,N_8901,N_8895);
xnor U9069 (N_9069,N_8903,N_8928);
and U9070 (N_9070,N_8986,N_8814);
or U9071 (N_9071,N_8870,N_8809);
or U9072 (N_9072,N_8861,N_8885);
nor U9073 (N_9073,N_8936,N_8950);
or U9074 (N_9074,N_8882,N_8867);
nor U9075 (N_9075,N_8916,N_8864);
and U9076 (N_9076,N_8924,N_8888);
nor U9077 (N_9077,N_8940,N_8992);
nor U9078 (N_9078,N_8921,N_8838);
nor U9079 (N_9079,N_8975,N_8998);
and U9080 (N_9080,N_8802,N_8909);
nand U9081 (N_9081,N_8933,N_8982);
and U9082 (N_9082,N_8868,N_8830);
xor U9083 (N_9083,N_8847,N_8803);
and U9084 (N_9084,N_8953,N_8880);
or U9085 (N_9085,N_8962,N_8937);
nor U9086 (N_9086,N_8846,N_8938);
nand U9087 (N_9087,N_8817,N_8874);
nand U9088 (N_9088,N_8825,N_8993);
and U9089 (N_9089,N_8843,N_8805);
nor U9090 (N_9090,N_8807,N_8889);
or U9091 (N_9091,N_8935,N_8863);
and U9092 (N_9092,N_8871,N_8973);
nor U9093 (N_9093,N_8854,N_8855);
xor U9094 (N_9094,N_8970,N_8876);
and U9095 (N_9095,N_8988,N_8866);
nand U9096 (N_9096,N_8881,N_8862);
and U9097 (N_9097,N_8840,N_8842);
nor U9098 (N_9098,N_8902,N_8948);
xor U9099 (N_9099,N_8932,N_8812);
nor U9100 (N_9100,N_8864,N_8962);
or U9101 (N_9101,N_8861,N_8835);
nor U9102 (N_9102,N_8979,N_8955);
xnor U9103 (N_9103,N_8801,N_8864);
and U9104 (N_9104,N_8933,N_8945);
nand U9105 (N_9105,N_8825,N_8966);
and U9106 (N_9106,N_8890,N_8954);
nand U9107 (N_9107,N_8902,N_8895);
xnor U9108 (N_9108,N_8902,N_8928);
nand U9109 (N_9109,N_8957,N_8971);
and U9110 (N_9110,N_8830,N_8846);
or U9111 (N_9111,N_8968,N_8823);
nor U9112 (N_9112,N_8983,N_8990);
or U9113 (N_9113,N_8874,N_8948);
xor U9114 (N_9114,N_8876,N_8893);
nand U9115 (N_9115,N_8899,N_8911);
or U9116 (N_9116,N_8858,N_8902);
xnor U9117 (N_9117,N_8905,N_8985);
and U9118 (N_9118,N_8918,N_8843);
nor U9119 (N_9119,N_8819,N_8850);
or U9120 (N_9120,N_8903,N_8854);
xnor U9121 (N_9121,N_8945,N_8827);
nor U9122 (N_9122,N_8901,N_8842);
and U9123 (N_9123,N_8937,N_8985);
and U9124 (N_9124,N_8894,N_8892);
nor U9125 (N_9125,N_8904,N_8990);
nand U9126 (N_9126,N_8872,N_8865);
nor U9127 (N_9127,N_8814,N_8854);
or U9128 (N_9128,N_8984,N_8935);
nor U9129 (N_9129,N_8825,N_8889);
nor U9130 (N_9130,N_8837,N_8910);
and U9131 (N_9131,N_8858,N_8947);
xnor U9132 (N_9132,N_8896,N_8852);
or U9133 (N_9133,N_8941,N_8885);
nand U9134 (N_9134,N_8864,N_8924);
nor U9135 (N_9135,N_8996,N_8879);
or U9136 (N_9136,N_8810,N_8881);
and U9137 (N_9137,N_8884,N_8969);
or U9138 (N_9138,N_8878,N_8870);
and U9139 (N_9139,N_8935,N_8925);
and U9140 (N_9140,N_8896,N_8928);
and U9141 (N_9141,N_8896,N_8851);
nor U9142 (N_9142,N_8891,N_8880);
nor U9143 (N_9143,N_8887,N_8942);
nor U9144 (N_9144,N_8913,N_8860);
nand U9145 (N_9145,N_8835,N_8848);
nand U9146 (N_9146,N_8853,N_8887);
nand U9147 (N_9147,N_8854,N_8902);
xnor U9148 (N_9148,N_8900,N_8888);
and U9149 (N_9149,N_8911,N_8873);
or U9150 (N_9150,N_8870,N_8943);
or U9151 (N_9151,N_8831,N_8868);
nor U9152 (N_9152,N_8951,N_8843);
nand U9153 (N_9153,N_8828,N_8873);
xnor U9154 (N_9154,N_8855,N_8919);
nor U9155 (N_9155,N_8872,N_8882);
and U9156 (N_9156,N_8836,N_8972);
nor U9157 (N_9157,N_8903,N_8824);
and U9158 (N_9158,N_8838,N_8933);
nand U9159 (N_9159,N_8845,N_8967);
xor U9160 (N_9160,N_8954,N_8951);
or U9161 (N_9161,N_8958,N_8831);
nand U9162 (N_9162,N_8972,N_8947);
nor U9163 (N_9163,N_8958,N_8976);
or U9164 (N_9164,N_8931,N_8842);
nor U9165 (N_9165,N_8987,N_8831);
or U9166 (N_9166,N_8897,N_8887);
nor U9167 (N_9167,N_8857,N_8893);
and U9168 (N_9168,N_8886,N_8945);
nor U9169 (N_9169,N_8903,N_8988);
nor U9170 (N_9170,N_8894,N_8981);
and U9171 (N_9171,N_8876,N_8902);
and U9172 (N_9172,N_8871,N_8950);
and U9173 (N_9173,N_8906,N_8817);
or U9174 (N_9174,N_8868,N_8925);
and U9175 (N_9175,N_8831,N_8928);
or U9176 (N_9176,N_8994,N_8932);
and U9177 (N_9177,N_8992,N_8906);
nor U9178 (N_9178,N_8862,N_8907);
nor U9179 (N_9179,N_8999,N_8997);
nand U9180 (N_9180,N_8995,N_8864);
xor U9181 (N_9181,N_8951,N_8952);
and U9182 (N_9182,N_8910,N_8930);
and U9183 (N_9183,N_8816,N_8955);
nor U9184 (N_9184,N_8847,N_8943);
and U9185 (N_9185,N_8874,N_8877);
and U9186 (N_9186,N_8912,N_8859);
and U9187 (N_9187,N_8833,N_8851);
nor U9188 (N_9188,N_8832,N_8879);
nor U9189 (N_9189,N_8893,N_8990);
or U9190 (N_9190,N_8919,N_8869);
nor U9191 (N_9191,N_8897,N_8861);
xnor U9192 (N_9192,N_8849,N_8967);
and U9193 (N_9193,N_8880,N_8868);
or U9194 (N_9194,N_8893,N_8965);
xor U9195 (N_9195,N_8848,N_8963);
or U9196 (N_9196,N_8812,N_8935);
nand U9197 (N_9197,N_8864,N_8958);
nand U9198 (N_9198,N_8990,N_8905);
nor U9199 (N_9199,N_8915,N_8894);
and U9200 (N_9200,N_9137,N_9159);
and U9201 (N_9201,N_9102,N_9031);
or U9202 (N_9202,N_9038,N_9053);
and U9203 (N_9203,N_9016,N_9029);
and U9204 (N_9204,N_9041,N_9186);
nor U9205 (N_9205,N_9122,N_9093);
nor U9206 (N_9206,N_9149,N_9005);
or U9207 (N_9207,N_9063,N_9034);
and U9208 (N_9208,N_9067,N_9074);
nor U9209 (N_9209,N_9071,N_9019);
nor U9210 (N_9210,N_9023,N_9014);
nand U9211 (N_9211,N_9124,N_9142);
or U9212 (N_9212,N_9037,N_9198);
nor U9213 (N_9213,N_9151,N_9009);
and U9214 (N_9214,N_9128,N_9166);
nand U9215 (N_9215,N_9013,N_9158);
xnor U9216 (N_9216,N_9082,N_9148);
nand U9217 (N_9217,N_9086,N_9135);
nor U9218 (N_9218,N_9160,N_9015);
and U9219 (N_9219,N_9105,N_9152);
and U9220 (N_9220,N_9043,N_9182);
xor U9221 (N_9221,N_9069,N_9104);
and U9222 (N_9222,N_9101,N_9130);
or U9223 (N_9223,N_9116,N_9052);
xor U9224 (N_9224,N_9134,N_9024);
or U9225 (N_9225,N_9188,N_9164);
or U9226 (N_9226,N_9125,N_9193);
xnor U9227 (N_9227,N_9042,N_9099);
or U9228 (N_9228,N_9039,N_9068);
nor U9229 (N_9229,N_9073,N_9021);
and U9230 (N_9230,N_9051,N_9036);
and U9231 (N_9231,N_9094,N_9006);
and U9232 (N_9232,N_9095,N_9055);
nor U9233 (N_9233,N_9110,N_9180);
nand U9234 (N_9234,N_9194,N_9129);
nand U9235 (N_9235,N_9106,N_9044);
and U9236 (N_9236,N_9155,N_9062);
and U9237 (N_9237,N_9167,N_9022);
nand U9238 (N_9238,N_9061,N_9000);
or U9239 (N_9239,N_9181,N_9177);
nor U9240 (N_9240,N_9045,N_9027);
and U9241 (N_9241,N_9169,N_9119);
or U9242 (N_9242,N_9084,N_9191);
nand U9243 (N_9243,N_9057,N_9187);
and U9244 (N_9244,N_9070,N_9143);
nand U9245 (N_9245,N_9126,N_9168);
or U9246 (N_9246,N_9098,N_9199);
or U9247 (N_9247,N_9107,N_9046);
and U9248 (N_9248,N_9111,N_9144);
nor U9249 (N_9249,N_9179,N_9025);
xor U9250 (N_9250,N_9088,N_9035);
nor U9251 (N_9251,N_9060,N_9140);
and U9252 (N_9252,N_9189,N_9097);
nand U9253 (N_9253,N_9058,N_9049);
or U9254 (N_9254,N_9017,N_9112);
and U9255 (N_9255,N_9004,N_9108);
xnor U9256 (N_9256,N_9087,N_9103);
xor U9257 (N_9257,N_9145,N_9026);
nand U9258 (N_9258,N_9141,N_9075);
and U9259 (N_9259,N_9118,N_9007);
nor U9260 (N_9260,N_9048,N_9184);
nand U9261 (N_9261,N_9020,N_9056);
and U9262 (N_9262,N_9150,N_9173);
xor U9263 (N_9263,N_9011,N_9132);
and U9264 (N_9264,N_9090,N_9138);
nand U9265 (N_9265,N_9065,N_9092);
and U9266 (N_9266,N_9001,N_9047);
nor U9267 (N_9267,N_9050,N_9096);
xor U9268 (N_9268,N_9109,N_9157);
or U9269 (N_9269,N_9139,N_9127);
nand U9270 (N_9270,N_9161,N_9113);
or U9271 (N_9271,N_9059,N_9040);
xor U9272 (N_9272,N_9030,N_9171);
xor U9273 (N_9273,N_9170,N_9028);
nand U9274 (N_9274,N_9174,N_9081);
nand U9275 (N_9275,N_9076,N_9175);
and U9276 (N_9276,N_9121,N_9080);
nand U9277 (N_9277,N_9078,N_9178);
and U9278 (N_9278,N_9032,N_9115);
nor U9279 (N_9279,N_9133,N_9146);
and U9280 (N_9280,N_9196,N_9131);
nor U9281 (N_9281,N_9018,N_9154);
and U9282 (N_9282,N_9123,N_9054);
nor U9283 (N_9283,N_9192,N_9089);
and U9284 (N_9284,N_9079,N_9156);
and U9285 (N_9285,N_9120,N_9190);
nand U9286 (N_9286,N_9185,N_9163);
or U9287 (N_9287,N_9183,N_9114);
or U9288 (N_9288,N_9064,N_9091);
xor U9289 (N_9289,N_9072,N_9153);
nor U9290 (N_9290,N_9172,N_9195);
xnor U9291 (N_9291,N_9100,N_9176);
xnor U9292 (N_9292,N_9165,N_9083);
or U9293 (N_9293,N_9162,N_9003);
xnor U9294 (N_9294,N_9010,N_9077);
nor U9295 (N_9295,N_9066,N_9136);
or U9296 (N_9296,N_9002,N_9008);
or U9297 (N_9297,N_9085,N_9197);
nand U9298 (N_9298,N_9147,N_9012);
xor U9299 (N_9299,N_9033,N_9117);
and U9300 (N_9300,N_9163,N_9130);
nand U9301 (N_9301,N_9096,N_9024);
and U9302 (N_9302,N_9105,N_9087);
nand U9303 (N_9303,N_9020,N_9095);
and U9304 (N_9304,N_9050,N_9124);
and U9305 (N_9305,N_9126,N_9086);
nor U9306 (N_9306,N_9119,N_9099);
or U9307 (N_9307,N_9124,N_9081);
nand U9308 (N_9308,N_9118,N_9045);
xnor U9309 (N_9309,N_9038,N_9198);
nand U9310 (N_9310,N_9128,N_9154);
or U9311 (N_9311,N_9185,N_9149);
and U9312 (N_9312,N_9110,N_9194);
and U9313 (N_9313,N_9077,N_9083);
nor U9314 (N_9314,N_9195,N_9041);
and U9315 (N_9315,N_9060,N_9011);
nand U9316 (N_9316,N_9032,N_9002);
and U9317 (N_9317,N_9119,N_9138);
nand U9318 (N_9318,N_9092,N_9087);
and U9319 (N_9319,N_9175,N_9111);
and U9320 (N_9320,N_9094,N_9157);
nor U9321 (N_9321,N_9193,N_9010);
nand U9322 (N_9322,N_9007,N_9090);
and U9323 (N_9323,N_9092,N_9182);
and U9324 (N_9324,N_9196,N_9123);
nor U9325 (N_9325,N_9050,N_9066);
nand U9326 (N_9326,N_9144,N_9073);
and U9327 (N_9327,N_9077,N_9067);
and U9328 (N_9328,N_9043,N_9029);
or U9329 (N_9329,N_9148,N_9093);
nor U9330 (N_9330,N_9169,N_9035);
nor U9331 (N_9331,N_9035,N_9006);
nand U9332 (N_9332,N_9154,N_9196);
nand U9333 (N_9333,N_9063,N_9090);
or U9334 (N_9334,N_9173,N_9031);
or U9335 (N_9335,N_9002,N_9051);
nor U9336 (N_9336,N_9122,N_9159);
and U9337 (N_9337,N_9069,N_9171);
xor U9338 (N_9338,N_9062,N_9079);
and U9339 (N_9339,N_9084,N_9139);
or U9340 (N_9340,N_9061,N_9019);
nor U9341 (N_9341,N_9171,N_9028);
nor U9342 (N_9342,N_9009,N_9139);
nand U9343 (N_9343,N_9077,N_9011);
nor U9344 (N_9344,N_9199,N_9025);
nand U9345 (N_9345,N_9044,N_9147);
xnor U9346 (N_9346,N_9050,N_9138);
nor U9347 (N_9347,N_9171,N_9106);
nor U9348 (N_9348,N_9156,N_9058);
nor U9349 (N_9349,N_9174,N_9173);
or U9350 (N_9350,N_9117,N_9065);
or U9351 (N_9351,N_9047,N_9014);
and U9352 (N_9352,N_9061,N_9018);
nand U9353 (N_9353,N_9012,N_9096);
nand U9354 (N_9354,N_9169,N_9024);
nand U9355 (N_9355,N_9098,N_9197);
and U9356 (N_9356,N_9071,N_9185);
and U9357 (N_9357,N_9128,N_9074);
and U9358 (N_9358,N_9149,N_9167);
and U9359 (N_9359,N_9023,N_9017);
nor U9360 (N_9360,N_9097,N_9095);
xor U9361 (N_9361,N_9198,N_9191);
and U9362 (N_9362,N_9198,N_9174);
nor U9363 (N_9363,N_9070,N_9125);
and U9364 (N_9364,N_9016,N_9187);
or U9365 (N_9365,N_9050,N_9188);
or U9366 (N_9366,N_9122,N_9153);
xnor U9367 (N_9367,N_9101,N_9118);
and U9368 (N_9368,N_9157,N_9070);
and U9369 (N_9369,N_9058,N_9007);
and U9370 (N_9370,N_9117,N_9046);
and U9371 (N_9371,N_9102,N_9058);
nand U9372 (N_9372,N_9166,N_9050);
and U9373 (N_9373,N_9180,N_9087);
or U9374 (N_9374,N_9075,N_9089);
nor U9375 (N_9375,N_9005,N_9100);
xnor U9376 (N_9376,N_9138,N_9147);
nor U9377 (N_9377,N_9125,N_9115);
xnor U9378 (N_9378,N_9172,N_9117);
xnor U9379 (N_9379,N_9096,N_9155);
or U9380 (N_9380,N_9059,N_9007);
nor U9381 (N_9381,N_9016,N_9060);
and U9382 (N_9382,N_9081,N_9181);
nor U9383 (N_9383,N_9175,N_9191);
nor U9384 (N_9384,N_9174,N_9046);
and U9385 (N_9385,N_9103,N_9044);
or U9386 (N_9386,N_9147,N_9168);
and U9387 (N_9387,N_9188,N_9072);
and U9388 (N_9388,N_9056,N_9069);
or U9389 (N_9389,N_9160,N_9193);
or U9390 (N_9390,N_9078,N_9189);
nand U9391 (N_9391,N_9199,N_9131);
or U9392 (N_9392,N_9063,N_9021);
or U9393 (N_9393,N_9005,N_9072);
nand U9394 (N_9394,N_9000,N_9124);
or U9395 (N_9395,N_9163,N_9156);
xor U9396 (N_9396,N_9171,N_9006);
and U9397 (N_9397,N_9000,N_9054);
or U9398 (N_9398,N_9013,N_9140);
and U9399 (N_9399,N_9000,N_9197);
nand U9400 (N_9400,N_9383,N_9244);
nor U9401 (N_9401,N_9233,N_9391);
and U9402 (N_9402,N_9259,N_9350);
and U9403 (N_9403,N_9255,N_9281);
nor U9404 (N_9404,N_9396,N_9295);
or U9405 (N_9405,N_9330,N_9238);
or U9406 (N_9406,N_9333,N_9338);
nand U9407 (N_9407,N_9357,N_9326);
nand U9408 (N_9408,N_9279,N_9272);
xnor U9409 (N_9409,N_9215,N_9349);
nand U9410 (N_9410,N_9390,N_9247);
xor U9411 (N_9411,N_9271,N_9223);
or U9412 (N_9412,N_9206,N_9309);
nand U9413 (N_9413,N_9341,N_9353);
xor U9414 (N_9414,N_9200,N_9251);
or U9415 (N_9415,N_9228,N_9235);
and U9416 (N_9416,N_9297,N_9211);
nand U9417 (N_9417,N_9278,N_9313);
or U9418 (N_9418,N_9254,N_9242);
nor U9419 (N_9419,N_9340,N_9393);
and U9420 (N_9420,N_9336,N_9343);
or U9421 (N_9421,N_9241,N_9323);
xor U9422 (N_9422,N_9231,N_9319);
or U9423 (N_9423,N_9257,N_9377);
and U9424 (N_9424,N_9225,N_9214);
nor U9425 (N_9425,N_9335,N_9258);
or U9426 (N_9426,N_9370,N_9269);
and U9427 (N_9427,N_9266,N_9203);
nand U9428 (N_9428,N_9221,N_9290);
nand U9429 (N_9429,N_9380,N_9232);
nor U9430 (N_9430,N_9287,N_9366);
or U9431 (N_9431,N_9318,N_9372);
or U9432 (N_9432,N_9240,N_9360);
nor U9433 (N_9433,N_9212,N_9256);
xor U9434 (N_9434,N_9347,N_9358);
nor U9435 (N_9435,N_9219,N_9369);
nor U9436 (N_9436,N_9312,N_9220);
xnor U9437 (N_9437,N_9314,N_9374);
nand U9438 (N_9438,N_9344,N_9275);
nor U9439 (N_9439,N_9284,N_9315);
nand U9440 (N_9440,N_9261,N_9305);
nor U9441 (N_9441,N_9299,N_9389);
nor U9442 (N_9442,N_9302,N_9332);
and U9443 (N_9443,N_9252,N_9268);
nor U9444 (N_9444,N_9348,N_9253);
or U9445 (N_9445,N_9245,N_9294);
and U9446 (N_9446,N_9250,N_9216);
and U9447 (N_9447,N_9375,N_9243);
or U9448 (N_9448,N_9337,N_9345);
or U9449 (N_9449,N_9329,N_9361);
nor U9450 (N_9450,N_9381,N_9207);
or U9451 (N_9451,N_9288,N_9236);
nor U9452 (N_9452,N_9291,N_9386);
and U9453 (N_9453,N_9282,N_9267);
nor U9454 (N_9454,N_9384,N_9303);
nor U9455 (N_9455,N_9316,N_9289);
nand U9456 (N_9456,N_9246,N_9308);
nor U9457 (N_9457,N_9388,N_9224);
and U9458 (N_9458,N_9292,N_9382);
and U9459 (N_9459,N_9356,N_9234);
and U9460 (N_9460,N_9277,N_9300);
nand U9461 (N_9461,N_9296,N_9230);
nand U9462 (N_9462,N_9365,N_9210);
nor U9463 (N_9463,N_9229,N_9354);
nand U9464 (N_9464,N_9274,N_9368);
nand U9465 (N_9465,N_9227,N_9395);
nor U9466 (N_9466,N_9392,N_9276);
nand U9467 (N_9467,N_9248,N_9283);
or U9468 (N_9468,N_9398,N_9352);
nor U9469 (N_9469,N_9367,N_9311);
and U9470 (N_9470,N_9222,N_9325);
or U9471 (N_9471,N_9327,N_9273);
nor U9472 (N_9472,N_9218,N_9342);
nand U9473 (N_9473,N_9201,N_9237);
and U9474 (N_9474,N_9397,N_9208);
nor U9475 (N_9475,N_9293,N_9286);
or U9476 (N_9476,N_9331,N_9239);
xor U9477 (N_9477,N_9376,N_9378);
nand U9478 (N_9478,N_9394,N_9324);
nor U9479 (N_9479,N_9217,N_9209);
nor U9480 (N_9480,N_9285,N_9204);
and U9481 (N_9481,N_9310,N_9322);
or U9482 (N_9482,N_9298,N_9379);
nor U9483 (N_9483,N_9359,N_9351);
nand U9484 (N_9484,N_9263,N_9355);
nand U9485 (N_9485,N_9262,N_9280);
and U9486 (N_9486,N_9328,N_9249);
nor U9487 (N_9487,N_9264,N_9385);
and U9488 (N_9488,N_9265,N_9339);
nand U9489 (N_9489,N_9321,N_9205);
or U9490 (N_9490,N_9301,N_9306);
and U9491 (N_9491,N_9346,N_9387);
or U9492 (N_9492,N_9334,N_9371);
nor U9493 (N_9493,N_9213,N_9362);
or U9494 (N_9494,N_9364,N_9307);
nand U9495 (N_9495,N_9399,N_9363);
or U9496 (N_9496,N_9260,N_9304);
nand U9497 (N_9497,N_9373,N_9226);
and U9498 (N_9498,N_9270,N_9317);
or U9499 (N_9499,N_9202,N_9320);
nand U9500 (N_9500,N_9242,N_9394);
nand U9501 (N_9501,N_9289,N_9267);
nor U9502 (N_9502,N_9366,N_9362);
xor U9503 (N_9503,N_9212,N_9292);
nor U9504 (N_9504,N_9301,N_9335);
or U9505 (N_9505,N_9200,N_9280);
or U9506 (N_9506,N_9330,N_9225);
and U9507 (N_9507,N_9361,N_9330);
and U9508 (N_9508,N_9255,N_9216);
or U9509 (N_9509,N_9329,N_9233);
nor U9510 (N_9510,N_9267,N_9367);
and U9511 (N_9511,N_9268,N_9376);
nand U9512 (N_9512,N_9243,N_9209);
nand U9513 (N_9513,N_9261,N_9224);
or U9514 (N_9514,N_9384,N_9310);
or U9515 (N_9515,N_9226,N_9261);
and U9516 (N_9516,N_9203,N_9268);
nor U9517 (N_9517,N_9289,N_9209);
or U9518 (N_9518,N_9236,N_9320);
nor U9519 (N_9519,N_9243,N_9373);
or U9520 (N_9520,N_9390,N_9243);
nand U9521 (N_9521,N_9367,N_9242);
and U9522 (N_9522,N_9276,N_9343);
nor U9523 (N_9523,N_9223,N_9350);
nand U9524 (N_9524,N_9239,N_9284);
nand U9525 (N_9525,N_9370,N_9271);
nor U9526 (N_9526,N_9247,N_9375);
nor U9527 (N_9527,N_9398,N_9293);
nand U9528 (N_9528,N_9228,N_9290);
nor U9529 (N_9529,N_9385,N_9393);
or U9530 (N_9530,N_9330,N_9259);
or U9531 (N_9531,N_9295,N_9369);
nor U9532 (N_9532,N_9360,N_9325);
or U9533 (N_9533,N_9337,N_9325);
nor U9534 (N_9534,N_9228,N_9395);
or U9535 (N_9535,N_9322,N_9247);
nand U9536 (N_9536,N_9275,N_9365);
nor U9537 (N_9537,N_9251,N_9371);
and U9538 (N_9538,N_9228,N_9202);
nor U9539 (N_9539,N_9291,N_9264);
xnor U9540 (N_9540,N_9201,N_9211);
nor U9541 (N_9541,N_9341,N_9337);
or U9542 (N_9542,N_9208,N_9273);
or U9543 (N_9543,N_9234,N_9294);
and U9544 (N_9544,N_9300,N_9375);
nand U9545 (N_9545,N_9367,N_9286);
nor U9546 (N_9546,N_9329,N_9387);
or U9547 (N_9547,N_9368,N_9373);
xnor U9548 (N_9548,N_9287,N_9377);
nand U9549 (N_9549,N_9269,N_9314);
nor U9550 (N_9550,N_9235,N_9349);
or U9551 (N_9551,N_9338,N_9360);
or U9552 (N_9552,N_9354,N_9340);
nand U9553 (N_9553,N_9385,N_9386);
and U9554 (N_9554,N_9289,N_9328);
nor U9555 (N_9555,N_9289,N_9353);
and U9556 (N_9556,N_9307,N_9283);
nor U9557 (N_9557,N_9396,N_9382);
or U9558 (N_9558,N_9296,N_9286);
and U9559 (N_9559,N_9259,N_9224);
nor U9560 (N_9560,N_9221,N_9359);
and U9561 (N_9561,N_9290,N_9235);
nor U9562 (N_9562,N_9399,N_9325);
or U9563 (N_9563,N_9267,N_9321);
and U9564 (N_9564,N_9256,N_9249);
or U9565 (N_9565,N_9267,N_9279);
nor U9566 (N_9566,N_9242,N_9217);
or U9567 (N_9567,N_9268,N_9275);
and U9568 (N_9568,N_9378,N_9264);
xor U9569 (N_9569,N_9260,N_9363);
or U9570 (N_9570,N_9294,N_9270);
or U9571 (N_9571,N_9218,N_9387);
nand U9572 (N_9572,N_9339,N_9299);
or U9573 (N_9573,N_9271,N_9243);
and U9574 (N_9574,N_9221,N_9243);
or U9575 (N_9575,N_9245,N_9372);
nand U9576 (N_9576,N_9333,N_9287);
nor U9577 (N_9577,N_9287,N_9276);
and U9578 (N_9578,N_9374,N_9327);
or U9579 (N_9579,N_9233,N_9228);
nor U9580 (N_9580,N_9253,N_9219);
and U9581 (N_9581,N_9352,N_9300);
nand U9582 (N_9582,N_9291,N_9254);
or U9583 (N_9583,N_9294,N_9233);
nor U9584 (N_9584,N_9338,N_9276);
xor U9585 (N_9585,N_9202,N_9217);
xnor U9586 (N_9586,N_9206,N_9384);
nand U9587 (N_9587,N_9202,N_9307);
and U9588 (N_9588,N_9331,N_9246);
or U9589 (N_9589,N_9275,N_9238);
nor U9590 (N_9590,N_9357,N_9366);
nand U9591 (N_9591,N_9336,N_9303);
and U9592 (N_9592,N_9262,N_9354);
xnor U9593 (N_9593,N_9325,N_9209);
xor U9594 (N_9594,N_9350,N_9327);
nand U9595 (N_9595,N_9274,N_9221);
or U9596 (N_9596,N_9365,N_9314);
or U9597 (N_9597,N_9355,N_9309);
and U9598 (N_9598,N_9298,N_9234);
or U9599 (N_9599,N_9243,N_9366);
nor U9600 (N_9600,N_9477,N_9497);
nand U9601 (N_9601,N_9539,N_9418);
or U9602 (N_9602,N_9462,N_9408);
and U9603 (N_9603,N_9547,N_9435);
and U9604 (N_9604,N_9523,N_9470);
nor U9605 (N_9605,N_9426,N_9591);
and U9606 (N_9606,N_9583,N_9549);
nand U9607 (N_9607,N_9489,N_9402);
or U9608 (N_9608,N_9537,N_9444);
and U9609 (N_9609,N_9527,N_9595);
nor U9610 (N_9610,N_9585,N_9438);
xnor U9611 (N_9611,N_9479,N_9504);
nand U9612 (N_9612,N_9560,N_9453);
xor U9613 (N_9613,N_9581,N_9490);
or U9614 (N_9614,N_9498,N_9421);
or U9615 (N_9615,N_9545,N_9409);
xnor U9616 (N_9616,N_9534,N_9507);
nand U9617 (N_9617,N_9553,N_9599);
or U9618 (N_9618,N_9519,N_9546);
and U9619 (N_9619,N_9503,N_9562);
nand U9620 (N_9620,N_9405,N_9416);
xnor U9621 (N_9621,N_9428,N_9509);
or U9622 (N_9622,N_9411,N_9568);
or U9623 (N_9623,N_9434,N_9455);
or U9624 (N_9624,N_9563,N_9437);
or U9625 (N_9625,N_9517,N_9508);
nor U9626 (N_9626,N_9433,N_9541);
nor U9627 (N_9627,N_9430,N_9424);
or U9628 (N_9628,N_9513,N_9485);
and U9629 (N_9629,N_9447,N_9524);
or U9630 (N_9630,N_9557,N_9461);
nor U9631 (N_9631,N_9420,N_9594);
or U9632 (N_9632,N_9593,N_9448);
and U9633 (N_9633,N_9582,N_9528);
nand U9634 (N_9634,N_9456,N_9592);
nor U9635 (N_9635,N_9505,N_9464);
xnor U9636 (N_9636,N_9514,N_9400);
or U9637 (N_9637,N_9457,N_9445);
or U9638 (N_9638,N_9506,N_9484);
or U9639 (N_9639,N_9515,N_9413);
or U9640 (N_9640,N_9443,N_9414);
and U9641 (N_9641,N_9530,N_9551);
nor U9642 (N_9642,N_9531,N_9510);
xnor U9643 (N_9643,N_9440,N_9454);
and U9644 (N_9644,N_9425,N_9565);
or U9645 (N_9645,N_9441,N_9522);
or U9646 (N_9646,N_9422,N_9495);
and U9647 (N_9647,N_9406,N_9521);
and U9648 (N_9648,N_9431,N_9487);
or U9649 (N_9649,N_9597,N_9566);
xor U9650 (N_9650,N_9561,N_9478);
nor U9651 (N_9651,N_9575,N_9550);
or U9652 (N_9652,N_9476,N_9493);
nand U9653 (N_9653,N_9442,N_9542);
nand U9654 (N_9654,N_9589,N_9412);
or U9655 (N_9655,N_9452,N_9446);
nand U9656 (N_9656,N_9463,N_9427);
nor U9657 (N_9657,N_9459,N_9469);
or U9658 (N_9658,N_9450,N_9598);
or U9659 (N_9659,N_9483,N_9520);
nand U9660 (N_9660,N_9518,N_9574);
xor U9661 (N_9661,N_9587,N_9540);
and U9662 (N_9662,N_9410,N_9558);
or U9663 (N_9663,N_9492,N_9475);
and U9664 (N_9664,N_9584,N_9499);
nand U9665 (N_9665,N_9404,N_9525);
and U9666 (N_9666,N_9488,N_9576);
and U9667 (N_9667,N_9555,N_9596);
or U9668 (N_9668,N_9466,N_9407);
nand U9669 (N_9669,N_9544,N_9480);
and U9670 (N_9670,N_9559,N_9419);
xnor U9671 (N_9671,N_9468,N_9580);
nand U9672 (N_9672,N_9556,N_9588);
nand U9673 (N_9673,N_9482,N_9578);
nand U9674 (N_9674,N_9496,N_9533);
and U9675 (N_9675,N_9564,N_9512);
xor U9676 (N_9676,N_9465,N_9481);
nand U9677 (N_9677,N_9538,N_9429);
nor U9678 (N_9678,N_9532,N_9573);
nor U9679 (N_9679,N_9567,N_9494);
or U9680 (N_9680,N_9449,N_9526);
nand U9681 (N_9681,N_9577,N_9569);
nand U9682 (N_9682,N_9571,N_9586);
and U9683 (N_9683,N_9536,N_9460);
and U9684 (N_9684,N_9579,N_9516);
or U9685 (N_9685,N_9535,N_9423);
nor U9686 (N_9686,N_9417,N_9572);
or U9687 (N_9687,N_9474,N_9491);
xor U9688 (N_9688,N_9554,N_9458);
and U9689 (N_9689,N_9548,N_9590);
and U9690 (N_9690,N_9570,N_9436);
or U9691 (N_9691,N_9401,N_9486);
or U9692 (N_9692,N_9511,N_9552);
or U9693 (N_9693,N_9451,N_9501);
xor U9694 (N_9694,N_9502,N_9500);
nand U9695 (N_9695,N_9473,N_9472);
and U9696 (N_9696,N_9439,N_9432);
nor U9697 (N_9697,N_9543,N_9471);
or U9698 (N_9698,N_9467,N_9403);
xor U9699 (N_9699,N_9415,N_9529);
and U9700 (N_9700,N_9402,N_9593);
nand U9701 (N_9701,N_9426,N_9520);
and U9702 (N_9702,N_9585,N_9543);
nand U9703 (N_9703,N_9453,N_9563);
nand U9704 (N_9704,N_9571,N_9493);
nand U9705 (N_9705,N_9413,N_9451);
or U9706 (N_9706,N_9500,N_9572);
and U9707 (N_9707,N_9584,N_9526);
or U9708 (N_9708,N_9513,N_9425);
nor U9709 (N_9709,N_9430,N_9550);
or U9710 (N_9710,N_9461,N_9492);
or U9711 (N_9711,N_9566,N_9456);
nor U9712 (N_9712,N_9571,N_9415);
nor U9713 (N_9713,N_9580,N_9445);
xnor U9714 (N_9714,N_9598,N_9495);
or U9715 (N_9715,N_9404,N_9457);
nor U9716 (N_9716,N_9536,N_9459);
or U9717 (N_9717,N_9553,N_9416);
and U9718 (N_9718,N_9520,N_9501);
or U9719 (N_9719,N_9460,N_9487);
or U9720 (N_9720,N_9455,N_9413);
nor U9721 (N_9721,N_9462,N_9515);
nor U9722 (N_9722,N_9517,N_9473);
or U9723 (N_9723,N_9420,N_9568);
xor U9724 (N_9724,N_9505,N_9547);
nor U9725 (N_9725,N_9465,N_9487);
nand U9726 (N_9726,N_9545,N_9483);
and U9727 (N_9727,N_9440,N_9599);
and U9728 (N_9728,N_9440,N_9508);
and U9729 (N_9729,N_9478,N_9419);
and U9730 (N_9730,N_9503,N_9521);
nor U9731 (N_9731,N_9465,N_9511);
nand U9732 (N_9732,N_9556,N_9566);
nand U9733 (N_9733,N_9463,N_9552);
or U9734 (N_9734,N_9414,N_9425);
nand U9735 (N_9735,N_9568,N_9496);
nand U9736 (N_9736,N_9431,N_9531);
nand U9737 (N_9737,N_9412,N_9422);
nand U9738 (N_9738,N_9410,N_9509);
and U9739 (N_9739,N_9483,N_9413);
or U9740 (N_9740,N_9589,N_9484);
or U9741 (N_9741,N_9409,N_9483);
and U9742 (N_9742,N_9465,N_9401);
nor U9743 (N_9743,N_9498,N_9419);
nor U9744 (N_9744,N_9574,N_9577);
nor U9745 (N_9745,N_9534,N_9597);
or U9746 (N_9746,N_9599,N_9449);
and U9747 (N_9747,N_9598,N_9524);
nand U9748 (N_9748,N_9552,N_9568);
nor U9749 (N_9749,N_9540,N_9461);
and U9750 (N_9750,N_9513,N_9570);
xnor U9751 (N_9751,N_9572,N_9447);
xor U9752 (N_9752,N_9481,N_9555);
and U9753 (N_9753,N_9493,N_9475);
or U9754 (N_9754,N_9486,N_9499);
nand U9755 (N_9755,N_9533,N_9502);
nand U9756 (N_9756,N_9559,N_9561);
nor U9757 (N_9757,N_9403,N_9483);
or U9758 (N_9758,N_9590,N_9491);
xor U9759 (N_9759,N_9444,N_9404);
nor U9760 (N_9760,N_9519,N_9480);
and U9761 (N_9761,N_9428,N_9583);
or U9762 (N_9762,N_9560,N_9448);
and U9763 (N_9763,N_9549,N_9477);
or U9764 (N_9764,N_9523,N_9464);
nor U9765 (N_9765,N_9457,N_9534);
nor U9766 (N_9766,N_9569,N_9579);
xnor U9767 (N_9767,N_9493,N_9450);
nand U9768 (N_9768,N_9504,N_9543);
nor U9769 (N_9769,N_9414,N_9483);
nor U9770 (N_9770,N_9591,N_9549);
xor U9771 (N_9771,N_9405,N_9571);
nor U9772 (N_9772,N_9475,N_9433);
nor U9773 (N_9773,N_9565,N_9584);
and U9774 (N_9774,N_9520,N_9406);
and U9775 (N_9775,N_9428,N_9573);
and U9776 (N_9776,N_9545,N_9538);
or U9777 (N_9777,N_9420,N_9477);
nand U9778 (N_9778,N_9407,N_9468);
nor U9779 (N_9779,N_9447,N_9543);
nand U9780 (N_9780,N_9443,N_9566);
and U9781 (N_9781,N_9482,N_9542);
or U9782 (N_9782,N_9487,N_9569);
nand U9783 (N_9783,N_9435,N_9529);
and U9784 (N_9784,N_9564,N_9553);
xnor U9785 (N_9785,N_9503,N_9573);
or U9786 (N_9786,N_9566,N_9590);
and U9787 (N_9787,N_9589,N_9523);
nand U9788 (N_9788,N_9414,N_9481);
and U9789 (N_9789,N_9554,N_9468);
xor U9790 (N_9790,N_9403,N_9419);
and U9791 (N_9791,N_9526,N_9414);
and U9792 (N_9792,N_9482,N_9493);
or U9793 (N_9793,N_9585,N_9450);
or U9794 (N_9794,N_9491,N_9444);
and U9795 (N_9795,N_9523,N_9501);
xor U9796 (N_9796,N_9540,N_9513);
and U9797 (N_9797,N_9464,N_9590);
nor U9798 (N_9798,N_9423,N_9552);
nand U9799 (N_9799,N_9433,N_9427);
nor U9800 (N_9800,N_9716,N_9728);
or U9801 (N_9801,N_9726,N_9612);
nor U9802 (N_9802,N_9784,N_9712);
or U9803 (N_9803,N_9686,N_9794);
nand U9804 (N_9804,N_9654,N_9638);
nand U9805 (N_9805,N_9600,N_9697);
nor U9806 (N_9806,N_9674,N_9744);
nand U9807 (N_9807,N_9700,N_9608);
or U9808 (N_9808,N_9771,N_9785);
and U9809 (N_9809,N_9635,N_9657);
or U9810 (N_9810,N_9611,N_9756);
and U9811 (N_9811,N_9607,N_9609);
nor U9812 (N_9812,N_9768,N_9779);
or U9813 (N_9813,N_9725,N_9737);
nor U9814 (N_9814,N_9741,N_9732);
nand U9815 (N_9815,N_9798,N_9621);
nor U9816 (N_9816,N_9791,N_9778);
xor U9817 (N_9817,N_9776,N_9708);
nand U9818 (N_9818,N_9619,N_9618);
xor U9819 (N_9819,N_9636,N_9615);
nor U9820 (N_9820,N_9671,N_9706);
and U9821 (N_9821,N_9714,N_9705);
xor U9822 (N_9822,N_9695,N_9665);
nor U9823 (N_9823,N_9722,N_9675);
and U9824 (N_9824,N_9724,N_9682);
and U9825 (N_9825,N_9614,N_9684);
and U9826 (N_9826,N_9797,N_9662);
nand U9827 (N_9827,N_9777,N_9749);
and U9828 (N_9828,N_9641,N_9625);
or U9829 (N_9829,N_9666,N_9623);
xor U9830 (N_9830,N_9775,N_9759);
nor U9831 (N_9831,N_9670,N_9651);
nand U9832 (N_9832,N_9783,N_9742);
nand U9833 (N_9833,N_9796,N_9605);
or U9834 (N_9834,N_9650,N_9613);
xor U9835 (N_9835,N_9626,N_9703);
xnor U9836 (N_9836,N_9720,N_9718);
nor U9837 (N_9837,N_9751,N_9753);
or U9838 (N_9838,N_9743,N_9734);
nand U9839 (N_9839,N_9745,N_9750);
xnor U9840 (N_9840,N_9669,N_9663);
nand U9841 (N_9841,N_9680,N_9606);
or U9842 (N_9842,N_9661,N_9693);
nand U9843 (N_9843,N_9761,N_9676);
nand U9844 (N_9844,N_9793,N_9601);
and U9845 (N_9845,N_9685,N_9748);
nor U9846 (N_9846,N_9723,N_9755);
and U9847 (N_9847,N_9770,N_9766);
nand U9848 (N_9848,N_9640,N_9648);
nand U9849 (N_9849,N_9790,N_9781);
or U9850 (N_9850,N_9692,N_9704);
and U9851 (N_9851,N_9795,N_9707);
and U9852 (N_9852,N_9696,N_9788);
nor U9853 (N_9853,N_9717,N_9653);
nand U9854 (N_9854,N_9645,N_9763);
or U9855 (N_9855,N_9735,N_9736);
and U9856 (N_9856,N_9715,N_9644);
or U9857 (N_9857,N_9780,N_9721);
nor U9858 (N_9858,N_9627,N_9694);
nor U9859 (N_9859,N_9729,N_9760);
or U9860 (N_9860,N_9639,N_9698);
nor U9861 (N_9861,N_9632,N_9667);
nand U9862 (N_9862,N_9604,N_9690);
or U9863 (N_9863,N_9634,N_9799);
or U9864 (N_9864,N_9792,N_9655);
and U9865 (N_9865,N_9758,N_9767);
or U9866 (N_9866,N_9649,N_9711);
and U9867 (N_9867,N_9789,N_9643);
nand U9868 (N_9868,N_9691,N_9658);
and U9869 (N_9869,N_9746,N_9630);
nand U9870 (N_9870,N_9774,N_9687);
or U9871 (N_9871,N_9660,N_9629);
nor U9872 (N_9872,N_9701,N_9659);
nand U9873 (N_9873,N_9622,N_9664);
nand U9874 (N_9874,N_9769,N_9620);
and U9875 (N_9875,N_9754,N_9709);
or U9876 (N_9876,N_9731,N_9652);
and U9877 (N_9877,N_9610,N_9673);
and U9878 (N_9878,N_9762,N_9699);
nand U9879 (N_9879,N_9727,N_9668);
nand U9880 (N_9880,N_9656,N_9677);
nor U9881 (N_9881,N_9757,N_9739);
and U9882 (N_9882,N_9738,N_9679);
nand U9883 (N_9883,N_9787,N_9782);
and U9884 (N_9884,N_9772,N_9764);
or U9885 (N_9885,N_9733,N_9672);
nor U9886 (N_9886,N_9681,N_9631);
or U9887 (N_9887,N_9642,N_9710);
and U9888 (N_9888,N_9752,N_9683);
nor U9889 (N_9889,N_9719,N_9773);
xnor U9890 (N_9890,N_9617,N_9628);
and U9891 (N_9891,N_9647,N_9689);
and U9892 (N_9892,N_9786,N_9633);
or U9893 (N_9893,N_9702,N_9624);
and U9894 (N_9894,N_9730,N_9713);
and U9895 (N_9895,N_9765,N_9678);
nor U9896 (N_9896,N_9688,N_9603);
nand U9897 (N_9897,N_9646,N_9616);
nand U9898 (N_9898,N_9602,N_9637);
or U9899 (N_9899,N_9747,N_9740);
or U9900 (N_9900,N_9605,N_9672);
nand U9901 (N_9901,N_9728,N_9721);
nand U9902 (N_9902,N_9732,N_9776);
or U9903 (N_9903,N_9755,N_9779);
nand U9904 (N_9904,N_9617,N_9690);
nand U9905 (N_9905,N_9738,N_9762);
nor U9906 (N_9906,N_9799,N_9692);
nand U9907 (N_9907,N_9670,N_9732);
and U9908 (N_9908,N_9651,N_9623);
and U9909 (N_9909,N_9651,N_9790);
and U9910 (N_9910,N_9715,N_9626);
and U9911 (N_9911,N_9728,N_9723);
nor U9912 (N_9912,N_9746,N_9622);
and U9913 (N_9913,N_9760,N_9712);
or U9914 (N_9914,N_9713,N_9732);
nor U9915 (N_9915,N_9633,N_9788);
or U9916 (N_9916,N_9628,N_9741);
xnor U9917 (N_9917,N_9623,N_9773);
or U9918 (N_9918,N_9618,N_9650);
and U9919 (N_9919,N_9665,N_9757);
and U9920 (N_9920,N_9613,N_9664);
nand U9921 (N_9921,N_9626,N_9681);
and U9922 (N_9922,N_9635,N_9660);
and U9923 (N_9923,N_9661,N_9674);
nor U9924 (N_9924,N_9639,N_9697);
or U9925 (N_9925,N_9636,N_9651);
nor U9926 (N_9926,N_9629,N_9783);
nor U9927 (N_9927,N_9702,N_9731);
nand U9928 (N_9928,N_9647,N_9675);
nand U9929 (N_9929,N_9635,N_9636);
nand U9930 (N_9930,N_9649,N_9724);
or U9931 (N_9931,N_9610,N_9758);
and U9932 (N_9932,N_9680,N_9783);
and U9933 (N_9933,N_9670,N_9784);
nor U9934 (N_9934,N_9767,N_9653);
or U9935 (N_9935,N_9739,N_9614);
xor U9936 (N_9936,N_9759,N_9662);
or U9937 (N_9937,N_9783,N_9723);
or U9938 (N_9938,N_9726,N_9775);
nand U9939 (N_9939,N_9740,N_9636);
and U9940 (N_9940,N_9637,N_9707);
xor U9941 (N_9941,N_9643,N_9707);
or U9942 (N_9942,N_9779,N_9665);
and U9943 (N_9943,N_9711,N_9776);
nor U9944 (N_9944,N_9734,N_9607);
nand U9945 (N_9945,N_9635,N_9639);
nor U9946 (N_9946,N_9778,N_9632);
and U9947 (N_9947,N_9772,N_9616);
nand U9948 (N_9948,N_9620,N_9779);
or U9949 (N_9949,N_9685,N_9660);
xnor U9950 (N_9950,N_9699,N_9722);
nor U9951 (N_9951,N_9625,N_9753);
nor U9952 (N_9952,N_9712,N_9680);
and U9953 (N_9953,N_9694,N_9735);
or U9954 (N_9954,N_9651,N_9615);
nand U9955 (N_9955,N_9707,N_9679);
nor U9956 (N_9956,N_9753,N_9717);
nor U9957 (N_9957,N_9720,N_9790);
nor U9958 (N_9958,N_9632,N_9630);
or U9959 (N_9959,N_9622,N_9683);
and U9960 (N_9960,N_9728,N_9738);
nor U9961 (N_9961,N_9779,N_9684);
and U9962 (N_9962,N_9766,N_9769);
or U9963 (N_9963,N_9740,N_9715);
nor U9964 (N_9964,N_9621,N_9601);
nor U9965 (N_9965,N_9631,N_9669);
nand U9966 (N_9966,N_9790,N_9751);
and U9967 (N_9967,N_9759,N_9796);
and U9968 (N_9968,N_9713,N_9767);
and U9969 (N_9969,N_9743,N_9703);
or U9970 (N_9970,N_9671,N_9745);
or U9971 (N_9971,N_9707,N_9793);
xor U9972 (N_9972,N_9779,N_9788);
and U9973 (N_9973,N_9766,N_9717);
nor U9974 (N_9974,N_9673,N_9749);
or U9975 (N_9975,N_9766,N_9646);
xnor U9976 (N_9976,N_9618,N_9694);
nor U9977 (N_9977,N_9686,N_9684);
nor U9978 (N_9978,N_9726,N_9671);
and U9979 (N_9979,N_9708,N_9686);
nor U9980 (N_9980,N_9666,N_9681);
and U9981 (N_9981,N_9731,N_9693);
and U9982 (N_9982,N_9765,N_9626);
nand U9983 (N_9983,N_9738,N_9773);
and U9984 (N_9984,N_9733,N_9624);
nor U9985 (N_9985,N_9694,N_9679);
xnor U9986 (N_9986,N_9681,N_9660);
xnor U9987 (N_9987,N_9767,N_9749);
and U9988 (N_9988,N_9638,N_9647);
nand U9989 (N_9989,N_9793,N_9652);
or U9990 (N_9990,N_9788,N_9684);
xor U9991 (N_9991,N_9656,N_9601);
nor U9992 (N_9992,N_9645,N_9655);
nor U9993 (N_9993,N_9630,N_9667);
xnor U9994 (N_9994,N_9780,N_9795);
nand U9995 (N_9995,N_9778,N_9642);
or U9996 (N_9996,N_9681,N_9735);
nor U9997 (N_9997,N_9702,N_9733);
or U9998 (N_9998,N_9691,N_9776);
xnor U9999 (N_9999,N_9639,N_9714);
or UO_0 (O_0,N_9893,N_9994);
and UO_1 (O_1,N_9972,N_9882);
nand UO_2 (O_2,N_9896,N_9951);
nor UO_3 (O_3,N_9849,N_9886);
nand UO_4 (O_4,N_9906,N_9862);
nor UO_5 (O_5,N_9873,N_9954);
xnor UO_6 (O_6,N_9913,N_9923);
nor UO_7 (O_7,N_9991,N_9957);
nand UO_8 (O_8,N_9993,N_9979);
nor UO_9 (O_9,N_9949,N_9945);
or UO_10 (O_10,N_9952,N_9915);
and UO_11 (O_11,N_9897,N_9927);
and UO_12 (O_12,N_9956,N_9961);
nand UO_13 (O_13,N_9844,N_9816);
or UO_14 (O_14,N_9801,N_9872);
nand UO_15 (O_15,N_9982,N_9924);
and UO_16 (O_16,N_9988,N_9852);
or UO_17 (O_17,N_9825,N_9970);
nand UO_18 (O_18,N_9997,N_9854);
xnor UO_19 (O_19,N_9916,N_9880);
nor UO_20 (O_20,N_9920,N_9863);
or UO_21 (O_21,N_9909,N_9936);
nor UO_22 (O_22,N_9941,N_9912);
nand UO_23 (O_23,N_9937,N_9884);
nand UO_24 (O_24,N_9855,N_9901);
or UO_25 (O_25,N_9881,N_9898);
xor UO_26 (O_26,N_9865,N_9959);
or UO_27 (O_27,N_9958,N_9889);
and UO_28 (O_28,N_9966,N_9831);
or UO_29 (O_29,N_9903,N_9823);
nor UO_30 (O_30,N_9826,N_9877);
and UO_31 (O_31,N_9996,N_9984);
nor UO_32 (O_32,N_9907,N_9942);
nor UO_33 (O_33,N_9931,N_9803);
and UO_34 (O_34,N_9960,N_9832);
or UO_35 (O_35,N_9922,N_9870);
nor UO_36 (O_36,N_9814,N_9928);
nand UO_37 (O_37,N_9890,N_9861);
or UO_38 (O_38,N_9919,N_9910);
nand UO_39 (O_39,N_9895,N_9995);
nand UO_40 (O_40,N_9947,N_9847);
nor UO_41 (O_41,N_9977,N_9869);
nor UO_42 (O_42,N_9804,N_9841);
nand UO_43 (O_43,N_9967,N_9867);
nor UO_44 (O_44,N_9811,N_9953);
and UO_45 (O_45,N_9874,N_9858);
nor UO_46 (O_46,N_9899,N_9808);
nand UO_47 (O_47,N_9815,N_9948);
nor UO_48 (O_48,N_9836,N_9879);
nand UO_49 (O_49,N_9838,N_9932);
nand UO_50 (O_50,N_9935,N_9914);
nand UO_51 (O_51,N_9926,N_9868);
or UO_52 (O_52,N_9859,N_9888);
nor UO_53 (O_53,N_9835,N_9843);
xnor UO_54 (O_54,N_9946,N_9908);
or UO_55 (O_55,N_9990,N_9817);
and UO_56 (O_56,N_9851,N_9940);
or UO_57 (O_57,N_9998,N_9891);
nor UO_58 (O_58,N_9860,N_9864);
nor UO_59 (O_59,N_9921,N_9819);
and UO_60 (O_60,N_9813,N_9837);
and UO_61 (O_61,N_9800,N_9939);
xor UO_62 (O_62,N_9878,N_9887);
nand UO_63 (O_63,N_9812,N_9976);
or UO_64 (O_64,N_9980,N_9856);
and UO_65 (O_65,N_9840,N_9969);
nand UO_66 (O_66,N_9974,N_9938);
nor UO_67 (O_67,N_9999,N_9929);
and UO_68 (O_68,N_9930,N_9845);
and UO_69 (O_69,N_9934,N_9950);
nor UO_70 (O_70,N_9985,N_9883);
and UO_71 (O_71,N_9986,N_9821);
or UO_72 (O_72,N_9802,N_9902);
or UO_73 (O_73,N_9871,N_9992);
or UO_74 (O_74,N_9978,N_9827);
nor UO_75 (O_75,N_9820,N_9943);
and UO_76 (O_76,N_9833,N_9866);
nand UO_77 (O_77,N_9809,N_9964);
nand UO_78 (O_78,N_9830,N_9981);
nand UO_79 (O_79,N_9822,N_9857);
and UO_80 (O_80,N_9824,N_9839);
xor UO_81 (O_81,N_9963,N_9846);
nor UO_82 (O_82,N_9829,N_9989);
nor UO_83 (O_83,N_9892,N_9876);
nand UO_84 (O_84,N_9885,N_9828);
nand UO_85 (O_85,N_9917,N_9894);
nor UO_86 (O_86,N_9944,N_9962);
and UO_87 (O_87,N_9810,N_9900);
nand UO_88 (O_88,N_9975,N_9983);
and UO_89 (O_89,N_9918,N_9973);
or UO_90 (O_90,N_9818,N_9875);
nor UO_91 (O_91,N_9955,N_9925);
nor UO_92 (O_92,N_9905,N_9807);
nand UO_93 (O_93,N_9911,N_9933);
or UO_94 (O_94,N_9805,N_9987);
nand UO_95 (O_95,N_9965,N_9971);
nand UO_96 (O_96,N_9834,N_9848);
nand UO_97 (O_97,N_9853,N_9850);
and UO_98 (O_98,N_9968,N_9842);
nand UO_99 (O_99,N_9904,N_9806);
or UO_100 (O_100,N_9808,N_9970);
and UO_101 (O_101,N_9832,N_9913);
or UO_102 (O_102,N_9909,N_9913);
nor UO_103 (O_103,N_9889,N_9924);
or UO_104 (O_104,N_9839,N_9991);
nor UO_105 (O_105,N_9974,N_9843);
or UO_106 (O_106,N_9861,N_9885);
and UO_107 (O_107,N_9806,N_9853);
and UO_108 (O_108,N_9812,N_9934);
or UO_109 (O_109,N_9941,N_9945);
nand UO_110 (O_110,N_9840,N_9872);
and UO_111 (O_111,N_9828,N_9865);
nor UO_112 (O_112,N_9851,N_9888);
or UO_113 (O_113,N_9824,N_9985);
nand UO_114 (O_114,N_9848,N_9999);
and UO_115 (O_115,N_9802,N_9976);
or UO_116 (O_116,N_9845,N_9896);
and UO_117 (O_117,N_9959,N_9926);
xnor UO_118 (O_118,N_9920,N_9862);
nand UO_119 (O_119,N_9832,N_9978);
xor UO_120 (O_120,N_9851,N_9924);
nand UO_121 (O_121,N_9946,N_9846);
nand UO_122 (O_122,N_9889,N_9850);
nor UO_123 (O_123,N_9937,N_9928);
nand UO_124 (O_124,N_9903,N_9837);
or UO_125 (O_125,N_9899,N_9823);
or UO_126 (O_126,N_9920,N_9841);
or UO_127 (O_127,N_9913,N_9853);
nor UO_128 (O_128,N_9995,N_9912);
and UO_129 (O_129,N_9883,N_9921);
or UO_130 (O_130,N_9926,N_9931);
nor UO_131 (O_131,N_9852,N_9842);
and UO_132 (O_132,N_9957,N_9814);
or UO_133 (O_133,N_9838,N_9825);
nand UO_134 (O_134,N_9956,N_9896);
nor UO_135 (O_135,N_9939,N_9840);
nand UO_136 (O_136,N_9866,N_9950);
and UO_137 (O_137,N_9864,N_9831);
and UO_138 (O_138,N_9966,N_9990);
and UO_139 (O_139,N_9823,N_9830);
and UO_140 (O_140,N_9812,N_9826);
nand UO_141 (O_141,N_9878,N_9926);
xnor UO_142 (O_142,N_9985,N_9809);
nand UO_143 (O_143,N_9883,N_9849);
or UO_144 (O_144,N_9956,N_9826);
xor UO_145 (O_145,N_9887,N_9957);
and UO_146 (O_146,N_9939,N_9907);
and UO_147 (O_147,N_9858,N_9867);
nor UO_148 (O_148,N_9977,N_9905);
nor UO_149 (O_149,N_9801,N_9882);
and UO_150 (O_150,N_9889,N_9925);
nand UO_151 (O_151,N_9920,N_9909);
nand UO_152 (O_152,N_9890,N_9866);
and UO_153 (O_153,N_9888,N_9810);
nor UO_154 (O_154,N_9929,N_9851);
nand UO_155 (O_155,N_9946,N_9975);
and UO_156 (O_156,N_9923,N_9962);
nor UO_157 (O_157,N_9822,N_9978);
or UO_158 (O_158,N_9892,N_9896);
and UO_159 (O_159,N_9860,N_9964);
nand UO_160 (O_160,N_9849,N_9828);
nand UO_161 (O_161,N_9857,N_9890);
nor UO_162 (O_162,N_9995,N_9873);
xor UO_163 (O_163,N_9899,N_9834);
or UO_164 (O_164,N_9862,N_9852);
or UO_165 (O_165,N_9949,N_9964);
or UO_166 (O_166,N_9904,N_9983);
or UO_167 (O_167,N_9903,N_9855);
nor UO_168 (O_168,N_9826,N_9878);
or UO_169 (O_169,N_9844,N_9988);
or UO_170 (O_170,N_9852,N_9830);
nand UO_171 (O_171,N_9866,N_9904);
and UO_172 (O_172,N_9973,N_9943);
and UO_173 (O_173,N_9924,N_9886);
and UO_174 (O_174,N_9906,N_9801);
nand UO_175 (O_175,N_9875,N_9939);
nor UO_176 (O_176,N_9987,N_9819);
or UO_177 (O_177,N_9814,N_9917);
nor UO_178 (O_178,N_9942,N_9951);
or UO_179 (O_179,N_9953,N_9861);
xnor UO_180 (O_180,N_9874,N_9913);
nand UO_181 (O_181,N_9826,N_9833);
nor UO_182 (O_182,N_9870,N_9914);
and UO_183 (O_183,N_9937,N_9995);
or UO_184 (O_184,N_9920,N_9823);
nand UO_185 (O_185,N_9855,N_9956);
and UO_186 (O_186,N_9932,N_9935);
xor UO_187 (O_187,N_9902,N_9978);
nand UO_188 (O_188,N_9912,N_9826);
nor UO_189 (O_189,N_9965,N_9960);
and UO_190 (O_190,N_9968,N_9941);
and UO_191 (O_191,N_9973,N_9993);
nand UO_192 (O_192,N_9835,N_9955);
or UO_193 (O_193,N_9857,N_9988);
and UO_194 (O_194,N_9951,N_9918);
and UO_195 (O_195,N_9830,N_9991);
xnor UO_196 (O_196,N_9997,N_9882);
or UO_197 (O_197,N_9882,N_9906);
or UO_198 (O_198,N_9931,N_9873);
or UO_199 (O_199,N_9988,N_9865);
or UO_200 (O_200,N_9865,N_9878);
nor UO_201 (O_201,N_9887,N_9868);
nand UO_202 (O_202,N_9864,N_9857);
nor UO_203 (O_203,N_9962,N_9981);
or UO_204 (O_204,N_9920,N_9964);
nor UO_205 (O_205,N_9877,N_9812);
xor UO_206 (O_206,N_9943,N_9859);
or UO_207 (O_207,N_9861,N_9945);
xor UO_208 (O_208,N_9857,N_9894);
nor UO_209 (O_209,N_9816,N_9914);
and UO_210 (O_210,N_9810,N_9856);
nand UO_211 (O_211,N_9854,N_9963);
nand UO_212 (O_212,N_9833,N_9888);
or UO_213 (O_213,N_9905,N_9863);
nand UO_214 (O_214,N_9817,N_9898);
xnor UO_215 (O_215,N_9838,N_9806);
nor UO_216 (O_216,N_9891,N_9941);
and UO_217 (O_217,N_9873,N_9906);
and UO_218 (O_218,N_9960,N_9822);
nand UO_219 (O_219,N_9948,N_9859);
nand UO_220 (O_220,N_9962,N_9992);
or UO_221 (O_221,N_9957,N_9899);
nor UO_222 (O_222,N_9939,N_9813);
xnor UO_223 (O_223,N_9896,N_9905);
nor UO_224 (O_224,N_9882,N_9862);
and UO_225 (O_225,N_9842,N_9803);
or UO_226 (O_226,N_9955,N_9951);
and UO_227 (O_227,N_9872,N_9933);
nand UO_228 (O_228,N_9812,N_9971);
nand UO_229 (O_229,N_9802,N_9914);
and UO_230 (O_230,N_9858,N_9814);
nor UO_231 (O_231,N_9979,N_9972);
nor UO_232 (O_232,N_9859,N_9923);
and UO_233 (O_233,N_9961,N_9948);
nand UO_234 (O_234,N_9839,N_9884);
and UO_235 (O_235,N_9872,N_9810);
nand UO_236 (O_236,N_9869,N_9836);
and UO_237 (O_237,N_9808,N_9923);
nor UO_238 (O_238,N_9945,N_9852);
or UO_239 (O_239,N_9927,N_9968);
xnor UO_240 (O_240,N_9967,N_9864);
or UO_241 (O_241,N_9939,N_9977);
or UO_242 (O_242,N_9943,N_9858);
nor UO_243 (O_243,N_9901,N_9933);
nor UO_244 (O_244,N_9919,N_9951);
and UO_245 (O_245,N_9913,N_9846);
or UO_246 (O_246,N_9827,N_9903);
nor UO_247 (O_247,N_9927,N_9857);
or UO_248 (O_248,N_9925,N_9834);
nand UO_249 (O_249,N_9878,N_9961);
nand UO_250 (O_250,N_9959,N_9929);
or UO_251 (O_251,N_9905,N_9825);
and UO_252 (O_252,N_9822,N_9889);
and UO_253 (O_253,N_9905,N_9982);
xnor UO_254 (O_254,N_9850,N_9962);
nand UO_255 (O_255,N_9842,N_9958);
nor UO_256 (O_256,N_9861,N_9888);
xor UO_257 (O_257,N_9927,N_9830);
or UO_258 (O_258,N_9980,N_9940);
and UO_259 (O_259,N_9940,N_9868);
nand UO_260 (O_260,N_9933,N_9950);
and UO_261 (O_261,N_9859,N_9919);
or UO_262 (O_262,N_9996,N_9805);
nor UO_263 (O_263,N_9841,N_9955);
or UO_264 (O_264,N_9827,N_9830);
nor UO_265 (O_265,N_9818,N_9978);
and UO_266 (O_266,N_9839,N_9987);
nand UO_267 (O_267,N_9937,N_9914);
and UO_268 (O_268,N_9919,N_9841);
nand UO_269 (O_269,N_9908,N_9984);
and UO_270 (O_270,N_9984,N_9945);
xnor UO_271 (O_271,N_9951,N_9884);
or UO_272 (O_272,N_9915,N_9992);
nor UO_273 (O_273,N_9827,N_9817);
and UO_274 (O_274,N_9812,N_9840);
and UO_275 (O_275,N_9973,N_9850);
or UO_276 (O_276,N_9801,N_9854);
xor UO_277 (O_277,N_9883,N_9881);
and UO_278 (O_278,N_9825,N_9885);
or UO_279 (O_279,N_9910,N_9932);
or UO_280 (O_280,N_9823,N_9866);
xor UO_281 (O_281,N_9888,N_9900);
nor UO_282 (O_282,N_9968,N_9959);
xor UO_283 (O_283,N_9842,N_9881);
nand UO_284 (O_284,N_9803,N_9960);
and UO_285 (O_285,N_9998,N_9840);
nor UO_286 (O_286,N_9823,N_9977);
xor UO_287 (O_287,N_9973,N_9951);
or UO_288 (O_288,N_9962,N_9862);
xor UO_289 (O_289,N_9922,N_9832);
nand UO_290 (O_290,N_9957,N_9976);
nand UO_291 (O_291,N_9846,N_9929);
xnor UO_292 (O_292,N_9947,N_9910);
nor UO_293 (O_293,N_9959,N_9978);
and UO_294 (O_294,N_9864,N_9992);
xor UO_295 (O_295,N_9969,N_9865);
or UO_296 (O_296,N_9959,N_9821);
nor UO_297 (O_297,N_9921,N_9836);
xnor UO_298 (O_298,N_9836,N_9827);
or UO_299 (O_299,N_9846,N_9899);
and UO_300 (O_300,N_9886,N_9819);
and UO_301 (O_301,N_9940,N_9820);
and UO_302 (O_302,N_9822,N_9957);
nor UO_303 (O_303,N_9923,N_9902);
or UO_304 (O_304,N_9849,N_9877);
or UO_305 (O_305,N_9874,N_9942);
or UO_306 (O_306,N_9990,N_9803);
and UO_307 (O_307,N_9857,N_9972);
nor UO_308 (O_308,N_9968,N_9954);
xor UO_309 (O_309,N_9963,N_9806);
or UO_310 (O_310,N_9912,N_9886);
or UO_311 (O_311,N_9952,N_9817);
nand UO_312 (O_312,N_9907,N_9976);
or UO_313 (O_313,N_9889,N_9997);
nand UO_314 (O_314,N_9806,N_9973);
nand UO_315 (O_315,N_9845,N_9944);
nand UO_316 (O_316,N_9836,N_9989);
or UO_317 (O_317,N_9859,N_9946);
and UO_318 (O_318,N_9939,N_9956);
nor UO_319 (O_319,N_9933,N_9894);
nand UO_320 (O_320,N_9883,N_9908);
or UO_321 (O_321,N_9852,N_9993);
and UO_322 (O_322,N_9992,N_9942);
or UO_323 (O_323,N_9917,N_9925);
and UO_324 (O_324,N_9821,N_9999);
or UO_325 (O_325,N_9940,N_9972);
xnor UO_326 (O_326,N_9812,N_9994);
nor UO_327 (O_327,N_9908,N_9903);
nand UO_328 (O_328,N_9819,N_9941);
and UO_329 (O_329,N_9892,N_9848);
and UO_330 (O_330,N_9957,N_9924);
nand UO_331 (O_331,N_9873,N_9974);
or UO_332 (O_332,N_9988,N_9866);
and UO_333 (O_333,N_9835,N_9839);
nor UO_334 (O_334,N_9914,N_9846);
nor UO_335 (O_335,N_9917,N_9885);
and UO_336 (O_336,N_9910,N_9840);
nand UO_337 (O_337,N_9882,N_9831);
nand UO_338 (O_338,N_9844,N_9913);
or UO_339 (O_339,N_9871,N_9976);
nand UO_340 (O_340,N_9835,N_9892);
nor UO_341 (O_341,N_9953,N_9852);
nor UO_342 (O_342,N_9865,N_9912);
nand UO_343 (O_343,N_9821,N_9939);
nand UO_344 (O_344,N_9894,N_9948);
xnor UO_345 (O_345,N_9866,N_9940);
xor UO_346 (O_346,N_9999,N_9918);
and UO_347 (O_347,N_9863,N_9882);
xnor UO_348 (O_348,N_9971,N_9946);
nand UO_349 (O_349,N_9942,N_9860);
nor UO_350 (O_350,N_9871,N_9950);
nor UO_351 (O_351,N_9941,N_9905);
nand UO_352 (O_352,N_9887,N_9856);
and UO_353 (O_353,N_9870,N_9987);
or UO_354 (O_354,N_9806,N_9881);
nor UO_355 (O_355,N_9896,N_9996);
nor UO_356 (O_356,N_9908,N_9844);
nand UO_357 (O_357,N_9942,N_9933);
nor UO_358 (O_358,N_9816,N_9884);
nor UO_359 (O_359,N_9806,N_9941);
or UO_360 (O_360,N_9946,N_9944);
nand UO_361 (O_361,N_9801,N_9822);
xor UO_362 (O_362,N_9998,N_9959);
or UO_363 (O_363,N_9812,N_9913);
nand UO_364 (O_364,N_9814,N_9919);
nor UO_365 (O_365,N_9884,N_9835);
and UO_366 (O_366,N_9910,N_9887);
nor UO_367 (O_367,N_9906,N_9805);
and UO_368 (O_368,N_9845,N_9897);
and UO_369 (O_369,N_9881,N_9965);
or UO_370 (O_370,N_9809,N_9956);
nand UO_371 (O_371,N_9952,N_9950);
or UO_372 (O_372,N_9891,N_9904);
or UO_373 (O_373,N_9913,N_9982);
and UO_374 (O_374,N_9988,N_9973);
xor UO_375 (O_375,N_9992,N_9826);
nand UO_376 (O_376,N_9868,N_9880);
xor UO_377 (O_377,N_9971,N_9917);
and UO_378 (O_378,N_9890,N_9805);
nand UO_379 (O_379,N_9951,N_9975);
nand UO_380 (O_380,N_9958,N_9831);
and UO_381 (O_381,N_9912,N_9874);
nand UO_382 (O_382,N_9876,N_9930);
nor UO_383 (O_383,N_9889,N_9968);
and UO_384 (O_384,N_9984,N_9839);
nand UO_385 (O_385,N_9812,N_9999);
xnor UO_386 (O_386,N_9964,N_9946);
nand UO_387 (O_387,N_9894,N_9973);
nand UO_388 (O_388,N_9828,N_9880);
or UO_389 (O_389,N_9858,N_9929);
or UO_390 (O_390,N_9996,N_9989);
and UO_391 (O_391,N_9908,N_9937);
or UO_392 (O_392,N_9974,N_9847);
nor UO_393 (O_393,N_9925,N_9823);
nor UO_394 (O_394,N_9981,N_9827);
nand UO_395 (O_395,N_9930,N_9934);
and UO_396 (O_396,N_9959,N_9897);
or UO_397 (O_397,N_9842,N_9860);
nor UO_398 (O_398,N_9879,N_9867);
or UO_399 (O_399,N_9810,N_9828);
nand UO_400 (O_400,N_9949,N_9960);
nand UO_401 (O_401,N_9987,N_9958);
xor UO_402 (O_402,N_9961,N_9922);
nand UO_403 (O_403,N_9844,N_9802);
nand UO_404 (O_404,N_9982,N_9859);
nand UO_405 (O_405,N_9964,N_9865);
nor UO_406 (O_406,N_9922,N_9927);
nor UO_407 (O_407,N_9952,N_9865);
and UO_408 (O_408,N_9971,N_9958);
and UO_409 (O_409,N_9904,N_9858);
or UO_410 (O_410,N_9951,N_9971);
nand UO_411 (O_411,N_9875,N_9915);
nand UO_412 (O_412,N_9872,N_9921);
nor UO_413 (O_413,N_9854,N_9956);
and UO_414 (O_414,N_9859,N_9800);
nand UO_415 (O_415,N_9956,N_9943);
and UO_416 (O_416,N_9984,N_9866);
xor UO_417 (O_417,N_9933,N_9806);
xnor UO_418 (O_418,N_9881,N_9974);
nor UO_419 (O_419,N_9959,N_9919);
nand UO_420 (O_420,N_9892,N_9959);
nor UO_421 (O_421,N_9943,N_9833);
nor UO_422 (O_422,N_9948,N_9958);
xor UO_423 (O_423,N_9942,N_9943);
xnor UO_424 (O_424,N_9852,N_9898);
nor UO_425 (O_425,N_9960,N_9908);
nand UO_426 (O_426,N_9914,N_9850);
and UO_427 (O_427,N_9971,N_9892);
nor UO_428 (O_428,N_9808,N_9872);
and UO_429 (O_429,N_9947,N_9854);
nand UO_430 (O_430,N_9937,N_9912);
nand UO_431 (O_431,N_9967,N_9835);
or UO_432 (O_432,N_9810,N_9998);
nor UO_433 (O_433,N_9947,N_9884);
and UO_434 (O_434,N_9835,N_9847);
or UO_435 (O_435,N_9957,N_9960);
or UO_436 (O_436,N_9971,N_9969);
and UO_437 (O_437,N_9912,N_9834);
nor UO_438 (O_438,N_9983,N_9831);
and UO_439 (O_439,N_9916,N_9970);
and UO_440 (O_440,N_9960,N_9966);
xnor UO_441 (O_441,N_9850,N_9947);
and UO_442 (O_442,N_9862,N_9947);
and UO_443 (O_443,N_9901,N_9948);
nand UO_444 (O_444,N_9851,N_9814);
nand UO_445 (O_445,N_9864,N_9846);
nor UO_446 (O_446,N_9960,N_9894);
nor UO_447 (O_447,N_9832,N_9844);
xnor UO_448 (O_448,N_9837,N_9834);
nand UO_449 (O_449,N_9886,N_9906);
and UO_450 (O_450,N_9934,N_9843);
or UO_451 (O_451,N_9896,N_9868);
nor UO_452 (O_452,N_9907,N_9974);
and UO_453 (O_453,N_9926,N_9869);
and UO_454 (O_454,N_9937,N_9887);
nor UO_455 (O_455,N_9869,N_9979);
nand UO_456 (O_456,N_9939,N_9962);
and UO_457 (O_457,N_9829,N_9847);
or UO_458 (O_458,N_9915,N_9963);
nor UO_459 (O_459,N_9966,N_9914);
nand UO_460 (O_460,N_9948,N_9913);
and UO_461 (O_461,N_9914,N_9822);
nor UO_462 (O_462,N_9980,N_9801);
nor UO_463 (O_463,N_9857,N_9892);
or UO_464 (O_464,N_9819,N_9996);
nor UO_465 (O_465,N_9801,N_9805);
nor UO_466 (O_466,N_9888,N_9863);
nand UO_467 (O_467,N_9900,N_9860);
or UO_468 (O_468,N_9806,N_9916);
or UO_469 (O_469,N_9822,N_9848);
nor UO_470 (O_470,N_9993,N_9904);
or UO_471 (O_471,N_9933,N_9992);
nand UO_472 (O_472,N_9837,N_9920);
or UO_473 (O_473,N_9813,N_9973);
nand UO_474 (O_474,N_9908,N_9813);
nand UO_475 (O_475,N_9828,N_9850);
nor UO_476 (O_476,N_9932,N_9845);
or UO_477 (O_477,N_9905,N_9915);
nand UO_478 (O_478,N_9857,N_9975);
or UO_479 (O_479,N_9942,N_9900);
and UO_480 (O_480,N_9826,N_9925);
nand UO_481 (O_481,N_9841,N_9974);
nand UO_482 (O_482,N_9975,N_9904);
or UO_483 (O_483,N_9943,N_9958);
and UO_484 (O_484,N_9982,N_9960);
nor UO_485 (O_485,N_9921,N_9948);
xnor UO_486 (O_486,N_9829,N_9995);
and UO_487 (O_487,N_9993,N_9865);
or UO_488 (O_488,N_9954,N_9859);
xnor UO_489 (O_489,N_9961,N_9931);
nor UO_490 (O_490,N_9809,N_9890);
nor UO_491 (O_491,N_9995,N_9988);
and UO_492 (O_492,N_9911,N_9988);
nand UO_493 (O_493,N_9879,N_9892);
or UO_494 (O_494,N_9923,N_9944);
and UO_495 (O_495,N_9969,N_9902);
nor UO_496 (O_496,N_9855,N_9912);
or UO_497 (O_497,N_9893,N_9819);
or UO_498 (O_498,N_9825,N_9880);
nand UO_499 (O_499,N_9882,N_9889);
nor UO_500 (O_500,N_9908,N_9975);
xor UO_501 (O_501,N_9941,N_9870);
nor UO_502 (O_502,N_9847,N_9909);
nand UO_503 (O_503,N_9932,N_9884);
nand UO_504 (O_504,N_9896,N_9836);
or UO_505 (O_505,N_9982,N_9973);
or UO_506 (O_506,N_9919,N_9892);
nor UO_507 (O_507,N_9988,N_9813);
nor UO_508 (O_508,N_9894,N_9910);
nand UO_509 (O_509,N_9951,N_9986);
nand UO_510 (O_510,N_9804,N_9922);
nor UO_511 (O_511,N_9820,N_9827);
or UO_512 (O_512,N_9968,N_9839);
or UO_513 (O_513,N_9828,N_9968);
and UO_514 (O_514,N_9876,N_9971);
or UO_515 (O_515,N_9927,N_9855);
xor UO_516 (O_516,N_9850,N_9888);
and UO_517 (O_517,N_9898,N_9989);
or UO_518 (O_518,N_9819,N_9983);
or UO_519 (O_519,N_9891,N_9893);
and UO_520 (O_520,N_9995,N_9820);
nand UO_521 (O_521,N_9973,N_9827);
nand UO_522 (O_522,N_9973,N_9869);
nand UO_523 (O_523,N_9884,N_9873);
and UO_524 (O_524,N_9948,N_9932);
nand UO_525 (O_525,N_9859,N_9918);
and UO_526 (O_526,N_9902,N_9997);
and UO_527 (O_527,N_9950,N_9987);
nand UO_528 (O_528,N_9978,N_9945);
and UO_529 (O_529,N_9893,N_9956);
or UO_530 (O_530,N_9955,N_9927);
and UO_531 (O_531,N_9926,N_9990);
nand UO_532 (O_532,N_9916,N_9909);
nor UO_533 (O_533,N_9908,N_9837);
and UO_534 (O_534,N_9872,N_9878);
nor UO_535 (O_535,N_9843,N_9995);
nand UO_536 (O_536,N_9864,N_9805);
xnor UO_537 (O_537,N_9928,N_9910);
and UO_538 (O_538,N_9847,N_9869);
nor UO_539 (O_539,N_9944,N_9854);
nor UO_540 (O_540,N_9913,N_9932);
nand UO_541 (O_541,N_9941,N_9964);
nand UO_542 (O_542,N_9959,N_9874);
nand UO_543 (O_543,N_9831,N_9875);
and UO_544 (O_544,N_9812,N_9804);
and UO_545 (O_545,N_9927,N_9893);
nor UO_546 (O_546,N_9806,N_9977);
or UO_547 (O_547,N_9826,N_9993);
nand UO_548 (O_548,N_9922,N_9875);
nand UO_549 (O_549,N_9864,N_9895);
and UO_550 (O_550,N_9849,N_9940);
and UO_551 (O_551,N_9990,N_9895);
and UO_552 (O_552,N_9852,N_9936);
and UO_553 (O_553,N_9926,N_9886);
nor UO_554 (O_554,N_9973,N_9853);
nor UO_555 (O_555,N_9946,N_9844);
nor UO_556 (O_556,N_9920,N_9835);
xnor UO_557 (O_557,N_9847,N_9984);
and UO_558 (O_558,N_9985,N_9875);
nor UO_559 (O_559,N_9926,N_9887);
and UO_560 (O_560,N_9899,N_9977);
and UO_561 (O_561,N_9860,N_9910);
nor UO_562 (O_562,N_9956,N_9845);
or UO_563 (O_563,N_9939,N_9886);
nor UO_564 (O_564,N_9955,N_9984);
nor UO_565 (O_565,N_9985,N_9837);
nor UO_566 (O_566,N_9869,N_9944);
xnor UO_567 (O_567,N_9953,N_9894);
nor UO_568 (O_568,N_9939,N_9869);
xnor UO_569 (O_569,N_9959,N_9883);
and UO_570 (O_570,N_9917,N_9825);
or UO_571 (O_571,N_9907,N_9887);
nand UO_572 (O_572,N_9891,N_9804);
nand UO_573 (O_573,N_9976,N_9820);
and UO_574 (O_574,N_9829,N_9996);
nand UO_575 (O_575,N_9919,N_9831);
and UO_576 (O_576,N_9837,N_9803);
nor UO_577 (O_577,N_9825,N_9896);
nand UO_578 (O_578,N_9896,N_9977);
nor UO_579 (O_579,N_9919,N_9992);
nor UO_580 (O_580,N_9999,N_9959);
nand UO_581 (O_581,N_9804,N_9913);
or UO_582 (O_582,N_9973,N_9854);
nand UO_583 (O_583,N_9809,N_9955);
and UO_584 (O_584,N_9980,N_9985);
nor UO_585 (O_585,N_9915,N_9818);
or UO_586 (O_586,N_9988,N_9972);
and UO_587 (O_587,N_9997,N_9945);
nor UO_588 (O_588,N_9939,N_9828);
and UO_589 (O_589,N_9884,N_9910);
nor UO_590 (O_590,N_9828,N_9924);
or UO_591 (O_591,N_9822,N_9983);
and UO_592 (O_592,N_9930,N_9984);
and UO_593 (O_593,N_9932,N_9908);
or UO_594 (O_594,N_9960,N_9906);
or UO_595 (O_595,N_9943,N_9941);
nor UO_596 (O_596,N_9987,N_9875);
nand UO_597 (O_597,N_9902,N_9929);
xnor UO_598 (O_598,N_9805,N_9834);
xnor UO_599 (O_599,N_9884,N_9992);
or UO_600 (O_600,N_9994,N_9806);
nand UO_601 (O_601,N_9924,N_9818);
or UO_602 (O_602,N_9835,N_9856);
and UO_603 (O_603,N_9963,N_9828);
xnor UO_604 (O_604,N_9925,N_9920);
and UO_605 (O_605,N_9888,N_9885);
and UO_606 (O_606,N_9835,N_9813);
and UO_607 (O_607,N_9969,N_9895);
and UO_608 (O_608,N_9826,N_9994);
nand UO_609 (O_609,N_9856,N_9821);
xnor UO_610 (O_610,N_9844,N_9956);
or UO_611 (O_611,N_9879,N_9941);
or UO_612 (O_612,N_9821,N_9916);
nand UO_613 (O_613,N_9900,N_9894);
and UO_614 (O_614,N_9989,N_9912);
nor UO_615 (O_615,N_9914,N_9910);
nand UO_616 (O_616,N_9886,N_9827);
nor UO_617 (O_617,N_9831,N_9884);
nor UO_618 (O_618,N_9959,N_9855);
nor UO_619 (O_619,N_9864,N_9984);
xor UO_620 (O_620,N_9966,N_9807);
nor UO_621 (O_621,N_9887,N_9857);
nand UO_622 (O_622,N_9840,N_9884);
nand UO_623 (O_623,N_9896,N_9870);
nor UO_624 (O_624,N_9986,N_9845);
and UO_625 (O_625,N_9995,N_9966);
and UO_626 (O_626,N_9989,N_9927);
or UO_627 (O_627,N_9931,N_9963);
and UO_628 (O_628,N_9804,N_9889);
nand UO_629 (O_629,N_9816,N_9934);
nor UO_630 (O_630,N_9966,N_9868);
nor UO_631 (O_631,N_9877,N_9913);
xor UO_632 (O_632,N_9806,N_9974);
and UO_633 (O_633,N_9960,N_9940);
nand UO_634 (O_634,N_9902,N_9810);
nor UO_635 (O_635,N_9891,N_9884);
nand UO_636 (O_636,N_9939,N_9960);
xnor UO_637 (O_637,N_9941,N_9821);
xor UO_638 (O_638,N_9921,N_9874);
xor UO_639 (O_639,N_9880,N_9848);
nor UO_640 (O_640,N_9820,N_9966);
nor UO_641 (O_641,N_9908,N_9841);
nand UO_642 (O_642,N_9843,N_9884);
or UO_643 (O_643,N_9923,N_9970);
nor UO_644 (O_644,N_9831,N_9805);
nor UO_645 (O_645,N_9881,N_9866);
nand UO_646 (O_646,N_9911,N_9843);
nand UO_647 (O_647,N_9944,N_9982);
and UO_648 (O_648,N_9863,N_9985);
nand UO_649 (O_649,N_9904,N_9961);
or UO_650 (O_650,N_9865,N_9855);
nor UO_651 (O_651,N_9941,N_9936);
nand UO_652 (O_652,N_9803,N_9844);
nand UO_653 (O_653,N_9957,N_9894);
nand UO_654 (O_654,N_9807,N_9844);
and UO_655 (O_655,N_9852,N_9888);
or UO_656 (O_656,N_9848,N_9974);
nor UO_657 (O_657,N_9936,N_9899);
and UO_658 (O_658,N_9853,N_9876);
xnor UO_659 (O_659,N_9913,N_9965);
and UO_660 (O_660,N_9933,N_9871);
or UO_661 (O_661,N_9930,N_9980);
and UO_662 (O_662,N_9941,N_9901);
nor UO_663 (O_663,N_9967,N_9820);
nor UO_664 (O_664,N_9809,N_9978);
nor UO_665 (O_665,N_9919,N_9921);
nor UO_666 (O_666,N_9814,N_9951);
nand UO_667 (O_667,N_9957,N_9989);
and UO_668 (O_668,N_9868,N_9844);
nor UO_669 (O_669,N_9906,N_9808);
and UO_670 (O_670,N_9887,N_9849);
or UO_671 (O_671,N_9938,N_9899);
or UO_672 (O_672,N_9830,N_9820);
xnor UO_673 (O_673,N_9994,N_9907);
nor UO_674 (O_674,N_9903,N_9854);
or UO_675 (O_675,N_9867,N_9939);
and UO_676 (O_676,N_9858,N_9970);
and UO_677 (O_677,N_9878,N_9886);
or UO_678 (O_678,N_9811,N_9968);
nand UO_679 (O_679,N_9976,N_9808);
nor UO_680 (O_680,N_9968,N_9862);
or UO_681 (O_681,N_9890,N_9902);
and UO_682 (O_682,N_9804,N_9982);
nor UO_683 (O_683,N_9993,N_9978);
nor UO_684 (O_684,N_9967,N_9828);
nand UO_685 (O_685,N_9911,N_9867);
nor UO_686 (O_686,N_9809,N_9939);
and UO_687 (O_687,N_9844,N_9920);
or UO_688 (O_688,N_9849,N_9931);
nor UO_689 (O_689,N_9868,N_9920);
nand UO_690 (O_690,N_9852,N_9879);
or UO_691 (O_691,N_9877,N_9809);
xor UO_692 (O_692,N_9947,N_9846);
nand UO_693 (O_693,N_9822,N_9872);
or UO_694 (O_694,N_9876,N_9813);
or UO_695 (O_695,N_9954,N_9809);
or UO_696 (O_696,N_9820,N_9854);
nand UO_697 (O_697,N_9817,N_9881);
and UO_698 (O_698,N_9804,N_9960);
and UO_699 (O_699,N_9959,N_9957);
nor UO_700 (O_700,N_9994,N_9851);
nand UO_701 (O_701,N_9843,N_9976);
and UO_702 (O_702,N_9917,N_9938);
nor UO_703 (O_703,N_9926,N_9885);
nor UO_704 (O_704,N_9916,N_9975);
nor UO_705 (O_705,N_9828,N_9937);
nor UO_706 (O_706,N_9879,N_9968);
nand UO_707 (O_707,N_9989,N_9931);
nand UO_708 (O_708,N_9866,N_9958);
or UO_709 (O_709,N_9971,N_9938);
and UO_710 (O_710,N_9926,N_9801);
nor UO_711 (O_711,N_9923,N_9883);
nor UO_712 (O_712,N_9896,N_9819);
and UO_713 (O_713,N_9867,N_9980);
nand UO_714 (O_714,N_9975,N_9837);
xor UO_715 (O_715,N_9935,N_9818);
xnor UO_716 (O_716,N_9846,N_9863);
xnor UO_717 (O_717,N_9868,N_9840);
nand UO_718 (O_718,N_9806,N_9842);
or UO_719 (O_719,N_9903,N_9921);
and UO_720 (O_720,N_9897,N_9972);
nor UO_721 (O_721,N_9821,N_9840);
nor UO_722 (O_722,N_9900,N_9917);
or UO_723 (O_723,N_9929,N_9817);
nor UO_724 (O_724,N_9961,N_9801);
xnor UO_725 (O_725,N_9991,N_9879);
and UO_726 (O_726,N_9825,N_9959);
nor UO_727 (O_727,N_9900,N_9914);
or UO_728 (O_728,N_9933,N_9855);
and UO_729 (O_729,N_9866,N_9927);
and UO_730 (O_730,N_9860,N_9801);
nand UO_731 (O_731,N_9805,N_9946);
and UO_732 (O_732,N_9978,N_9989);
and UO_733 (O_733,N_9904,N_9890);
nor UO_734 (O_734,N_9826,N_9963);
and UO_735 (O_735,N_9995,N_9981);
nor UO_736 (O_736,N_9810,N_9962);
and UO_737 (O_737,N_9939,N_9879);
nor UO_738 (O_738,N_9927,N_9996);
nand UO_739 (O_739,N_9883,N_9830);
nor UO_740 (O_740,N_9847,N_9866);
and UO_741 (O_741,N_9991,N_9924);
and UO_742 (O_742,N_9993,N_9954);
nand UO_743 (O_743,N_9847,N_9953);
nor UO_744 (O_744,N_9902,N_9925);
or UO_745 (O_745,N_9852,N_9829);
nand UO_746 (O_746,N_9839,N_9996);
nand UO_747 (O_747,N_9828,N_9888);
or UO_748 (O_748,N_9931,N_9862);
or UO_749 (O_749,N_9996,N_9947);
nor UO_750 (O_750,N_9976,N_9826);
nor UO_751 (O_751,N_9827,N_9863);
and UO_752 (O_752,N_9934,N_9901);
nand UO_753 (O_753,N_9876,N_9865);
nor UO_754 (O_754,N_9995,N_9969);
nand UO_755 (O_755,N_9851,N_9988);
nor UO_756 (O_756,N_9855,N_9828);
and UO_757 (O_757,N_9904,N_9982);
or UO_758 (O_758,N_9990,N_9835);
nand UO_759 (O_759,N_9981,N_9876);
and UO_760 (O_760,N_9815,N_9975);
nand UO_761 (O_761,N_9807,N_9884);
and UO_762 (O_762,N_9815,N_9956);
nand UO_763 (O_763,N_9845,N_9898);
and UO_764 (O_764,N_9870,N_9875);
or UO_765 (O_765,N_9901,N_9964);
nand UO_766 (O_766,N_9835,N_9824);
xor UO_767 (O_767,N_9848,N_9888);
nor UO_768 (O_768,N_9869,N_9855);
or UO_769 (O_769,N_9846,N_9995);
nand UO_770 (O_770,N_9873,N_9872);
nor UO_771 (O_771,N_9861,N_9895);
or UO_772 (O_772,N_9887,N_9809);
nor UO_773 (O_773,N_9861,N_9851);
nand UO_774 (O_774,N_9921,N_9811);
xnor UO_775 (O_775,N_9932,N_9820);
and UO_776 (O_776,N_9953,N_9929);
nor UO_777 (O_777,N_9861,N_9803);
or UO_778 (O_778,N_9925,N_9845);
nor UO_779 (O_779,N_9854,N_9885);
nand UO_780 (O_780,N_9851,N_9911);
xor UO_781 (O_781,N_9934,N_9817);
and UO_782 (O_782,N_9962,N_9915);
nand UO_783 (O_783,N_9825,N_9864);
nand UO_784 (O_784,N_9858,N_9850);
nand UO_785 (O_785,N_9938,N_9901);
and UO_786 (O_786,N_9825,N_9945);
nand UO_787 (O_787,N_9982,N_9955);
nor UO_788 (O_788,N_9872,N_9820);
nor UO_789 (O_789,N_9931,N_9816);
nor UO_790 (O_790,N_9853,N_9970);
nor UO_791 (O_791,N_9910,N_9806);
or UO_792 (O_792,N_9890,N_9839);
or UO_793 (O_793,N_9981,N_9857);
and UO_794 (O_794,N_9922,N_9848);
nand UO_795 (O_795,N_9926,N_9849);
and UO_796 (O_796,N_9933,N_9905);
or UO_797 (O_797,N_9967,N_9936);
and UO_798 (O_798,N_9921,N_9887);
xor UO_799 (O_799,N_9974,N_9918);
or UO_800 (O_800,N_9948,N_9803);
nor UO_801 (O_801,N_9864,N_9862);
or UO_802 (O_802,N_9949,N_9976);
or UO_803 (O_803,N_9824,N_9897);
nor UO_804 (O_804,N_9870,N_9986);
or UO_805 (O_805,N_9858,N_9875);
nand UO_806 (O_806,N_9848,N_9898);
or UO_807 (O_807,N_9820,N_9871);
nor UO_808 (O_808,N_9885,N_9991);
nand UO_809 (O_809,N_9880,N_9850);
or UO_810 (O_810,N_9930,N_9999);
xnor UO_811 (O_811,N_9912,N_9905);
nand UO_812 (O_812,N_9978,N_9912);
nor UO_813 (O_813,N_9964,N_9839);
and UO_814 (O_814,N_9850,N_9851);
nand UO_815 (O_815,N_9935,N_9969);
or UO_816 (O_816,N_9862,N_9973);
nand UO_817 (O_817,N_9862,N_9824);
or UO_818 (O_818,N_9815,N_9940);
nand UO_819 (O_819,N_9872,N_9875);
and UO_820 (O_820,N_9880,N_9973);
nand UO_821 (O_821,N_9883,N_9915);
nor UO_822 (O_822,N_9927,N_9939);
nand UO_823 (O_823,N_9986,N_9846);
nor UO_824 (O_824,N_9973,N_9963);
and UO_825 (O_825,N_9858,N_9899);
nor UO_826 (O_826,N_9951,N_9872);
and UO_827 (O_827,N_9937,N_9916);
and UO_828 (O_828,N_9958,N_9995);
nand UO_829 (O_829,N_9930,N_9983);
or UO_830 (O_830,N_9942,N_9990);
or UO_831 (O_831,N_9988,N_9859);
or UO_832 (O_832,N_9968,N_9815);
xnor UO_833 (O_833,N_9985,N_9811);
nand UO_834 (O_834,N_9937,N_9956);
nor UO_835 (O_835,N_9954,N_9804);
nor UO_836 (O_836,N_9880,N_9944);
or UO_837 (O_837,N_9800,N_9957);
or UO_838 (O_838,N_9830,N_9843);
nor UO_839 (O_839,N_9950,N_9911);
and UO_840 (O_840,N_9949,N_9857);
nand UO_841 (O_841,N_9915,N_9910);
or UO_842 (O_842,N_9886,N_9883);
nor UO_843 (O_843,N_9918,N_9924);
or UO_844 (O_844,N_9896,N_9860);
or UO_845 (O_845,N_9971,N_9891);
xnor UO_846 (O_846,N_9945,N_9989);
or UO_847 (O_847,N_9876,N_9828);
xor UO_848 (O_848,N_9979,N_9872);
or UO_849 (O_849,N_9939,N_9988);
nand UO_850 (O_850,N_9974,N_9969);
and UO_851 (O_851,N_9992,N_9834);
and UO_852 (O_852,N_9979,N_9966);
and UO_853 (O_853,N_9881,N_9963);
and UO_854 (O_854,N_9832,N_9930);
nand UO_855 (O_855,N_9912,N_9961);
nor UO_856 (O_856,N_9888,N_9971);
nand UO_857 (O_857,N_9991,N_9880);
and UO_858 (O_858,N_9914,N_9942);
nand UO_859 (O_859,N_9912,N_9889);
and UO_860 (O_860,N_9881,N_9900);
nor UO_861 (O_861,N_9913,N_9871);
xnor UO_862 (O_862,N_9905,N_9885);
nand UO_863 (O_863,N_9836,N_9817);
nand UO_864 (O_864,N_9930,N_9997);
and UO_865 (O_865,N_9896,N_9861);
nor UO_866 (O_866,N_9874,N_9929);
and UO_867 (O_867,N_9823,N_9943);
nand UO_868 (O_868,N_9916,N_9984);
nor UO_869 (O_869,N_9868,N_9909);
or UO_870 (O_870,N_9866,N_9929);
nand UO_871 (O_871,N_9918,N_9905);
nand UO_872 (O_872,N_9800,N_9815);
nor UO_873 (O_873,N_9851,N_9986);
nand UO_874 (O_874,N_9971,N_9832);
or UO_875 (O_875,N_9904,N_9883);
nand UO_876 (O_876,N_9906,N_9897);
nand UO_877 (O_877,N_9830,N_9859);
and UO_878 (O_878,N_9982,N_9907);
or UO_879 (O_879,N_9888,N_9886);
nor UO_880 (O_880,N_9865,N_9867);
xnor UO_881 (O_881,N_9935,N_9806);
nor UO_882 (O_882,N_9951,N_9949);
and UO_883 (O_883,N_9840,N_9953);
nand UO_884 (O_884,N_9827,N_9803);
xor UO_885 (O_885,N_9856,N_9878);
nand UO_886 (O_886,N_9998,N_9928);
and UO_887 (O_887,N_9828,N_9944);
or UO_888 (O_888,N_9909,N_9895);
nor UO_889 (O_889,N_9802,N_9986);
nand UO_890 (O_890,N_9814,N_9921);
xor UO_891 (O_891,N_9842,N_9973);
nand UO_892 (O_892,N_9882,N_9856);
nand UO_893 (O_893,N_9895,N_9946);
and UO_894 (O_894,N_9941,N_9955);
nand UO_895 (O_895,N_9890,N_9870);
nor UO_896 (O_896,N_9996,N_9935);
and UO_897 (O_897,N_9942,N_9939);
xor UO_898 (O_898,N_9836,N_9929);
nor UO_899 (O_899,N_9940,N_9919);
or UO_900 (O_900,N_9871,N_9929);
nand UO_901 (O_901,N_9999,N_9802);
nand UO_902 (O_902,N_9871,N_9926);
nand UO_903 (O_903,N_9868,N_9941);
nor UO_904 (O_904,N_9807,N_9868);
and UO_905 (O_905,N_9919,N_9835);
and UO_906 (O_906,N_9991,N_9844);
or UO_907 (O_907,N_9994,N_9968);
or UO_908 (O_908,N_9983,N_9988);
nand UO_909 (O_909,N_9828,N_9953);
nand UO_910 (O_910,N_9957,N_9831);
and UO_911 (O_911,N_9856,N_9845);
and UO_912 (O_912,N_9811,N_9808);
nor UO_913 (O_913,N_9901,N_9918);
and UO_914 (O_914,N_9914,N_9899);
nand UO_915 (O_915,N_9842,N_9964);
nand UO_916 (O_916,N_9933,N_9877);
nand UO_917 (O_917,N_9906,N_9859);
or UO_918 (O_918,N_9947,N_9981);
nor UO_919 (O_919,N_9925,N_9940);
or UO_920 (O_920,N_9930,N_9837);
nand UO_921 (O_921,N_9876,N_9921);
xnor UO_922 (O_922,N_9962,N_9818);
or UO_923 (O_923,N_9898,N_9812);
nor UO_924 (O_924,N_9852,N_9895);
and UO_925 (O_925,N_9871,N_9932);
xnor UO_926 (O_926,N_9921,N_9867);
nor UO_927 (O_927,N_9866,N_9985);
or UO_928 (O_928,N_9876,N_9824);
nand UO_929 (O_929,N_9830,N_9970);
xnor UO_930 (O_930,N_9836,N_9800);
nor UO_931 (O_931,N_9809,N_9970);
xnor UO_932 (O_932,N_9903,N_9955);
and UO_933 (O_933,N_9900,N_9965);
nor UO_934 (O_934,N_9884,N_9930);
nand UO_935 (O_935,N_9856,N_9853);
xor UO_936 (O_936,N_9903,N_9977);
nor UO_937 (O_937,N_9986,N_9873);
or UO_938 (O_938,N_9991,N_9860);
or UO_939 (O_939,N_9989,N_9929);
nor UO_940 (O_940,N_9948,N_9873);
nor UO_941 (O_941,N_9902,N_9834);
nor UO_942 (O_942,N_9810,N_9838);
or UO_943 (O_943,N_9964,N_9998);
or UO_944 (O_944,N_9928,N_9849);
nand UO_945 (O_945,N_9994,N_9871);
nand UO_946 (O_946,N_9907,N_9828);
and UO_947 (O_947,N_9873,N_9892);
or UO_948 (O_948,N_9808,N_9981);
nand UO_949 (O_949,N_9912,N_9898);
xor UO_950 (O_950,N_9842,N_9814);
nor UO_951 (O_951,N_9902,N_9820);
or UO_952 (O_952,N_9929,N_9854);
and UO_953 (O_953,N_9936,N_9905);
xnor UO_954 (O_954,N_9801,N_9859);
xnor UO_955 (O_955,N_9937,N_9929);
nand UO_956 (O_956,N_9871,N_9971);
nand UO_957 (O_957,N_9923,N_9976);
xnor UO_958 (O_958,N_9959,N_9818);
nor UO_959 (O_959,N_9837,N_9974);
and UO_960 (O_960,N_9814,N_9986);
or UO_961 (O_961,N_9893,N_9983);
and UO_962 (O_962,N_9892,N_9836);
or UO_963 (O_963,N_9940,N_9971);
and UO_964 (O_964,N_9823,N_9948);
or UO_965 (O_965,N_9839,N_9938);
xor UO_966 (O_966,N_9965,N_9832);
and UO_967 (O_967,N_9801,N_9851);
nor UO_968 (O_968,N_9821,N_9841);
or UO_969 (O_969,N_9992,N_9886);
and UO_970 (O_970,N_9949,N_9824);
nand UO_971 (O_971,N_9803,N_9921);
nand UO_972 (O_972,N_9852,N_9809);
and UO_973 (O_973,N_9981,N_9819);
nand UO_974 (O_974,N_9933,N_9879);
and UO_975 (O_975,N_9821,N_9854);
or UO_976 (O_976,N_9877,N_9820);
and UO_977 (O_977,N_9901,N_9884);
or UO_978 (O_978,N_9965,N_9939);
xor UO_979 (O_979,N_9979,N_9893);
or UO_980 (O_980,N_9963,N_9895);
nand UO_981 (O_981,N_9825,N_9960);
xor UO_982 (O_982,N_9805,N_9912);
and UO_983 (O_983,N_9828,N_9974);
and UO_984 (O_984,N_9988,N_9948);
and UO_985 (O_985,N_9992,N_9843);
nand UO_986 (O_986,N_9980,N_9946);
xor UO_987 (O_987,N_9994,N_9942);
or UO_988 (O_988,N_9863,N_9866);
and UO_989 (O_989,N_9992,N_9880);
and UO_990 (O_990,N_9872,N_9864);
or UO_991 (O_991,N_9977,N_9894);
or UO_992 (O_992,N_9886,N_9892);
and UO_993 (O_993,N_9839,N_9828);
and UO_994 (O_994,N_9884,N_9955);
nor UO_995 (O_995,N_9959,N_9882);
nor UO_996 (O_996,N_9835,N_9949);
nand UO_997 (O_997,N_9904,N_9885);
or UO_998 (O_998,N_9887,N_9855);
xnor UO_999 (O_999,N_9882,N_9988);
xor UO_1000 (O_1000,N_9953,N_9981);
and UO_1001 (O_1001,N_9955,N_9976);
nor UO_1002 (O_1002,N_9933,N_9880);
and UO_1003 (O_1003,N_9882,N_9995);
or UO_1004 (O_1004,N_9838,N_9918);
nor UO_1005 (O_1005,N_9974,N_9867);
or UO_1006 (O_1006,N_9841,N_9913);
nand UO_1007 (O_1007,N_9894,N_9972);
and UO_1008 (O_1008,N_9936,N_9842);
nor UO_1009 (O_1009,N_9887,N_9903);
nor UO_1010 (O_1010,N_9825,N_9833);
or UO_1011 (O_1011,N_9886,N_9981);
or UO_1012 (O_1012,N_9973,N_9920);
nand UO_1013 (O_1013,N_9911,N_9920);
nand UO_1014 (O_1014,N_9923,N_9876);
xnor UO_1015 (O_1015,N_9891,N_9820);
nand UO_1016 (O_1016,N_9811,N_9905);
xor UO_1017 (O_1017,N_9855,N_9932);
or UO_1018 (O_1018,N_9957,N_9856);
and UO_1019 (O_1019,N_9871,N_9817);
and UO_1020 (O_1020,N_9806,N_9871);
nand UO_1021 (O_1021,N_9870,N_9853);
and UO_1022 (O_1022,N_9973,N_9987);
or UO_1023 (O_1023,N_9836,N_9822);
and UO_1024 (O_1024,N_9963,N_9975);
and UO_1025 (O_1025,N_9995,N_9834);
or UO_1026 (O_1026,N_9950,N_9830);
nand UO_1027 (O_1027,N_9963,N_9857);
nor UO_1028 (O_1028,N_9967,N_9868);
and UO_1029 (O_1029,N_9948,N_9841);
xnor UO_1030 (O_1030,N_9969,N_9872);
or UO_1031 (O_1031,N_9952,N_9955);
nor UO_1032 (O_1032,N_9880,N_9818);
nor UO_1033 (O_1033,N_9874,N_9839);
xnor UO_1034 (O_1034,N_9847,N_9806);
nand UO_1035 (O_1035,N_9873,N_9825);
xnor UO_1036 (O_1036,N_9805,N_9839);
or UO_1037 (O_1037,N_9940,N_9901);
nand UO_1038 (O_1038,N_9892,N_9883);
and UO_1039 (O_1039,N_9998,N_9973);
nand UO_1040 (O_1040,N_9898,N_9891);
and UO_1041 (O_1041,N_9832,N_9840);
and UO_1042 (O_1042,N_9951,N_9864);
or UO_1043 (O_1043,N_9988,N_9879);
and UO_1044 (O_1044,N_9891,N_9934);
and UO_1045 (O_1045,N_9800,N_9833);
nand UO_1046 (O_1046,N_9936,N_9868);
or UO_1047 (O_1047,N_9885,N_9996);
or UO_1048 (O_1048,N_9934,N_9910);
and UO_1049 (O_1049,N_9921,N_9861);
nand UO_1050 (O_1050,N_9989,N_9925);
and UO_1051 (O_1051,N_9922,N_9836);
nor UO_1052 (O_1052,N_9940,N_9934);
or UO_1053 (O_1053,N_9858,N_9882);
and UO_1054 (O_1054,N_9800,N_9890);
or UO_1055 (O_1055,N_9867,N_9889);
or UO_1056 (O_1056,N_9985,N_9872);
and UO_1057 (O_1057,N_9849,N_9924);
and UO_1058 (O_1058,N_9854,N_9968);
and UO_1059 (O_1059,N_9873,N_9804);
and UO_1060 (O_1060,N_9998,N_9874);
nand UO_1061 (O_1061,N_9909,N_9819);
nor UO_1062 (O_1062,N_9884,N_9996);
nand UO_1063 (O_1063,N_9862,N_9849);
and UO_1064 (O_1064,N_9804,N_9978);
nand UO_1065 (O_1065,N_9833,N_9945);
or UO_1066 (O_1066,N_9905,N_9965);
or UO_1067 (O_1067,N_9987,N_9919);
or UO_1068 (O_1068,N_9937,N_9854);
nand UO_1069 (O_1069,N_9989,N_9827);
nand UO_1070 (O_1070,N_9879,N_9832);
nand UO_1071 (O_1071,N_9806,N_9821);
and UO_1072 (O_1072,N_9995,N_9931);
and UO_1073 (O_1073,N_9969,N_9833);
nand UO_1074 (O_1074,N_9899,N_9828);
nand UO_1075 (O_1075,N_9803,N_9939);
or UO_1076 (O_1076,N_9871,N_9939);
nor UO_1077 (O_1077,N_9924,N_9844);
nand UO_1078 (O_1078,N_9868,N_9938);
or UO_1079 (O_1079,N_9952,N_9962);
or UO_1080 (O_1080,N_9865,N_9894);
nor UO_1081 (O_1081,N_9967,N_9838);
or UO_1082 (O_1082,N_9805,N_9840);
or UO_1083 (O_1083,N_9908,N_9838);
xor UO_1084 (O_1084,N_9942,N_9967);
nand UO_1085 (O_1085,N_9811,N_9941);
and UO_1086 (O_1086,N_9809,N_9844);
or UO_1087 (O_1087,N_9841,N_9848);
nor UO_1088 (O_1088,N_9960,N_9953);
or UO_1089 (O_1089,N_9865,N_9874);
or UO_1090 (O_1090,N_9876,N_9823);
and UO_1091 (O_1091,N_9915,N_9893);
and UO_1092 (O_1092,N_9931,N_9930);
or UO_1093 (O_1093,N_9809,N_9820);
nand UO_1094 (O_1094,N_9900,N_9973);
nand UO_1095 (O_1095,N_9978,N_9907);
or UO_1096 (O_1096,N_9913,N_9862);
and UO_1097 (O_1097,N_9865,N_9911);
or UO_1098 (O_1098,N_9869,N_9810);
nand UO_1099 (O_1099,N_9803,N_9807);
or UO_1100 (O_1100,N_9964,N_9806);
nand UO_1101 (O_1101,N_9872,N_9992);
nand UO_1102 (O_1102,N_9977,N_9881);
or UO_1103 (O_1103,N_9807,N_9901);
nor UO_1104 (O_1104,N_9971,N_9814);
xnor UO_1105 (O_1105,N_9975,N_9999);
or UO_1106 (O_1106,N_9835,N_9969);
nand UO_1107 (O_1107,N_9830,N_9890);
xor UO_1108 (O_1108,N_9811,N_9967);
and UO_1109 (O_1109,N_9996,N_9933);
xnor UO_1110 (O_1110,N_9949,N_9827);
and UO_1111 (O_1111,N_9971,N_9972);
nor UO_1112 (O_1112,N_9975,N_9932);
and UO_1113 (O_1113,N_9994,N_9844);
nor UO_1114 (O_1114,N_9996,N_9997);
and UO_1115 (O_1115,N_9868,N_9937);
or UO_1116 (O_1116,N_9915,N_9953);
and UO_1117 (O_1117,N_9944,N_9827);
xnor UO_1118 (O_1118,N_9897,N_9914);
and UO_1119 (O_1119,N_9892,N_9881);
xnor UO_1120 (O_1120,N_9999,N_9867);
nand UO_1121 (O_1121,N_9933,N_9835);
xnor UO_1122 (O_1122,N_9973,N_9824);
xnor UO_1123 (O_1123,N_9954,N_9843);
nand UO_1124 (O_1124,N_9865,N_9892);
nor UO_1125 (O_1125,N_9936,N_9806);
xnor UO_1126 (O_1126,N_9901,N_9843);
nor UO_1127 (O_1127,N_9984,N_9807);
or UO_1128 (O_1128,N_9923,N_9904);
and UO_1129 (O_1129,N_9997,N_9901);
nor UO_1130 (O_1130,N_9831,N_9947);
nor UO_1131 (O_1131,N_9907,N_9956);
or UO_1132 (O_1132,N_9803,N_9919);
nand UO_1133 (O_1133,N_9934,N_9917);
or UO_1134 (O_1134,N_9889,N_9838);
nand UO_1135 (O_1135,N_9929,N_9951);
or UO_1136 (O_1136,N_9973,N_9944);
nor UO_1137 (O_1137,N_9812,N_9947);
or UO_1138 (O_1138,N_9893,N_9815);
and UO_1139 (O_1139,N_9874,N_9829);
or UO_1140 (O_1140,N_9819,N_9926);
and UO_1141 (O_1141,N_9818,N_9895);
nor UO_1142 (O_1142,N_9978,N_9857);
and UO_1143 (O_1143,N_9808,N_9988);
nand UO_1144 (O_1144,N_9879,N_9986);
nor UO_1145 (O_1145,N_9911,N_9915);
or UO_1146 (O_1146,N_9978,N_9865);
nand UO_1147 (O_1147,N_9994,N_9982);
nor UO_1148 (O_1148,N_9898,N_9923);
or UO_1149 (O_1149,N_9822,N_9840);
xor UO_1150 (O_1150,N_9950,N_9995);
nor UO_1151 (O_1151,N_9946,N_9818);
nor UO_1152 (O_1152,N_9884,N_9975);
nand UO_1153 (O_1153,N_9923,N_9884);
nand UO_1154 (O_1154,N_9927,N_9884);
or UO_1155 (O_1155,N_9961,N_9957);
or UO_1156 (O_1156,N_9973,N_9990);
xor UO_1157 (O_1157,N_9993,N_9989);
or UO_1158 (O_1158,N_9887,N_9822);
and UO_1159 (O_1159,N_9810,N_9929);
nor UO_1160 (O_1160,N_9863,N_9854);
and UO_1161 (O_1161,N_9836,N_9813);
or UO_1162 (O_1162,N_9823,N_9904);
and UO_1163 (O_1163,N_9922,N_9919);
or UO_1164 (O_1164,N_9806,N_9837);
and UO_1165 (O_1165,N_9970,N_9879);
xnor UO_1166 (O_1166,N_9840,N_9878);
or UO_1167 (O_1167,N_9877,N_9988);
nand UO_1168 (O_1168,N_9834,N_9923);
nand UO_1169 (O_1169,N_9846,N_9841);
nand UO_1170 (O_1170,N_9879,N_9875);
nor UO_1171 (O_1171,N_9903,N_9995);
and UO_1172 (O_1172,N_9825,N_9854);
or UO_1173 (O_1173,N_9865,N_9818);
and UO_1174 (O_1174,N_9820,N_9978);
and UO_1175 (O_1175,N_9934,N_9814);
xnor UO_1176 (O_1176,N_9890,N_9895);
nand UO_1177 (O_1177,N_9878,N_9813);
xnor UO_1178 (O_1178,N_9872,N_9869);
xor UO_1179 (O_1179,N_9950,N_9982);
xnor UO_1180 (O_1180,N_9967,N_9964);
nor UO_1181 (O_1181,N_9912,N_9821);
or UO_1182 (O_1182,N_9836,N_9912);
nand UO_1183 (O_1183,N_9944,N_9901);
and UO_1184 (O_1184,N_9980,N_9911);
and UO_1185 (O_1185,N_9966,N_9869);
or UO_1186 (O_1186,N_9956,N_9857);
and UO_1187 (O_1187,N_9876,N_9819);
nand UO_1188 (O_1188,N_9920,N_9904);
nand UO_1189 (O_1189,N_9865,N_9938);
xor UO_1190 (O_1190,N_9883,N_9998);
nor UO_1191 (O_1191,N_9828,N_9866);
xor UO_1192 (O_1192,N_9949,N_9952);
nand UO_1193 (O_1193,N_9834,N_9851);
or UO_1194 (O_1194,N_9999,N_9830);
and UO_1195 (O_1195,N_9877,N_9885);
or UO_1196 (O_1196,N_9825,N_9962);
and UO_1197 (O_1197,N_9877,N_9968);
nand UO_1198 (O_1198,N_9932,N_9942);
and UO_1199 (O_1199,N_9823,N_9985);
nand UO_1200 (O_1200,N_9896,N_9902);
nor UO_1201 (O_1201,N_9806,N_9965);
or UO_1202 (O_1202,N_9824,N_9828);
and UO_1203 (O_1203,N_9969,N_9820);
or UO_1204 (O_1204,N_9983,N_9931);
and UO_1205 (O_1205,N_9974,N_9949);
or UO_1206 (O_1206,N_9901,N_9859);
nor UO_1207 (O_1207,N_9951,N_9853);
nand UO_1208 (O_1208,N_9867,N_9963);
xor UO_1209 (O_1209,N_9948,N_9843);
nor UO_1210 (O_1210,N_9852,N_9942);
or UO_1211 (O_1211,N_9895,N_9874);
nand UO_1212 (O_1212,N_9966,N_9994);
nor UO_1213 (O_1213,N_9925,N_9935);
or UO_1214 (O_1214,N_9991,N_9889);
nand UO_1215 (O_1215,N_9925,N_9851);
xnor UO_1216 (O_1216,N_9895,N_9809);
or UO_1217 (O_1217,N_9991,N_9918);
nor UO_1218 (O_1218,N_9955,N_9938);
and UO_1219 (O_1219,N_9930,N_9918);
and UO_1220 (O_1220,N_9867,N_9940);
nand UO_1221 (O_1221,N_9937,N_9856);
or UO_1222 (O_1222,N_9910,N_9850);
or UO_1223 (O_1223,N_9801,N_9818);
and UO_1224 (O_1224,N_9970,N_9942);
nor UO_1225 (O_1225,N_9824,N_9972);
nor UO_1226 (O_1226,N_9877,N_9974);
nand UO_1227 (O_1227,N_9871,N_9881);
nor UO_1228 (O_1228,N_9892,N_9980);
or UO_1229 (O_1229,N_9850,N_9968);
nand UO_1230 (O_1230,N_9962,N_9967);
or UO_1231 (O_1231,N_9811,N_9910);
nor UO_1232 (O_1232,N_9880,N_9805);
nand UO_1233 (O_1233,N_9971,N_9925);
nand UO_1234 (O_1234,N_9847,N_9821);
or UO_1235 (O_1235,N_9988,N_9856);
and UO_1236 (O_1236,N_9808,N_9876);
and UO_1237 (O_1237,N_9989,N_9987);
and UO_1238 (O_1238,N_9861,N_9883);
and UO_1239 (O_1239,N_9915,N_9988);
or UO_1240 (O_1240,N_9818,N_9987);
nand UO_1241 (O_1241,N_9988,N_9943);
or UO_1242 (O_1242,N_9839,N_9870);
and UO_1243 (O_1243,N_9919,N_9978);
nand UO_1244 (O_1244,N_9828,N_9969);
and UO_1245 (O_1245,N_9998,N_9954);
and UO_1246 (O_1246,N_9946,N_9950);
or UO_1247 (O_1247,N_9825,N_9900);
nor UO_1248 (O_1248,N_9816,N_9832);
xnor UO_1249 (O_1249,N_9897,N_9835);
nand UO_1250 (O_1250,N_9948,N_9995);
nor UO_1251 (O_1251,N_9923,N_9955);
nor UO_1252 (O_1252,N_9959,N_9901);
and UO_1253 (O_1253,N_9965,N_9836);
and UO_1254 (O_1254,N_9810,N_9972);
nand UO_1255 (O_1255,N_9853,N_9839);
and UO_1256 (O_1256,N_9848,N_9803);
or UO_1257 (O_1257,N_9845,N_9911);
nand UO_1258 (O_1258,N_9990,N_9916);
nand UO_1259 (O_1259,N_9846,N_9840);
nor UO_1260 (O_1260,N_9942,N_9820);
nor UO_1261 (O_1261,N_9909,N_9855);
or UO_1262 (O_1262,N_9916,N_9847);
or UO_1263 (O_1263,N_9818,N_9847);
nor UO_1264 (O_1264,N_9956,N_9931);
nor UO_1265 (O_1265,N_9808,N_9860);
nor UO_1266 (O_1266,N_9959,N_9974);
nand UO_1267 (O_1267,N_9886,N_9830);
or UO_1268 (O_1268,N_9957,N_9985);
nand UO_1269 (O_1269,N_9912,N_9976);
nand UO_1270 (O_1270,N_9967,N_9825);
nand UO_1271 (O_1271,N_9815,N_9868);
and UO_1272 (O_1272,N_9909,N_9905);
or UO_1273 (O_1273,N_9917,N_9947);
nor UO_1274 (O_1274,N_9868,N_9850);
nor UO_1275 (O_1275,N_9899,N_9852);
nor UO_1276 (O_1276,N_9877,N_9995);
nor UO_1277 (O_1277,N_9827,N_9864);
or UO_1278 (O_1278,N_9908,N_9921);
nor UO_1279 (O_1279,N_9987,N_9913);
and UO_1280 (O_1280,N_9964,N_9870);
nand UO_1281 (O_1281,N_9865,N_9944);
nand UO_1282 (O_1282,N_9889,N_9978);
and UO_1283 (O_1283,N_9990,N_9804);
nor UO_1284 (O_1284,N_9882,N_9876);
and UO_1285 (O_1285,N_9802,N_9890);
or UO_1286 (O_1286,N_9946,N_9883);
and UO_1287 (O_1287,N_9852,N_9901);
xor UO_1288 (O_1288,N_9996,N_9833);
nand UO_1289 (O_1289,N_9869,N_9845);
or UO_1290 (O_1290,N_9981,N_9914);
nand UO_1291 (O_1291,N_9939,N_9822);
or UO_1292 (O_1292,N_9932,N_9875);
nor UO_1293 (O_1293,N_9858,N_9960);
nand UO_1294 (O_1294,N_9862,N_9907);
nand UO_1295 (O_1295,N_9831,N_9895);
or UO_1296 (O_1296,N_9876,N_9960);
and UO_1297 (O_1297,N_9939,N_9959);
and UO_1298 (O_1298,N_9916,N_9931);
or UO_1299 (O_1299,N_9944,N_9971);
xor UO_1300 (O_1300,N_9885,N_9957);
or UO_1301 (O_1301,N_9960,N_9901);
or UO_1302 (O_1302,N_9968,N_9873);
or UO_1303 (O_1303,N_9859,N_9876);
nand UO_1304 (O_1304,N_9840,N_9890);
nand UO_1305 (O_1305,N_9921,N_9801);
or UO_1306 (O_1306,N_9975,N_9851);
nor UO_1307 (O_1307,N_9871,N_9816);
nand UO_1308 (O_1308,N_9947,N_9982);
and UO_1309 (O_1309,N_9909,N_9978);
nand UO_1310 (O_1310,N_9862,N_9937);
xnor UO_1311 (O_1311,N_9873,N_9839);
or UO_1312 (O_1312,N_9978,N_9914);
nor UO_1313 (O_1313,N_9950,N_9988);
and UO_1314 (O_1314,N_9849,N_9818);
and UO_1315 (O_1315,N_9826,N_9861);
or UO_1316 (O_1316,N_9897,N_9962);
or UO_1317 (O_1317,N_9853,N_9890);
or UO_1318 (O_1318,N_9816,N_9982);
nor UO_1319 (O_1319,N_9807,N_9985);
or UO_1320 (O_1320,N_9925,N_9976);
nor UO_1321 (O_1321,N_9972,N_9823);
and UO_1322 (O_1322,N_9894,N_9989);
or UO_1323 (O_1323,N_9835,N_9875);
nand UO_1324 (O_1324,N_9884,N_9967);
or UO_1325 (O_1325,N_9952,N_9901);
and UO_1326 (O_1326,N_9942,N_9821);
nor UO_1327 (O_1327,N_9926,N_9862);
or UO_1328 (O_1328,N_9804,N_9929);
nand UO_1329 (O_1329,N_9955,N_9962);
and UO_1330 (O_1330,N_9959,N_9911);
nand UO_1331 (O_1331,N_9915,N_9824);
or UO_1332 (O_1332,N_9995,N_9880);
or UO_1333 (O_1333,N_9814,N_9863);
nor UO_1334 (O_1334,N_9898,N_9956);
nand UO_1335 (O_1335,N_9962,N_9974);
nand UO_1336 (O_1336,N_9854,N_9936);
nor UO_1337 (O_1337,N_9919,N_9801);
and UO_1338 (O_1338,N_9857,N_9991);
nand UO_1339 (O_1339,N_9966,N_9893);
or UO_1340 (O_1340,N_9992,N_9817);
nor UO_1341 (O_1341,N_9936,N_9973);
and UO_1342 (O_1342,N_9850,N_9950);
or UO_1343 (O_1343,N_9835,N_9947);
xor UO_1344 (O_1344,N_9993,N_9912);
nand UO_1345 (O_1345,N_9914,N_9972);
and UO_1346 (O_1346,N_9974,N_9830);
or UO_1347 (O_1347,N_9868,N_9984);
and UO_1348 (O_1348,N_9966,N_9916);
or UO_1349 (O_1349,N_9947,N_9838);
nor UO_1350 (O_1350,N_9851,N_9828);
nand UO_1351 (O_1351,N_9801,N_9910);
xnor UO_1352 (O_1352,N_9940,N_9941);
nand UO_1353 (O_1353,N_9976,N_9944);
and UO_1354 (O_1354,N_9955,N_9987);
nand UO_1355 (O_1355,N_9862,N_9881);
xnor UO_1356 (O_1356,N_9815,N_9806);
and UO_1357 (O_1357,N_9848,N_9839);
xnor UO_1358 (O_1358,N_9914,N_9962);
nand UO_1359 (O_1359,N_9995,N_9822);
and UO_1360 (O_1360,N_9932,N_9896);
and UO_1361 (O_1361,N_9930,N_9924);
nand UO_1362 (O_1362,N_9814,N_9878);
and UO_1363 (O_1363,N_9929,N_9828);
or UO_1364 (O_1364,N_9968,N_9841);
nand UO_1365 (O_1365,N_9857,N_9825);
xor UO_1366 (O_1366,N_9996,N_9847);
or UO_1367 (O_1367,N_9976,N_9870);
and UO_1368 (O_1368,N_9934,N_9925);
xor UO_1369 (O_1369,N_9851,N_9983);
and UO_1370 (O_1370,N_9983,N_9928);
and UO_1371 (O_1371,N_9930,N_9816);
and UO_1372 (O_1372,N_9986,N_9978);
nor UO_1373 (O_1373,N_9893,N_9838);
nor UO_1374 (O_1374,N_9905,N_9992);
or UO_1375 (O_1375,N_9994,N_9845);
and UO_1376 (O_1376,N_9867,N_9982);
xor UO_1377 (O_1377,N_9876,N_9983);
nor UO_1378 (O_1378,N_9887,N_9988);
nand UO_1379 (O_1379,N_9814,N_9914);
nor UO_1380 (O_1380,N_9938,N_9860);
or UO_1381 (O_1381,N_9873,N_9901);
or UO_1382 (O_1382,N_9806,N_9879);
nand UO_1383 (O_1383,N_9926,N_9938);
or UO_1384 (O_1384,N_9951,N_9841);
and UO_1385 (O_1385,N_9831,N_9878);
nand UO_1386 (O_1386,N_9966,N_9930);
or UO_1387 (O_1387,N_9931,N_9914);
nor UO_1388 (O_1388,N_9937,N_9936);
nor UO_1389 (O_1389,N_9823,N_9847);
and UO_1390 (O_1390,N_9971,N_9905);
and UO_1391 (O_1391,N_9997,N_9818);
or UO_1392 (O_1392,N_9987,N_9997);
or UO_1393 (O_1393,N_9977,N_9910);
nor UO_1394 (O_1394,N_9837,N_9809);
nand UO_1395 (O_1395,N_9941,N_9803);
or UO_1396 (O_1396,N_9941,N_9807);
nor UO_1397 (O_1397,N_9841,N_9874);
xnor UO_1398 (O_1398,N_9939,N_9964);
xnor UO_1399 (O_1399,N_9881,N_9843);
or UO_1400 (O_1400,N_9945,N_9890);
nand UO_1401 (O_1401,N_9939,N_9925);
nor UO_1402 (O_1402,N_9850,N_9902);
nor UO_1403 (O_1403,N_9928,N_9984);
xnor UO_1404 (O_1404,N_9858,N_9841);
nand UO_1405 (O_1405,N_9963,N_9819);
nor UO_1406 (O_1406,N_9932,N_9993);
nand UO_1407 (O_1407,N_9860,N_9985);
and UO_1408 (O_1408,N_9857,N_9926);
and UO_1409 (O_1409,N_9847,N_9807);
xnor UO_1410 (O_1410,N_9868,N_9898);
xnor UO_1411 (O_1411,N_9844,N_9923);
and UO_1412 (O_1412,N_9901,N_9862);
nand UO_1413 (O_1413,N_9906,N_9946);
or UO_1414 (O_1414,N_9986,N_9826);
nand UO_1415 (O_1415,N_9897,N_9801);
xor UO_1416 (O_1416,N_9961,N_9873);
or UO_1417 (O_1417,N_9800,N_9868);
and UO_1418 (O_1418,N_9916,N_9998);
nand UO_1419 (O_1419,N_9839,N_9927);
and UO_1420 (O_1420,N_9800,N_9867);
or UO_1421 (O_1421,N_9824,N_9975);
and UO_1422 (O_1422,N_9906,N_9865);
nand UO_1423 (O_1423,N_9824,N_9809);
xnor UO_1424 (O_1424,N_9941,N_9992);
xnor UO_1425 (O_1425,N_9851,N_9883);
nor UO_1426 (O_1426,N_9923,N_9975);
nor UO_1427 (O_1427,N_9884,N_9877);
nand UO_1428 (O_1428,N_9991,N_9886);
nor UO_1429 (O_1429,N_9853,N_9919);
nor UO_1430 (O_1430,N_9830,N_9861);
and UO_1431 (O_1431,N_9806,N_9827);
nor UO_1432 (O_1432,N_9963,N_9985);
nor UO_1433 (O_1433,N_9952,N_9932);
and UO_1434 (O_1434,N_9980,N_9965);
nand UO_1435 (O_1435,N_9940,N_9915);
or UO_1436 (O_1436,N_9994,N_9905);
nand UO_1437 (O_1437,N_9873,N_9834);
nor UO_1438 (O_1438,N_9832,N_9929);
and UO_1439 (O_1439,N_9877,N_9898);
and UO_1440 (O_1440,N_9921,N_9870);
and UO_1441 (O_1441,N_9833,N_9878);
nor UO_1442 (O_1442,N_9835,N_9992);
or UO_1443 (O_1443,N_9820,N_9983);
or UO_1444 (O_1444,N_9951,N_9992);
nor UO_1445 (O_1445,N_9826,N_9823);
nor UO_1446 (O_1446,N_9911,N_9816);
or UO_1447 (O_1447,N_9822,N_9842);
or UO_1448 (O_1448,N_9931,N_9820);
nand UO_1449 (O_1449,N_9977,N_9828);
and UO_1450 (O_1450,N_9845,N_9968);
and UO_1451 (O_1451,N_9945,N_9952);
nor UO_1452 (O_1452,N_9877,N_9946);
and UO_1453 (O_1453,N_9841,N_9900);
nor UO_1454 (O_1454,N_9804,N_9837);
nor UO_1455 (O_1455,N_9876,N_9829);
nor UO_1456 (O_1456,N_9802,N_9875);
and UO_1457 (O_1457,N_9838,N_9903);
and UO_1458 (O_1458,N_9827,N_9929);
or UO_1459 (O_1459,N_9848,N_9942);
nand UO_1460 (O_1460,N_9802,N_9983);
xnor UO_1461 (O_1461,N_9892,N_9826);
nor UO_1462 (O_1462,N_9915,N_9842);
or UO_1463 (O_1463,N_9818,N_9890);
and UO_1464 (O_1464,N_9954,N_9858);
nand UO_1465 (O_1465,N_9861,N_9825);
and UO_1466 (O_1466,N_9880,N_9906);
or UO_1467 (O_1467,N_9978,N_9936);
and UO_1468 (O_1468,N_9999,N_9925);
nor UO_1469 (O_1469,N_9950,N_9990);
and UO_1470 (O_1470,N_9947,N_9848);
nand UO_1471 (O_1471,N_9819,N_9982);
nand UO_1472 (O_1472,N_9879,N_9973);
nand UO_1473 (O_1473,N_9818,N_9907);
nor UO_1474 (O_1474,N_9970,N_9945);
nor UO_1475 (O_1475,N_9807,N_9964);
nand UO_1476 (O_1476,N_9900,N_9958);
xnor UO_1477 (O_1477,N_9842,N_9872);
nor UO_1478 (O_1478,N_9929,N_9850);
or UO_1479 (O_1479,N_9946,N_9831);
or UO_1480 (O_1480,N_9807,N_9809);
nand UO_1481 (O_1481,N_9933,N_9946);
or UO_1482 (O_1482,N_9816,N_9818);
nor UO_1483 (O_1483,N_9995,N_9951);
or UO_1484 (O_1484,N_9931,N_9808);
and UO_1485 (O_1485,N_9969,N_9861);
and UO_1486 (O_1486,N_9822,N_9825);
nand UO_1487 (O_1487,N_9951,N_9875);
nor UO_1488 (O_1488,N_9960,N_9891);
xor UO_1489 (O_1489,N_9981,N_9831);
nor UO_1490 (O_1490,N_9925,N_9871);
nand UO_1491 (O_1491,N_9801,N_9883);
xor UO_1492 (O_1492,N_9969,N_9997);
nand UO_1493 (O_1493,N_9887,N_9934);
nand UO_1494 (O_1494,N_9932,N_9972);
nor UO_1495 (O_1495,N_9809,N_9944);
xnor UO_1496 (O_1496,N_9941,N_9995);
nor UO_1497 (O_1497,N_9951,N_9972);
nor UO_1498 (O_1498,N_9985,N_9878);
or UO_1499 (O_1499,N_9920,N_9901);
endmodule