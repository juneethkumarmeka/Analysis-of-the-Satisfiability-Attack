module basic_1500_15000_2000_15_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_1007,In_15);
or U1 (N_1,In_624,In_317);
xnor U2 (N_2,In_955,In_722);
or U3 (N_3,In_193,In_1306);
or U4 (N_4,In_804,In_417);
and U5 (N_5,In_358,In_3);
and U6 (N_6,In_54,In_1066);
or U7 (N_7,In_553,In_1405);
or U8 (N_8,In_983,In_1132);
and U9 (N_9,In_1087,In_503);
and U10 (N_10,In_461,In_492);
or U11 (N_11,In_780,In_1240);
or U12 (N_12,In_467,In_1068);
and U13 (N_13,In_177,In_717);
and U14 (N_14,In_1412,In_1138);
or U15 (N_15,In_96,In_622);
or U16 (N_16,In_950,In_607);
and U17 (N_17,In_39,In_189);
and U18 (N_18,In_816,In_221);
or U19 (N_19,In_336,In_677);
and U20 (N_20,In_604,In_1444);
and U21 (N_21,In_1318,In_1472);
xor U22 (N_22,In_850,In_835);
xor U23 (N_23,In_443,In_897);
nor U24 (N_24,In_1070,In_362);
or U25 (N_25,In_172,In_99);
xor U26 (N_26,In_1226,In_847);
or U27 (N_27,In_1057,In_646);
and U28 (N_28,In_206,In_222);
and U29 (N_29,In_1120,In_86);
or U30 (N_30,In_473,In_396);
nand U31 (N_31,In_185,In_1462);
and U32 (N_32,In_13,In_261);
and U33 (N_33,In_342,In_912);
xnor U34 (N_34,In_346,In_602);
and U35 (N_35,In_77,In_56);
nor U36 (N_36,In_877,In_1229);
nor U37 (N_37,In_989,In_1383);
xnor U38 (N_38,In_125,In_1496);
nand U39 (N_39,In_203,In_991);
xnor U40 (N_40,In_240,In_855);
nand U41 (N_41,In_628,In_1029);
xnor U42 (N_42,In_1117,In_630);
or U43 (N_43,In_80,In_1458);
nand U44 (N_44,In_1113,In_1036);
or U45 (N_45,In_739,In_851);
and U46 (N_46,In_1220,In_719);
and U47 (N_47,In_19,In_946);
and U48 (N_48,In_545,In_64);
or U49 (N_49,In_1034,In_139);
nor U50 (N_50,In_814,In_378);
nand U51 (N_51,In_369,In_482);
and U52 (N_52,In_759,In_1297);
nand U53 (N_53,In_270,In_149);
or U54 (N_54,In_665,In_238);
nor U55 (N_55,In_481,In_701);
and U56 (N_56,In_600,In_340);
nand U57 (N_57,In_913,In_1050);
or U58 (N_58,In_1244,In_640);
nand U59 (N_59,In_1468,In_1475);
nor U60 (N_60,In_1321,In_1353);
and U61 (N_61,In_401,In_7);
and U62 (N_62,In_612,In_598);
nand U63 (N_63,In_1079,In_1393);
nor U64 (N_64,In_1379,In_244);
nor U65 (N_65,In_988,In_144);
nor U66 (N_66,In_499,In_310);
nor U67 (N_67,In_1122,In_100);
nor U68 (N_68,In_813,In_1249);
nand U69 (N_69,In_351,In_10);
xnor U70 (N_70,In_159,In_936);
nand U71 (N_71,In_60,In_583);
nand U72 (N_72,In_1455,In_1267);
nand U73 (N_73,In_822,In_1433);
nor U74 (N_74,In_1337,In_446);
nor U75 (N_75,In_879,In_1390);
nand U76 (N_76,In_196,In_343);
xor U77 (N_77,In_275,In_366);
nor U78 (N_78,In_166,In_263);
nor U79 (N_79,In_1416,In_252);
nand U80 (N_80,In_668,In_315);
or U81 (N_81,In_382,In_994);
nor U82 (N_82,In_1016,In_954);
or U83 (N_83,In_757,In_1241);
nor U84 (N_84,In_1237,In_610);
and U85 (N_85,In_1258,In_1478);
and U86 (N_86,In_682,In_680);
or U87 (N_87,In_899,In_25);
nor U88 (N_88,In_1056,In_292);
nor U89 (N_89,In_30,In_1340);
and U90 (N_90,In_1260,In_241);
nand U91 (N_91,In_48,In_357);
or U92 (N_92,In_1217,In_1364);
xor U93 (N_93,In_324,In_675);
xor U94 (N_94,In_1310,In_632);
or U95 (N_95,In_517,In_471);
nand U96 (N_96,In_760,In_738);
and U97 (N_97,In_614,In_423);
or U98 (N_98,In_264,In_1439);
or U99 (N_99,In_1362,In_200);
nand U100 (N_100,In_255,In_1319);
xnor U101 (N_101,In_393,In_645);
and U102 (N_102,In_634,In_1428);
or U103 (N_103,In_114,In_724);
nor U104 (N_104,In_1161,In_654);
nor U105 (N_105,In_845,In_1219);
xnor U106 (N_106,In_692,In_1228);
nand U107 (N_107,In_367,In_1127);
and U108 (N_108,In_447,In_601);
nand U109 (N_109,In_1320,In_1130);
and U110 (N_110,In_1373,In_1247);
and U111 (N_111,In_704,In_697);
nor U112 (N_112,In_45,In_307);
and U113 (N_113,In_844,In_771);
or U114 (N_114,In_440,In_1135);
nand U115 (N_115,In_1252,In_18);
nand U116 (N_116,In_171,In_1427);
and U117 (N_117,In_237,In_78);
nor U118 (N_118,In_1104,In_1180);
nor U119 (N_119,In_1111,In_1043);
or U120 (N_120,In_463,In_79);
nand U121 (N_121,In_773,In_1346);
or U122 (N_122,In_1191,In_1261);
or U123 (N_123,In_1401,In_158);
or U124 (N_124,In_1304,In_165);
and U125 (N_125,In_702,In_885);
and U126 (N_126,In_176,In_1243);
or U127 (N_127,In_348,In_987);
or U128 (N_128,In_993,In_1095);
nand U129 (N_129,In_948,In_647);
nor U130 (N_130,In_548,In_1133);
or U131 (N_131,In_860,In_1227);
or U132 (N_132,In_297,In_454);
xor U133 (N_133,In_1316,In_1372);
nand U134 (N_134,In_190,In_1403);
or U135 (N_135,In_468,In_391);
nor U136 (N_136,In_1285,In_934);
and U137 (N_137,In_91,In_1188);
or U138 (N_138,In_428,In_1162);
and U139 (N_139,In_1268,In_1042);
or U140 (N_140,In_865,In_1266);
or U141 (N_141,In_671,In_1305);
and U142 (N_142,In_1051,In_713);
nor U143 (N_143,In_82,In_429);
nor U144 (N_144,In_737,In_872);
and U145 (N_145,In_643,In_497);
and U146 (N_146,In_41,In_1435);
xnor U147 (N_147,In_689,In_599);
nor U148 (N_148,In_389,In_123);
and U149 (N_149,In_1485,In_1361);
or U150 (N_150,In_1011,In_1420);
nand U151 (N_151,In_873,In_910);
nand U152 (N_152,In_696,In_1271);
and U153 (N_153,In_810,In_1015);
nor U154 (N_154,In_145,In_1174);
nand U155 (N_155,In_333,In_652);
or U156 (N_156,In_909,In_280);
or U157 (N_157,In_1441,In_323);
nand U158 (N_158,In_731,In_431);
nand U159 (N_159,In_586,In_1296);
xnor U160 (N_160,In_354,In_66);
nand U161 (N_161,In_735,In_313);
xor U162 (N_162,In_146,In_1445);
and U163 (N_163,In_1024,In_707);
nor U164 (N_164,In_422,In_450);
and U165 (N_165,In_706,In_136);
nor U166 (N_166,In_188,In_65);
xnor U167 (N_167,In_1169,In_1131);
nor U168 (N_168,In_304,In_558);
nor U169 (N_169,In_282,In_435);
nor U170 (N_170,In_1473,In_711);
nand U171 (N_171,In_901,In_57);
nand U172 (N_172,In_939,In_83);
nor U173 (N_173,In_488,In_819);
nand U174 (N_174,In_220,In_720);
or U175 (N_175,In_1023,In_1457);
or U176 (N_176,In_449,In_1397);
nor U177 (N_177,In_225,In_526);
nand U178 (N_178,In_131,In_1239);
nor U179 (N_179,In_1425,In_1067);
nor U180 (N_180,In_831,In_1436);
and U181 (N_181,In_808,In_637);
and U182 (N_182,In_26,In_8);
nor U183 (N_183,In_809,In_1380);
and U184 (N_184,In_1317,In_1215);
nand U185 (N_185,In_444,In_1018);
nand U186 (N_186,In_1109,In_1012);
nand U187 (N_187,In_1286,In_1146);
nor U188 (N_188,In_1308,In_807);
or U189 (N_189,In_1218,In_195);
nor U190 (N_190,In_876,In_736);
or U191 (N_191,In_953,In_615);
and U192 (N_192,In_337,In_734);
and U193 (N_193,In_1335,In_356);
nor U194 (N_194,In_900,In_260);
and U195 (N_195,In_53,In_314);
and U196 (N_196,In_1126,In_477);
nand U197 (N_197,In_1288,In_664);
nor U198 (N_198,In_888,In_565);
and U199 (N_199,In_439,In_1437);
xor U200 (N_200,In_1028,In_981);
nor U201 (N_201,In_984,In_515);
and U202 (N_202,In_688,In_1214);
nor U203 (N_203,In_636,In_148);
or U204 (N_204,In_300,In_1384);
and U205 (N_205,In_1287,In_779);
nor U206 (N_206,In_920,In_533);
nor U207 (N_207,In_725,In_75);
and U208 (N_208,In_1086,In_208);
or U209 (N_209,In_1008,In_1369);
or U210 (N_210,In_17,In_386);
nor U211 (N_211,In_996,In_162);
nand U212 (N_212,In_613,In_432);
nand U213 (N_213,In_588,In_1482);
and U214 (N_214,In_529,In_1470);
and U215 (N_215,In_124,In_320);
nor U216 (N_216,In_498,In_922);
or U217 (N_217,In_1303,In_1498);
or U218 (N_218,In_718,In_93);
or U219 (N_219,In_364,In_424);
nand U220 (N_220,In_1031,In_522);
or U221 (N_221,In_1178,In_1114);
or U222 (N_222,In_782,In_334);
nand U223 (N_223,In_288,In_254);
and U224 (N_224,In_1115,In_1005);
nand U225 (N_225,In_55,In_1495);
nand U226 (N_226,In_960,In_1484);
xnor U227 (N_227,In_1269,In_1155);
and U228 (N_228,In_1238,In_11);
nand U229 (N_229,In_730,In_50);
nand U230 (N_230,In_698,In_1233);
nor U231 (N_231,In_575,In_1391);
nor U232 (N_232,In_452,In_486);
or U233 (N_233,In_1449,In_1476);
xor U234 (N_234,In_906,In_1366);
nor U235 (N_235,In_308,In_29);
nand U236 (N_236,In_377,In_669);
xnor U237 (N_237,In_1058,In_319);
and U238 (N_238,In_217,In_205);
or U239 (N_239,In_1329,In_284);
and U240 (N_240,In_426,In_619);
xnor U241 (N_241,In_1469,In_49);
nor U242 (N_242,In_95,In_705);
nor U243 (N_243,In_410,In_1082);
nor U244 (N_244,In_101,In_418);
xnor U245 (N_245,In_1448,In_213);
xor U246 (N_246,In_1325,In_1078);
or U247 (N_247,In_1466,In_1017);
xnor U248 (N_248,In_1338,In_562);
or U249 (N_249,In_122,In_1387);
nand U250 (N_250,In_778,In_107);
or U251 (N_251,In_311,In_1374);
nand U252 (N_252,In_1084,In_249);
or U253 (N_253,In_327,In_69);
nand U254 (N_254,In_1112,In_1276);
or U255 (N_255,In_1370,In_925);
or U256 (N_256,In_714,In_233);
nor U257 (N_257,In_67,In_1302);
nand U258 (N_258,In_258,In_798);
and U259 (N_259,In_1004,In_1153);
and U260 (N_260,In_1163,In_539);
or U261 (N_261,In_801,In_1207);
and U262 (N_262,In_1460,In_44);
or U263 (N_263,In_866,In_456);
or U264 (N_264,In_512,In_1002);
or U265 (N_265,In_1110,In_1356);
nor U266 (N_266,In_579,In_178);
nand U267 (N_267,In_708,In_1407);
nand U268 (N_268,In_937,In_974);
and U269 (N_269,In_928,In_802);
and U270 (N_270,In_384,In_580);
or U271 (N_271,In_863,In_700);
and U272 (N_272,In_1290,In_202);
nand U273 (N_273,In_113,In_803);
nand U274 (N_274,In_1211,In_1328);
nor U275 (N_275,In_40,In_880);
nor U276 (N_276,In_658,In_427);
and U277 (N_277,In_1280,In_137);
nand U278 (N_278,In_965,In_929);
or U279 (N_279,In_1025,In_1279);
or U280 (N_280,In_1432,In_1020);
and U281 (N_281,In_694,In_1254);
and U282 (N_282,In_1388,In_820);
nand U283 (N_283,In_678,In_1422);
nand U284 (N_284,In_861,In_608);
nand U285 (N_285,In_1242,In_889);
nor U286 (N_286,In_651,In_1019);
and U287 (N_287,In_777,In_1201);
or U288 (N_288,In_296,In_584);
and U289 (N_289,In_1499,In_187);
and U290 (N_290,In_1168,In_1000);
nand U291 (N_291,In_127,In_1093);
xnor U292 (N_292,In_849,In_1);
or U293 (N_293,In_554,In_672);
nand U294 (N_294,In_893,In_46);
or U295 (N_295,In_715,In_1077);
and U296 (N_296,In_359,In_236);
nor U297 (N_297,In_1404,In_374);
nand U298 (N_298,In_753,In_1322);
nor U299 (N_299,In_138,In_103);
or U300 (N_300,In_1144,In_226);
or U301 (N_301,In_952,In_1481);
or U302 (N_302,In_246,In_650);
nand U303 (N_303,In_457,In_1486);
nand U304 (N_304,In_1124,In_1143);
or U305 (N_305,In_1172,In_52);
nor U306 (N_306,In_1063,In_504);
or U307 (N_307,In_881,In_1368);
nand U308 (N_308,In_977,In_500);
nand U309 (N_309,In_116,In_505);
nor U310 (N_310,In_478,In_1136);
xnor U311 (N_311,In_433,In_430);
and U312 (N_312,In_997,In_390);
nand U313 (N_313,In_420,In_1193);
xor U314 (N_314,In_243,In_381);
nor U315 (N_315,In_1152,In_117);
or U316 (N_316,In_1053,In_1141);
and U317 (N_317,In_1300,In_1467);
and U318 (N_318,In_521,In_1206);
nor U319 (N_319,In_1440,In_963);
and U320 (N_320,In_1105,In_531);
nor U321 (N_321,In_230,In_1293);
nand U322 (N_322,In_277,In_578);
nor U323 (N_323,In_170,In_279);
xor U324 (N_324,In_918,In_0);
and U325 (N_325,In_1332,In_289);
nand U326 (N_326,In_886,In_514);
or U327 (N_327,In_1209,In_520);
nor U328 (N_328,In_774,In_161);
nand U329 (N_329,In_1097,In_594);
nand U330 (N_330,In_527,In_1071);
or U331 (N_331,In_685,In_33);
or U332 (N_332,In_1176,In_1424);
and U333 (N_333,In_405,In_903);
nand U334 (N_334,In_815,In_1157);
nor U335 (N_335,In_837,In_84);
or U336 (N_336,In_829,In_676);
xor U337 (N_337,In_1116,In_1224);
and U338 (N_338,In_1147,In_1001);
xnor U339 (N_339,In_787,In_940);
nand U340 (N_340,In_540,In_400);
nand U341 (N_341,In_616,In_834);
nand U342 (N_342,In_419,In_765);
nand U343 (N_343,In_1107,In_1182);
xor U344 (N_344,In_490,In_1336);
or U345 (N_345,In_878,In_415);
xnor U346 (N_346,In_1396,In_458);
nand U347 (N_347,In_394,In_218);
xor U348 (N_348,In_569,In_180);
and U349 (N_349,In_1376,In_181);
nor U350 (N_350,In_566,In_1076);
or U351 (N_351,In_1434,In_154);
nor U352 (N_352,In_824,In_541);
and U353 (N_353,In_789,In_1159);
or U354 (N_354,In_535,In_1489);
and U355 (N_355,In_1171,In_85);
nand U356 (N_356,In_644,In_194);
xnor U357 (N_357,In_979,In_322);
or U358 (N_358,In_530,In_1186);
and U359 (N_359,In_1274,In_16);
nor U360 (N_360,In_756,In_1072);
and U361 (N_361,In_1378,In_413);
nor U362 (N_362,In_510,In_1045);
nand U363 (N_363,In_1041,In_931);
or U364 (N_364,In_968,In_110);
nand U365 (N_365,In_1208,In_408);
nor U366 (N_366,In_1118,In_1375);
and U367 (N_367,In_1343,In_466);
or U368 (N_368,In_1301,In_235);
and U369 (N_369,In_1483,In_331);
and U370 (N_370,In_1101,In_462);
or U371 (N_371,In_999,In_1006);
and U372 (N_372,In_383,In_716);
nor U373 (N_373,In_796,In_199);
xnor U374 (N_374,In_784,In_582);
nand U375 (N_375,In_1426,In_309);
or U376 (N_376,In_51,In_1044);
nor U377 (N_377,In_88,In_128);
nor U378 (N_378,In_32,In_2);
nor U379 (N_379,In_355,In_1327);
nand U380 (N_380,In_465,In_479);
or U381 (N_381,In_751,In_215);
and U382 (N_382,In_932,In_484);
or U383 (N_383,In_1281,In_776);
nor U384 (N_384,In_1234,In_231);
nand U385 (N_385,In_299,In_684);
or U386 (N_386,In_421,In_763);
nand U387 (N_387,In_224,In_414);
or U388 (N_388,In_61,In_76);
nand U389 (N_389,In_92,In_755);
nor U390 (N_390,In_63,In_1463);
nand U391 (N_391,In_892,In_794);
and U392 (N_392,In_972,In_980);
or U393 (N_393,In_1395,In_248);
nor U394 (N_394,In_287,In_133);
nand U395 (N_395,In_740,In_617);
or U396 (N_396,In_890,In_1221);
nand U397 (N_397,In_1394,In_1350);
and U398 (N_398,In_480,In_818);
xnor U399 (N_399,In_1264,In_1265);
nand U400 (N_400,In_6,In_469);
or U401 (N_401,In_1245,In_821);
and U402 (N_402,In_347,In_112);
or U403 (N_403,In_805,In_1365);
and U404 (N_404,In_1413,In_1456);
nand U405 (N_405,In_869,In_1014);
or U406 (N_406,In_961,In_1289);
nand U407 (N_407,In_1179,In_1357);
nor U408 (N_408,In_1085,In_1190);
xor U409 (N_409,In_1282,In_27);
and U410 (N_410,In_1106,In_268);
or U411 (N_411,In_896,In_129);
or U412 (N_412,In_552,In_674);
and U413 (N_413,In_1270,In_693);
and U414 (N_414,In_1194,In_1073);
nand U415 (N_415,In_967,In_326);
and U416 (N_416,In_1040,In_251);
nand U417 (N_417,In_219,In_1345);
nor U418 (N_418,In_38,In_549);
nor U419 (N_419,In_155,In_352);
or U420 (N_420,In_1342,In_1339);
nor U421 (N_421,In_792,In_1200);
nand U422 (N_422,In_570,In_387);
and U423 (N_423,In_403,In_1415);
nand U424 (N_424,In_1213,In_1490);
nor U425 (N_425,In_164,In_22);
or U426 (N_426,In_551,In_135);
nor U427 (N_427,In_1398,In_1400);
and U428 (N_428,In_1263,In_68);
and U429 (N_429,In_281,In_1236);
or U430 (N_430,In_325,In_841);
and U431 (N_431,In_550,In_1096);
xor U432 (N_432,In_978,In_1223);
or U433 (N_433,In_1069,In_212);
and U434 (N_434,In_269,In_1351);
nand U435 (N_435,In_204,In_507);
or U436 (N_436,In_111,In_1352);
or U437 (N_437,In_302,In_1360);
nand U438 (N_438,In_791,In_924);
nand U439 (N_439,In_1430,In_524);
or U440 (N_440,In_1102,In_797);
nand U441 (N_441,In_843,In_295);
and U442 (N_442,In_303,In_769);
or U443 (N_443,In_595,In_721);
nand U444 (N_444,In_970,In_43);
or U445 (N_445,In_1294,In_795);
and U446 (N_446,In_1283,In_9);
and U447 (N_447,In_1326,In_670);
and U448 (N_448,In_376,In_1148);
nor U449 (N_449,In_338,In_1185);
nand U450 (N_450,In_1421,In_1442);
nor U451 (N_451,In_312,In_259);
nand U452 (N_452,In_663,In_72);
and U453 (N_453,In_157,In_817);
and U454 (N_454,In_1037,In_151);
or U455 (N_455,In_1443,In_656);
nor U456 (N_456,In_276,In_1021);
and U457 (N_457,In_360,In_1222);
nand U458 (N_458,In_908,In_848);
nand U459 (N_459,In_790,In_611);
nand U460 (N_460,In_1108,In_1202);
and U461 (N_461,In_605,In_898);
nand U462 (N_462,In_140,In_1103);
or U463 (N_463,In_621,In_294);
and U464 (N_464,In_770,In_102);
and U465 (N_465,In_168,In_945);
xnor U466 (N_466,In_105,In_1091);
nand U467 (N_467,In_653,In_732);
and U468 (N_468,In_555,In_97);
nand U469 (N_469,In_661,In_286);
nor U470 (N_470,In_1386,In_126);
xnor U471 (N_471,In_1480,In_1088);
or U472 (N_472,In_576,In_830);
and U473 (N_473,In_862,In_1100);
nand U474 (N_474,In_710,In_935);
nor U475 (N_475,In_345,In_662);
and U476 (N_476,In_70,In_250);
nand U477 (N_477,In_1027,In_1477);
or U478 (N_478,In_1248,In_1464);
and U479 (N_479,In_856,In_464);
nor U480 (N_480,In_655,In_1454);
nand U481 (N_481,In_494,In_975);
and U482 (N_482,In_641,In_470);
nand U483 (N_483,In_733,In_455);
and U484 (N_484,In_1198,In_686);
nand U485 (N_485,In_1140,In_556);
xnor U486 (N_486,In_927,In_130);
and U487 (N_487,In_546,In_832);
or U488 (N_488,In_772,In_1173);
and U489 (N_489,In_58,In_626);
nor U490 (N_490,In_1491,In_916);
nor U491 (N_491,In_160,In_589);
or U492 (N_492,In_1341,In_1013);
nor U493 (N_493,In_748,In_635);
nand U494 (N_494,In_228,In_859);
xor U495 (N_495,In_373,In_854);
and U496 (N_496,In_867,In_174);
or U497 (N_497,In_47,In_1035);
and U498 (N_498,In_1312,In_506);
nor U499 (N_499,In_214,In_372);
nor U500 (N_500,In_585,In_852);
nor U501 (N_501,In_1246,In_1164);
and U502 (N_502,In_353,In_673);
or U503 (N_503,In_581,In_256);
or U504 (N_504,In_823,In_1094);
nor U505 (N_505,In_175,In_754);
and U506 (N_506,In_919,In_853);
nand U507 (N_507,In_547,In_472);
and U508 (N_508,In_34,In_328);
or U509 (N_509,In_385,In_609);
nor U510 (N_510,In_329,In_1061);
and U511 (N_511,In_926,In_964);
and U512 (N_512,In_887,In_907);
nor U513 (N_513,In_679,In_1177);
or U514 (N_514,In_758,In_5);
xnor U515 (N_515,In_37,In_411);
and U516 (N_516,In_1392,In_560);
nor U517 (N_517,In_321,In_1026);
or U518 (N_518,In_828,In_1417);
xnor U519 (N_519,In_152,In_475);
nor U520 (N_520,In_659,In_474);
xnor U521 (N_521,In_842,In_1196);
or U522 (N_522,In_271,In_1154);
xor U523 (N_523,In_460,In_1052);
nand U524 (N_524,In_1402,In_606);
or U525 (N_525,In_836,In_891);
xor U526 (N_526,In_573,In_209);
nand U527 (N_527,In_1235,In_409);
xnor U528 (N_528,In_742,In_1183);
or U529 (N_529,In_211,In_559);
nand U530 (N_530,In_253,In_120);
nand U531 (N_531,In_593,In_745);
xor U532 (N_532,In_1359,In_1408);
and U533 (N_533,In_1151,In_59);
and U534 (N_534,In_192,In_501);
and U535 (N_535,In_150,In_20);
nor U536 (N_536,In_257,In_266);
nand U537 (N_537,In_245,In_509);
or U538 (N_538,In_783,In_316);
xnor U539 (N_539,In_712,In_169);
or U540 (N_540,In_274,In_639);
nor U541 (N_541,In_242,In_603);
nor U542 (N_542,In_1331,In_538);
and U543 (N_543,In_1048,In_528);
nand U544 (N_544,In_523,In_1358);
xor U545 (N_545,In_108,In_143);
nand U546 (N_546,In_1446,In_207);
nand U547 (N_547,In_642,In_163);
and U548 (N_548,In_71,In_184);
nor U549 (N_549,In_201,In_833);
nor U550 (N_550,In_827,In_21);
or U551 (N_551,In_511,In_398);
nand U552 (N_552,In_1459,In_298);
nor U553 (N_553,In_923,In_1277);
or U554 (N_554,In_884,In_445);
and U555 (N_555,In_365,In_567);
nor U556 (N_556,In_1251,In_534);
nand U557 (N_557,In_564,In_1210);
nand U558 (N_558,In_1291,In_1431);
or U559 (N_559,In_917,In_476);
and U560 (N_560,In_1089,In_436);
and U561 (N_561,In_285,In_434);
nor U562 (N_562,In_412,In_544);
and U563 (N_563,In_825,In_1059);
nand U564 (N_564,In_90,In_1074);
and U565 (N_565,In_516,In_167);
nand U566 (N_566,In_1129,In_89);
nand U567 (N_567,In_191,In_683);
and U568 (N_568,In_747,In_762);
nand U569 (N_569,In_775,In_1165);
xor U570 (N_570,In_638,In_1203);
nand U571 (N_571,In_1046,In_868);
nand U572 (N_572,In_94,In_1205);
nand U573 (N_573,In_73,In_1349);
nand U574 (N_574,In_1160,In_1175);
nor U575 (N_575,In_561,In_330);
nand U576 (N_576,In_1354,In_633);
nand U577 (N_577,In_451,In_938);
nand U578 (N_578,In_691,In_727);
nor U579 (N_579,In_1170,In_508);
nor U580 (N_580,In_1487,In_1314);
nand U581 (N_581,In_404,In_1465);
or U582 (N_582,In_930,In_915);
nor U583 (N_583,In_141,In_749);
nand U584 (N_584,In_1324,In_625);
or U585 (N_585,In_951,In_1275);
or U586 (N_586,In_800,In_1080);
and U587 (N_587,In_459,In_741);
nor U588 (N_588,In_489,In_1121);
and U589 (N_589,In_681,In_1429);
nor U590 (N_590,In_687,In_132);
xor U591 (N_591,In_1299,In_998);
nor U592 (N_592,In_631,In_262);
and U593 (N_593,In_379,In_1414);
xnor U594 (N_594,In_1158,In_1039);
nor U595 (N_595,In_563,In_1295);
and U596 (N_596,In_239,In_272);
xor U597 (N_597,In_947,In_437);
and U598 (N_598,In_349,In_1181);
and U599 (N_599,In_42,In_31);
and U600 (N_600,In_992,In_183);
nor U601 (N_601,In_596,In_438);
nor U602 (N_602,In_870,In_1399);
nand U603 (N_603,In_1452,In_198);
nor U604 (N_604,In_623,In_493);
nor U605 (N_605,In_491,In_1255);
nand U606 (N_606,In_1347,In_1030);
or U607 (N_607,In_806,In_1389);
nor U608 (N_608,In_119,In_1334);
nand U609 (N_609,In_1192,In_657);
nor U610 (N_610,In_28,In_995);
nor U611 (N_611,In_723,In_227);
nor U612 (N_612,In_1410,In_874);
xor U613 (N_613,In_858,In_416);
nand U614 (N_614,In_905,In_557);
or U615 (N_615,In_267,In_1493);
nor U616 (N_616,In_290,In_1292);
nor U617 (N_617,In_388,In_441);
nor U618 (N_618,In_1232,In_12);
and U619 (N_619,In_1333,In_1166);
nor U620 (N_620,In_306,In_1257);
xor U621 (N_621,In_1125,In_990);
and U622 (N_622,In_1038,In_332);
nand U623 (N_623,In_966,In_1381);
nand U624 (N_624,In_1055,In_1212);
nand U625 (N_625,In_425,In_1075);
xnor U626 (N_626,In_1259,In_752);
and U627 (N_627,In_4,In_895);
nand U628 (N_628,In_1184,In_293);
xnor U629 (N_629,In_448,In_532);
or U630 (N_630,In_1010,In_1479);
or U631 (N_631,In_1330,In_406);
nor U632 (N_632,In_666,In_962);
and U633 (N_633,In_703,In_911);
and U634 (N_634,In_1447,In_210);
nor U635 (N_635,In_442,In_1060);
nand U636 (N_636,In_1311,In_24);
or U637 (N_637,In_1156,In_115);
nand U638 (N_638,In_1423,In_1216);
or U639 (N_639,In_106,In_883);
and U640 (N_640,In_1497,In_537);
and U641 (N_641,In_781,In_620);
or U642 (N_642,In_87,In_153);
xor U643 (N_643,In_1256,In_1262);
and U644 (N_644,In_1461,In_1099);
or U645 (N_645,In_921,In_375);
xor U646 (N_646,In_1298,In_147);
nor U647 (N_647,In_982,In_971);
or U648 (N_648,In_216,In_1047);
xor U649 (N_649,In_914,In_104);
or U650 (N_650,In_1062,In_695);
and U651 (N_651,In_496,In_1123);
or U652 (N_652,In_483,In_247);
and U653 (N_653,In_1199,In_986);
and U654 (N_654,In_976,In_392);
and U655 (N_655,In_785,In_1385);
nand U656 (N_656,In_956,In_1250);
nor U657 (N_657,In_957,In_812);
nor U658 (N_658,In_1418,In_649);
or U659 (N_659,In_943,In_648);
nand U660 (N_660,In_959,In_363);
nand U661 (N_661,In_283,In_399);
nand U662 (N_662,In_402,In_1145);
or U663 (N_663,In_1187,In_495);
nand U664 (N_664,In_571,In_942);
xor U665 (N_665,In_453,In_1090);
nor U666 (N_666,In_902,In_1438);
or U667 (N_667,In_1142,In_371);
nand U668 (N_668,In_1377,In_592);
nand U669 (N_669,In_1065,In_182);
nand U670 (N_670,In_629,In_1315);
nand U671 (N_671,In_525,In_1273);
xor U672 (N_672,In_840,In_339);
or U673 (N_673,In_291,In_36);
and U674 (N_674,In_699,In_1009);
xor U675 (N_675,In_572,In_1230);
nand U676 (N_676,In_1137,In_944);
or U677 (N_677,In_1409,In_743);
or U678 (N_678,In_904,In_766);
or U679 (N_679,In_341,In_318);
nor U680 (N_680,In_1225,In_941);
nor U681 (N_681,In_1453,In_109);
or U682 (N_682,In_380,In_23);
or U683 (N_683,In_871,In_1344);
nand U684 (N_684,In_973,In_660);
xor U685 (N_685,In_361,In_591);
or U686 (N_686,In_587,In_1128);
and U687 (N_687,In_519,In_857);
and U688 (N_688,In_969,In_265);
and U689 (N_689,In_1411,In_395);
and U690 (N_690,In_1406,In_397);
and U691 (N_691,In_1471,In_407);
nand U692 (N_692,In_1092,In_767);
xor U693 (N_693,In_1049,In_502);
nor U694 (N_694,In_1003,In_568);
or U695 (N_695,In_368,In_933);
or U696 (N_696,In_14,In_746);
nor U697 (N_697,In_1363,In_882);
and U698 (N_698,In_864,In_786);
nor U699 (N_699,In_536,In_846);
or U700 (N_700,In_811,In_1419);
nor U701 (N_701,In_597,In_1197);
and U702 (N_702,In_1382,In_1189);
nor U703 (N_703,In_350,In_1278);
nor U704 (N_704,In_1371,In_335);
and U705 (N_705,In_1309,In_1451);
nand U706 (N_706,In_799,In_1033);
or U707 (N_707,In_118,In_81);
nor U708 (N_708,In_761,In_1313);
nor U709 (N_709,In_35,In_958);
or U710 (N_710,In_543,In_764);
or U711 (N_711,In_728,In_1167);
nor U712 (N_712,In_1307,In_788);
and U713 (N_713,In_1204,In_62);
nor U714 (N_714,In_1022,In_826);
or U715 (N_715,In_709,In_590);
or U716 (N_716,In_1323,In_186);
and U717 (N_717,In_197,In_179);
nand U718 (N_718,In_750,In_577);
or U719 (N_719,In_618,In_690);
nor U720 (N_720,In_793,In_1488);
nor U721 (N_721,In_98,In_729);
nand U722 (N_722,In_894,In_1494);
and U723 (N_723,In_518,In_1134);
nand U724 (N_724,In_1348,In_1450);
and U725 (N_725,In_301,In_1081);
and U726 (N_726,In_1098,In_1195);
and U727 (N_727,In_838,In_1231);
and U728 (N_728,In_370,In_1367);
nand U729 (N_729,In_744,In_1284);
or U730 (N_730,In_985,In_74);
or U731 (N_731,In_344,In_121);
xnor U732 (N_732,In_949,In_134);
or U733 (N_733,In_1083,In_1054);
nand U734 (N_734,In_273,In_1139);
nand U735 (N_735,In_542,In_1150);
and U736 (N_736,In_1355,In_1064);
and U737 (N_737,In_223,In_1474);
and U738 (N_738,In_875,In_1149);
and U739 (N_739,In_627,In_229);
xnor U740 (N_740,In_305,In_278);
nand U741 (N_741,In_232,In_234);
nand U742 (N_742,In_485,In_574);
or U743 (N_743,In_173,In_768);
nor U744 (N_744,In_1032,In_1253);
and U745 (N_745,In_142,In_1492);
or U746 (N_746,In_1119,In_726);
xnor U747 (N_747,In_156,In_839);
nor U748 (N_748,In_487,In_513);
nor U749 (N_749,In_1272,In_667);
nor U750 (N_750,In_173,In_258);
and U751 (N_751,In_198,In_1303);
nand U752 (N_752,In_1492,In_1478);
nand U753 (N_753,In_156,In_1146);
or U754 (N_754,In_159,In_1113);
nand U755 (N_755,In_702,In_420);
and U756 (N_756,In_702,In_599);
and U757 (N_757,In_210,In_855);
nand U758 (N_758,In_739,In_1001);
xnor U759 (N_759,In_974,In_1008);
nor U760 (N_760,In_287,In_1151);
nand U761 (N_761,In_1435,In_11);
nand U762 (N_762,In_1178,In_1007);
and U763 (N_763,In_845,In_747);
and U764 (N_764,In_417,In_27);
nand U765 (N_765,In_448,In_188);
nand U766 (N_766,In_771,In_220);
and U767 (N_767,In_1341,In_1057);
nand U768 (N_768,In_937,In_1060);
nor U769 (N_769,In_1026,In_1458);
xor U770 (N_770,In_1145,In_787);
or U771 (N_771,In_473,In_1443);
nor U772 (N_772,In_1190,In_1042);
nand U773 (N_773,In_432,In_1224);
nand U774 (N_774,In_969,In_213);
xnor U775 (N_775,In_816,In_601);
nand U776 (N_776,In_911,In_68);
nor U777 (N_777,In_851,In_1374);
xnor U778 (N_778,In_71,In_1122);
nand U779 (N_779,In_1205,In_1335);
nand U780 (N_780,In_1101,In_1004);
nand U781 (N_781,In_1475,In_1434);
nand U782 (N_782,In_363,In_671);
nor U783 (N_783,In_452,In_891);
nor U784 (N_784,In_1326,In_726);
nor U785 (N_785,In_1312,In_1440);
nand U786 (N_786,In_870,In_901);
or U787 (N_787,In_448,In_203);
nor U788 (N_788,In_1168,In_1394);
and U789 (N_789,In_1147,In_884);
or U790 (N_790,In_969,In_974);
and U791 (N_791,In_877,In_303);
nand U792 (N_792,In_1327,In_444);
xor U793 (N_793,In_873,In_956);
xor U794 (N_794,In_1294,In_1230);
and U795 (N_795,In_1088,In_714);
or U796 (N_796,In_1294,In_256);
or U797 (N_797,In_667,In_1113);
or U798 (N_798,In_310,In_324);
and U799 (N_799,In_1207,In_147);
and U800 (N_800,In_1435,In_57);
xor U801 (N_801,In_1114,In_1281);
nand U802 (N_802,In_966,In_137);
and U803 (N_803,In_1012,In_1431);
or U804 (N_804,In_1143,In_1310);
or U805 (N_805,In_1458,In_1065);
and U806 (N_806,In_617,In_1091);
nand U807 (N_807,In_134,In_1340);
nand U808 (N_808,In_785,In_532);
nor U809 (N_809,In_101,In_1292);
nand U810 (N_810,In_1310,In_41);
nor U811 (N_811,In_602,In_264);
nor U812 (N_812,In_515,In_362);
nand U813 (N_813,In_1056,In_651);
or U814 (N_814,In_1026,In_1191);
nor U815 (N_815,In_1391,In_600);
nor U816 (N_816,In_353,In_1425);
nand U817 (N_817,In_820,In_634);
xnor U818 (N_818,In_1369,In_926);
and U819 (N_819,In_526,In_68);
nor U820 (N_820,In_1186,In_1338);
nand U821 (N_821,In_230,In_1006);
or U822 (N_822,In_552,In_341);
nand U823 (N_823,In_1122,In_553);
nor U824 (N_824,In_624,In_1245);
or U825 (N_825,In_290,In_711);
or U826 (N_826,In_1114,In_112);
or U827 (N_827,In_759,In_543);
or U828 (N_828,In_1224,In_1142);
or U829 (N_829,In_1050,In_849);
and U830 (N_830,In_881,In_642);
nand U831 (N_831,In_139,In_1230);
nand U832 (N_832,In_1356,In_1243);
nand U833 (N_833,In_20,In_571);
and U834 (N_834,In_731,In_302);
nor U835 (N_835,In_1487,In_936);
nor U836 (N_836,In_716,In_166);
nand U837 (N_837,In_310,In_1219);
nand U838 (N_838,In_1485,In_1016);
and U839 (N_839,In_1386,In_959);
or U840 (N_840,In_98,In_671);
nand U841 (N_841,In_123,In_1203);
xnor U842 (N_842,In_583,In_1229);
nor U843 (N_843,In_594,In_1338);
nor U844 (N_844,In_1353,In_1163);
nor U845 (N_845,In_35,In_1496);
nor U846 (N_846,In_53,In_942);
nand U847 (N_847,In_212,In_1248);
or U848 (N_848,In_1453,In_432);
and U849 (N_849,In_693,In_1038);
nand U850 (N_850,In_113,In_185);
nor U851 (N_851,In_1269,In_340);
xnor U852 (N_852,In_1275,In_355);
and U853 (N_853,In_1297,In_27);
xnor U854 (N_854,In_57,In_263);
or U855 (N_855,In_809,In_640);
nor U856 (N_856,In_258,In_992);
xnor U857 (N_857,In_980,In_786);
nor U858 (N_858,In_744,In_119);
or U859 (N_859,In_481,In_354);
nand U860 (N_860,In_1393,In_279);
nor U861 (N_861,In_546,In_1463);
nand U862 (N_862,In_424,In_365);
or U863 (N_863,In_731,In_326);
nor U864 (N_864,In_434,In_1226);
nor U865 (N_865,In_1251,In_436);
and U866 (N_866,In_44,In_250);
nand U867 (N_867,In_1334,In_938);
nor U868 (N_868,In_729,In_766);
nor U869 (N_869,In_1462,In_1478);
or U870 (N_870,In_1056,In_212);
or U871 (N_871,In_944,In_112);
or U872 (N_872,In_275,In_34);
or U873 (N_873,In_1352,In_1218);
or U874 (N_874,In_1216,In_462);
and U875 (N_875,In_1000,In_921);
or U876 (N_876,In_174,In_762);
or U877 (N_877,In_820,In_697);
or U878 (N_878,In_417,In_552);
nor U879 (N_879,In_1018,In_334);
or U880 (N_880,In_456,In_896);
and U881 (N_881,In_609,In_625);
nand U882 (N_882,In_1125,In_76);
nand U883 (N_883,In_727,In_1479);
nand U884 (N_884,In_494,In_701);
nor U885 (N_885,In_342,In_417);
nor U886 (N_886,In_395,In_1315);
xnor U887 (N_887,In_1343,In_699);
or U888 (N_888,In_398,In_1293);
and U889 (N_889,In_1043,In_23);
and U890 (N_890,In_197,In_1465);
and U891 (N_891,In_1293,In_778);
nand U892 (N_892,In_387,In_1304);
nor U893 (N_893,In_952,In_717);
or U894 (N_894,In_239,In_440);
and U895 (N_895,In_801,In_203);
and U896 (N_896,In_449,In_1364);
xor U897 (N_897,In_1183,In_884);
xnor U898 (N_898,In_322,In_128);
xnor U899 (N_899,In_554,In_321);
nand U900 (N_900,In_174,In_1032);
and U901 (N_901,In_0,In_276);
and U902 (N_902,In_516,In_1469);
and U903 (N_903,In_981,In_1271);
or U904 (N_904,In_753,In_481);
xnor U905 (N_905,In_16,In_732);
nor U906 (N_906,In_1151,In_920);
or U907 (N_907,In_1047,In_530);
nor U908 (N_908,In_1383,In_218);
and U909 (N_909,In_299,In_980);
or U910 (N_910,In_1268,In_902);
xor U911 (N_911,In_796,In_616);
and U912 (N_912,In_828,In_762);
or U913 (N_913,In_612,In_1187);
and U914 (N_914,In_146,In_784);
and U915 (N_915,In_610,In_1398);
nor U916 (N_916,In_1360,In_1075);
or U917 (N_917,In_77,In_1152);
nand U918 (N_918,In_1095,In_913);
or U919 (N_919,In_1350,In_881);
xor U920 (N_920,In_1156,In_1249);
or U921 (N_921,In_1228,In_548);
nor U922 (N_922,In_885,In_1490);
nor U923 (N_923,In_327,In_1209);
or U924 (N_924,In_1484,In_52);
and U925 (N_925,In_140,In_606);
or U926 (N_926,In_345,In_1126);
or U927 (N_927,In_18,In_1492);
nand U928 (N_928,In_47,In_328);
nand U929 (N_929,In_925,In_302);
and U930 (N_930,In_777,In_1067);
or U931 (N_931,In_76,In_442);
xor U932 (N_932,In_998,In_14);
xnor U933 (N_933,In_769,In_390);
or U934 (N_934,In_168,In_1405);
and U935 (N_935,In_1105,In_1140);
nand U936 (N_936,In_211,In_855);
nor U937 (N_937,In_317,In_696);
nand U938 (N_938,In_750,In_1364);
nand U939 (N_939,In_649,In_373);
nand U940 (N_940,In_151,In_1277);
and U941 (N_941,In_1216,In_428);
nor U942 (N_942,In_28,In_627);
or U943 (N_943,In_1231,In_1062);
or U944 (N_944,In_1356,In_4);
nor U945 (N_945,In_795,In_868);
and U946 (N_946,In_1299,In_1175);
and U947 (N_947,In_161,In_510);
xnor U948 (N_948,In_642,In_975);
nand U949 (N_949,In_432,In_388);
nand U950 (N_950,In_1468,In_643);
and U951 (N_951,In_714,In_352);
nand U952 (N_952,In_817,In_330);
nor U953 (N_953,In_857,In_1284);
nor U954 (N_954,In_668,In_162);
nor U955 (N_955,In_154,In_432);
nand U956 (N_956,In_1249,In_1136);
xor U957 (N_957,In_871,In_110);
and U958 (N_958,In_971,In_553);
and U959 (N_959,In_208,In_1398);
or U960 (N_960,In_1139,In_272);
nor U961 (N_961,In_1449,In_1070);
nor U962 (N_962,In_379,In_1290);
or U963 (N_963,In_215,In_1083);
or U964 (N_964,In_1340,In_825);
nand U965 (N_965,In_64,In_1095);
nand U966 (N_966,In_1394,In_133);
or U967 (N_967,In_742,In_366);
nand U968 (N_968,In_205,In_914);
nand U969 (N_969,In_1105,In_1006);
and U970 (N_970,In_1453,In_740);
nor U971 (N_971,In_1312,In_131);
and U972 (N_972,In_982,In_850);
nand U973 (N_973,In_1220,In_507);
xnor U974 (N_974,In_829,In_909);
xnor U975 (N_975,In_859,In_1088);
or U976 (N_976,In_1212,In_912);
or U977 (N_977,In_619,In_1233);
nor U978 (N_978,In_1095,In_43);
nor U979 (N_979,In_658,In_1305);
nor U980 (N_980,In_883,In_1229);
nor U981 (N_981,In_1333,In_1234);
and U982 (N_982,In_1246,In_1357);
nor U983 (N_983,In_160,In_242);
nand U984 (N_984,In_1006,In_441);
or U985 (N_985,In_1103,In_860);
and U986 (N_986,In_152,In_714);
nor U987 (N_987,In_48,In_354);
and U988 (N_988,In_403,In_839);
and U989 (N_989,In_1320,In_1422);
nand U990 (N_990,In_1196,In_666);
nand U991 (N_991,In_1386,In_409);
xnor U992 (N_992,In_1117,In_666);
or U993 (N_993,In_1162,In_1165);
nor U994 (N_994,In_724,In_9);
or U995 (N_995,In_1092,In_1166);
nand U996 (N_996,In_1364,In_189);
or U997 (N_997,In_33,In_1431);
and U998 (N_998,In_771,In_68);
or U999 (N_999,In_1210,In_181);
nor U1000 (N_1000,N_729,N_652);
nand U1001 (N_1001,N_192,N_433);
and U1002 (N_1002,N_670,N_738);
nand U1003 (N_1003,N_444,N_757);
xor U1004 (N_1004,N_285,N_100);
and U1005 (N_1005,N_804,N_482);
nand U1006 (N_1006,N_199,N_774);
and U1007 (N_1007,N_68,N_142);
and U1008 (N_1008,N_337,N_559);
and U1009 (N_1009,N_853,N_555);
or U1010 (N_1010,N_826,N_892);
nor U1011 (N_1011,N_56,N_353);
nand U1012 (N_1012,N_301,N_47);
nor U1013 (N_1013,N_924,N_576);
nand U1014 (N_1014,N_131,N_707);
nand U1015 (N_1015,N_264,N_417);
nor U1016 (N_1016,N_858,N_538);
or U1017 (N_1017,N_401,N_709);
and U1018 (N_1018,N_318,N_935);
or U1019 (N_1019,N_876,N_728);
and U1020 (N_1020,N_389,N_393);
nand U1021 (N_1021,N_244,N_21);
nor U1022 (N_1022,N_296,N_78);
and U1023 (N_1023,N_309,N_613);
or U1024 (N_1024,N_771,N_537);
or U1025 (N_1025,N_690,N_878);
and U1026 (N_1026,N_750,N_569);
nand U1027 (N_1027,N_772,N_281);
nand U1028 (N_1028,N_788,N_390);
xor U1029 (N_1029,N_66,N_907);
and U1030 (N_1030,N_777,N_455);
nor U1031 (N_1031,N_38,N_879);
nor U1032 (N_1032,N_332,N_120);
and U1033 (N_1033,N_122,N_730);
nand U1034 (N_1034,N_67,N_64);
nand U1035 (N_1035,N_282,N_779);
nand U1036 (N_1036,N_500,N_840);
and U1037 (N_1037,N_564,N_351);
nand U1038 (N_1038,N_240,N_780);
xor U1039 (N_1039,N_813,N_571);
and U1040 (N_1040,N_151,N_894);
nand U1041 (N_1041,N_355,N_827);
and U1042 (N_1042,N_74,N_228);
or U1043 (N_1043,N_653,N_620);
or U1044 (N_1044,N_783,N_803);
xnor U1045 (N_1045,N_300,N_499);
nand U1046 (N_1046,N_60,N_243);
and U1047 (N_1047,N_502,N_460);
or U1048 (N_1048,N_823,N_609);
xnor U1049 (N_1049,N_394,N_81);
xnor U1050 (N_1050,N_964,N_617);
nor U1051 (N_1051,N_7,N_668);
or U1052 (N_1052,N_648,N_548);
nand U1053 (N_1053,N_48,N_104);
nor U1054 (N_1054,N_345,N_687);
and U1055 (N_1055,N_540,N_268);
nand U1056 (N_1056,N_622,N_927);
nand U1057 (N_1057,N_226,N_970);
and U1058 (N_1058,N_890,N_114);
and U1059 (N_1059,N_657,N_820);
and U1060 (N_1060,N_658,N_517);
nand U1061 (N_1061,N_539,N_515);
nor U1062 (N_1062,N_125,N_546);
nor U1063 (N_1063,N_516,N_407);
and U1064 (N_1064,N_751,N_856);
xor U1065 (N_1065,N_615,N_526);
xor U1066 (N_1066,N_725,N_118);
nor U1067 (N_1067,N_427,N_972);
nand U1068 (N_1068,N_486,N_986);
or U1069 (N_1069,N_391,N_824);
or U1070 (N_1070,N_875,N_440);
nor U1071 (N_1071,N_900,N_676);
and U1072 (N_1072,N_736,N_694);
or U1073 (N_1073,N_134,N_380);
or U1074 (N_1074,N_156,N_714);
nor U1075 (N_1075,N_520,N_959);
nand U1076 (N_1076,N_895,N_831);
and U1077 (N_1077,N_600,N_587);
nand U1078 (N_1078,N_320,N_912);
or U1079 (N_1079,N_713,N_65);
or U1080 (N_1080,N_329,N_14);
nor U1081 (N_1081,N_53,N_932);
nor U1082 (N_1082,N_397,N_145);
nand U1083 (N_1083,N_975,N_384);
nor U1084 (N_1084,N_280,N_457);
and U1085 (N_1085,N_375,N_225);
nand U1086 (N_1086,N_553,N_825);
or U1087 (N_1087,N_365,N_160);
and U1088 (N_1088,N_313,N_193);
and U1089 (N_1089,N_669,N_230);
nor U1090 (N_1090,N_469,N_834);
nand U1091 (N_1091,N_987,N_643);
or U1092 (N_1092,N_425,N_437);
nor U1093 (N_1093,N_719,N_662);
or U1094 (N_1094,N_592,N_4);
and U1095 (N_1095,N_426,N_636);
and U1096 (N_1096,N_378,N_819);
and U1097 (N_1097,N_37,N_184);
and U1098 (N_1098,N_445,N_299);
or U1099 (N_1099,N_284,N_712);
nor U1100 (N_1100,N_412,N_494);
nand U1101 (N_1101,N_861,N_950);
and U1102 (N_1102,N_654,N_42);
and U1103 (N_1103,N_256,N_162);
or U1104 (N_1104,N_626,N_930);
nand U1105 (N_1105,N_829,N_101);
nand U1106 (N_1106,N_556,N_787);
xor U1107 (N_1107,N_852,N_597);
xor U1108 (N_1108,N_245,N_881);
and U1109 (N_1109,N_436,N_305);
or U1110 (N_1110,N_689,N_155);
and U1111 (N_1111,N_635,N_321);
nand U1112 (N_1112,N_168,N_58);
nand U1113 (N_1113,N_767,N_232);
and U1114 (N_1114,N_582,N_854);
nor U1115 (N_1115,N_490,N_73);
nand U1116 (N_1116,N_599,N_405);
or U1117 (N_1117,N_784,N_504);
and U1118 (N_1118,N_498,N_439);
or U1119 (N_1119,N_262,N_420);
nor U1120 (N_1120,N_949,N_186);
and U1121 (N_1121,N_678,N_450);
xor U1122 (N_1122,N_641,N_188);
nor U1123 (N_1123,N_550,N_395);
nand U1124 (N_1124,N_428,N_346);
nand U1125 (N_1125,N_373,N_998);
xor U1126 (N_1126,N_89,N_695);
nand U1127 (N_1127,N_740,N_19);
nor U1128 (N_1128,N_344,N_148);
nand U1129 (N_1129,N_107,N_413);
nor U1130 (N_1130,N_290,N_586);
or U1131 (N_1131,N_717,N_419);
nor U1132 (N_1132,N_61,N_704);
nor U1133 (N_1133,N_83,N_170);
nor U1134 (N_1134,N_567,N_942);
nor U1135 (N_1135,N_24,N_115);
xor U1136 (N_1136,N_288,N_706);
or U1137 (N_1137,N_454,N_589);
xor U1138 (N_1138,N_34,N_6);
and U1139 (N_1139,N_802,N_492);
and U1140 (N_1140,N_319,N_533);
xnor U1141 (N_1141,N_833,N_529);
nand U1142 (N_1142,N_431,N_625);
nor U1143 (N_1143,N_381,N_743);
or U1144 (N_1144,N_388,N_234);
and U1145 (N_1145,N_404,N_235);
and U1146 (N_1146,N_86,N_449);
xnor U1147 (N_1147,N_606,N_448);
xnor U1148 (N_1148,N_124,N_638);
or U1149 (N_1149,N_896,N_446);
xnor U1150 (N_1150,N_370,N_680);
nor U1151 (N_1151,N_749,N_790);
nor U1152 (N_1152,N_985,N_647);
nor U1153 (N_1153,N_205,N_874);
and U1154 (N_1154,N_286,N_8);
nor U1155 (N_1155,N_175,N_254);
nand U1156 (N_1156,N_399,N_700);
nand U1157 (N_1157,N_350,N_863);
nor U1158 (N_1158,N_877,N_276);
and U1159 (N_1159,N_266,N_493);
nand U1160 (N_1160,N_948,N_623);
nor U1161 (N_1161,N_882,N_503);
nor U1162 (N_1162,N_289,N_443);
nor U1163 (N_1163,N_32,N_521);
and U1164 (N_1164,N_675,N_781);
xnor U1165 (N_1165,N_776,N_541);
and U1166 (N_1166,N_846,N_222);
or U1167 (N_1167,N_651,N_965);
or U1168 (N_1168,N_485,N_45);
nor U1169 (N_1169,N_112,N_333);
or U1170 (N_1170,N_684,N_631);
xor U1171 (N_1171,N_75,N_176);
nor U1172 (N_1172,N_765,N_307);
nand U1173 (N_1173,N_462,N_737);
and U1174 (N_1174,N_123,N_614);
and U1175 (N_1175,N_483,N_797);
nand U1176 (N_1176,N_259,N_260);
xnor U1177 (N_1177,N_174,N_545);
and U1178 (N_1178,N_809,N_110);
and U1179 (N_1179,N_465,N_630);
or U1180 (N_1180,N_593,N_136);
and U1181 (N_1181,N_721,N_655);
nand U1182 (N_1182,N_835,N_855);
and U1183 (N_1183,N_837,N_656);
and U1184 (N_1184,N_920,N_28);
or U1185 (N_1185,N_430,N_796);
nand U1186 (N_1186,N_435,N_202);
and U1187 (N_1187,N_361,N_688);
or U1188 (N_1188,N_509,N_880);
or U1189 (N_1189,N_768,N_293);
nand U1190 (N_1190,N_302,N_782);
or U1191 (N_1191,N_869,N_308);
and U1192 (N_1192,N_158,N_660);
and U1193 (N_1193,N_88,N_514);
and U1194 (N_1194,N_720,N_996);
and U1195 (N_1195,N_505,N_672);
xor U1196 (N_1196,N_785,N_421);
nor U1197 (N_1197,N_255,N_627);
and U1198 (N_1198,N_328,N_872);
and U1199 (N_1199,N_558,N_868);
and U1200 (N_1200,N_1,N_974);
nand U1201 (N_1201,N_792,N_769);
or U1202 (N_1202,N_166,N_645);
xnor U1203 (N_1203,N_758,N_10);
and U1204 (N_1204,N_943,N_921);
or U1205 (N_1205,N_273,N_691);
and U1206 (N_1206,N_130,N_566);
nor U1207 (N_1207,N_29,N_117);
nand U1208 (N_1208,N_929,N_325);
xor U1209 (N_1209,N_632,N_696);
and U1210 (N_1210,N_178,N_54);
xnor U1211 (N_1211,N_96,N_291);
nand U1212 (N_1212,N_206,N_637);
nor U1213 (N_1213,N_251,N_955);
xor U1214 (N_1214,N_715,N_610);
nor U1215 (N_1215,N_572,N_212);
nand U1216 (N_1216,N_62,N_468);
nand U1217 (N_1217,N_966,N_800);
and U1218 (N_1218,N_588,N_640);
and U1219 (N_1219,N_993,N_973);
nor U1220 (N_1220,N_575,N_204);
and U1221 (N_1221,N_451,N_761);
nor U1222 (N_1222,N_795,N_140);
nor U1223 (N_1223,N_474,N_899);
and U1224 (N_1224,N_480,N_180);
or U1225 (N_1225,N_363,N_698);
and U1226 (N_1226,N_360,N_798);
or U1227 (N_1227,N_43,N_507);
nand U1228 (N_1228,N_536,N_411);
and U1229 (N_1229,N_988,N_999);
nor U1230 (N_1230,N_961,N_9);
nor U1231 (N_1231,N_138,N_778);
nor U1232 (N_1232,N_956,N_983);
or U1233 (N_1233,N_770,N_317);
nand U1234 (N_1234,N_946,N_732);
and U1235 (N_1235,N_137,N_11);
nand U1236 (N_1236,N_182,N_897);
nand U1237 (N_1237,N_547,N_242);
nor U1238 (N_1238,N_159,N_551);
and U1239 (N_1239,N_119,N_349);
nor U1240 (N_1240,N_164,N_338);
xor U1241 (N_1241,N_258,N_153);
or U1242 (N_1242,N_22,N_116);
and U1243 (N_1243,N_969,N_705);
and U1244 (N_1244,N_673,N_368);
nand U1245 (N_1245,N_362,N_710);
nor U1246 (N_1246,N_267,N_383);
and U1247 (N_1247,N_685,N_13);
or U1248 (N_1248,N_82,N_938);
or U1249 (N_1249,N_914,N_544);
nor U1250 (N_1250,N_220,N_44);
nor U1251 (N_1251,N_377,N_607);
nand U1252 (N_1252,N_697,N_463);
nor U1253 (N_1253,N_594,N_239);
or U1254 (N_1254,N_584,N_667);
or U1255 (N_1255,N_940,N_98);
and U1256 (N_1256,N_141,N_99);
nor U1257 (N_1257,N_39,N_724);
nor U1258 (N_1258,N_917,N_198);
or U1259 (N_1259,N_731,N_557);
nor U1260 (N_1260,N_165,N_901);
nor U1261 (N_1261,N_671,N_708);
or U1262 (N_1262,N_379,N_808);
or U1263 (N_1263,N_931,N_133);
xor U1264 (N_1264,N_441,N_570);
xor U1265 (N_1265,N_811,N_311);
nand U1266 (N_1266,N_560,N_801);
or U1267 (N_1267,N_315,N_423);
nor U1268 (N_1268,N_911,N_272);
nor U1269 (N_1269,N_686,N_756);
or U1270 (N_1270,N_518,N_2);
and U1271 (N_1271,N_354,N_200);
and U1272 (N_1272,N_250,N_995);
nand U1273 (N_1273,N_523,N_257);
and U1274 (N_1274,N_214,N_794);
or U1275 (N_1275,N_722,N_295);
or U1276 (N_1276,N_866,N_902);
or U1277 (N_1277,N_663,N_976);
or U1278 (N_1278,N_665,N_984);
or U1279 (N_1279,N_147,N_734);
nand U1280 (N_1280,N_945,N_554);
nor U1281 (N_1281,N_522,N_69);
nor U1282 (N_1282,N_885,N_893);
nand U1283 (N_1283,N_314,N_292);
nor U1284 (N_1284,N_487,N_579);
nand U1285 (N_1285,N_102,N_922);
nor U1286 (N_1286,N_848,N_113);
xor U1287 (N_1287,N_603,N_598);
and U1288 (N_1288,N_20,N_424);
nand U1289 (N_1289,N_699,N_386);
or U1290 (N_1290,N_126,N_236);
nand U1291 (N_1291,N_532,N_919);
nor U1292 (N_1292,N_471,N_408);
xor U1293 (N_1293,N_591,N_601);
and U1294 (N_1294,N_674,N_310);
and U1295 (N_1295,N_447,N_464);
nand U1296 (N_1296,N_549,N_847);
or U1297 (N_1297,N_477,N_838);
and U1298 (N_1298,N_644,N_530);
xnor U1299 (N_1299,N_211,N_832);
nand U1300 (N_1300,N_596,N_191);
nor U1301 (N_1301,N_619,N_903);
and U1302 (N_1302,N_479,N_94);
or U1303 (N_1303,N_957,N_331);
xnor U1304 (N_1304,N_303,N_163);
nor U1305 (N_1305,N_595,N_789);
xor U1306 (N_1306,N_461,N_79);
xor U1307 (N_1307,N_238,N_371);
nor U1308 (N_1308,N_527,N_229);
nand U1309 (N_1309,N_342,N_71);
or U1310 (N_1310,N_585,N_746);
or U1311 (N_1311,N_343,N_452);
xnor U1312 (N_1312,N_372,N_519);
nand U1313 (N_1313,N_602,N_481);
nor U1314 (N_1314,N_128,N_865);
or U1315 (N_1315,N_227,N_843);
or U1316 (N_1316,N_535,N_563);
xnor U1317 (N_1317,N_666,N_573);
nor U1318 (N_1318,N_958,N_991);
nand U1319 (N_1319,N_279,N_543);
and U1320 (N_1320,N_358,N_745);
or U1321 (N_1321,N_52,N_941);
nor U1322 (N_1322,N_219,N_859);
nand U1323 (N_1323,N_978,N_703);
nor U1324 (N_1324,N_822,N_97);
nor U1325 (N_1325,N_422,N_839);
and U1326 (N_1326,N_992,N_936);
or U1327 (N_1327,N_135,N_891);
nand U1328 (N_1328,N_628,N_764);
nand U1329 (N_1329,N_248,N_981);
nor U1330 (N_1330,N_616,N_348);
xor U1331 (N_1331,N_979,N_618);
or U1332 (N_1332,N_341,N_77);
nor U1333 (N_1333,N_997,N_106);
or U1334 (N_1334,N_265,N_581);
or U1335 (N_1335,N_842,N_762);
or U1336 (N_1336,N_85,N_287);
nor U1337 (N_1337,N_884,N_187);
and U1338 (N_1338,N_962,N_467);
and U1339 (N_1339,N_817,N_35);
or U1340 (N_1340,N_629,N_217);
or U1341 (N_1341,N_400,N_830);
and U1342 (N_1342,N_791,N_409);
or U1343 (N_1343,N_76,N_814);
or U1344 (N_1344,N_806,N_864);
or U1345 (N_1345,N_194,N_501);
nor U1346 (N_1346,N_171,N_197);
or U1347 (N_1347,N_752,N_369);
nand U1348 (N_1348,N_634,N_429);
nand U1349 (N_1349,N_590,N_488);
and U1350 (N_1350,N_508,N_951);
nand U1351 (N_1351,N_913,N_818);
nand U1352 (N_1352,N_72,N_473);
or U1353 (N_1353,N_111,N_415);
nand U1354 (N_1354,N_18,N_298);
nor U1355 (N_1355,N_860,N_108);
or U1356 (N_1356,N_366,N_249);
nor U1357 (N_1357,N_718,N_271);
nor U1358 (N_1358,N_132,N_867);
nor U1359 (N_1359,N_915,N_442);
xnor U1360 (N_1360,N_763,N_524);
nor U1361 (N_1361,N_661,N_513);
or U1362 (N_1362,N_149,N_172);
nand U1363 (N_1363,N_968,N_624);
nand U1364 (N_1364,N_453,N_203);
and U1365 (N_1365,N_971,N_744);
nand U1366 (N_1366,N_491,N_711);
or U1367 (N_1367,N_27,N_977);
or U1368 (N_1368,N_210,N_177);
or U1369 (N_1369,N_387,N_816);
or U1370 (N_1370,N_646,N_916);
nor U1371 (N_1371,N_306,N_621);
nand U1372 (N_1372,N_799,N_857);
and U1373 (N_1373,N_608,N_475);
xor U1374 (N_1374,N_679,N_91);
or U1375 (N_1375,N_432,N_456);
xnor U1376 (N_1376,N_270,N_46);
or U1377 (N_1377,N_12,N_190);
and U1378 (N_1378,N_506,N_726);
nor U1379 (N_1379,N_478,N_278);
nor U1380 (N_1380,N_15,N_980);
and U1381 (N_1381,N_723,N_953);
or U1382 (N_1382,N_334,N_41);
nand U1383 (N_1383,N_497,N_905);
or U1384 (N_1384,N_990,N_870);
and U1385 (N_1385,N_611,N_173);
nand U1386 (N_1386,N_146,N_129);
nor U1387 (N_1387,N_36,N_735);
xor U1388 (N_1388,N_871,N_406);
or U1389 (N_1389,N_476,N_807);
nor U1390 (N_1390,N_80,N_759);
nand U1391 (N_1391,N_0,N_416);
or U1392 (N_1392,N_574,N_484);
or U1393 (N_1393,N_207,N_283);
xor U1394 (N_1394,N_753,N_873);
nand U1395 (N_1395,N_189,N_90);
nor U1396 (N_1396,N_364,N_495);
and U1397 (N_1397,N_459,N_909);
or U1398 (N_1398,N_755,N_747);
nand U1399 (N_1399,N_324,N_323);
nor U1400 (N_1400,N_340,N_470);
nand U1401 (N_1401,N_862,N_376);
or U1402 (N_1402,N_326,N_583);
nand U1403 (N_1403,N_327,N_367);
nand U1404 (N_1404,N_139,N_167);
xor U1405 (N_1405,N_396,N_604);
nand U1406 (N_1406,N_51,N_954);
nand U1407 (N_1407,N_741,N_944);
xnor U1408 (N_1408,N_196,N_294);
nand U1409 (N_1409,N_231,N_928);
nor U1410 (N_1410,N_26,N_568);
nor U1411 (N_1411,N_70,N_677);
nor U1412 (N_1412,N_359,N_923);
or U1413 (N_1413,N_682,N_253);
nand U1414 (N_1414,N_466,N_561);
and U1415 (N_1415,N_414,N_25);
or U1416 (N_1416,N_33,N_93);
or U1417 (N_1417,N_664,N_103);
and U1418 (N_1418,N_312,N_5);
and U1419 (N_1419,N_815,N_181);
nand U1420 (N_1420,N_639,N_926);
nor U1421 (N_1421,N_92,N_304);
nand U1422 (N_1422,N_150,N_952);
or U1423 (N_1423,N_269,N_908);
or U1424 (N_1424,N_947,N_385);
and U1425 (N_1425,N_316,N_716);
nor U1426 (N_1426,N_934,N_49);
nand U1427 (N_1427,N_16,N_392);
and U1428 (N_1428,N_336,N_775);
nor U1429 (N_1429,N_213,N_143);
xor U1430 (N_1430,N_418,N_733);
nand U1431 (N_1431,N_510,N_221);
or U1432 (N_1432,N_208,N_261);
nor U1433 (N_1433,N_215,N_933);
or U1434 (N_1434,N_805,N_374);
or U1435 (N_1435,N_152,N_458);
xnor U1436 (N_1436,N_322,N_169);
xnor U1437 (N_1437,N_434,N_201);
nor U1438 (N_1438,N_531,N_223);
nand U1439 (N_1439,N_512,N_109);
and U1440 (N_1440,N_773,N_216);
xnor U1441 (N_1441,N_55,N_95);
and U1442 (N_1442,N_154,N_402);
and U1443 (N_1443,N_127,N_793);
or U1444 (N_1444,N_766,N_844);
nand U1445 (N_1445,N_489,N_23);
nor U1446 (N_1446,N_339,N_889);
nand U1447 (N_1447,N_252,N_963);
xnor U1448 (N_1448,N_812,N_496);
nor U1449 (N_1449,N_534,N_382);
or U1450 (N_1450,N_275,N_17);
and U1451 (N_1451,N_939,N_605);
and U1452 (N_1452,N_195,N_681);
nor U1453 (N_1453,N_994,N_982);
nor U1454 (N_1454,N_850,N_565);
or U1455 (N_1455,N_330,N_562);
nor U1456 (N_1456,N_828,N_233);
or U1457 (N_1457,N_580,N_179);
xor U1458 (N_1458,N_528,N_335);
nor U1459 (N_1459,N_209,N_786);
nand U1460 (N_1460,N_224,N_851);
nand U1461 (N_1461,N_760,N_633);
and U1462 (N_1462,N_748,N_183);
xnor U1463 (N_1463,N_356,N_84);
nand U1464 (N_1464,N_525,N_904);
nor U1465 (N_1465,N_821,N_925);
nor U1466 (N_1466,N_841,N_237);
or U1467 (N_1467,N_87,N_277);
or U1468 (N_1468,N_121,N_403);
or U1469 (N_1469,N_247,N_888);
nand U1470 (N_1470,N_577,N_692);
nor U1471 (N_1471,N_63,N_883);
or U1472 (N_1472,N_910,N_650);
and U1473 (N_1473,N_739,N_727);
xnor U1474 (N_1474,N_810,N_472);
or U1475 (N_1475,N_246,N_887);
nand U1476 (N_1476,N_989,N_31);
nand U1477 (N_1477,N_683,N_157);
or U1478 (N_1478,N_578,N_357);
and U1479 (N_1479,N_886,N_410);
nand U1480 (N_1480,N_754,N_161);
xor U1481 (N_1481,N_659,N_347);
or U1482 (N_1482,N_274,N_960);
nor U1483 (N_1483,N_612,N_967);
nand U1484 (N_1484,N_241,N_693);
xnor U1485 (N_1485,N_40,N_742);
nor U1486 (N_1486,N_144,N_845);
and U1487 (N_1487,N_918,N_30);
nand U1488 (N_1488,N_702,N_263);
and U1489 (N_1489,N_105,N_185);
or U1490 (N_1490,N_849,N_649);
nor U1491 (N_1491,N_906,N_50);
nor U1492 (N_1492,N_59,N_297);
xor U1493 (N_1493,N_398,N_898);
or U1494 (N_1494,N_642,N_701);
or U1495 (N_1495,N_438,N_352);
nor U1496 (N_1496,N_511,N_937);
nor U1497 (N_1497,N_57,N_3);
xor U1498 (N_1498,N_836,N_218);
nand U1499 (N_1499,N_552,N_542);
and U1500 (N_1500,N_971,N_916);
nor U1501 (N_1501,N_201,N_321);
nor U1502 (N_1502,N_257,N_772);
and U1503 (N_1503,N_268,N_770);
nand U1504 (N_1504,N_654,N_161);
or U1505 (N_1505,N_702,N_126);
nand U1506 (N_1506,N_921,N_591);
or U1507 (N_1507,N_214,N_944);
and U1508 (N_1508,N_304,N_695);
nand U1509 (N_1509,N_130,N_516);
nor U1510 (N_1510,N_471,N_29);
and U1511 (N_1511,N_249,N_488);
nor U1512 (N_1512,N_835,N_201);
and U1513 (N_1513,N_345,N_561);
or U1514 (N_1514,N_681,N_483);
nor U1515 (N_1515,N_989,N_356);
or U1516 (N_1516,N_806,N_303);
and U1517 (N_1517,N_918,N_81);
or U1518 (N_1518,N_309,N_494);
nor U1519 (N_1519,N_828,N_359);
or U1520 (N_1520,N_4,N_777);
or U1521 (N_1521,N_581,N_714);
or U1522 (N_1522,N_419,N_156);
nor U1523 (N_1523,N_917,N_837);
nor U1524 (N_1524,N_207,N_808);
or U1525 (N_1525,N_310,N_374);
and U1526 (N_1526,N_866,N_69);
nor U1527 (N_1527,N_502,N_936);
nor U1528 (N_1528,N_470,N_192);
nand U1529 (N_1529,N_588,N_131);
nor U1530 (N_1530,N_267,N_740);
or U1531 (N_1531,N_199,N_390);
nor U1532 (N_1532,N_558,N_150);
and U1533 (N_1533,N_924,N_920);
xnor U1534 (N_1534,N_943,N_475);
xor U1535 (N_1535,N_93,N_567);
and U1536 (N_1536,N_77,N_12);
nand U1537 (N_1537,N_632,N_43);
nor U1538 (N_1538,N_589,N_314);
xnor U1539 (N_1539,N_71,N_720);
nand U1540 (N_1540,N_138,N_204);
nand U1541 (N_1541,N_288,N_129);
xnor U1542 (N_1542,N_16,N_203);
nor U1543 (N_1543,N_175,N_986);
nor U1544 (N_1544,N_304,N_759);
or U1545 (N_1545,N_589,N_662);
and U1546 (N_1546,N_846,N_842);
nand U1547 (N_1547,N_851,N_431);
nor U1548 (N_1548,N_918,N_520);
and U1549 (N_1549,N_410,N_181);
and U1550 (N_1550,N_402,N_996);
nand U1551 (N_1551,N_771,N_11);
xnor U1552 (N_1552,N_528,N_244);
and U1553 (N_1553,N_332,N_790);
xor U1554 (N_1554,N_802,N_386);
nor U1555 (N_1555,N_494,N_846);
nand U1556 (N_1556,N_346,N_30);
nor U1557 (N_1557,N_856,N_696);
nor U1558 (N_1558,N_174,N_600);
nor U1559 (N_1559,N_746,N_402);
nand U1560 (N_1560,N_970,N_216);
nor U1561 (N_1561,N_506,N_497);
or U1562 (N_1562,N_25,N_835);
or U1563 (N_1563,N_843,N_325);
xnor U1564 (N_1564,N_540,N_445);
nand U1565 (N_1565,N_373,N_891);
or U1566 (N_1566,N_859,N_231);
xnor U1567 (N_1567,N_224,N_985);
nor U1568 (N_1568,N_681,N_695);
or U1569 (N_1569,N_306,N_648);
or U1570 (N_1570,N_180,N_307);
nor U1571 (N_1571,N_873,N_929);
and U1572 (N_1572,N_734,N_813);
nor U1573 (N_1573,N_772,N_605);
nor U1574 (N_1574,N_135,N_675);
nor U1575 (N_1575,N_725,N_349);
nand U1576 (N_1576,N_573,N_892);
nand U1577 (N_1577,N_120,N_794);
and U1578 (N_1578,N_189,N_478);
nor U1579 (N_1579,N_655,N_489);
nor U1580 (N_1580,N_38,N_445);
nand U1581 (N_1581,N_27,N_579);
nor U1582 (N_1582,N_728,N_622);
xnor U1583 (N_1583,N_564,N_49);
nor U1584 (N_1584,N_105,N_221);
or U1585 (N_1585,N_125,N_235);
nor U1586 (N_1586,N_539,N_357);
nor U1587 (N_1587,N_703,N_395);
or U1588 (N_1588,N_783,N_425);
xor U1589 (N_1589,N_706,N_875);
nor U1590 (N_1590,N_310,N_50);
and U1591 (N_1591,N_831,N_515);
and U1592 (N_1592,N_581,N_189);
or U1593 (N_1593,N_457,N_173);
xor U1594 (N_1594,N_373,N_387);
and U1595 (N_1595,N_884,N_258);
nor U1596 (N_1596,N_647,N_63);
nand U1597 (N_1597,N_268,N_44);
xor U1598 (N_1598,N_584,N_386);
or U1599 (N_1599,N_726,N_72);
nand U1600 (N_1600,N_789,N_573);
nand U1601 (N_1601,N_46,N_42);
nand U1602 (N_1602,N_486,N_796);
and U1603 (N_1603,N_322,N_10);
nor U1604 (N_1604,N_45,N_326);
nor U1605 (N_1605,N_705,N_588);
nor U1606 (N_1606,N_995,N_62);
nor U1607 (N_1607,N_564,N_247);
nand U1608 (N_1608,N_937,N_660);
nand U1609 (N_1609,N_181,N_776);
nor U1610 (N_1610,N_669,N_362);
nor U1611 (N_1611,N_286,N_417);
xnor U1612 (N_1612,N_921,N_972);
nand U1613 (N_1613,N_301,N_525);
nand U1614 (N_1614,N_606,N_993);
nand U1615 (N_1615,N_936,N_525);
or U1616 (N_1616,N_271,N_894);
nor U1617 (N_1617,N_390,N_329);
nor U1618 (N_1618,N_16,N_119);
nand U1619 (N_1619,N_953,N_405);
nand U1620 (N_1620,N_6,N_744);
nor U1621 (N_1621,N_5,N_359);
nor U1622 (N_1622,N_488,N_5);
nand U1623 (N_1623,N_518,N_558);
nand U1624 (N_1624,N_30,N_107);
nor U1625 (N_1625,N_30,N_188);
nand U1626 (N_1626,N_334,N_840);
nor U1627 (N_1627,N_716,N_836);
or U1628 (N_1628,N_566,N_757);
nand U1629 (N_1629,N_42,N_363);
nor U1630 (N_1630,N_264,N_225);
and U1631 (N_1631,N_647,N_642);
nand U1632 (N_1632,N_660,N_103);
or U1633 (N_1633,N_831,N_858);
nor U1634 (N_1634,N_774,N_235);
and U1635 (N_1635,N_505,N_309);
nor U1636 (N_1636,N_648,N_595);
nor U1637 (N_1637,N_150,N_498);
and U1638 (N_1638,N_65,N_825);
nor U1639 (N_1639,N_150,N_973);
and U1640 (N_1640,N_242,N_497);
nand U1641 (N_1641,N_641,N_265);
or U1642 (N_1642,N_935,N_323);
nor U1643 (N_1643,N_567,N_24);
or U1644 (N_1644,N_73,N_683);
and U1645 (N_1645,N_403,N_883);
or U1646 (N_1646,N_764,N_153);
nand U1647 (N_1647,N_721,N_601);
nor U1648 (N_1648,N_361,N_655);
and U1649 (N_1649,N_9,N_650);
nor U1650 (N_1650,N_248,N_917);
and U1651 (N_1651,N_764,N_480);
and U1652 (N_1652,N_815,N_751);
or U1653 (N_1653,N_572,N_529);
nor U1654 (N_1654,N_931,N_535);
or U1655 (N_1655,N_557,N_407);
nand U1656 (N_1656,N_911,N_180);
xor U1657 (N_1657,N_997,N_421);
nand U1658 (N_1658,N_873,N_973);
nand U1659 (N_1659,N_755,N_881);
nor U1660 (N_1660,N_885,N_634);
nand U1661 (N_1661,N_266,N_21);
and U1662 (N_1662,N_414,N_352);
or U1663 (N_1663,N_941,N_903);
xor U1664 (N_1664,N_859,N_488);
and U1665 (N_1665,N_656,N_421);
and U1666 (N_1666,N_709,N_167);
nor U1667 (N_1667,N_705,N_80);
or U1668 (N_1668,N_167,N_344);
nor U1669 (N_1669,N_700,N_752);
or U1670 (N_1670,N_73,N_328);
and U1671 (N_1671,N_654,N_254);
xor U1672 (N_1672,N_570,N_579);
and U1673 (N_1673,N_587,N_243);
and U1674 (N_1674,N_563,N_140);
nor U1675 (N_1675,N_125,N_113);
nand U1676 (N_1676,N_560,N_58);
nand U1677 (N_1677,N_18,N_436);
and U1678 (N_1678,N_138,N_433);
and U1679 (N_1679,N_509,N_735);
or U1680 (N_1680,N_337,N_953);
nand U1681 (N_1681,N_742,N_388);
or U1682 (N_1682,N_315,N_586);
or U1683 (N_1683,N_182,N_719);
nand U1684 (N_1684,N_222,N_680);
nor U1685 (N_1685,N_337,N_393);
xor U1686 (N_1686,N_739,N_561);
xnor U1687 (N_1687,N_208,N_677);
xnor U1688 (N_1688,N_278,N_894);
nand U1689 (N_1689,N_128,N_607);
nor U1690 (N_1690,N_636,N_563);
xor U1691 (N_1691,N_336,N_995);
nor U1692 (N_1692,N_815,N_386);
and U1693 (N_1693,N_210,N_951);
or U1694 (N_1694,N_551,N_283);
and U1695 (N_1695,N_571,N_206);
nor U1696 (N_1696,N_166,N_997);
and U1697 (N_1697,N_989,N_743);
or U1698 (N_1698,N_423,N_777);
xor U1699 (N_1699,N_390,N_985);
nor U1700 (N_1700,N_658,N_972);
and U1701 (N_1701,N_214,N_551);
nor U1702 (N_1702,N_537,N_146);
and U1703 (N_1703,N_375,N_508);
and U1704 (N_1704,N_488,N_897);
and U1705 (N_1705,N_447,N_52);
nand U1706 (N_1706,N_816,N_900);
or U1707 (N_1707,N_119,N_330);
and U1708 (N_1708,N_951,N_54);
and U1709 (N_1709,N_96,N_311);
nand U1710 (N_1710,N_825,N_915);
or U1711 (N_1711,N_736,N_592);
nand U1712 (N_1712,N_822,N_369);
and U1713 (N_1713,N_447,N_497);
nor U1714 (N_1714,N_348,N_907);
nor U1715 (N_1715,N_729,N_413);
or U1716 (N_1716,N_197,N_783);
and U1717 (N_1717,N_645,N_473);
or U1718 (N_1718,N_601,N_84);
or U1719 (N_1719,N_499,N_478);
and U1720 (N_1720,N_861,N_773);
nand U1721 (N_1721,N_821,N_723);
nand U1722 (N_1722,N_669,N_65);
and U1723 (N_1723,N_194,N_206);
and U1724 (N_1724,N_983,N_481);
nor U1725 (N_1725,N_758,N_363);
nand U1726 (N_1726,N_482,N_795);
nor U1727 (N_1727,N_75,N_634);
and U1728 (N_1728,N_563,N_513);
and U1729 (N_1729,N_178,N_619);
nand U1730 (N_1730,N_993,N_336);
and U1731 (N_1731,N_929,N_494);
xor U1732 (N_1732,N_478,N_927);
xor U1733 (N_1733,N_382,N_523);
nor U1734 (N_1734,N_603,N_887);
and U1735 (N_1735,N_753,N_152);
nor U1736 (N_1736,N_191,N_998);
xor U1737 (N_1737,N_176,N_960);
and U1738 (N_1738,N_62,N_431);
nor U1739 (N_1739,N_144,N_234);
and U1740 (N_1740,N_851,N_286);
and U1741 (N_1741,N_681,N_329);
nor U1742 (N_1742,N_442,N_516);
or U1743 (N_1743,N_821,N_835);
or U1744 (N_1744,N_814,N_630);
or U1745 (N_1745,N_123,N_159);
and U1746 (N_1746,N_797,N_501);
or U1747 (N_1747,N_141,N_270);
and U1748 (N_1748,N_263,N_46);
nor U1749 (N_1749,N_100,N_184);
or U1750 (N_1750,N_136,N_985);
or U1751 (N_1751,N_70,N_793);
nand U1752 (N_1752,N_738,N_293);
and U1753 (N_1753,N_732,N_710);
nand U1754 (N_1754,N_311,N_681);
and U1755 (N_1755,N_936,N_926);
or U1756 (N_1756,N_649,N_685);
xnor U1757 (N_1757,N_793,N_618);
or U1758 (N_1758,N_720,N_93);
and U1759 (N_1759,N_868,N_975);
and U1760 (N_1760,N_443,N_144);
xor U1761 (N_1761,N_583,N_956);
nand U1762 (N_1762,N_235,N_421);
or U1763 (N_1763,N_825,N_393);
and U1764 (N_1764,N_329,N_74);
and U1765 (N_1765,N_413,N_357);
nor U1766 (N_1766,N_741,N_866);
nor U1767 (N_1767,N_563,N_670);
or U1768 (N_1768,N_17,N_189);
nand U1769 (N_1769,N_831,N_990);
nand U1770 (N_1770,N_487,N_377);
xnor U1771 (N_1771,N_68,N_21);
nor U1772 (N_1772,N_61,N_883);
and U1773 (N_1773,N_871,N_467);
and U1774 (N_1774,N_73,N_304);
or U1775 (N_1775,N_586,N_630);
nor U1776 (N_1776,N_420,N_220);
nor U1777 (N_1777,N_932,N_776);
nor U1778 (N_1778,N_221,N_773);
nor U1779 (N_1779,N_445,N_229);
or U1780 (N_1780,N_307,N_336);
nor U1781 (N_1781,N_701,N_480);
or U1782 (N_1782,N_228,N_622);
nor U1783 (N_1783,N_527,N_100);
or U1784 (N_1784,N_170,N_169);
nor U1785 (N_1785,N_753,N_288);
xnor U1786 (N_1786,N_702,N_955);
and U1787 (N_1787,N_702,N_768);
nand U1788 (N_1788,N_515,N_47);
nand U1789 (N_1789,N_809,N_586);
and U1790 (N_1790,N_525,N_456);
or U1791 (N_1791,N_891,N_66);
nand U1792 (N_1792,N_820,N_765);
nor U1793 (N_1793,N_376,N_386);
or U1794 (N_1794,N_92,N_983);
xnor U1795 (N_1795,N_53,N_424);
nor U1796 (N_1796,N_409,N_526);
and U1797 (N_1797,N_685,N_616);
and U1798 (N_1798,N_89,N_314);
xor U1799 (N_1799,N_9,N_512);
nor U1800 (N_1800,N_485,N_227);
or U1801 (N_1801,N_357,N_208);
nand U1802 (N_1802,N_177,N_199);
nor U1803 (N_1803,N_198,N_331);
and U1804 (N_1804,N_956,N_91);
or U1805 (N_1805,N_0,N_312);
nand U1806 (N_1806,N_472,N_980);
nor U1807 (N_1807,N_501,N_982);
nand U1808 (N_1808,N_285,N_695);
xor U1809 (N_1809,N_980,N_850);
xor U1810 (N_1810,N_614,N_777);
xnor U1811 (N_1811,N_537,N_396);
and U1812 (N_1812,N_968,N_507);
or U1813 (N_1813,N_425,N_951);
nand U1814 (N_1814,N_774,N_797);
nand U1815 (N_1815,N_243,N_969);
nand U1816 (N_1816,N_769,N_289);
nand U1817 (N_1817,N_923,N_927);
nand U1818 (N_1818,N_403,N_274);
xnor U1819 (N_1819,N_889,N_277);
and U1820 (N_1820,N_708,N_10);
or U1821 (N_1821,N_601,N_94);
or U1822 (N_1822,N_57,N_904);
nand U1823 (N_1823,N_156,N_792);
or U1824 (N_1824,N_791,N_356);
nand U1825 (N_1825,N_134,N_862);
and U1826 (N_1826,N_711,N_874);
xnor U1827 (N_1827,N_584,N_638);
or U1828 (N_1828,N_519,N_156);
and U1829 (N_1829,N_991,N_91);
and U1830 (N_1830,N_675,N_151);
nor U1831 (N_1831,N_265,N_123);
xor U1832 (N_1832,N_836,N_4);
or U1833 (N_1833,N_941,N_315);
nand U1834 (N_1834,N_997,N_252);
nand U1835 (N_1835,N_959,N_5);
or U1836 (N_1836,N_216,N_342);
and U1837 (N_1837,N_52,N_748);
and U1838 (N_1838,N_935,N_486);
nand U1839 (N_1839,N_325,N_714);
and U1840 (N_1840,N_392,N_257);
and U1841 (N_1841,N_657,N_181);
xor U1842 (N_1842,N_184,N_94);
or U1843 (N_1843,N_315,N_68);
and U1844 (N_1844,N_133,N_630);
or U1845 (N_1845,N_186,N_369);
and U1846 (N_1846,N_174,N_378);
and U1847 (N_1847,N_971,N_459);
nand U1848 (N_1848,N_330,N_642);
or U1849 (N_1849,N_546,N_835);
nor U1850 (N_1850,N_544,N_516);
nor U1851 (N_1851,N_29,N_345);
or U1852 (N_1852,N_463,N_757);
xnor U1853 (N_1853,N_224,N_560);
nor U1854 (N_1854,N_566,N_56);
and U1855 (N_1855,N_202,N_876);
nand U1856 (N_1856,N_608,N_844);
xor U1857 (N_1857,N_411,N_348);
nor U1858 (N_1858,N_273,N_68);
or U1859 (N_1859,N_827,N_32);
nand U1860 (N_1860,N_248,N_585);
and U1861 (N_1861,N_970,N_89);
and U1862 (N_1862,N_211,N_598);
xor U1863 (N_1863,N_905,N_243);
or U1864 (N_1864,N_290,N_983);
and U1865 (N_1865,N_74,N_906);
nand U1866 (N_1866,N_649,N_138);
and U1867 (N_1867,N_260,N_782);
and U1868 (N_1868,N_34,N_897);
or U1869 (N_1869,N_178,N_213);
or U1870 (N_1870,N_584,N_147);
or U1871 (N_1871,N_767,N_366);
and U1872 (N_1872,N_735,N_560);
xor U1873 (N_1873,N_926,N_72);
or U1874 (N_1874,N_258,N_338);
nor U1875 (N_1875,N_475,N_537);
nor U1876 (N_1876,N_224,N_338);
nand U1877 (N_1877,N_480,N_686);
nand U1878 (N_1878,N_691,N_481);
or U1879 (N_1879,N_715,N_739);
xor U1880 (N_1880,N_398,N_490);
nor U1881 (N_1881,N_172,N_961);
nor U1882 (N_1882,N_810,N_920);
and U1883 (N_1883,N_292,N_317);
nand U1884 (N_1884,N_504,N_314);
nand U1885 (N_1885,N_138,N_915);
nor U1886 (N_1886,N_600,N_802);
nand U1887 (N_1887,N_655,N_320);
or U1888 (N_1888,N_768,N_283);
or U1889 (N_1889,N_471,N_822);
and U1890 (N_1890,N_335,N_297);
nand U1891 (N_1891,N_139,N_158);
nor U1892 (N_1892,N_997,N_843);
nand U1893 (N_1893,N_727,N_127);
or U1894 (N_1894,N_39,N_515);
and U1895 (N_1895,N_282,N_621);
nor U1896 (N_1896,N_472,N_522);
or U1897 (N_1897,N_435,N_467);
nand U1898 (N_1898,N_401,N_762);
and U1899 (N_1899,N_221,N_125);
nor U1900 (N_1900,N_396,N_535);
nor U1901 (N_1901,N_0,N_667);
xor U1902 (N_1902,N_805,N_52);
nand U1903 (N_1903,N_303,N_260);
nor U1904 (N_1904,N_66,N_397);
nand U1905 (N_1905,N_962,N_848);
and U1906 (N_1906,N_335,N_482);
and U1907 (N_1907,N_353,N_40);
or U1908 (N_1908,N_820,N_457);
or U1909 (N_1909,N_17,N_863);
nand U1910 (N_1910,N_92,N_942);
nand U1911 (N_1911,N_745,N_929);
xor U1912 (N_1912,N_435,N_571);
or U1913 (N_1913,N_933,N_957);
nand U1914 (N_1914,N_836,N_740);
nor U1915 (N_1915,N_977,N_646);
nand U1916 (N_1916,N_801,N_227);
nor U1917 (N_1917,N_538,N_469);
nand U1918 (N_1918,N_445,N_812);
and U1919 (N_1919,N_763,N_228);
or U1920 (N_1920,N_840,N_192);
nand U1921 (N_1921,N_120,N_878);
or U1922 (N_1922,N_217,N_172);
nand U1923 (N_1923,N_731,N_889);
and U1924 (N_1924,N_49,N_371);
or U1925 (N_1925,N_273,N_262);
and U1926 (N_1926,N_853,N_678);
and U1927 (N_1927,N_199,N_561);
or U1928 (N_1928,N_928,N_255);
or U1929 (N_1929,N_223,N_192);
and U1930 (N_1930,N_981,N_219);
nor U1931 (N_1931,N_216,N_818);
nor U1932 (N_1932,N_203,N_436);
and U1933 (N_1933,N_767,N_31);
nand U1934 (N_1934,N_972,N_818);
xor U1935 (N_1935,N_376,N_863);
xor U1936 (N_1936,N_126,N_36);
xnor U1937 (N_1937,N_394,N_740);
nand U1938 (N_1938,N_104,N_791);
xor U1939 (N_1939,N_917,N_577);
or U1940 (N_1940,N_213,N_860);
and U1941 (N_1941,N_121,N_897);
or U1942 (N_1942,N_203,N_807);
or U1943 (N_1943,N_627,N_149);
and U1944 (N_1944,N_337,N_753);
or U1945 (N_1945,N_235,N_882);
xnor U1946 (N_1946,N_383,N_744);
nor U1947 (N_1947,N_697,N_973);
or U1948 (N_1948,N_846,N_895);
nor U1949 (N_1949,N_818,N_265);
and U1950 (N_1950,N_985,N_434);
nor U1951 (N_1951,N_748,N_611);
nand U1952 (N_1952,N_716,N_64);
nand U1953 (N_1953,N_21,N_597);
nand U1954 (N_1954,N_779,N_734);
or U1955 (N_1955,N_94,N_810);
nand U1956 (N_1956,N_453,N_230);
and U1957 (N_1957,N_560,N_79);
nand U1958 (N_1958,N_948,N_79);
nand U1959 (N_1959,N_465,N_724);
and U1960 (N_1960,N_606,N_412);
or U1961 (N_1961,N_401,N_481);
xor U1962 (N_1962,N_775,N_332);
xnor U1963 (N_1963,N_288,N_639);
xor U1964 (N_1964,N_535,N_1);
nand U1965 (N_1965,N_330,N_875);
nand U1966 (N_1966,N_924,N_15);
xnor U1967 (N_1967,N_611,N_247);
nand U1968 (N_1968,N_362,N_295);
and U1969 (N_1969,N_339,N_628);
nor U1970 (N_1970,N_858,N_832);
nand U1971 (N_1971,N_302,N_295);
nor U1972 (N_1972,N_318,N_928);
and U1973 (N_1973,N_474,N_870);
and U1974 (N_1974,N_759,N_52);
nand U1975 (N_1975,N_626,N_600);
and U1976 (N_1976,N_108,N_578);
nor U1977 (N_1977,N_713,N_622);
nor U1978 (N_1978,N_972,N_19);
nand U1979 (N_1979,N_42,N_128);
or U1980 (N_1980,N_790,N_879);
nand U1981 (N_1981,N_603,N_650);
and U1982 (N_1982,N_621,N_256);
nand U1983 (N_1983,N_97,N_107);
and U1984 (N_1984,N_486,N_392);
nand U1985 (N_1985,N_743,N_577);
and U1986 (N_1986,N_976,N_883);
nand U1987 (N_1987,N_464,N_27);
or U1988 (N_1988,N_574,N_598);
or U1989 (N_1989,N_458,N_197);
or U1990 (N_1990,N_61,N_69);
nand U1991 (N_1991,N_163,N_186);
xor U1992 (N_1992,N_158,N_13);
or U1993 (N_1993,N_479,N_931);
or U1994 (N_1994,N_170,N_85);
and U1995 (N_1995,N_320,N_777);
nand U1996 (N_1996,N_554,N_677);
or U1997 (N_1997,N_470,N_234);
and U1998 (N_1998,N_572,N_327);
xor U1999 (N_1999,N_547,N_395);
nor U2000 (N_2000,N_1129,N_1442);
xor U2001 (N_2001,N_1887,N_1773);
nand U2002 (N_2002,N_1635,N_1600);
nand U2003 (N_2003,N_1058,N_1257);
xnor U2004 (N_2004,N_1333,N_1860);
nor U2005 (N_2005,N_1493,N_1593);
nand U2006 (N_2006,N_1694,N_1060);
xor U2007 (N_2007,N_1581,N_1548);
nor U2008 (N_2008,N_1578,N_1701);
nand U2009 (N_2009,N_1680,N_1262);
and U2010 (N_2010,N_1774,N_1647);
nor U2011 (N_2011,N_1859,N_1185);
nand U2012 (N_2012,N_1758,N_1072);
or U2013 (N_2013,N_1220,N_1959);
nand U2014 (N_2014,N_1381,N_1208);
nor U2015 (N_2015,N_1321,N_1173);
nand U2016 (N_2016,N_1083,N_1681);
nand U2017 (N_2017,N_1102,N_1078);
nand U2018 (N_2018,N_1624,N_1994);
and U2019 (N_2019,N_1122,N_1944);
and U2020 (N_2020,N_1753,N_1157);
and U2021 (N_2021,N_1455,N_1249);
nor U2022 (N_2022,N_1534,N_1799);
nand U2023 (N_2023,N_1491,N_1747);
and U2024 (N_2024,N_1268,N_1974);
or U2025 (N_2025,N_1383,N_1246);
nor U2026 (N_2026,N_1477,N_1226);
nor U2027 (N_2027,N_1948,N_1672);
or U2028 (N_2028,N_1530,N_1025);
nand U2029 (N_2029,N_1167,N_1481);
or U2030 (N_2030,N_1568,N_1588);
or U2031 (N_2031,N_1721,N_1320);
nor U2032 (N_2032,N_1404,N_1825);
and U2033 (N_2033,N_1334,N_1685);
or U2034 (N_2034,N_1158,N_1499);
or U2035 (N_2035,N_1171,N_1750);
and U2036 (N_2036,N_1931,N_1990);
nor U2037 (N_2037,N_1437,N_1461);
nor U2038 (N_2038,N_1095,N_1292);
nand U2039 (N_2039,N_1483,N_1506);
and U2040 (N_2040,N_1682,N_1756);
and U2041 (N_2041,N_1143,N_1676);
and U2042 (N_2042,N_1263,N_1550);
nand U2043 (N_2043,N_1638,N_1772);
nand U2044 (N_2044,N_1553,N_1179);
or U2045 (N_2045,N_1340,N_1947);
xor U2046 (N_2046,N_1920,N_1536);
and U2047 (N_2047,N_1401,N_1514);
nand U2048 (N_2048,N_1669,N_1807);
or U2049 (N_2049,N_1659,N_1402);
xnor U2050 (N_2050,N_1011,N_1443);
nand U2051 (N_2051,N_1365,N_1995);
or U2052 (N_2052,N_1728,N_1511);
nand U2053 (N_2053,N_1003,N_1020);
or U2054 (N_2054,N_1832,N_1719);
or U2055 (N_2055,N_1159,N_1956);
nor U2056 (N_2056,N_1771,N_1776);
nand U2057 (N_2057,N_1643,N_1561);
nand U2058 (N_2058,N_1252,N_1923);
and U2059 (N_2059,N_1196,N_1356);
or U2060 (N_2060,N_1325,N_1068);
and U2061 (N_2061,N_1501,N_1720);
nand U2062 (N_2062,N_1114,N_1762);
or U2063 (N_2063,N_1890,N_1833);
nor U2064 (N_2064,N_1057,N_1961);
or U2065 (N_2065,N_1070,N_1378);
or U2066 (N_2066,N_1801,N_1871);
nand U2067 (N_2067,N_1282,N_1535);
xnor U2068 (N_2068,N_1693,N_1949);
or U2069 (N_2069,N_1526,N_1836);
nand U2070 (N_2070,N_1872,N_1022);
and U2071 (N_2071,N_1877,N_1140);
or U2072 (N_2072,N_1579,N_1782);
nand U2073 (N_2073,N_1665,N_1010);
and U2074 (N_2074,N_1644,N_1136);
and U2075 (N_2075,N_1864,N_1898);
and U2076 (N_2076,N_1465,N_1075);
or U2077 (N_2077,N_1970,N_1894);
nand U2078 (N_2078,N_1690,N_1323);
nand U2079 (N_2079,N_1658,N_1538);
xnor U2080 (N_2080,N_1373,N_1398);
and U2081 (N_2081,N_1188,N_1101);
and U2082 (N_2082,N_1130,N_1521);
or U2083 (N_2083,N_1251,N_1951);
or U2084 (N_2084,N_1086,N_1395);
or U2085 (N_2085,N_1955,N_1827);
or U2086 (N_2086,N_1903,N_1397);
and U2087 (N_2087,N_1926,N_1525);
nand U2088 (N_2088,N_1794,N_1749);
or U2089 (N_2089,N_1004,N_1627);
and U2090 (N_2090,N_1908,N_1983);
or U2091 (N_2091,N_1494,N_1766);
and U2092 (N_2092,N_1213,N_1107);
nor U2093 (N_2093,N_1940,N_1376);
nor U2094 (N_2094,N_1123,N_1989);
and U2095 (N_2095,N_1834,N_1326);
nand U2096 (N_2096,N_1718,N_1973);
or U2097 (N_2097,N_1456,N_1472);
and U2098 (N_2098,N_1524,N_1614);
or U2099 (N_2099,N_1988,N_1050);
nand U2100 (N_2100,N_1338,N_1375);
nor U2101 (N_2101,N_1116,N_1838);
nor U2102 (N_2102,N_1190,N_1419);
and U2103 (N_2103,N_1138,N_1270);
and U2104 (N_2104,N_1181,N_1977);
or U2105 (N_2105,N_1119,N_1717);
xor U2106 (N_2106,N_1929,N_1054);
xor U2107 (N_2107,N_1163,N_1307);
nand U2108 (N_2108,N_1350,N_1784);
xnor U2109 (N_2109,N_1653,N_1967);
xnor U2110 (N_2110,N_1002,N_1149);
or U2111 (N_2111,N_1556,N_1291);
nor U2112 (N_2112,N_1731,N_1780);
nand U2113 (N_2113,N_1469,N_1045);
nand U2114 (N_2114,N_1222,N_1869);
and U2115 (N_2115,N_1424,N_1473);
nand U2116 (N_2116,N_1539,N_1080);
nand U2117 (N_2117,N_1839,N_1508);
or U2118 (N_2118,N_1622,N_1372);
nand U2119 (N_2119,N_1269,N_1632);
and U2120 (N_2120,N_1374,N_1710);
xnor U2121 (N_2121,N_1266,N_1031);
and U2122 (N_2122,N_1065,N_1904);
or U2123 (N_2123,N_1607,N_1626);
nor U2124 (N_2124,N_1309,N_1432);
or U2125 (N_2125,N_1633,N_1905);
and U2126 (N_2126,N_1178,N_1862);
nor U2127 (N_2127,N_1815,N_1552);
nor U2128 (N_2128,N_1428,N_1889);
and U2129 (N_2129,N_1620,N_1554);
or U2130 (N_2130,N_1283,N_1162);
nand U2131 (N_2131,N_1744,N_1357);
nand U2132 (N_2132,N_1751,N_1657);
nand U2133 (N_2133,N_1301,N_1921);
nand U2134 (N_2134,N_1980,N_1699);
and U2135 (N_2135,N_1788,N_1354);
nand U2136 (N_2136,N_1169,N_1892);
and U2137 (N_2137,N_1802,N_1950);
nand U2138 (N_2138,N_1924,N_1106);
and U2139 (N_2139,N_1144,N_1015);
or U2140 (N_2140,N_1186,N_1569);
nand U2141 (N_2141,N_1384,N_1998);
nor U2142 (N_2142,N_1727,N_1132);
and U2143 (N_2143,N_1368,N_1580);
nor U2144 (N_2144,N_1849,N_1230);
or U2145 (N_2145,N_1351,N_1881);
nand U2146 (N_2146,N_1233,N_1152);
or U2147 (N_2147,N_1987,N_1935);
xor U2148 (N_2148,N_1930,N_1822);
nor U2149 (N_2149,N_1891,N_1285);
nand U2150 (N_2150,N_1203,N_1012);
nor U2151 (N_2151,N_1901,N_1367);
xor U2152 (N_2152,N_1545,N_1558);
and U2153 (N_2153,N_1431,N_1434);
nor U2154 (N_2154,N_1147,N_1399);
xnor U2155 (N_2155,N_1958,N_1709);
xor U2156 (N_2156,N_1996,N_1359);
and U2157 (N_2157,N_1253,N_1243);
and U2158 (N_2158,N_1430,N_1021);
nand U2159 (N_2159,N_1039,N_1759);
or U2160 (N_2160,N_1444,N_1298);
or U2161 (N_2161,N_1606,N_1724);
nand U2162 (N_2162,N_1867,N_1209);
or U2163 (N_2163,N_1515,N_1512);
and U2164 (N_2164,N_1315,N_1571);
xor U2165 (N_2165,N_1168,N_1572);
and U2166 (N_2166,N_1407,N_1734);
nor U2167 (N_2167,N_1077,N_1616);
xnor U2168 (N_2168,N_1370,N_1532);
and U2169 (N_2169,N_1589,N_1599);
nand U2170 (N_2170,N_1245,N_1023);
or U2171 (N_2171,N_1284,N_1183);
and U2172 (N_2172,N_1646,N_1651);
nor U2173 (N_2173,N_1069,N_1343);
xnor U2174 (N_2174,N_1059,N_1071);
and U2175 (N_2175,N_1590,N_1198);
or U2176 (N_2176,N_1857,N_1886);
nor U2177 (N_2177,N_1715,N_1133);
and U2178 (N_2178,N_1382,N_1166);
nor U2179 (N_2179,N_1306,N_1618);
and U2180 (N_2180,N_1513,N_1033);
nor U2181 (N_2181,N_1331,N_1479);
nand U2182 (N_2182,N_1153,N_1703);
and U2183 (N_2183,N_1969,N_1668);
nor U2184 (N_2184,N_1797,N_1700);
or U2185 (N_2185,N_1229,N_1953);
nand U2186 (N_2186,N_1820,N_1936);
nor U2187 (N_2187,N_1805,N_1853);
and U2188 (N_2188,N_1986,N_1244);
nor U2189 (N_2189,N_1408,N_1108);
nor U2190 (N_2190,N_1981,N_1504);
nand U2191 (N_2191,N_1966,N_1206);
xnor U2192 (N_2192,N_1598,N_1517);
and U2193 (N_2193,N_1278,N_1195);
and U2194 (N_2194,N_1613,N_1870);
nor U2195 (N_2195,N_1850,N_1741);
nor U2196 (N_2196,N_1110,N_1276);
or U2197 (N_2197,N_1675,N_1174);
nor U2198 (N_2198,N_1748,N_1844);
nor U2199 (N_2199,N_1722,N_1621);
or U2200 (N_2200,N_1678,N_1848);
or U2201 (N_2201,N_1803,N_1705);
and U2202 (N_2202,N_1605,N_1319);
nor U2203 (N_2203,N_1451,N_1418);
nor U2204 (N_2204,N_1218,N_1063);
nand U2205 (N_2205,N_1507,N_1677);
nand U2206 (N_2206,N_1294,N_1938);
or U2207 (N_2207,N_1217,N_1236);
or U2208 (N_2208,N_1785,N_1649);
or U2209 (N_2209,N_1641,N_1363);
or U2210 (N_2210,N_1197,N_1429);
and U2211 (N_2211,N_1868,N_1317);
or U2212 (N_2212,N_1629,N_1313);
xor U2213 (N_2213,N_1855,N_1177);
and U2214 (N_2214,N_1001,N_1962);
and U2215 (N_2215,N_1449,N_1422);
nand U2216 (N_2216,N_1231,N_1735);
and U2217 (N_2217,N_1366,N_1349);
or U2218 (N_2218,N_1040,N_1737);
and U2219 (N_2219,N_1946,N_1876);
nor U2220 (N_2220,N_1380,N_1046);
nor U2221 (N_2221,N_1533,N_1126);
xnor U2222 (N_2222,N_1726,N_1330);
and U2223 (N_2223,N_1723,N_1255);
xor U2224 (N_2224,N_1189,N_1563);
or U2225 (N_2225,N_1085,N_1609);
xor U2226 (N_2226,N_1910,N_1851);
or U2227 (N_2227,N_1041,N_1982);
nor U2228 (N_2228,N_1683,N_1312);
nor U2229 (N_2229,N_1435,N_1076);
and U2230 (N_2230,N_1937,N_1463);
xnor U2231 (N_2231,N_1884,N_1852);
xnor U2232 (N_2232,N_1329,N_1939);
nor U2233 (N_2233,N_1302,N_1281);
nand U2234 (N_2234,N_1056,N_1035);
or U2235 (N_2235,N_1628,N_1297);
or U2236 (N_2236,N_1652,N_1656);
nor U2237 (N_2237,N_1201,N_1714);
or U2238 (N_2238,N_1207,N_1945);
and U2239 (N_2239,N_1725,N_1360);
nor U2240 (N_2240,N_1711,N_1248);
or U2241 (N_2241,N_1907,N_1492);
and U2242 (N_2242,N_1767,N_1342);
xnor U2243 (N_2243,N_1007,N_1089);
or U2244 (N_2244,N_1441,N_1345);
or U2245 (N_2245,N_1223,N_1663);
nor U2246 (N_2246,N_1642,N_1446);
nand U2247 (N_2247,N_1752,N_1810);
nor U2248 (N_2248,N_1586,N_1423);
and U2249 (N_2249,N_1991,N_1739);
and U2250 (N_2250,N_1490,N_1707);
nor U2251 (N_2251,N_1503,N_1567);
or U2252 (N_2252,N_1893,N_1030);
nor U2253 (N_2253,N_1165,N_1238);
nand U2254 (N_2254,N_1120,N_1671);
nor U2255 (N_2255,N_1564,N_1362);
xor U2256 (N_2256,N_1043,N_1537);
nor U2257 (N_2257,N_1170,N_1691);
and U2258 (N_2258,N_1648,N_1640);
or U2259 (N_2259,N_1470,N_1425);
or U2260 (N_2260,N_1505,N_1420);
nand U2261 (N_2261,N_1768,N_1639);
nand U2262 (N_2262,N_1034,N_1702);
or U2263 (N_2263,N_1295,N_1352);
nand U2264 (N_2264,N_1176,N_1061);
or U2265 (N_2265,N_1017,N_1666);
xor U2266 (N_2266,N_1300,N_1156);
nand U2267 (N_2267,N_1498,N_1142);
nand U2268 (N_2268,N_1879,N_1601);
and U2269 (N_2269,N_1228,N_1786);
or U2270 (N_2270,N_1105,N_1664);
or U2271 (N_2271,N_1919,N_1127);
nand U2272 (N_2272,N_1293,N_1496);
nor U2273 (N_2273,N_1760,N_1976);
or U2274 (N_2274,N_1286,N_1194);
nor U2275 (N_2275,N_1448,N_1670);
or U2276 (N_2276,N_1172,N_1414);
nand U2277 (N_2277,N_1846,N_1275);
or U2278 (N_2278,N_1305,N_1112);
and U2279 (N_2279,N_1592,N_1385);
nand U2280 (N_2280,N_1324,N_1912);
nand U2281 (N_2281,N_1712,N_1014);
nand U2282 (N_2282,N_1055,N_1510);
nor U2283 (N_2283,N_1817,N_1204);
and U2284 (N_2284,N_1497,N_1250);
or U2285 (N_2285,N_1617,N_1235);
and U2286 (N_2286,N_1073,N_1740);
nor U2287 (N_2287,N_1316,N_1091);
or U2288 (N_2288,N_1079,N_1933);
nor U2289 (N_2289,N_1775,N_1484);
or U2290 (N_2290,N_1916,N_1963);
and U2291 (N_2291,N_1742,N_1322);
nor U2292 (N_2292,N_1390,N_1387);
nor U2293 (N_2293,N_1013,N_1038);
nor U2294 (N_2294,N_1978,N_1733);
nand U2295 (N_2295,N_1746,N_1625);
nand U2296 (N_2296,N_1290,N_1103);
nand U2297 (N_2297,N_1093,N_1232);
and U2298 (N_2298,N_1769,N_1895);
xnor U2299 (N_2299,N_1518,N_1743);
nor U2300 (N_2300,N_1224,N_1090);
or U2301 (N_2301,N_1761,N_1234);
and U2302 (N_2302,N_1450,N_1814);
or U2303 (N_2303,N_1409,N_1225);
nand U2304 (N_2304,N_1464,N_1067);
or U2305 (N_2305,N_1485,N_1125);
and U2306 (N_2306,N_1979,N_1115);
nand U2307 (N_2307,N_1732,N_1335);
nor U2308 (N_2308,N_1328,N_1909);
nor U2309 (N_2309,N_1459,N_1109);
nor U2310 (N_2310,N_1151,N_1812);
nand U2311 (N_2311,N_1882,N_1866);
nor U2312 (N_2312,N_1928,N_1026);
or U2313 (N_2313,N_1098,N_1818);
nor U2314 (N_2314,N_1476,N_1457);
nand U2315 (N_2315,N_1288,N_1687);
or U2316 (N_2316,N_1081,N_1261);
and U2317 (N_2317,N_1828,N_1674);
nor U2318 (N_2318,N_1673,N_1154);
nor U2319 (N_2319,N_1242,N_1965);
nor U2320 (N_2320,N_1787,N_1911);
or U2321 (N_2321,N_1412,N_1544);
nor U2322 (N_2322,N_1934,N_1445);
and U2323 (N_2323,N_1689,N_1612);
nor U2324 (N_2324,N_1210,N_1264);
nor U2325 (N_2325,N_1371,N_1764);
or U2326 (N_2326,N_1800,N_1527);
and U2327 (N_2327,N_1557,N_1032);
or U2328 (N_2328,N_1161,N_1272);
xor U2329 (N_2329,N_1028,N_1062);
and U2330 (N_2330,N_1051,N_1917);
nand U2331 (N_2331,N_1792,N_1053);
nor U2332 (N_2332,N_1611,N_1662);
nand U2333 (N_2333,N_1755,N_1708);
nor U2334 (N_2334,N_1417,N_1466);
xor U2335 (N_2335,N_1280,N_1636);
nand U2336 (N_2336,N_1205,N_1826);
nor U2337 (N_2337,N_1808,N_1964);
nand U2338 (N_2338,N_1241,N_1303);
nor U2339 (N_2339,N_1757,N_1403);
or U2340 (N_2340,N_1576,N_1654);
nor U2341 (N_2341,N_1202,N_1922);
nand U2342 (N_2342,N_1440,N_1623);
nand U2343 (N_2343,N_1570,N_1645);
nor U2344 (N_2344,N_1856,N_1388);
nor U2345 (N_2345,N_1139,N_1842);
nand U2346 (N_2346,N_1259,N_1531);
nand U2347 (N_2347,N_1566,N_1555);
or U2348 (N_2348,N_1899,N_1631);
nor U2349 (N_2349,N_1471,N_1716);
and U2350 (N_2350,N_1873,N_1094);
and U2351 (N_2351,N_1415,N_1952);
and U2352 (N_2352,N_1124,N_1954);
or U2353 (N_2353,N_1861,N_1346);
nor U2354 (N_2354,N_1630,N_1522);
xor U2355 (N_2355,N_1468,N_1047);
nor U2356 (N_2356,N_1064,N_1829);
nor U2357 (N_2357,N_1216,N_1361);
and U2358 (N_2358,N_1247,N_1793);
nand U2359 (N_2359,N_1688,N_1379);
xor U2360 (N_2360,N_1968,N_1650);
nor U2361 (N_2361,N_1509,N_1005);
nor U2362 (N_2362,N_1239,N_1474);
nand U2363 (N_2363,N_1574,N_1128);
nand U2364 (N_2364,N_1655,N_1391);
and U2365 (N_2365,N_1480,N_1460);
or U2366 (N_2366,N_1896,N_1489);
or U2367 (N_2367,N_1192,N_1084);
xor U2368 (N_2368,N_1427,N_1837);
nand U2369 (N_2369,N_1809,N_1913);
nor U2370 (N_2370,N_1211,N_1018);
nor U2371 (N_2371,N_1679,N_1482);
nand U2372 (N_2372,N_1327,N_1118);
nor U2373 (N_2373,N_1187,N_1615);
and U2374 (N_2374,N_1344,N_1575);
or U2375 (N_2375,N_1540,N_1692);
nor U2376 (N_2376,N_1426,N_1393);
and U2377 (N_2377,N_1227,N_1155);
xnor U2378 (N_2378,N_1191,N_1289);
nor U2379 (N_2379,N_1215,N_1237);
nand U2380 (N_2380,N_1277,N_1500);
nand U2381 (N_2381,N_1847,N_1594);
nor U2382 (N_2382,N_1927,N_1273);
nand U2383 (N_2383,N_1583,N_1565);
or U2384 (N_2384,N_1475,N_1131);
nand U2385 (N_2385,N_1551,N_1560);
and U2386 (N_2386,N_1148,N_1897);
nor U2387 (N_2387,N_1405,N_1274);
and U2388 (N_2388,N_1821,N_1347);
and U2389 (N_2389,N_1591,N_1037);
nand U2390 (N_2390,N_1453,N_1008);
xnor U2391 (N_2391,N_1971,N_1394);
and U2392 (N_2392,N_1875,N_1137);
xor U2393 (N_2393,N_1845,N_1943);
and U2394 (N_2394,N_1695,N_1706);
nor U2395 (N_2395,N_1585,N_1914);
or U2396 (N_2396,N_1878,N_1097);
nor U2397 (N_2397,N_1738,N_1254);
xor U2398 (N_2398,N_1219,N_1637);
or U2399 (N_2399,N_1729,N_1487);
and U2400 (N_2400,N_1942,N_1549);
or U2401 (N_2401,N_1900,N_1212);
or U2402 (N_2402,N_1816,N_1660);
nor U2403 (N_2403,N_1100,N_1048);
nand U2404 (N_2404,N_1411,N_1495);
and U2405 (N_2405,N_1790,N_1164);
xor U2406 (N_2406,N_1182,N_1906);
nor U2407 (N_2407,N_1087,N_1713);
or U2408 (N_2408,N_1597,N_1146);
or U2409 (N_2409,N_1433,N_1027);
xor U2410 (N_2410,N_1813,N_1547);
or U2411 (N_2411,N_1529,N_1835);
nor U2412 (N_2412,N_1036,N_1364);
and U2413 (N_2413,N_1044,N_1256);
nand U2414 (N_2414,N_1462,N_1135);
or U2415 (N_2415,N_1406,N_1258);
nand U2416 (N_2416,N_1985,N_1796);
and U2417 (N_2417,N_1520,N_1193);
nor U2418 (N_2418,N_1042,N_1265);
and U2419 (N_2419,N_1602,N_1863);
nor U2420 (N_2420,N_1117,N_1999);
nor U2421 (N_2421,N_1634,N_1765);
nor U2422 (N_2422,N_1175,N_1113);
nand U2423 (N_2423,N_1436,N_1337);
or U2424 (N_2424,N_1299,N_1925);
nand U2425 (N_2425,N_1134,N_1369);
nand U2426 (N_2426,N_1488,N_1358);
or U2427 (N_2427,N_1355,N_1957);
or U2428 (N_2428,N_1918,N_1902);
nor U2429 (N_2429,N_1795,N_1543);
or U2430 (N_2430,N_1577,N_1377);
or U2431 (N_2431,N_1180,N_1467);
and U2432 (N_2432,N_1587,N_1972);
and U2433 (N_2433,N_1478,N_1318);
and U2434 (N_2434,N_1661,N_1145);
nor U2435 (N_2435,N_1019,N_1932);
and U2436 (N_2436,N_1573,N_1975);
nor U2437 (N_2437,N_1447,N_1854);
nand U2438 (N_2438,N_1562,N_1823);
and U2439 (N_2439,N_1271,N_1603);
and U2440 (N_2440,N_1696,N_1698);
nor U2441 (N_2441,N_1049,N_1960);
nand U2442 (N_2442,N_1074,N_1584);
nor U2443 (N_2443,N_1667,N_1883);
nor U2444 (N_2444,N_1778,N_1704);
nand U2445 (N_2445,N_1121,N_1619);
or U2446 (N_2446,N_1779,N_1066);
xor U2447 (N_2447,N_1610,N_1088);
and U2448 (N_2448,N_1546,N_1111);
or U2449 (N_2449,N_1353,N_1811);
or U2450 (N_2450,N_1184,N_1348);
nor U2451 (N_2451,N_1339,N_1806);
or U2452 (N_2452,N_1608,N_1596);
nand U2453 (N_2453,N_1410,N_1604);
xor U2454 (N_2454,N_1798,N_1885);
or U2455 (N_2455,N_1416,N_1824);
nand U2456 (N_2456,N_1684,N_1831);
nand U2457 (N_2457,N_1454,N_1009);
and U2458 (N_2458,N_1421,N_1000);
nor U2459 (N_2459,N_1804,N_1341);
or U2460 (N_2460,N_1016,N_1697);
nor U2461 (N_2461,N_1984,N_1199);
nor U2462 (N_2462,N_1096,N_1941);
nand U2463 (N_2463,N_1486,N_1915);
or U2464 (N_2464,N_1099,N_1542);
nor U2465 (N_2465,N_1841,N_1052);
or U2466 (N_2466,N_1843,N_1214);
nor U2467 (N_2467,N_1993,N_1783);
nand U2468 (N_2468,N_1686,N_1819);
xor U2469 (N_2469,N_1528,N_1858);
and U2470 (N_2470,N_1396,N_1439);
nand U2471 (N_2471,N_1736,N_1770);
nand U2472 (N_2472,N_1024,N_1314);
nor U2473 (N_2473,N_1413,N_1389);
nor U2474 (N_2474,N_1438,N_1559);
nand U2475 (N_2475,N_1595,N_1874);
nor U2476 (N_2476,N_1221,N_1458);
nand U2477 (N_2477,N_1332,N_1997);
nand U2478 (N_2478,N_1865,N_1200);
or U2479 (N_2479,N_1092,N_1279);
nand U2480 (N_2480,N_1400,N_1789);
nand U2481 (N_2481,N_1730,N_1888);
nor U2482 (N_2482,N_1519,N_1541);
and U2483 (N_2483,N_1781,N_1310);
nand U2484 (N_2484,N_1880,N_1992);
or U2485 (N_2485,N_1754,N_1240);
nand U2486 (N_2486,N_1304,N_1392);
and U2487 (N_2487,N_1150,N_1311);
or U2488 (N_2488,N_1452,N_1516);
nor U2489 (N_2489,N_1791,N_1260);
and U2490 (N_2490,N_1502,N_1777);
nand U2491 (N_2491,N_1082,N_1840);
nand U2492 (N_2492,N_1296,N_1287);
nand U2493 (N_2493,N_1745,N_1104);
and U2494 (N_2494,N_1029,N_1336);
nor U2495 (N_2495,N_1386,N_1141);
and U2496 (N_2496,N_1160,N_1582);
xnor U2497 (N_2497,N_1763,N_1308);
and U2498 (N_2498,N_1523,N_1267);
or U2499 (N_2499,N_1006,N_1830);
and U2500 (N_2500,N_1302,N_1376);
nor U2501 (N_2501,N_1324,N_1215);
and U2502 (N_2502,N_1398,N_1905);
nor U2503 (N_2503,N_1973,N_1403);
nor U2504 (N_2504,N_1610,N_1613);
nor U2505 (N_2505,N_1942,N_1014);
or U2506 (N_2506,N_1771,N_1697);
nor U2507 (N_2507,N_1531,N_1418);
nor U2508 (N_2508,N_1747,N_1204);
xnor U2509 (N_2509,N_1993,N_1772);
and U2510 (N_2510,N_1258,N_1051);
and U2511 (N_2511,N_1063,N_1624);
nand U2512 (N_2512,N_1886,N_1710);
and U2513 (N_2513,N_1113,N_1318);
and U2514 (N_2514,N_1803,N_1242);
and U2515 (N_2515,N_1658,N_1243);
or U2516 (N_2516,N_1338,N_1245);
nor U2517 (N_2517,N_1282,N_1032);
nor U2518 (N_2518,N_1000,N_1279);
or U2519 (N_2519,N_1508,N_1692);
nor U2520 (N_2520,N_1519,N_1943);
nand U2521 (N_2521,N_1432,N_1787);
nor U2522 (N_2522,N_1810,N_1342);
or U2523 (N_2523,N_1721,N_1678);
nor U2524 (N_2524,N_1883,N_1613);
and U2525 (N_2525,N_1152,N_1466);
xor U2526 (N_2526,N_1152,N_1782);
nor U2527 (N_2527,N_1135,N_1465);
and U2528 (N_2528,N_1406,N_1325);
nor U2529 (N_2529,N_1386,N_1172);
or U2530 (N_2530,N_1958,N_1891);
nand U2531 (N_2531,N_1839,N_1339);
or U2532 (N_2532,N_1761,N_1991);
nor U2533 (N_2533,N_1331,N_1912);
nor U2534 (N_2534,N_1313,N_1450);
xnor U2535 (N_2535,N_1235,N_1201);
and U2536 (N_2536,N_1472,N_1326);
and U2537 (N_2537,N_1951,N_1052);
nand U2538 (N_2538,N_1667,N_1698);
nor U2539 (N_2539,N_1830,N_1320);
or U2540 (N_2540,N_1464,N_1314);
nor U2541 (N_2541,N_1090,N_1830);
and U2542 (N_2542,N_1051,N_1322);
or U2543 (N_2543,N_1688,N_1575);
nor U2544 (N_2544,N_1630,N_1022);
xor U2545 (N_2545,N_1266,N_1861);
nor U2546 (N_2546,N_1661,N_1783);
nand U2547 (N_2547,N_1283,N_1199);
nor U2548 (N_2548,N_1901,N_1035);
or U2549 (N_2549,N_1850,N_1580);
nor U2550 (N_2550,N_1203,N_1147);
and U2551 (N_2551,N_1467,N_1582);
nand U2552 (N_2552,N_1976,N_1873);
nand U2553 (N_2553,N_1853,N_1922);
or U2554 (N_2554,N_1796,N_1613);
nand U2555 (N_2555,N_1959,N_1020);
or U2556 (N_2556,N_1625,N_1579);
or U2557 (N_2557,N_1639,N_1130);
or U2558 (N_2558,N_1679,N_1056);
and U2559 (N_2559,N_1886,N_1164);
and U2560 (N_2560,N_1922,N_1438);
nand U2561 (N_2561,N_1689,N_1771);
nand U2562 (N_2562,N_1991,N_1464);
nand U2563 (N_2563,N_1471,N_1306);
nor U2564 (N_2564,N_1099,N_1114);
nor U2565 (N_2565,N_1765,N_1995);
nand U2566 (N_2566,N_1312,N_1558);
and U2567 (N_2567,N_1061,N_1123);
nand U2568 (N_2568,N_1082,N_1921);
nor U2569 (N_2569,N_1338,N_1987);
or U2570 (N_2570,N_1695,N_1771);
and U2571 (N_2571,N_1103,N_1209);
and U2572 (N_2572,N_1608,N_1224);
nor U2573 (N_2573,N_1721,N_1869);
nand U2574 (N_2574,N_1207,N_1856);
nand U2575 (N_2575,N_1254,N_1508);
xnor U2576 (N_2576,N_1683,N_1400);
nand U2577 (N_2577,N_1806,N_1421);
nand U2578 (N_2578,N_1599,N_1485);
nand U2579 (N_2579,N_1338,N_1556);
nand U2580 (N_2580,N_1760,N_1036);
or U2581 (N_2581,N_1296,N_1858);
nor U2582 (N_2582,N_1029,N_1402);
or U2583 (N_2583,N_1476,N_1459);
nor U2584 (N_2584,N_1160,N_1743);
nand U2585 (N_2585,N_1732,N_1744);
and U2586 (N_2586,N_1616,N_1215);
xnor U2587 (N_2587,N_1036,N_1356);
nand U2588 (N_2588,N_1338,N_1772);
nor U2589 (N_2589,N_1464,N_1535);
nor U2590 (N_2590,N_1029,N_1871);
xor U2591 (N_2591,N_1208,N_1043);
nand U2592 (N_2592,N_1230,N_1221);
and U2593 (N_2593,N_1477,N_1814);
nand U2594 (N_2594,N_1283,N_1544);
nand U2595 (N_2595,N_1571,N_1263);
and U2596 (N_2596,N_1777,N_1679);
and U2597 (N_2597,N_1178,N_1049);
nand U2598 (N_2598,N_1670,N_1158);
and U2599 (N_2599,N_1590,N_1175);
nand U2600 (N_2600,N_1439,N_1644);
nand U2601 (N_2601,N_1915,N_1767);
and U2602 (N_2602,N_1446,N_1575);
or U2603 (N_2603,N_1650,N_1048);
and U2604 (N_2604,N_1068,N_1629);
and U2605 (N_2605,N_1347,N_1547);
nand U2606 (N_2606,N_1708,N_1551);
xor U2607 (N_2607,N_1203,N_1728);
nand U2608 (N_2608,N_1993,N_1041);
xnor U2609 (N_2609,N_1098,N_1298);
xor U2610 (N_2610,N_1405,N_1402);
and U2611 (N_2611,N_1106,N_1308);
nand U2612 (N_2612,N_1592,N_1038);
and U2613 (N_2613,N_1237,N_1396);
nor U2614 (N_2614,N_1026,N_1547);
and U2615 (N_2615,N_1153,N_1817);
and U2616 (N_2616,N_1079,N_1531);
and U2617 (N_2617,N_1925,N_1686);
nor U2618 (N_2618,N_1131,N_1718);
xor U2619 (N_2619,N_1444,N_1246);
and U2620 (N_2620,N_1095,N_1485);
or U2621 (N_2621,N_1505,N_1024);
nand U2622 (N_2622,N_1750,N_1996);
or U2623 (N_2623,N_1344,N_1908);
nand U2624 (N_2624,N_1836,N_1606);
nand U2625 (N_2625,N_1609,N_1280);
or U2626 (N_2626,N_1180,N_1298);
xor U2627 (N_2627,N_1176,N_1852);
nor U2628 (N_2628,N_1743,N_1639);
nand U2629 (N_2629,N_1089,N_1748);
nand U2630 (N_2630,N_1388,N_1941);
nor U2631 (N_2631,N_1008,N_1019);
xnor U2632 (N_2632,N_1515,N_1376);
nand U2633 (N_2633,N_1159,N_1839);
or U2634 (N_2634,N_1959,N_1103);
and U2635 (N_2635,N_1589,N_1502);
or U2636 (N_2636,N_1286,N_1568);
xnor U2637 (N_2637,N_1218,N_1261);
or U2638 (N_2638,N_1776,N_1874);
and U2639 (N_2639,N_1388,N_1153);
xor U2640 (N_2640,N_1815,N_1519);
nand U2641 (N_2641,N_1492,N_1444);
nor U2642 (N_2642,N_1606,N_1350);
or U2643 (N_2643,N_1718,N_1858);
and U2644 (N_2644,N_1691,N_1807);
nand U2645 (N_2645,N_1113,N_1209);
or U2646 (N_2646,N_1095,N_1192);
nand U2647 (N_2647,N_1562,N_1875);
and U2648 (N_2648,N_1394,N_1622);
and U2649 (N_2649,N_1872,N_1631);
nor U2650 (N_2650,N_1370,N_1341);
xor U2651 (N_2651,N_1155,N_1121);
nor U2652 (N_2652,N_1662,N_1312);
nor U2653 (N_2653,N_1364,N_1554);
nand U2654 (N_2654,N_1572,N_1204);
xor U2655 (N_2655,N_1810,N_1656);
nand U2656 (N_2656,N_1633,N_1461);
xnor U2657 (N_2657,N_1420,N_1133);
and U2658 (N_2658,N_1623,N_1359);
or U2659 (N_2659,N_1928,N_1439);
or U2660 (N_2660,N_1917,N_1121);
nor U2661 (N_2661,N_1298,N_1771);
and U2662 (N_2662,N_1706,N_1200);
nand U2663 (N_2663,N_1466,N_1179);
nand U2664 (N_2664,N_1966,N_1993);
xor U2665 (N_2665,N_1596,N_1579);
xnor U2666 (N_2666,N_1202,N_1639);
nand U2667 (N_2667,N_1261,N_1300);
or U2668 (N_2668,N_1316,N_1980);
xnor U2669 (N_2669,N_1749,N_1014);
nor U2670 (N_2670,N_1786,N_1636);
nand U2671 (N_2671,N_1479,N_1997);
nand U2672 (N_2672,N_1880,N_1103);
or U2673 (N_2673,N_1172,N_1077);
nor U2674 (N_2674,N_1807,N_1002);
nand U2675 (N_2675,N_1447,N_1395);
or U2676 (N_2676,N_1357,N_1114);
and U2677 (N_2677,N_1677,N_1369);
xor U2678 (N_2678,N_1090,N_1432);
xor U2679 (N_2679,N_1419,N_1959);
or U2680 (N_2680,N_1532,N_1044);
nand U2681 (N_2681,N_1100,N_1306);
nor U2682 (N_2682,N_1683,N_1012);
or U2683 (N_2683,N_1748,N_1301);
xor U2684 (N_2684,N_1862,N_1430);
or U2685 (N_2685,N_1693,N_1432);
and U2686 (N_2686,N_1481,N_1893);
and U2687 (N_2687,N_1063,N_1438);
nand U2688 (N_2688,N_1702,N_1751);
or U2689 (N_2689,N_1259,N_1968);
and U2690 (N_2690,N_1165,N_1061);
xor U2691 (N_2691,N_1206,N_1374);
nand U2692 (N_2692,N_1185,N_1109);
nor U2693 (N_2693,N_1454,N_1408);
or U2694 (N_2694,N_1187,N_1332);
and U2695 (N_2695,N_1303,N_1464);
nor U2696 (N_2696,N_1846,N_1520);
nor U2697 (N_2697,N_1449,N_1796);
and U2698 (N_2698,N_1193,N_1798);
or U2699 (N_2699,N_1136,N_1046);
nand U2700 (N_2700,N_1098,N_1967);
nor U2701 (N_2701,N_1987,N_1230);
or U2702 (N_2702,N_1850,N_1313);
nor U2703 (N_2703,N_1600,N_1521);
nand U2704 (N_2704,N_1044,N_1517);
nand U2705 (N_2705,N_1130,N_1961);
or U2706 (N_2706,N_1127,N_1183);
and U2707 (N_2707,N_1223,N_1066);
and U2708 (N_2708,N_1038,N_1386);
xor U2709 (N_2709,N_1456,N_1902);
or U2710 (N_2710,N_1811,N_1820);
and U2711 (N_2711,N_1092,N_1065);
nand U2712 (N_2712,N_1457,N_1988);
or U2713 (N_2713,N_1071,N_1572);
nand U2714 (N_2714,N_1164,N_1725);
or U2715 (N_2715,N_1631,N_1466);
and U2716 (N_2716,N_1086,N_1036);
and U2717 (N_2717,N_1907,N_1267);
and U2718 (N_2718,N_1114,N_1126);
nor U2719 (N_2719,N_1615,N_1509);
nor U2720 (N_2720,N_1896,N_1368);
xor U2721 (N_2721,N_1289,N_1157);
and U2722 (N_2722,N_1324,N_1839);
nor U2723 (N_2723,N_1457,N_1497);
or U2724 (N_2724,N_1726,N_1418);
nor U2725 (N_2725,N_1372,N_1773);
nand U2726 (N_2726,N_1676,N_1683);
or U2727 (N_2727,N_1743,N_1420);
nand U2728 (N_2728,N_1914,N_1279);
nor U2729 (N_2729,N_1178,N_1033);
nand U2730 (N_2730,N_1090,N_1016);
and U2731 (N_2731,N_1451,N_1703);
nand U2732 (N_2732,N_1004,N_1112);
nand U2733 (N_2733,N_1961,N_1706);
nand U2734 (N_2734,N_1355,N_1280);
nand U2735 (N_2735,N_1298,N_1418);
or U2736 (N_2736,N_1144,N_1729);
and U2737 (N_2737,N_1543,N_1991);
nand U2738 (N_2738,N_1701,N_1626);
nor U2739 (N_2739,N_1548,N_1219);
xnor U2740 (N_2740,N_1618,N_1408);
nand U2741 (N_2741,N_1097,N_1765);
nand U2742 (N_2742,N_1253,N_1882);
xor U2743 (N_2743,N_1569,N_1257);
nand U2744 (N_2744,N_1920,N_1796);
and U2745 (N_2745,N_1205,N_1501);
or U2746 (N_2746,N_1171,N_1559);
or U2747 (N_2747,N_1837,N_1258);
xnor U2748 (N_2748,N_1222,N_1649);
nand U2749 (N_2749,N_1023,N_1544);
nor U2750 (N_2750,N_1850,N_1750);
xnor U2751 (N_2751,N_1602,N_1827);
and U2752 (N_2752,N_1560,N_1216);
and U2753 (N_2753,N_1256,N_1254);
and U2754 (N_2754,N_1045,N_1653);
and U2755 (N_2755,N_1680,N_1138);
and U2756 (N_2756,N_1688,N_1522);
nor U2757 (N_2757,N_1487,N_1693);
nand U2758 (N_2758,N_1279,N_1743);
nand U2759 (N_2759,N_1504,N_1933);
or U2760 (N_2760,N_1988,N_1191);
and U2761 (N_2761,N_1370,N_1188);
nand U2762 (N_2762,N_1058,N_1613);
nand U2763 (N_2763,N_1035,N_1522);
or U2764 (N_2764,N_1914,N_1561);
nor U2765 (N_2765,N_1712,N_1781);
xnor U2766 (N_2766,N_1921,N_1216);
nor U2767 (N_2767,N_1977,N_1737);
xnor U2768 (N_2768,N_1649,N_1500);
nand U2769 (N_2769,N_1957,N_1607);
xor U2770 (N_2770,N_1995,N_1804);
or U2771 (N_2771,N_1809,N_1336);
xnor U2772 (N_2772,N_1524,N_1908);
nand U2773 (N_2773,N_1979,N_1555);
and U2774 (N_2774,N_1312,N_1670);
and U2775 (N_2775,N_1766,N_1008);
xnor U2776 (N_2776,N_1728,N_1552);
and U2777 (N_2777,N_1105,N_1570);
nor U2778 (N_2778,N_1741,N_1742);
nor U2779 (N_2779,N_1388,N_1108);
nand U2780 (N_2780,N_1030,N_1741);
nor U2781 (N_2781,N_1597,N_1494);
nand U2782 (N_2782,N_1118,N_1717);
nor U2783 (N_2783,N_1562,N_1200);
or U2784 (N_2784,N_1761,N_1098);
and U2785 (N_2785,N_1201,N_1582);
nor U2786 (N_2786,N_1742,N_1540);
and U2787 (N_2787,N_1936,N_1054);
and U2788 (N_2788,N_1650,N_1838);
nor U2789 (N_2789,N_1210,N_1440);
and U2790 (N_2790,N_1165,N_1071);
nand U2791 (N_2791,N_1400,N_1248);
nor U2792 (N_2792,N_1612,N_1045);
nor U2793 (N_2793,N_1782,N_1972);
nor U2794 (N_2794,N_1957,N_1091);
nand U2795 (N_2795,N_1889,N_1127);
nand U2796 (N_2796,N_1719,N_1098);
nand U2797 (N_2797,N_1969,N_1576);
nor U2798 (N_2798,N_1227,N_1452);
xnor U2799 (N_2799,N_1747,N_1155);
nor U2800 (N_2800,N_1517,N_1841);
or U2801 (N_2801,N_1902,N_1576);
and U2802 (N_2802,N_1450,N_1453);
or U2803 (N_2803,N_1300,N_1999);
xor U2804 (N_2804,N_1499,N_1181);
and U2805 (N_2805,N_1015,N_1684);
xnor U2806 (N_2806,N_1118,N_1973);
nand U2807 (N_2807,N_1672,N_1390);
or U2808 (N_2808,N_1625,N_1203);
nor U2809 (N_2809,N_1843,N_1712);
nand U2810 (N_2810,N_1010,N_1707);
or U2811 (N_2811,N_1270,N_1427);
nor U2812 (N_2812,N_1350,N_1118);
and U2813 (N_2813,N_1124,N_1291);
or U2814 (N_2814,N_1509,N_1607);
or U2815 (N_2815,N_1437,N_1122);
or U2816 (N_2816,N_1528,N_1147);
or U2817 (N_2817,N_1071,N_1039);
or U2818 (N_2818,N_1185,N_1930);
nor U2819 (N_2819,N_1079,N_1317);
nand U2820 (N_2820,N_1031,N_1649);
or U2821 (N_2821,N_1867,N_1813);
nor U2822 (N_2822,N_1762,N_1411);
and U2823 (N_2823,N_1628,N_1555);
and U2824 (N_2824,N_1643,N_1239);
nand U2825 (N_2825,N_1690,N_1376);
nand U2826 (N_2826,N_1090,N_1247);
nor U2827 (N_2827,N_1580,N_1152);
nor U2828 (N_2828,N_1634,N_1973);
xnor U2829 (N_2829,N_1309,N_1516);
nand U2830 (N_2830,N_1183,N_1222);
and U2831 (N_2831,N_1232,N_1712);
and U2832 (N_2832,N_1422,N_1778);
and U2833 (N_2833,N_1929,N_1683);
or U2834 (N_2834,N_1050,N_1910);
or U2835 (N_2835,N_1765,N_1576);
and U2836 (N_2836,N_1228,N_1975);
nor U2837 (N_2837,N_1913,N_1992);
xor U2838 (N_2838,N_1628,N_1817);
nand U2839 (N_2839,N_1778,N_1806);
nand U2840 (N_2840,N_1929,N_1843);
xor U2841 (N_2841,N_1446,N_1580);
or U2842 (N_2842,N_1458,N_1873);
nand U2843 (N_2843,N_1699,N_1227);
xor U2844 (N_2844,N_1639,N_1960);
and U2845 (N_2845,N_1992,N_1405);
nand U2846 (N_2846,N_1424,N_1606);
and U2847 (N_2847,N_1692,N_1061);
and U2848 (N_2848,N_1604,N_1770);
or U2849 (N_2849,N_1464,N_1509);
nor U2850 (N_2850,N_1197,N_1165);
nand U2851 (N_2851,N_1143,N_1908);
nor U2852 (N_2852,N_1777,N_1601);
and U2853 (N_2853,N_1796,N_1056);
xnor U2854 (N_2854,N_1331,N_1924);
or U2855 (N_2855,N_1810,N_1976);
nand U2856 (N_2856,N_1094,N_1021);
and U2857 (N_2857,N_1387,N_1280);
nor U2858 (N_2858,N_1896,N_1458);
nand U2859 (N_2859,N_1768,N_1854);
or U2860 (N_2860,N_1234,N_1159);
xnor U2861 (N_2861,N_1569,N_1940);
nand U2862 (N_2862,N_1201,N_1877);
nand U2863 (N_2863,N_1266,N_1637);
xnor U2864 (N_2864,N_1266,N_1989);
or U2865 (N_2865,N_1466,N_1606);
nor U2866 (N_2866,N_1986,N_1622);
xor U2867 (N_2867,N_1353,N_1582);
nor U2868 (N_2868,N_1992,N_1997);
nor U2869 (N_2869,N_1984,N_1398);
and U2870 (N_2870,N_1481,N_1921);
nand U2871 (N_2871,N_1060,N_1565);
nand U2872 (N_2872,N_1487,N_1930);
and U2873 (N_2873,N_1969,N_1660);
or U2874 (N_2874,N_1389,N_1927);
and U2875 (N_2875,N_1442,N_1832);
xnor U2876 (N_2876,N_1783,N_1365);
or U2877 (N_2877,N_1057,N_1028);
or U2878 (N_2878,N_1581,N_1386);
and U2879 (N_2879,N_1231,N_1391);
nand U2880 (N_2880,N_1738,N_1146);
or U2881 (N_2881,N_1839,N_1010);
or U2882 (N_2882,N_1768,N_1772);
or U2883 (N_2883,N_1995,N_1674);
nor U2884 (N_2884,N_1017,N_1051);
nand U2885 (N_2885,N_1841,N_1206);
or U2886 (N_2886,N_1345,N_1284);
nand U2887 (N_2887,N_1568,N_1441);
xnor U2888 (N_2888,N_1686,N_1189);
and U2889 (N_2889,N_1834,N_1440);
or U2890 (N_2890,N_1234,N_1734);
nor U2891 (N_2891,N_1927,N_1391);
nand U2892 (N_2892,N_1637,N_1848);
nand U2893 (N_2893,N_1523,N_1100);
and U2894 (N_2894,N_1303,N_1175);
and U2895 (N_2895,N_1379,N_1739);
or U2896 (N_2896,N_1332,N_1673);
nand U2897 (N_2897,N_1667,N_1768);
xnor U2898 (N_2898,N_1311,N_1796);
xor U2899 (N_2899,N_1707,N_1786);
nand U2900 (N_2900,N_1428,N_1003);
xnor U2901 (N_2901,N_1633,N_1938);
or U2902 (N_2902,N_1494,N_1128);
nor U2903 (N_2903,N_1229,N_1678);
and U2904 (N_2904,N_1765,N_1251);
xor U2905 (N_2905,N_1362,N_1323);
or U2906 (N_2906,N_1209,N_1274);
nand U2907 (N_2907,N_1140,N_1110);
and U2908 (N_2908,N_1168,N_1407);
and U2909 (N_2909,N_1024,N_1032);
nand U2910 (N_2910,N_1670,N_1378);
nand U2911 (N_2911,N_1009,N_1676);
and U2912 (N_2912,N_1144,N_1640);
nor U2913 (N_2913,N_1090,N_1922);
and U2914 (N_2914,N_1400,N_1423);
or U2915 (N_2915,N_1680,N_1980);
and U2916 (N_2916,N_1566,N_1763);
nor U2917 (N_2917,N_1934,N_1114);
nor U2918 (N_2918,N_1390,N_1831);
and U2919 (N_2919,N_1211,N_1286);
and U2920 (N_2920,N_1017,N_1090);
nand U2921 (N_2921,N_1705,N_1727);
and U2922 (N_2922,N_1500,N_1547);
xor U2923 (N_2923,N_1093,N_1349);
and U2924 (N_2924,N_1039,N_1365);
nand U2925 (N_2925,N_1600,N_1974);
nand U2926 (N_2926,N_1734,N_1116);
and U2927 (N_2927,N_1660,N_1542);
and U2928 (N_2928,N_1717,N_1842);
or U2929 (N_2929,N_1256,N_1094);
nor U2930 (N_2930,N_1760,N_1228);
or U2931 (N_2931,N_1800,N_1949);
or U2932 (N_2932,N_1129,N_1518);
nor U2933 (N_2933,N_1563,N_1501);
nand U2934 (N_2934,N_1978,N_1625);
or U2935 (N_2935,N_1908,N_1972);
and U2936 (N_2936,N_1401,N_1850);
xnor U2937 (N_2937,N_1301,N_1760);
and U2938 (N_2938,N_1528,N_1141);
nor U2939 (N_2939,N_1650,N_1613);
or U2940 (N_2940,N_1012,N_1988);
or U2941 (N_2941,N_1820,N_1172);
and U2942 (N_2942,N_1204,N_1976);
nor U2943 (N_2943,N_1881,N_1776);
xnor U2944 (N_2944,N_1664,N_1507);
or U2945 (N_2945,N_1068,N_1503);
and U2946 (N_2946,N_1372,N_1448);
nor U2947 (N_2947,N_1640,N_1089);
nand U2948 (N_2948,N_1939,N_1036);
xor U2949 (N_2949,N_1830,N_1167);
or U2950 (N_2950,N_1984,N_1404);
xor U2951 (N_2951,N_1491,N_1395);
and U2952 (N_2952,N_1834,N_1357);
or U2953 (N_2953,N_1179,N_1064);
or U2954 (N_2954,N_1742,N_1353);
and U2955 (N_2955,N_1648,N_1382);
nor U2956 (N_2956,N_1833,N_1236);
nand U2957 (N_2957,N_1256,N_1013);
or U2958 (N_2958,N_1889,N_1459);
and U2959 (N_2959,N_1490,N_1949);
and U2960 (N_2960,N_1265,N_1098);
and U2961 (N_2961,N_1407,N_1722);
or U2962 (N_2962,N_1870,N_1227);
nand U2963 (N_2963,N_1786,N_1803);
and U2964 (N_2964,N_1324,N_1411);
or U2965 (N_2965,N_1213,N_1625);
and U2966 (N_2966,N_1196,N_1036);
and U2967 (N_2967,N_1549,N_1307);
nand U2968 (N_2968,N_1229,N_1226);
or U2969 (N_2969,N_1980,N_1814);
nor U2970 (N_2970,N_1608,N_1311);
xnor U2971 (N_2971,N_1520,N_1788);
or U2972 (N_2972,N_1182,N_1963);
nor U2973 (N_2973,N_1377,N_1465);
and U2974 (N_2974,N_1297,N_1681);
or U2975 (N_2975,N_1144,N_1658);
nor U2976 (N_2976,N_1168,N_1934);
nand U2977 (N_2977,N_1022,N_1120);
or U2978 (N_2978,N_1065,N_1252);
or U2979 (N_2979,N_1460,N_1392);
xor U2980 (N_2980,N_1635,N_1723);
nor U2981 (N_2981,N_1811,N_1616);
nor U2982 (N_2982,N_1293,N_1118);
nand U2983 (N_2983,N_1593,N_1414);
or U2984 (N_2984,N_1718,N_1270);
nor U2985 (N_2985,N_1472,N_1835);
or U2986 (N_2986,N_1909,N_1573);
nor U2987 (N_2987,N_1064,N_1863);
and U2988 (N_2988,N_1392,N_1913);
and U2989 (N_2989,N_1904,N_1770);
or U2990 (N_2990,N_1861,N_1088);
or U2991 (N_2991,N_1719,N_1435);
nor U2992 (N_2992,N_1492,N_1039);
or U2993 (N_2993,N_1623,N_1269);
and U2994 (N_2994,N_1622,N_1614);
or U2995 (N_2995,N_1941,N_1314);
and U2996 (N_2996,N_1214,N_1059);
or U2997 (N_2997,N_1645,N_1899);
nor U2998 (N_2998,N_1042,N_1179);
or U2999 (N_2999,N_1592,N_1922);
nor U3000 (N_3000,N_2935,N_2835);
xor U3001 (N_3001,N_2489,N_2267);
or U3002 (N_3002,N_2378,N_2506);
nand U3003 (N_3003,N_2830,N_2241);
nand U3004 (N_3004,N_2049,N_2588);
nor U3005 (N_3005,N_2953,N_2023);
nand U3006 (N_3006,N_2372,N_2688);
and U3007 (N_3007,N_2577,N_2018);
and U3008 (N_3008,N_2030,N_2594);
and U3009 (N_3009,N_2986,N_2949);
or U3010 (N_3010,N_2075,N_2041);
or U3011 (N_3011,N_2676,N_2723);
and U3012 (N_3012,N_2832,N_2358);
and U3013 (N_3013,N_2786,N_2463);
xor U3014 (N_3014,N_2735,N_2653);
and U3015 (N_3015,N_2199,N_2509);
nand U3016 (N_3016,N_2504,N_2557);
nand U3017 (N_3017,N_2122,N_2687);
or U3018 (N_3018,N_2206,N_2966);
nand U3019 (N_3019,N_2955,N_2065);
or U3020 (N_3020,N_2188,N_2814);
and U3021 (N_3021,N_2348,N_2231);
or U3022 (N_3022,N_2565,N_2598);
nor U3023 (N_3023,N_2856,N_2502);
nand U3024 (N_3024,N_2131,N_2712);
nor U3025 (N_3025,N_2535,N_2649);
and U3026 (N_3026,N_2238,N_2984);
nor U3027 (N_3027,N_2548,N_2683);
nor U3028 (N_3028,N_2024,N_2938);
or U3029 (N_3029,N_2056,N_2756);
and U3030 (N_3030,N_2335,N_2518);
nor U3031 (N_3031,N_2957,N_2774);
nand U3032 (N_3032,N_2717,N_2446);
nor U3033 (N_3033,N_2132,N_2442);
and U3034 (N_3034,N_2225,N_2083);
nand U3035 (N_3035,N_2314,N_2211);
nand U3036 (N_3036,N_2531,N_2483);
and U3037 (N_3037,N_2675,N_2583);
and U3038 (N_3038,N_2136,N_2316);
nor U3039 (N_3039,N_2793,N_2346);
nor U3040 (N_3040,N_2930,N_2118);
xnor U3041 (N_3041,N_2232,N_2001);
nand U3042 (N_3042,N_2377,N_2678);
or U3043 (N_3043,N_2362,N_2396);
nor U3044 (N_3044,N_2566,N_2494);
nand U3045 (N_3045,N_2264,N_2529);
and U3046 (N_3046,N_2920,N_2948);
nand U3047 (N_3047,N_2845,N_2226);
nand U3048 (N_3048,N_2542,N_2342);
xnor U3049 (N_3049,N_2848,N_2445);
nor U3050 (N_3050,N_2960,N_2080);
nand U3051 (N_3051,N_2787,N_2640);
and U3052 (N_3052,N_2855,N_2724);
and U3053 (N_3053,N_2886,N_2981);
nand U3054 (N_3054,N_2230,N_2792);
xnor U3055 (N_3055,N_2561,N_2987);
nor U3056 (N_3056,N_2631,N_2769);
nand U3057 (N_3057,N_2618,N_2757);
xnor U3058 (N_3058,N_2659,N_2991);
and U3059 (N_3059,N_2105,N_2842);
and U3060 (N_3060,N_2242,N_2759);
nor U3061 (N_3061,N_2027,N_2785);
or U3062 (N_3062,N_2202,N_2309);
and U3063 (N_3063,N_2375,N_2718);
nor U3064 (N_3064,N_2976,N_2526);
nand U3065 (N_3065,N_2809,N_2498);
nand U3066 (N_3066,N_2743,N_2534);
nand U3067 (N_3067,N_2682,N_2628);
nor U3068 (N_3068,N_2604,N_2720);
nor U3069 (N_3069,N_2304,N_2197);
nor U3070 (N_3070,N_2635,N_2175);
nand U3071 (N_3071,N_2081,N_2591);
nor U3072 (N_3072,N_2694,N_2416);
and U3073 (N_3073,N_2982,N_2258);
nor U3074 (N_3074,N_2484,N_2662);
or U3075 (N_3075,N_2877,N_2725);
nor U3076 (N_3076,N_2052,N_2731);
or U3077 (N_3077,N_2990,N_2137);
xnor U3078 (N_3078,N_2871,N_2183);
nor U3079 (N_3079,N_2825,N_2904);
nand U3080 (N_3080,N_2589,N_2352);
or U3081 (N_3081,N_2611,N_2807);
nand U3082 (N_3082,N_2946,N_2019);
xor U3083 (N_3083,N_2317,N_2324);
nand U3084 (N_3084,N_2382,N_2089);
xnor U3085 (N_3085,N_2550,N_2087);
or U3086 (N_3086,N_2745,N_2897);
nand U3087 (N_3087,N_2562,N_2360);
nor U3088 (N_3088,N_2798,N_2411);
and U3089 (N_3089,N_2189,N_2652);
and U3090 (N_3090,N_2564,N_2826);
nand U3091 (N_3091,N_2275,N_2100);
nand U3092 (N_3092,N_2071,N_2207);
xnor U3093 (N_3093,N_2738,N_2289);
nand U3094 (N_3094,N_2022,N_2468);
nand U3095 (N_3095,N_2859,N_2808);
and U3096 (N_3096,N_2302,N_2501);
and U3097 (N_3097,N_2008,N_2811);
nand U3098 (N_3098,N_2334,N_2488);
nand U3099 (N_3099,N_2657,N_2002);
nand U3100 (N_3100,N_2954,N_2777);
and U3101 (N_3101,N_2580,N_2124);
xor U3102 (N_3102,N_2250,N_2166);
and U3103 (N_3103,N_2702,N_2729);
and U3104 (N_3104,N_2394,N_2726);
or U3105 (N_3105,N_2854,N_2074);
nor U3106 (N_3106,N_2921,N_2244);
or U3107 (N_3107,N_2940,N_2069);
or U3108 (N_3108,N_2029,N_2595);
nand U3109 (N_3109,N_2721,N_2764);
nor U3110 (N_3110,N_2407,N_2666);
or U3111 (N_3111,N_2812,N_2670);
nand U3112 (N_3112,N_2767,N_2697);
or U3113 (N_3113,N_2109,N_2404);
and U3114 (N_3114,N_2704,N_2647);
and U3115 (N_3115,N_2963,N_2097);
xor U3116 (N_3116,N_2354,N_2055);
and U3117 (N_3117,N_2999,N_2444);
and U3118 (N_3118,N_2406,N_2117);
or U3119 (N_3119,N_2418,N_2283);
nor U3120 (N_3120,N_2545,N_2454);
and U3121 (N_3121,N_2385,N_2297);
nand U3122 (N_3122,N_2715,N_2210);
nand U3123 (N_3123,N_2381,N_2365);
nor U3124 (N_3124,N_2186,N_2923);
nand U3125 (N_3125,N_2867,N_2600);
and U3126 (N_3126,N_2651,N_2200);
nor U3127 (N_3127,N_2632,N_2369);
or U3128 (N_3128,N_2373,N_2751);
and U3129 (N_3129,N_2839,N_2638);
and U3130 (N_3130,N_2491,N_2338);
or U3131 (N_3131,N_2750,N_2451);
or U3132 (N_3132,N_2789,N_2235);
nand U3133 (N_3133,N_2332,N_2343);
or U3134 (N_3134,N_2891,N_2581);
or U3135 (N_3135,N_2644,N_2270);
or U3136 (N_3136,N_2695,N_2155);
and U3137 (N_3137,N_2943,N_2037);
nor U3138 (N_3138,N_2925,N_2661);
nand U3139 (N_3139,N_2858,N_2655);
nand U3140 (N_3140,N_2587,N_2179);
or U3141 (N_3141,N_2349,N_2933);
xor U3142 (N_3142,N_2433,N_2528);
nor U3143 (N_3143,N_2795,N_2350);
or U3144 (N_3144,N_2079,N_2778);
nand U3145 (N_3145,N_2578,N_2203);
nand U3146 (N_3146,N_2585,N_2298);
and U3147 (N_3147,N_2120,N_2601);
and U3148 (N_3148,N_2469,N_2552);
and U3149 (N_3149,N_2668,N_2490);
nor U3150 (N_3150,N_2328,N_2625);
nand U3151 (N_3151,N_2749,N_2277);
or U3152 (N_3152,N_2914,N_2493);
and U3153 (N_3153,N_2453,N_2850);
nor U3154 (N_3154,N_2614,N_2586);
nand U3155 (N_3155,N_2000,N_2234);
nor U3156 (N_3156,N_2172,N_2779);
xor U3157 (N_3157,N_2734,N_2046);
nor U3158 (N_3158,N_2541,N_2144);
or U3159 (N_3159,N_2971,N_2783);
nor U3160 (N_3160,N_2866,N_2692);
nor U3161 (N_3161,N_2916,N_2156);
and U3162 (N_3162,N_2123,N_2841);
and U3163 (N_3163,N_2829,N_2962);
nand U3164 (N_3164,N_2579,N_2428);
or U3165 (N_3165,N_2152,N_2634);
nand U3166 (N_3166,N_2608,N_2711);
nor U3167 (N_3167,N_2260,N_2573);
or U3168 (N_3168,N_2937,N_2708);
or U3169 (N_3169,N_2879,N_2395);
nor U3170 (N_3170,N_2673,N_2222);
xnor U3171 (N_3171,N_2843,N_2928);
nor U3172 (N_3172,N_2791,N_2758);
nor U3173 (N_3173,N_2319,N_2048);
nand U3174 (N_3174,N_2171,N_2831);
nor U3175 (N_3175,N_2414,N_2520);
nand U3176 (N_3176,N_2788,N_2538);
and U3177 (N_3177,N_2945,N_2471);
or U3178 (N_3178,N_2582,N_2015);
or U3179 (N_3179,N_2801,N_2714);
nand U3180 (N_3180,N_2180,N_2380);
nand U3181 (N_3181,N_2941,N_2950);
or U3182 (N_3182,N_2840,N_2153);
nand U3183 (N_3183,N_2178,N_2527);
nand U3184 (N_3184,N_2684,N_2457);
xnor U3185 (N_3185,N_2931,N_2429);
or U3186 (N_3186,N_2280,N_2393);
nor U3187 (N_3187,N_2784,N_2399);
xor U3188 (N_3188,N_2020,N_2384);
and U3189 (N_3189,N_2221,N_2663);
nand U3190 (N_3190,N_2392,N_2569);
or U3191 (N_3191,N_2803,N_2077);
nor U3192 (N_3192,N_2851,N_2370);
nor U3193 (N_3193,N_2567,N_2146);
nor U3194 (N_3194,N_2664,N_2432);
and U3195 (N_3195,N_2730,N_2129);
nor U3196 (N_3196,N_2965,N_2042);
xor U3197 (N_3197,N_2351,N_2093);
nor U3198 (N_3198,N_2255,N_2145);
or U3199 (N_3199,N_2101,N_2290);
nor U3200 (N_3200,N_2887,N_2278);
xor U3201 (N_3201,N_2417,N_2810);
or U3202 (N_3202,N_2727,N_2243);
nor U3203 (N_3203,N_2383,N_2165);
nor U3204 (N_3204,N_2820,N_2936);
and U3205 (N_3205,N_2882,N_2677);
and U3206 (N_3206,N_2794,N_2536);
nor U3207 (N_3207,N_2031,N_2617);
nor U3208 (N_3208,N_2464,N_2733);
or U3209 (N_3209,N_2053,N_2599);
nor U3210 (N_3210,N_2007,N_2613);
and U3211 (N_3211,N_2603,N_2696);
and U3212 (N_3212,N_2969,N_2888);
nor U3213 (N_3213,N_2766,N_2403);
nor U3214 (N_3214,N_2044,N_2646);
nor U3215 (N_3215,N_2782,N_2308);
xor U3216 (N_3216,N_2558,N_2274);
nor U3217 (N_3217,N_2112,N_2198);
xnor U3218 (N_3218,N_2689,N_2227);
or U3219 (N_3219,N_2742,N_2555);
or U3220 (N_3220,N_2134,N_2424);
or U3221 (N_3221,N_2514,N_2543);
and U3222 (N_3222,N_2674,N_2422);
and U3223 (N_3223,N_2896,N_2823);
or U3224 (N_3224,N_2205,N_2259);
or U3225 (N_3225,N_2447,N_2014);
xnor U3226 (N_3226,N_2420,N_2374);
and U3227 (N_3227,N_2271,N_2961);
nand U3228 (N_3228,N_2300,N_2237);
nor U3229 (N_3229,N_2698,N_2460);
nand U3230 (N_3230,N_2623,N_2461);
and U3231 (N_3231,N_2149,N_2884);
and U3232 (N_3232,N_2575,N_2775);
nor U3233 (N_3233,N_2465,N_2110);
and U3234 (N_3234,N_2063,N_2699);
nor U3235 (N_3235,N_2761,N_2844);
nor U3236 (N_3236,N_2253,N_2160);
nand U3237 (N_3237,N_2173,N_2728);
nand U3238 (N_3238,N_2540,N_2201);
nor U3239 (N_3239,N_2363,N_2658);
nand U3240 (N_3240,N_2492,N_2066);
xnor U3241 (N_3241,N_2138,N_2285);
nor U3242 (N_3242,N_2802,N_2609);
or U3243 (N_3243,N_2551,N_2980);
xor U3244 (N_3244,N_2997,N_2248);
xnor U3245 (N_3245,N_2905,N_2010);
nor U3246 (N_3246,N_2257,N_2003);
or U3247 (N_3247,N_2058,N_2240);
or U3248 (N_3248,N_2455,N_2681);
nand U3249 (N_3249,N_2246,N_2184);
or U3250 (N_3250,N_2032,N_2906);
nand U3251 (N_3251,N_2036,N_2108);
or U3252 (N_3252,N_2524,N_2357);
nand U3253 (N_3253,N_2894,N_2705);
nand U3254 (N_3254,N_2747,N_2443);
or U3255 (N_3255,N_2322,N_2883);
or U3256 (N_3256,N_2716,N_2435);
or U3257 (N_3257,N_2922,N_2306);
nor U3258 (N_3258,N_2553,N_2988);
nand U3259 (N_3259,N_2017,N_2115);
and U3260 (N_3260,N_2050,N_2310);
and U3261 (N_3261,N_2596,N_2126);
nor U3262 (N_3262,N_2161,N_2368);
and U3263 (N_3263,N_2560,N_2009);
or U3264 (N_3264,N_2078,N_2141);
nand U3265 (N_3265,N_2092,N_2806);
and U3266 (N_3266,N_2430,N_2286);
or U3267 (N_3267,N_2630,N_2437);
nor U3268 (N_3268,N_2336,N_2497);
nor U3269 (N_3269,N_2474,N_2685);
nor U3270 (N_3270,N_2864,N_2292);
nor U3271 (N_3271,N_2313,N_2983);
nor U3272 (N_3272,N_2568,N_2770);
and U3273 (N_3273,N_2939,N_2367);
nand U3274 (N_3274,N_2719,N_2318);
and U3275 (N_3275,N_2265,N_2084);
or U3276 (N_3276,N_2236,N_2846);
or U3277 (N_3277,N_2507,N_2998);
nor U3278 (N_3278,N_2194,N_2584);
nand U3279 (N_3279,N_2376,N_2174);
nand U3280 (N_3280,N_2499,N_2755);
or U3281 (N_3281,N_2626,N_2865);
nand U3282 (N_3282,N_2772,N_2261);
nor U3283 (N_3283,N_2401,N_2296);
and U3284 (N_3284,N_2590,N_2450);
nand U3285 (N_3285,N_2910,N_2642);
or U3286 (N_3286,N_2409,N_2934);
or U3287 (N_3287,N_2827,N_2072);
and U3288 (N_3288,N_2157,N_2517);
or U3289 (N_3289,N_2763,N_2091);
or U3290 (N_3290,N_2899,N_2119);
or U3291 (N_3291,N_2090,N_2660);
nand U3292 (N_3292,N_2216,N_2881);
nor U3293 (N_3293,N_2480,N_2907);
nand U3294 (N_3294,N_2639,N_2070);
or U3295 (N_3295,N_2819,N_2012);
and U3296 (N_3296,N_2154,N_2113);
and U3297 (N_3297,N_2752,N_2853);
or U3298 (N_3298,N_2177,N_2505);
nand U3299 (N_3299,N_2426,N_2958);
xnor U3300 (N_3300,N_2654,N_2870);
and U3301 (N_3301,N_2006,N_2592);
nand U3302 (N_3302,N_2780,N_2073);
and U3303 (N_3303,N_2797,N_2163);
xor U3304 (N_3304,N_2620,N_2389);
nand U3305 (N_3305,N_2047,N_2790);
or U3306 (N_3306,N_2095,N_2272);
or U3307 (N_3307,N_2068,N_2765);
or U3308 (N_3308,N_2423,N_2508);
and U3309 (N_3309,N_2722,N_2732);
nor U3310 (N_3310,N_2817,N_2345);
or U3311 (N_3311,N_2315,N_2521);
nor U3312 (N_3312,N_2397,N_2574);
and U3313 (N_3313,N_2834,N_2610);
nand U3314 (N_3314,N_2919,N_2546);
nand U3315 (N_3315,N_2467,N_2776);
nor U3316 (N_3316,N_2691,N_2636);
nor U3317 (N_3317,N_2762,N_2974);
nor U3318 (N_3318,N_2927,N_2294);
nor U3319 (N_3319,N_2158,N_2218);
and U3320 (N_3320,N_2539,N_2873);
nor U3321 (N_3321,N_2857,N_2475);
nand U3322 (N_3322,N_2929,N_2185);
nand U3323 (N_3323,N_2771,N_2256);
or U3324 (N_3324,N_2208,N_2192);
and U3325 (N_3325,N_2355,N_2513);
nor U3326 (N_3326,N_2693,N_2515);
xor U3327 (N_3327,N_2667,N_2325);
nor U3328 (N_3328,N_2710,N_2898);
nor U3329 (N_3329,N_2287,N_2059);
or U3330 (N_3330,N_2151,N_2804);
and U3331 (N_3331,N_2915,N_2076);
nand U3332 (N_3332,N_2458,N_2597);
or U3333 (N_3333,N_2082,N_2473);
nand U3334 (N_3334,N_2605,N_2537);
and U3335 (N_3335,N_2744,N_2947);
or U3336 (N_3336,N_2341,N_2709);
or U3337 (N_3337,N_2593,N_2833);
and U3338 (N_3338,N_2602,N_2837);
or U3339 (N_3339,N_2951,N_2104);
or U3340 (N_3340,N_2099,N_2706);
nor U3341 (N_3341,N_2427,N_2500);
xnor U3342 (N_3342,N_2554,N_2908);
nand U3343 (N_3343,N_2511,N_2627);
xnor U3344 (N_3344,N_2379,N_2522);
nand U3345 (N_3345,N_2239,N_2466);
nor U3346 (N_3346,N_2330,N_2893);
nand U3347 (N_3347,N_2822,N_2438);
or U3348 (N_3348,N_2876,N_2512);
nand U3349 (N_3349,N_2690,N_2441);
or U3350 (N_3350,N_2487,N_2641);
xor U3351 (N_3351,N_2193,N_2295);
or U3352 (N_3352,N_2972,N_2622);
or U3353 (N_3353,N_2043,N_2680);
and U3354 (N_3354,N_2781,N_2995);
or U3355 (N_3355,N_2805,N_2967);
nand U3356 (N_3356,N_2813,N_2167);
nor U3357 (N_3357,N_2224,N_2563);
and U3358 (N_3358,N_2836,N_2707);
and U3359 (N_3359,N_2523,N_2901);
nand U3360 (N_3360,N_2190,N_2143);
nor U3361 (N_3361,N_2989,N_2975);
or U3362 (N_3362,N_2364,N_2195);
or U3363 (N_3363,N_2016,N_2616);
nor U3364 (N_3364,N_2312,N_2878);
or U3365 (N_3365,N_2985,N_2533);
or U3366 (N_3366,N_2924,N_2114);
nand U3367 (N_3367,N_2572,N_2085);
or U3368 (N_3368,N_2273,N_2576);
and U3369 (N_3369,N_2170,N_2233);
nand U3370 (N_3370,N_2164,N_2860);
nor U3371 (N_3371,N_2214,N_2532);
nand U3372 (N_3372,N_2040,N_2861);
and U3373 (N_3373,N_2410,N_2880);
or U3374 (N_3374,N_2062,N_2021);
or U3375 (N_3375,N_2150,N_2067);
or U3376 (N_3376,N_2900,N_2251);
or U3377 (N_3377,N_2485,N_2223);
xor U3378 (N_3378,N_2992,N_2125);
nand U3379 (N_3379,N_2182,N_2247);
or U3380 (N_3380,N_2686,N_2094);
or U3381 (N_3381,N_2400,N_2419);
or U3382 (N_3382,N_2993,N_2215);
xor U3383 (N_3383,N_2821,N_2266);
nand U3384 (N_3384,N_2107,N_2863);
nand U3385 (N_3385,N_2979,N_2061);
or U3386 (N_3386,N_2434,N_2977);
and U3387 (N_3387,N_2282,N_2390);
nor U3388 (N_3388,N_2824,N_2703);
or U3389 (N_3389,N_2026,N_2456);
nor U3390 (N_3390,N_2964,N_2387);
nor U3391 (N_3391,N_2495,N_2746);
nand U3392 (N_3392,N_2168,N_2956);
nand U3393 (N_3393,N_2909,N_2337);
nand U3394 (N_3394,N_2060,N_2952);
or U3395 (N_3395,N_2741,N_2281);
xnor U3396 (N_3396,N_2339,N_2329);
or U3397 (N_3397,N_2994,N_2229);
or U3398 (N_3398,N_2978,N_2147);
xor U3399 (N_3399,N_2912,N_2800);
or U3400 (N_3400,N_2847,N_2353);
and U3401 (N_3401,N_2519,N_2918);
nand U3402 (N_3402,N_2503,N_2347);
or U3403 (N_3403,N_2176,N_2740);
or U3404 (N_3404,N_2748,N_2181);
nor U3405 (N_3405,N_2116,N_2799);
and U3406 (N_3406,N_2739,N_2665);
nand U3407 (N_3407,N_2701,N_2525);
and U3408 (N_3408,N_2263,N_2650);
xnor U3409 (N_3409,N_2405,N_2838);
xnor U3410 (N_3410,N_2633,N_2187);
or U3411 (N_3411,N_2025,N_2556);
nor U3412 (N_3412,N_2402,N_2034);
nor U3413 (N_3413,N_2902,N_2011);
xor U3414 (N_3414,N_2874,N_2968);
xnor U3415 (N_3415,N_2340,N_2544);
or U3416 (N_3416,N_2629,N_2486);
xnor U3417 (N_3417,N_2643,N_2816);
or U3418 (N_3418,N_2398,N_2098);
nand U3419 (N_3419,N_2425,N_2760);
and U3420 (N_3420,N_2415,N_2033);
and U3421 (N_3421,N_2913,N_2452);
xor U3422 (N_3422,N_2440,N_2219);
and U3423 (N_3423,N_2249,N_2481);
nand U3424 (N_3424,N_2459,N_2293);
or U3425 (N_3425,N_2773,N_2013);
nand U3426 (N_3426,N_2288,N_2892);
nand U3427 (N_3427,N_2103,N_2291);
nor U3428 (N_3428,N_2669,N_2331);
or U3429 (N_3429,N_2619,N_2262);
xor U3430 (N_3430,N_2344,N_2096);
nand U3431 (N_3431,N_2612,N_2621);
or U3432 (N_3432,N_2818,N_2478);
nand U3433 (N_3433,N_2038,N_2510);
nor U3434 (N_3434,N_2169,N_2359);
nand U3435 (N_3435,N_2615,N_2736);
nor U3436 (N_3436,N_2162,N_2142);
and U3437 (N_3437,N_2127,N_2889);
nand U3438 (N_3438,N_2140,N_2875);
xor U3439 (N_3439,N_2196,N_2106);
nand U3440 (N_3440,N_2996,N_2039);
or U3441 (N_3441,N_2869,N_2606);
nand U3442 (N_3442,N_2371,N_2391);
nand U3443 (N_3443,N_2570,N_2645);
or U3444 (N_3444,N_2852,N_2496);
or U3445 (N_3445,N_2472,N_2333);
and U3446 (N_3446,N_2672,N_2942);
nand U3447 (N_3447,N_2326,N_2148);
and U3448 (N_3448,N_2516,N_2559);
nand U3449 (N_3449,N_2045,N_2911);
or U3450 (N_3450,N_2815,N_2932);
nor U3451 (N_3451,N_2547,N_2305);
nor U3452 (N_3452,N_2220,N_2470);
and U3453 (N_3453,N_2035,N_2530);
nor U3454 (N_3454,N_2111,N_2204);
nand U3455 (N_3455,N_2269,N_2051);
nand U3456 (N_3456,N_2482,N_2607);
nor U3457 (N_3457,N_2436,N_2386);
and U3458 (N_3458,N_2449,N_2849);
nor U3459 (N_3459,N_2477,N_2299);
nor U3460 (N_3460,N_2872,N_2121);
and U3461 (N_3461,N_2624,N_2217);
xor U3462 (N_3462,N_2890,N_2301);
nor U3463 (N_3463,N_2276,N_2476);
nand U3464 (N_3464,N_2311,N_2135);
nand U3465 (N_3465,N_2753,N_2252);
nor U3466 (N_3466,N_2057,N_2284);
nand U3467 (N_3467,N_2321,N_2959);
nand U3468 (N_3468,N_2917,N_2970);
or U3469 (N_3469,N_2412,N_2209);
xor U3470 (N_3470,N_2828,N_2439);
nand U3471 (N_3471,N_2064,N_2213);
nor U3472 (N_3472,N_2549,N_2868);
nor U3473 (N_3473,N_2462,N_2130);
or U3474 (N_3474,N_2700,N_2005);
nor U3475 (N_3475,N_2086,N_2448);
or U3476 (N_3476,N_2327,N_2656);
or U3477 (N_3477,N_2479,N_2388);
or U3478 (N_3478,N_2737,N_2307);
nor U3479 (N_3479,N_2366,N_2088);
or U3480 (N_3480,N_2926,N_2139);
or U3481 (N_3481,N_2159,N_2796);
xnor U3482 (N_3482,N_2191,N_2228);
nor U3483 (N_3483,N_2133,N_2431);
nand U3484 (N_3484,N_2754,N_2323);
or U3485 (N_3485,N_2671,N_2571);
and U3486 (N_3486,N_2356,N_2973);
or U3487 (N_3487,N_2279,N_2028);
and U3488 (N_3488,N_2768,N_2413);
nand U3489 (N_3489,N_2408,N_2054);
nand U3490 (N_3490,N_2004,N_2903);
nand U3491 (N_3491,N_2885,N_2254);
or U3492 (N_3492,N_2128,N_2895);
xor U3493 (N_3493,N_2713,N_2679);
or U3494 (N_3494,N_2421,N_2102);
nor U3495 (N_3495,N_2637,N_2320);
nand U3496 (N_3496,N_2648,N_2944);
nand U3497 (N_3497,N_2303,N_2268);
or U3498 (N_3498,N_2212,N_2361);
nor U3499 (N_3499,N_2245,N_2862);
nand U3500 (N_3500,N_2416,N_2420);
and U3501 (N_3501,N_2329,N_2081);
nor U3502 (N_3502,N_2762,N_2635);
nor U3503 (N_3503,N_2952,N_2843);
nand U3504 (N_3504,N_2335,N_2769);
and U3505 (N_3505,N_2820,N_2918);
or U3506 (N_3506,N_2735,N_2786);
nand U3507 (N_3507,N_2552,N_2908);
nand U3508 (N_3508,N_2263,N_2663);
xor U3509 (N_3509,N_2049,N_2896);
or U3510 (N_3510,N_2162,N_2669);
nor U3511 (N_3511,N_2627,N_2735);
xnor U3512 (N_3512,N_2991,N_2336);
nor U3513 (N_3513,N_2171,N_2288);
nand U3514 (N_3514,N_2299,N_2556);
or U3515 (N_3515,N_2674,N_2990);
nor U3516 (N_3516,N_2774,N_2971);
nor U3517 (N_3517,N_2261,N_2753);
or U3518 (N_3518,N_2920,N_2085);
or U3519 (N_3519,N_2095,N_2332);
or U3520 (N_3520,N_2966,N_2367);
or U3521 (N_3521,N_2274,N_2778);
and U3522 (N_3522,N_2709,N_2784);
or U3523 (N_3523,N_2720,N_2282);
and U3524 (N_3524,N_2317,N_2399);
nand U3525 (N_3525,N_2835,N_2487);
nand U3526 (N_3526,N_2425,N_2306);
nor U3527 (N_3527,N_2496,N_2601);
nand U3528 (N_3528,N_2763,N_2274);
nand U3529 (N_3529,N_2043,N_2156);
or U3530 (N_3530,N_2716,N_2941);
or U3531 (N_3531,N_2001,N_2147);
and U3532 (N_3532,N_2651,N_2725);
or U3533 (N_3533,N_2213,N_2132);
and U3534 (N_3534,N_2345,N_2686);
and U3535 (N_3535,N_2848,N_2938);
nor U3536 (N_3536,N_2744,N_2380);
nor U3537 (N_3537,N_2631,N_2217);
xor U3538 (N_3538,N_2604,N_2575);
nor U3539 (N_3539,N_2231,N_2333);
and U3540 (N_3540,N_2859,N_2102);
nor U3541 (N_3541,N_2134,N_2592);
nor U3542 (N_3542,N_2453,N_2796);
nand U3543 (N_3543,N_2473,N_2622);
nor U3544 (N_3544,N_2241,N_2431);
and U3545 (N_3545,N_2828,N_2467);
nand U3546 (N_3546,N_2685,N_2346);
and U3547 (N_3547,N_2171,N_2269);
xor U3548 (N_3548,N_2396,N_2101);
or U3549 (N_3549,N_2149,N_2992);
and U3550 (N_3550,N_2719,N_2357);
and U3551 (N_3551,N_2031,N_2634);
nor U3552 (N_3552,N_2791,N_2400);
or U3553 (N_3553,N_2109,N_2891);
nand U3554 (N_3554,N_2248,N_2788);
xor U3555 (N_3555,N_2884,N_2183);
nand U3556 (N_3556,N_2606,N_2631);
or U3557 (N_3557,N_2928,N_2471);
or U3558 (N_3558,N_2453,N_2357);
nand U3559 (N_3559,N_2585,N_2566);
and U3560 (N_3560,N_2286,N_2508);
xnor U3561 (N_3561,N_2108,N_2084);
nand U3562 (N_3562,N_2620,N_2175);
xnor U3563 (N_3563,N_2119,N_2910);
or U3564 (N_3564,N_2464,N_2986);
or U3565 (N_3565,N_2746,N_2321);
nor U3566 (N_3566,N_2410,N_2589);
nor U3567 (N_3567,N_2780,N_2734);
or U3568 (N_3568,N_2730,N_2207);
nand U3569 (N_3569,N_2863,N_2085);
or U3570 (N_3570,N_2771,N_2150);
nor U3571 (N_3571,N_2883,N_2162);
and U3572 (N_3572,N_2979,N_2226);
and U3573 (N_3573,N_2537,N_2085);
nand U3574 (N_3574,N_2757,N_2124);
xor U3575 (N_3575,N_2661,N_2060);
nand U3576 (N_3576,N_2298,N_2386);
nor U3577 (N_3577,N_2065,N_2295);
nor U3578 (N_3578,N_2382,N_2509);
nand U3579 (N_3579,N_2822,N_2416);
nand U3580 (N_3580,N_2167,N_2617);
or U3581 (N_3581,N_2188,N_2397);
and U3582 (N_3582,N_2265,N_2270);
nor U3583 (N_3583,N_2535,N_2059);
or U3584 (N_3584,N_2904,N_2222);
nor U3585 (N_3585,N_2581,N_2099);
nor U3586 (N_3586,N_2284,N_2233);
nand U3587 (N_3587,N_2010,N_2796);
and U3588 (N_3588,N_2678,N_2531);
nor U3589 (N_3589,N_2021,N_2574);
nand U3590 (N_3590,N_2816,N_2656);
xor U3591 (N_3591,N_2232,N_2023);
and U3592 (N_3592,N_2933,N_2594);
and U3593 (N_3593,N_2128,N_2595);
nand U3594 (N_3594,N_2709,N_2893);
and U3595 (N_3595,N_2791,N_2044);
nor U3596 (N_3596,N_2314,N_2250);
nand U3597 (N_3597,N_2902,N_2997);
nor U3598 (N_3598,N_2675,N_2587);
nand U3599 (N_3599,N_2528,N_2003);
nor U3600 (N_3600,N_2926,N_2619);
xor U3601 (N_3601,N_2931,N_2319);
and U3602 (N_3602,N_2586,N_2713);
and U3603 (N_3603,N_2226,N_2709);
nand U3604 (N_3604,N_2663,N_2553);
xor U3605 (N_3605,N_2755,N_2846);
and U3606 (N_3606,N_2810,N_2815);
nand U3607 (N_3607,N_2669,N_2268);
nand U3608 (N_3608,N_2863,N_2773);
and U3609 (N_3609,N_2318,N_2801);
nand U3610 (N_3610,N_2636,N_2440);
nor U3611 (N_3611,N_2276,N_2836);
nand U3612 (N_3612,N_2021,N_2837);
nor U3613 (N_3613,N_2770,N_2570);
and U3614 (N_3614,N_2034,N_2575);
nand U3615 (N_3615,N_2405,N_2380);
nand U3616 (N_3616,N_2621,N_2617);
or U3617 (N_3617,N_2575,N_2308);
nand U3618 (N_3618,N_2932,N_2035);
nand U3619 (N_3619,N_2909,N_2853);
or U3620 (N_3620,N_2887,N_2760);
nand U3621 (N_3621,N_2079,N_2168);
nand U3622 (N_3622,N_2979,N_2895);
xnor U3623 (N_3623,N_2344,N_2323);
nor U3624 (N_3624,N_2015,N_2444);
nor U3625 (N_3625,N_2083,N_2252);
and U3626 (N_3626,N_2309,N_2790);
or U3627 (N_3627,N_2731,N_2264);
nor U3628 (N_3628,N_2858,N_2450);
nand U3629 (N_3629,N_2547,N_2177);
and U3630 (N_3630,N_2176,N_2408);
nor U3631 (N_3631,N_2150,N_2032);
and U3632 (N_3632,N_2592,N_2643);
nor U3633 (N_3633,N_2362,N_2426);
or U3634 (N_3634,N_2025,N_2439);
or U3635 (N_3635,N_2384,N_2667);
and U3636 (N_3636,N_2917,N_2778);
and U3637 (N_3637,N_2992,N_2918);
nor U3638 (N_3638,N_2332,N_2553);
nor U3639 (N_3639,N_2245,N_2728);
and U3640 (N_3640,N_2729,N_2811);
or U3641 (N_3641,N_2939,N_2275);
nor U3642 (N_3642,N_2799,N_2047);
nand U3643 (N_3643,N_2466,N_2337);
or U3644 (N_3644,N_2808,N_2710);
nand U3645 (N_3645,N_2626,N_2967);
nor U3646 (N_3646,N_2169,N_2051);
and U3647 (N_3647,N_2788,N_2661);
or U3648 (N_3648,N_2139,N_2719);
nor U3649 (N_3649,N_2782,N_2241);
nand U3650 (N_3650,N_2205,N_2089);
and U3651 (N_3651,N_2594,N_2379);
or U3652 (N_3652,N_2799,N_2844);
nand U3653 (N_3653,N_2262,N_2716);
or U3654 (N_3654,N_2082,N_2185);
or U3655 (N_3655,N_2287,N_2261);
nand U3656 (N_3656,N_2341,N_2951);
xor U3657 (N_3657,N_2379,N_2832);
nand U3658 (N_3658,N_2728,N_2985);
nor U3659 (N_3659,N_2395,N_2996);
and U3660 (N_3660,N_2472,N_2679);
nand U3661 (N_3661,N_2682,N_2315);
xnor U3662 (N_3662,N_2140,N_2769);
nand U3663 (N_3663,N_2357,N_2598);
nor U3664 (N_3664,N_2392,N_2208);
nand U3665 (N_3665,N_2028,N_2257);
nor U3666 (N_3666,N_2048,N_2306);
nand U3667 (N_3667,N_2601,N_2924);
and U3668 (N_3668,N_2305,N_2176);
and U3669 (N_3669,N_2630,N_2663);
nand U3670 (N_3670,N_2020,N_2802);
nand U3671 (N_3671,N_2947,N_2856);
nand U3672 (N_3672,N_2141,N_2083);
or U3673 (N_3673,N_2329,N_2303);
and U3674 (N_3674,N_2868,N_2809);
xor U3675 (N_3675,N_2313,N_2551);
nor U3676 (N_3676,N_2421,N_2137);
or U3677 (N_3677,N_2464,N_2517);
nand U3678 (N_3678,N_2271,N_2084);
nand U3679 (N_3679,N_2337,N_2239);
and U3680 (N_3680,N_2079,N_2995);
or U3681 (N_3681,N_2070,N_2486);
nand U3682 (N_3682,N_2546,N_2803);
or U3683 (N_3683,N_2195,N_2148);
nor U3684 (N_3684,N_2636,N_2293);
nor U3685 (N_3685,N_2799,N_2342);
nand U3686 (N_3686,N_2043,N_2635);
nand U3687 (N_3687,N_2452,N_2737);
or U3688 (N_3688,N_2699,N_2466);
nand U3689 (N_3689,N_2844,N_2020);
nor U3690 (N_3690,N_2972,N_2067);
and U3691 (N_3691,N_2193,N_2220);
and U3692 (N_3692,N_2727,N_2849);
xor U3693 (N_3693,N_2244,N_2594);
xnor U3694 (N_3694,N_2848,N_2013);
and U3695 (N_3695,N_2493,N_2255);
or U3696 (N_3696,N_2605,N_2999);
or U3697 (N_3697,N_2029,N_2448);
xor U3698 (N_3698,N_2000,N_2941);
and U3699 (N_3699,N_2824,N_2346);
or U3700 (N_3700,N_2595,N_2752);
xor U3701 (N_3701,N_2709,N_2509);
and U3702 (N_3702,N_2068,N_2594);
and U3703 (N_3703,N_2094,N_2804);
or U3704 (N_3704,N_2636,N_2816);
nor U3705 (N_3705,N_2289,N_2621);
and U3706 (N_3706,N_2126,N_2531);
nand U3707 (N_3707,N_2934,N_2303);
nand U3708 (N_3708,N_2350,N_2520);
and U3709 (N_3709,N_2242,N_2386);
and U3710 (N_3710,N_2248,N_2032);
xnor U3711 (N_3711,N_2973,N_2274);
or U3712 (N_3712,N_2412,N_2837);
nand U3713 (N_3713,N_2806,N_2159);
and U3714 (N_3714,N_2802,N_2176);
nand U3715 (N_3715,N_2400,N_2090);
or U3716 (N_3716,N_2516,N_2090);
nand U3717 (N_3717,N_2565,N_2002);
or U3718 (N_3718,N_2162,N_2258);
and U3719 (N_3719,N_2273,N_2424);
and U3720 (N_3720,N_2664,N_2746);
nor U3721 (N_3721,N_2611,N_2853);
xnor U3722 (N_3722,N_2365,N_2531);
or U3723 (N_3723,N_2946,N_2415);
or U3724 (N_3724,N_2031,N_2274);
and U3725 (N_3725,N_2221,N_2905);
xnor U3726 (N_3726,N_2578,N_2573);
or U3727 (N_3727,N_2470,N_2459);
or U3728 (N_3728,N_2722,N_2829);
nor U3729 (N_3729,N_2692,N_2468);
nand U3730 (N_3730,N_2824,N_2684);
nand U3731 (N_3731,N_2260,N_2869);
nand U3732 (N_3732,N_2247,N_2463);
nor U3733 (N_3733,N_2086,N_2270);
nand U3734 (N_3734,N_2387,N_2970);
and U3735 (N_3735,N_2475,N_2726);
nor U3736 (N_3736,N_2641,N_2600);
and U3737 (N_3737,N_2618,N_2073);
nor U3738 (N_3738,N_2360,N_2705);
nor U3739 (N_3739,N_2674,N_2068);
or U3740 (N_3740,N_2364,N_2584);
and U3741 (N_3741,N_2668,N_2665);
xor U3742 (N_3742,N_2599,N_2175);
and U3743 (N_3743,N_2247,N_2068);
nand U3744 (N_3744,N_2607,N_2015);
nor U3745 (N_3745,N_2038,N_2389);
and U3746 (N_3746,N_2722,N_2315);
and U3747 (N_3747,N_2146,N_2164);
xor U3748 (N_3748,N_2420,N_2058);
or U3749 (N_3749,N_2422,N_2453);
or U3750 (N_3750,N_2076,N_2306);
nand U3751 (N_3751,N_2944,N_2323);
and U3752 (N_3752,N_2574,N_2854);
or U3753 (N_3753,N_2584,N_2073);
nor U3754 (N_3754,N_2330,N_2363);
nand U3755 (N_3755,N_2602,N_2778);
or U3756 (N_3756,N_2540,N_2482);
nor U3757 (N_3757,N_2675,N_2340);
nand U3758 (N_3758,N_2467,N_2346);
and U3759 (N_3759,N_2680,N_2743);
nor U3760 (N_3760,N_2418,N_2765);
nor U3761 (N_3761,N_2984,N_2718);
nor U3762 (N_3762,N_2503,N_2049);
nand U3763 (N_3763,N_2999,N_2366);
and U3764 (N_3764,N_2314,N_2887);
or U3765 (N_3765,N_2678,N_2801);
and U3766 (N_3766,N_2988,N_2365);
or U3767 (N_3767,N_2093,N_2482);
or U3768 (N_3768,N_2506,N_2144);
or U3769 (N_3769,N_2104,N_2788);
or U3770 (N_3770,N_2360,N_2900);
nor U3771 (N_3771,N_2153,N_2578);
and U3772 (N_3772,N_2499,N_2066);
nor U3773 (N_3773,N_2183,N_2730);
and U3774 (N_3774,N_2521,N_2163);
and U3775 (N_3775,N_2831,N_2796);
nor U3776 (N_3776,N_2972,N_2388);
nand U3777 (N_3777,N_2707,N_2057);
or U3778 (N_3778,N_2741,N_2251);
nor U3779 (N_3779,N_2417,N_2932);
and U3780 (N_3780,N_2072,N_2257);
and U3781 (N_3781,N_2083,N_2176);
nor U3782 (N_3782,N_2955,N_2290);
or U3783 (N_3783,N_2655,N_2533);
nand U3784 (N_3784,N_2254,N_2198);
and U3785 (N_3785,N_2990,N_2898);
nand U3786 (N_3786,N_2939,N_2574);
and U3787 (N_3787,N_2361,N_2023);
xor U3788 (N_3788,N_2046,N_2408);
nor U3789 (N_3789,N_2436,N_2431);
nor U3790 (N_3790,N_2268,N_2461);
and U3791 (N_3791,N_2188,N_2702);
and U3792 (N_3792,N_2473,N_2234);
and U3793 (N_3793,N_2627,N_2161);
or U3794 (N_3794,N_2586,N_2628);
nor U3795 (N_3795,N_2685,N_2537);
and U3796 (N_3796,N_2799,N_2829);
or U3797 (N_3797,N_2315,N_2783);
nor U3798 (N_3798,N_2339,N_2411);
and U3799 (N_3799,N_2633,N_2141);
or U3800 (N_3800,N_2229,N_2702);
nand U3801 (N_3801,N_2209,N_2634);
or U3802 (N_3802,N_2631,N_2717);
nor U3803 (N_3803,N_2950,N_2045);
nor U3804 (N_3804,N_2904,N_2394);
nor U3805 (N_3805,N_2865,N_2059);
nor U3806 (N_3806,N_2343,N_2278);
and U3807 (N_3807,N_2928,N_2249);
and U3808 (N_3808,N_2825,N_2100);
xor U3809 (N_3809,N_2309,N_2466);
nor U3810 (N_3810,N_2330,N_2341);
and U3811 (N_3811,N_2834,N_2478);
nand U3812 (N_3812,N_2743,N_2915);
and U3813 (N_3813,N_2481,N_2463);
and U3814 (N_3814,N_2918,N_2151);
and U3815 (N_3815,N_2542,N_2446);
or U3816 (N_3816,N_2056,N_2551);
nor U3817 (N_3817,N_2149,N_2875);
and U3818 (N_3818,N_2662,N_2807);
or U3819 (N_3819,N_2030,N_2352);
and U3820 (N_3820,N_2866,N_2222);
xor U3821 (N_3821,N_2503,N_2229);
nor U3822 (N_3822,N_2540,N_2500);
or U3823 (N_3823,N_2958,N_2583);
and U3824 (N_3824,N_2033,N_2692);
and U3825 (N_3825,N_2952,N_2142);
or U3826 (N_3826,N_2662,N_2441);
or U3827 (N_3827,N_2646,N_2747);
or U3828 (N_3828,N_2657,N_2926);
and U3829 (N_3829,N_2277,N_2084);
and U3830 (N_3830,N_2047,N_2202);
nand U3831 (N_3831,N_2599,N_2457);
nor U3832 (N_3832,N_2608,N_2363);
and U3833 (N_3833,N_2884,N_2901);
or U3834 (N_3834,N_2944,N_2527);
nand U3835 (N_3835,N_2338,N_2272);
nor U3836 (N_3836,N_2985,N_2530);
and U3837 (N_3837,N_2987,N_2830);
nor U3838 (N_3838,N_2090,N_2569);
nor U3839 (N_3839,N_2562,N_2298);
nand U3840 (N_3840,N_2223,N_2553);
xor U3841 (N_3841,N_2802,N_2374);
xnor U3842 (N_3842,N_2388,N_2027);
nand U3843 (N_3843,N_2639,N_2850);
nor U3844 (N_3844,N_2286,N_2333);
or U3845 (N_3845,N_2971,N_2698);
nor U3846 (N_3846,N_2501,N_2933);
and U3847 (N_3847,N_2435,N_2157);
nor U3848 (N_3848,N_2107,N_2731);
or U3849 (N_3849,N_2538,N_2863);
xnor U3850 (N_3850,N_2226,N_2557);
and U3851 (N_3851,N_2014,N_2266);
nor U3852 (N_3852,N_2569,N_2888);
or U3853 (N_3853,N_2179,N_2039);
or U3854 (N_3854,N_2768,N_2175);
and U3855 (N_3855,N_2986,N_2704);
nor U3856 (N_3856,N_2446,N_2798);
and U3857 (N_3857,N_2820,N_2523);
xor U3858 (N_3858,N_2187,N_2902);
nor U3859 (N_3859,N_2320,N_2944);
or U3860 (N_3860,N_2229,N_2320);
nor U3861 (N_3861,N_2665,N_2246);
or U3862 (N_3862,N_2329,N_2109);
or U3863 (N_3863,N_2061,N_2641);
nand U3864 (N_3864,N_2027,N_2113);
or U3865 (N_3865,N_2446,N_2587);
nor U3866 (N_3866,N_2585,N_2709);
and U3867 (N_3867,N_2310,N_2711);
or U3868 (N_3868,N_2185,N_2833);
and U3869 (N_3869,N_2557,N_2752);
or U3870 (N_3870,N_2713,N_2335);
or U3871 (N_3871,N_2690,N_2008);
and U3872 (N_3872,N_2154,N_2516);
or U3873 (N_3873,N_2350,N_2524);
nor U3874 (N_3874,N_2040,N_2703);
or U3875 (N_3875,N_2021,N_2691);
nand U3876 (N_3876,N_2751,N_2616);
and U3877 (N_3877,N_2915,N_2266);
and U3878 (N_3878,N_2240,N_2973);
nand U3879 (N_3879,N_2744,N_2087);
nor U3880 (N_3880,N_2231,N_2305);
nor U3881 (N_3881,N_2616,N_2775);
or U3882 (N_3882,N_2464,N_2613);
nand U3883 (N_3883,N_2732,N_2821);
xor U3884 (N_3884,N_2165,N_2450);
or U3885 (N_3885,N_2967,N_2774);
and U3886 (N_3886,N_2973,N_2529);
nand U3887 (N_3887,N_2442,N_2194);
and U3888 (N_3888,N_2386,N_2115);
and U3889 (N_3889,N_2580,N_2715);
nor U3890 (N_3890,N_2488,N_2487);
nor U3891 (N_3891,N_2371,N_2283);
nand U3892 (N_3892,N_2564,N_2034);
and U3893 (N_3893,N_2965,N_2630);
or U3894 (N_3894,N_2024,N_2292);
and U3895 (N_3895,N_2706,N_2389);
or U3896 (N_3896,N_2707,N_2508);
nor U3897 (N_3897,N_2615,N_2866);
xor U3898 (N_3898,N_2111,N_2254);
nand U3899 (N_3899,N_2524,N_2138);
nand U3900 (N_3900,N_2789,N_2539);
nor U3901 (N_3901,N_2955,N_2698);
or U3902 (N_3902,N_2910,N_2779);
and U3903 (N_3903,N_2882,N_2447);
or U3904 (N_3904,N_2820,N_2022);
or U3905 (N_3905,N_2796,N_2627);
or U3906 (N_3906,N_2119,N_2449);
or U3907 (N_3907,N_2304,N_2119);
nand U3908 (N_3908,N_2398,N_2695);
nor U3909 (N_3909,N_2414,N_2972);
nor U3910 (N_3910,N_2706,N_2869);
nor U3911 (N_3911,N_2588,N_2465);
xor U3912 (N_3912,N_2488,N_2930);
or U3913 (N_3913,N_2292,N_2662);
nor U3914 (N_3914,N_2455,N_2655);
and U3915 (N_3915,N_2877,N_2314);
and U3916 (N_3916,N_2846,N_2899);
or U3917 (N_3917,N_2206,N_2344);
and U3918 (N_3918,N_2029,N_2582);
or U3919 (N_3919,N_2567,N_2191);
nor U3920 (N_3920,N_2073,N_2434);
nand U3921 (N_3921,N_2046,N_2761);
nor U3922 (N_3922,N_2168,N_2393);
nand U3923 (N_3923,N_2092,N_2163);
nor U3924 (N_3924,N_2599,N_2573);
nand U3925 (N_3925,N_2246,N_2666);
and U3926 (N_3926,N_2156,N_2748);
or U3927 (N_3927,N_2390,N_2549);
and U3928 (N_3928,N_2663,N_2326);
nand U3929 (N_3929,N_2497,N_2384);
nor U3930 (N_3930,N_2163,N_2218);
nor U3931 (N_3931,N_2330,N_2988);
and U3932 (N_3932,N_2890,N_2991);
and U3933 (N_3933,N_2959,N_2202);
xnor U3934 (N_3934,N_2688,N_2726);
xnor U3935 (N_3935,N_2843,N_2773);
nand U3936 (N_3936,N_2750,N_2979);
or U3937 (N_3937,N_2422,N_2765);
or U3938 (N_3938,N_2064,N_2961);
and U3939 (N_3939,N_2560,N_2573);
and U3940 (N_3940,N_2338,N_2064);
nand U3941 (N_3941,N_2634,N_2010);
or U3942 (N_3942,N_2948,N_2494);
nor U3943 (N_3943,N_2855,N_2906);
and U3944 (N_3944,N_2618,N_2279);
nor U3945 (N_3945,N_2492,N_2151);
nand U3946 (N_3946,N_2851,N_2966);
xnor U3947 (N_3947,N_2542,N_2960);
and U3948 (N_3948,N_2460,N_2439);
nor U3949 (N_3949,N_2954,N_2185);
and U3950 (N_3950,N_2999,N_2357);
nor U3951 (N_3951,N_2853,N_2554);
nand U3952 (N_3952,N_2592,N_2571);
and U3953 (N_3953,N_2360,N_2992);
or U3954 (N_3954,N_2271,N_2503);
or U3955 (N_3955,N_2260,N_2079);
nand U3956 (N_3956,N_2971,N_2654);
and U3957 (N_3957,N_2637,N_2309);
xor U3958 (N_3958,N_2726,N_2806);
nor U3959 (N_3959,N_2025,N_2931);
xor U3960 (N_3960,N_2513,N_2883);
nand U3961 (N_3961,N_2794,N_2842);
or U3962 (N_3962,N_2815,N_2887);
or U3963 (N_3963,N_2983,N_2936);
or U3964 (N_3964,N_2355,N_2606);
nand U3965 (N_3965,N_2535,N_2669);
and U3966 (N_3966,N_2485,N_2133);
nor U3967 (N_3967,N_2895,N_2122);
and U3968 (N_3968,N_2746,N_2485);
and U3969 (N_3969,N_2192,N_2500);
or U3970 (N_3970,N_2302,N_2994);
nand U3971 (N_3971,N_2427,N_2931);
xor U3972 (N_3972,N_2144,N_2589);
and U3973 (N_3973,N_2262,N_2684);
nor U3974 (N_3974,N_2237,N_2003);
nor U3975 (N_3975,N_2926,N_2233);
xor U3976 (N_3976,N_2584,N_2160);
or U3977 (N_3977,N_2791,N_2274);
xnor U3978 (N_3978,N_2172,N_2516);
nor U3979 (N_3979,N_2918,N_2430);
nor U3980 (N_3980,N_2208,N_2041);
or U3981 (N_3981,N_2035,N_2484);
nor U3982 (N_3982,N_2148,N_2791);
nor U3983 (N_3983,N_2752,N_2001);
or U3984 (N_3984,N_2320,N_2538);
xnor U3985 (N_3985,N_2398,N_2472);
nand U3986 (N_3986,N_2285,N_2379);
nor U3987 (N_3987,N_2562,N_2482);
nor U3988 (N_3988,N_2788,N_2197);
and U3989 (N_3989,N_2375,N_2732);
or U3990 (N_3990,N_2320,N_2848);
nor U3991 (N_3991,N_2904,N_2002);
xor U3992 (N_3992,N_2677,N_2177);
or U3993 (N_3993,N_2822,N_2917);
nand U3994 (N_3994,N_2484,N_2395);
or U3995 (N_3995,N_2108,N_2864);
xor U3996 (N_3996,N_2101,N_2039);
and U3997 (N_3997,N_2318,N_2531);
xnor U3998 (N_3998,N_2893,N_2856);
nand U3999 (N_3999,N_2898,N_2789);
nor U4000 (N_4000,N_3833,N_3456);
nor U4001 (N_4001,N_3662,N_3786);
nor U4002 (N_4002,N_3700,N_3371);
and U4003 (N_4003,N_3637,N_3432);
nand U4004 (N_4004,N_3244,N_3028);
xor U4005 (N_4005,N_3962,N_3723);
nor U4006 (N_4006,N_3642,N_3128);
nand U4007 (N_4007,N_3204,N_3035);
nor U4008 (N_4008,N_3799,N_3965);
nand U4009 (N_4009,N_3331,N_3695);
nor U4010 (N_4010,N_3278,N_3241);
nand U4011 (N_4011,N_3831,N_3923);
nand U4012 (N_4012,N_3918,N_3068);
nand U4013 (N_4013,N_3215,N_3102);
or U4014 (N_4014,N_3400,N_3195);
and U4015 (N_4015,N_3980,N_3552);
nor U4016 (N_4016,N_3622,N_3271);
nor U4017 (N_4017,N_3142,N_3766);
or U4018 (N_4018,N_3040,N_3222);
nand U4019 (N_4019,N_3607,N_3060);
and U4020 (N_4020,N_3237,N_3977);
and U4021 (N_4021,N_3365,N_3879);
nor U4022 (N_4022,N_3186,N_3652);
and U4023 (N_4023,N_3210,N_3517);
nand U4024 (N_4024,N_3732,N_3540);
nor U4025 (N_4025,N_3947,N_3995);
nand U4026 (N_4026,N_3105,N_3683);
nor U4027 (N_4027,N_3321,N_3903);
xnor U4028 (N_4028,N_3049,N_3409);
and U4029 (N_4029,N_3134,N_3940);
nand U4030 (N_4030,N_3182,N_3985);
or U4031 (N_4031,N_3735,N_3263);
or U4032 (N_4032,N_3260,N_3258);
and U4033 (N_4033,N_3538,N_3789);
xor U4034 (N_4034,N_3870,N_3151);
nor U4035 (N_4035,N_3959,N_3532);
nor U4036 (N_4036,N_3803,N_3248);
or U4037 (N_4037,N_3184,N_3283);
nor U4038 (N_4038,N_3467,N_3763);
or U4039 (N_4039,N_3508,N_3385);
xor U4040 (N_4040,N_3911,N_3058);
nor U4041 (N_4041,N_3307,N_3793);
or U4042 (N_4042,N_3707,N_3595);
or U4043 (N_4043,N_3692,N_3869);
nand U4044 (N_4044,N_3664,N_3447);
nor U4045 (N_4045,N_3576,N_3915);
nor U4046 (N_4046,N_3649,N_3927);
xnor U4047 (N_4047,N_3890,N_3380);
and U4048 (N_4048,N_3505,N_3840);
and U4049 (N_4049,N_3991,N_3535);
xnor U4050 (N_4050,N_3668,N_3953);
xnor U4051 (N_4051,N_3477,N_3641);
or U4052 (N_4052,N_3116,N_3451);
or U4053 (N_4053,N_3929,N_3069);
and U4054 (N_4054,N_3197,N_3312);
and U4055 (N_4055,N_3620,N_3575);
nand U4056 (N_4056,N_3476,N_3526);
nand U4057 (N_4057,N_3085,N_3234);
xnor U4058 (N_4058,N_3511,N_3292);
and U4059 (N_4059,N_3531,N_3850);
nor U4060 (N_4060,N_3804,N_3956);
nand U4061 (N_4061,N_3917,N_3338);
and U4062 (N_4062,N_3439,N_3482);
nand U4063 (N_4063,N_3568,N_3320);
and U4064 (N_4064,N_3080,N_3103);
or U4065 (N_4065,N_3277,N_3284);
or U4066 (N_4066,N_3126,N_3772);
and U4067 (N_4067,N_3893,N_3632);
nor U4068 (N_4068,N_3427,N_3486);
and U4069 (N_4069,N_3254,N_3589);
nand U4070 (N_4070,N_3809,N_3823);
and U4071 (N_4071,N_3319,N_3377);
nand U4072 (N_4072,N_3359,N_3416);
nand U4073 (N_4073,N_3480,N_3553);
nor U4074 (N_4074,N_3408,N_3557);
and U4075 (N_4075,N_3618,N_3906);
or U4076 (N_4076,N_3226,N_3188);
xor U4077 (N_4077,N_3458,N_3031);
and U4078 (N_4078,N_3998,N_3871);
nand U4079 (N_4079,N_3691,N_3086);
or U4080 (N_4080,N_3779,N_3328);
or U4081 (N_4081,N_3584,N_3073);
and U4082 (N_4082,N_3737,N_3136);
and U4083 (N_4083,N_3560,N_3370);
or U4084 (N_4084,N_3685,N_3897);
xor U4085 (N_4085,N_3717,N_3183);
nand U4086 (N_4086,N_3884,N_3079);
nor U4087 (N_4087,N_3462,N_3302);
nand U4088 (N_4088,N_3812,N_3084);
nand U4089 (N_4089,N_3951,N_3017);
nand U4090 (N_4090,N_3654,N_3094);
or U4091 (N_4091,N_3386,N_3533);
nor U4092 (N_4092,N_3898,N_3597);
nor U4093 (N_4093,N_3418,N_3381);
nor U4094 (N_4094,N_3656,N_3971);
xnor U4095 (N_4095,N_3153,N_3144);
or U4096 (N_4096,N_3600,N_3115);
and U4097 (N_4097,N_3473,N_3718);
xor U4098 (N_4098,N_3154,N_3122);
and U4099 (N_4099,N_3817,N_3521);
nor U4100 (N_4100,N_3164,N_3888);
and U4101 (N_4101,N_3537,N_3363);
nand U4102 (N_4102,N_3714,N_3438);
or U4103 (N_4103,N_3016,N_3921);
or U4104 (N_4104,N_3033,N_3748);
nand U4105 (N_4105,N_3376,N_3163);
and U4106 (N_4106,N_3420,N_3070);
and U4107 (N_4107,N_3894,N_3635);
or U4108 (N_4108,N_3670,N_3099);
and U4109 (N_4109,N_3751,N_3601);
xnor U4110 (N_4110,N_3912,N_3372);
nand U4111 (N_4111,N_3639,N_3491);
nand U4112 (N_4112,N_3324,N_3348);
and U4113 (N_4113,N_3908,N_3587);
and U4114 (N_4114,N_3463,N_3095);
or U4115 (N_4115,N_3876,N_3326);
nand U4116 (N_4116,N_3562,N_3738);
and U4117 (N_4117,N_3082,N_3332);
and U4118 (N_4118,N_3148,N_3768);
or U4119 (N_4119,N_3716,N_3863);
nor U4120 (N_4120,N_3556,N_3149);
nor U4121 (N_4121,N_3034,N_3913);
or U4122 (N_4122,N_3075,N_3228);
or U4123 (N_4123,N_3047,N_3820);
or U4124 (N_4124,N_3225,N_3452);
or U4125 (N_4125,N_3293,N_3968);
and U4126 (N_4126,N_3807,N_3954);
nand U4127 (N_4127,N_3446,N_3131);
xnor U4128 (N_4128,N_3811,N_3881);
nor U4129 (N_4129,N_3265,N_3591);
xor U4130 (N_4130,N_3443,N_3431);
and U4131 (N_4131,N_3202,N_3629);
or U4132 (N_4132,N_3794,N_3140);
nor U4133 (N_4133,N_3536,N_3887);
nand U4134 (N_4134,N_3993,N_3663);
nor U4135 (N_4135,N_3698,N_3529);
xor U4136 (N_4136,N_3203,N_3755);
nand U4137 (N_4137,N_3496,N_3773);
nand U4138 (N_4138,N_3403,N_3383);
nand U4139 (N_4139,N_3527,N_3349);
nand U4140 (N_4140,N_3395,N_3001);
and U4141 (N_4141,N_3355,N_3873);
nand U4142 (N_4142,N_3185,N_3907);
nor U4143 (N_4143,N_3752,N_3741);
or U4144 (N_4144,N_3118,N_3657);
or U4145 (N_4145,N_3350,N_3343);
or U4146 (N_4146,N_3390,N_3740);
or U4147 (N_4147,N_3147,N_3050);
or U4148 (N_4148,N_3964,N_3327);
xor U4149 (N_4149,N_3586,N_3747);
or U4150 (N_4150,N_3235,N_3734);
nor U4151 (N_4151,N_3242,N_3819);
nand U4152 (N_4152,N_3139,N_3112);
nand U4153 (N_4153,N_3445,N_3711);
and U4154 (N_4154,N_3598,N_3757);
or U4155 (N_4155,N_3571,N_3979);
nor U4156 (N_4156,N_3989,N_3880);
and U4157 (N_4157,N_3674,N_3301);
and U4158 (N_4158,N_3628,N_3141);
nor U4159 (N_4159,N_3750,N_3217);
or U4160 (N_4160,N_3563,N_3208);
and U4161 (N_4161,N_3676,N_3725);
or U4162 (N_4162,N_3659,N_3855);
or U4163 (N_4163,N_3178,N_3868);
nor U4164 (N_4164,N_3209,N_3398);
nor U4165 (N_4165,N_3981,N_3155);
or U4166 (N_4166,N_3366,N_3437);
or U4167 (N_4167,N_3514,N_3938);
nand U4168 (N_4168,N_3885,N_3191);
or U4169 (N_4169,N_3719,N_3973);
xnor U4170 (N_4170,N_3159,N_3125);
nor U4171 (N_4171,N_3479,N_3950);
nand U4172 (N_4172,N_3680,N_3667);
or U4173 (N_4173,N_3090,N_3650);
or U4174 (N_4174,N_3594,N_3269);
and U4175 (N_4175,N_3024,N_3490);
or U4176 (N_4176,N_3252,N_3986);
nand U4177 (N_4177,N_3828,N_3678);
nand U4178 (N_4178,N_3852,N_3513);
or U4179 (N_4179,N_3106,N_3032);
nand U4180 (N_4180,N_3026,N_3375);
xnor U4181 (N_4181,N_3822,N_3502);
nor U4182 (N_4182,N_3449,N_3276);
nand U4183 (N_4183,N_3459,N_3334);
nor U4184 (N_4184,N_3404,N_3193);
nor U4185 (N_4185,N_3818,N_3150);
nor U4186 (N_4186,N_3045,N_3410);
nand U4187 (N_4187,N_3158,N_3646);
or U4188 (N_4188,N_3645,N_3722);
and U4189 (N_4189,N_3081,N_3997);
nor U4190 (N_4190,N_3506,N_3984);
nor U4191 (N_4191,N_3815,N_3624);
nand U4192 (N_4192,N_3129,N_3928);
and U4193 (N_4193,N_3296,N_3264);
or U4194 (N_4194,N_3883,N_3078);
and U4195 (N_4195,N_3567,N_3961);
nand U4196 (N_4196,N_3644,N_3247);
nand U4197 (N_4197,N_3920,N_3021);
or U4198 (N_4198,N_3936,N_3742);
xnor U4199 (N_4199,N_3119,N_3097);
or U4200 (N_4200,N_3565,N_3392);
xnor U4201 (N_4201,N_3262,N_3539);
or U4202 (N_4202,N_3192,N_3616);
or U4203 (N_4203,N_3874,N_3466);
or U4204 (N_4204,N_3207,N_3056);
nor U4205 (N_4205,N_3574,N_3764);
xor U4206 (N_4206,N_3935,N_3417);
and U4207 (N_4207,N_3165,N_3945);
xor U4208 (N_4208,N_3621,N_3011);
nor U4209 (N_4209,N_3487,N_3922);
nand U4210 (N_4210,N_3858,N_3176);
nand U4211 (N_4211,N_3559,N_3914);
nand U4212 (N_4212,N_3651,N_3053);
nor U4213 (N_4213,N_3702,N_3104);
or U4214 (N_4214,N_3402,N_3608);
or U4215 (N_4215,N_3859,N_3469);
xor U4216 (N_4216,N_3713,N_3708);
nand U4217 (N_4217,N_3933,N_3937);
or U4218 (N_4218,N_3289,N_3323);
nand U4219 (N_4219,N_3522,N_3453);
nor U4220 (N_4220,N_3925,N_3109);
nand U4221 (N_4221,N_3317,N_3633);
xnor U4222 (N_4222,N_3810,N_3825);
nor U4223 (N_4223,N_3329,N_3108);
nor U4224 (N_4224,N_3232,N_3904);
or U4225 (N_4225,N_3788,N_3133);
and U4226 (N_4226,N_3123,N_3223);
nor U4227 (N_4227,N_3290,N_3579);
xnor U4228 (N_4228,N_3944,N_3093);
and U4229 (N_4229,N_3351,N_3072);
and U4230 (N_4230,N_3845,N_3967);
and U4231 (N_4231,N_3839,N_3932);
nor U4232 (N_4232,N_3166,N_3515);
xor U4233 (N_4233,N_3267,N_3975);
or U4234 (N_4234,N_3569,N_3573);
nor U4235 (N_4235,N_3780,N_3025);
or U4236 (N_4236,N_3543,N_3795);
xnor U4237 (N_4237,N_3778,N_3062);
or U4238 (N_4238,N_3239,N_3805);
or U4239 (N_4239,N_3982,N_3860);
and U4240 (N_4240,N_3541,N_3304);
xnor U4241 (N_4241,N_3394,N_3457);
nand U4242 (N_4242,N_3229,N_3160);
and U4243 (N_4243,N_3826,N_3064);
nor U4244 (N_4244,N_3096,N_3137);
or U4245 (N_4245,N_3423,N_3340);
nand U4246 (N_4246,N_3038,N_3127);
nor U4247 (N_4247,N_3948,N_3117);
nand U4248 (N_4248,N_3369,N_3291);
nand U4249 (N_4249,N_3547,N_3609);
nor U4250 (N_4250,N_3983,N_3441);
and U4251 (N_4251,N_3460,N_3444);
nand U4252 (N_4252,N_3275,N_3952);
nor U4253 (N_4253,N_3083,N_3864);
nor U4254 (N_4254,N_3548,N_3009);
and U4255 (N_4255,N_3900,N_3132);
and U4256 (N_4256,N_3684,N_3987);
or U4257 (N_4257,N_3030,N_3806);
and U4258 (N_4258,N_3114,N_3509);
nor U4259 (N_4259,N_3055,N_3824);
and U4260 (N_4260,N_3311,N_3753);
and U4261 (N_4261,N_3554,N_3798);
nor U4262 (N_4262,N_3648,N_3610);
and U4263 (N_4263,N_3528,N_3675);
xor U4264 (N_4264,N_3309,N_3617);
xor U4265 (N_4265,N_3801,N_3227);
nor U4266 (N_4266,N_3524,N_3057);
and U4267 (N_4267,N_3715,N_3054);
nor U4268 (N_4268,N_3838,N_3036);
nand U4269 (N_4269,N_3942,N_3875);
nand U4270 (N_4270,N_3401,N_3274);
or U4271 (N_4271,N_3318,N_3802);
nor U4272 (N_4272,N_3358,N_3337);
xnor U4273 (N_4273,N_3414,N_3424);
and U4274 (N_4274,N_3280,N_3672);
nor U4275 (N_4275,N_3739,N_3796);
nand U4276 (N_4276,N_3044,N_3577);
nand U4277 (N_4277,N_3145,N_3357);
and U4278 (N_4278,N_3266,N_3919);
and U4279 (N_4279,N_3306,N_3168);
nor U4280 (N_4280,N_3493,N_3976);
nand U4281 (N_4281,N_3316,N_3848);
and U4282 (N_4282,N_3010,N_3161);
or U4283 (N_4283,N_3762,N_3902);
xor U4284 (N_4284,N_3626,N_3623);
nor U4285 (N_4285,N_3924,N_3816);
nand U4286 (N_4286,N_3214,N_3857);
nand U4287 (N_4287,N_3405,N_3743);
and U4288 (N_4288,N_3240,N_3555);
nand U4289 (N_4289,N_3023,N_3604);
or U4290 (N_4290,N_3257,N_3581);
nor U4291 (N_4291,N_3978,N_3974);
and U4292 (N_4292,N_3882,N_3736);
or U4293 (N_4293,N_3504,N_3934);
or U4294 (N_4294,N_3245,N_3500);
and U4295 (N_4295,N_3250,N_3867);
or U4296 (N_4296,N_3889,N_3428);
or U4297 (N_4297,N_3483,N_3042);
nand U4298 (N_4298,N_3614,N_3322);
nor U4299 (N_4299,N_3842,N_3733);
nor U4300 (N_4300,N_3298,N_3230);
and U4301 (N_4301,N_3211,N_3957);
nor U4302 (N_4302,N_3963,N_3611);
or U4303 (N_4303,N_3249,N_3679);
nand U4304 (N_4304,N_3666,N_3696);
or U4305 (N_4305,N_3588,N_3744);
or U4306 (N_4306,N_3846,N_3220);
xor U4307 (N_4307,N_3018,N_3730);
nand U4308 (N_4308,N_3558,N_3785);
nor U4309 (N_4309,N_3782,N_3014);
and U4310 (N_4310,N_3005,N_3728);
nor U4311 (N_4311,N_3135,N_3865);
and U4312 (N_4312,N_3710,N_3749);
xor U4313 (N_4313,N_3771,N_3368);
or U4314 (N_4314,N_3305,N_3759);
nand U4315 (N_4315,N_3653,N_3100);
nor U4316 (N_4316,N_3905,N_3465);
and U4317 (N_4317,N_3325,N_3512);
nand U4318 (N_4318,N_3143,N_3157);
nor U4319 (N_4319,N_3236,N_3570);
and U4320 (N_4320,N_3724,N_3287);
or U4321 (N_4321,N_3687,N_3546);
and U4322 (N_4322,N_3854,N_3255);
xor U4323 (N_4323,N_3808,N_3448);
nand U4324 (N_4324,N_3489,N_3545);
or U4325 (N_4325,N_3146,N_3703);
nor U4326 (N_4326,N_3847,N_3167);
and U4327 (N_4327,N_3494,N_3273);
nand U4328 (N_4328,N_3039,N_3425);
and U4329 (N_4329,N_3761,N_3374);
nand U4330 (N_4330,N_3243,N_3484);
nand U4331 (N_4331,N_3549,N_3180);
or U4332 (N_4332,N_3955,N_3534);
and U4333 (N_4333,N_3216,N_3200);
and U4334 (N_4334,N_3690,N_3499);
or U4335 (N_4335,N_3397,N_3174);
nand U4336 (N_4336,N_3205,N_3530);
and U4337 (N_4337,N_3261,N_3124);
nand U4338 (N_4338,N_3943,N_3877);
nor U4339 (N_4339,N_3688,N_3442);
nand U4340 (N_4340,N_3345,N_3272);
nor U4341 (N_4341,N_3303,N_3152);
or U4342 (N_4342,N_3721,N_3636);
nor U4343 (N_4343,N_3171,N_3110);
nand U4344 (N_4344,N_3022,N_3411);
or U4345 (N_4345,N_3660,N_3781);
nand U4346 (N_4346,N_3827,N_3926);
or U4347 (N_4347,N_3189,N_3655);
xnor U4348 (N_4348,N_3065,N_3378);
or U4349 (N_4349,N_3091,N_3561);
nand U4350 (N_4350,N_3231,N_3407);
nor U4351 (N_4351,N_3516,N_3475);
or U4352 (N_4352,N_3800,N_3966);
nand U4353 (N_4353,N_3027,N_3603);
nor U4354 (N_4354,N_3294,N_3834);
and U4355 (N_4355,N_3396,N_3002);
or U4356 (N_4356,N_3288,N_3492);
and U4357 (N_4357,N_3787,N_3130);
or U4358 (N_4358,N_3916,N_3886);
nand U4359 (N_4359,N_3941,N_3472);
nor U4360 (N_4360,N_3583,N_3899);
or U4361 (N_4361,N_3760,N_3791);
nor U4362 (N_4362,N_3605,N_3455);
and U4363 (N_4363,N_3238,N_3813);
xor U4364 (N_4364,N_3003,N_3098);
nand U4365 (N_4365,N_3281,N_3783);
or U4366 (N_4366,N_3170,N_3580);
or U4367 (N_4367,N_3497,N_3221);
nor U4368 (N_4368,N_3896,N_3996);
and U4369 (N_4369,N_3784,N_3364);
nand U4370 (N_4370,N_3246,N_3849);
nand U4371 (N_4371,N_3585,N_3593);
or U4372 (N_4372,N_3615,N_3862);
or U4373 (N_4373,N_3720,N_3313);
nand U4374 (N_4374,N_3756,N_3892);
or U4375 (N_4375,N_3335,N_3088);
nand U4376 (N_4376,N_3468,N_3121);
and U4377 (N_4377,N_3361,N_3029);
nand U4378 (N_4378,N_3406,N_3156);
nand U4379 (N_4379,N_3640,N_3602);
xor U4380 (N_4380,N_3596,N_3689);
nor U4381 (N_4381,N_3300,N_3990);
or U4382 (N_4382,N_3485,N_3770);
xnor U4383 (N_4383,N_3471,N_3797);
nor U4384 (N_4384,N_3341,N_3774);
nand U4385 (N_4385,N_3190,N_3510);
nor U4386 (N_4386,N_3454,N_3518);
or U4387 (N_4387,N_3379,N_3046);
or U4388 (N_4388,N_3041,N_3910);
xnor U4389 (N_4389,N_3767,N_3891);
xnor U4390 (N_4390,N_3436,N_3347);
nand U4391 (N_4391,N_3638,N_3067);
or U4392 (N_4392,N_3399,N_3330);
nand U4393 (N_4393,N_3061,N_3895);
and U4394 (N_4394,N_3074,N_3111);
or U4395 (N_4395,N_3949,N_3107);
xnor U4396 (N_4396,N_3259,N_3089);
or U4397 (N_4397,N_3422,N_3087);
and U4398 (N_4398,N_3285,N_3829);
nor U4399 (N_4399,N_3551,N_3630);
nand U4400 (N_4400,N_3572,N_3013);
nand U4401 (N_4401,N_3172,N_3619);
nor U4402 (N_4402,N_3853,N_3353);
nand U4403 (N_4403,N_3665,N_3051);
xor U4404 (N_4404,N_3286,N_3387);
nor U4405 (N_4405,N_3769,N_3019);
xnor U4406 (N_4406,N_3412,N_3194);
and U4407 (N_4407,N_3196,N_3206);
nor U4408 (N_4408,N_3790,N_3474);
xnor U4409 (N_4409,N_3212,N_3999);
nor U4410 (N_4410,N_3909,N_3542);
and U4411 (N_4411,N_3169,N_3419);
and U4412 (N_4412,N_3199,N_3625);
and U4413 (N_4413,N_3861,N_3478);
xnor U4414 (N_4414,N_3213,N_3590);
nor U4415 (N_4415,N_3000,N_3843);
xor U4416 (N_4416,N_3413,N_3498);
or U4417 (N_4417,N_3661,N_3279);
and U4418 (N_4418,N_3175,N_3382);
or U4419 (N_4419,N_3373,N_3308);
nand U4420 (N_4420,N_3344,N_3181);
nor U4421 (N_4421,N_3113,N_3647);
and U4422 (N_4422,N_3878,N_3004);
nor U4423 (N_4423,N_3931,N_3972);
nand U4424 (N_4424,N_3037,N_3697);
xnor U4425 (N_4425,N_3671,N_3681);
nor U4426 (N_4426,N_3314,N_3901);
nor U4427 (N_4427,N_3077,N_3356);
and U4428 (N_4428,N_3270,N_3727);
and U4429 (N_4429,N_3352,N_3219);
nor U4430 (N_4430,N_3007,N_3837);
nor U4431 (N_4431,N_3775,N_3835);
xor U4432 (N_4432,N_3832,N_3354);
or U4433 (N_4433,N_3592,N_3694);
and U4434 (N_4434,N_3523,N_3415);
nor U4435 (N_4435,N_3450,N_3495);
and U4436 (N_4436,N_3699,N_3520);
nor U4437 (N_4437,N_3939,N_3076);
or U4438 (N_4438,N_3006,N_3179);
or U4439 (N_4439,N_3673,N_3063);
nor U4440 (N_4440,N_3440,N_3464);
nor U4441 (N_4441,N_3362,N_3613);
xnor U4442 (N_4442,N_3310,N_3336);
nor U4443 (N_4443,N_3960,N_3519);
and U4444 (N_4444,N_3434,N_3187);
and U4445 (N_4445,N_3503,N_3992);
nand U4446 (N_4446,N_3969,N_3389);
nor U4447 (N_4447,N_3564,N_3282);
nor U4448 (N_4448,N_3712,N_3224);
nor U4449 (N_4449,N_3643,N_3233);
nor U4450 (N_4450,N_3704,N_3393);
or U4451 (N_4451,N_3339,N_3008);
or U4452 (N_4452,N_3501,N_3295);
nand U4453 (N_4453,N_3844,N_3872);
nor U4454 (N_4454,N_3836,N_3970);
nor U4455 (N_4455,N_3268,N_3792);
or U4456 (N_4456,N_3821,N_3856);
xor U4457 (N_4457,N_3384,N_3430);
nand U4458 (N_4458,N_3391,N_3729);
nand U4459 (N_4459,N_3627,N_3612);
and U4460 (N_4460,N_3015,N_3253);
nor U4461 (N_4461,N_3682,N_3566);
and U4462 (N_4462,N_3120,N_3066);
nand U4463 (N_4463,N_3525,N_3841);
nand U4464 (N_4464,N_3048,N_3256);
or U4465 (N_4465,N_3658,N_3433);
and U4466 (N_4466,N_3669,N_3582);
or U4467 (N_4467,N_3745,N_3092);
nand U4468 (N_4468,N_3830,N_3631);
or U4469 (N_4469,N_3346,N_3043);
or U4470 (N_4470,N_3946,N_3481);
and U4471 (N_4471,N_3634,N_3544);
nand U4472 (N_4472,N_3866,N_3550);
and U4473 (N_4473,N_3851,N_3367);
or U4474 (N_4474,N_3814,N_3333);
or U4475 (N_4475,N_3388,N_3746);
nor U4476 (N_4476,N_3071,N_3930);
nor U4477 (N_4477,N_3677,N_3758);
nor U4478 (N_4478,N_3765,N_3435);
xnor U4479 (N_4479,N_3218,N_3429);
xnor U4480 (N_4480,N_3360,N_3101);
nor U4481 (N_4481,N_3701,N_3052);
and U4482 (N_4482,N_3177,N_3297);
and U4483 (N_4483,N_3777,N_3162);
or U4484 (N_4484,N_3606,N_3299);
nand U4485 (N_4485,N_3426,N_3693);
and U4486 (N_4486,N_3059,N_3470);
xor U4487 (N_4487,N_3342,N_3726);
nand U4488 (N_4488,N_3731,N_3705);
and U4489 (N_4489,N_3251,N_3599);
nand U4490 (N_4490,N_3686,N_3198);
and U4491 (N_4491,N_3578,N_3988);
nand U4492 (N_4492,N_3201,N_3461);
and U4493 (N_4493,N_3173,N_3706);
or U4494 (N_4494,N_3776,N_3020);
and U4495 (N_4495,N_3709,N_3507);
and U4496 (N_4496,N_3315,N_3958);
nand U4497 (N_4497,N_3138,N_3012);
or U4498 (N_4498,N_3994,N_3421);
nor U4499 (N_4499,N_3754,N_3488);
or U4500 (N_4500,N_3260,N_3161);
and U4501 (N_4501,N_3819,N_3121);
and U4502 (N_4502,N_3932,N_3680);
and U4503 (N_4503,N_3635,N_3427);
and U4504 (N_4504,N_3755,N_3066);
nor U4505 (N_4505,N_3338,N_3094);
nor U4506 (N_4506,N_3516,N_3405);
nor U4507 (N_4507,N_3216,N_3693);
or U4508 (N_4508,N_3747,N_3692);
nor U4509 (N_4509,N_3324,N_3743);
nor U4510 (N_4510,N_3555,N_3094);
and U4511 (N_4511,N_3526,N_3411);
and U4512 (N_4512,N_3241,N_3160);
nand U4513 (N_4513,N_3459,N_3010);
nand U4514 (N_4514,N_3711,N_3834);
or U4515 (N_4515,N_3009,N_3720);
or U4516 (N_4516,N_3989,N_3075);
nand U4517 (N_4517,N_3927,N_3896);
or U4518 (N_4518,N_3354,N_3305);
nor U4519 (N_4519,N_3382,N_3467);
and U4520 (N_4520,N_3742,N_3836);
and U4521 (N_4521,N_3387,N_3182);
or U4522 (N_4522,N_3883,N_3349);
nand U4523 (N_4523,N_3568,N_3718);
nor U4524 (N_4524,N_3465,N_3563);
nand U4525 (N_4525,N_3173,N_3970);
and U4526 (N_4526,N_3024,N_3999);
nand U4527 (N_4527,N_3444,N_3660);
or U4528 (N_4528,N_3405,N_3602);
or U4529 (N_4529,N_3895,N_3675);
and U4530 (N_4530,N_3977,N_3434);
and U4531 (N_4531,N_3789,N_3704);
or U4532 (N_4532,N_3961,N_3074);
nor U4533 (N_4533,N_3970,N_3694);
nor U4534 (N_4534,N_3230,N_3536);
or U4535 (N_4535,N_3565,N_3130);
nor U4536 (N_4536,N_3822,N_3407);
and U4537 (N_4537,N_3797,N_3395);
xnor U4538 (N_4538,N_3284,N_3962);
nor U4539 (N_4539,N_3978,N_3126);
nand U4540 (N_4540,N_3736,N_3126);
or U4541 (N_4541,N_3015,N_3980);
nor U4542 (N_4542,N_3311,N_3195);
and U4543 (N_4543,N_3851,N_3321);
nand U4544 (N_4544,N_3872,N_3593);
and U4545 (N_4545,N_3273,N_3553);
or U4546 (N_4546,N_3043,N_3214);
nor U4547 (N_4547,N_3387,N_3844);
and U4548 (N_4548,N_3652,N_3150);
or U4549 (N_4549,N_3956,N_3344);
xnor U4550 (N_4550,N_3397,N_3531);
nand U4551 (N_4551,N_3040,N_3618);
or U4552 (N_4552,N_3325,N_3153);
and U4553 (N_4553,N_3590,N_3448);
and U4554 (N_4554,N_3941,N_3837);
xnor U4555 (N_4555,N_3624,N_3699);
and U4556 (N_4556,N_3637,N_3741);
nand U4557 (N_4557,N_3950,N_3398);
nand U4558 (N_4558,N_3880,N_3626);
and U4559 (N_4559,N_3192,N_3506);
nor U4560 (N_4560,N_3869,N_3165);
nand U4561 (N_4561,N_3460,N_3409);
or U4562 (N_4562,N_3946,N_3693);
nand U4563 (N_4563,N_3783,N_3999);
and U4564 (N_4564,N_3189,N_3599);
and U4565 (N_4565,N_3601,N_3895);
or U4566 (N_4566,N_3541,N_3165);
or U4567 (N_4567,N_3803,N_3471);
or U4568 (N_4568,N_3307,N_3147);
and U4569 (N_4569,N_3239,N_3647);
and U4570 (N_4570,N_3082,N_3229);
nand U4571 (N_4571,N_3904,N_3251);
nand U4572 (N_4572,N_3821,N_3324);
nor U4573 (N_4573,N_3304,N_3203);
or U4574 (N_4574,N_3917,N_3577);
and U4575 (N_4575,N_3809,N_3267);
or U4576 (N_4576,N_3704,N_3726);
and U4577 (N_4577,N_3208,N_3785);
nor U4578 (N_4578,N_3509,N_3082);
or U4579 (N_4579,N_3127,N_3304);
and U4580 (N_4580,N_3304,N_3965);
nor U4581 (N_4581,N_3384,N_3813);
nor U4582 (N_4582,N_3559,N_3684);
nor U4583 (N_4583,N_3153,N_3106);
or U4584 (N_4584,N_3741,N_3384);
or U4585 (N_4585,N_3913,N_3154);
nor U4586 (N_4586,N_3991,N_3160);
or U4587 (N_4587,N_3090,N_3947);
nor U4588 (N_4588,N_3912,N_3306);
xor U4589 (N_4589,N_3332,N_3669);
xnor U4590 (N_4590,N_3324,N_3824);
or U4591 (N_4591,N_3881,N_3608);
or U4592 (N_4592,N_3916,N_3773);
and U4593 (N_4593,N_3099,N_3776);
nor U4594 (N_4594,N_3789,N_3411);
and U4595 (N_4595,N_3562,N_3805);
nor U4596 (N_4596,N_3245,N_3984);
or U4597 (N_4597,N_3312,N_3557);
nor U4598 (N_4598,N_3543,N_3944);
nor U4599 (N_4599,N_3336,N_3026);
nor U4600 (N_4600,N_3036,N_3628);
or U4601 (N_4601,N_3946,N_3716);
and U4602 (N_4602,N_3203,N_3484);
or U4603 (N_4603,N_3019,N_3270);
or U4604 (N_4604,N_3869,N_3911);
nand U4605 (N_4605,N_3127,N_3717);
xor U4606 (N_4606,N_3958,N_3345);
nand U4607 (N_4607,N_3129,N_3998);
nor U4608 (N_4608,N_3177,N_3755);
nor U4609 (N_4609,N_3550,N_3340);
or U4610 (N_4610,N_3299,N_3008);
or U4611 (N_4611,N_3401,N_3778);
nand U4612 (N_4612,N_3993,N_3219);
and U4613 (N_4613,N_3968,N_3569);
nand U4614 (N_4614,N_3553,N_3334);
nand U4615 (N_4615,N_3028,N_3466);
and U4616 (N_4616,N_3982,N_3304);
and U4617 (N_4617,N_3113,N_3597);
and U4618 (N_4618,N_3219,N_3558);
nor U4619 (N_4619,N_3198,N_3031);
or U4620 (N_4620,N_3451,N_3484);
nand U4621 (N_4621,N_3025,N_3442);
xnor U4622 (N_4622,N_3578,N_3274);
nand U4623 (N_4623,N_3234,N_3243);
nand U4624 (N_4624,N_3570,N_3412);
nor U4625 (N_4625,N_3418,N_3608);
nand U4626 (N_4626,N_3867,N_3172);
or U4627 (N_4627,N_3560,N_3397);
nand U4628 (N_4628,N_3515,N_3950);
nor U4629 (N_4629,N_3166,N_3503);
and U4630 (N_4630,N_3035,N_3103);
nand U4631 (N_4631,N_3049,N_3378);
and U4632 (N_4632,N_3441,N_3307);
and U4633 (N_4633,N_3841,N_3063);
or U4634 (N_4634,N_3492,N_3330);
or U4635 (N_4635,N_3700,N_3563);
nand U4636 (N_4636,N_3043,N_3690);
xnor U4637 (N_4637,N_3241,N_3229);
or U4638 (N_4638,N_3572,N_3986);
nand U4639 (N_4639,N_3792,N_3181);
or U4640 (N_4640,N_3095,N_3596);
xnor U4641 (N_4641,N_3048,N_3397);
nand U4642 (N_4642,N_3188,N_3594);
nor U4643 (N_4643,N_3698,N_3594);
nand U4644 (N_4644,N_3817,N_3468);
nand U4645 (N_4645,N_3714,N_3337);
or U4646 (N_4646,N_3733,N_3171);
nand U4647 (N_4647,N_3855,N_3922);
nor U4648 (N_4648,N_3933,N_3660);
nand U4649 (N_4649,N_3549,N_3320);
and U4650 (N_4650,N_3018,N_3163);
or U4651 (N_4651,N_3216,N_3729);
and U4652 (N_4652,N_3770,N_3973);
nor U4653 (N_4653,N_3479,N_3212);
xnor U4654 (N_4654,N_3142,N_3963);
and U4655 (N_4655,N_3238,N_3201);
nor U4656 (N_4656,N_3541,N_3207);
nor U4657 (N_4657,N_3572,N_3442);
xor U4658 (N_4658,N_3851,N_3313);
or U4659 (N_4659,N_3541,N_3881);
xor U4660 (N_4660,N_3659,N_3427);
nor U4661 (N_4661,N_3543,N_3394);
and U4662 (N_4662,N_3662,N_3282);
nor U4663 (N_4663,N_3211,N_3755);
or U4664 (N_4664,N_3603,N_3659);
nand U4665 (N_4665,N_3813,N_3447);
or U4666 (N_4666,N_3872,N_3854);
nor U4667 (N_4667,N_3402,N_3748);
or U4668 (N_4668,N_3580,N_3781);
and U4669 (N_4669,N_3535,N_3027);
nor U4670 (N_4670,N_3620,N_3150);
nand U4671 (N_4671,N_3748,N_3703);
and U4672 (N_4672,N_3859,N_3958);
xor U4673 (N_4673,N_3658,N_3772);
nor U4674 (N_4674,N_3279,N_3192);
nor U4675 (N_4675,N_3213,N_3922);
nand U4676 (N_4676,N_3827,N_3079);
nor U4677 (N_4677,N_3610,N_3796);
and U4678 (N_4678,N_3672,N_3816);
nand U4679 (N_4679,N_3684,N_3900);
or U4680 (N_4680,N_3285,N_3668);
xnor U4681 (N_4681,N_3881,N_3354);
or U4682 (N_4682,N_3742,N_3733);
and U4683 (N_4683,N_3452,N_3102);
and U4684 (N_4684,N_3707,N_3740);
nor U4685 (N_4685,N_3835,N_3330);
xnor U4686 (N_4686,N_3804,N_3430);
and U4687 (N_4687,N_3844,N_3914);
nand U4688 (N_4688,N_3590,N_3940);
or U4689 (N_4689,N_3225,N_3592);
xnor U4690 (N_4690,N_3380,N_3785);
or U4691 (N_4691,N_3877,N_3955);
nand U4692 (N_4692,N_3698,N_3868);
or U4693 (N_4693,N_3213,N_3795);
and U4694 (N_4694,N_3943,N_3879);
xnor U4695 (N_4695,N_3643,N_3236);
or U4696 (N_4696,N_3424,N_3608);
nor U4697 (N_4697,N_3944,N_3355);
or U4698 (N_4698,N_3714,N_3744);
or U4699 (N_4699,N_3686,N_3849);
nand U4700 (N_4700,N_3859,N_3183);
nor U4701 (N_4701,N_3385,N_3376);
nand U4702 (N_4702,N_3632,N_3536);
and U4703 (N_4703,N_3050,N_3242);
nand U4704 (N_4704,N_3452,N_3994);
nor U4705 (N_4705,N_3780,N_3204);
nand U4706 (N_4706,N_3662,N_3869);
or U4707 (N_4707,N_3044,N_3617);
nor U4708 (N_4708,N_3982,N_3141);
and U4709 (N_4709,N_3393,N_3517);
and U4710 (N_4710,N_3694,N_3365);
nand U4711 (N_4711,N_3188,N_3417);
nand U4712 (N_4712,N_3316,N_3718);
or U4713 (N_4713,N_3754,N_3736);
or U4714 (N_4714,N_3512,N_3510);
nor U4715 (N_4715,N_3481,N_3153);
nor U4716 (N_4716,N_3515,N_3481);
or U4717 (N_4717,N_3331,N_3298);
nor U4718 (N_4718,N_3072,N_3849);
nand U4719 (N_4719,N_3039,N_3447);
nand U4720 (N_4720,N_3690,N_3823);
or U4721 (N_4721,N_3077,N_3398);
xnor U4722 (N_4722,N_3531,N_3376);
nand U4723 (N_4723,N_3061,N_3055);
nor U4724 (N_4724,N_3096,N_3087);
nand U4725 (N_4725,N_3627,N_3243);
or U4726 (N_4726,N_3834,N_3436);
nor U4727 (N_4727,N_3379,N_3436);
nor U4728 (N_4728,N_3353,N_3204);
nor U4729 (N_4729,N_3733,N_3215);
and U4730 (N_4730,N_3677,N_3354);
and U4731 (N_4731,N_3314,N_3196);
or U4732 (N_4732,N_3723,N_3661);
and U4733 (N_4733,N_3622,N_3292);
or U4734 (N_4734,N_3789,N_3199);
nand U4735 (N_4735,N_3914,N_3145);
nand U4736 (N_4736,N_3361,N_3597);
nor U4737 (N_4737,N_3378,N_3645);
or U4738 (N_4738,N_3934,N_3016);
or U4739 (N_4739,N_3915,N_3631);
nor U4740 (N_4740,N_3428,N_3789);
or U4741 (N_4741,N_3452,N_3864);
nor U4742 (N_4742,N_3382,N_3759);
nor U4743 (N_4743,N_3786,N_3635);
nand U4744 (N_4744,N_3589,N_3757);
and U4745 (N_4745,N_3499,N_3233);
nand U4746 (N_4746,N_3767,N_3778);
or U4747 (N_4747,N_3166,N_3913);
nand U4748 (N_4748,N_3948,N_3851);
nor U4749 (N_4749,N_3712,N_3235);
xor U4750 (N_4750,N_3812,N_3192);
or U4751 (N_4751,N_3415,N_3942);
and U4752 (N_4752,N_3874,N_3767);
nand U4753 (N_4753,N_3680,N_3601);
or U4754 (N_4754,N_3815,N_3223);
nor U4755 (N_4755,N_3105,N_3453);
xnor U4756 (N_4756,N_3653,N_3407);
nor U4757 (N_4757,N_3022,N_3961);
xnor U4758 (N_4758,N_3735,N_3829);
nand U4759 (N_4759,N_3436,N_3626);
or U4760 (N_4760,N_3628,N_3266);
nand U4761 (N_4761,N_3138,N_3949);
or U4762 (N_4762,N_3684,N_3156);
or U4763 (N_4763,N_3907,N_3823);
or U4764 (N_4764,N_3794,N_3539);
and U4765 (N_4765,N_3034,N_3523);
or U4766 (N_4766,N_3707,N_3135);
nand U4767 (N_4767,N_3416,N_3915);
xor U4768 (N_4768,N_3925,N_3605);
and U4769 (N_4769,N_3315,N_3799);
and U4770 (N_4770,N_3137,N_3819);
or U4771 (N_4771,N_3841,N_3982);
nor U4772 (N_4772,N_3620,N_3066);
nand U4773 (N_4773,N_3198,N_3526);
or U4774 (N_4774,N_3519,N_3081);
nor U4775 (N_4775,N_3432,N_3589);
xnor U4776 (N_4776,N_3784,N_3948);
nand U4777 (N_4777,N_3957,N_3554);
nand U4778 (N_4778,N_3503,N_3743);
nor U4779 (N_4779,N_3594,N_3904);
nand U4780 (N_4780,N_3199,N_3583);
and U4781 (N_4781,N_3471,N_3841);
or U4782 (N_4782,N_3610,N_3652);
nor U4783 (N_4783,N_3891,N_3084);
and U4784 (N_4784,N_3909,N_3935);
and U4785 (N_4785,N_3328,N_3282);
and U4786 (N_4786,N_3030,N_3854);
nor U4787 (N_4787,N_3201,N_3243);
nor U4788 (N_4788,N_3031,N_3651);
nand U4789 (N_4789,N_3108,N_3142);
and U4790 (N_4790,N_3845,N_3774);
or U4791 (N_4791,N_3320,N_3596);
and U4792 (N_4792,N_3232,N_3550);
or U4793 (N_4793,N_3044,N_3451);
nand U4794 (N_4794,N_3372,N_3105);
and U4795 (N_4795,N_3840,N_3870);
or U4796 (N_4796,N_3615,N_3959);
and U4797 (N_4797,N_3793,N_3787);
nand U4798 (N_4798,N_3448,N_3543);
nand U4799 (N_4799,N_3184,N_3471);
or U4800 (N_4800,N_3813,N_3473);
nor U4801 (N_4801,N_3917,N_3620);
and U4802 (N_4802,N_3431,N_3610);
and U4803 (N_4803,N_3163,N_3408);
or U4804 (N_4804,N_3896,N_3023);
nor U4805 (N_4805,N_3006,N_3385);
nor U4806 (N_4806,N_3419,N_3438);
or U4807 (N_4807,N_3182,N_3415);
xor U4808 (N_4808,N_3021,N_3322);
nand U4809 (N_4809,N_3118,N_3185);
and U4810 (N_4810,N_3063,N_3551);
nand U4811 (N_4811,N_3204,N_3406);
or U4812 (N_4812,N_3656,N_3890);
xnor U4813 (N_4813,N_3806,N_3662);
nand U4814 (N_4814,N_3436,N_3054);
nand U4815 (N_4815,N_3833,N_3693);
xor U4816 (N_4816,N_3103,N_3269);
and U4817 (N_4817,N_3068,N_3732);
or U4818 (N_4818,N_3015,N_3785);
and U4819 (N_4819,N_3577,N_3986);
nor U4820 (N_4820,N_3237,N_3674);
nor U4821 (N_4821,N_3412,N_3088);
nor U4822 (N_4822,N_3545,N_3398);
xor U4823 (N_4823,N_3063,N_3521);
and U4824 (N_4824,N_3026,N_3478);
and U4825 (N_4825,N_3079,N_3490);
nand U4826 (N_4826,N_3417,N_3605);
or U4827 (N_4827,N_3761,N_3157);
and U4828 (N_4828,N_3510,N_3399);
and U4829 (N_4829,N_3266,N_3895);
or U4830 (N_4830,N_3759,N_3966);
nor U4831 (N_4831,N_3889,N_3127);
and U4832 (N_4832,N_3921,N_3706);
nand U4833 (N_4833,N_3663,N_3082);
and U4834 (N_4834,N_3790,N_3428);
nor U4835 (N_4835,N_3301,N_3450);
nand U4836 (N_4836,N_3803,N_3305);
or U4837 (N_4837,N_3801,N_3968);
nor U4838 (N_4838,N_3940,N_3956);
nand U4839 (N_4839,N_3070,N_3328);
nor U4840 (N_4840,N_3886,N_3955);
xnor U4841 (N_4841,N_3668,N_3396);
nor U4842 (N_4842,N_3501,N_3959);
or U4843 (N_4843,N_3091,N_3639);
nand U4844 (N_4844,N_3588,N_3037);
nand U4845 (N_4845,N_3035,N_3407);
and U4846 (N_4846,N_3543,N_3830);
nor U4847 (N_4847,N_3328,N_3206);
xor U4848 (N_4848,N_3639,N_3658);
or U4849 (N_4849,N_3201,N_3393);
or U4850 (N_4850,N_3112,N_3210);
and U4851 (N_4851,N_3226,N_3618);
and U4852 (N_4852,N_3854,N_3285);
or U4853 (N_4853,N_3958,N_3161);
or U4854 (N_4854,N_3266,N_3758);
or U4855 (N_4855,N_3432,N_3934);
nand U4856 (N_4856,N_3502,N_3763);
or U4857 (N_4857,N_3283,N_3340);
nand U4858 (N_4858,N_3917,N_3764);
nand U4859 (N_4859,N_3982,N_3498);
nand U4860 (N_4860,N_3047,N_3861);
and U4861 (N_4861,N_3096,N_3462);
nor U4862 (N_4862,N_3924,N_3462);
and U4863 (N_4863,N_3902,N_3746);
xor U4864 (N_4864,N_3045,N_3844);
xor U4865 (N_4865,N_3356,N_3257);
or U4866 (N_4866,N_3990,N_3121);
and U4867 (N_4867,N_3628,N_3486);
or U4868 (N_4868,N_3109,N_3582);
nand U4869 (N_4869,N_3863,N_3046);
nor U4870 (N_4870,N_3019,N_3207);
nor U4871 (N_4871,N_3208,N_3086);
xnor U4872 (N_4872,N_3951,N_3679);
nand U4873 (N_4873,N_3830,N_3792);
nor U4874 (N_4874,N_3837,N_3761);
xor U4875 (N_4875,N_3697,N_3532);
or U4876 (N_4876,N_3187,N_3271);
nand U4877 (N_4877,N_3747,N_3003);
or U4878 (N_4878,N_3978,N_3503);
and U4879 (N_4879,N_3631,N_3714);
and U4880 (N_4880,N_3075,N_3188);
and U4881 (N_4881,N_3753,N_3472);
xor U4882 (N_4882,N_3741,N_3744);
nand U4883 (N_4883,N_3601,N_3761);
nand U4884 (N_4884,N_3455,N_3421);
xor U4885 (N_4885,N_3393,N_3348);
and U4886 (N_4886,N_3854,N_3652);
nand U4887 (N_4887,N_3281,N_3798);
and U4888 (N_4888,N_3234,N_3346);
and U4889 (N_4889,N_3491,N_3312);
or U4890 (N_4890,N_3816,N_3751);
xor U4891 (N_4891,N_3233,N_3400);
and U4892 (N_4892,N_3179,N_3657);
xnor U4893 (N_4893,N_3877,N_3565);
nor U4894 (N_4894,N_3880,N_3435);
nand U4895 (N_4895,N_3158,N_3064);
nand U4896 (N_4896,N_3139,N_3206);
nand U4897 (N_4897,N_3392,N_3225);
and U4898 (N_4898,N_3194,N_3155);
nand U4899 (N_4899,N_3360,N_3951);
and U4900 (N_4900,N_3810,N_3430);
and U4901 (N_4901,N_3349,N_3855);
or U4902 (N_4902,N_3461,N_3385);
xnor U4903 (N_4903,N_3558,N_3782);
and U4904 (N_4904,N_3309,N_3225);
nand U4905 (N_4905,N_3188,N_3394);
and U4906 (N_4906,N_3072,N_3163);
nand U4907 (N_4907,N_3906,N_3542);
nand U4908 (N_4908,N_3354,N_3938);
nor U4909 (N_4909,N_3389,N_3161);
nand U4910 (N_4910,N_3695,N_3438);
nand U4911 (N_4911,N_3046,N_3887);
and U4912 (N_4912,N_3316,N_3878);
and U4913 (N_4913,N_3527,N_3554);
or U4914 (N_4914,N_3014,N_3631);
or U4915 (N_4915,N_3328,N_3641);
nand U4916 (N_4916,N_3301,N_3836);
nand U4917 (N_4917,N_3989,N_3149);
or U4918 (N_4918,N_3091,N_3740);
nand U4919 (N_4919,N_3382,N_3496);
and U4920 (N_4920,N_3330,N_3475);
nand U4921 (N_4921,N_3951,N_3332);
xor U4922 (N_4922,N_3260,N_3666);
or U4923 (N_4923,N_3212,N_3060);
and U4924 (N_4924,N_3703,N_3617);
or U4925 (N_4925,N_3960,N_3004);
nand U4926 (N_4926,N_3140,N_3905);
and U4927 (N_4927,N_3686,N_3009);
and U4928 (N_4928,N_3100,N_3216);
or U4929 (N_4929,N_3206,N_3797);
nand U4930 (N_4930,N_3642,N_3161);
nor U4931 (N_4931,N_3337,N_3042);
or U4932 (N_4932,N_3515,N_3360);
nor U4933 (N_4933,N_3460,N_3535);
and U4934 (N_4934,N_3000,N_3604);
and U4935 (N_4935,N_3596,N_3459);
and U4936 (N_4936,N_3215,N_3233);
nand U4937 (N_4937,N_3146,N_3847);
and U4938 (N_4938,N_3168,N_3275);
nor U4939 (N_4939,N_3220,N_3288);
or U4940 (N_4940,N_3543,N_3593);
and U4941 (N_4941,N_3717,N_3903);
and U4942 (N_4942,N_3508,N_3115);
and U4943 (N_4943,N_3620,N_3948);
and U4944 (N_4944,N_3955,N_3651);
xnor U4945 (N_4945,N_3023,N_3907);
and U4946 (N_4946,N_3636,N_3733);
and U4947 (N_4947,N_3377,N_3971);
xor U4948 (N_4948,N_3794,N_3939);
nand U4949 (N_4949,N_3470,N_3365);
nand U4950 (N_4950,N_3147,N_3059);
nand U4951 (N_4951,N_3578,N_3192);
and U4952 (N_4952,N_3583,N_3098);
xor U4953 (N_4953,N_3257,N_3194);
nand U4954 (N_4954,N_3776,N_3973);
nand U4955 (N_4955,N_3116,N_3162);
nand U4956 (N_4956,N_3025,N_3470);
nand U4957 (N_4957,N_3271,N_3845);
xnor U4958 (N_4958,N_3809,N_3820);
and U4959 (N_4959,N_3886,N_3005);
or U4960 (N_4960,N_3140,N_3062);
and U4961 (N_4961,N_3466,N_3884);
nand U4962 (N_4962,N_3203,N_3941);
nor U4963 (N_4963,N_3788,N_3271);
nor U4964 (N_4964,N_3413,N_3935);
and U4965 (N_4965,N_3718,N_3311);
nor U4966 (N_4966,N_3950,N_3594);
or U4967 (N_4967,N_3229,N_3578);
and U4968 (N_4968,N_3018,N_3659);
or U4969 (N_4969,N_3614,N_3098);
nor U4970 (N_4970,N_3810,N_3523);
and U4971 (N_4971,N_3792,N_3772);
nor U4972 (N_4972,N_3526,N_3034);
and U4973 (N_4973,N_3663,N_3956);
nor U4974 (N_4974,N_3129,N_3024);
and U4975 (N_4975,N_3640,N_3158);
nor U4976 (N_4976,N_3737,N_3632);
xnor U4977 (N_4977,N_3331,N_3768);
and U4978 (N_4978,N_3728,N_3396);
nor U4979 (N_4979,N_3794,N_3370);
and U4980 (N_4980,N_3735,N_3365);
xnor U4981 (N_4981,N_3685,N_3642);
and U4982 (N_4982,N_3624,N_3054);
or U4983 (N_4983,N_3476,N_3496);
or U4984 (N_4984,N_3829,N_3233);
or U4985 (N_4985,N_3793,N_3929);
or U4986 (N_4986,N_3363,N_3843);
nand U4987 (N_4987,N_3254,N_3495);
and U4988 (N_4988,N_3428,N_3163);
or U4989 (N_4989,N_3801,N_3954);
nand U4990 (N_4990,N_3053,N_3611);
nor U4991 (N_4991,N_3509,N_3280);
nor U4992 (N_4992,N_3784,N_3902);
nor U4993 (N_4993,N_3356,N_3383);
or U4994 (N_4994,N_3899,N_3788);
and U4995 (N_4995,N_3004,N_3738);
and U4996 (N_4996,N_3337,N_3699);
nor U4997 (N_4997,N_3654,N_3942);
and U4998 (N_4998,N_3215,N_3797);
and U4999 (N_4999,N_3502,N_3222);
xnor U5000 (N_5000,N_4746,N_4330);
nand U5001 (N_5001,N_4027,N_4081);
nor U5002 (N_5002,N_4151,N_4362);
xor U5003 (N_5003,N_4324,N_4458);
and U5004 (N_5004,N_4024,N_4054);
nand U5005 (N_5005,N_4492,N_4471);
nor U5006 (N_5006,N_4956,N_4602);
and U5007 (N_5007,N_4754,N_4539);
and U5008 (N_5008,N_4398,N_4581);
or U5009 (N_5009,N_4600,N_4144);
nor U5010 (N_5010,N_4283,N_4409);
nor U5011 (N_5011,N_4040,N_4023);
and U5012 (N_5012,N_4293,N_4031);
or U5013 (N_5013,N_4604,N_4466);
xor U5014 (N_5014,N_4046,N_4993);
nor U5015 (N_5015,N_4473,N_4617);
nor U5016 (N_5016,N_4937,N_4109);
nand U5017 (N_5017,N_4171,N_4227);
nor U5018 (N_5018,N_4459,N_4947);
or U5019 (N_5019,N_4340,N_4176);
xnor U5020 (N_5020,N_4035,N_4018);
xnor U5021 (N_5021,N_4851,N_4463);
or U5022 (N_5022,N_4958,N_4977);
nor U5023 (N_5023,N_4590,N_4796);
and U5024 (N_5024,N_4509,N_4478);
nor U5025 (N_5025,N_4136,N_4964);
and U5026 (N_5026,N_4211,N_4990);
or U5027 (N_5027,N_4260,N_4702);
nor U5028 (N_5028,N_4195,N_4598);
and U5029 (N_5029,N_4716,N_4767);
xor U5030 (N_5030,N_4676,N_4788);
and U5031 (N_5031,N_4436,N_4631);
xnor U5032 (N_5032,N_4460,N_4221);
and U5033 (N_5033,N_4942,N_4725);
and U5034 (N_5034,N_4935,N_4419);
xor U5035 (N_5035,N_4808,N_4430);
nand U5036 (N_5036,N_4072,N_4969);
nand U5037 (N_5037,N_4428,N_4665);
nor U5038 (N_5038,N_4254,N_4675);
nor U5039 (N_5039,N_4306,N_4913);
or U5040 (N_5040,N_4143,N_4500);
and U5041 (N_5041,N_4295,N_4216);
nor U5042 (N_5042,N_4495,N_4313);
nand U5043 (N_5043,N_4597,N_4455);
nor U5044 (N_5044,N_4548,N_4641);
and U5045 (N_5045,N_4100,N_4535);
or U5046 (N_5046,N_4710,N_4231);
nand U5047 (N_5047,N_4950,N_4779);
nor U5048 (N_5048,N_4257,N_4824);
or U5049 (N_5049,N_4606,N_4513);
nor U5050 (N_5050,N_4250,N_4294);
nand U5051 (N_5051,N_4396,N_4467);
nand U5052 (N_5052,N_4524,N_4367);
nand U5053 (N_5053,N_4738,N_4593);
nand U5054 (N_5054,N_4859,N_4288);
nand U5055 (N_5055,N_4213,N_4968);
nor U5056 (N_5056,N_4538,N_4265);
nand U5057 (N_5057,N_4233,N_4762);
and U5058 (N_5058,N_4029,N_4642);
or U5059 (N_5059,N_4579,N_4658);
and U5060 (N_5060,N_4925,N_4749);
nand U5061 (N_5061,N_4536,N_4476);
nand U5062 (N_5062,N_4025,N_4487);
nand U5063 (N_5063,N_4517,N_4899);
nand U5064 (N_5064,N_4315,N_4668);
or U5065 (N_5065,N_4255,N_4994);
nor U5066 (N_5066,N_4192,N_4044);
xor U5067 (N_5067,N_4416,N_4532);
and U5068 (N_5068,N_4425,N_4089);
and U5069 (N_5069,N_4888,N_4483);
nand U5070 (N_5070,N_4618,N_4045);
nor U5071 (N_5071,N_4972,N_4032);
and U5072 (N_5072,N_4744,N_4621);
xor U5073 (N_5073,N_4502,N_4101);
and U5074 (N_5074,N_4690,N_4472);
or U5075 (N_5075,N_4301,N_4526);
and U5076 (N_5076,N_4686,N_4026);
and U5077 (N_5077,N_4141,N_4804);
and U5078 (N_5078,N_4574,N_4713);
nor U5079 (N_5079,N_4060,N_4612);
nor U5080 (N_5080,N_4407,N_4012);
or U5081 (N_5081,N_4527,N_4567);
and U5082 (N_5082,N_4393,N_4893);
and U5083 (N_5083,N_4701,N_4599);
nor U5084 (N_5084,N_4922,N_4875);
and U5085 (N_5085,N_4773,N_4534);
or U5086 (N_5086,N_4537,N_4772);
or U5087 (N_5087,N_4501,N_4789);
nand U5088 (N_5088,N_4154,N_4733);
nor U5089 (N_5089,N_4672,N_4943);
and U5090 (N_5090,N_4783,N_4058);
or U5091 (N_5091,N_4004,N_4659);
and U5092 (N_5092,N_4855,N_4902);
xor U5093 (N_5093,N_4203,N_4333);
or U5094 (N_5094,N_4242,N_4774);
and U5095 (N_5095,N_4441,N_4812);
or U5096 (N_5096,N_4322,N_4303);
nor U5097 (N_5097,N_4670,N_4128);
and U5098 (N_5098,N_4966,N_4437);
or U5099 (N_5099,N_4368,N_4785);
nor U5100 (N_5100,N_4087,N_4861);
nor U5101 (N_5101,N_4155,N_4841);
nand U5102 (N_5102,N_4243,N_4415);
nor U5103 (N_5103,N_4892,N_4818);
or U5104 (N_5104,N_4369,N_4830);
xnor U5105 (N_5105,N_4989,N_4280);
nor U5106 (N_5106,N_4119,N_4829);
nand U5107 (N_5107,N_4177,N_4167);
or U5108 (N_5108,N_4022,N_4560);
and U5109 (N_5109,N_4669,N_4199);
or U5110 (N_5110,N_4692,N_4279);
nor U5111 (N_5111,N_4955,N_4585);
nand U5112 (N_5112,N_4055,N_4099);
nor U5113 (N_5113,N_4652,N_4169);
nor U5114 (N_5114,N_4435,N_4533);
nand U5115 (N_5115,N_4433,N_4912);
xnor U5116 (N_5116,N_4803,N_4857);
nand U5117 (N_5117,N_4186,N_4520);
nand U5118 (N_5118,N_4247,N_4223);
or U5119 (N_5119,N_4846,N_4939);
nand U5120 (N_5120,N_4831,N_4782);
or U5121 (N_5121,N_4129,N_4225);
or U5122 (N_5122,N_4619,N_4571);
nor U5123 (N_5123,N_4959,N_4062);
and U5124 (N_5124,N_4663,N_4148);
nand U5125 (N_5125,N_4292,N_4781);
or U5126 (N_5126,N_4936,N_4603);
nand U5127 (N_5127,N_4008,N_4575);
or U5128 (N_5128,N_4919,N_4084);
nand U5129 (N_5129,N_4165,N_4391);
xor U5130 (N_5130,N_4696,N_4275);
and U5131 (N_5131,N_4317,N_4891);
or U5132 (N_5132,N_4684,N_4777);
and U5133 (N_5133,N_4039,N_4797);
and U5134 (N_5134,N_4798,N_4107);
nor U5135 (N_5135,N_4735,N_4237);
or U5136 (N_5136,N_4354,N_4518);
nand U5137 (N_5137,N_4193,N_4314);
and U5138 (N_5138,N_4941,N_4140);
nand U5139 (N_5139,N_4461,N_4270);
or U5140 (N_5140,N_4775,N_4664);
nor U5141 (N_5141,N_4852,N_4146);
or U5142 (N_5142,N_4346,N_4302);
or U5143 (N_5143,N_4836,N_4932);
and U5144 (N_5144,N_4553,N_4699);
nand U5145 (N_5145,N_4508,N_4352);
nand U5146 (N_5146,N_4871,N_4776);
nor U5147 (N_5147,N_4312,N_4378);
and U5148 (N_5148,N_4421,N_4927);
nand U5149 (N_5149,N_4823,N_4429);
xnor U5150 (N_5150,N_4503,N_4863);
nand U5151 (N_5151,N_4931,N_4510);
and U5152 (N_5152,N_4271,N_4630);
nor U5153 (N_5153,N_4244,N_4149);
nor U5154 (N_5154,N_4150,N_4651);
nand U5155 (N_5155,N_4423,N_4856);
and U5156 (N_5156,N_4261,N_4468);
and U5157 (N_5157,N_4486,N_4923);
or U5158 (N_5158,N_4731,N_4066);
xor U5159 (N_5159,N_4674,N_4870);
nand U5160 (N_5160,N_4632,N_4883);
nor U5161 (N_5161,N_4805,N_4895);
xor U5162 (N_5162,N_4616,N_4813);
nand U5163 (N_5163,N_4918,N_4714);
or U5164 (N_5164,N_4137,N_4086);
and U5165 (N_5165,N_4505,N_4605);
nand U5166 (N_5166,N_4679,N_4700);
xnor U5167 (N_5167,N_4715,N_4240);
nand U5168 (N_5168,N_4007,N_4273);
nor U5169 (N_5169,N_4357,N_4438);
nand U5170 (N_5170,N_4729,N_4440);
nand U5171 (N_5171,N_4906,N_4626);
nor U5172 (N_5172,N_4952,N_4291);
nor U5173 (N_5173,N_4807,N_4342);
xor U5174 (N_5174,N_4979,N_4426);
nor U5175 (N_5175,N_4728,N_4077);
nand U5176 (N_5176,N_4564,N_4142);
nor U5177 (N_5177,N_4189,N_4145);
or U5178 (N_5178,N_4904,N_4277);
nor U5179 (N_5179,N_4845,N_4061);
xnor U5180 (N_5180,N_4310,N_4236);
and U5181 (N_5181,N_4547,N_4439);
and U5182 (N_5182,N_4982,N_4938);
nand U5183 (N_5183,N_4516,N_4083);
xnor U5184 (N_5184,N_4238,N_4057);
nand U5185 (N_5185,N_4256,N_4860);
or U5186 (N_5186,N_4975,N_4953);
nor U5187 (N_5187,N_4311,N_4724);
nand U5188 (N_5188,N_4981,N_4643);
nand U5189 (N_5189,N_4052,N_4706);
or U5190 (N_5190,N_4214,N_4200);
and U5191 (N_5191,N_4278,N_4542);
nor U5192 (N_5192,N_4105,N_4924);
nand U5193 (N_5193,N_4349,N_4992);
and U5194 (N_5194,N_4205,N_4645);
xor U5195 (N_5195,N_4331,N_4673);
and U5196 (N_5196,N_4771,N_4622);
xor U5197 (N_5197,N_4954,N_4047);
nor U5198 (N_5198,N_4188,N_4898);
nand U5199 (N_5199,N_4562,N_4911);
xor U5200 (N_5200,N_4147,N_4443);
nand U5201 (N_5201,N_4065,N_4795);
xnor U5202 (N_5202,N_4489,N_4496);
nor U5203 (N_5203,N_4561,N_4850);
and U5204 (N_5204,N_4965,N_4793);
or U5205 (N_5205,N_4131,N_4817);
xnor U5206 (N_5206,N_4565,N_4041);
and U5207 (N_5207,N_4786,N_4093);
nor U5208 (N_5208,N_4736,N_4138);
nand U5209 (N_5209,N_4764,N_4945);
nor U5210 (N_5210,N_4474,N_4384);
or U5211 (N_5211,N_4338,N_4720);
nand U5212 (N_5212,N_4076,N_4098);
nor U5213 (N_5213,N_4197,N_4739);
nor U5214 (N_5214,N_4647,N_4000);
or U5215 (N_5215,N_4479,N_4082);
or U5216 (N_5216,N_4090,N_4530);
and U5217 (N_5217,N_4688,N_4218);
and U5218 (N_5218,N_4760,N_4896);
xnor U5219 (N_5219,N_4529,N_4194);
nor U5220 (N_5220,N_4334,N_4753);
or U5221 (N_5221,N_4592,N_4634);
nand U5222 (N_5222,N_4068,N_4163);
nor U5223 (N_5223,N_4017,N_4070);
or U5224 (N_5224,N_4103,N_4794);
or U5225 (N_5225,N_4828,N_4971);
or U5226 (N_5226,N_4718,N_4206);
nor U5227 (N_5227,N_4963,N_4414);
nand U5228 (N_5228,N_4970,N_4452);
or U5229 (N_5229,N_4497,N_4589);
and U5230 (N_5230,N_4212,N_4108);
nand U5231 (N_5231,N_4464,N_4268);
nand U5232 (N_5232,N_4417,N_4269);
or U5233 (N_5233,N_4230,N_4578);
xnor U5234 (N_5234,N_4873,N_4974);
nor U5235 (N_5235,N_4499,N_4318);
nor U5236 (N_5236,N_4405,N_4412);
or U5237 (N_5237,N_4390,N_4327);
xnor U5238 (N_5238,N_4759,N_4262);
nor U5239 (N_5239,N_4872,N_4201);
nand U5240 (N_5240,N_4389,N_4563);
or U5241 (N_5241,N_4667,N_4876);
and U5242 (N_5242,N_4678,N_4940);
or U5243 (N_5243,N_4125,N_4601);
nor U5244 (N_5244,N_4595,N_4910);
nor U5245 (N_5245,N_4071,N_4682);
nor U5246 (N_5246,N_4697,N_4849);
nor U5247 (N_5247,N_4448,N_4111);
xnor U5248 (N_5248,N_4722,N_4434);
or U5249 (N_5249,N_4800,N_4835);
xnor U5250 (N_5250,N_4451,N_4894);
nor U5251 (N_5251,N_4006,N_4360);
or U5252 (N_5252,N_4826,N_4868);
and U5253 (N_5253,N_4329,N_4921);
xor U5254 (N_5254,N_4465,N_4853);
xor U5255 (N_5255,N_4116,N_4741);
xnor U5256 (N_5256,N_4558,N_4625);
or U5257 (N_5257,N_4064,N_4987);
nand U5258 (N_5258,N_4839,N_4220);
nor U5259 (N_5259,N_4747,N_4687);
nand U5260 (N_5260,N_4693,N_4030);
and U5261 (N_5261,N_4249,N_4088);
and U5262 (N_5262,N_4662,N_4930);
or U5263 (N_5263,N_4991,N_4984);
nor U5264 (N_5264,N_4209,N_4259);
nor U5265 (N_5265,N_4726,N_4048);
and U5266 (N_5266,N_4063,N_4049);
nor U5267 (N_5267,N_4420,N_4778);
and U5268 (N_5268,N_4926,N_4934);
nand U5269 (N_5269,N_4862,N_4594);
xor U5270 (N_5270,N_4162,N_4226);
nand U5271 (N_5271,N_4115,N_4258);
xor U5272 (N_5272,N_4708,N_4610);
nand U5273 (N_5273,N_4251,N_4297);
nand U5274 (N_5274,N_4763,N_4059);
nand U5275 (N_5275,N_4769,N_4705);
nand U5276 (N_5276,N_4091,N_4576);
and U5277 (N_5277,N_4881,N_4586);
nor U5278 (N_5278,N_4043,N_4765);
nor U5279 (N_5279,N_4557,N_4611);
nand U5280 (N_5280,N_4944,N_4445);
xor U5281 (N_5281,N_4350,N_4078);
xnor U5282 (N_5282,N_4998,N_4050);
nand U5283 (N_5283,N_4624,N_4118);
nor U5284 (N_5284,N_4210,N_4021);
xor U5285 (N_5285,N_4252,N_4792);
or U5286 (N_5286,N_4395,N_4752);
and U5287 (N_5287,N_4106,N_4323);
nand U5288 (N_5288,N_4347,N_4909);
nand U5289 (N_5289,N_4392,N_4422);
and U5290 (N_5290,N_4388,N_4507);
nand U5291 (N_5291,N_4184,N_4766);
nor U5292 (N_5292,N_4181,N_4654);
and U5293 (N_5293,N_4168,N_4999);
and U5294 (N_5294,N_4164,N_4638);
and U5295 (N_5295,N_4858,N_4572);
nor U5296 (N_5296,N_4305,N_4307);
or U5297 (N_5297,N_4867,N_4477);
and U5298 (N_5298,N_4020,N_4325);
nor U5299 (N_5299,N_4158,N_4245);
and U5300 (N_5300,N_4656,N_4637);
nand U5301 (N_5301,N_4289,N_4504);
or U5302 (N_5302,N_4740,N_4094);
and U5303 (N_5303,N_4351,N_4629);
and U5304 (N_5304,N_4880,N_4232);
nor U5305 (N_5305,N_4336,N_4374);
nand U5306 (N_5306,N_4446,N_4811);
nor U5307 (N_5307,N_4494,N_4207);
and U5308 (N_5308,N_4928,N_4636);
nand U5309 (N_5309,N_4838,N_4370);
xor U5310 (N_5310,N_4995,N_4366);
nor U5311 (N_5311,N_4707,N_4387);
xor U5312 (N_5312,N_4758,N_4727);
or U5313 (N_5313,N_4453,N_4515);
and U5314 (N_5314,N_4635,N_4646);
nor U5315 (N_5315,N_4903,N_4432);
or U5316 (N_5316,N_4135,N_4755);
xnor U5317 (N_5317,N_4545,N_4973);
and U5318 (N_5318,N_4092,N_4484);
nor U5319 (N_5319,N_4879,N_4957);
and U5320 (N_5320,N_4229,N_4885);
nor U5321 (N_5321,N_4110,N_4819);
nand U5322 (N_5322,N_4588,N_4555);
and U5323 (N_5323,N_4397,N_4519);
xor U5324 (N_5324,N_4770,N_4003);
xor U5325 (N_5325,N_4816,N_4345);
nand U5326 (N_5326,N_4608,N_4485);
nand U5327 (N_5327,N_4821,N_4614);
nand U5328 (N_5328,N_4152,N_4228);
or U5329 (N_5329,N_4217,N_4001);
and U5330 (N_5330,N_4551,N_4447);
or U5331 (N_5331,N_4402,N_4449);
nor U5332 (N_5332,N_4413,N_4096);
nor U5333 (N_5333,N_4272,N_4840);
xnor U5334 (N_5334,N_4948,N_4399);
nor U5335 (N_5335,N_4239,N_4287);
or U5336 (N_5336,N_4666,N_4469);
or U5337 (N_5337,N_4920,N_4337);
nand U5338 (N_5338,N_4790,N_4385);
nor U5339 (N_5339,N_4967,N_4640);
and U5340 (N_5340,N_4386,N_4607);
or U5341 (N_5341,N_4525,N_4187);
and U5342 (N_5342,N_4719,N_4717);
and U5343 (N_5343,N_4011,N_4224);
nand U5344 (N_5344,N_4801,N_4178);
or U5345 (N_5345,N_4120,N_4681);
and U5346 (N_5346,N_4761,N_4274);
nor U5347 (N_5347,N_4380,N_4219);
or U5348 (N_5348,N_4822,N_4890);
nor U5349 (N_5349,N_4907,N_4976);
xnor U5350 (N_5350,N_4596,N_4431);
and U5351 (N_5351,N_4365,N_4016);
nor U5352 (N_5352,N_4677,N_4915);
nand U5353 (N_5353,N_4157,N_4577);
nor U5354 (N_5354,N_4865,N_4263);
or U5355 (N_5355,N_4986,N_4377);
and U5356 (N_5356,N_4056,N_4751);
and U5357 (N_5357,N_4285,N_4491);
nand U5358 (N_5358,N_4361,N_4121);
nor U5359 (N_5359,N_4359,N_4053);
and U5360 (N_5360,N_4456,N_4627);
xnor U5361 (N_5361,N_4810,N_4657);
xor U5362 (N_5362,N_4332,N_4475);
or U5363 (N_5363,N_4013,N_4364);
nand U5364 (N_5364,N_4037,N_4134);
nor U5365 (N_5365,N_4833,N_4034);
and U5366 (N_5366,N_4756,N_4540);
nand U5367 (N_5367,N_4653,N_4712);
nor U5368 (N_5368,N_4587,N_4356);
nand U5369 (N_5369,N_4709,N_4884);
and U5370 (N_5370,N_4886,N_4582);
or U5371 (N_5371,N_4546,N_4549);
nor U5372 (N_5372,N_4339,N_4123);
xor U5373 (N_5373,N_4570,N_4127);
nor U5374 (N_5374,N_4284,N_4511);
or U5375 (N_5375,N_4787,N_4848);
and U5376 (N_5376,N_4097,N_4248);
or U5377 (N_5377,N_4411,N_4300);
nor U5378 (N_5378,N_4182,N_4757);
and U5379 (N_5379,N_4124,N_4372);
nand U5380 (N_5380,N_4132,N_4490);
or U5381 (N_5381,N_4689,N_4117);
or U5382 (N_5382,N_4566,N_4961);
nor U5383 (N_5383,N_4512,N_4069);
or U5384 (N_5384,N_4427,N_4085);
nor U5385 (N_5385,N_4996,N_4639);
nor U5386 (N_5386,N_4073,N_4363);
nand U5387 (N_5387,N_4208,N_4102);
or U5388 (N_5388,N_4933,N_4394);
nand U5389 (N_5389,N_4694,N_4522);
and U5390 (N_5390,N_4745,N_4286);
nor U5391 (N_5391,N_4202,N_4015);
and U5392 (N_5392,N_4698,N_4929);
nand U5393 (N_5393,N_4308,N_4376);
or U5394 (N_5394,N_4355,N_4172);
xor U5395 (N_5395,N_4344,N_4410);
nand U5396 (N_5396,N_4482,N_4552);
and U5397 (N_5397,N_4159,N_4620);
and U5398 (N_5398,N_4014,N_4591);
nor U5399 (N_5399,N_4832,N_4042);
nor U5400 (N_5400,N_4568,N_4309);
and U5401 (N_5401,N_4887,N_4051);
nor U5402 (N_5402,N_4978,N_4290);
nand U5403 (N_5403,N_4541,N_4341);
nand U5404 (N_5404,N_4074,N_4408);
and U5405 (N_5405,N_4153,N_4175);
nand U5406 (N_5406,N_4842,N_4914);
nand U5407 (N_5407,N_4866,N_4401);
or U5408 (N_5408,N_4983,N_4156);
and U5409 (N_5409,N_4951,N_4264);
nand U5410 (N_5410,N_4916,N_4253);
and U5411 (N_5411,N_4843,N_4234);
nor U5412 (N_5412,N_4276,N_4375);
and U5413 (N_5413,N_4130,N_4655);
nor U5414 (N_5414,N_4784,N_4854);
nor U5415 (N_5415,N_4481,N_4864);
nor U5416 (N_5416,N_4316,N_4457);
or U5417 (N_5417,N_4400,N_4648);
xnor U5418 (N_5418,N_4633,N_4623);
xnor U5419 (N_5419,N_4079,N_4166);
nand U5420 (N_5420,N_4695,N_4442);
nand U5421 (N_5421,N_4556,N_4246);
nor U5422 (N_5422,N_4038,N_4196);
or U5423 (N_5423,N_4946,N_4185);
or U5424 (N_5424,N_4573,N_4768);
or U5425 (N_5425,N_4241,N_4814);
nor U5426 (N_5426,N_4002,N_4296);
nor U5427 (N_5427,N_4721,N_4113);
nand U5428 (N_5428,N_4962,N_4321);
or U5429 (N_5429,N_4523,N_4837);
nor U5430 (N_5430,N_4075,N_4615);
nor U5431 (N_5431,N_4348,N_4470);
nor U5432 (N_5432,N_4005,N_4780);
or U5433 (N_5433,N_4901,N_4703);
xor U5434 (N_5434,N_4730,N_4874);
nand U5435 (N_5435,N_4869,N_4320);
nand U5436 (N_5436,N_4917,N_4985);
or U5437 (N_5437,N_4514,N_4878);
nor U5438 (N_5438,N_4889,N_4298);
nor U5439 (N_5439,N_4748,N_4183);
and U5440 (N_5440,N_4877,N_4133);
xor U5441 (N_5441,N_4095,N_4028);
nor U5442 (N_5442,N_4173,N_4750);
nand U5443 (N_5443,N_4528,N_4114);
and U5444 (N_5444,N_4980,N_4649);
nor U5445 (N_5445,N_4480,N_4161);
and U5446 (N_5446,N_4583,N_4009);
nand U5447 (N_5447,N_4791,N_4949);
or U5448 (N_5448,N_4960,N_4554);
nand U5449 (N_5449,N_4997,N_4190);
nand U5450 (N_5450,N_4613,N_4450);
or U5451 (N_5451,N_4418,N_4905);
xnor U5452 (N_5452,N_4806,N_4844);
nand U5453 (N_5453,N_4010,N_4506);
and U5454 (N_5454,N_4174,N_4019);
nor U5455 (N_5455,N_4660,N_4382);
or U5456 (N_5456,N_4282,N_4266);
xor U5457 (N_5457,N_4454,N_4825);
nand U5458 (N_5458,N_4033,N_4683);
nor U5459 (N_5459,N_4424,N_4122);
nand U5460 (N_5460,N_4488,N_4820);
nand U5461 (N_5461,N_4691,N_4650);
nor U5462 (N_5462,N_4988,N_4737);
or U5463 (N_5463,N_4531,N_4799);
nor U5464 (N_5464,N_4685,N_4815);
nand U5465 (N_5465,N_4104,N_4406);
nand U5466 (N_5466,N_4304,N_4543);
nand U5467 (N_5467,N_4734,N_4550);
nor U5468 (N_5468,N_4379,N_4462);
nand U5469 (N_5469,N_4802,N_4371);
nand U5470 (N_5470,N_4809,N_4198);
and U5471 (N_5471,N_4299,N_4584);
nor U5472 (N_5472,N_4170,N_4222);
or U5473 (N_5473,N_4358,N_4180);
or U5474 (N_5474,N_4444,N_4139);
nor U5475 (N_5475,N_4080,N_4281);
and U5476 (N_5476,N_4493,N_4711);
or U5477 (N_5477,N_4644,N_4559);
and U5478 (N_5478,N_4544,N_4235);
nand U5479 (N_5479,N_4882,N_4383);
and U5480 (N_5480,N_4834,N_4661);
nor U5481 (N_5481,N_4723,N_4373);
nor U5482 (N_5482,N_4908,N_4521);
and U5483 (N_5483,N_4743,N_4569);
nor U5484 (N_5484,N_4897,N_4704);
nand U5485 (N_5485,N_4067,N_4732);
nor U5486 (N_5486,N_4160,N_4847);
nor U5487 (N_5487,N_4191,N_4609);
and U5488 (N_5488,N_4827,N_4328);
or U5489 (N_5489,N_4680,N_4343);
and U5490 (N_5490,N_4319,N_4403);
and U5491 (N_5491,N_4580,N_4900);
and U5492 (N_5492,N_4671,N_4353);
nand U5493 (N_5493,N_4381,N_4404);
nor U5494 (N_5494,N_4126,N_4179);
nand U5495 (N_5495,N_4204,N_4335);
and U5496 (N_5496,N_4215,N_4112);
or U5497 (N_5497,N_4036,N_4267);
nand U5498 (N_5498,N_4326,N_4628);
nor U5499 (N_5499,N_4742,N_4498);
or U5500 (N_5500,N_4267,N_4683);
and U5501 (N_5501,N_4133,N_4827);
or U5502 (N_5502,N_4211,N_4819);
and U5503 (N_5503,N_4285,N_4474);
and U5504 (N_5504,N_4718,N_4816);
nand U5505 (N_5505,N_4588,N_4886);
nand U5506 (N_5506,N_4364,N_4577);
nor U5507 (N_5507,N_4448,N_4702);
nand U5508 (N_5508,N_4673,N_4641);
xor U5509 (N_5509,N_4754,N_4513);
and U5510 (N_5510,N_4293,N_4367);
and U5511 (N_5511,N_4205,N_4867);
and U5512 (N_5512,N_4805,N_4902);
and U5513 (N_5513,N_4564,N_4830);
and U5514 (N_5514,N_4888,N_4512);
and U5515 (N_5515,N_4326,N_4923);
and U5516 (N_5516,N_4196,N_4125);
nor U5517 (N_5517,N_4104,N_4459);
nand U5518 (N_5518,N_4856,N_4589);
nand U5519 (N_5519,N_4178,N_4783);
nor U5520 (N_5520,N_4505,N_4453);
nor U5521 (N_5521,N_4961,N_4172);
xor U5522 (N_5522,N_4295,N_4979);
or U5523 (N_5523,N_4433,N_4735);
and U5524 (N_5524,N_4806,N_4949);
nor U5525 (N_5525,N_4873,N_4685);
nand U5526 (N_5526,N_4173,N_4769);
or U5527 (N_5527,N_4451,N_4060);
nand U5528 (N_5528,N_4520,N_4996);
or U5529 (N_5529,N_4115,N_4571);
and U5530 (N_5530,N_4081,N_4435);
or U5531 (N_5531,N_4180,N_4651);
xnor U5532 (N_5532,N_4355,N_4056);
and U5533 (N_5533,N_4759,N_4178);
or U5534 (N_5534,N_4771,N_4133);
xor U5535 (N_5535,N_4878,N_4331);
xnor U5536 (N_5536,N_4242,N_4753);
or U5537 (N_5537,N_4057,N_4424);
nor U5538 (N_5538,N_4058,N_4568);
nand U5539 (N_5539,N_4329,N_4960);
and U5540 (N_5540,N_4782,N_4108);
nand U5541 (N_5541,N_4926,N_4909);
or U5542 (N_5542,N_4055,N_4862);
nor U5543 (N_5543,N_4395,N_4501);
nor U5544 (N_5544,N_4733,N_4515);
and U5545 (N_5545,N_4421,N_4527);
or U5546 (N_5546,N_4288,N_4884);
or U5547 (N_5547,N_4141,N_4508);
nor U5548 (N_5548,N_4242,N_4857);
and U5549 (N_5549,N_4922,N_4369);
or U5550 (N_5550,N_4867,N_4154);
xnor U5551 (N_5551,N_4482,N_4066);
and U5552 (N_5552,N_4608,N_4057);
xnor U5553 (N_5553,N_4535,N_4039);
or U5554 (N_5554,N_4048,N_4775);
and U5555 (N_5555,N_4323,N_4779);
or U5556 (N_5556,N_4546,N_4611);
xnor U5557 (N_5557,N_4677,N_4070);
and U5558 (N_5558,N_4211,N_4857);
and U5559 (N_5559,N_4654,N_4144);
and U5560 (N_5560,N_4895,N_4268);
or U5561 (N_5561,N_4862,N_4835);
and U5562 (N_5562,N_4993,N_4052);
nor U5563 (N_5563,N_4952,N_4364);
nand U5564 (N_5564,N_4243,N_4562);
nor U5565 (N_5565,N_4389,N_4833);
or U5566 (N_5566,N_4507,N_4172);
and U5567 (N_5567,N_4217,N_4209);
nand U5568 (N_5568,N_4471,N_4910);
nor U5569 (N_5569,N_4176,N_4425);
and U5570 (N_5570,N_4598,N_4891);
xnor U5571 (N_5571,N_4878,N_4052);
nor U5572 (N_5572,N_4511,N_4824);
nand U5573 (N_5573,N_4420,N_4696);
or U5574 (N_5574,N_4625,N_4756);
or U5575 (N_5575,N_4334,N_4516);
nor U5576 (N_5576,N_4112,N_4607);
or U5577 (N_5577,N_4643,N_4145);
or U5578 (N_5578,N_4348,N_4253);
nor U5579 (N_5579,N_4385,N_4408);
and U5580 (N_5580,N_4879,N_4055);
and U5581 (N_5581,N_4532,N_4373);
and U5582 (N_5582,N_4298,N_4644);
or U5583 (N_5583,N_4499,N_4530);
or U5584 (N_5584,N_4170,N_4620);
or U5585 (N_5585,N_4681,N_4520);
nand U5586 (N_5586,N_4474,N_4620);
xor U5587 (N_5587,N_4538,N_4482);
or U5588 (N_5588,N_4255,N_4546);
nand U5589 (N_5589,N_4313,N_4006);
nor U5590 (N_5590,N_4818,N_4247);
and U5591 (N_5591,N_4118,N_4433);
or U5592 (N_5592,N_4573,N_4286);
nor U5593 (N_5593,N_4509,N_4703);
nor U5594 (N_5594,N_4682,N_4976);
or U5595 (N_5595,N_4181,N_4258);
and U5596 (N_5596,N_4390,N_4571);
nor U5597 (N_5597,N_4004,N_4278);
nor U5598 (N_5598,N_4983,N_4261);
nand U5599 (N_5599,N_4841,N_4196);
nand U5600 (N_5600,N_4092,N_4268);
xor U5601 (N_5601,N_4855,N_4112);
nand U5602 (N_5602,N_4464,N_4511);
nor U5603 (N_5603,N_4691,N_4974);
nand U5604 (N_5604,N_4772,N_4122);
nor U5605 (N_5605,N_4537,N_4604);
and U5606 (N_5606,N_4948,N_4123);
or U5607 (N_5607,N_4396,N_4260);
and U5608 (N_5608,N_4203,N_4803);
and U5609 (N_5609,N_4039,N_4568);
or U5610 (N_5610,N_4855,N_4788);
or U5611 (N_5611,N_4007,N_4037);
and U5612 (N_5612,N_4192,N_4988);
nand U5613 (N_5613,N_4058,N_4274);
xnor U5614 (N_5614,N_4680,N_4670);
nand U5615 (N_5615,N_4357,N_4242);
nand U5616 (N_5616,N_4014,N_4420);
or U5617 (N_5617,N_4670,N_4054);
xnor U5618 (N_5618,N_4757,N_4056);
nor U5619 (N_5619,N_4785,N_4202);
or U5620 (N_5620,N_4532,N_4351);
nor U5621 (N_5621,N_4009,N_4291);
nor U5622 (N_5622,N_4350,N_4962);
nand U5623 (N_5623,N_4490,N_4588);
nor U5624 (N_5624,N_4250,N_4318);
or U5625 (N_5625,N_4498,N_4690);
and U5626 (N_5626,N_4478,N_4821);
nor U5627 (N_5627,N_4500,N_4006);
xnor U5628 (N_5628,N_4291,N_4197);
xor U5629 (N_5629,N_4334,N_4037);
or U5630 (N_5630,N_4428,N_4449);
and U5631 (N_5631,N_4775,N_4041);
nand U5632 (N_5632,N_4345,N_4418);
xnor U5633 (N_5633,N_4865,N_4475);
nand U5634 (N_5634,N_4216,N_4860);
nand U5635 (N_5635,N_4278,N_4273);
xnor U5636 (N_5636,N_4986,N_4856);
and U5637 (N_5637,N_4232,N_4212);
xor U5638 (N_5638,N_4112,N_4021);
nand U5639 (N_5639,N_4300,N_4867);
xnor U5640 (N_5640,N_4178,N_4620);
or U5641 (N_5641,N_4776,N_4668);
nand U5642 (N_5642,N_4341,N_4431);
and U5643 (N_5643,N_4111,N_4906);
or U5644 (N_5644,N_4259,N_4572);
and U5645 (N_5645,N_4247,N_4064);
or U5646 (N_5646,N_4934,N_4319);
xnor U5647 (N_5647,N_4299,N_4297);
or U5648 (N_5648,N_4439,N_4737);
and U5649 (N_5649,N_4981,N_4205);
xor U5650 (N_5650,N_4707,N_4909);
and U5651 (N_5651,N_4988,N_4402);
nor U5652 (N_5652,N_4462,N_4941);
and U5653 (N_5653,N_4944,N_4003);
or U5654 (N_5654,N_4387,N_4004);
xor U5655 (N_5655,N_4810,N_4644);
and U5656 (N_5656,N_4435,N_4345);
nor U5657 (N_5657,N_4613,N_4318);
and U5658 (N_5658,N_4272,N_4430);
or U5659 (N_5659,N_4044,N_4412);
or U5660 (N_5660,N_4415,N_4060);
and U5661 (N_5661,N_4882,N_4182);
or U5662 (N_5662,N_4014,N_4027);
and U5663 (N_5663,N_4298,N_4963);
or U5664 (N_5664,N_4697,N_4580);
and U5665 (N_5665,N_4149,N_4360);
nand U5666 (N_5666,N_4273,N_4464);
xnor U5667 (N_5667,N_4266,N_4605);
or U5668 (N_5668,N_4517,N_4729);
nand U5669 (N_5669,N_4770,N_4561);
and U5670 (N_5670,N_4124,N_4218);
and U5671 (N_5671,N_4652,N_4679);
nor U5672 (N_5672,N_4069,N_4148);
and U5673 (N_5673,N_4019,N_4630);
nor U5674 (N_5674,N_4591,N_4208);
and U5675 (N_5675,N_4614,N_4658);
nand U5676 (N_5676,N_4987,N_4167);
xnor U5677 (N_5677,N_4167,N_4893);
nor U5678 (N_5678,N_4402,N_4475);
xnor U5679 (N_5679,N_4439,N_4444);
or U5680 (N_5680,N_4489,N_4349);
nor U5681 (N_5681,N_4385,N_4134);
nor U5682 (N_5682,N_4556,N_4824);
or U5683 (N_5683,N_4542,N_4339);
or U5684 (N_5684,N_4601,N_4395);
nand U5685 (N_5685,N_4811,N_4671);
nand U5686 (N_5686,N_4206,N_4979);
or U5687 (N_5687,N_4841,N_4481);
and U5688 (N_5688,N_4176,N_4875);
nor U5689 (N_5689,N_4902,N_4631);
xnor U5690 (N_5690,N_4049,N_4082);
nand U5691 (N_5691,N_4096,N_4736);
nor U5692 (N_5692,N_4077,N_4988);
nor U5693 (N_5693,N_4682,N_4655);
and U5694 (N_5694,N_4718,N_4679);
or U5695 (N_5695,N_4654,N_4165);
and U5696 (N_5696,N_4953,N_4611);
nor U5697 (N_5697,N_4211,N_4082);
or U5698 (N_5698,N_4515,N_4584);
xnor U5699 (N_5699,N_4747,N_4001);
nand U5700 (N_5700,N_4142,N_4690);
xnor U5701 (N_5701,N_4365,N_4677);
or U5702 (N_5702,N_4992,N_4746);
nor U5703 (N_5703,N_4681,N_4037);
nand U5704 (N_5704,N_4564,N_4827);
nor U5705 (N_5705,N_4979,N_4251);
or U5706 (N_5706,N_4086,N_4804);
or U5707 (N_5707,N_4898,N_4057);
nand U5708 (N_5708,N_4184,N_4912);
nand U5709 (N_5709,N_4914,N_4653);
or U5710 (N_5710,N_4286,N_4739);
nor U5711 (N_5711,N_4044,N_4941);
nand U5712 (N_5712,N_4561,N_4702);
and U5713 (N_5713,N_4887,N_4609);
or U5714 (N_5714,N_4059,N_4076);
nor U5715 (N_5715,N_4228,N_4000);
xnor U5716 (N_5716,N_4368,N_4208);
xor U5717 (N_5717,N_4101,N_4483);
nand U5718 (N_5718,N_4126,N_4148);
and U5719 (N_5719,N_4216,N_4742);
or U5720 (N_5720,N_4679,N_4917);
xnor U5721 (N_5721,N_4252,N_4152);
and U5722 (N_5722,N_4938,N_4265);
nor U5723 (N_5723,N_4389,N_4035);
nand U5724 (N_5724,N_4463,N_4103);
nand U5725 (N_5725,N_4539,N_4315);
and U5726 (N_5726,N_4257,N_4008);
nand U5727 (N_5727,N_4764,N_4136);
xnor U5728 (N_5728,N_4446,N_4188);
or U5729 (N_5729,N_4542,N_4437);
nor U5730 (N_5730,N_4935,N_4291);
or U5731 (N_5731,N_4671,N_4042);
nor U5732 (N_5732,N_4174,N_4719);
and U5733 (N_5733,N_4573,N_4812);
or U5734 (N_5734,N_4491,N_4776);
nand U5735 (N_5735,N_4912,N_4068);
nor U5736 (N_5736,N_4220,N_4976);
nor U5737 (N_5737,N_4511,N_4050);
or U5738 (N_5738,N_4095,N_4988);
nand U5739 (N_5739,N_4395,N_4088);
xnor U5740 (N_5740,N_4419,N_4407);
nand U5741 (N_5741,N_4729,N_4565);
nand U5742 (N_5742,N_4848,N_4327);
nand U5743 (N_5743,N_4208,N_4552);
and U5744 (N_5744,N_4497,N_4421);
xor U5745 (N_5745,N_4304,N_4504);
xnor U5746 (N_5746,N_4515,N_4451);
nor U5747 (N_5747,N_4798,N_4836);
xor U5748 (N_5748,N_4765,N_4788);
nand U5749 (N_5749,N_4502,N_4179);
nor U5750 (N_5750,N_4189,N_4423);
or U5751 (N_5751,N_4581,N_4570);
and U5752 (N_5752,N_4364,N_4763);
nand U5753 (N_5753,N_4640,N_4679);
or U5754 (N_5754,N_4050,N_4512);
nor U5755 (N_5755,N_4753,N_4718);
xor U5756 (N_5756,N_4573,N_4039);
nand U5757 (N_5757,N_4710,N_4019);
or U5758 (N_5758,N_4314,N_4339);
nand U5759 (N_5759,N_4602,N_4361);
nand U5760 (N_5760,N_4011,N_4036);
nand U5761 (N_5761,N_4618,N_4583);
nor U5762 (N_5762,N_4682,N_4605);
nor U5763 (N_5763,N_4880,N_4292);
nor U5764 (N_5764,N_4830,N_4693);
xnor U5765 (N_5765,N_4588,N_4384);
xor U5766 (N_5766,N_4374,N_4521);
nor U5767 (N_5767,N_4980,N_4361);
and U5768 (N_5768,N_4974,N_4116);
xor U5769 (N_5769,N_4585,N_4543);
and U5770 (N_5770,N_4816,N_4078);
xor U5771 (N_5771,N_4559,N_4921);
xor U5772 (N_5772,N_4136,N_4847);
nor U5773 (N_5773,N_4209,N_4920);
or U5774 (N_5774,N_4403,N_4884);
nand U5775 (N_5775,N_4850,N_4798);
nand U5776 (N_5776,N_4084,N_4030);
or U5777 (N_5777,N_4721,N_4414);
or U5778 (N_5778,N_4862,N_4316);
xnor U5779 (N_5779,N_4393,N_4068);
and U5780 (N_5780,N_4049,N_4729);
and U5781 (N_5781,N_4815,N_4010);
or U5782 (N_5782,N_4321,N_4486);
or U5783 (N_5783,N_4061,N_4642);
nand U5784 (N_5784,N_4044,N_4437);
and U5785 (N_5785,N_4452,N_4223);
or U5786 (N_5786,N_4583,N_4933);
and U5787 (N_5787,N_4438,N_4786);
and U5788 (N_5788,N_4838,N_4224);
nor U5789 (N_5789,N_4421,N_4275);
nor U5790 (N_5790,N_4300,N_4523);
nor U5791 (N_5791,N_4897,N_4635);
nand U5792 (N_5792,N_4178,N_4853);
nor U5793 (N_5793,N_4899,N_4788);
and U5794 (N_5794,N_4549,N_4496);
and U5795 (N_5795,N_4573,N_4833);
nor U5796 (N_5796,N_4671,N_4842);
nand U5797 (N_5797,N_4292,N_4590);
nor U5798 (N_5798,N_4692,N_4139);
nor U5799 (N_5799,N_4599,N_4585);
or U5800 (N_5800,N_4037,N_4194);
nand U5801 (N_5801,N_4463,N_4621);
nand U5802 (N_5802,N_4680,N_4548);
nand U5803 (N_5803,N_4021,N_4497);
nand U5804 (N_5804,N_4295,N_4015);
nor U5805 (N_5805,N_4815,N_4089);
nor U5806 (N_5806,N_4854,N_4473);
nor U5807 (N_5807,N_4411,N_4408);
nand U5808 (N_5808,N_4510,N_4239);
or U5809 (N_5809,N_4909,N_4236);
nor U5810 (N_5810,N_4268,N_4659);
or U5811 (N_5811,N_4258,N_4016);
nand U5812 (N_5812,N_4389,N_4929);
nor U5813 (N_5813,N_4098,N_4250);
or U5814 (N_5814,N_4580,N_4556);
nand U5815 (N_5815,N_4257,N_4175);
nor U5816 (N_5816,N_4964,N_4178);
and U5817 (N_5817,N_4761,N_4970);
nand U5818 (N_5818,N_4568,N_4856);
xor U5819 (N_5819,N_4759,N_4825);
and U5820 (N_5820,N_4274,N_4014);
nand U5821 (N_5821,N_4261,N_4329);
or U5822 (N_5822,N_4065,N_4730);
nor U5823 (N_5823,N_4358,N_4079);
and U5824 (N_5824,N_4400,N_4645);
and U5825 (N_5825,N_4191,N_4006);
nand U5826 (N_5826,N_4661,N_4954);
nand U5827 (N_5827,N_4687,N_4865);
and U5828 (N_5828,N_4269,N_4952);
and U5829 (N_5829,N_4129,N_4404);
nor U5830 (N_5830,N_4304,N_4282);
xor U5831 (N_5831,N_4302,N_4953);
xor U5832 (N_5832,N_4014,N_4390);
and U5833 (N_5833,N_4714,N_4814);
and U5834 (N_5834,N_4552,N_4788);
nand U5835 (N_5835,N_4369,N_4943);
nand U5836 (N_5836,N_4965,N_4174);
or U5837 (N_5837,N_4895,N_4606);
nand U5838 (N_5838,N_4298,N_4106);
and U5839 (N_5839,N_4307,N_4310);
and U5840 (N_5840,N_4301,N_4474);
or U5841 (N_5841,N_4017,N_4158);
and U5842 (N_5842,N_4315,N_4699);
or U5843 (N_5843,N_4314,N_4073);
nand U5844 (N_5844,N_4581,N_4339);
nor U5845 (N_5845,N_4433,N_4361);
nor U5846 (N_5846,N_4577,N_4865);
or U5847 (N_5847,N_4433,N_4291);
or U5848 (N_5848,N_4065,N_4072);
nor U5849 (N_5849,N_4169,N_4581);
nand U5850 (N_5850,N_4349,N_4776);
nor U5851 (N_5851,N_4799,N_4645);
and U5852 (N_5852,N_4957,N_4943);
nor U5853 (N_5853,N_4321,N_4109);
or U5854 (N_5854,N_4698,N_4159);
and U5855 (N_5855,N_4544,N_4182);
or U5856 (N_5856,N_4935,N_4613);
nor U5857 (N_5857,N_4001,N_4879);
nor U5858 (N_5858,N_4875,N_4981);
or U5859 (N_5859,N_4925,N_4362);
nand U5860 (N_5860,N_4482,N_4585);
and U5861 (N_5861,N_4663,N_4715);
and U5862 (N_5862,N_4971,N_4153);
nand U5863 (N_5863,N_4554,N_4683);
nand U5864 (N_5864,N_4343,N_4250);
and U5865 (N_5865,N_4675,N_4659);
or U5866 (N_5866,N_4964,N_4328);
nand U5867 (N_5867,N_4023,N_4134);
or U5868 (N_5868,N_4303,N_4481);
nand U5869 (N_5869,N_4145,N_4152);
or U5870 (N_5870,N_4680,N_4787);
or U5871 (N_5871,N_4904,N_4415);
and U5872 (N_5872,N_4318,N_4905);
and U5873 (N_5873,N_4072,N_4293);
xnor U5874 (N_5874,N_4864,N_4621);
xnor U5875 (N_5875,N_4446,N_4357);
or U5876 (N_5876,N_4041,N_4653);
or U5877 (N_5877,N_4002,N_4865);
and U5878 (N_5878,N_4740,N_4628);
xor U5879 (N_5879,N_4289,N_4399);
or U5880 (N_5880,N_4614,N_4404);
and U5881 (N_5881,N_4951,N_4547);
nor U5882 (N_5882,N_4537,N_4952);
nor U5883 (N_5883,N_4001,N_4032);
nor U5884 (N_5884,N_4941,N_4566);
nand U5885 (N_5885,N_4886,N_4570);
and U5886 (N_5886,N_4670,N_4222);
nor U5887 (N_5887,N_4433,N_4631);
nand U5888 (N_5888,N_4952,N_4408);
and U5889 (N_5889,N_4021,N_4979);
or U5890 (N_5890,N_4897,N_4479);
nor U5891 (N_5891,N_4144,N_4862);
and U5892 (N_5892,N_4030,N_4174);
nor U5893 (N_5893,N_4807,N_4619);
nand U5894 (N_5894,N_4618,N_4869);
nand U5895 (N_5895,N_4273,N_4939);
nand U5896 (N_5896,N_4628,N_4373);
xnor U5897 (N_5897,N_4250,N_4446);
or U5898 (N_5898,N_4205,N_4585);
nand U5899 (N_5899,N_4977,N_4583);
nor U5900 (N_5900,N_4934,N_4200);
nor U5901 (N_5901,N_4682,N_4093);
nand U5902 (N_5902,N_4443,N_4087);
or U5903 (N_5903,N_4518,N_4622);
and U5904 (N_5904,N_4497,N_4355);
and U5905 (N_5905,N_4042,N_4842);
xnor U5906 (N_5906,N_4465,N_4171);
nor U5907 (N_5907,N_4112,N_4311);
xnor U5908 (N_5908,N_4293,N_4039);
and U5909 (N_5909,N_4774,N_4173);
and U5910 (N_5910,N_4888,N_4116);
nor U5911 (N_5911,N_4338,N_4246);
and U5912 (N_5912,N_4906,N_4903);
and U5913 (N_5913,N_4594,N_4271);
nor U5914 (N_5914,N_4204,N_4804);
xor U5915 (N_5915,N_4688,N_4999);
and U5916 (N_5916,N_4449,N_4742);
nor U5917 (N_5917,N_4013,N_4287);
nand U5918 (N_5918,N_4591,N_4402);
nand U5919 (N_5919,N_4204,N_4764);
xor U5920 (N_5920,N_4279,N_4203);
nor U5921 (N_5921,N_4384,N_4424);
or U5922 (N_5922,N_4821,N_4382);
nor U5923 (N_5923,N_4494,N_4239);
and U5924 (N_5924,N_4478,N_4956);
nand U5925 (N_5925,N_4865,N_4552);
nand U5926 (N_5926,N_4144,N_4360);
and U5927 (N_5927,N_4316,N_4431);
or U5928 (N_5928,N_4906,N_4697);
and U5929 (N_5929,N_4146,N_4372);
and U5930 (N_5930,N_4051,N_4573);
or U5931 (N_5931,N_4311,N_4141);
nand U5932 (N_5932,N_4533,N_4810);
nand U5933 (N_5933,N_4485,N_4932);
and U5934 (N_5934,N_4621,N_4587);
and U5935 (N_5935,N_4947,N_4661);
nand U5936 (N_5936,N_4850,N_4550);
xor U5937 (N_5937,N_4710,N_4058);
nor U5938 (N_5938,N_4322,N_4406);
or U5939 (N_5939,N_4104,N_4951);
xnor U5940 (N_5940,N_4087,N_4974);
nand U5941 (N_5941,N_4260,N_4617);
nand U5942 (N_5942,N_4198,N_4360);
and U5943 (N_5943,N_4948,N_4744);
xor U5944 (N_5944,N_4926,N_4081);
nor U5945 (N_5945,N_4465,N_4997);
nand U5946 (N_5946,N_4033,N_4532);
and U5947 (N_5947,N_4255,N_4928);
or U5948 (N_5948,N_4236,N_4999);
nand U5949 (N_5949,N_4291,N_4881);
nor U5950 (N_5950,N_4372,N_4312);
and U5951 (N_5951,N_4973,N_4586);
nor U5952 (N_5952,N_4971,N_4447);
nor U5953 (N_5953,N_4668,N_4745);
and U5954 (N_5954,N_4311,N_4424);
or U5955 (N_5955,N_4525,N_4728);
or U5956 (N_5956,N_4635,N_4226);
nor U5957 (N_5957,N_4480,N_4956);
and U5958 (N_5958,N_4464,N_4535);
or U5959 (N_5959,N_4479,N_4586);
or U5960 (N_5960,N_4719,N_4907);
nor U5961 (N_5961,N_4206,N_4883);
nor U5962 (N_5962,N_4545,N_4069);
xor U5963 (N_5963,N_4963,N_4991);
or U5964 (N_5964,N_4319,N_4909);
or U5965 (N_5965,N_4987,N_4479);
nand U5966 (N_5966,N_4675,N_4375);
nand U5967 (N_5967,N_4981,N_4851);
nor U5968 (N_5968,N_4710,N_4540);
nor U5969 (N_5969,N_4358,N_4969);
or U5970 (N_5970,N_4710,N_4373);
nor U5971 (N_5971,N_4721,N_4971);
xor U5972 (N_5972,N_4391,N_4680);
nand U5973 (N_5973,N_4970,N_4218);
xor U5974 (N_5974,N_4486,N_4579);
or U5975 (N_5975,N_4171,N_4463);
or U5976 (N_5976,N_4332,N_4913);
nor U5977 (N_5977,N_4720,N_4044);
xor U5978 (N_5978,N_4785,N_4231);
or U5979 (N_5979,N_4740,N_4447);
nand U5980 (N_5980,N_4261,N_4309);
or U5981 (N_5981,N_4386,N_4075);
nor U5982 (N_5982,N_4517,N_4977);
and U5983 (N_5983,N_4991,N_4472);
nor U5984 (N_5984,N_4561,N_4546);
and U5985 (N_5985,N_4164,N_4769);
nor U5986 (N_5986,N_4570,N_4610);
xor U5987 (N_5987,N_4446,N_4286);
nand U5988 (N_5988,N_4179,N_4592);
nand U5989 (N_5989,N_4626,N_4085);
nand U5990 (N_5990,N_4207,N_4225);
nand U5991 (N_5991,N_4267,N_4519);
and U5992 (N_5992,N_4153,N_4392);
or U5993 (N_5993,N_4519,N_4253);
or U5994 (N_5994,N_4432,N_4224);
or U5995 (N_5995,N_4691,N_4512);
nand U5996 (N_5996,N_4703,N_4829);
nand U5997 (N_5997,N_4592,N_4213);
or U5998 (N_5998,N_4626,N_4317);
and U5999 (N_5999,N_4121,N_4546);
or U6000 (N_6000,N_5692,N_5397);
nor U6001 (N_6001,N_5388,N_5502);
and U6002 (N_6002,N_5578,N_5566);
nand U6003 (N_6003,N_5574,N_5365);
or U6004 (N_6004,N_5894,N_5945);
nor U6005 (N_6005,N_5083,N_5164);
nor U6006 (N_6006,N_5102,N_5690);
and U6007 (N_6007,N_5707,N_5678);
nand U6008 (N_6008,N_5295,N_5022);
nor U6009 (N_6009,N_5158,N_5637);
nor U6010 (N_6010,N_5401,N_5227);
nor U6011 (N_6011,N_5186,N_5673);
or U6012 (N_6012,N_5434,N_5374);
xnor U6013 (N_6013,N_5344,N_5988);
nor U6014 (N_6014,N_5127,N_5252);
and U6015 (N_6015,N_5904,N_5551);
nand U6016 (N_6016,N_5340,N_5552);
xnor U6017 (N_6017,N_5855,N_5954);
nor U6018 (N_6018,N_5483,N_5949);
nor U6019 (N_6019,N_5579,N_5752);
xnor U6020 (N_6020,N_5473,N_5203);
xor U6021 (N_6021,N_5644,N_5605);
nor U6022 (N_6022,N_5096,N_5646);
nand U6023 (N_6023,N_5947,N_5216);
nor U6024 (N_6024,N_5970,N_5492);
nand U6025 (N_6025,N_5071,N_5940);
or U6026 (N_6026,N_5178,N_5453);
nand U6027 (N_6027,N_5895,N_5980);
nor U6028 (N_6028,N_5070,N_5156);
xor U6029 (N_6029,N_5586,N_5345);
and U6030 (N_6030,N_5284,N_5881);
nor U6031 (N_6031,N_5769,N_5181);
or U6032 (N_6032,N_5258,N_5132);
and U6033 (N_6033,N_5400,N_5779);
or U6034 (N_6034,N_5763,N_5982);
nand U6035 (N_6035,N_5405,N_5268);
nand U6036 (N_6036,N_5333,N_5890);
xor U6037 (N_6037,N_5470,N_5963);
and U6038 (N_6038,N_5974,N_5997);
and U6039 (N_6039,N_5038,N_5462);
xnor U6040 (N_6040,N_5231,N_5078);
or U6041 (N_6041,N_5817,N_5170);
or U6042 (N_6042,N_5802,N_5047);
and U6043 (N_6043,N_5282,N_5680);
nor U6044 (N_6044,N_5564,N_5745);
and U6045 (N_6045,N_5059,N_5439);
and U6046 (N_6046,N_5206,N_5064);
nor U6047 (N_6047,N_5917,N_5384);
nor U6048 (N_6048,N_5557,N_5264);
nand U6049 (N_6049,N_5792,N_5062);
nor U6050 (N_6050,N_5674,N_5145);
xor U6051 (N_6051,N_5539,N_5836);
and U6052 (N_6052,N_5577,N_5977);
and U6053 (N_6053,N_5202,N_5727);
nor U6054 (N_6054,N_5677,N_5919);
and U6055 (N_6055,N_5499,N_5100);
or U6056 (N_6056,N_5920,N_5985);
xnor U6057 (N_6057,N_5060,N_5438);
nand U6058 (N_6058,N_5337,N_5278);
or U6059 (N_6059,N_5590,N_5274);
nor U6060 (N_6060,N_5850,N_5781);
xor U6061 (N_6061,N_5251,N_5714);
nor U6062 (N_6062,N_5343,N_5689);
nor U6063 (N_6063,N_5010,N_5839);
and U6064 (N_6064,N_5444,N_5381);
nand U6065 (N_6065,N_5654,N_5331);
nor U6066 (N_6066,N_5632,N_5230);
and U6067 (N_6067,N_5496,N_5994);
or U6068 (N_6068,N_5554,N_5139);
and U6069 (N_6069,N_5751,N_5157);
nand U6070 (N_6070,N_5187,N_5131);
nor U6071 (N_6071,N_5531,N_5615);
nor U6072 (N_6072,N_5873,N_5511);
and U6073 (N_6073,N_5032,N_5332);
and U6074 (N_6074,N_5767,N_5854);
and U6075 (N_6075,N_5599,N_5978);
nand U6076 (N_6076,N_5141,N_5961);
nor U6077 (N_6077,N_5744,N_5236);
or U6078 (N_6078,N_5076,N_5087);
nand U6079 (N_6079,N_5442,N_5428);
xnor U6080 (N_6080,N_5510,N_5056);
nor U6081 (N_6081,N_5080,N_5199);
nand U6082 (N_6082,N_5097,N_5778);
or U6083 (N_6083,N_5204,N_5923);
nor U6084 (N_6084,N_5451,N_5645);
or U6085 (N_6085,N_5772,N_5477);
nor U6086 (N_6086,N_5706,N_5596);
and U6087 (N_6087,N_5372,N_5447);
xor U6088 (N_6088,N_5184,N_5570);
nand U6089 (N_6089,N_5541,N_5475);
nor U6090 (N_6090,N_5800,N_5804);
nor U6091 (N_6091,N_5829,N_5696);
and U6092 (N_6092,N_5350,N_5443);
and U6093 (N_6093,N_5816,N_5602);
nand U6094 (N_6094,N_5063,N_5369);
nor U6095 (N_6095,N_5305,N_5731);
nand U6096 (N_6096,N_5247,N_5207);
and U6097 (N_6097,N_5611,N_5858);
nor U6098 (N_6098,N_5323,N_5346);
nand U6099 (N_6099,N_5082,N_5105);
nand U6100 (N_6100,N_5983,N_5277);
nor U6101 (N_6101,N_5889,N_5315);
or U6102 (N_6102,N_5634,N_5065);
and U6103 (N_6103,N_5360,N_5279);
or U6104 (N_6104,N_5281,N_5094);
xnor U6105 (N_6105,N_5630,N_5776);
nand U6106 (N_6106,N_5042,N_5747);
xor U6107 (N_6107,N_5553,N_5385);
nand U6108 (N_6108,N_5999,N_5521);
nand U6109 (N_6109,N_5799,N_5973);
and U6110 (N_6110,N_5777,N_5716);
and U6111 (N_6111,N_5414,N_5148);
or U6112 (N_6112,N_5253,N_5780);
or U6113 (N_6113,N_5943,N_5785);
nor U6114 (N_6114,N_5418,N_5756);
nor U6115 (N_6115,N_5652,N_5831);
nand U6116 (N_6116,N_5957,N_5807);
nor U6117 (N_6117,N_5612,N_5500);
nand U6118 (N_6118,N_5921,N_5594);
nor U6119 (N_6119,N_5250,N_5812);
nand U6120 (N_6120,N_5995,N_5606);
xor U6121 (N_6121,N_5840,N_5754);
nand U6122 (N_6122,N_5495,N_5497);
nand U6123 (N_6123,N_5432,N_5725);
nor U6124 (N_6124,N_5006,N_5240);
nand U6125 (N_6125,N_5618,N_5458);
nand U6126 (N_6126,N_5710,N_5522);
nand U6127 (N_6127,N_5998,N_5478);
nor U6128 (N_6128,N_5121,N_5694);
or U6129 (N_6129,N_5433,N_5249);
and U6130 (N_6130,N_5311,N_5712);
or U6131 (N_6131,N_5143,N_5964);
nand U6132 (N_6132,N_5271,N_5519);
nand U6133 (N_6133,N_5662,N_5797);
nor U6134 (N_6134,N_5878,N_5790);
or U6135 (N_6135,N_5025,N_5693);
nand U6136 (N_6136,N_5313,N_5708);
or U6137 (N_6137,N_5852,N_5560);
and U6138 (N_6138,N_5445,N_5933);
or U6139 (N_6139,N_5061,N_5530);
or U6140 (N_6140,N_5325,N_5969);
or U6141 (N_6141,N_5736,N_5114);
or U6142 (N_6142,N_5762,N_5944);
and U6143 (N_6143,N_5174,N_5823);
nor U6144 (N_6144,N_5228,N_5135);
nor U6145 (N_6145,N_5989,N_5591);
nor U6146 (N_6146,N_5613,N_5024);
nor U6147 (N_6147,N_5704,N_5622);
and U6148 (N_6148,N_5351,N_5563);
or U6149 (N_6149,N_5967,N_5293);
nand U6150 (N_6150,N_5050,N_5086);
xor U6151 (N_6151,N_5270,N_5406);
and U6152 (N_6152,N_5358,N_5175);
xnor U6153 (N_6153,N_5932,N_5292);
nand U6154 (N_6154,N_5986,N_5155);
nand U6155 (N_6155,N_5324,N_5225);
and U6156 (N_6156,N_5391,N_5821);
or U6157 (N_6157,N_5614,N_5066);
nor U6158 (N_6158,N_5387,N_5830);
nor U6159 (N_6159,N_5865,N_5609);
or U6160 (N_6160,N_5291,N_5179);
nor U6161 (N_6161,N_5740,N_5242);
nand U6162 (N_6162,N_5440,N_5520);
nor U6163 (N_6163,N_5111,N_5755);
or U6164 (N_6164,N_5421,N_5911);
nor U6165 (N_6165,N_5209,N_5866);
nor U6166 (N_6166,N_5898,N_5805);
or U6167 (N_6167,N_5877,N_5631);
nor U6168 (N_6168,N_5198,N_5843);
and U6169 (N_6169,N_5359,N_5410);
nand U6170 (N_6170,N_5922,N_5454);
or U6171 (N_6171,N_5294,N_5180);
nand U6172 (N_6172,N_5208,N_5261);
nor U6173 (N_6173,N_5600,N_5941);
and U6174 (N_6174,N_5424,N_5925);
nor U6175 (N_6175,N_5394,N_5806);
xnor U6176 (N_6176,N_5525,N_5482);
and U6177 (N_6177,N_5057,N_5221);
nand U6178 (N_6178,N_5547,N_5163);
or U6179 (N_6179,N_5263,N_5137);
nor U6180 (N_6180,N_5770,N_5017);
nor U6181 (N_6181,N_5758,N_5460);
and U6182 (N_6182,N_5205,N_5856);
or U6183 (N_6183,N_5196,N_5962);
or U6184 (N_6184,N_5589,N_5214);
or U6185 (N_6185,N_5162,N_5548);
nand U6186 (N_6186,N_5784,N_5699);
nor U6187 (N_6187,N_5182,N_5368);
or U6188 (N_6188,N_5757,N_5820);
nor U6189 (N_6189,N_5195,N_5075);
or U6190 (N_6190,N_5996,N_5713);
and U6191 (N_6191,N_5328,N_5789);
nand U6192 (N_6192,N_5626,N_5090);
nor U6193 (N_6193,N_5367,N_5003);
and U6194 (N_6194,N_5608,N_5504);
nand U6195 (N_6195,N_5824,N_5415);
xor U6196 (N_6196,N_5771,N_5452);
xor U6197 (N_6197,N_5335,N_5640);
nor U6198 (N_6198,N_5660,N_5938);
nor U6199 (N_6199,N_5134,N_5506);
or U6200 (N_6200,N_5857,N_5297);
nand U6201 (N_6201,N_5761,N_5582);
or U6202 (N_6202,N_5826,N_5691);
or U6203 (N_6203,N_5389,N_5378);
and U6204 (N_6204,N_5039,N_5798);
nor U6205 (N_6205,N_5124,N_5927);
and U6206 (N_6206,N_5349,N_5948);
nor U6207 (N_6207,N_5628,N_5112);
xor U6208 (N_6208,N_5069,N_5882);
and U6209 (N_6209,N_5011,N_5098);
and U6210 (N_6210,N_5138,N_5675);
nor U6211 (N_6211,N_5471,N_5012);
or U6212 (N_6212,N_5639,N_5741);
nand U6213 (N_6213,N_5379,N_5649);
and U6214 (N_6214,N_5053,N_5067);
nand U6215 (N_6215,N_5285,N_5946);
and U6216 (N_6216,N_5565,N_5016);
or U6217 (N_6217,N_5441,N_5259);
and U6218 (N_6218,N_5347,N_5126);
and U6219 (N_6219,N_5643,N_5931);
or U6220 (N_6220,N_5910,N_5241);
xor U6221 (N_6221,N_5903,N_5666);
nor U6222 (N_6222,N_5077,N_5524);
or U6223 (N_6223,N_5152,N_5197);
nor U6224 (N_6224,N_5383,N_5908);
or U6225 (N_6225,N_5031,N_5376);
or U6226 (N_6226,N_5863,N_5701);
or U6227 (N_6227,N_5987,N_5867);
xor U6228 (N_6228,N_5584,N_5334);
or U6229 (N_6229,N_5048,N_5795);
and U6230 (N_6230,N_5142,N_5033);
nor U6231 (N_6231,N_5382,N_5348);
and U6232 (N_6232,N_5226,N_5884);
nor U6233 (N_6233,N_5262,N_5538);
nor U6234 (N_6234,N_5448,N_5296);
and U6235 (N_6235,N_5133,N_5773);
or U6236 (N_6236,N_5853,N_5507);
and U6237 (N_6237,N_5220,N_5869);
or U6238 (N_6238,N_5309,N_5750);
xor U6239 (N_6239,N_5341,N_5935);
nor U6240 (N_6240,N_5575,N_5118);
nand U6241 (N_6241,N_5559,N_5572);
and U6242 (N_6242,N_5629,N_5194);
nand U6243 (N_6243,N_5561,N_5267);
or U6244 (N_6244,N_5366,N_5153);
nor U6245 (N_6245,N_5861,N_5419);
nand U6246 (N_6246,N_5664,N_5353);
xor U6247 (N_6247,N_5796,N_5667);
and U6248 (N_6248,N_5212,N_5847);
and U6249 (N_6249,N_5647,N_5373);
nand U6250 (N_6250,N_5123,N_5321);
nor U6251 (N_6251,N_5312,N_5446);
nor U6252 (N_6252,N_5891,N_5034);
nand U6253 (N_6253,N_5233,N_5975);
or U6254 (N_6254,N_5167,N_5607);
or U6255 (N_6255,N_5408,N_5425);
nand U6256 (N_6256,N_5088,N_5669);
or U6257 (N_6257,N_5390,N_5543);
nand U6258 (N_6258,N_5362,N_5166);
or U6259 (N_6259,N_5573,N_5981);
nand U6260 (N_6260,N_5015,N_5571);
and U6261 (N_6261,N_5794,N_5339);
or U6262 (N_6262,N_5912,N_5879);
or U6263 (N_6263,N_5165,N_5306);
nand U6264 (N_6264,N_5909,N_5416);
or U6265 (N_6265,N_5528,N_5642);
or U6266 (N_6266,N_5841,N_5984);
nor U6267 (N_6267,N_5467,N_5972);
nand U6268 (N_6268,N_5505,N_5396);
nor U6269 (N_6269,N_5803,N_5715);
xor U6270 (N_6270,N_5223,N_5775);
and U6271 (N_6271,N_5356,N_5283);
and U6272 (N_6272,N_5929,N_5304);
and U6273 (N_6273,N_5827,N_5030);
nand U6274 (N_6274,N_5449,N_5310);
and U6275 (N_6275,N_5392,N_5256);
nor U6276 (N_6276,N_5875,N_5301);
or U6277 (N_6277,N_5160,N_5663);
or U6278 (N_6278,N_5682,N_5318);
xor U6279 (N_6279,N_5481,N_5044);
xor U6280 (N_6280,N_5567,N_5215);
and U6281 (N_6281,N_5239,N_5966);
nor U6282 (N_6282,N_5526,N_5968);
nand U6283 (N_6283,N_5110,N_5730);
or U6284 (N_6284,N_5000,N_5176);
nor U6285 (N_6285,N_5657,N_5939);
nand U6286 (N_6286,N_5107,N_5058);
and U6287 (N_6287,N_5201,N_5487);
and U6288 (N_6288,N_5951,N_5783);
nor U6289 (N_6289,N_5793,N_5009);
xnor U6290 (N_6290,N_5509,N_5257);
nor U6291 (N_6291,N_5172,N_5423);
xor U6292 (N_6292,N_5737,N_5275);
and U6293 (N_6293,N_5742,N_5464);
and U6294 (N_6294,N_5409,N_5870);
or U6295 (N_6295,N_5217,N_5246);
or U6296 (N_6296,N_5330,N_5237);
nor U6297 (N_6297,N_5229,N_5849);
and U6298 (N_6298,N_5928,N_5398);
nand U6299 (N_6299,N_5595,N_5659);
and U6300 (N_6300,N_5658,N_5914);
nand U6301 (N_6301,N_5913,N_5864);
and U6302 (N_6302,N_5036,N_5749);
nor U6303 (N_6303,N_5120,N_5684);
or U6304 (N_6304,N_5638,N_5248);
nand U6305 (N_6305,N_5814,N_5876);
nand U6306 (N_6306,N_5558,N_5289);
xor U6307 (N_6307,N_5043,N_5185);
nor U6308 (N_6308,N_5598,N_5859);
and U6309 (N_6309,N_5013,N_5883);
nand U6310 (N_6310,N_5791,N_5403);
nor U6311 (N_6311,N_5683,N_5211);
and U6312 (N_6312,N_5052,N_5085);
or U6313 (N_6313,N_5544,N_5900);
xnor U6314 (N_6314,N_5748,N_5971);
nand U6315 (N_6315,N_5430,N_5676);
nor U6316 (N_6316,N_5380,N_5218);
nand U6317 (N_6317,N_5045,N_5906);
nor U6318 (N_6318,N_5485,N_5768);
nor U6319 (N_6319,N_5934,N_5844);
xnor U6320 (N_6320,N_5177,N_5355);
xor U6321 (N_6321,N_5342,N_5193);
xnor U6322 (N_6322,N_5838,N_5314);
or U6323 (N_6323,N_5641,N_5517);
and U6324 (N_6324,N_5041,N_5159);
nor U6325 (N_6325,N_5616,N_5183);
or U6326 (N_6326,N_5101,N_5422);
xor U6327 (N_6327,N_5244,N_5371);
xor U6328 (N_6328,N_5670,N_5463);
and U6329 (N_6329,N_5329,N_5672);
and U6330 (N_6330,N_5412,N_5224);
nor U6331 (N_6331,N_5149,N_5860);
nor U6332 (N_6332,N_5918,N_5357);
and U6333 (N_6333,N_5535,N_5534);
nor U6334 (N_6334,N_5549,N_5104);
xor U6335 (N_6335,N_5782,N_5735);
and U6336 (N_6336,N_5990,N_5722);
or U6337 (N_6337,N_5480,N_5188);
nand U6338 (N_6338,N_5386,N_5627);
or U6339 (N_6339,N_5848,N_5465);
nor U6340 (N_6340,N_5395,N_5498);
xnor U6341 (N_6341,N_5760,N_5037);
nor U6342 (N_6342,N_5697,N_5581);
or U6343 (N_6343,N_5222,N_5592);
and U6344 (N_6344,N_5488,N_5635);
nand U6345 (N_6345,N_5455,N_5393);
nand U6346 (N_6346,N_5173,N_5260);
nand U6347 (N_6347,N_5837,N_5508);
and U6348 (N_6348,N_5266,N_5150);
nand U6349 (N_6349,N_5835,N_5788);
nor U6350 (N_6350,N_5597,N_5468);
nand U6351 (N_6351,N_5265,N_5020);
or U6352 (N_6352,N_5068,N_5113);
xor U6353 (N_6353,N_5007,N_5720);
xor U6354 (N_6354,N_5897,N_5702);
or U6355 (N_6355,N_5129,N_5550);
nand U6356 (N_6356,N_5512,N_5916);
or U6357 (N_6357,N_5810,N_5436);
and U6358 (N_6358,N_5992,N_5746);
or U6359 (N_6359,N_5437,N_5461);
nor U6360 (N_6360,N_5326,N_5363);
or U6361 (N_6361,N_5955,N_5494);
nand U6362 (N_6362,N_5404,N_5456);
or U6363 (N_6363,N_5516,N_5536);
and U6364 (N_6364,N_5021,N_5420);
or U6365 (N_6365,N_5122,N_5930);
nor U6366 (N_6366,N_5842,N_5942);
nand U6367 (N_6367,N_5079,N_5650);
xnor U6368 (N_6368,N_5486,N_5109);
or U6369 (N_6369,N_5093,N_5718);
nand U6370 (N_6370,N_5950,N_5621);
and U6371 (N_6371,N_5014,N_5317);
xor U6372 (N_6372,N_5026,N_5307);
and U6373 (N_6373,N_5472,N_5617);
or U6374 (N_6374,N_5308,N_5555);
and U6375 (N_6375,N_5546,N_5288);
or U6376 (N_6376,N_5399,N_5302);
nor U6377 (N_6377,N_5336,N_5213);
nand U6378 (N_6378,N_5029,N_5046);
xnor U6379 (N_6379,N_5084,N_5729);
and U6380 (N_6380,N_5035,N_5759);
nor U6381 (N_6381,N_5092,N_5833);
and U6382 (N_6382,N_5431,N_5103);
and U6383 (N_6383,N_5880,N_5818);
and U6384 (N_6384,N_5834,N_5907);
nor U6385 (N_6385,N_5601,N_5845);
nor U6386 (N_6386,N_5106,N_5411);
or U6387 (N_6387,N_5040,N_5168);
or U6388 (N_6388,N_5190,N_5116);
and U6389 (N_6389,N_5892,N_5280);
and U6390 (N_6390,N_5001,N_5765);
and U6391 (N_6391,N_5825,N_5273);
nand U6392 (N_6392,N_5095,N_5809);
nor U6393 (N_6393,N_5562,N_5991);
or U6394 (N_6394,N_5698,N_5154);
nand U6395 (N_6395,N_5300,N_5924);
nand U6396 (N_6396,N_5377,N_5518);
xor U6397 (N_6397,N_5953,N_5739);
nor U6398 (N_6398,N_5287,N_5665);
or U6399 (N_6399,N_5625,N_5624);
nand U6400 (N_6400,N_5542,N_5888);
and U6401 (N_6401,N_5005,N_5886);
and U6402 (N_6402,N_5588,N_5901);
xnor U6403 (N_6403,N_5243,N_5656);
nor U6404 (N_6404,N_5091,N_5619);
xnor U6405 (N_6405,N_5636,N_5537);
and U6406 (N_6406,N_5717,N_5099);
nor U6407 (N_6407,N_5234,N_5681);
nand U6408 (N_6408,N_5620,N_5457);
and U6409 (N_6409,N_5171,N_5051);
or U6410 (N_6410,N_5476,N_5532);
nand U6411 (N_6411,N_5290,N_5719);
and U6412 (N_6412,N_5724,N_5479);
or U6413 (N_6413,N_5115,N_5603);
xor U6414 (N_6414,N_5899,N_5686);
and U6415 (N_6415,N_5254,N_5733);
or U6416 (N_6416,N_5125,N_5764);
nor U6417 (N_6417,N_5721,N_5862);
and U6418 (N_6418,N_5633,N_5354);
or U6419 (N_6419,N_5832,N_5576);
nand U6420 (N_6420,N_5370,N_5958);
and U6421 (N_6421,N_5074,N_5753);
or U6422 (N_6422,N_5286,N_5671);
or U6423 (N_6423,N_5569,N_5688);
and U6424 (N_6424,N_5685,N_5872);
and U6425 (N_6425,N_5711,N_5965);
or U6426 (N_6426,N_5435,N_5527);
xnor U6427 (N_6427,N_5811,N_5556);
and U6428 (N_6428,N_5322,N_5728);
and U6429 (N_6429,N_5466,N_5151);
xor U6430 (N_6430,N_5130,N_5072);
and U6431 (N_6431,N_5269,N_5587);
nor U6432 (N_6432,N_5902,N_5361);
or U6433 (N_6433,N_5402,N_5668);
and U6434 (N_6434,N_5298,N_5474);
nor U6435 (N_6435,N_5514,N_5993);
nand U6436 (N_6436,N_5593,N_5846);
or U6437 (N_6437,N_5513,N_5008);
xor U6438 (N_6438,N_5004,N_5338);
nor U6439 (N_6439,N_5956,N_5709);
or U6440 (N_6440,N_5407,N_5427);
or U6441 (N_6441,N_5235,N_5734);
and U6442 (N_6442,N_5503,N_5580);
or U6443 (N_6443,N_5952,N_5027);
nor U6444 (N_6444,N_5238,N_5469);
xor U6445 (N_6445,N_5490,N_5073);
nor U6446 (N_6446,N_5018,N_5002);
or U6447 (N_6447,N_5726,N_5146);
nand U6448 (N_6448,N_5200,N_5926);
and U6449 (N_6449,N_5417,N_5738);
or U6450 (N_6450,N_5459,N_5501);
and U6451 (N_6451,N_5585,N_5489);
or U6452 (N_6452,N_5245,N_5255);
or U6453 (N_6453,N_5054,N_5189);
xor U6454 (N_6454,N_5959,N_5413);
xnor U6455 (N_6455,N_5484,N_5874);
nand U6456 (N_6456,N_5529,N_5905);
or U6457 (N_6457,N_5327,N_5960);
or U6458 (N_6458,N_5868,N_5316);
nand U6459 (N_6459,N_5937,N_5732);
xnor U6460 (N_6460,N_5936,N_5787);
or U6461 (N_6461,N_5700,N_5896);
nand U6462 (N_6462,N_5191,N_5979);
or U6463 (N_6463,N_5819,N_5108);
nor U6464 (N_6464,N_5055,N_5232);
or U6465 (N_6465,N_5450,N_5117);
nor U6466 (N_6466,N_5915,N_5140);
xor U6467 (N_6467,N_5851,N_5272);
nand U6468 (N_6468,N_5128,N_5161);
nand U6469 (N_6469,N_5493,N_5893);
nor U6470 (N_6470,N_5610,N_5648);
nand U6471 (N_6471,N_5545,N_5303);
and U6472 (N_6472,N_5822,N_5523);
xor U6473 (N_6473,N_5887,N_5655);
nand U6474 (N_6474,N_5604,N_5192);
and U6475 (N_6475,N_5089,N_5429);
or U6476 (N_6476,N_5976,N_5375);
and U6477 (N_6477,N_5144,N_5491);
or U6478 (N_6478,N_5081,N_5147);
xor U6479 (N_6479,N_5540,N_5885);
nor U6480 (N_6480,N_5568,N_5815);
or U6481 (N_6481,N_5299,N_5743);
or U6482 (N_6482,N_5705,N_5687);
or U6483 (N_6483,N_5583,N_5703);
nor U6484 (N_6484,N_5774,N_5352);
and U6485 (N_6485,N_5515,N_5801);
and U6486 (N_6486,N_5210,N_5679);
xnor U6487 (N_6487,N_5320,N_5808);
nand U6488 (N_6488,N_5828,N_5049);
nand U6489 (N_6489,N_5023,N_5695);
and U6490 (N_6490,N_5364,N_5276);
or U6491 (N_6491,N_5219,N_5019);
or U6492 (N_6492,N_5028,N_5623);
or U6493 (N_6493,N_5813,N_5653);
and U6494 (N_6494,N_5766,N_5871);
nand U6495 (N_6495,N_5651,N_5533);
nor U6496 (N_6496,N_5136,N_5319);
and U6497 (N_6497,N_5661,N_5786);
xor U6498 (N_6498,N_5119,N_5723);
or U6499 (N_6499,N_5426,N_5169);
nor U6500 (N_6500,N_5857,N_5134);
or U6501 (N_6501,N_5653,N_5498);
nor U6502 (N_6502,N_5929,N_5611);
or U6503 (N_6503,N_5246,N_5654);
nand U6504 (N_6504,N_5239,N_5681);
nor U6505 (N_6505,N_5709,N_5946);
xor U6506 (N_6506,N_5683,N_5620);
nand U6507 (N_6507,N_5533,N_5657);
nand U6508 (N_6508,N_5863,N_5919);
and U6509 (N_6509,N_5618,N_5866);
nor U6510 (N_6510,N_5650,N_5706);
nand U6511 (N_6511,N_5334,N_5007);
or U6512 (N_6512,N_5235,N_5871);
nor U6513 (N_6513,N_5111,N_5062);
nand U6514 (N_6514,N_5903,N_5326);
and U6515 (N_6515,N_5637,N_5538);
nand U6516 (N_6516,N_5664,N_5215);
xnor U6517 (N_6517,N_5859,N_5733);
xnor U6518 (N_6518,N_5817,N_5167);
nor U6519 (N_6519,N_5189,N_5292);
or U6520 (N_6520,N_5374,N_5127);
nor U6521 (N_6521,N_5569,N_5670);
nand U6522 (N_6522,N_5467,N_5050);
nand U6523 (N_6523,N_5728,N_5480);
nand U6524 (N_6524,N_5605,N_5960);
and U6525 (N_6525,N_5168,N_5519);
xnor U6526 (N_6526,N_5891,N_5078);
or U6527 (N_6527,N_5540,N_5351);
nand U6528 (N_6528,N_5120,N_5839);
nand U6529 (N_6529,N_5748,N_5683);
and U6530 (N_6530,N_5455,N_5127);
or U6531 (N_6531,N_5173,N_5836);
nand U6532 (N_6532,N_5478,N_5426);
nor U6533 (N_6533,N_5699,N_5377);
nor U6534 (N_6534,N_5707,N_5052);
xor U6535 (N_6535,N_5701,N_5905);
nand U6536 (N_6536,N_5059,N_5449);
nor U6537 (N_6537,N_5573,N_5887);
and U6538 (N_6538,N_5529,N_5527);
nor U6539 (N_6539,N_5700,N_5377);
and U6540 (N_6540,N_5925,N_5045);
nor U6541 (N_6541,N_5606,N_5006);
nor U6542 (N_6542,N_5493,N_5865);
nor U6543 (N_6543,N_5725,N_5495);
nor U6544 (N_6544,N_5969,N_5330);
nor U6545 (N_6545,N_5202,N_5816);
or U6546 (N_6546,N_5949,N_5081);
xor U6547 (N_6547,N_5446,N_5093);
nor U6548 (N_6548,N_5627,N_5008);
nand U6549 (N_6549,N_5610,N_5783);
nand U6550 (N_6550,N_5676,N_5366);
nor U6551 (N_6551,N_5779,N_5288);
nand U6552 (N_6552,N_5839,N_5228);
nand U6553 (N_6553,N_5873,N_5228);
nor U6554 (N_6554,N_5839,N_5394);
nand U6555 (N_6555,N_5258,N_5482);
nand U6556 (N_6556,N_5837,N_5400);
nand U6557 (N_6557,N_5477,N_5498);
and U6558 (N_6558,N_5551,N_5572);
nor U6559 (N_6559,N_5787,N_5756);
or U6560 (N_6560,N_5270,N_5238);
nor U6561 (N_6561,N_5873,N_5794);
and U6562 (N_6562,N_5967,N_5020);
and U6563 (N_6563,N_5001,N_5150);
and U6564 (N_6564,N_5600,N_5443);
nor U6565 (N_6565,N_5066,N_5988);
and U6566 (N_6566,N_5980,N_5376);
nor U6567 (N_6567,N_5583,N_5887);
nor U6568 (N_6568,N_5608,N_5034);
xor U6569 (N_6569,N_5743,N_5566);
nand U6570 (N_6570,N_5751,N_5810);
nand U6571 (N_6571,N_5102,N_5094);
nor U6572 (N_6572,N_5923,N_5633);
xnor U6573 (N_6573,N_5518,N_5619);
nor U6574 (N_6574,N_5684,N_5069);
nor U6575 (N_6575,N_5292,N_5019);
and U6576 (N_6576,N_5284,N_5063);
nor U6577 (N_6577,N_5488,N_5026);
nor U6578 (N_6578,N_5498,N_5200);
nand U6579 (N_6579,N_5179,N_5422);
nor U6580 (N_6580,N_5182,N_5924);
nand U6581 (N_6581,N_5432,N_5203);
nand U6582 (N_6582,N_5503,N_5359);
and U6583 (N_6583,N_5326,N_5770);
and U6584 (N_6584,N_5895,N_5495);
and U6585 (N_6585,N_5145,N_5159);
nand U6586 (N_6586,N_5034,N_5423);
or U6587 (N_6587,N_5514,N_5647);
and U6588 (N_6588,N_5250,N_5762);
or U6589 (N_6589,N_5108,N_5248);
and U6590 (N_6590,N_5699,N_5573);
or U6591 (N_6591,N_5876,N_5658);
and U6592 (N_6592,N_5829,N_5231);
nand U6593 (N_6593,N_5547,N_5855);
nand U6594 (N_6594,N_5044,N_5666);
xor U6595 (N_6595,N_5599,N_5595);
xnor U6596 (N_6596,N_5201,N_5421);
or U6597 (N_6597,N_5808,N_5722);
nor U6598 (N_6598,N_5405,N_5737);
nor U6599 (N_6599,N_5636,N_5343);
and U6600 (N_6600,N_5391,N_5802);
nor U6601 (N_6601,N_5782,N_5338);
or U6602 (N_6602,N_5051,N_5559);
and U6603 (N_6603,N_5221,N_5547);
or U6604 (N_6604,N_5007,N_5928);
nand U6605 (N_6605,N_5879,N_5860);
and U6606 (N_6606,N_5806,N_5752);
xnor U6607 (N_6607,N_5614,N_5212);
or U6608 (N_6608,N_5315,N_5784);
and U6609 (N_6609,N_5565,N_5647);
and U6610 (N_6610,N_5638,N_5300);
and U6611 (N_6611,N_5943,N_5293);
nor U6612 (N_6612,N_5834,N_5748);
or U6613 (N_6613,N_5230,N_5781);
xnor U6614 (N_6614,N_5143,N_5711);
or U6615 (N_6615,N_5482,N_5876);
nor U6616 (N_6616,N_5950,N_5317);
or U6617 (N_6617,N_5979,N_5088);
xnor U6618 (N_6618,N_5941,N_5516);
nand U6619 (N_6619,N_5521,N_5136);
or U6620 (N_6620,N_5050,N_5280);
nand U6621 (N_6621,N_5680,N_5473);
or U6622 (N_6622,N_5461,N_5088);
nand U6623 (N_6623,N_5211,N_5580);
and U6624 (N_6624,N_5321,N_5429);
and U6625 (N_6625,N_5489,N_5153);
or U6626 (N_6626,N_5878,N_5615);
or U6627 (N_6627,N_5161,N_5600);
and U6628 (N_6628,N_5170,N_5964);
nor U6629 (N_6629,N_5067,N_5481);
xnor U6630 (N_6630,N_5925,N_5100);
nand U6631 (N_6631,N_5277,N_5917);
or U6632 (N_6632,N_5390,N_5053);
nor U6633 (N_6633,N_5874,N_5430);
and U6634 (N_6634,N_5930,N_5995);
or U6635 (N_6635,N_5727,N_5225);
nand U6636 (N_6636,N_5455,N_5836);
or U6637 (N_6637,N_5574,N_5956);
or U6638 (N_6638,N_5120,N_5308);
or U6639 (N_6639,N_5746,N_5075);
nor U6640 (N_6640,N_5173,N_5383);
and U6641 (N_6641,N_5304,N_5540);
nor U6642 (N_6642,N_5821,N_5635);
and U6643 (N_6643,N_5194,N_5451);
xor U6644 (N_6644,N_5610,N_5890);
nor U6645 (N_6645,N_5156,N_5901);
nand U6646 (N_6646,N_5440,N_5782);
nor U6647 (N_6647,N_5478,N_5043);
and U6648 (N_6648,N_5247,N_5912);
or U6649 (N_6649,N_5836,N_5258);
nand U6650 (N_6650,N_5667,N_5611);
and U6651 (N_6651,N_5491,N_5504);
nor U6652 (N_6652,N_5175,N_5330);
nor U6653 (N_6653,N_5421,N_5364);
nor U6654 (N_6654,N_5554,N_5494);
nand U6655 (N_6655,N_5210,N_5704);
or U6656 (N_6656,N_5578,N_5358);
or U6657 (N_6657,N_5815,N_5875);
or U6658 (N_6658,N_5468,N_5092);
and U6659 (N_6659,N_5239,N_5180);
nor U6660 (N_6660,N_5355,N_5011);
xor U6661 (N_6661,N_5065,N_5730);
or U6662 (N_6662,N_5941,N_5233);
nand U6663 (N_6663,N_5428,N_5947);
nand U6664 (N_6664,N_5755,N_5201);
and U6665 (N_6665,N_5737,N_5359);
or U6666 (N_6666,N_5873,N_5994);
nor U6667 (N_6667,N_5415,N_5267);
and U6668 (N_6668,N_5853,N_5031);
nand U6669 (N_6669,N_5401,N_5882);
nand U6670 (N_6670,N_5309,N_5663);
nand U6671 (N_6671,N_5446,N_5017);
nor U6672 (N_6672,N_5651,N_5092);
or U6673 (N_6673,N_5909,N_5226);
and U6674 (N_6674,N_5460,N_5934);
nand U6675 (N_6675,N_5847,N_5802);
nand U6676 (N_6676,N_5563,N_5400);
and U6677 (N_6677,N_5006,N_5150);
nand U6678 (N_6678,N_5337,N_5349);
and U6679 (N_6679,N_5939,N_5589);
nor U6680 (N_6680,N_5619,N_5921);
nor U6681 (N_6681,N_5637,N_5287);
nand U6682 (N_6682,N_5294,N_5298);
and U6683 (N_6683,N_5630,N_5141);
and U6684 (N_6684,N_5644,N_5184);
and U6685 (N_6685,N_5122,N_5787);
and U6686 (N_6686,N_5264,N_5243);
or U6687 (N_6687,N_5714,N_5765);
and U6688 (N_6688,N_5208,N_5985);
nand U6689 (N_6689,N_5388,N_5812);
and U6690 (N_6690,N_5278,N_5401);
or U6691 (N_6691,N_5383,N_5483);
and U6692 (N_6692,N_5511,N_5423);
xor U6693 (N_6693,N_5182,N_5303);
nor U6694 (N_6694,N_5148,N_5445);
nor U6695 (N_6695,N_5214,N_5045);
or U6696 (N_6696,N_5258,N_5465);
or U6697 (N_6697,N_5851,N_5227);
nand U6698 (N_6698,N_5834,N_5435);
nor U6699 (N_6699,N_5158,N_5426);
nor U6700 (N_6700,N_5790,N_5247);
and U6701 (N_6701,N_5182,N_5619);
xnor U6702 (N_6702,N_5566,N_5801);
and U6703 (N_6703,N_5529,N_5548);
and U6704 (N_6704,N_5440,N_5849);
or U6705 (N_6705,N_5896,N_5472);
or U6706 (N_6706,N_5614,N_5795);
nor U6707 (N_6707,N_5890,N_5115);
or U6708 (N_6708,N_5857,N_5577);
and U6709 (N_6709,N_5791,N_5621);
or U6710 (N_6710,N_5618,N_5754);
nor U6711 (N_6711,N_5699,N_5338);
and U6712 (N_6712,N_5013,N_5459);
xnor U6713 (N_6713,N_5551,N_5611);
or U6714 (N_6714,N_5369,N_5938);
or U6715 (N_6715,N_5297,N_5199);
nand U6716 (N_6716,N_5401,N_5605);
and U6717 (N_6717,N_5459,N_5089);
or U6718 (N_6718,N_5206,N_5604);
and U6719 (N_6719,N_5388,N_5165);
and U6720 (N_6720,N_5691,N_5149);
and U6721 (N_6721,N_5887,N_5380);
and U6722 (N_6722,N_5772,N_5136);
nand U6723 (N_6723,N_5022,N_5784);
and U6724 (N_6724,N_5262,N_5178);
or U6725 (N_6725,N_5389,N_5386);
or U6726 (N_6726,N_5321,N_5709);
xnor U6727 (N_6727,N_5990,N_5775);
and U6728 (N_6728,N_5566,N_5417);
and U6729 (N_6729,N_5153,N_5442);
and U6730 (N_6730,N_5209,N_5631);
or U6731 (N_6731,N_5256,N_5491);
nor U6732 (N_6732,N_5615,N_5205);
xor U6733 (N_6733,N_5285,N_5309);
nor U6734 (N_6734,N_5663,N_5992);
nor U6735 (N_6735,N_5342,N_5139);
nand U6736 (N_6736,N_5620,N_5837);
nand U6737 (N_6737,N_5694,N_5064);
xor U6738 (N_6738,N_5298,N_5918);
xor U6739 (N_6739,N_5470,N_5641);
nand U6740 (N_6740,N_5953,N_5241);
and U6741 (N_6741,N_5515,N_5462);
xor U6742 (N_6742,N_5911,N_5969);
nand U6743 (N_6743,N_5138,N_5921);
nor U6744 (N_6744,N_5857,N_5451);
xor U6745 (N_6745,N_5939,N_5218);
or U6746 (N_6746,N_5386,N_5228);
and U6747 (N_6747,N_5558,N_5822);
nand U6748 (N_6748,N_5249,N_5978);
or U6749 (N_6749,N_5139,N_5655);
nand U6750 (N_6750,N_5004,N_5043);
nand U6751 (N_6751,N_5156,N_5289);
nor U6752 (N_6752,N_5970,N_5782);
and U6753 (N_6753,N_5819,N_5039);
nand U6754 (N_6754,N_5034,N_5432);
and U6755 (N_6755,N_5414,N_5804);
nor U6756 (N_6756,N_5753,N_5427);
or U6757 (N_6757,N_5388,N_5615);
and U6758 (N_6758,N_5444,N_5926);
nor U6759 (N_6759,N_5640,N_5837);
nand U6760 (N_6760,N_5138,N_5142);
and U6761 (N_6761,N_5482,N_5241);
nand U6762 (N_6762,N_5404,N_5953);
nor U6763 (N_6763,N_5603,N_5681);
or U6764 (N_6764,N_5694,N_5654);
xor U6765 (N_6765,N_5735,N_5390);
nor U6766 (N_6766,N_5635,N_5631);
nand U6767 (N_6767,N_5338,N_5690);
xnor U6768 (N_6768,N_5575,N_5578);
xnor U6769 (N_6769,N_5037,N_5407);
or U6770 (N_6770,N_5875,N_5656);
nor U6771 (N_6771,N_5955,N_5207);
nand U6772 (N_6772,N_5205,N_5425);
nor U6773 (N_6773,N_5314,N_5531);
and U6774 (N_6774,N_5511,N_5616);
nor U6775 (N_6775,N_5950,N_5411);
nand U6776 (N_6776,N_5855,N_5398);
and U6777 (N_6777,N_5447,N_5496);
nor U6778 (N_6778,N_5918,N_5340);
xnor U6779 (N_6779,N_5813,N_5560);
or U6780 (N_6780,N_5940,N_5134);
nand U6781 (N_6781,N_5556,N_5445);
and U6782 (N_6782,N_5620,N_5192);
nor U6783 (N_6783,N_5886,N_5936);
nor U6784 (N_6784,N_5838,N_5952);
or U6785 (N_6785,N_5611,N_5775);
nand U6786 (N_6786,N_5967,N_5240);
xnor U6787 (N_6787,N_5172,N_5048);
and U6788 (N_6788,N_5696,N_5128);
nand U6789 (N_6789,N_5750,N_5086);
nand U6790 (N_6790,N_5819,N_5851);
nand U6791 (N_6791,N_5498,N_5997);
or U6792 (N_6792,N_5900,N_5848);
and U6793 (N_6793,N_5197,N_5884);
and U6794 (N_6794,N_5282,N_5536);
and U6795 (N_6795,N_5648,N_5211);
or U6796 (N_6796,N_5800,N_5279);
or U6797 (N_6797,N_5755,N_5122);
nand U6798 (N_6798,N_5828,N_5041);
xor U6799 (N_6799,N_5423,N_5887);
xnor U6800 (N_6800,N_5620,N_5833);
or U6801 (N_6801,N_5798,N_5703);
nand U6802 (N_6802,N_5974,N_5023);
xor U6803 (N_6803,N_5694,N_5195);
nor U6804 (N_6804,N_5464,N_5342);
or U6805 (N_6805,N_5707,N_5881);
nor U6806 (N_6806,N_5614,N_5016);
nor U6807 (N_6807,N_5070,N_5455);
and U6808 (N_6808,N_5871,N_5812);
nand U6809 (N_6809,N_5766,N_5449);
nand U6810 (N_6810,N_5457,N_5743);
nor U6811 (N_6811,N_5916,N_5272);
and U6812 (N_6812,N_5783,N_5102);
or U6813 (N_6813,N_5456,N_5491);
nand U6814 (N_6814,N_5512,N_5231);
nand U6815 (N_6815,N_5129,N_5228);
or U6816 (N_6816,N_5436,N_5124);
xor U6817 (N_6817,N_5049,N_5560);
or U6818 (N_6818,N_5730,N_5157);
or U6819 (N_6819,N_5350,N_5534);
nand U6820 (N_6820,N_5148,N_5463);
nor U6821 (N_6821,N_5138,N_5109);
nand U6822 (N_6822,N_5027,N_5760);
and U6823 (N_6823,N_5360,N_5088);
and U6824 (N_6824,N_5155,N_5999);
and U6825 (N_6825,N_5211,N_5548);
nor U6826 (N_6826,N_5702,N_5368);
or U6827 (N_6827,N_5087,N_5770);
nand U6828 (N_6828,N_5053,N_5507);
nor U6829 (N_6829,N_5492,N_5480);
or U6830 (N_6830,N_5456,N_5361);
nand U6831 (N_6831,N_5858,N_5134);
or U6832 (N_6832,N_5424,N_5586);
nor U6833 (N_6833,N_5049,N_5120);
and U6834 (N_6834,N_5626,N_5997);
nand U6835 (N_6835,N_5970,N_5748);
or U6836 (N_6836,N_5293,N_5113);
or U6837 (N_6837,N_5454,N_5471);
and U6838 (N_6838,N_5439,N_5601);
nand U6839 (N_6839,N_5147,N_5428);
nor U6840 (N_6840,N_5649,N_5846);
nor U6841 (N_6841,N_5984,N_5152);
and U6842 (N_6842,N_5057,N_5905);
nor U6843 (N_6843,N_5462,N_5538);
nand U6844 (N_6844,N_5896,N_5096);
and U6845 (N_6845,N_5504,N_5758);
xnor U6846 (N_6846,N_5823,N_5474);
and U6847 (N_6847,N_5316,N_5746);
or U6848 (N_6848,N_5497,N_5294);
xor U6849 (N_6849,N_5619,N_5791);
or U6850 (N_6850,N_5934,N_5665);
nor U6851 (N_6851,N_5031,N_5927);
xor U6852 (N_6852,N_5967,N_5739);
nand U6853 (N_6853,N_5289,N_5929);
nor U6854 (N_6854,N_5630,N_5775);
and U6855 (N_6855,N_5248,N_5755);
nor U6856 (N_6856,N_5935,N_5182);
or U6857 (N_6857,N_5211,N_5760);
xnor U6858 (N_6858,N_5848,N_5261);
or U6859 (N_6859,N_5303,N_5152);
nand U6860 (N_6860,N_5165,N_5965);
xor U6861 (N_6861,N_5826,N_5322);
nand U6862 (N_6862,N_5808,N_5715);
nor U6863 (N_6863,N_5119,N_5549);
or U6864 (N_6864,N_5400,N_5621);
or U6865 (N_6865,N_5230,N_5880);
and U6866 (N_6866,N_5749,N_5111);
nand U6867 (N_6867,N_5866,N_5295);
nor U6868 (N_6868,N_5389,N_5437);
and U6869 (N_6869,N_5131,N_5065);
nand U6870 (N_6870,N_5077,N_5340);
nand U6871 (N_6871,N_5441,N_5603);
or U6872 (N_6872,N_5922,N_5443);
and U6873 (N_6873,N_5652,N_5774);
and U6874 (N_6874,N_5880,N_5912);
and U6875 (N_6875,N_5556,N_5741);
xnor U6876 (N_6876,N_5184,N_5495);
xnor U6877 (N_6877,N_5479,N_5940);
nand U6878 (N_6878,N_5323,N_5988);
nor U6879 (N_6879,N_5202,N_5757);
and U6880 (N_6880,N_5148,N_5558);
and U6881 (N_6881,N_5976,N_5296);
or U6882 (N_6882,N_5782,N_5688);
nand U6883 (N_6883,N_5102,N_5215);
nor U6884 (N_6884,N_5227,N_5915);
or U6885 (N_6885,N_5222,N_5362);
and U6886 (N_6886,N_5468,N_5447);
and U6887 (N_6887,N_5794,N_5842);
nor U6888 (N_6888,N_5015,N_5189);
and U6889 (N_6889,N_5768,N_5680);
and U6890 (N_6890,N_5220,N_5820);
nand U6891 (N_6891,N_5764,N_5013);
nand U6892 (N_6892,N_5622,N_5733);
and U6893 (N_6893,N_5369,N_5800);
or U6894 (N_6894,N_5640,N_5477);
and U6895 (N_6895,N_5886,N_5849);
and U6896 (N_6896,N_5869,N_5015);
nor U6897 (N_6897,N_5265,N_5961);
and U6898 (N_6898,N_5429,N_5555);
or U6899 (N_6899,N_5213,N_5248);
nand U6900 (N_6900,N_5671,N_5284);
or U6901 (N_6901,N_5748,N_5749);
and U6902 (N_6902,N_5650,N_5071);
nor U6903 (N_6903,N_5402,N_5389);
xor U6904 (N_6904,N_5696,N_5156);
nand U6905 (N_6905,N_5833,N_5081);
nor U6906 (N_6906,N_5933,N_5306);
or U6907 (N_6907,N_5045,N_5327);
nor U6908 (N_6908,N_5196,N_5380);
nand U6909 (N_6909,N_5356,N_5398);
nor U6910 (N_6910,N_5544,N_5483);
nand U6911 (N_6911,N_5235,N_5449);
nor U6912 (N_6912,N_5582,N_5443);
and U6913 (N_6913,N_5225,N_5845);
and U6914 (N_6914,N_5759,N_5895);
and U6915 (N_6915,N_5427,N_5342);
xnor U6916 (N_6916,N_5050,N_5588);
or U6917 (N_6917,N_5691,N_5576);
and U6918 (N_6918,N_5307,N_5122);
or U6919 (N_6919,N_5481,N_5212);
nor U6920 (N_6920,N_5665,N_5779);
or U6921 (N_6921,N_5599,N_5427);
or U6922 (N_6922,N_5851,N_5531);
nor U6923 (N_6923,N_5584,N_5770);
and U6924 (N_6924,N_5301,N_5649);
nand U6925 (N_6925,N_5232,N_5328);
nand U6926 (N_6926,N_5006,N_5332);
and U6927 (N_6927,N_5742,N_5596);
xnor U6928 (N_6928,N_5399,N_5795);
and U6929 (N_6929,N_5359,N_5084);
nand U6930 (N_6930,N_5797,N_5493);
or U6931 (N_6931,N_5347,N_5258);
nand U6932 (N_6932,N_5064,N_5944);
nand U6933 (N_6933,N_5895,N_5049);
nor U6934 (N_6934,N_5481,N_5013);
xor U6935 (N_6935,N_5814,N_5023);
nor U6936 (N_6936,N_5460,N_5657);
xnor U6937 (N_6937,N_5901,N_5513);
or U6938 (N_6938,N_5601,N_5382);
nand U6939 (N_6939,N_5814,N_5045);
nand U6940 (N_6940,N_5869,N_5534);
and U6941 (N_6941,N_5382,N_5352);
or U6942 (N_6942,N_5309,N_5740);
nand U6943 (N_6943,N_5202,N_5129);
or U6944 (N_6944,N_5103,N_5854);
xor U6945 (N_6945,N_5166,N_5701);
and U6946 (N_6946,N_5658,N_5041);
and U6947 (N_6947,N_5075,N_5135);
and U6948 (N_6948,N_5850,N_5416);
or U6949 (N_6949,N_5901,N_5747);
and U6950 (N_6950,N_5051,N_5386);
or U6951 (N_6951,N_5444,N_5333);
nand U6952 (N_6952,N_5305,N_5415);
nor U6953 (N_6953,N_5106,N_5776);
or U6954 (N_6954,N_5350,N_5805);
and U6955 (N_6955,N_5364,N_5580);
nand U6956 (N_6956,N_5458,N_5896);
or U6957 (N_6957,N_5847,N_5813);
or U6958 (N_6958,N_5407,N_5192);
and U6959 (N_6959,N_5711,N_5716);
nor U6960 (N_6960,N_5048,N_5385);
nand U6961 (N_6961,N_5225,N_5634);
xnor U6962 (N_6962,N_5619,N_5242);
nand U6963 (N_6963,N_5614,N_5498);
nand U6964 (N_6964,N_5520,N_5478);
nor U6965 (N_6965,N_5868,N_5360);
or U6966 (N_6966,N_5859,N_5148);
or U6967 (N_6967,N_5477,N_5079);
and U6968 (N_6968,N_5859,N_5510);
and U6969 (N_6969,N_5954,N_5750);
or U6970 (N_6970,N_5084,N_5808);
nor U6971 (N_6971,N_5380,N_5857);
or U6972 (N_6972,N_5243,N_5085);
nor U6973 (N_6973,N_5650,N_5623);
or U6974 (N_6974,N_5105,N_5242);
xnor U6975 (N_6975,N_5042,N_5602);
nor U6976 (N_6976,N_5169,N_5459);
xnor U6977 (N_6977,N_5600,N_5924);
nor U6978 (N_6978,N_5326,N_5215);
nand U6979 (N_6979,N_5532,N_5257);
or U6980 (N_6980,N_5965,N_5188);
or U6981 (N_6981,N_5720,N_5556);
or U6982 (N_6982,N_5658,N_5494);
and U6983 (N_6983,N_5507,N_5194);
nor U6984 (N_6984,N_5558,N_5201);
and U6985 (N_6985,N_5794,N_5868);
or U6986 (N_6986,N_5953,N_5415);
xnor U6987 (N_6987,N_5054,N_5297);
or U6988 (N_6988,N_5310,N_5888);
nand U6989 (N_6989,N_5710,N_5539);
and U6990 (N_6990,N_5384,N_5567);
nand U6991 (N_6991,N_5653,N_5328);
or U6992 (N_6992,N_5560,N_5987);
or U6993 (N_6993,N_5112,N_5800);
nor U6994 (N_6994,N_5297,N_5597);
and U6995 (N_6995,N_5274,N_5262);
or U6996 (N_6996,N_5949,N_5024);
and U6997 (N_6997,N_5636,N_5546);
nor U6998 (N_6998,N_5797,N_5137);
or U6999 (N_6999,N_5424,N_5154);
nor U7000 (N_7000,N_6118,N_6396);
nand U7001 (N_7001,N_6910,N_6376);
xor U7002 (N_7002,N_6007,N_6377);
and U7003 (N_7003,N_6086,N_6035);
xor U7004 (N_7004,N_6976,N_6730);
xnor U7005 (N_7005,N_6145,N_6224);
nor U7006 (N_7006,N_6471,N_6223);
nand U7007 (N_7007,N_6925,N_6555);
and U7008 (N_7008,N_6785,N_6257);
nand U7009 (N_7009,N_6983,N_6921);
xnor U7010 (N_7010,N_6809,N_6543);
or U7011 (N_7011,N_6315,N_6758);
nor U7012 (N_7012,N_6311,N_6703);
or U7013 (N_7013,N_6738,N_6905);
and U7014 (N_7014,N_6652,N_6161);
and U7015 (N_7015,N_6830,N_6904);
nand U7016 (N_7016,N_6680,N_6177);
or U7017 (N_7017,N_6822,N_6919);
and U7018 (N_7018,N_6528,N_6316);
nand U7019 (N_7019,N_6185,N_6868);
nand U7020 (N_7020,N_6916,N_6172);
or U7021 (N_7021,N_6599,N_6023);
and U7022 (N_7022,N_6737,N_6426);
nand U7023 (N_7023,N_6724,N_6792);
and U7024 (N_7024,N_6212,N_6256);
nor U7025 (N_7025,N_6998,N_6295);
nand U7026 (N_7026,N_6800,N_6337);
or U7027 (N_7027,N_6339,N_6138);
and U7028 (N_7028,N_6974,N_6382);
xnor U7029 (N_7029,N_6441,N_6187);
and U7030 (N_7030,N_6650,N_6777);
xnor U7031 (N_7031,N_6038,N_6569);
nand U7032 (N_7032,N_6099,N_6860);
and U7033 (N_7033,N_6550,N_6851);
nand U7034 (N_7034,N_6318,N_6207);
or U7035 (N_7035,N_6649,N_6701);
nand U7036 (N_7036,N_6957,N_6663);
nand U7037 (N_7037,N_6373,N_6620);
nor U7038 (N_7038,N_6358,N_6116);
xnor U7039 (N_7039,N_6900,N_6580);
nor U7040 (N_7040,N_6022,N_6829);
nor U7041 (N_7041,N_6855,N_6661);
nand U7042 (N_7042,N_6962,N_6516);
or U7043 (N_7043,N_6319,N_6763);
nor U7044 (N_7044,N_6492,N_6981);
and U7045 (N_7045,N_6158,N_6310);
or U7046 (N_7046,N_6191,N_6385);
or U7047 (N_7047,N_6840,N_6400);
or U7048 (N_7048,N_6206,N_6759);
nand U7049 (N_7049,N_6352,N_6253);
or U7050 (N_7050,N_6888,N_6596);
and U7051 (N_7051,N_6869,N_6784);
nor U7052 (N_7052,N_6130,N_6727);
or U7053 (N_7053,N_6065,N_6183);
nand U7054 (N_7054,N_6530,N_6806);
nand U7055 (N_7055,N_6936,N_6720);
nand U7056 (N_7056,N_6370,N_6912);
xor U7057 (N_7057,N_6141,N_6564);
or U7058 (N_7058,N_6458,N_6693);
nand U7059 (N_7059,N_6163,N_6837);
nor U7060 (N_7060,N_6406,N_6390);
nand U7061 (N_7061,N_6278,N_6131);
and U7062 (N_7062,N_6789,N_6895);
nor U7063 (N_7063,N_6250,N_6866);
nor U7064 (N_7064,N_6005,N_6695);
and U7065 (N_7065,N_6323,N_6155);
or U7066 (N_7066,N_6536,N_6330);
nand U7067 (N_7067,N_6051,N_6624);
xor U7068 (N_7068,N_6827,N_6526);
and U7069 (N_7069,N_6646,N_6261);
nand U7070 (N_7070,N_6314,N_6044);
or U7071 (N_7071,N_6908,N_6768);
xor U7072 (N_7072,N_6014,N_6032);
or U7073 (N_7073,N_6036,N_6419);
nand U7074 (N_7074,N_6560,N_6941);
nand U7075 (N_7075,N_6479,N_6101);
and U7076 (N_7076,N_6380,N_6274);
nor U7077 (N_7077,N_6689,N_6075);
or U7078 (N_7078,N_6710,N_6752);
or U7079 (N_7079,N_6520,N_6234);
and U7080 (N_7080,N_6462,N_6003);
nor U7081 (N_7081,N_6864,N_6457);
nor U7082 (N_7082,N_6772,N_6285);
or U7083 (N_7083,N_6579,N_6736);
nor U7084 (N_7084,N_6084,N_6168);
and U7085 (N_7085,N_6142,N_6948);
and U7086 (N_7086,N_6272,N_6364);
xor U7087 (N_7087,N_6808,N_6412);
xnor U7088 (N_7088,N_6688,N_6898);
nand U7089 (N_7089,N_6276,N_6843);
nand U7090 (N_7090,N_6016,N_6991);
nor U7091 (N_7091,N_6095,N_6133);
nor U7092 (N_7092,N_6934,N_6371);
or U7093 (N_7093,N_6993,N_6399);
nor U7094 (N_7094,N_6498,N_6748);
or U7095 (N_7095,N_6445,N_6271);
nor U7096 (N_7096,N_6870,N_6711);
nor U7097 (N_7097,N_6657,N_6388);
nand U7098 (N_7098,N_6113,N_6039);
nor U7099 (N_7099,N_6436,N_6556);
and U7100 (N_7100,N_6106,N_6205);
and U7101 (N_7101,N_6119,N_6514);
nand U7102 (N_7102,N_6653,N_6287);
nor U7103 (N_7103,N_6728,N_6629);
xor U7104 (N_7104,N_6774,N_6665);
and U7105 (N_7105,N_6346,N_6140);
nor U7106 (N_7106,N_6553,N_6424);
or U7107 (N_7107,N_6668,N_6963);
or U7108 (N_7108,N_6659,N_6715);
nand U7109 (N_7109,N_6117,N_6940);
nand U7110 (N_7110,N_6488,N_6590);
nor U7111 (N_7111,N_6468,N_6392);
nor U7112 (N_7112,N_6899,N_6719);
and U7113 (N_7113,N_6494,N_6486);
nor U7114 (N_7114,N_6745,N_6021);
and U7115 (N_7115,N_6561,N_6574);
or U7116 (N_7116,N_6078,N_6121);
and U7117 (N_7117,N_6831,N_6322);
nand U7118 (N_7118,N_6066,N_6911);
nand U7119 (N_7119,N_6173,N_6317);
or U7120 (N_7120,N_6398,N_6211);
nor U7121 (N_7121,N_6004,N_6418);
and U7122 (N_7122,N_6167,N_6055);
nand U7123 (N_7123,N_6175,N_6935);
xor U7124 (N_7124,N_6684,N_6291);
and U7125 (N_7125,N_6702,N_6679);
or U7126 (N_7126,N_6918,N_6028);
and U7127 (N_7127,N_6722,N_6781);
or U7128 (N_7128,N_6577,N_6930);
or U7129 (N_7129,N_6633,N_6862);
nor U7130 (N_7130,N_6273,N_6415);
and U7131 (N_7131,N_6944,N_6350);
xor U7132 (N_7132,N_6013,N_6334);
nand U7133 (N_7133,N_6447,N_6296);
or U7134 (N_7134,N_6074,N_6549);
nand U7135 (N_7135,N_6237,N_6456);
nand U7136 (N_7136,N_6959,N_6926);
or U7137 (N_7137,N_6776,N_6128);
or U7138 (N_7138,N_6241,N_6773);
nor U7139 (N_7139,N_6631,N_6662);
nand U7140 (N_7140,N_6188,N_6402);
and U7141 (N_7141,N_6416,N_6181);
nor U7142 (N_7142,N_6157,N_6923);
and U7143 (N_7143,N_6303,N_6239);
nand U7144 (N_7144,N_6306,N_6203);
nor U7145 (N_7145,N_6533,N_6793);
nand U7146 (N_7146,N_6089,N_6593);
nor U7147 (N_7147,N_6980,N_6780);
nor U7148 (N_7148,N_6651,N_6029);
nor U7149 (N_7149,N_6717,N_6884);
nor U7150 (N_7150,N_6664,N_6299);
nand U7151 (N_7151,N_6761,N_6443);
xor U7152 (N_7152,N_6425,N_6401);
or U7153 (N_7153,N_6849,N_6775);
nor U7154 (N_7154,N_6875,N_6685);
nor U7155 (N_7155,N_6159,N_6361);
or U7156 (N_7156,N_6542,N_6420);
nand U7157 (N_7157,N_6277,N_6369);
nand U7158 (N_7158,N_6790,N_6585);
nand U7159 (N_7159,N_6613,N_6137);
and U7160 (N_7160,N_6938,N_6641);
nand U7161 (N_7161,N_6833,N_6753);
or U7162 (N_7162,N_6491,N_6026);
xor U7163 (N_7163,N_6069,N_6521);
nor U7164 (N_7164,N_6623,N_6920);
xor U7165 (N_7165,N_6439,N_6076);
nor U7166 (N_7166,N_6913,N_6050);
nand U7167 (N_7167,N_6474,N_6942);
xor U7168 (N_7168,N_6674,N_6472);
nand U7169 (N_7169,N_6068,N_6325);
or U7170 (N_7170,N_6970,N_6270);
nor U7171 (N_7171,N_6791,N_6698);
or U7172 (N_7172,N_6015,N_6512);
nor U7173 (N_7173,N_6129,N_6867);
or U7174 (N_7174,N_6372,N_6890);
nand U7175 (N_7175,N_6081,N_6885);
or U7176 (N_7176,N_6294,N_6554);
or U7177 (N_7177,N_6927,N_6150);
nand U7178 (N_7178,N_6483,N_6395);
or U7179 (N_7179,N_6576,N_6109);
nor U7180 (N_7180,N_6857,N_6058);
nor U7181 (N_7181,N_6464,N_6850);
nor U7182 (N_7182,N_6986,N_6732);
nand U7183 (N_7183,N_6265,N_6949);
and U7184 (N_7184,N_6783,N_6421);
nor U7185 (N_7185,N_6969,N_6985);
and U7186 (N_7186,N_6838,N_6033);
nor U7187 (N_7187,N_6972,N_6009);
nor U7188 (N_7188,N_6437,N_6627);
and U7189 (N_7189,N_6281,N_6766);
xnor U7190 (N_7190,N_6539,N_6892);
nand U7191 (N_7191,N_6328,N_6891);
and U7192 (N_7192,N_6854,N_6359);
nand U7193 (N_7193,N_6386,N_6880);
nand U7194 (N_7194,N_6135,N_6476);
or U7195 (N_7195,N_6151,N_6490);
and U7196 (N_7196,N_6523,N_6154);
or U7197 (N_7197,N_6214,N_6489);
and U7198 (N_7198,N_6097,N_6625);
xnor U7199 (N_7199,N_6202,N_6677);
nand U7200 (N_7200,N_6017,N_6782);
nor U7201 (N_7201,N_6813,N_6723);
nor U7202 (N_7202,N_6360,N_6108);
nor U7203 (N_7203,N_6345,N_6606);
xor U7204 (N_7204,N_6951,N_6072);
and U7205 (N_7205,N_6102,N_6225);
xnor U7206 (N_7206,N_6267,N_6966);
nand U7207 (N_7207,N_6511,N_6454);
nor U7208 (N_7208,N_6324,N_6654);
xnor U7209 (N_7209,N_6453,N_6902);
and U7210 (N_7210,N_6997,N_6552);
nor U7211 (N_7211,N_6292,N_6242);
xnor U7212 (N_7212,N_6482,N_6194);
nor U7213 (N_7213,N_6882,N_6990);
nand U7214 (N_7214,N_6823,N_6182);
nand U7215 (N_7215,N_6010,N_6197);
or U7216 (N_7216,N_6587,N_6031);
xnor U7217 (N_7217,N_6193,N_6280);
and U7218 (N_7218,N_6391,N_6034);
nor U7219 (N_7219,N_6500,N_6466);
and U7220 (N_7220,N_6956,N_6048);
and U7221 (N_7221,N_6538,N_6465);
nand U7222 (N_7222,N_6704,N_6356);
xnor U7223 (N_7223,N_6939,N_6933);
and U7224 (N_7224,N_6308,N_6534);
nand U7225 (N_7225,N_6778,N_6025);
or U7226 (N_7226,N_6407,N_6405);
and U7227 (N_7227,N_6355,N_6820);
nor U7228 (N_7228,N_6977,N_6252);
and U7229 (N_7229,N_6731,N_6545);
nand U7230 (N_7230,N_6896,N_6826);
and U7231 (N_7231,N_6609,N_6215);
xor U7232 (N_7232,N_6622,N_6189);
or U7233 (N_7233,N_6871,N_6873);
or U7234 (N_7234,N_6507,N_6501);
nor U7235 (N_7235,N_6563,N_6716);
nand U7236 (N_7236,N_6463,N_6403);
nor U7237 (N_7237,N_6053,N_6041);
nor U7238 (N_7238,N_6847,N_6856);
or U7239 (N_7239,N_6100,N_6136);
and U7240 (N_7240,N_6379,N_6779);
and U7241 (N_7241,N_6825,N_6572);
or U7242 (N_7242,N_6945,N_6814);
nor U7243 (N_7243,N_6247,N_6149);
and U7244 (N_7244,N_6043,N_6219);
or U7245 (N_7245,N_6146,N_6897);
nand U7246 (N_7246,N_6414,N_6030);
nor U7247 (N_7247,N_6460,N_6529);
or U7248 (N_7248,N_6164,N_6115);
and U7249 (N_7249,N_6960,N_6012);
nor U7250 (N_7250,N_6519,N_6383);
nand U7251 (N_7251,N_6709,N_6060);
nand U7252 (N_7252,N_6708,N_6289);
nand U7253 (N_7253,N_6192,N_6469);
or U7254 (N_7254,N_6132,N_6746);
and U7255 (N_7255,N_6687,N_6600);
xor U7256 (N_7256,N_6799,N_6660);
nand U7257 (N_7257,N_6608,N_6208);
and U7258 (N_7258,N_6839,N_6374);
nand U7259 (N_7259,N_6351,N_6932);
and U7260 (N_7260,N_6505,N_6741);
xor U7261 (N_7261,N_6236,N_6389);
and U7262 (N_7262,N_6874,N_6297);
nand U7263 (N_7263,N_6527,N_6221);
nand U7264 (N_7264,N_6063,N_6755);
nand U7265 (N_7265,N_6094,N_6751);
nor U7266 (N_7266,N_6690,N_6994);
or U7267 (N_7267,N_6964,N_6255);
xnor U7268 (N_7268,N_6714,N_6901);
nor U7269 (N_7269,N_6584,N_6264);
or U7270 (N_7270,N_6618,N_6636);
xnor U7271 (N_7271,N_6626,N_6096);
nor U7272 (N_7272,N_6947,N_6548);
or U7273 (N_7273,N_6275,N_6435);
or U7274 (N_7274,N_6816,N_6162);
and U7275 (N_7275,N_6513,N_6557);
and U7276 (N_7276,N_6305,N_6551);
and U7277 (N_7277,N_6293,N_6312);
nor U7278 (N_7278,N_6655,N_6152);
and U7279 (N_7279,N_6546,N_6331);
nand U7280 (N_7280,N_6493,N_6644);
and U7281 (N_7281,N_6672,N_6988);
xor U7282 (N_7282,N_6982,N_6509);
xor U7283 (N_7283,N_6589,N_6842);
nand U7284 (N_7284,N_6802,N_6125);
xor U7285 (N_7285,N_6886,N_6450);
nor U7286 (N_7286,N_6226,N_6446);
nand U7287 (N_7287,N_6228,N_6971);
nor U7288 (N_7288,N_6368,N_6190);
and U7289 (N_7289,N_6669,N_6670);
nand U7290 (N_7290,N_6818,N_6694);
nand U7291 (N_7291,N_6767,N_6567);
and U7292 (N_7292,N_6931,N_6647);
xnor U7293 (N_7293,N_6353,N_6643);
nand U7294 (N_7294,N_6721,N_6423);
nor U7295 (N_7295,N_6571,N_6544);
and U7296 (N_7296,N_6645,N_6090);
xor U7297 (N_7297,N_6262,N_6667);
or U7298 (N_7298,N_6565,N_6558);
nor U7299 (N_7299,N_6245,N_6616);
nor U7300 (N_7300,N_6087,N_6001);
and U7301 (N_7301,N_6834,N_6455);
nand U7302 (N_7302,N_6054,N_6628);
and U7303 (N_7303,N_6251,N_6384);
nand U7304 (N_7304,N_6605,N_6467);
or U7305 (N_7305,N_6110,N_6123);
nand U7306 (N_7306,N_6438,N_6357);
and U7307 (N_7307,N_6307,N_6770);
nor U7308 (N_7308,N_6968,N_6592);
nor U7309 (N_7309,N_6760,N_6747);
and U7310 (N_7310,N_6686,N_6475);
xnor U7311 (N_7311,N_6794,N_6841);
xnor U7312 (N_7312,N_6678,N_6953);
nor U7313 (N_7313,N_6091,N_6805);
or U7314 (N_7314,N_6697,N_6691);
xnor U7315 (N_7315,N_6865,N_6165);
nand U7316 (N_7316,N_6713,N_6321);
and U7317 (N_7317,N_6568,N_6967);
nor U7318 (N_7318,N_6008,N_6344);
and U7319 (N_7319,N_6996,N_6040);
nor U7320 (N_7320,N_6754,N_6617);
nand U7321 (N_7321,N_6266,N_6451);
and U7322 (N_7322,N_6583,N_6954);
nor U7323 (N_7323,N_6578,N_6676);
nor U7324 (N_7324,N_6700,N_6952);
xor U7325 (N_7325,N_6046,N_6349);
or U7326 (N_7326,N_6581,N_6877);
xnor U7327 (N_7327,N_6430,N_6431);
or U7328 (N_7328,N_6122,N_6883);
and U7329 (N_7329,N_6893,N_6473);
xor U7330 (N_7330,N_6566,N_6478);
and U7331 (N_7331,N_6810,N_6699);
nand U7332 (N_7332,N_6531,N_6320);
nand U7333 (N_7333,N_6216,N_6153);
and U7334 (N_7334,N_6057,N_6409);
nor U7335 (N_7335,N_6607,N_6744);
and U7336 (N_7336,N_6301,N_6160);
or U7337 (N_7337,N_6124,N_6047);
nand U7338 (N_7338,N_6532,N_6365);
nor U7339 (N_7339,N_6333,N_6946);
xnor U7340 (N_7340,N_6470,N_6411);
nand U7341 (N_7341,N_6804,N_6378);
and U7342 (N_7342,N_6448,N_6481);
xnor U7343 (N_7343,N_6696,N_6230);
xor U7344 (N_7344,N_6503,N_6749);
and U7345 (N_7345,N_6978,N_6598);
nand U7346 (N_7346,N_6638,N_6329);
or U7347 (N_7347,N_6615,N_6632);
nor U7348 (N_7348,N_6218,N_6750);
nand U7349 (N_7349,N_6120,N_6496);
nand U7350 (N_7350,N_6706,N_6619);
nand U7351 (N_7351,N_6903,N_6449);
or U7352 (N_7352,N_6510,N_6906);
nand U7353 (N_7353,N_6683,N_6950);
nand U7354 (N_7354,N_6147,N_6232);
or U7355 (N_7355,N_6440,N_6027);
nor U7356 (N_7356,N_6186,N_6397);
or U7357 (N_7357,N_6268,N_6354);
xnor U7358 (N_7358,N_6082,N_6248);
and U7359 (N_7359,N_6037,N_6195);
and U7360 (N_7360,N_6098,N_6852);
nand U7361 (N_7361,N_6914,N_6071);
xor U7362 (N_7362,N_6302,N_6807);
and U7363 (N_7363,N_6070,N_6595);
nand U7364 (N_7364,N_6541,N_6844);
nor U7365 (N_7365,N_6588,N_6853);
and U7366 (N_7366,N_6433,N_6811);
nor U7367 (N_7367,N_6929,N_6362);
or U7368 (N_7368,N_6169,N_6114);
nand U7369 (N_7369,N_6300,N_6367);
nand U7370 (N_7370,N_6594,N_6858);
nor U7371 (N_7371,N_6249,N_6144);
nand U7372 (N_7372,N_6410,N_6611);
and U7373 (N_7373,N_6073,N_6056);
nor U7374 (N_7374,N_6803,N_6083);
nand U7375 (N_7375,N_6943,N_6006);
nor U7376 (N_7376,N_6126,N_6878);
nor U7377 (N_7377,N_6304,N_6042);
or U7378 (N_7378,N_6635,N_6432);
or U7379 (N_7379,N_6269,N_6341);
xor U7380 (N_7380,N_6681,N_6288);
or U7381 (N_7381,N_6085,N_6832);
nand U7382 (N_7382,N_6601,N_6771);
nand U7383 (N_7383,N_6497,N_6915);
and U7384 (N_7384,N_6517,N_6176);
nor U7385 (N_7385,N_6427,N_6061);
and U7386 (N_7386,N_6178,N_6522);
nor U7387 (N_7387,N_6111,N_6917);
and U7388 (N_7388,N_6434,N_6879);
nand U7389 (N_7389,N_6077,N_6387);
nand U7390 (N_7390,N_6143,N_6452);
nor U7391 (N_7391,N_6444,N_6059);
or U7392 (N_7392,N_6286,N_6313);
nand U7393 (N_7393,N_6103,N_6712);
and U7394 (N_7394,N_6928,N_6965);
xor U7395 (N_7395,N_6734,N_6170);
nand U7396 (N_7396,N_6375,N_6705);
xnor U7397 (N_7397,N_6537,N_6326);
xnor U7398 (N_7398,N_6506,N_6020);
or U7399 (N_7399,N_6787,N_6562);
and U7400 (N_7400,N_6614,N_6417);
nand U7401 (N_7401,N_6134,N_6642);
and U7402 (N_7402,N_6999,N_6062);
nand U7403 (N_7403,N_6235,N_6336);
or U7404 (N_7404,N_6675,N_6909);
nand U7405 (N_7405,N_6797,N_6756);
and U7406 (N_7406,N_6524,N_6637);
or U7407 (N_7407,N_6260,N_6610);
nand U7408 (N_7408,N_6284,N_6582);
xor U7409 (N_7409,N_6762,N_6198);
nor U7410 (N_7410,N_6347,N_6210);
nor U7411 (N_7411,N_6861,N_6508);
and U7412 (N_7412,N_6002,N_6045);
and U7413 (N_7413,N_6332,N_6340);
nand U7414 (N_7414,N_6682,N_6283);
nor U7415 (N_7415,N_6656,N_6666);
nor U7416 (N_7416,N_6575,N_6105);
nand U7417 (N_7417,N_6428,N_6639);
and U7418 (N_7418,N_6671,N_6729);
and U7419 (N_7419,N_6079,N_6067);
or U7420 (N_7420,N_6742,N_6394);
nand U7421 (N_7421,N_6798,N_6204);
nor U7422 (N_7422,N_6796,N_6995);
nand U7423 (N_7423,N_6240,N_6835);
xnor U7424 (N_7424,N_6570,N_6740);
or U7425 (N_7425,N_6217,N_6764);
or U7426 (N_7426,N_6525,N_6973);
nor U7427 (N_7427,N_6591,N_6889);
nor U7428 (N_7428,N_6184,N_6640);
or U7429 (N_7429,N_6000,N_6630);
or U7430 (N_7430,N_6243,N_6733);
xnor U7431 (N_7431,N_6648,N_6166);
nand U7432 (N_7432,N_6634,N_6180);
and U7433 (N_7433,N_6229,N_6757);
nand U7434 (N_7434,N_6238,N_6499);
nor U7435 (N_7435,N_6139,N_6812);
xnor U7436 (N_7436,N_6343,N_6201);
nor U7437 (N_7437,N_6979,N_6707);
nor U7438 (N_7438,N_6815,N_6393);
and U7439 (N_7439,N_6876,N_6801);
nand U7440 (N_7440,N_6559,N_6586);
nand U7441 (N_7441,N_6718,N_6233);
nand U7442 (N_7442,N_6363,N_6196);
or U7443 (N_7443,N_6658,N_6603);
nand U7444 (N_7444,N_6612,N_6597);
nor U7445 (N_7445,N_6156,N_6937);
and U7446 (N_7446,N_6259,N_6817);
nand U7447 (N_7447,N_6327,N_6765);
and U7448 (N_7448,N_6298,N_6429);
or U7449 (N_7449,N_6961,N_6335);
or U7450 (N_7450,N_6872,N_6819);
nor U7451 (N_7451,N_6200,N_6573);
nand U7452 (N_7452,N_6052,N_6024);
and U7453 (N_7453,N_6282,N_6127);
xnor U7454 (N_7454,N_6171,N_6213);
and U7455 (N_7455,N_6955,N_6019);
and U7456 (N_7456,N_6845,N_6064);
and U7457 (N_7457,N_6413,N_6739);
or U7458 (N_7458,N_6907,N_6726);
nor U7459 (N_7459,N_6863,N_6673);
or U7460 (N_7460,N_6477,N_6254);
nand U7461 (N_7461,N_6246,N_6104);
nor U7462 (N_7462,N_6992,N_6209);
or U7463 (N_7463,N_6836,N_6989);
and U7464 (N_7464,N_6824,N_6309);
nor U7465 (N_7465,N_6604,N_6887);
or U7466 (N_7466,N_6922,N_6018);
and U7467 (N_7467,N_6011,N_6828);
or U7468 (N_7468,N_6515,N_6540);
nor U7469 (N_7469,N_6487,N_6484);
or U7470 (N_7470,N_6220,N_6148);
or U7471 (N_7471,N_6459,N_6342);
and U7472 (N_7472,N_6080,N_6848);
nand U7473 (N_7473,N_6338,N_6366);
and U7474 (N_7474,N_6894,N_6199);
nand U7475 (N_7475,N_6692,N_6422);
xnor U7476 (N_7476,N_6174,N_6786);
nand U7477 (N_7477,N_6924,N_6485);
and U7478 (N_7478,N_6788,N_6495);
nor U7479 (N_7479,N_6461,N_6502);
and U7480 (N_7480,N_6602,N_6735);
and U7481 (N_7481,N_6263,N_6621);
xor U7482 (N_7482,N_6987,N_6518);
or U7483 (N_7483,N_6480,N_6769);
nor U7484 (N_7484,N_6258,N_6975);
nor U7485 (N_7485,N_6958,N_6795);
or U7486 (N_7486,N_6093,N_6290);
nor U7487 (N_7487,N_6279,N_6984);
or U7488 (N_7488,N_6222,N_6881);
and U7489 (N_7489,N_6535,N_6179);
or U7490 (N_7490,N_6547,N_6846);
xnor U7491 (N_7491,N_6227,N_6049);
nor U7492 (N_7492,N_6107,N_6112);
or U7493 (N_7493,N_6092,N_6404);
nor U7494 (N_7494,N_6442,N_6504);
xnor U7495 (N_7495,N_6348,N_6408);
or U7496 (N_7496,N_6725,N_6821);
and U7497 (N_7497,N_6381,N_6231);
and U7498 (N_7498,N_6743,N_6859);
nor U7499 (N_7499,N_6088,N_6244);
nor U7500 (N_7500,N_6704,N_6054);
and U7501 (N_7501,N_6931,N_6319);
nand U7502 (N_7502,N_6641,N_6959);
nor U7503 (N_7503,N_6637,N_6669);
and U7504 (N_7504,N_6995,N_6695);
nor U7505 (N_7505,N_6880,N_6244);
and U7506 (N_7506,N_6633,N_6257);
or U7507 (N_7507,N_6997,N_6017);
or U7508 (N_7508,N_6450,N_6225);
and U7509 (N_7509,N_6634,N_6694);
xor U7510 (N_7510,N_6734,N_6470);
and U7511 (N_7511,N_6123,N_6809);
and U7512 (N_7512,N_6809,N_6829);
nand U7513 (N_7513,N_6121,N_6071);
nor U7514 (N_7514,N_6653,N_6370);
nor U7515 (N_7515,N_6748,N_6528);
nor U7516 (N_7516,N_6071,N_6667);
or U7517 (N_7517,N_6461,N_6407);
or U7518 (N_7518,N_6506,N_6833);
nor U7519 (N_7519,N_6384,N_6239);
or U7520 (N_7520,N_6005,N_6275);
nand U7521 (N_7521,N_6606,N_6577);
nor U7522 (N_7522,N_6205,N_6262);
xnor U7523 (N_7523,N_6578,N_6858);
or U7524 (N_7524,N_6597,N_6834);
nand U7525 (N_7525,N_6104,N_6201);
nand U7526 (N_7526,N_6945,N_6618);
and U7527 (N_7527,N_6900,N_6192);
nand U7528 (N_7528,N_6562,N_6457);
or U7529 (N_7529,N_6310,N_6009);
and U7530 (N_7530,N_6960,N_6356);
and U7531 (N_7531,N_6625,N_6972);
nand U7532 (N_7532,N_6256,N_6669);
xnor U7533 (N_7533,N_6393,N_6271);
or U7534 (N_7534,N_6242,N_6732);
and U7535 (N_7535,N_6608,N_6042);
xnor U7536 (N_7536,N_6361,N_6049);
nand U7537 (N_7537,N_6473,N_6517);
or U7538 (N_7538,N_6060,N_6840);
or U7539 (N_7539,N_6467,N_6194);
and U7540 (N_7540,N_6267,N_6802);
and U7541 (N_7541,N_6348,N_6244);
nor U7542 (N_7542,N_6809,N_6979);
nor U7543 (N_7543,N_6489,N_6538);
nand U7544 (N_7544,N_6434,N_6374);
nand U7545 (N_7545,N_6640,N_6683);
nor U7546 (N_7546,N_6453,N_6719);
nor U7547 (N_7547,N_6547,N_6493);
or U7548 (N_7548,N_6394,N_6034);
or U7549 (N_7549,N_6682,N_6051);
or U7550 (N_7550,N_6204,N_6505);
nand U7551 (N_7551,N_6524,N_6489);
nand U7552 (N_7552,N_6710,N_6451);
nand U7553 (N_7553,N_6011,N_6912);
nand U7554 (N_7554,N_6050,N_6853);
and U7555 (N_7555,N_6031,N_6173);
nor U7556 (N_7556,N_6513,N_6864);
and U7557 (N_7557,N_6580,N_6554);
nor U7558 (N_7558,N_6619,N_6348);
and U7559 (N_7559,N_6512,N_6920);
xor U7560 (N_7560,N_6058,N_6976);
nand U7561 (N_7561,N_6733,N_6480);
or U7562 (N_7562,N_6249,N_6624);
nand U7563 (N_7563,N_6529,N_6465);
nand U7564 (N_7564,N_6687,N_6408);
nor U7565 (N_7565,N_6269,N_6791);
nand U7566 (N_7566,N_6538,N_6105);
nor U7567 (N_7567,N_6807,N_6706);
nor U7568 (N_7568,N_6724,N_6615);
and U7569 (N_7569,N_6942,N_6456);
nor U7570 (N_7570,N_6751,N_6547);
nor U7571 (N_7571,N_6926,N_6505);
nor U7572 (N_7572,N_6879,N_6945);
or U7573 (N_7573,N_6967,N_6422);
nor U7574 (N_7574,N_6766,N_6484);
and U7575 (N_7575,N_6855,N_6562);
or U7576 (N_7576,N_6263,N_6066);
or U7577 (N_7577,N_6704,N_6458);
xnor U7578 (N_7578,N_6183,N_6840);
and U7579 (N_7579,N_6719,N_6313);
nor U7580 (N_7580,N_6866,N_6264);
and U7581 (N_7581,N_6771,N_6375);
nand U7582 (N_7582,N_6629,N_6926);
nand U7583 (N_7583,N_6286,N_6495);
nand U7584 (N_7584,N_6546,N_6444);
xor U7585 (N_7585,N_6024,N_6582);
or U7586 (N_7586,N_6468,N_6492);
or U7587 (N_7587,N_6040,N_6806);
and U7588 (N_7588,N_6919,N_6697);
xor U7589 (N_7589,N_6859,N_6598);
xnor U7590 (N_7590,N_6333,N_6987);
or U7591 (N_7591,N_6732,N_6749);
and U7592 (N_7592,N_6053,N_6455);
xor U7593 (N_7593,N_6728,N_6925);
xnor U7594 (N_7594,N_6283,N_6217);
nand U7595 (N_7595,N_6737,N_6397);
nand U7596 (N_7596,N_6310,N_6692);
or U7597 (N_7597,N_6719,N_6109);
nand U7598 (N_7598,N_6924,N_6900);
or U7599 (N_7599,N_6084,N_6299);
and U7600 (N_7600,N_6898,N_6509);
nor U7601 (N_7601,N_6105,N_6154);
xnor U7602 (N_7602,N_6823,N_6591);
or U7603 (N_7603,N_6804,N_6267);
and U7604 (N_7604,N_6117,N_6757);
xnor U7605 (N_7605,N_6700,N_6486);
nor U7606 (N_7606,N_6079,N_6837);
and U7607 (N_7607,N_6691,N_6386);
or U7608 (N_7608,N_6573,N_6653);
nand U7609 (N_7609,N_6903,N_6493);
nor U7610 (N_7610,N_6146,N_6572);
and U7611 (N_7611,N_6703,N_6481);
nand U7612 (N_7612,N_6488,N_6235);
nor U7613 (N_7613,N_6061,N_6648);
nor U7614 (N_7614,N_6204,N_6396);
or U7615 (N_7615,N_6265,N_6067);
nor U7616 (N_7616,N_6877,N_6156);
nand U7617 (N_7617,N_6811,N_6259);
nor U7618 (N_7618,N_6968,N_6463);
and U7619 (N_7619,N_6649,N_6170);
and U7620 (N_7620,N_6368,N_6320);
nand U7621 (N_7621,N_6561,N_6249);
and U7622 (N_7622,N_6100,N_6001);
xor U7623 (N_7623,N_6402,N_6759);
and U7624 (N_7624,N_6125,N_6183);
or U7625 (N_7625,N_6576,N_6030);
and U7626 (N_7626,N_6546,N_6303);
and U7627 (N_7627,N_6308,N_6413);
nand U7628 (N_7628,N_6013,N_6997);
or U7629 (N_7629,N_6963,N_6669);
xnor U7630 (N_7630,N_6339,N_6382);
nor U7631 (N_7631,N_6952,N_6240);
nor U7632 (N_7632,N_6893,N_6022);
and U7633 (N_7633,N_6198,N_6488);
nand U7634 (N_7634,N_6603,N_6513);
xor U7635 (N_7635,N_6276,N_6974);
or U7636 (N_7636,N_6160,N_6224);
nor U7637 (N_7637,N_6695,N_6434);
nand U7638 (N_7638,N_6917,N_6853);
xnor U7639 (N_7639,N_6992,N_6174);
nor U7640 (N_7640,N_6521,N_6848);
or U7641 (N_7641,N_6515,N_6397);
and U7642 (N_7642,N_6561,N_6784);
nand U7643 (N_7643,N_6955,N_6805);
and U7644 (N_7644,N_6070,N_6425);
nand U7645 (N_7645,N_6460,N_6545);
or U7646 (N_7646,N_6337,N_6925);
nor U7647 (N_7647,N_6400,N_6063);
xor U7648 (N_7648,N_6094,N_6615);
and U7649 (N_7649,N_6045,N_6039);
xnor U7650 (N_7650,N_6892,N_6227);
or U7651 (N_7651,N_6955,N_6032);
nor U7652 (N_7652,N_6222,N_6323);
nand U7653 (N_7653,N_6335,N_6324);
xnor U7654 (N_7654,N_6497,N_6156);
and U7655 (N_7655,N_6457,N_6499);
xnor U7656 (N_7656,N_6545,N_6072);
nor U7657 (N_7657,N_6557,N_6850);
or U7658 (N_7658,N_6645,N_6809);
or U7659 (N_7659,N_6422,N_6436);
or U7660 (N_7660,N_6035,N_6904);
xnor U7661 (N_7661,N_6799,N_6487);
nor U7662 (N_7662,N_6609,N_6733);
and U7663 (N_7663,N_6080,N_6862);
and U7664 (N_7664,N_6068,N_6617);
nand U7665 (N_7665,N_6762,N_6019);
nand U7666 (N_7666,N_6368,N_6867);
xor U7667 (N_7667,N_6078,N_6260);
nand U7668 (N_7668,N_6370,N_6548);
and U7669 (N_7669,N_6519,N_6938);
and U7670 (N_7670,N_6719,N_6953);
or U7671 (N_7671,N_6765,N_6810);
or U7672 (N_7672,N_6127,N_6607);
nor U7673 (N_7673,N_6796,N_6836);
and U7674 (N_7674,N_6577,N_6944);
or U7675 (N_7675,N_6275,N_6225);
nand U7676 (N_7676,N_6275,N_6085);
nand U7677 (N_7677,N_6306,N_6561);
nand U7678 (N_7678,N_6675,N_6516);
nand U7679 (N_7679,N_6987,N_6250);
nor U7680 (N_7680,N_6938,N_6143);
xnor U7681 (N_7681,N_6250,N_6902);
nor U7682 (N_7682,N_6969,N_6414);
and U7683 (N_7683,N_6020,N_6066);
nand U7684 (N_7684,N_6225,N_6939);
and U7685 (N_7685,N_6606,N_6548);
nand U7686 (N_7686,N_6629,N_6017);
nor U7687 (N_7687,N_6174,N_6772);
and U7688 (N_7688,N_6670,N_6278);
xnor U7689 (N_7689,N_6366,N_6816);
xnor U7690 (N_7690,N_6403,N_6566);
nand U7691 (N_7691,N_6830,N_6675);
nand U7692 (N_7692,N_6396,N_6213);
or U7693 (N_7693,N_6985,N_6062);
and U7694 (N_7694,N_6790,N_6991);
nand U7695 (N_7695,N_6479,N_6098);
nand U7696 (N_7696,N_6913,N_6462);
or U7697 (N_7697,N_6787,N_6085);
and U7698 (N_7698,N_6441,N_6453);
nor U7699 (N_7699,N_6827,N_6867);
nand U7700 (N_7700,N_6512,N_6317);
nand U7701 (N_7701,N_6409,N_6872);
xnor U7702 (N_7702,N_6547,N_6359);
nand U7703 (N_7703,N_6422,N_6160);
and U7704 (N_7704,N_6156,N_6367);
nand U7705 (N_7705,N_6257,N_6895);
and U7706 (N_7706,N_6601,N_6704);
or U7707 (N_7707,N_6692,N_6596);
or U7708 (N_7708,N_6208,N_6958);
nand U7709 (N_7709,N_6246,N_6114);
or U7710 (N_7710,N_6163,N_6559);
and U7711 (N_7711,N_6041,N_6655);
nor U7712 (N_7712,N_6987,N_6101);
or U7713 (N_7713,N_6573,N_6354);
nand U7714 (N_7714,N_6434,N_6502);
nor U7715 (N_7715,N_6737,N_6673);
and U7716 (N_7716,N_6581,N_6541);
nor U7717 (N_7717,N_6636,N_6496);
nor U7718 (N_7718,N_6901,N_6318);
nor U7719 (N_7719,N_6852,N_6518);
or U7720 (N_7720,N_6664,N_6166);
nor U7721 (N_7721,N_6020,N_6178);
nor U7722 (N_7722,N_6792,N_6886);
or U7723 (N_7723,N_6441,N_6495);
or U7724 (N_7724,N_6062,N_6567);
nor U7725 (N_7725,N_6760,N_6930);
xnor U7726 (N_7726,N_6068,N_6790);
nor U7727 (N_7727,N_6078,N_6043);
nor U7728 (N_7728,N_6098,N_6485);
nand U7729 (N_7729,N_6408,N_6400);
xor U7730 (N_7730,N_6451,N_6237);
nor U7731 (N_7731,N_6022,N_6908);
nor U7732 (N_7732,N_6305,N_6401);
nor U7733 (N_7733,N_6624,N_6938);
nor U7734 (N_7734,N_6584,N_6897);
or U7735 (N_7735,N_6863,N_6342);
nor U7736 (N_7736,N_6340,N_6620);
or U7737 (N_7737,N_6549,N_6062);
nor U7738 (N_7738,N_6463,N_6365);
and U7739 (N_7739,N_6293,N_6572);
nor U7740 (N_7740,N_6293,N_6440);
nor U7741 (N_7741,N_6430,N_6087);
xor U7742 (N_7742,N_6575,N_6583);
or U7743 (N_7743,N_6058,N_6045);
nor U7744 (N_7744,N_6425,N_6602);
and U7745 (N_7745,N_6102,N_6717);
nand U7746 (N_7746,N_6549,N_6661);
and U7747 (N_7747,N_6489,N_6468);
nand U7748 (N_7748,N_6110,N_6191);
and U7749 (N_7749,N_6612,N_6829);
or U7750 (N_7750,N_6332,N_6520);
or U7751 (N_7751,N_6796,N_6406);
nand U7752 (N_7752,N_6808,N_6659);
nand U7753 (N_7753,N_6324,N_6523);
or U7754 (N_7754,N_6319,N_6087);
nand U7755 (N_7755,N_6962,N_6396);
nor U7756 (N_7756,N_6916,N_6676);
nand U7757 (N_7757,N_6749,N_6635);
nor U7758 (N_7758,N_6162,N_6922);
xnor U7759 (N_7759,N_6430,N_6924);
nor U7760 (N_7760,N_6816,N_6583);
xnor U7761 (N_7761,N_6031,N_6405);
and U7762 (N_7762,N_6036,N_6460);
and U7763 (N_7763,N_6053,N_6600);
nand U7764 (N_7764,N_6492,N_6949);
or U7765 (N_7765,N_6520,N_6061);
and U7766 (N_7766,N_6017,N_6949);
or U7767 (N_7767,N_6253,N_6087);
xor U7768 (N_7768,N_6886,N_6287);
or U7769 (N_7769,N_6353,N_6862);
nand U7770 (N_7770,N_6724,N_6698);
nand U7771 (N_7771,N_6144,N_6411);
or U7772 (N_7772,N_6360,N_6862);
xor U7773 (N_7773,N_6438,N_6352);
nand U7774 (N_7774,N_6693,N_6316);
or U7775 (N_7775,N_6175,N_6191);
nand U7776 (N_7776,N_6209,N_6666);
and U7777 (N_7777,N_6142,N_6282);
or U7778 (N_7778,N_6855,N_6214);
and U7779 (N_7779,N_6192,N_6884);
nor U7780 (N_7780,N_6117,N_6069);
or U7781 (N_7781,N_6424,N_6427);
nand U7782 (N_7782,N_6540,N_6513);
xor U7783 (N_7783,N_6898,N_6209);
nand U7784 (N_7784,N_6061,N_6160);
or U7785 (N_7785,N_6975,N_6837);
nor U7786 (N_7786,N_6033,N_6780);
nand U7787 (N_7787,N_6586,N_6268);
xor U7788 (N_7788,N_6485,N_6779);
xnor U7789 (N_7789,N_6072,N_6986);
nand U7790 (N_7790,N_6138,N_6399);
xnor U7791 (N_7791,N_6648,N_6733);
nor U7792 (N_7792,N_6299,N_6088);
or U7793 (N_7793,N_6566,N_6837);
nand U7794 (N_7794,N_6352,N_6807);
and U7795 (N_7795,N_6293,N_6727);
nand U7796 (N_7796,N_6710,N_6745);
and U7797 (N_7797,N_6242,N_6837);
nand U7798 (N_7798,N_6075,N_6992);
or U7799 (N_7799,N_6108,N_6747);
nor U7800 (N_7800,N_6368,N_6533);
nor U7801 (N_7801,N_6348,N_6627);
nor U7802 (N_7802,N_6117,N_6070);
nand U7803 (N_7803,N_6220,N_6817);
and U7804 (N_7804,N_6390,N_6481);
nor U7805 (N_7805,N_6448,N_6647);
and U7806 (N_7806,N_6945,N_6259);
and U7807 (N_7807,N_6855,N_6017);
or U7808 (N_7808,N_6310,N_6811);
and U7809 (N_7809,N_6981,N_6483);
and U7810 (N_7810,N_6215,N_6966);
or U7811 (N_7811,N_6398,N_6939);
nand U7812 (N_7812,N_6383,N_6154);
nor U7813 (N_7813,N_6385,N_6935);
nand U7814 (N_7814,N_6345,N_6631);
xor U7815 (N_7815,N_6302,N_6869);
and U7816 (N_7816,N_6521,N_6074);
nor U7817 (N_7817,N_6772,N_6106);
nand U7818 (N_7818,N_6768,N_6468);
nor U7819 (N_7819,N_6605,N_6366);
nor U7820 (N_7820,N_6536,N_6581);
or U7821 (N_7821,N_6452,N_6809);
nor U7822 (N_7822,N_6596,N_6377);
nor U7823 (N_7823,N_6185,N_6229);
xor U7824 (N_7824,N_6991,N_6985);
xor U7825 (N_7825,N_6446,N_6135);
xnor U7826 (N_7826,N_6618,N_6559);
nor U7827 (N_7827,N_6559,N_6797);
or U7828 (N_7828,N_6217,N_6046);
nand U7829 (N_7829,N_6675,N_6548);
or U7830 (N_7830,N_6507,N_6667);
and U7831 (N_7831,N_6509,N_6334);
or U7832 (N_7832,N_6380,N_6507);
and U7833 (N_7833,N_6981,N_6334);
nor U7834 (N_7834,N_6074,N_6978);
nand U7835 (N_7835,N_6825,N_6877);
xor U7836 (N_7836,N_6412,N_6698);
nor U7837 (N_7837,N_6342,N_6952);
or U7838 (N_7838,N_6067,N_6813);
nor U7839 (N_7839,N_6605,N_6552);
nand U7840 (N_7840,N_6344,N_6043);
nand U7841 (N_7841,N_6541,N_6933);
and U7842 (N_7842,N_6949,N_6237);
and U7843 (N_7843,N_6993,N_6927);
nor U7844 (N_7844,N_6917,N_6143);
nand U7845 (N_7845,N_6417,N_6802);
or U7846 (N_7846,N_6200,N_6044);
or U7847 (N_7847,N_6942,N_6541);
or U7848 (N_7848,N_6861,N_6846);
or U7849 (N_7849,N_6505,N_6465);
or U7850 (N_7850,N_6918,N_6505);
or U7851 (N_7851,N_6372,N_6811);
or U7852 (N_7852,N_6593,N_6300);
nand U7853 (N_7853,N_6348,N_6433);
or U7854 (N_7854,N_6594,N_6183);
nor U7855 (N_7855,N_6102,N_6841);
nand U7856 (N_7856,N_6676,N_6405);
nand U7857 (N_7857,N_6118,N_6291);
or U7858 (N_7858,N_6639,N_6777);
nand U7859 (N_7859,N_6467,N_6206);
and U7860 (N_7860,N_6205,N_6834);
and U7861 (N_7861,N_6883,N_6030);
nor U7862 (N_7862,N_6944,N_6766);
nor U7863 (N_7863,N_6635,N_6325);
or U7864 (N_7864,N_6149,N_6828);
or U7865 (N_7865,N_6145,N_6174);
nand U7866 (N_7866,N_6512,N_6403);
and U7867 (N_7867,N_6747,N_6267);
and U7868 (N_7868,N_6184,N_6000);
nand U7869 (N_7869,N_6366,N_6927);
and U7870 (N_7870,N_6660,N_6670);
or U7871 (N_7871,N_6176,N_6364);
nor U7872 (N_7872,N_6530,N_6478);
nor U7873 (N_7873,N_6916,N_6101);
nand U7874 (N_7874,N_6885,N_6718);
or U7875 (N_7875,N_6974,N_6512);
nor U7876 (N_7876,N_6548,N_6112);
nand U7877 (N_7877,N_6166,N_6921);
and U7878 (N_7878,N_6144,N_6456);
nand U7879 (N_7879,N_6136,N_6030);
or U7880 (N_7880,N_6813,N_6665);
or U7881 (N_7881,N_6101,N_6553);
xnor U7882 (N_7882,N_6839,N_6723);
nor U7883 (N_7883,N_6956,N_6120);
or U7884 (N_7884,N_6730,N_6795);
nor U7885 (N_7885,N_6476,N_6251);
and U7886 (N_7886,N_6151,N_6236);
nand U7887 (N_7887,N_6081,N_6726);
nand U7888 (N_7888,N_6171,N_6834);
or U7889 (N_7889,N_6357,N_6756);
and U7890 (N_7890,N_6420,N_6323);
nor U7891 (N_7891,N_6642,N_6469);
or U7892 (N_7892,N_6739,N_6429);
and U7893 (N_7893,N_6933,N_6623);
or U7894 (N_7894,N_6274,N_6876);
and U7895 (N_7895,N_6230,N_6358);
nor U7896 (N_7896,N_6097,N_6444);
and U7897 (N_7897,N_6977,N_6753);
nand U7898 (N_7898,N_6104,N_6807);
and U7899 (N_7899,N_6701,N_6804);
and U7900 (N_7900,N_6598,N_6841);
nand U7901 (N_7901,N_6350,N_6544);
nand U7902 (N_7902,N_6216,N_6282);
or U7903 (N_7903,N_6249,N_6952);
and U7904 (N_7904,N_6461,N_6161);
nand U7905 (N_7905,N_6568,N_6938);
xor U7906 (N_7906,N_6253,N_6297);
nand U7907 (N_7907,N_6603,N_6987);
nor U7908 (N_7908,N_6140,N_6767);
or U7909 (N_7909,N_6856,N_6543);
and U7910 (N_7910,N_6834,N_6439);
and U7911 (N_7911,N_6812,N_6301);
nand U7912 (N_7912,N_6525,N_6540);
nand U7913 (N_7913,N_6818,N_6369);
nor U7914 (N_7914,N_6124,N_6471);
nand U7915 (N_7915,N_6751,N_6610);
nor U7916 (N_7916,N_6798,N_6452);
and U7917 (N_7917,N_6322,N_6340);
or U7918 (N_7918,N_6573,N_6771);
or U7919 (N_7919,N_6220,N_6150);
and U7920 (N_7920,N_6871,N_6291);
or U7921 (N_7921,N_6553,N_6276);
nand U7922 (N_7922,N_6297,N_6130);
and U7923 (N_7923,N_6144,N_6174);
nor U7924 (N_7924,N_6372,N_6670);
or U7925 (N_7925,N_6665,N_6660);
nand U7926 (N_7926,N_6591,N_6189);
nand U7927 (N_7927,N_6667,N_6599);
nand U7928 (N_7928,N_6576,N_6424);
nand U7929 (N_7929,N_6560,N_6536);
nor U7930 (N_7930,N_6414,N_6307);
or U7931 (N_7931,N_6074,N_6717);
nand U7932 (N_7932,N_6956,N_6539);
nor U7933 (N_7933,N_6816,N_6134);
xnor U7934 (N_7934,N_6764,N_6316);
xor U7935 (N_7935,N_6218,N_6743);
xor U7936 (N_7936,N_6251,N_6258);
nor U7937 (N_7937,N_6259,N_6246);
nand U7938 (N_7938,N_6953,N_6655);
and U7939 (N_7939,N_6453,N_6946);
or U7940 (N_7940,N_6075,N_6716);
nor U7941 (N_7941,N_6980,N_6883);
nor U7942 (N_7942,N_6543,N_6020);
nand U7943 (N_7943,N_6046,N_6158);
nor U7944 (N_7944,N_6874,N_6871);
nor U7945 (N_7945,N_6929,N_6164);
nand U7946 (N_7946,N_6673,N_6353);
nand U7947 (N_7947,N_6380,N_6711);
nand U7948 (N_7948,N_6633,N_6552);
nand U7949 (N_7949,N_6303,N_6388);
nor U7950 (N_7950,N_6681,N_6509);
nand U7951 (N_7951,N_6553,N_6844);
and U7952 (N_7952,N_6005,N_6656);
nand U7953 (N_7953,N_6052,N_6385);
and U7954 (N_7954,N_6942,N_6373);
nand U7955 (N_7955,N_6450,N_6757);
and U7956 (N_7956,N_6845,N_6789);
or U7957 (N_7957,N_6456,N_6418);
nand U7958 (N_7958,N_6918,N_6170);
nand U7959 (N_7959,N_6368,N_6081);
xor U7960 (N_7960,N_6243,N_6184);
and U7961 (N_7961,N_6950,N_6892);
xnor U7962 (N_7962,N_6880,N_6629);
nand U7963 (N_7963,N_6638,N_6073);
xnor U7964 (N_7964,N_6873,N_6280);
xnor U7965 (N_7965,N_6627,N_6314);
nand U7966 (N_7966,N_6456,N_6275);
nor U7967 (N_7967,N_6780,N_6445);
xor U7968 (N_7968,N_6684,N_6900);
nand U7969 (N_7969,N_6504,N_6351);
and U7970 (N_7970,N_6589,N_6618);
nor U7971 (N_7971,N_6106,N_6459);
nand U7972 (N_7972,N_6631,N_6399);
nor U7973 (N_7973,N_6274,N_6053);
nand U7974 (N_7974,N_6263,N_6739);
nor U7975 (N_7975,N_6819,N_6756);
nor U7976 (N_7976,N_6372,N_6932);
and U7977 (N_7977,N_6767,N_6295);
and U7978 (N_7978,N_6108,N_6202);
nor U7979 (N_7979,N_6610,N_6671);
or U7980 (N_7980,N_6093,N_6073);
nor U7981 (N_7981,N_6216,N_6158);
nor U7982 (N_7982,N_6565,N_6632);
nand U7983 (N_7983,N_6835,N_6697);
and U7984 (N_7984,N_6854,N_6714);
and U7985 (N_7985,N_6521,N_6980);
nor U7986 (N_7986,N_6129,N_6980);
nand U7987 (N_7987,N_6188,N_6737);
nand U7988 (N_7988,N_6547,N_6398);
nand U7989 (N_7989,N_6978,N_6623);
nor U7990 (N_7990,N_6716,N_6538);
or U7991 (N_7991,N_6334,N_6527);
nand U7992 (N_7992,N_6793,N_6589);
xor U7993 (N_7993,N_6256,N_6460);
xor U7994 (N_7994,N_6861,N_6887);
and U7995 (N_7995,N_6279,N_6093);
and U7996 (N_7996,N_6573,N_6809);
and U7997 (N_7997,N_6511,N_6974);
nand U7998 (N_7998,N_6622,N_6913);
and U7999 (N_7999,N_6275,N_6514);
or U8000 (N_8000,N_7062,N_7229);
and U8001 (N_8001,N_7988,N_7742);
or U8002 (N_8002,N_7943,N_7236);
and U8003 (N_8003,N_7293,N_7531);
and U8004 (N_8004,N_7775,N_7434);
nor U8005 (N_8005,N_7838,N_7431);
or U8006 (N_8006,N_7342,N_7803);
and U8007 (N_8007,N_7926,N_7797);
or U8008 (N_8008,N_7100,N_7762);
and U8009 (N_8009,N_7520,N_7880);
nor U8010 (N_8010,N_7966,N_7864);
xnor U8011 (N_8011,N_7045,N_7599);
nand U8012 (N_8012,N_7121,N_7693);
nand U8013 (N_8013,N_7020,N_7708);
and U8014 (N_8014,N_7581,N_7899);
nand U8015 (N_8015,N_7211,N_7189);
or U8016 (N_8016,N_7458,N_7980);
nor U8017 (N_8017,N_7035,N_7150);
nand U8018 (N_8018,N_7554,N_7560);
nor U8019 (N_8019,N_7927,N_7230);
nor U8020 (N_8020,N_7848,N_7874);
and U8021 (N_8021,N_7796,N_7265);
or U8022 (N_8022,N_7183,N_7378);
and U8023 (N_8023,N_7091,N_7276);
xor U8024 (N_8024,N_7260,N_7930);
or U8025 (N_8025,N_7303,N_7688);
or U8026 (N_8026,N_7615,N_7248);
or U8027 (N_8027,N_7094,N_7125);
nor U8028 (N_8028,N_7627,N_7791);
nand U8029 (N_8029,N_7534,N_7559);
or U8030 (N_8030,N_7733,N_7630);
or U8031 (N_8031,N_7883,N_7277);
and U8032 (N_8032,N_7590,N_7290);
or U8033 (N_8033,N_7116,N_7916);
and U8034 (N_8034,N_7625,N_7356);
nand U8035 (N_8035,N_7237,N_7405);
or U8036 (N_8036,N_7141,N_7096);
nand U8037 (N_8037,N_7895,N_7146);
and U8038 (N_8038,N_7389,N_7368);
nor U8039 (N_8039,N_7903,N_7370);
nand U8040 (N_8040,N_7021,N_7729);
and U8041 (N_8041,N_7462,N_7649);
or U8042 (N_8042,N_7427,N_7078);
nor U8043 (N_8043,N_7801,N_7437);
or U8044 (N_8044,N_7780,N_7337);
and U8045 (N_8045,N_7993,N_7933);
nor U8046 (N_8046,N_7586,N_7511);
nor U8047 (N_8047,N_7213,N_7812);
xnor U8048 (N_8048,N_7810,N_7242);
and U8049 (N_8049,N_7584,N_7460);
xor U8050 (N_8050,N_7129,N_7232);
and U8051 (N_8051,N_7203,N_7744);
nand U8052 (N_8052,N_7962,N_7798);
nor U8053 (N_8053,N_7524,N_7117);
nand U8054 (N_8054,N_7906,N_7996);
or U8055 (N_8055,N_7030,N_7098);
or U8056 (N_8056,N_7367,N_7765);
or U8057 (N_8057,N_7093,N_7132);
or U8058 (N_8058,N_7081,N_7432);
nand U8059 (N_8059,N_7335,N_7365);
nor U8060 (N_8060,N_7829,N_7738);
or U8061 (N_8061,N_7860,N_7598);
nor U8062 (N_8062,N_7792,N_7366);
or U8063 (N_8063,N_7015,N_7071);
or U8064 (N_8064,N_7907,N_7683);
and U8065 (N_8065,N_7942,N_7173);
or U8066 (N_8066,N_7573,N_7143);
and U8067 (N_8067,N_7244,N_7059);
nand U8068 (N_8068,N_7650,N_7503);
xor U8069 (N_8069,N_7959,N_7270);
nand U8070 (N_8070,N_7299,N_7522);
and U8071 (N_8071,N_7338,N_7710);
and U8072 (N_8072,N_7164,N_7137);
and U8073 (N_8073,N_7602,N_7336);
nor U8074 (N_8074,N_7928,N_7558);
nand U8075 (N_8075,N_7357,N_7379);
nand U8076 (N_8076,N_7392,N_7140);
and U8077 (N_8077,N_7752,N_7169);
or U8078 (N_8078,N_7994,N_7058);
or U8079 (N_8079,N_7414,N_7970);
or U8080 (N_8080,N_7038,N_7313);
and U8081 (N_8081,N_7890,N_7361);
nor U8082 (N_8082,N_7159,N_7477);
or U8083 (N_8083,N_7817,N_7861);
and U8084 (N_8084,N_7888,N_7539);
and U8085 (N_8085,N_7102,N_7662);
or U8086 (N_8086,N_7341,N_7893);
or U8087 (N_8087,N_7429,N_7291);
and U8088 (N_8088,N_7536,N_7799);
nand U8089 (N_8089,N_7023,N_7223);
and U8090 (N_8090,N_7761,N_7428);
and U8091 (N_8091,N_7974,N_7448);
nor U8092 (N_8092,N_7482,N_7605);
or U8093 (N_8093,N_7517,N_7263);
xor U8094 (N_8094,N_7543,N_7334);
nand U8095 (N_8095,N_7013,N_7174);
and U8096 (N_8096,N_7447,N_7523);
nand U8097 (N_8097,N_7629,N_7672);
and U8098 (N_8098,N_7495,N_7734);
nor U8099 (N_8099,N_7452,N_7190);
or U8100 (N_8100,N_7148,N_7922);
nand U8101 (N_8101,N_7162,N_7931);
or U8102 (N_8102,N_7727,N_7051);
nor U8103 (N_8103,N_7939,N_7748);
nand U8104 (N_8104,N_7494,N_7967);
nand U8105 (N_8105,N_7623,N_7288);
or U8106 (N_8106,N_7006,N_7900);
nand U8107 (N_8107,N_7409,N_7467);
nor U8108 (N_8108,N_7202,N_7294);
nor U8109 (N_8109,N_7885,N_7420);
and U8110 (N_8110,N_7069,N_7756);
nand U8111 (N_8111,N_7663,N_7915);
nand U8112 (N_8112,N_7018,N_7725);
nand U8113 (N_8113,N_7846,N_7561);
nor U8114 (N_8114,N_7677,N_7144);
and U8115 (N_8115,N_7610,N_7016);
nor U8116 (N_8116,N_7250,N_7325);
nor U8117 (N_8117,N_7283,N_7564);
and U8118 (N_8118,N_7346,N_7519);
or U8119 (N_8119,N_7323,N_7530);
nand U8120 (N_8120,N_7921,N_7101);
xnor U8121 (N_8121,N_7444,N_7743);
or U8122 (N_8122,N_7876,N_7269);
or U8123 (N_8123,N_7235,N_7377);
nand U8124 (N_8124,N_7925,N_7295);
or U8125 (N_8125,N_7212,N_7318);
and U8126 (N_8126,N_7853,N_7234);
nand U8127 (N_8127,N_7156,N_7579);
xnor U8128 (N_8128,N_7296,N_7594);
and U8129 (N_8129,N_7972,N_7454);
nor U8130 (N_8130,N_7619,N_7858);
and U8131 (N_8131,N_7737,N_7122);
xor U8132 (N_8132,N_7439,N_7596);
and U8133 (N_8133,N_7443,N_7687);
nor U8134 (N_8134,N_7685,N_7867);
nand U8135 (N_8135,N_7066,N_7612);
and U8136 (N_8136,N_7225,N_7360);
nor U8137 (N_8137,N_7655,N_7975);
nand U8138 (N_8138,N_7175,N_7279);
or U8139 (N_8139,N_7292,N_7833);
and U8140 (N_8140,N_7582,N_7772);
nor U8141 (N_8141,N_7553,N_7637);
or U8142 (N_8142,N_7842,N_7750);
nand U8143 (N_8143,N_7606,N_7453);
or U8144 (N_8144,N_7246,N_7375);
or U8145 (N_8145,N_7284,N_7597);
nor U8146 (N_8146,N_7157,N_7938);
or U8147 (N_8147,N_7992,N_7851);
and U8148 (N_8148,N_7466,N_7852);
nand U8149 (N_8149,N_7971,N_7344);
nand U8150 (N_8150,N_7953,N_7546);
nand U8151 (N_8151,N_7345,N_7948);
or U8152 (N_8152,N_7741,N_7954);
xnor U8153 (N_8153,N_7376,N_7919);
and U8154 (N_8154,N_7527,N_7032);
nor U8155 (N_8155,N_7754,N_7542);
and U8156 (N_8156,N_7824,N_7976);
nor U8157 (N_8157,N_7047,N_7347);
and U8158 (N_8158,N_7825,N_7287);
nand U8159 (N_8159,N_7418,N_7407);
nor U8160 (N_8160,N_7875,N_7484);
or U8161 (N_8161,N_7784,N_7968);
nor U8162 (N_8162,N_7210,N_7843);
nand U8163 (N_8163,N_7363,N_7600);
and U8164 (N_8164,N_7831,N_7326);
or U8165 (N_8165,N_7163,N_7856);
nand U8166 (N_8166,N_7340,N_7358);
and U8167 (N_8167,N_7396,N_7349);
xor U8168 (N_8168,N_7089,N_7406);
nor U8169 (N_8169,N_7816,N_7421);
or U8170 (N_8170,N_7312,N_7412);
nor U8171 (N_8171,N_7736,N_7866);
nor U8172 (N_8172,N_7635,N_7771);
xor U8173 (N_8173,N_7509,N_7548);
or U8174 (N_8174,N_7574,N_7311);
and U8175 (N_8175,N_7551,N_7383);
xnor U8176 (N_8176,N_7881,N_7097);
xor U8177 (N_8177,N_7024,N_7304);
and U8178 (N_8178,N_7695,N_7809);
and U8179 (N_8179,N_7485,N_7684);
nor U8180 (N_8180,N_7869,N_7104);
and U8181 (N_8181,N_7892,N_7656);
or U8182 (N_8182,N_7835,N_7155);
nor U8183 (N_8183,N_7702,N_7721);
nand U8184 (N_8184,N_7221,N_7497);
nand U8185 (N_8185,N_7747,N_7187);
and U8186 (N_8186,N_7981,N_7528);
or U8187 (N_8187,N_7192,N_7195);
nand U8188 (N_8188,N_7067,N_7647);
and U8189 (N_8189,N_7233,N_7332);
nor U8190 (N_8190,N_7158,N_7348);
or U8191 (N_8191,N_7438,N_7001);
or U8192 (N_8192,N_7130,N_7779);
nand U8193 (N_8193,N_7254,N_7219);
nand U8194 (N_8194,N_7675,N_7673);
or U8195 (N_8195,N_7639,N_7425);
or U8196 (N_8196,N_7424,N_7740);
xnor U8197 (N_8197,N_7070,N_7354);
and U8198 (N_8198,N_7877,N_7128);
nor U8199 (N_8199,N_7956,N_7372);
nor U8200 (N_8200,N_7778,N_7442);
nor U8201 (N_8201,N_7142,N_7570);
nor U8202 (N_8202,N_7714,N_7136);
xnor U8203 (N_8203,N_7651,N_7138);
and U8204 (N_8204,N_7124,N_7944);
and U8205 (N_8205,N_7243,N_7355);
or U8206 (N_8206,N_7196,N_7904);
nand U8207 (N_8207,N_7696,N_7440);
nand U8208 (N_8208,N_7267,N_7398);
and U8209 (N_8209,N_7513,N_7153);
and U8210 (N_8210,N_7215,N_7955);
or U8211 (N_8211,N_7674,N_7588);
nor U8212 (N_8212,N_7819,N_7682);
and U8213 (N_8213,N_7764,N_7510);
nand U8214 (N_8214,N_7505,N_7571);
xnor U8215 (N_8215,N_7583,N_7618);
nor U8216 (N_8216,N_7218,N_7172);
xor U8217 (N_8217,N_7364,N_7697);
nor U8218 (N_8218,N_7133,N_7611);
nand U8219 (N_8219,N_7808,N_7302);
and U8220 (N_8220,N_7847,N_7704);
nand U8221 (N_8221,N_7728,N_7834);
nor U8222 (N_8222,N_7010,N_7671);
nand U8223 (N_8223,N_7855,N_7565);
or U8224 (N_8224,N_7533,N_7952);
and U8225 (N_8225,N_7821,N_7214);
nand U8226 (N_8226,N_7152,N_7592);
nor U8227 (N_8227,N_7836,N_7964);
xor U8228 (N_8228,N_7065,N_7206);
nor U8229 (N_8229,N_7430,N_7076);
nand U8230 (N_8230,N_7415,N_7545);
nor U8231 (N_8231,N_7788,N_7508);
or U8232 (N_8232,N_7487,N_7620);
and U8233 (N_8233,N_7423,N_7562);
nor U8234 (N_8234,N_7550,N_7908);
and U8235 (N_8235,N_7924,N_7755);
or U8236 (N_8236,N_7987,N_7151);
or U8237 (N_8237,N_7465,N_7666);
and U8238 (N_8238,N_7207,N_7608);
nor U8239 (N_8239,N_7205,N_7170);
or U8240 (N_8240,N_7028,N_7055);
nor U8241 (N_8241,N_7009,N_7521);
nand U8242 (N_8242,N_7087,N_7555);
and U8243 (N_8243,N_7476,N_7947);
xnor U8244 (N_8244,N_7567,N_7787);
and U8245 (N_8245,N_7631,N_7227);
or U8246 (N_8246,N_7113,N_7770);
and U8247 (N_8247,N_7258,N_7217);
nand U8248 (N_8248,N_7636,N_7918);
nand U8249 (N_8249,N_7641,N_7958);
nor U8250 (N_8250,N_7879,N_7445);
nor U8251 (N_8251,N_7910,N_7168);
or U8252 (N_8252,N_7665,N_7413);
or U8253 (N_8253,N_7251,N_7488);
nand U8254 (N_8254,N_7621,N_7397);
and U8255 (N_8255,N_7123,N_7374);
or U8256 (N_8256,N_7676,N_7607);
or U8257 (N_8257,N_7231,N_7540);
and U8258 (N_8258,N_7359,N_7802);
and U8259 (N_8259,N_7969,N_7126);
and U8260 (N_8260,N_7498,N_7758);
xor U8261 (N_8261,N_7095,N_7046);
or U8262 (N_8262,N_7241,N_7837);
and U8263 (N_8263,N_7297,N_7468);
nand U8264 (N_8264,N_7135,N_7282);
and U8265 (N_8265,N_7257,N_7049);
nand U8266 (N_8266,N_7316,N_7456);
nor U8267 (N_8267,N_7811,N_7481);
or U8268 (N_8268,N_7896,N_7701);
or U8269 (N_8269,N_7331,N_7723);
xnor U8270 (N_8270,N_7614,N_7891);
and U8271 (N_8271,N_7735,N_7262);
and U8272 (N_8272,N_7199,N_7746);
nand U8273 (N_8273,N_7705,N_7934);
or U8274 (N_8274,N_7694,N_7785);
nand U8275 (N_8275,N_7563,N_7616);
and U8276 (N_8276,N_7617,N_7624);
and U8277 (N_8277,N_7362,N_7381);
nand U8278 (N_8278,N_7111,N_7857);
nor U8279 (N_8279,N_7960,N_7391);
or U8280 (N_8280,N_7670,N_7781);
nand U8281 (N_8281,N_7459,N_7228);
xnor U8282 (N_8282,N_7327,N_7790);
nor U8283 (N_8283,N_7706,N_7403);
nand U8284 (N_8284,N_7859,N_7986);
and U8285 (N_8285,N_7208,N_7769);
or U8286 (N_8286,N_7216,N_7587);
or U8287 (N_8287,N_7713,N_7854);
nor U8288 (N_8288,N_7092,N_7632);
and U8289 (N_8289,N_7793,N_7305);
nor U8290 (N_8290,N_7469,N_7898);
nand U8291 (N_8291,N_7449,N_7913);
nand U8292 (N_8292,N_7593,N_7106);
nand U8293 (N_8293,N_7000,N_7640);
and U8294 (N_8294,N_7180,N_7507);
nor U8295 (N_8295,N_7491,N_7518);
nand U8296 (N_8296,N_7814,N_7917);
xor U8297 (N_8297,N_7450,N_7300);
and U8298 (N_8298,N_7201,N_7086);
or U8299 (N_8299,N_7572,N_7777);
or U8300 (N_8300,N_7176,N_7063);
and U8301 (N_8301,N_7978,N_7805);
nor U8302 (N_8302,N_7185,N_7451);
xor U8303 (N_8303,N_7249,N_7794);
nand U8304 (N_8304,N_7060,N_7002);
nor U8305 (N_8305,N_7646,N_7399);
and U8306 (N_8306,N_7820,N_7390);
or U8307 (N_8307,N_7134,N_7274);
nor U8308 (N_8308,N_7184,N_7167);
nor U8309 (N_8309,N_7845,N_7373);
nor U8310 (N_8310,N_7400,N_7654);
and U8311 (N_8311,N_7680,N_7753);
nor U8312 (N_8312,N_7731,N_7935);
xor U8313 (N_8313,N_7514,N_7998);
nand U8314 (N_8314,N_7333,N_7471);
nor U8315 (N_8315,N_7800,N_7658);
nand U8316 (N_8316,N_7818,N_7884);
nand U8317 (N_8317,N_7751,N_7268);
or U8318 (N_8318,N_7490,N_7863);
or U8319 (N_8319,N_7317,N_7679);
xnor U8320 (N_8320,N_7011,N_7648);
or U8321 (N_8321,N_7749,N_7064);
nor U8322 (N_8322,N_7017,N_7999);
nand U8323 (N_8323,N_7862,N_7120);
and U8324 (N_8324,N_7669,N_7384);
and U8325 (N_8325,N_7711,N_7394);
and U8326 (N_8326,N_7003,N_7989);
nor U8327 (N_8327,N_7541,N_7515);
and U8328 (N_8328,N_7763,N_7052);
nor U8329 (N_8329,N_7131,N_7516);
nand U8330 (N_8330,N_7827,N_7767);
nand U8331 (N_8331,N_7961,N_7147);
and U8332 (N_8332,N_7027,N_7273);
nor U8333 (N_8333,N_7386,N_7480);
or U8334 (N_8334,N_7692,N_7191);
and U8335 (N_8335,N_7473,N_7871);
xor U8336 (N_8336,N_7774,N_7983);
or U8337 (N_8337,N_7209,N_7526);
xor U8338 (N_8338,N_7114,N_7048);
nor U8339 (N_8339,N_7689,N_7882);
and U8340 (N_8340,N_7105,N_7188);
or U8341 (N_8341,N_7865,N_7436);
nor U8342 (N_8342,N_7990,N_7224);
nand U8343 (N_8343,N_7039,N_7298);
nor U8344 (N_8344,N_7040,N_7849);
nor U8345 (N_8345,N_7160,N_7929);
and U8346 (N_8346,N_7609,N_7760);
and U8347 (N_8347,N_7309,N_7280);
or U8348 (N_8348,N_7461,N_7850);
nand U8349 (N_8349,N_7029,N_7878);
nor U8350 (N_8350,N_7433,N_7252);
and U8351 (N_8351,N_7700,N_7826);
nor U8352 (N_8352,N_7773,N_7946);
xnor U8353 (N_8353,N_7053,N_7417);
and U8354 (N_8354,N_7319,N_7603);
and U8355 (N_8355,N_7901,N_7532);
and U8356 (N_8356,N_7073,N_7902);
and U8357 (N_8357,N_7984,N_7455);
and U8358 (N_8358,N_7912,N_7678);
nor U8359 (N_8359,N_7239,N_7538);
nand U8360 (N_8360,N_7278,N_7082);
and U8361 (N_8361,N_7652,N_7084);
or U8362 (N_8362,N_7139,N_7289);
nor U8363 (N_8363,N_7044,N_7350);
nand U8364 (N_8364,N_7719,N_7932);
and U8365 (N_8365,N_7645,N_7965);
xnor U8366 (N_8366,N_7807,N_7822);
nor U8367 (N_8367,N_7256,N_7036);
or U8368 (N_8368,N_7535,N_7795);
nor U8369 (N_8369,N_7037,N_7281);
nand U8370 (N_8370,N_7077,N_7310);
xor U8371 (N_8371,N_7568,N_7977);
or U8372 (N_8372,N_7475,N_7005);
and U8373 (N_8373,N_7200,N_7261);
nor U8374 (N_8374,N_7759,N_7591);
nand U8375 (N_8375,N_7569,N_7470);
or U8376 (N_8376,N_7985,N_7557);
or U8377 (N_8377,N_7887,N_7642);
and U8378 (N_8378,N_7745,N_7698);
nor U8379 (N_8379,N_7489,N_7395);
and U8380 (N_8380,N_7501,N_7782);
xor U8381 (N_8381,N_7840,N_7198);
and U8382 (N_8382,N_7668,N_7393);
nand U8383 (N_8383,N_7112,N_7628);
and U8384 (N_8384,N_7492,N_7329);
nor U8385 (N_8385,N_7074,N_7506);
nand U8386 (N_8386,N_7963,N_7633);
nor U8387 (N_8387,N_7496,N_7410);
xor U8388 (N_8388,N_7979,N_7720);
nor U8389 (N_8389,N_7245,N_7766);
and U8390 (N_8390,N_7786,N_7712);
nand U8391 (N_8391,N_7686,N_7008);
nor U8392 (N_8392,N_7718,N_7474);
or U8393 (N_8393,N_7991,N_7870);
or U8394 (N_8394,N_7401,N_7054);
nor U8395 (N_8395,N_7108,N_7982);
or U8396 (N_8396,N_7957,N_7352);
and U8397 (N_8397,N_7119,N_7285);
or U8398 (N_8398,N_7703,N_7149);
or U8399 (N_8399,N_7315,N_7330);
nor U8400 (N_8400,N_7457,N_7806);
nand U8401 (N_8401,N_7079,N_7830);
and U8402 (N_8402,N_7380,N_7578);
nand U8403 (N_8403,N_7691,N_7525);
nor U8404 (N_8404,N_7499,N_7324);
or U8405 (N_8405,N_7643,N_7951);
or U8406 (N_8406,N_7446,N_7783);
nor U8407 (N_8407,N_7657,N_7041);
nand U8408 (N_8408,N_7815,N_7544);
nor U8409 (N_8409,N_7844,N_7699);
or U8410 (N_8410,N_7661,N_7080);
and U8411 (N_8411,N_7547,N_7240);
nand U8412 (N_8412,N_7050,N_7973);
nand U8413 (N_8413,N_7644,N_7681);
xnor U8414 (N_8414,N_7388,N_7115);
nor U8415 (N_8415,N_7014,N_7667);
and U8416 (N_8416,N_7385,N_7099);
nor U8417 (N_8417,N_7118,N_7945);
nor U8418 (N_8418,N_7556,N_7033);
nor U8419 (N_8419,N_7272,N_7264);
nor U8420 (N_8420,N_7589,N_7823);
nor U8421 (N_8421,N_7813,N_7909);
nand U8422 (N_8422,N_7937,N_7369);
nor U8423 (N_8423,N_7911,N_7690);
nand U8424 (N_8424,N_7613,N_7601);
or U8425 (N_8425,N_7472,N_7905);
nand U8426 (N_8426,N_7306,N_7997);
nand U8427 (N_8427,N_7411,N_7920);
and U8428 (N_8428,N_7075,N_7634);
nor U8429 (N_8429,N_7730,N_7301);
nand U8430 (N_8430,N_7638,N_7253);
xnor U8431 (N_8431,N_7321,N_7441);
xnor U8432 (N_8432,N_7426,N_7416);
and U8433 (N_8433,N_7716,N_7186);
and U8434 (N_8434,N_7259,N_7757);
nor U8435 (N_8435,N_7166,N_7178);
and U8436 (N_8436,N_7022,N_7575);
and U8437 (N_8437,N_7950,N_7504);
nand U8438 (N_8438,N_7088,N_7220);
and U8439 (N_8439,N_7328,N_7664);
nand U8440 (N_8440,N_7387,N_7182);
or U8441 (N_8441,N_7371,N_7042);
nand U8442 (N_8442,N_7083,N_7537);
or U8443 (N_8443,N_7109,N_7732);
nand U8444 (N_8444,N_7886,N_7314);
xor U8445 (N_8445,N_7897,N_7804);
nand U8446 (N_8446,N_7715,N_7726);
or U8447 (N_8447,N_7353,N_7320);
and U8448 (N_8448,N_7841,N_7653);
nand U8449 (N_8449,N_7419,N_7549);
or U8450 (N_8450,N_7404,N_7483);
nand U8451 (N_8451,N_7512,N_7709);
nand U8452 (N_8452,N_7193,N_7154);
nand U8453 (N_8453,N_7308,N_7408);
or U8454 (N_8454,N_7255,N_7402);
nand U8455 (N_8455,N_7351,N_7161);
or U8456 (N_8456,N_7832,N_7343);
nand U8457 (N_8457,N_7464,N_7026);
nand U8458 (N_8458,N_7145,N_7577);
nand U8459 (N_8459,N_7872,N_7940);
or U8460 (N_8460,N_7322,N_7072);
nand U8461 (N_8461,N_7576,N_7103);
or U8462 (N_8462,N_7204,N_7339);
xnor U8463 (N_8463,N_7768,N_7286);
xor U8464 (N_8464,N_7271,N_7085);
nand U8465 (N_8465,N_7622,N_7995);
xor U8466 (N_8466,N_7238,N_7660);
and U8467 (N_8467,N_7435,N_7941);
or U8468 (N_8468,N_7659,N_7585);
nor U8469 (N_8469,N_7061,N_7478);
or U8470 (N_8470,N_7486,N_7717);
nand U8471 (N_8471,N_7595,N_7266);
nor U8472 (N_8472,N_7056,N_7107);
and U8473 (N_8473,N_7171,N_7034);
xnor U8474 (N_8474,N_7194,N_7177);
or U8475 (N_8475,N_7894,N_7868);
and U8476 (N_8476,N_7165,N_7604);
or U8477 (N_8477,N_7626,N_7566);
xor U8478 (N_8478,N_7090,N_7043);
nand U8479 (N_8479,N_7019,N_7479);
and U8480 (N_8480,N_7226,N_7382);
nor U8481 (N_8481,N_7181,N_7949);
nor U8482 (N_8482,N_7722,N_7004);
nor U8483 (N_8483,N_7529,N_7789);
or U8484 (N_8484,N_7936,N_7422);
nand U8485 (N_8485,N_7463,N_7500);
nand U8486 (N_8486,N_7197,N_7776);
or U8487 (N_8487,N_7307,N_7031);
or U8488 (N_8488,N_7914,N_7828);
nor U8489 (N_8489,N_7110,N_7068);
or U8490 (N_8490,N_7057,N_7873);
and U8491 (N_8491,N_7724,N_7502);
or U8492 (N_8492,N_7179,N_7580);
or U8493 (N_8493,N_7247,N_7923);
or U8494 (N_8494,N_7222,N_7839);
nor U8495 (N_8495,N_7012,N_7493);
or U8496 (N_8496,N_7025,N_7707);
nand U8497 (N_8497,N_7739,N_7127);
and U8498 (N_8498,N_7889,N_7552);
and U8499 (N_8499,N_7007,N_7275);
nor U8500 (N_8500,N_7707,N_7329);
nor U8501 (N_8501,N_7793,N_7285);
or U8502 (N_8502,N_7458,N_7757);
and U8503 (N_8503,N_7269,N_7026);
and U8504 (N_8504,N_7101,N_7022);
and U8505 (N_8505,N_7217,N_7656);
or U8506 (N_8506,N_7285,N_7947);
nor U8507 (N_8507,N_7929,N_7832);
nand U8508 (N_8508,N_7113,N_7562);
and U8509 (N_8509,N_7092,N_7309);
and U8510 (N_8510,N_7192,N_7856);
or U8511 (N_8511,N_7141,N_7812);
nor U8512 (N_8512,N_7246,N_7870);
nand U8513 (N_8513,N_7983,N_7517);
and U8514 (N_8514,N_7692,N_7687);
xnor U8515 (N_8515,N_7512,N_7048);
nand U8516 (N_8516,N_7516,N_7594);
nand U8517 (N_8517,N_7965,N_7292);
nor U8518 (N_8518,N_7575,N_7534);
nand U8519 (N_8519,N_7045,N_7476);
nor U8520 (N_8520,N_7661,N_7040);
or U8521 (N_8521,N_7802,N_7653);
or U8522 (N_8522,N_7795,N_7599);
nor U8523 (N_8523,N_7061,N_7111);
nor U8524 (N_8524,N_7243,N_7548);
and U8525 (N_8525,N_7731,N_7184);
or U8526 (N_8526,N_7779,N_7104);
nand U8527 (N_8527,N_7824,N_7360);
nand U8528 (N_8528,N_7231,N_7565);
nand U8529 (N_8529,N_7941,N_7841);
nand U8530 (N_8530,N_7033,N_7655);
nor U8531 (N_8531,N_7093,N_7431);
and U8532 (N_8532,N_7053,N_7549);
or U8533 (N_8533,N_7286,N_7436);
nand U8534 (N_8534,N_7979,N_7537);
and U8535 (N_8535,N_7147,N_7470);
or U8536 (N_8536,N_7133,N_7945);
or U8537 (N_8537,N_7052,N_7254);
and U8538 (N_8538,N_7828,N_7768);
and U8539 (N_8539,N_7498,N_7336);
xnor U8540 (N_8540,N_7145,N_7547);
and U8541 (N_8541,N_7303,N_7901);
xor U8542 (N_8542,N_7803,N_7439);
and U8543 (N_8543,N_7783,N_7616);
and U8544 (N_8544,N_7775,N_7193);
and U8545 (N_8545,N_7258,N_7665);
nor U8546 (N_8546,N_7800,N_7157);
and U8547 (N_8547,N_7583,N_7117);
nand U8548 (N_8548,N_7418,N_7447);
nor U8549 (N_8549,N_7321,N_7106);
and U8550 (N_8550,N_7978,N_7603);
xnor U8551 (N_8551,N_7780,N_7003);
or U8552 (N_8552,N_7273,N_7825);
xor U8553 (N_8553,N_7321,N_7961);
or U8554 (N_8554,N_7034,N_7836);
nor U8555 (N_8555,N_7303,N_7804);
or U8556 (N_8556,N_7503,N_7223);
or U8557 (N_8557,N_7159,N_7348);
or U8558 (N_8558,N_7363,N_7462);
and U8559 (N_8559,N_7216,N_7381);
or U8560 (N_8560,N_7650,N_7851);
and U8561 (N_8561,N_7509,N_7062);
or U8562 (N_8562,N_7873,N_7026);
nor U8563 (N_8563,N_7696,N_7846);
nor U8564 (N_8564,N_7167,N_7929);
xnor U8565 (N_8565,N_7907,N_7049);
nand U8566 (N_8566,N_7459,N_7486);
nand U8567 (N_8567,N_7480,N_7740);
and U8568 (N_8568,N_7938,N_7426);
nand U8569 (N_8569,N_7585,N_7353);
or U8570 (N_8570,N_7871,N_7600);
nand U8571 (N_8571,N_7579,N_7683);
nor U8572 (N_8572,N_7910,N_7490);
nand U8573 (N_8573,N_7177,N_7800);
nand U8574 (N_8574,N_7258,N_7925);
or U8575 (N_8575,N_7011,N_7724);
nand U8576 (N_8576,N_7494,N_7009);
nand U8577 (N_8577,N_7760,N_7347);
or U8578 (N_8578,N_7770,N_7042);
or U8579 (N_8579,N_7065,N_7482);
nor U8580 (N_8580,N_7816,N_7937);
nor U8581 (N_8581,N_7333,N_7447);
nand U8582 (N_8582,N_7777,N_7617);
nand U8583 (N_8583,N_7982,N_7691);
or U8584 (N_8584,N_7949,N_7751);
xnor U8585 (N_8585,N_7833,N_7271);
nor U8586 (N_8586,N_7118,N_7327);
xor U8587 (N_8587,N_7653,N_7480);
or U8588 (N_8588,N_7570,N_7654);
nand U8589 (N_8589,N_7578,N_7911);
or U8590 (N_8590,N_7612,N_7556);
or U8591 (N_8591,N_7485,N_7237);
or U8592 (N_8592,N_7319,N_7477);
nor U8593 (N_8593,N_7884,N_7874);
nand U8594 (N_8594,N_7265,N_7530);
or U8595 (N_8595,N_7957,N_7308);
nor U8596 (N_8596,N_7930,N_7006);
nor U8597 (N_8597,N_7108,N_7472);
and U8598 (N_8598,N_7694,N_7075);
and U8599 (N_8599,N_7977,N_7565);
nor U8600 (N_8600,N_7551,N_7629);
xor U8601 (N_8601,N_7980,N_7940);
and U8602 (N_8602,N_7423,N_7249);
or U8603 (N_8603,N_7318,N_7457);
or U8604 (N_8604,N_7101,N_7526);
nand U8605 (N_8605,N_7447,N_7069);
or U8606 (N_8606,N_7242,N_7820);
nor U8607 (N_8607,N_7884,N_7859);
or U8608 (N_8608,N_7467,N_7839);
nor U8609 (N_8609,N_7393,N_7321);
nor U8610 (N_8610,N_7597,N_7368);
or U8611 (N_8611,N_7419,N_7139);
and U8612 (N_8612,N_7839,N_7646);
nand U8613 (N_8613,N_7347,N_7030);
or U8614 (N_8614,N_7112,N_7370);
or U8615 (N_8615,N_7124,N_7743);
xnor U8616 (N_8616,N_7887,N_7622);
nor U8617 (N_8617,N_7852,N_7455);
and U8618 (N_8618,N_7850,N_7244);
xnor U8619 (N_8619,N_7525,N_7766);
or U8620 (N_8620,N_7283,N_7076);
nand U8621 (N_8621,N_7775,N_7813);
nand U8622 (N_8622,N_7501,N_7319);
nor U8623 (N_8623,N_7686,N_7617);
nand U8624 (N_8624,N_7809,N_7637);
and U8625 (N_8625,N_7827,N_7137);
and U8626 (N_8626,N_7792,N_7550);
or U8627 (N_8627,N_7612,N_7310);
nor U8628 (N_8628,N_7565,N_7409);
nor U8629 (N_8629,N_7563,N_7299);
nor U8630 (N_8630,N_7218,N_7888);
or U8631 (N_8631,N_7285,N_7496);
or U8632 (N_8632,N_7894,N_7316);
or U8633 (N_8633,N_7880,N_7555);
and U8634 (N_8634,N_7311,N_7224);
nand U8635 (N_8635,N_7655,N_7325);
and U8636 (N_8636,N_7514,N_7910);
nand U8637 (N_8637,N_7986,N_7170);
nor U8638 (N_8638,N_7022,N_7231);
nand U8639 (N_8639,N_7315,N_7055);
xor U8640 (N_8640,N_7785,N_7000);
nor U8641 (N_8641,N_7242,N_7978);
or U8642 (N_8642,N_7439,N_7442);
nor U8643 (N_8643,N_7147,N_7723);
nand U8644 (N_8644,N_7799,N_7592);
nand U8645 (N_8645,N_7080,N_7836);
nor U8646 (N_8646,N_7236,N_7982);
nor U8647 (N_8647,N_7217,N_7136);
and U8648 (N_8648,N_7262,N_7988);
nand U8649 (N_8649,N_7807,N_7213);
nand U8650 (N_8650,N_7967,N_7878);
or U8651 (N_8651,N_7213,N_7051);
nor U8652 (N_8652,N_7865,N_7052);
or U8653 (N_8653,N_7091,N_7269);
nand U8654 (N_8654,N_7445,N_7912);
xor U8655 (N_8655,N_7756,N_7074);
nor U8656 (N_8656,N_7742,N_7475);
and U8657 (N_8657,N_7155,N_7948);
xnor U8658 (N_8658,N_7137,N_7820);
or U8659 (N_8659,N_7767,N_7530);
xnor U8660 (N_8660,N_7654,N_7600);
and U8661 (N_8661,N_7921,N_7419);
xor U8662 (N_8662,N_7023,N_7187);
xor U8663 (N_8663,N_7076,N_7279);
nand U8664 (N_8664,N_7969,N_7813);
and U8665 (N_8665,N_7459,N_7774);
and U8666 (N_8666,N_7599,N_7756);
or U8667 (N_8667,N_7569,N_7477);
and U8668 (N_8668,N_7228,N_7596);
or U8669 (N_8669,N_7055,N_7699);
or U8670 (N_8670,N_7606,N_7467);
or U8671 (N_8671,N_7701,N_7219);
or U8672 (N_8672,N_7719,N_7507);
nor U8673 (N_8673,N_7496,N_7955);
or U8674 (N_8674,N_7806,N_7227);
or U8675 (N_8675,N_7344,N_7256);
or U8676 (N_8676,N_7127,N_7874);
nor U8677 (N_8677,N_7598,N_7139);
and U8678 (N_8678,N_7130,N_7066);
nor U8679 (N_8679,N_7323,N_7809);
and U8680 (N_8680,N_7510,N_7739);
nand U8681 (N_8681,N_7355,N_7552);
and U8682 (N_8682,N_7497,N_7254);
nand U8683 (N_8683,N_7582,N_7909);
nor U8684 (N_8684,N_7279,N_7150);
and U8685 (N_8685,N_7966,N_7939);
and U8686 (N_8686,N_7011,N_7463);
nor U8687 (N_8687,N_7781,N_7499);
nor U8688 (N_8688,N_7141,N_7625);
or U8689 (N_8689,N_7845,N_7476);
or U8690 (N_8690,N_7936,N_7592);
xor U8691 (N_8691,N_7962,N_7617);
or U8692 (N_8692,N_7633,N_7704);
and U8693 (N_8693,N_7512,N_7871);
nand U8694 (N_8694,N_7460,N_7657);
nand U8695 (N_8695,N_7738,N_7662);
or U8696 (N_8696,N_7850,N_7969);
or U8697 (N_8697,N_7847,N_7376);
nand U8698 (N_8698,N_7026,N_7263);
nor U8699 (N_8699,N_7020,N_7036);
or U8700 (N_8700,N_7929,N_7881);
and U8701 (N_8701,N_7248,N_7813);
nand U8702 (N_8702,N_7154,N_7511);
xor U8703 (N_8703,N_7375,N_7182);
nand U8704 (N_8704,N_7381,N_7357);
nor U8705 (N_8705,N_7326,N_7997);
or U8706 (N_8706,N_7188,N_7472);
nand U8707 (N_8707,N_7061,N_7543);
and U8708 (N_8708,N_7119,N_7175);
and U8709 (N_8709,N_7828,N_7766);
and U8710 (N_8710,N_7685,N_7491);
xnor U8711 (N_8711,N_7030,N_7768);
nand U8712 (N_8712,N_7069,N_7220);
xor U8713 (N_8713,N_7178,N_7933);
xor U8714 (N_8714,N_7997,N_7371);
and U8715 (N_8715,N_7790,N_7221);
nand U8716 (N_8716,N_7430,N_7132);
or U8717 (N_8717,N_7730,N_7467);
nor U8718 (N_8718,N_7326,N_7027);
nand U8719 (N_8719,N_7394,N_7110);
and U8720 (N_8720,N_7743,N_7140);
and U8721 (N_8721,N_7089,N_7662);
or U8722 (N_8722,N_7337,N_7032);
nor U8723 (N_8723,N_7398,N_7252);
or U8724 (N_8724,N_7789,N_7871);
or U8725 (N_8725,N_7278,N_7200);
and U8726 (N_8726,N_7494,N_7163);
or U8727 (N_8727,N_7511,N_7343);
xnor U8728 (N_8728,N_7937,N_7015);
nor U8729 (N_8729,N_7655,N_7473);
or U8730 (N_8730,N_7841,N_7673);
and U8731 (N_8731,N_7142,N_7386);
and U8732 (N_8732,N_7365,N_7701);
nand U8733 (N_8733,N_7294,N_7667);
nand U8734 (N_8734,N_7302,N_7284);
nor U8735 (N_8735,N_7323,N_7798);
or U8736 (N_8736,N_7488,N_7988);
xor U8737 (N_8737,N_7475,N_7073);
nor U8738 (N_8738,N_7334,N_7660);
and U8739 (N_8739,N_7124,N_7487);
nand U8740 (N_8740,N_7640,N_7016);
nand U8741 (N_8741,N_7361,N_7158);
or U8742 (N_8742,N_7067,N_7028);
nand U8743 (N_8743,N_7646,N_7644);
nand U8744 (N_8744,N_7922,N_7509);
and U8745 (N_8745,N_7932,N_7226);
nor U8746 (N_8746,N_7894,N_7297);
or U8747 (N_8747,N_7867,N_7526);
nor U8748 (N_8748,N_7782,N_7647);
xor U8749 (N_8749,N_7421,N_7656);
and U8750 (N_8750,N_7475,N_7535);
or U8751 (N_8751,N_7947,N_7430);
nand U8752 (N_8752,N_7766,N_7936);
or U8753 (N_8753,N_7640,N_7326);
nand U8754 (N_8754,N_7700,N_7283);
and U8755 (N_8755,N_7757,N_7207);
or U8756 (N_8756,N_7149,N_7034);
xnor U8757 (N_8757,N_7462,N_7451);
and U8758 (N_8758,N_7345,N_7159);
nor U8759 (N_8759,N_7078,N_7895);
nor U8760 (N_8760,N_7334,N_7568);
nand U8761 (N_8761,N_7206,N_7594);
or U8762 (N_8762,N_7498,N_7593);
or U8763 (N_8763,N_7051,N_7083);
nand U8764 (N_8764,N_7374,N_7172);
nor U8765 (N_8765,N_7623,N_7313);
or U8766 (N_8766,N_7258,N_7411);
and U8767 (N_8767,N_7381,N_7268);
or U8768 (N_8768,N_7928,N_7989);
nand U8769 (N_8769,N_7607,N_7415);
or U8770 (N_8770,N_7437,N_7278);
nor U8771 (N_8771,N_7094,N_7242);
nand U8772 (N_8772,N_7385,N_7491);
and U8773 (N_8773,N_7626,N_7438);
and U8774 (N_8774,N_7362,N_7531);
or U8775 (N_8775,N_7222,N_7278);
and U8776 (N_8776,N_7230,N_7675);
and U8777 (N_8777,N_7637,N_7451);
and U8778 (N_8778,N_7554,N_7940);
and U8779 (N_8779,N_7332,N_7140);
nor U8780 (N_8780,N_7116,N_7104);
nand U8781 (N_8781,N_7185,N_7748);
xnor U8782 (N_8782,N_7376,N_7590);
or U8783 (N_8783,N_7739,N_7808);
nand U8784 (N_8784,N_7336,N_7616);
nor U8785 (N_8785,N_7140,N_7982);
xnor U8786 (N_8786,N_7009,N_7233);
nor U8787 (N_8787,N_7564,N_7230);
or U8788 (N_8788,N_7174,N_7289);
xnor U8789 (N_8789,N_7622,N_7708);
or U8790 (N_8790,N_7073,N_7361);
or U8791 (N_8791,N_7357,N_7286);
nand U8792 (N_8792,N_7858,N_7526);
nand U8793 (N_8793,N_7030,N_7375);
nand U8794 (N_8794,N_7119,N_7813);
nand U8795 (N_8795,N_7168,N_7749);
xnor U8796 (N_8796,N_7357,N_7401);
or U8797 (N_8797,N_7113,N_7876);
or U8798 (N_8798,N_7324,N_7621);
nand U8799 (N_8799,N_7435,N_7049);
or U8800 (N_8800,N_7156,N_7961);
nand U8801 (N_8801,N_7459,N_7143);
nand U8802 (N_8802,N_7930,N_7141);
nor U8803 (N_8803,N_7583,N_7250);
nand U8804 (N_8804,N_7600,N_7170);
and U8805 (N_8805,N_7810,N_7910);
xor U8806 (N_8806,N_7630,N_7656);
nand U8807 (N_8807,N_7556,N_7713);
nor U8808 (N_8808,N_7328,N_7599);
or U8809 (N_8809,N_7596,N_7347);
and U8810 (N_8810,N_7270,N_7100);
or U8811 (N_8811,N_7794,N_7371);
nor U8812 (N_8812,N_7157,N_7009);
nor U8813 (N_8813,N_7859,N_7702);
or U8814 (N_8814,N_7590,N_7243);
nand U8815 (N_8815,N_7759,N_7560);
xnor U8816 (N_8816,N_7648,N_7396);
xnor U8817 (N_8817,N_7052,N_7168);
or U8818 (N_8818,N_7793,N_7487);
and U8819 (N_8819,N_7783,N_7078);
and U8820 (N_8820,N_7789,N_7539);
and U8821 (N_8821,N_7768,N_7492);
and U8822 (N_8822,N_7193,N_7992);
nand U8823 (N_8823,N_7341,N_7827);
or U8824 (N_8824,N_7271,N_7783);
nor U8825 (N_8825,N_7132,N_7760);
xnor U8826 (N_8826,N_7243,N_7539);
nand U8827 (N_8827,N_7638,N_7939);
xor U8828 (N_8828,N_7347,N_7009);
or U8829 (N_8829,N_7352,N_7054);
nand U8830 (N_8830,N_7360,N_7369);
nor U8831 (N_8831,N_7652,N_7660);
nor U8832 (N_8832,N_7153,N_7610);
nor U8833 (N_8833,N_7669,N_7166);
and U8834 (N_8834,N_7069,N_7108);
and U8835 (N_8835,N_7123,N_7654);
and U8836 (N_8836,N_7300,N_7830);
nor U8837 (N_8837,N_7759,N_7284);
or U8838 (N_8838,N_7346,N_7150);
or U8839 (N_8839,N_7145,N_7350);
or U8840 (N_8840,N_7163,N_7194);
nand U8841 (N_8841,N_7612,N_7880);
nand U8842 (N_8842,N_7932,N_7691);
or U8843 (N_8843,N_7669,N_7057);
and U8844 (N_8844,N_7554,N_7097);
nand U8845 (N_8845,N_7491,N_7678);
nor U8846 (N_8846,N_7392,N_7630);
nor U8847 (N_8847,N_7999,N_7458);
nor U8848 (N_8848,N_7716,N_7357);
nand U8849 (N_8849,N_7046,N_7491);
and U8850 (N_8850,N_7563,N_7515);
nand U8851 (N_8851,N_7777,N_7053);
nor U8852 (N_8852,N_7246,N_7597);
nand U8853 (N_8853,N_7450,N_7896);
and U8854 (N_8854,N_7531,N_7084);
or U8855 (N_8855,N_7828,N_7888);
nand U8856 (N_8856,N_7130,N_7961);
nor U8857 (N_8857,N_7260,N_7475);
nand U8858 (N_8858,N_7859,N_7456);
or U8859 (N_8859,N_7451,N_7626);
nand U8860 (N_8860,N_7602,N_7540);
nor U8861 (N_8861,N_7273,N_7732);
nor U8862 (N_8862,N_7436,N_7546);
nor U8863 (N_8863,N_7150,N_7184);
or U8864 (N_8864,N_7089,N_7480);
nor U8865 (N_8865,N_7839,N_7684);
xor U8866 (N_8866,N_7399,N_7486);
or U8867 (N_8867,N_7179,N_7734);
or U8868 (N_8868,N_7842,N_7831);
and U8869 (N_8869,N_7355,N_7578);
nor U8870 (N_8870,N_7040,N_7779);
nor U8871 (N_8871,N_7420,N_7414);
nor U8872 (N_8872,N_7472,N_7221);
and U8873 (N_8873,N_7113,N_7542);
nand U8874 (N_8874,N_7831,N_7103);
or U8875 (N_8875,N_7510,N_7016);
and U8876 (N_8876,N_7794,N_7725);
nand U8877 (N_8877,N_7198,N_7206);
or U8878 (N_8878,N_7531,N_7862);
nand U8879 (N_8879,N_7405,N_7618);
and U8880 (N_8880,N_7320,N_7044);
xor U8881 (N_8881,N_7238,N_7472);
nand U8882 (N_8882,N_7450,N_7142);
and U8883 (N_8883,N_7646,N_7294);
nor U8884 (N_8884,N_7215,N_7285);
or U8885 (N_8885,N_7772,N_7485);
and U8886 (N_8886,N_7890,N_7792);
nor U8887 (N_8887,N_7329,N_7448);
or U8888 (N_8888,N_7898,N_7343);
or U8889 (N_8889,N_7299,N_7221);
nor U8890 (N_8890,N_7623,N_7578);
or U8891 (N_8891,N_7772,N_7909);
nor U8892 (N_8892,N_7403,N_7228);
nand U8893 (N_8893,N_7139,N_7015);
nor U8894 (N_8894,N_7028,N_7503);
and U8895 (N_8895,N_7929,N_7754);
nor U8896 (N_8896,N_7875,N_7202);
or U8897 (N_8897,N_7970,N_7341);
nand U8898 (N_8898,N_7194,N_7178);
nand U8899 (N_8899,N_7443,N_7868);
and U8900 (N_8900,N_7050,N_7179);
or U8901 (N_8901,N_7081,N_7125);
nor U8902 (N_8902,N_7995,N_7436);
nand U8903 (N_8903,N_7350,N_7742);
xor U8904 (N_8904,N_7594,N_7945);
nor U8905 (N_8905,N_7941,N_7119);
nand U8906 (N_8906,N_7499,N_7801);
nor U8907 (N_8907,N_7559,N_7029);
nand U8908 (N_8908,N_7524,N_7904);
and U8909 (N_8909,N_7889,N_7054);
nand U8910 (N_8910,N_7943,N_7429);
nand U8911 (N_8911,N_7429,N_7449);
nor U8912 (N_8912,N_7426,N_7205);
nand U8913 (N_8913,N_7512,N_7029);
xnor U8914 (N_8914,N_7343,N_7910);
nor U8915 (N_8915,N_7482,N_7498);
xnor U8916 (N_8916,N_7282,N_7924);
and U8917 (N_8917,N_7045,N_7819);
and U8918 (N_8918,N_7136,N_7656);
or U8919 (N_8919,N_7319,N_7816);
xor U8920 (N_8920,N_7903,N_7547);
nand U8921 (N_8921,N_7872,N_7421);
and U8922 (N_8922,N_7274,N_7147);
or U8923 (N_8923,N_7778,N_7687);
or U8924 (N_8924,N_7509,N_7222);
and U8925 (N_8925,N_7338,N_7226);
or U8926 (N_8926,N_7559,N_7377);
nor U8927 (N_8927,N_7435,N_7683);
and U8928 (N_8928,N_7166,N_7602);
nor U8929 (N_8929,N_7681,N_7395);
or U8930 (N_8930,N_7854,N_7841);
nor U8931 (N_8931,N_7892,N_7712);
nor U8932 (N_8932,N_7605,N_7812);
nor U8933 (N_8933,N_7537,N_7406);
xor U8934 (N_8934,N_7979,N_7819);
nand U8935 (N_8935,N_7202,N_7298);
xnor U8936 (N_8936,N_7795,N_7978);
nor U8937 (N_8937,N_7219,N_7025);
and U8938 (N_8938,N_7074,N_7229);
nor U8939 (N_8939,N_7082,N_7753);
xnor U8940 (N_8940,N_7053,N_7812);
or U8941 (N_8941,N_7430,N_7637);
or U8942 (N_8942,N_7699,N_7135);
or U8943 (N_8943,N_7763,N_7036);
nor U8944 (N_8944,N_7204,N_7594);
or U8945 (N_8945,N_7147,N_7081);
nand U8946 (N_8946,N_7539,N_7437);
and U8947 (N_8947,N_7443,N_7772);
or U8948 (N_8948,N_7203,N_7089);
nor U8949 (N_8949,N_7997,N_7743);
xor U8950 (N_8950,N_7184,N_7739);
and U8951 (N_8951,N_7936,N_7081);
nor U8952 (N_8952,N_7933,N_7643);
nor U8953 (N_8953,N_7461,N_7166);
nand U8954 (N_8954,N_7196,N_7663);
and U8955 (N_8955,N_7989,N_7987);
or U8956 (N_8956,N_7483,N_7357);
xor U8957 (N_8957,N_7357,N_7983);
or U8958 (N_8958,N_7804,N_7517);
or U8959 (N_8959,N_7434,N_7799);
and U8960 (N_8960,N_7324,N_7356);
nand U8961 (N_8961,N_7186,N_7261);
or U8962 (N_8962,N_7608,N_7056);
and U8963 (N_8963,N_7549,N_7433);
and U8964 (N_8964,N_7937,N_7320);
nand U8965 (N_8965,N_7000,N_7599);
nand U8966 (N_8966,N_7255,N_7464);
nor U8967 (N_8967,N_7080,N_7057);
nor U8968 (N_8968,N_7599,N_7716);
and U8969 (N_8969,N_7088,N_7019);
and U8970 (N_8970,N_7100,N_7483);
nand U8971 (N_8971,N_7690,N_7763);
nand U8972 (N_8972,N_7565,N_7345);
nand U8973 (N_8973,N_7238,N_7004);
nand U8974 (N_8974,N_7086,N_7625);
nand U8975 (N_8975,N_7004,N_7900);
nand U8976 (N_8976,N_7164,N_7302);
or U8977 (N_8977,N_7157,N_7315);
nor U8978 (N_8978,N_7794,N_7262);
and U8979 (N_8979,N_7538,N_7641);
or U8980 (N_8980,N_7692,N_7928);
or U8981 (N_8981,N_7468,N_7241);
or U8982 (N_8982,N_7878,N_7429);
nand U8983 (N_8983,N_7979,N_7302);
or U8984 (N_8984,N_7192,N_7682);
and U8985 (N_8985,N_7099,N_7508);
nand U8986 (N_8986,N_7141,N_7457);
nand U8987 (N_8987,N_7657,N_7301);
or U8988 (N_8988,N_7985,N_7758);
or U8989 (N_8989,N_7688,N_7791);
nand U8990 (N_8990,N_7571,N_7542);
nor U8991 (N_8991,N_7425,N_7061);
and U8992 (N_8992,N_7124,N_7544);
nor U8993 (N_8993,N_7070,N_7382);
and U8994 (N_8994,N_7254,N_7302);
nand U8995 (N_8995,N_7637,N_7766);
nor U8996 (N_8996,N_7185,N_7267);
and U8997 (N_8997,N_7185,N_7022);
nand U8998 (N_8998,N_7300,N_7329);
nand U8999 (N_8999,N_7430,N_7097);
and U9000 (N_9000,N_8589,N_8247);
nand U9001 (N_9001,N_8685,N_8532);
or U9002 (N_9002,N_8785,N_8106);
nand U9003 (N_9003,N_8397,N_8241);
nor U9004 (N_9004,N_8217,N_8859);
xnor U9005 (N_9005,N_8238,N_8497);
or U9006 (N_9006,N_8839,N_8662);
nand U9007 (N_9007,N_8439,N_8700);
nor U9008 (N_9008,N_8597,N_8009);
or U9009 (N_9009,N_8516,N_8572);
or U9010 (N_9010,N_8774,N_8014);
xor U9011 (N_9011,N_8707,N_8153);
nor U9012 (N_9012,N_8187,N_8354);
nand U9013 (N_9013,N_8942,N_8491);
nor U9014 (N_9014,N_8133,N_8436);
nor U9015 (N_9015,N_8146,N_8568);
and U9016 (N_9016,N_8547,N_8297);
nand U9017 (N_9017,N_8914,N_8664);
xor U9018 (N_9018,N_8824,N_8886);
nand U9019 (N_9019,N_8968,N_8470);
or U9020 (N_9020,N_8925,N_8251);
or U9021 (N_9021,N_8038,N_8699);
or U9022 (N_9022,N_8538,N_8602);
nand U9023 (N_9023,N_8035,N_8503);
nor U9024 (N_9024,N_8471,N_8459);
nor U9025 (N_9025,N_8412,N_8943);
nor U9026 (N_9026,N_8273,N_8402);
nor U9027 (N_9027,N_8884,N_8403);
or U9028 (N_9028,N_8766,N_8825);
or U9029 (N_9029,N_8642,N_8213);
nor U9030 (N_9030,N_8335,N_8831);
and U9031 (N_9031,N_8566,N_8904);
nor U9032 (N_9032,N_8789,N_8716);
and U9033 (N_9033,N_8544,N_8132);
nand U9034 (N_9034,N_8546,N_8718);
nand U9035 (N_9035,N_8940,N_8793);
or U9036 (N_9036,N_8350,N_8620);
xor U9037 (N_9037,N_8137,N_8918);
and U9038 (N_9038,N_8446,N_8261);
nor U9039 (N_9039,N_8314,N_8590);
nor U9040 (N_9040,N_8042,N_8263);
nor U9041 (N_9041,N_8696,N_8433);
and U9042 (N_9042,N_8603,N_8582);
and U9043 (N_9043,N_8573,N_8254);
xnor U9044 (N_9044,N_8521,N_8967);
and U9045 (N_9045,N_8265,N_8299);
nand U9046 (N_9046,N_8026,N_8478);
or U9047 (N_9047,N_8746,N_8847);
nor U9048 (N_9048,N_8311,N_8910);
nor U9049 (N_9049,N_8370,N_8322);
xnor U9050 (N_9050,N_8577,N_8670);
and U9051 (N_9051,N_8535,N_8448);
and U9052 (N_9052,N_8358,N_8690);
and U9053 (N_9053,N_8072,N_8821);
or U9054 (N_9054,N_8644,N_8632);
and U9055 (N_9055,N_8180,N_8906);
xor U9056 (N_9056,N_8722,N_8103);
nand U9057 (N_9057,N_8396,N_8932);
nor U9058 (N_9058,N_8159,N_8430);
nand U9059 (N_9059,N_8554,N_8239);
nor U9060 (N_9060,N_8958,N_8729);
xnor U9061 (N_9061,N_8861,N_8426);
or U9062 (N_9062,N_8731,N_8684);
and U9063 (N_9063,N_8449,N_8329);
nor U9064 (N_9064,N_8024,N_8078);
or U9065 (N_9065,N_8246,N_8605);
nand U9066 (N_9066,N_8594,N_8668);
and U9067 (N_9067,N_8807,N_8899);
and U9068 (N_9068,N_8306,N_8303);
nand U9069 (N_9069,N_8182,N_8530);
and U9070 (N_9070,N_8541,N_8081);
or U9071 (N_9071,N_8252,N_8977);
and U9072 (N_9072,N_8117,N_8666);
and U9073 (N_9073,N_8327,N_8211);
and U9074 (N_9074,N_8628,N_8361);
or U9075 (N_9075,N_8293,N_8665);
nand U9076 (N_9076,N_8695,N_8074);
nor U9077 (N_9077,N_8416,N_8274);
nor U9078 (N_9078,N_8488,N_8971);
nor U9079 (N_9079,N_8498,N_8333);
nor U9080 (N_9080,N_8156,N_8797);
or U9081 (N_9081,N_8836,N_8870);
nand U9082 (N_9082,N_8601,N_8184);
nand U9083 (N_9083,N_8984,N_8704);
and U9084 (N_9084,N_8121,N_8320);
nand U9085 (N_9085,N_8075,N_8619);
nand U9086 (N_9086,N_8893,N_8673);
and U9087 (N_9087,N_8931,N_8805);
nor U9088 (N_9088,N_8959,N_8413);
and U9089 (N_9089,N_8260,N_8876);
nand U9090 (N_9090,N_8130,N_8466);
and U9091 (N_9091,N_8703,N_8759);
and U9092 (N_9092,N_8688,N_8202);
or U9093 (N_9093,N_8866,N_8450);
xor U9094 (N_9094,N_8083,N_8862);
nand U9095 (N_9095,N_8321,N_8525);
nor U9096 (N_9096,N_8843,N_8504);
nand U9097 (N_9097,N_8339,N_8622);
nand U9098 (N_9098,N_8835,N_8855);
nor U9099 (N_9099,N_8816,N_8970);
nand U9100 (N_9100,N_8697,N_8909);
or U9101 (N_9101,N_8745,N_8576);
nor U9102 (N_9102,N_8016,N_8828);
nor U9103 (N_9103,N_8302,N_8633);
or U9104 (N_9104,N_8519,N_8419);
and U9105 (N_9105,N_8868,N_8496);
nand U9106 (N_9106,N_8489,N_8853);
and U9107 (N_9107,N_8938,N_8750);
and U9108 (N_9108,N_8658,N_8134);
and U9109 (N_9109,N_8002,N_8772);
and U9110 (N_9110,N_8410,N_8988);
xnor U9111 (N_9111,N_8371,N_8362);
nand U9112 (N_9112,N_8343,N_8262);
xor U9113 (N_9113,N_8054,N_8815);
and U9114 (N_9114,N_8879,N_8983);
or U9115 (N_9115,N_8656,N_8860);
or U9116 (N_9116,N_8098,N_8513);
nor U9117 (N_9117,N_8721,N_8025);
and U9118 (N_9118,N_8972,N_8948);
nor U9119 (N_9119,N_8481,N_8288);
or U9120 (N_9120,N_8041,N_8553);
or U9121 (N_9121,N_8279,N_8749);
nand U9122 (N_9122,N_8381,N_8142);
nor U9123 (N_9123,N_8787,N_8874);
and U9124 (N_9124,N_8065,N_8015);
nor U9125 (N_9125,N_8119,N_8800);
nand U9126 (N_9126,N_8116,N_8349);
nor U9127 (N_9127,N_8719,N_8534);
or U9128 (N_9128,N_8593,N_8753);
nand U9129 (N_9129,N_8890,N_8526);
nor U9130 (N_9130,N_8201,N_8708);
and U9131 (N_9131,N_8198,N_8806);
or U9132 (N_9132,N_8369,N_8441);
xor U9133 (N_9133,N_8483,N_8732);
nor U9134 (N_9134,N_8230,N_8648);
nor U9135 (N_9135,N_8013,N_8200);
nor U9136 (N_9136,N_8484,N_8851);
or U9137 (N_9137,N_8376,N_8372);
or U9138 (N_9138,N_8487,N_8779);
or U9139 (N_9139,N_8640,N_8404);
and U9140 (N_9140,N_8267,N_8231);
xnor U9141 (N_9141,N_8569,N_8913);
nand U9142 (N_9142,N_8555,N_8196);
nand U9143 (N_9143,N_8928,N_8469);
nor U9144 (N_9144,N_8340,N_8924);
nand U9145 (N_9145,N_8889,N_8296);
and U9146 (N_9146,N_8687,N_8570);
nand U9147 (N_9147,N_8706,N_8011);
or U9148 (N_9148,N_8627,N_8395);
xnor U9149 (N_9149,N_8768,N_8990);
nand U9150 (N_9150,N_8680,N_8389);
nand U9151 (N_9151,N_8060,N_8586);
or U9152 (N_9152,N_8170,N_8794);
nor U9153 (N_9153,N_8945,N_8624);
and U9154 (N_9154,N_8391,N_8552);
or U9155 (N_9155,N_8382,N_8752);
or U9156 (N_9156,N_8682,N_8677);
nor U9157 (N_9157,N_8244,N_8558);
or U9158 (N_9158,N_8438,N_8423);
or U9159 (N_9159,N_8390,N_8715);
and U9160 (N_9160,N_8638,N_8177);
nor U9161 (N_9161,N_8937,N_8819);
and U9162 (N_9162,N_8653,N_8224);
nand U9163 (N_9163,N_8457,N_8309);
xor U9164 (N_9164,N_8255,N_8877);
nand U9165 (N_9165,N_8148,N_8092);
nor U9166 (N_9166,N_8277,N_8891);
or U9167 (N_9167,N_8218,N_8604);
nor U9168 (N_9168,N_8975,N_8406);
nor U9169 (N_9169,N_8456,N_8451);
nand U9170 (N_9170,N_8784,N_8220);
xor U9171 (N_9171,N_8115,N_8637);
nor U9172 (N_9172,N_8319,N_8803);
and U9173 (N_9173,N_8888,N_8935);
nor U9174 (N_9174,N_8947,N_8055);
nand U9175 (N_9175,N_8344,N_8878);
or U9176 (N_9176,N_8674,N_8233);
nand U9177 (N_9177,N_8834,N_8592);
xor U9178 (N_9178,N_8829,N_8776);
nor U9179 (N_9179,N_8561,N_8240);
and U9180 (N_9180,N_8974,N_8867);
and U9181 (N_9181,N_8109,N_8956);
nand U9182 (N_9182,N_8997,N_8986);
nor U9183 (N_9183,N_8671,N_8926);
or U9184 (N_9184,N_8048,N_8623);
nor U9185 (N_9185,N_8463,N_8268);
nand U9186 (N_9186,N_8307,N_8502);
or U9187 (N_9187,N_8388,N_8650);
and U9188 (N_9188,N_8095,N_8737);
nand U9189 (N_9189,N_8005,N_8363);
xor U9190 (N_9190,N_8961,N_8540);
nor U9191 (N_9191,N_8581,N_8352);
xnor U9192 (N_9192,N_8373,N_8565);
and U9193 (N_9193,N_8635,N_8822);
nor U9194 (N_9194,N_8085,N_8995);
or U9195 (N_9195,N_8023,N_8675);
nand U9196 (N_9196,N_8346,N_8848);
nor U9197 (N_9197,N_8248,N_8814);
or U9198 (N_9198,N_8162,N_8809);
nor U9199 (N_9199,N_8567,N_8813);
nand U9200 (N_9200,N_8840,N_8705);
or U9201 (N_9201,N_8222,N_8799);
or U9202 (N_9202,N_8464,N_8377);
or U9203 (N_9203,N_8885,N_8102);
xor U9204 (N_9204,N_8571,N_8712);
nand U9205 (N_9205,N_8392,N_8325);
nand U9206 (N_9206,N_8923,N_8844);
and U9207 (N_9207,N_8122,N_8740);
nand U9208 (N_9208,N_8387,N_8149);
nor U9209 (N_9209,N_8963,N_8077);
nor U9210 (N_9210,N_8154,N_8667);
and U9211 (N_9211,N_8892,N_8398);
xor U9212 (N_9212,N_8097,N_8061);
or U9213 (N_9213,N_8533,N_8140);
nand U9214 (N_9214,N_8930,N_8973);
xnor U9215 (N_9215,N_8003,N_8786);
xor U9216 (N_9216,N_8120,N_8345);
xnor U9217 (N_9217,N_8294,N_8017);
nand U9218 (N_9218,N_8950,N_8318);
or U9219 (N_9219,N_8756,N_8384);
nand U9220 (N_9220,N_8617,N_8127);
and U9221 (N_9221,N_8754,N_8903);
nand U9222 (N_9222,N_8429,N_8506);
or U9223 (N_9223,N_8138,N_8071);
nor U9224 (N_9224,N_8219,N_8427);
nor U9225 (N_9225,N_8164,N_8175);
nand U9226 (N_9226,N_8068,N_8812);
or U9227 (N_9227,N_8452,N_8804);
nand U9228 (N_9228,N_8278,N_8724);
xnor U9229 (N_9229,N_8486,N_8052);
and U9230 (N_9230,N_8315,N_8039);
or U9231 (N_9231,N_8720,N_8713);
nor U9232 (N_9232,N_8698,N_8528);
xnor U9233 (N_9233,N_8147,N_8043);
xor U9234 (N_9234,N_8099,N_8036);
and U9235 (N_9235,N_8953,N_8336);
and U9236 (N_9236,N_8905,N_8801);
nor U9237 (N_9237,N_8215,N_8560);
nor U9238 (N_9238,N_8911,N_8292);
nor U9239 (N_9239,N_8357,N_8225);
nand U9240 (N_9240,N_8764,N_8190);
xor U9241 (N_9241,N_8442,N_8195);
and U9242 (N_9242,N_8778,N_8505);
nor U9243 (N_9243,N_8790,N_8181);
and U9244 (N_9244,N_8987,N_8992);
nand U9245 (N_9245,N_8508,N_8204);
xor U9246 (N_9246,N_8155,N_8123);
or U9247 (N_9247,N_8701,N_8500);
nand U9248 (N_9248,N_8286,N_8751);
nand U9249 (N_9249,N_8902,N_8270);
nand U9250 (N_9250,N_8460,N_8385);
nor U9251 (N_9251,N_8735,N_8976);
nand U9252 (N_9252,N_8414,N_8520);
nand U9253 (N_9253,N_8837,N_8331);
nand U9254 (N_9254,N_8762,N_8771);
or U9255 (N_9255,N_8356,N_8151);
nand U9256 (N_9256,N_8050,N_8069);
nand U9257 (N_9257,N_8205,N_8145);
and U9258 (N_9258,N_8418,N_8305);
or U9259 (N_9259,N_8129,N_8514);
and U9260 (N_9260,N_8587,N_8474);
nand U9261 (N_9261,N_8743,N_8375);
or U9262 (N_9262,N_8453,N_8490);
xor U9263 (N_9263,N_8609,N_8511);
xor U9264 (N_9264,N_8782,N_8432);
nor U9265 (N_9265,N_8539,N_8872);
nand U9266 (N_9266,N_8507,N_8324);
or U9267 (N_9267,N_8264,N_8135);
nor U9268 (N_9268,N_8818,N_8157);
nand U9269 (N_9269,N_8018,N_8199);
nand U9270 (N_9270,N_8266,N_8304);
nand U9271 (N_9271,N_8606,N_8854);
nor U9272 (N_9272,N_8780,N_8317);
and U9273 (N_9273,N_8019,N_8501);
nand U9274 (N_9274,N_8034,N_8598);
and U9275 (N_9275,N_8841,N_8168);
or U9276 (N_9276,N_8982,N_8351);
nand U9277 (N_9277,N_8447,N_8733);
xor U9278 (N_9278,N_8249,N_8143);
nand U9279 (N_9279,N_8536,N_8871);
or U9280 (N_9280,N_8634,N_8179);
nand U9281 (N_9281,N_8066,N_8059);
and U9282 (N_9282,N_8091,N_8517);
nand U9283 (N_9283,N_8300,N_8367);
or U9284 (N_9284,N_8022,N_8028);
nor U9285 (N_9285,N_8941,N_8461);
or U9286 (N_9286,N_8951,N_8400);
xor U9287 (N_9287,N_8214,N_8237);
and U9288 (N_9288,N_8939,N_8747);
or U9289 (N_9289,N_8607,N_8082);
and U9290 (N_9290,N_8725,N_8070);
or U9291 (N_9291,N_8613,N_8921);
or U9292 (N_9292,N_8655,N_8915);
nor U9293 (N_9293,N_8796,N_8394);
or U9294 (N_9294,N_8473,N_8944);
nand U9295 (N_9295,N_8313,N_8462);
and U9296 (N_9296,N_8010,N_8887);
nor U9297 (N_9297,N_8284,N_8518);
or U9298 (N_9298,N_8647,N_8485);
nor U9299 (N_9299,N_8599,N_8171);
and U9300 (N_9300,N_8272,N_8849);
nor U9301 (N_9301,N_8857,N_8527);
and U9302 (N_9302,N_8679,N_8291);
nand U9303 (N_9303,N_8591,N_8999);
nor U9304 (N_9304,N_8046,N_8657);
nor U9305 (N_9305,N_8229,N_8386);
nand U9306 (N_9306,N_8901,N_8374);
and U9307 (N_9307,N_8194,N_8775);
nand U9308 (N_9308,N_8985,N_8104);
nand U9309 (N_9309,N_8649,N_8420);
nor U9310 (N_9310,N_8777,N_8580);
nand U9311 (N_9311,N_8206,N_8158);
xor U9312 (N_9312,N_8087,N_8476);
nor U9313 (N_9313,N_8960,N_8257);
nand U9314 (N_9314,N_8833,N_8323);
xnor U9315 (N_9315,N_8838,N_8614);
nor U9316 (N_9316,N_8118,N_8223);
and U9317 (N_9317,N_8949,N_8730);
nor U9318 (N_9318,N_8437,N_8186);
nor U9319 (N_9319,N_8669,N_8636);
or U9320 (N_9320,N_8191,N_8101);
xor U9321 (N_9321,N_8826,N_8643);
xor U9322 (N_9322,N_8165,N_8978);
nand U9323 (N_9323,N_8531,N_8062);
or U9324 (N_9324,N_8900,N_8625);
and U9325 (N_9325,N_8672,N_8342);
nand U9326 (N_9326,N_8894,N_8676);
nor U9327 (N_9327,N_8160,N_8711);
nand U9328 (N_9328,N_8269,N_8758);
nor U9329 (N_9329,N_8608,N_8610);
nand U9330 (N_9330,N_8250,N_8810);
and U9331 (N_9331,N_8966,N_8334);
nand U9332 (N_9332,N_8310,N_8600);
xnor U9333 (N_9333,N_8094,N_8480);
xor U9334 (N_9334,N_8049,N_8341);
nor U9335 (N_9335,N_8864,N_8290);
nand U9336 (N_9336,N_8033,N_8316);
and U9337 (N_9337,N_8629,N_8896);
nor U9338 (N_9338,N_8053,N_8209);
and U9339 (N_9339,N_8051,N_8128);
xnor U9340 (N_9340,N_8090,N_8916);
nor U9341 (N_9341,N_8969,N_8898);
or U9342 (N_9342,N_8652,N_8285);
nand U9343 (N_9343,N_8631,N_8193);
nor U9344 (N_9344,N_8755,N_8616);
nor U9345 (N_9345,N_8301,N_8981);
nand U9346 (N_9346,N_8692,N_8236);
nand U9347 (N_9347,N_8611,N_8739);
nand U9348 (N_9348,N_8686,N_8742);
or U9349 (N_9349,N_8359,N_8980);
or U9350 (N_9350,N_8817,N_8152);
or U9351 (N_9351,N_8783,N_8492);
nor U9352 (N_9352,N_8773,N_8086);
nand U9353 (N_9353,N_8588,N_8365);
nor U9354 (N_9354,N_8630,N_8258);
nor U9355 (N_9355,N_8031,N_8691);
and U9356 (N_9356,N_8208,N_8020);
nand U9357 (N_9357,N_8523,N_8475);
nand U9358 (N_9358,N_8595,N_8056);
nor U9359 (N_9359,N_8654,N_8661);
or U9360 (N_9360,N_8173,N_8559);
nand U9361 (N_9361,N_8702,N_8161);
and U9362 (N_9362,N_8431,N_8612);
nand U9363 (N_9363,N_8144,N_8934);
or U9364 (N_9364,N_8563,N_8422);
and U9365 (N_9365,N_8421,N_8651);
nand U9366 (N_9366,N_8873,N_8936);
and U9367 (N_9367,N_8998,N_8100);
or U9368 (N_9368,N_8364,N_8232);
or U9369 (N_9369,N_8626,N_8378);
or U9370 (N_9370,N_8348,N_8126);
or U9371 (N_9371,N_8467,N_8929);
nand U9372 (N_9372,N_8615,N_8477);
nor U9373 (N_9373,N_8407,N_8820);
nand U9374 (N_9374,N_8096,N_8618);
and U9375 (N_9375,N_8113,N_8079);
or U9376 (N_9376,N_8047,N_8827);
nor U9377 (N_9377,N_8338,N_8174);
and U9378 (N_9378,N_8908,N_8681);
and U9379 (N_9379,N_8808,N_8761);
or U9380 (N_9380,N_8522,N_8207);
nor U9381 (N_9381,N_8032,N_8326);
or U9382 (N_9382,N_8283,N_8089);
and U9383 (N_9383,N_8007,N_8548);
and U9384 (N_9384,N_8166,N_8012);
or U9385 (N_9385,N_8869,N_8289);
and U9386 (N_9386,N_8366,N_8842);
nor U9387 (N_9387,N_8424,N_8596);
and U9388 (N_9388,N_8399,N_8802);
nor U9389 (N_9389,N_8646,N_8434);
or U9390 (N_9390,N_8578,N_8203);
or U9391 (N_9391,N_8280,N_8188);
nand U9392 (N_9392,N_8259,N_8245);
nand U9393 (N_9393,N_8337,N_8212);
nor U9394 (N_9394,N_8411,N_8445);
nand U9395 (N_9395,N_8993,N_8221);
and U9396 (N_9396,N_8858,N_8763);
nand U9397 (N_9397,N_8380,N_8564);
xnor U9398 (N_9398,N_8183,N_8178);
or U9399 (N_9399,N_8131,N_8881);
or U9400 (N_9400,N_8659,N_8883);
nor U9401 (N_9401,N_8465,N_8111);
or U9402 (N_9402,N_8425,N_8714);
and U9403 (N_9403,N_8328,N_8845);
and U9404 (N_9404,N_8176,N_8040);
or U9405 (N_9405,N_8063,N_8922);
and U9406 (N_9406,N_8493,N_8748);
and U9407 (N_9407,N_8726,N_8927);
or U9408 (N_9408,N_8458,N_8006);
nand U9409 (N_9409,N_8917,N_8996);
nor U9410 (N_9410,N_8717,N_8830);
nor U9411 (N_9411,N_8585,N_8863);
and U9412 (N_9412,N_8537,N_8639);
and U9413 (N_9413,N_8964,N_8989);
nand U9414 (N_9414,N_8192,N_8645);
nor U9415 (N_9415,N_8791,N_8004);
and U9416 (N_9416,N_8689,N_8955);
and U9417 (N_9417,N_8744,N_8515);
or U9418 (N_9418,N_8045,N_8169);
nor U9419 (N_9419,N_8124,N_8562);
xnor U9420 (N_9420,N_8621,N_8027);
nand U9421 (N_9421,N_8393,N_8865);
nor U9422 (N_9422,N_8556,N_8355);
nor U9423 (N_9423,N_8308,N_8275);
and U9424 (N_9424,N_8415,N_8727);
nand U9425 (N_9425,N_8112,N_8295);
nand U9426 (N_9426,N_8472,N_8058);
and U9427 (N_9427,N_8347,N_8736);
and U9428 (N_9428,N_8545,N_8660);
and U9429 (N_9429,N_8443,N_8440);
nor U9430 (N_9430,N_8454,N_8912);
nor U9431 (N_9431,N_8907,N_8543);
nand U9432 (N_9432,N_8788,N_8683);
nor U9433 (N_9433,N_8850,N_8379);
and U9434 (N_9434,N_8029,N_8228);
or U9435 (N_9435,N_8076,N_8979);
nor U9436 (N_9436,N_8678,N_8575);
nor U9437 (N_9437,N_8852,N_8084);
nand U9438 (N_9438,N_8216,N_8769);
nand U9439 (N_9439,N_8455,N_8723);
nand U9440 (N_9440,N_8281,N_8067);
and U9441 (N_9441,N_8882,N_8210);
or U9442 (N_9442,N_8125,N_8494);
nor U9443 (N_9443,N_8920,N_8479);
nand U9444 (N_9444,N_8312,N_8197);
nand U9445 (N_9445,N_8435,N_8542);
and U9446 (N_9446,N_8509,N_8163);
nor U9447 (N_9447,N_8405,N_8172);
nor U9448 (N_9448,N_8846,N_8080);
nor U9449 (N_9449,N_8954,N_8811);
and U9450 (N_9450,N_8332,N_8551);
nor U9451 (N_9451,N_8495,N_8510);
nand U9452 (N_9452,N_8141,N_8136);
nor U9453 (N_9453,N_8710,N_8428);
or U9454 (N_9454,N_8583,N_8298);
nor U9455 (N_9455,N_8353,N_8895);
nor U9456 (N_9456,N_8287,N_8057);
and U9457 (N_9457,N_8037,N_8417);
and U9458 (N_9458,N_8167,N_8088);
or U9459 (N_9459,N_8952,N_8073);
nor U9460 (N_9460,N_8897,N_8957);
nand U9461 (N_9461,N_8757,N_8021);
nand U9462 (N_9462,N_8933,N_8962);
and U9463 (N_9463,N_8741,N_8641);
or U9464 (N_9464,N_8767,N_8064);
nor U9465 (N_9465,N_8919,N_8512);
xnor U9466 (N_9466,N_8107,N_8242);
nor U9467 (N_9467,N_8000,N_8253);
and U9468 (N_9468,N_8549,N_8738);
nor U9469 (N_9469,N_8368,N_8770);
or U9470 (N_9470,N_8584,N_8781);
nand U9471 (N_9471,N_8044,N_8408);
nor U9472 (N_9472,N_8832,N_8282);
nor U9473 (N_9473,N_8765,N_8150);
nand U9474 (N_9474,N_8524,N_8574);
nand U9475 (N_9475,N_8734,N_8482);
or U9476 (N_9476,N_8139,N_8001);
xor U9477 (N_9477,N_8360,N_8189);
and U9478 (N_9478,N_8256,N_8798);
and U9479 (N_9479,N_8235,N_8693);
and U9480 (N_9480,N_8994,N_8795);
xor U9481 (N_9481,N_8856,N_8105);
nor U9482 (N_9482,N_8709,N_8880);
nand U9483 (N_9483,N_8243,N_8409);
nor U9484 (N_9484,N_8694,N_8468);
nor U9485 (N_9485,N_8226,N_8185);
or U9486 (N_9486,N_8276,N_8227);
or U9487 (N_9487,N_8444,N_8383);
nand U9488 (N_9488,N_8946,N_8875);
xor U9489 (N_9489,N_8110,N_8499);
nand U9490 (N_9490,N_8823,N_8114);
nand U9491 (N_9491,N_8557,N_8965);
or U9492 (N_9492,N_8728,N_8529);
nor U9493 (N_9493,N_8991,N_8401);
xor U9494 (N_9494,N_8030,N_8234);
nand U9495 (N_9495,N_8330,N_8550);
or U9496 (N_9496,N_8792,N_8760);
nand U9497 (N_9497,N_8108,N_8093);
and U9498 (N_9498,N_8579,N_8008);
nand U9499 (N_9499,N_8271,N_8663);
and U9500 (N_9500,N_8472,N_8646);
nand U9501 (N_9501,N_8861,N_8393);
and U9502 (N_9502,N_8373,N_8518);
and U9503 (N_9503,N_8029,N_8785);
or U9504 (N_9504,N_8930,N_8308);
and U9505 (N_9505,N_8767,N_8386);
and U9506 (N_9506,N_8982,N_8236);
or U9507 (N_9507,N_8412,N_8770);
nand U9508 (N_9508,N_8934,N_8644);
nand U9509 (N_9509,N_8447,N_8207);
nand U9510 (N_9510,N_8529,N_8730);
and U9511 (N_9511,N_8329,N_8050);
nand U9512 (N_9512,N_8208,N_8113);
or U9513 (N_9513,N_8584,N_8495);
nor U9514 (N_9514,N_8370,N_8888);
or U9515 (N_9515,N_8748,N_8120);
and U9516 (N_9516,N_8633,N_8547);
nand U9517 (N_9517,N_8850,N_8706);
or U9518 (N_9518,N_8779,N_8785);
or U9519 (N_9519,N_8756,N_8491);
and U9520 (N_9520,N_8343,N_8602);
nand U9521 (N_9521,N_8969,N_8011);
nor U9522 (N_9522,N_8297,N_8399);
and U9523 (N_9523,N_8205,N_8968);
or U9524 (N_9524,N_8352,N_8707);
xor U9525 (N_9525,N_8091,N_8309);
nor U9526 (N_9526,N_8393,N_8302);
and U9527 (N_9527,N_8778,N_8027);
or U9528 (N_9528,N_8730,N_8235);
nor U9529 (N_9529,N_8450,N_8455);
or U9530 (N_9530,N_8584,N_8396);
or U9531 (N_9531,N_8575,N_8552);
or U9532 (N_9532,N_8564,N_8833);
and U9533 (N_9533,N_8120,N_8525);
and U9534 (N_9534,N_8831,N_8918);
or U9535 (N_9535,N_8806,N_8290);
and U9536 (N_9536,N_8425,N_8212);
nor U9537 (N_9537,N_8435,N_8989);
and U9538 (N_9538,N_8852,N_8029);
nand U9539 (N_9539,N_8135,N_8183);
or U9540 (N_9540,N_8910,N_8997);
and U9541 (N_9541,N_8736,N_8875);
and U9542 (N_9542,N_8414,N_8642);
nand U9543 (N_9543,N_8532,N_8517);
and U9544 (N_9544,N_8500,N_8400);
nand U9545 (N_9545,N_8536,N_8476);
xnor U9546 (N_9546,N_8958,N_8378);
nand U9547 (N_9547,N_8420,N_8451);
and U9548 (N_9548,N_8459,N_8410);
and U9549 (N_9549,N_8995,N_8939);
or U9550 (N_9550,N_8434,N_8992);
nor U9551 (N_9551,N_8227,N_8666);
or U9552 (N_9552,N_8164,N_8757);
nor U9553 (N_9553,N_8223,N_8833);
and U9554 (N_9554,N_8717,N_8212);
and U9555 (N_9555,N_8830,N_8575);
or U9556 (N_9556,N_8860,N_8926);
or U9557 (N_9557,N_8814,N_8886);
nand U9558 (N_9558,N_8739,N_8271);
xor U9559 (N_9559,N_8752,N_8113);
and U9560 (N_9560,N_8126,N_8185);
nand U9561 (N_9561,N_8288,N_8405);
and U9562 (N_9562,N_8086,N_8896);
nor U9563 (N_9563,N_8242,N_8108);
xor U9564 (N_9564,N_8497,N_8299);
and U9565 (N_9565,N_8797,N_8782);
and U9566 (N_9566,N_8469,N_8584);
nor U9567 (N_9567,N_8351,N_8173);
and U9568 (N_9568,N_8091,N_8297);
nand U9569 (N_9569,N_8301,N_8341);
or U9570 (N_9570,N_8136,N_8299);
nand U9571 (N_9571,N_8635,N_8756);
or U9572 (N_9572,N_8390,N_8595);
nor U9573 (N_9573,N_8273,N_8357);
or U9574 (N_9574,N_8922,N_8235);
nor U9575 (N_9575,N_8390,N_8876);
or U9576 (N_9576,N_8749,N_8454);
and U9577 (N_9577,N_8505,N_8671);
nor U9578 (N_9578,N_8211,N_8150);
nand U9579 (N_9579,N_8830,N_8257);
and U9580 (N_9580,N_8461,N_8244);
and U9581 (N_9581,N_8717,N_8135);
nor U9582 (N_9582,N_8884,N_8418);
or U9583 (N_9583,N_8272,N_8098);
or U9584 (N_9584,N_8467,N_8297);
and U9585 (N_9585,N_8323,N_8645);
or U9586 (N_9586,N_8106,N_8753);
or U9587 (N_9587,N_8286,N_8919);
nand U9588 (N_9588,N_8025,N_8089);
nor U9589 (N_9589,N_8974,N_8436);
and U9590 (N_9590,N_8447,N_8049);
nand U9591 (N_9591,N_8832,N_8312);
nor U9592 (N_9592,N_8032,N_8838);
nand U9593 (N_9593,N_8374,N_8171);
nor U9594 (N_9594,N_8309,N_8889);
or U9595 (N_9595,N_8422,N_8806);
and U9596 (N_9596,N_8697,N_8032);
xor U9597 (N_9597,N_8280,N_8655);
nand U9598 (N_9598,N_8333,N_8982);
nor U9599 (N_9599,N_8993,N_8202);
xor U9600 (N_9600,N_8819,N_8735);
nor U9601 (N_9601,N_8204,N_8342);
nor U9602 (N_9602,N_8215,N_8286);
and U9603 (N_9603,N_8210,N_8711);
xor U9604 (N_9604,N_8962,N_8199);
nand U9605 (N_9605,N_8391,N_8660);
nand U9606 (N_9606,N_8895,N_8301);
and U9607 (N_9607,N_8233,N_8361);
and U9608 (N_9608,N_8736,N_8621);
or U9609 (N_9609,N_8278,N_8965);
nand U9610 (N_9610,N_8407,N_8287);
nand U9611 (N_9611,N_8856,N_8864);
nor U9612 (N_9612,N_8313,N_8862);
xnor U9613 (N_9613,N_8847,N_8687);
nand U9614 (N_9614,N_8375,N_8710);
or U9615 (N_9615,N_8019,N_8695);
and U9616 (N_9616,N_8555,N_8277);
xor U9617 (N_9617,N_8218,N_8329);
and U9618 (N_9618,N_8647,N_8938);
xor U9619 (N_9619,N_8071,N_8648);
nand U9620 (N_9620,N_8948,N_8564);
or U9621 (N_9621,N_8334,N_8585);
and U9622 (N_9622,N_8730,N_8511);
or U9623 (N_9623,N_8489,N_8087);
or U9624 (N_9624,N_8347,N_8066);
and U9625 (N_9625,N_8755,N_8542);
nor U9626 (N_9626,N_8199,N_8790);
nor U9627 (N_9627,N_8326,N_8140);
or U9628 (N_9628,N_8440,N_8175);
or U9629 (N_9629,N_8060,N_8037);
and U9630 (N_9630,N_8266,N_8760);
or U9631 (N_9631,N_8092,N_8397);
or U9632 (N_9632,N_8623,N_8851);
xnor U9633 (N_9633,N_8375,N_8272);
nor U9634 (N_9634,N_8366,N_8959);
and U9635 (N_9635,N_8425,N_8704);
and U9636 (N_9636,N_8310,N_8289);
or U9637 (N_9637,N_8169,N_8930);
and U9638 (N_9638,N_8724,N_8445);
nand U9639 (N_9639,N_8630,N_8804);
nand U9640 (N_9640,N_8595,N_8360);
nor U9641 (N_9641,N_8041,N_8176);
and U9642 (N_9642,N_8730,N_8776);
nor U9643 (N_9643,N_8048,N_8809);
xor U9644 (N_9644,N_8631,N_8394);
nor U9645 (N_9645,N_8913,N_8951);
or U9646 (N_9646,N_8139,N_8294);
nand U9647 (N_9647,N_8010,N_8115);
or U9648 (N_9648,N_8662,N_8205);
nand U9649 (N_9649,N_8687,N_8521);
nand U9650 (N_9650,N_8111,N_8459);
nand U9651 (N_9651,N_8651,N_8412);
nand U9652 (N_9652,N_8364,N_8200);
xnor U9653 (N_9653,N_8982,N_8303);
and U9654 (N_9654,N_8888,N_8371);
xor U9655 (N_9655,N_8382,N_8403);
nor U9656 (N_9656,N_8910,N_8212);
and U9657 (N_9657,N_8888,N_8989);
nor U9658 (N_9658,N_8854,N_8475);
or U9659 (N_9659,N_8599,N_8644);
nor U9660 (N_9660,N_8847,N_8994);
nor U9661 (N_9661,N_8008,N_8842);
nand U9662 (N_9662,N_8020,N_8002);
nand U9663 (N_9663,N_8184,N_8372);
and U9664 (N_9664,N_8561,N_8872);
and U9665 (N_9665,N_8078,N_8952);
and U9666 (N_9666,N_8277,N_8964);
and U9667 (N_9667,N_8767,N_8512);
and U9668 (N_9668,N_8853,N_8339);
nor U9669 (N_9669,N_8942,N_8378);
and U9670 (N_9670,N_8112,N_8455);
or U9671 (N_9671,N_8115,N_8764);
nor U9672 (N_9672,N_8599,N_8463);
and U9673 (N_9673,N_8060,N_8134);
and U9674 (N_9674,N_8463,N_8700);
nor U9675 (N_9675,N_8599,N_8568);
nand U9676 (N_9676,N_8889,N_8842);
or U9677 (N_9677,N_8017,N_8953);
and U9678 (N_9678,N_8256,N_8156);
nand U9679 (N_9679,N_8000,N_8142);
or U9680 (N_9680,N_8023,N_8609);
nand U9681 (N_9681,N_8064,N_8222);
nand U9682 (N_9682,N_8577,N_8419);
nor U9683 (N_9683,N_8731,N_8761);
and U9684 (N_9684,N_8237,N_8881);
nand U9685 (N_9685,N_8957,N_8254);
nand U9686 (N_9686,N_8812,N_8448);
or U9687 (N_9687,N_8388,N_8834);
and U9688 (N_9688,N_8153,N_8732);
nand U9689 (N_9689,N_8931,N_8700);
and U9690 (N_9690,N_8712,N_8115);
xor U9691 (N_9691,N_8971,N_8093);
nand U9692 (N_9692,N_8730,N_8840);
nand U9693 (N_9693,N_8140,N_8702);
nor U9694 (N_9694,N_8280,N_8099);
nor U9695 (N_9695,N_8690,N_8808);
nor U9696 (N_9696,N_8356,N_8963);
nand U9697 (N_9697,N_8705,N_8347);
and U9698 (N_9698,N_8765,N_8609);
xnor U9699 (N_9699,N_8502,N_8507);
and U9700 (N_9700,N_8308,N_8862);
or U9701 (N_9701,N_8656,N_8466);
nor U9702 (N_9702,N_8167,N_8703);
or U9703 (N_9703,N_8124,N_8037);
and U9704 (N_9704,N_8696,N_8278);
and U9705 (N_9705,N_8160,N_8655);
xnor U9706 (N_9706,N_8251,N_8249);
nand U9707 (N_9707,N_8298,N_8457);
or U9708 (N_9708,N_8382,N_8451);
nor U9709 (N_9709,N_8723,N_8002);
nor U9710 (N_9710,N_8439,N_8568);
and U9711 (N_9711,N_8990,N_8891);
nor U9712 (N_9712,N_8375,N_8693);
nor U9713 (N_9713,N_8519,N_8866);
nor U9714 (N_9714,N_8325,N_8222);
nor U9715 (N_9715,N_8484,N_8245);
nand U9716 (N_9716,N_8952,N_8658);
nand U9717 (N_9717,N_8290,N_8695);
and U9718 (N_9718,N_8211,N_8820);
nand U9719 (N_9719,N_8643,N_8210);
nand U9720 (N_9720,N_8206,N_8892);
nand U9721 (N_9721,N_8413,N_8828);
and U9722 (N_9722,N_8713,N_8798);
nand U9723 (N_9723,N_8288,N_8054);
nand U9724 (N_9724,N_8863,N_8749);
or U9725 (N_9725,N_8481,N_8270);
nor U9726 (N_9726,N_8899,N_8411);
and U9727 (N_9727,N_8126,N_8506);
and U9728 (N_9728,N_8311,N_8079);
nand U9729 (N_9729,N_8079,N_8087);
and U9730 (N_9730,N_8345,N_8895);
nand U9731 (N_9731,N_8629,N_8329);
nor U9732 (N_9732,N_8425,N_8099);
and U9733 (N_9733,N_8502,N_8511);
or U9734 (N_9734,N_8966,N_8134);
or U9735 (N_9735,N_8970,N_8239);
nand U9736 (N_9736,N_8583,N_8910);
xor U9737 (N_9737,N_8889,N_8052);
or U9738 (N_9738,N_8727,N_8879);
and U9739 (N_9739,N_8284,N_8157);
nor U9740 (N_9740,N_8490,N_8268);
and U9741 (N_9741,N_8234,N_8971);
nor U9742 (N_9742,N_8328,N_8839);
and U9743 (N_9743,N_8094,N_8470);
and U9744 (N_9744,N_8166,N_8903);
nor U9745 (N_9745,N_8298,N_8721);
nand U9746 (N_9746,N_8224,N_8515);
nand U9747 (N_9747,N_8473,N_8364);
nand U9748 (N_9748,N_8701,N_8322);
nand U9749 (N_9749,N_8120,N_8858);
and U9750 (N_9750,N_8714,N_8407);
xor U9751 (N_9751,N_8064,N_8892);
or U9752 (N_9752,N_8774,N_8706);
nor U9753 (N_9753,N_8050,N_8484);
nand U9754 (N_9754,N_8639,N_8876);
or U9755 (N_9755,N_8337,N_8627);
or U9756 (N_9756,N_8615,N_8427);
and U9757 (N_9757,N_8564,N_8568);
xor U9758 (N_9758,N_8105,N_8134);
nor U9759 (N_9759,N_8198,N_8391);
nor U9760 (N_9760,N_8689,N_8584);
and U9761 (N_9761,N_8291,N_8415);
nand U9762 (N_9762,N_8299,N_8900);
nor U9763 (N_9763,N_8646,N_8328);
nand U9764 (N_9764,N_8149,N_8840);
and U9765 (N_9765,N_8782,N_8213);
nor U9766 (N_9766,N_8401,N_8322);
or U9767 (N_9767,N_8972,N_8584);
and U9768 (N_9768,N_8425,N_8667);
nand U9769 (N_9769,N_8500,N_8081);
or U9770 (N_9770,N_8907,N_8874);
xor U9771 (N_9771,N_8266,N_8267);
nand U9772 (N_9772,N_8913,N_8922);
nand U9773 (N_9773,N_8632,N_8346);
nor U9774 (N_9774,N_8240,N_8507);
xnor U9775 (N_9775,N_8962,N_8179);
nand U9776 (N_9776,N_8621,N_8325);
and U9777 (N_9777,N_8977,N_8103);
nand U9778 (N_9778,N_8991,N_8302);
nand U9779 (N_9779,N_8726,N_8801);
nor U9780 (N_9780,N_8873,N_8372);
nor U9781 (N_9781,N_8243,N_8738);
and U9782 (N_9782,N_8390,N_8418);
or U9783 (N_9783,N_8050,N_8582);
nand U9784 (N_9784,N_8792,N_8874);
nor U9785 (N_9785,N_8912,N_8132);
and U9786 (N_9786,N_8143,N_8818);
or U9787 (N_9787,N_8158,N_8917);
nand U9788 (N_9788,N_8808,N_8314);
nand U9789 (N_9789,N_8095,N_8314);
and U9790 (N_9790,N_8704,N_8364);
nor U9791 (N_9791,N_8244,N_8946);
nor U9792 (N_9792,N_8817,N_8276);
or U9793 (N_9793,N_8361,N_8870);
nand U9794 (N_9794,N_8040,N_8262);
nand U9795 (N_9795,N_8277,N_8462);
and U9796 (N_9796,N_8549,N_8550);
nand U9797 (N_9797,N_8792,N_8130);
nand U9798 (N_9798,N_8440,N_8097);
xnor U9799 (N_9799,N_8340,N_8182);
or U9800 (N_9800,N_8397,N_8254);
and U9801 (N_9801,N_8920,N_8184);
nor U9802 (N_9802,N_8342,N_8054);
or U9803 (N_9803,N_8553,N_8540);
nand U9804 (N_9804,N_8897,N_8374);
or U9805 (N_9805,N_8597,N_8192);
xnor U9806 (N_9806,N_8893,N_8404);
and U9807 (N_9807,N_8355,N_8122);
or U9808 (N_9808,N_8713,N_8124);
nand U9809 (N_9809,N_8126,N_8897);
or U9810 (N_9810,N_8080,N_8779);
nand U9811 (N_9811,N_8615,N_8145);
or U9812 (N_9812,N_8225,N_8364);
and U9813 (N_9813,N_8498,N_8156);
nor U9814 (N_9814,N_8466,N_8486);
or U9815 (N_9815,N_8003,N_8512);
nor U9816 (N_9816,N_8471,N_8702);
and U9817 (N_9817,N_8840,N_8435);
nand U9818 (N_9818,N_8108,N_8809);
and U9819 (N_9819,N_8267,N_8893);
xnor U9820 (N_9820,N_8381,N_8359);
nor U9821 (N_9821,N_8173,N_8097);
and U9822 (N_9822,N_8270,N_8998);
nor U9823 (N_9823,N_8522,N_8109);
nor U9824 (N_9824,N_8235,N_8015);
nand U9825 (N_9825,N_8443,N_8462);
nand U9826 (N_9826,N_8650,N_8068);
and U9827 (N_9827,N_8789,N_8753);
nor U9828 (N_9828,N_8071,N_8619);
nor U9829 (N_9829,N_8041,N_8878);
xnor U9830 (N_9830,N_8000,N_8819);
nor U9831 (N_9831,N_8838,N_8891);
xnor U9832 (N_9832,N_8402,N_8432);
nor U9833 (N_9833,N_8601,N_8980);
or U9834 (N_9834,N_8980,N_8042);
and U9835 (N_9835,N_8594,N_8670);
or U9836 (N_9836,N_8364,N_8222);
nor U9837 (N_9837,N_8634,N_8478);
or U9838 (N_9838,N_8735,N_8045);
xor U9839 (N_9839,N_8415,N_8558);
and U9840 (N_9840,N_8979,N_8573);
or U9841 (N_9841,N_8535,N_8753);
or U9842 (N_9842,N_8083,N_8285);
xor U9843 (N_9843,N_8295,N_8741);
or U9844 (N_9844,N_8730,N_8594);
and U9845 (N_9845,N_8740,N_8892);
nand U9846 (N_9846,N_8718,N_8473);
nor U9847 (N_9847,N_8555,N_8982);
nor U9848 (N_9848,N_8816,N_8648);
or U9849 (N_9849,N_8540,N_8921);
and U9850 (N_9850,N_8731,N_8840);
nor U9851 (N_9851,N_8111,N_8170);
nor U9852 (N_9852,N_8078,N_8613);
nand U9853 (N_9853,N_8040,N_8849);
and U9854 (N_9854,N_8892,N_8513);
nor U9855 (N_9855,N_8916,N_8628);
or U9856 (N_9856,N_8706,N_8185);
and U9857 (N_9857,N_8953,N_8905);
xor U9858 (N_9858,N_8293,N_8013);
or U9859 (N_9859,N_8571,N_8532);
and U9860 (N_9860,N_8141,N_8665);
nand U9861 (N_9861,N_8365,N_8606);
or U9862 (N_9862,N_8561,N_8805);
and U9863 (N_9863,N_8545,N_8111);
and U9864 (N_9864,N_8460,N_8459);
and U9865 (N_9865,N_8671,N_8795);
xor U9866 (N_9866,N_8998,N_8063);
or U9867 (N_9867,N_8487,N_8778);
and U9868 (N_9868,N_8597,N_8740);
and U9869 (N_9869,N_8770,N_8147);
nor U9870 (N_9870,N_8978,N_8870);
nor U9871 (N_9871,N_8136,N_8898);
nand U9872 (N_9872,N_8918,N_8575);
nand U9873 (N_9873,N_8935,N_8218);
nand U9874 (N_9874,N_8431,N_8820);
xnor U9875 (N_9875,N_8857,N_8938);
nand U9876 (N_9876,N_8274,N_8856);
or U9877 (N_9877,N_8570,N_8041);
nor U9878 (N_9878,N_8501,N_8452);
or U9879 (N_9879,N_8341,N_8349);
or U9880 (N_9880,N_8448,N_8767);
and U9881 (N_9881,N_8223,N_8585);
xnor U9882 (N_9882,N_8487,N_8428);
or U9883 (N_9883,N_8275,N_8004);
or U9884 (N_9884,N_8562,N_8029);
or U9885 (N_9885,N_8109,N_8066);
nand U9886 (N_9886,N_8088,N_8766);
or U9887 (N_9887,N_8399,N_8235);
nor U9888 (N_9888,N_8731,N_8949);
nand U9889 (N_9889,N_8346,N_8326);
nor U9890 (N_9890,N_8377,N_8469);
xnor U9891 (N_9891,N_8141,N_8976);
nor U9892 (N_9892,N_8804,N_8404);
nor U9893 (N_9893,N_8495,N_8977);
nor U9894 (N_9894,N_8682,N_8768);
xnor U9895 (N_9895,N_8722,N_8893);
and U9896 (N_9896,N_8867,N_8366);
and U9897 (N_9897,N_8683,N_8502);
nor U9898 (N_9898,N_8834,N_8116);
and U9899 (N_9899,N_8647,N_8560);
and U9900 (N_9900,N_8949,N_8226);
nor U9901 (N_9901,N_8115,N_8947);
or U9902 (N_9902,N_8427,N_8861);
and U9903 (N_9903,N_8910,N_8601);
nand U9904 (N_9904,N_8012,N_8961);
or U9905 (N_9905,N_8727,N_8648);
nand U9906 (N_9906,N_8341,N_8029);
and U9907 (N_9907,N_8926,N_8965);
or U9908 (N_9908,N_8050,N_8567);
or U9909 (N_9909,N_8857,N_8257);
or U9910 (N_9910,N_8985,N_8562);
nand U9911 (N_9911,N_8102,N_8604);
nor U9912 (N_9912,N_8375,N_8576);
nand U9913 (N_9913,N_8888,N_8719);
nor U9914 (N_9914,N_8695,N_8931);
nor U9915 (N_9915,N_8371,N_8066);
or U9916 (N_9916,N_8468,N_8601);
nor U9917 (N_9917,N_8707,N_8673);
and U9918 (N_9918,N_8438,N_8481);
nor U9919 (N_9919,N_8730,N_8589);
nand U9920 (N_9920,N_8742,N_8368);
nand U9921 (N_9921,N_8816,N_8036);
nand U9922 (N_9922,N_8123,N_8629);
nand U9923 (N_9923,N_8257,N_8797);
and U9924 (N_9924,N_8005,N_8543);
or U9925 (N_9925,N_8723,N_8226);
nand U9926 (N_9926,N_8880,N_8016);
nor U9927 (N_9927,N_8869,N_8405);
nand U9928 (N_9928,N_8046,N_8248);
or U9929 (N_9929,N_8722,N_8640);
or U9930 (N_9930,N_8911,N_8727);
nand U9931 (N_9931,N_8159,N_8256);
or U9932 (N_9932,N_8519,N_8403);
or U9933 (N_9933,N_8941,N_8511);
nor U9934 (N_9934,N_8837,N_8760);
or U9935 (N_9935,N_8086,N_8052);
or U9936 (N_9936,N_8122,N_8363);
or U9937 (N_9937,N_8343,N_8679);
or U9938 (N_9938,N_8591,N_8160);
nor U9939 (N_9939,N_8388,N_8029);
xor U9940 (N_9940,N_8948,N_8365);
nand U9941 (N_9941,N_8643,N_8496);
nand U9942 (N_9942,N_8270,N_8828);
or U9943 (N_9943,N_8320,N_8692);
nor U9944 (N_9944,N_8008,N_8887);
nor U9945 (N_9945,N_8057,N_8884);
nand U9946 (N_9946,N_8896,N_8541);
nand U9947 (N_9947,N_8278,N_8608);
nand U9948 (N_9948,N_8427,N_8657);
and U9949 (N_9949,N_8652,N_8492);
or U9950 (N_9950,N_8266,N_8387);
and U9951 (N_9951,N_8299,N_8215);
nand U9952 (N_9952,N_8515,N_8098);
nor U9953 (N_9953,N_8979,N_8681);
nand U9954 (N_9954,N_8078,N_8274);
xor U9955 (N_9955,N_8342,N_8989);
or U9956 (N_9956,N_8307,N_8254);
xor U9957 (N_9957,N_8952,N_8572);
and U9958 (N_9958,N_8195,N_8230);
nor U9959 (N_9959,N_8315,N_8235);
or U9960 (N_9960,N_8024,N_8501);
nand U9961 (N_9961,N_8835,N_8671);
nand U9962 (N_9962,N_8658,N_8295);
nor U9963 (N_9963,N_8330,N_8775);
and U9964 (N_9964,N_8520,N_8560);
nor U9965 (N_9965,N_8866,N_8040);
or U9966 (N_9966,N_8789,N_8122);
or U9967 (N_9967,N_8968,N_8919);
or U9968 (N_9968,N_8191,N_8967);
nand U9969 (N_9969,N_8308,N_8313);
or U9970 (N_9970,N_8236,N_8826);
nor U9971 (N_9971,N_8572,N_8789);
xor U9972 (N_9972,N_8535,N_8865);
xnor U9973 (N_9973,N_8211,N_8411);
and U9974 (N_9974,N_8449,N_8587);
or U9975 (N_9975,N_8493,N_8803);
xor U9976 (N_9976,N_8088,N_8876);
nor U9977 (N_9977,N_8493,N_8975);
and U9978 (N_9978,N_8802,N_8323);
and U9979 (N_9979,N_8131,N_8686);
and U9980 (N_9980,N_8258,N_8447);
and U9981 (N_9981,N_8400,N_8613);
or U9982 (N_9982,N_8348,N_8677);
and U9983 (N_9983,N_8916,N_8154);
or U9984 (N_9984,N_8844,N_8906);
nor U9985 (N_9985,N_8801,N_8943);
xnor U9986 (N_9986,N_8570,N_8162);
and U9987 (N_9987,N_8532,N_8547);
nand U9988 (N_9988,N_8686,N_8885);
or U9989 (N_9989,N_8956,N_8558);
nand U9990 (N_9990,N_8116,N_8012);
or U9991 (N_9991,N_8935,N_8743);
or U9992 (N_9992,N_8273,N_8741);
or U9993 (N_9993,N_8894,N_8437);
and U9994 (N_9994,N_8594,N_8304);
xor U9995 (N_9995,N_8854,N_8495);
or U9996 (N_9996,N_8568,N_8536);
nand U9997 (N_9997,N_8562,N_8156);
and U9998 (N_9998,N_8248,N_8436);
nor U9999 (N_9999,N_8591,N_8165);
and U10000 (N_10000,N_9649,N_9014);
nor U10001 (N_10001,N_9909,N_9538);
nor U10002 (N_10002,N_9494,N_9485);
nor U10003 (N_10003,N_9934,N_9498);
and U10004 (N_10004,N_9563,N_9639);
and U10005 (N_10005,N_9381,N_9711);
and U10006 (N_10006,N_9378,N_9841);
nor U10007 (N_10007,N_9020,N_9578);
or U10008 (N_10008,N_9113,N_9447);
nand U10009 (N_10009,N_9532,N_9663);
nand U10010 (N_10010,N_9998,N_9674);
nand U10011 (N_10011,N_9009,N_9181);
nand U10012 (N_10012,N_9268,N_9997);
or U10013 (N_10013,N_9428,N_9673);
nor U10014 (N_10014,N_9296,N_9005);
nand U10015 (N_10015,N_9486,N_9777);
nand U10016 (N_10016,N_9341,N_9408);
xor U10017 (N_10017,N_9662,N_9921);
nand U10018 (N_10018,N_9317,N_9753);
or U10019 (N_10019,N_9101,N_9714);
and U10020 (N_10020,N_9034,N_9374);
or U10021 (N_10021,N_9307,N_9470);
or U10022 (N_10022,N_9106,N_9624);
and U10023 (N_10023,N_9876,N_9877);
or U10024 (N_10024,N_9367,N_9806);
or U10025 (N_10025,N_9281,N_9242);
nand U10026 (N_10026,N_9245,N_9458);
and U10027 (N_10027,N_9868,N_9569);
and U10028 (N_10028,N_9069,N_9683);
nor U10029 (N_10029,N_9555,N_9985);
and U10030 (N_10030,N_9748,N_9346);
nand U10031 (N_10031,N_9339,N_9442);
or U10032 (N_10032,N_9475,N_9235);
nand U10033 (N_10033,N_9795,N_9140);
nor U10034 (N_10034,N_9298,N_9309);
nand U10035 (N_10035,N_9037,N_9954);
and U10036 (N_10036,N_9716,N_9501);
or U10037 (N_10037,N_9616,N_9200);
nand U10038 (N_10038,N_9659,N_9945);
nand U10039 (N_10039,N_9786,N_9450);
nand U10040 (N_10040,N_9459,N_9647);
or U10041 (N_10041,N_9646,N_9580);
nor U10042 (N_10042,N_9070,N_9903);
or U10043 (N_10043,N_9397,N_9404);
nand U10044 (N_10044,N_9276,N_9520);
or U10045 (N_10045,N_9991,N_9935);
and U10046 (N_10046,N_9093,N_9222);
or U10047 (N_10047,N_9204,N_9155);
or U10048 (N_10048,N_9967,N_9544);
or U10049 (N_10049,N_9180,N_9051);
or U10050 (N_10050,N_9696,N_9363);
and U10051 (N_10051,N_9349,N_9384);
nor U10052 (N_10052,N_9210,N_9084);
and U10053 (N_10053,N_9698,N_9418);
and U10054 (N_10054,N_9249,N_9358);
nand U10055 (N_10055,N_9875,N_9291);
nand U10056 (N_10056,N_9534,N_9267);
or U10057 (N_10057,N_9856,N_9852);
nand U10058 (N_10058,N_9133,N_9926);
xor U10059 (N_10059,N_9566,N_9496);
nand U10060 (N_10060,N_9816,N_9743);
nand U10061 (N_10061,N_9600,N_9894);
nor U10062 (N_10062,N_9526,N_9798);
and U10063 (N_10063,N_9148,N_9282);
nor U10064 (N_10064,N_9587,N_9247);
nand U10065 (N_10065,N_9482,N_9310);
xnor U10066 (N_10066,N_9817,N_9197);
nor U10067 (N_10067,N_9451,N_9509);
xnor U10068 (N_10068,N_9656,N_9900);
nand U10069 (N_10069,N_9278,N_9539);
nand U10070 (N_10070,N_9283,N_9059);
and U10071 (N_10071,N_9726,N_9541);
nor U10072 (N_10072,N_9957,N_9527);
nor U10073 (N_10073,N_9045,N_9433);
and U10074 (N_10074,N_9866,N_9170);
xnor U10075 (N_10075,N_9749,N_9046);
or U10076 (N_10076,N_9254,N_9831);
and U10077 (N_10077,N_9388,N_9734);
and U10078 (N_10078,N_9038,N_9585);
or U10079 (N_10079,N_9925,N_9444);
and U10080 (N_10080,N_9859,N_9350);
and U10081 (N_10081,N_9635,N_9620);
xnor U10082 (N_10082,N_9231,N_9375);
nand U10083 (N_10083,N_9599,N_9581);
nor U10084 (N_10084,N_9809,N_9007);
nor U10085 (N_10085,N_9636,N_9724);
nand U10086 (N_10086,N_9637,N_9631);
nor U10087 (N_10087,N_9577,N_9697);
nor U10088 (N_10088,N_9454,N_9503);
or U10089 (N_10089,N_9739,N_9685);
and U10090 (N_10090,N_9568,N_9941);
xnor U10091 (N_10091,N_9778,N_9386);
and U10092 (N_10092,N_9025,N_9571);
nor U10093 (N_10093,N_9011,N_9864);
and U10094 (N_10094,N_9978,N_9699);
or U10095 (N_10095,N_9125,N_9732);
nand U10096 (N_10096,N_9560,N_9744);
nand U10097 (N_10097,N_9071,N_9962);
and U10098 (N_10098,N_9615,N_9331);
or U10099 (N_10099,N_9187,N_9373);
and U10100 (N_10100,N_9729,N_9913);
xnor U10101 (N_10101,N_9361,N_9145);
or U10102 (N_10102,N_9193,N_9480);
and U10103 (N_10103,N_9337,N_9653);
nor U10104 (N_10104,N_9285,N_9015);
or U10105 (N_10105,N_9522,N_9703);
nor U10106 (N_10106,N_9948,N_9413);
and U10107 (N_10107,N_9471,N_9351);
nand U10108 (N_10108,N_9535,N_9460);
nor U10109 (N_10109,N_9003,N_9694);
nand U10110 (N_10110,N_9754,N_9314);
nand U10111 (N_10111,N_9944,N_9030);
or U10112 (N_10112,N_9968,N_9202);
and U10113 (N_10113,N_9583,N_9336);
nor U10114 (N_10114,N_9543,N_9862);
and U10115 (N_10115,N_9256,N_9255);
or U10116 (N_10116,N_9359,N_9312);
xor U10117 (N_10117,N_9320,N_9313);
nand U10118 (N_10118,N_9239,N_9040);
and U10119 (N_10119,N_9556,N_9820);
nand U10120 (N_10120,N_9474,N_9099);
nor U10121 (N_10121,N_9369,N_9623);
or U10122 (N_10122,N_9784,N_9243);
nand U10123 (N_10123,N_9722,N_9209);
nand U10124 (N_10124,N_9406,N_9700);
or U10125 (N_10125,N_9995,N_9452);
or U10126 (N_10126,N_9608,N_9244);
nor U10127 (N_10127,N_9865,N_9758);
nand U10128 (N_10128,N_9213,N_9299);
nand U10129 (N_10129,N_9063,N_9171);
or U10130 (N_10130,N_9780,N_9735);
nand U10131 (N_10131,N_9016,N_9504);
nand U10132 (N_10132,N_9969,N_9105);
nor U10133 (N_10133,N_9676,N_9379);
xnor U10134 (N_10134,N_9169,N_9114);
nand U10135 (N_10135,N_9372,N_9497);
nand U10136 (N_10136,N_9860,N_9545);
nand U10137 (N_10137,N_9727,N_9073);
nand U10138 (N_10138,N_9602,N_9770);
nor U10139 (N_10139,N_9690,N_9469);
nor U10140 (N_10140,N_9164,N_9253);
and U10141 (N_10141,N_9645,N_9746);
nor U10142 (N_10142,N_9064,N_9088);
or U10143 (N_10143,N_9211,N_9153);
nand U10144 (N_10144,N_9043,N_9248);
or U10145 (N_10145,N_9225,N_9082);
or U10146 (N_10146,N_9018,N_9672);
nor U10147 (N_10147,N_9787,N_9885);
or U10148 (N_10148,N_9939,N_9733);
xnor U10149 (N_10149,N_9455,N_9465);
or U10150 (N_10150,N_9146,N_9869);
xor U10151 (N_10151,N_9610,N_9707);
or U10152 (N_10152,N_9399,N_9912);
and U10153 (N_10153,N_9606,N_9223);
nor U10154 (N_10154,N_9110,N_9265);
xor U10155 (N_10155,N_9271,N_9915);
nand U10156 (N_10156,N_9149,N_9449);
nand U10157 (N_10157,N_9609,N_9670);
nand U10158 (N_10158,N_9290,N_9956);
nor U10159 (N_10159,N_9483,N_9713);
nand U10160 (N_10160,N_9429,N_9029);
and U10161 (N_10161,N_9226,N_9318);
nor U10162 (N_10162,N_9316,N_9490);
and U10163 (N_10163,N_9144,N_9546);
nor U10164 (N_10164,N_9232,N_9679);
or U10165 (N_10165,N_9742,N_9289);
xnor U10166 (N_10166,N_9523,N_9489);
nor U10167 (N_10167,N_9216,N_9717);
nor U10168 (N_10168,N_9371,N_9633);
nor U10169 (N_10169,N_9584,N_9705);
or U10170 (N_10170,N_9837,N_9757);
xor U10171 (N_10171,N_9184,N_9812);
xor U10172 (N_10172,N_9319,N_9022);
or U10173 (N_10173,N_9960,N_9120);
nand U10174 (N_10174,N_9619,N_9559);
or U10175 (N_10175,N_9500,N_9215);
nand U10176 (N_10176,N_9198,N_9785);
nand U10177 (N_10177,N_9557,N_9330);
and U10178 (N_10178,N_9078,N_9026);
nand U10179 (N_10179,N_9052,N_9905);
xor U10180 (N_10180,N_9075,N_9325);
nor U10181 (N_10181,N_9701,N_9807);
xor U10182 (N_10182,N_9661,N_9094);
xnor U10183 (N_10183,N_9838,N_9775);
nor U10184 (N_10184,N_9626,N_9230);
xnor U10185 (N_10185,N_9421,N_9463);
nand U10186 (N_10186,N_9828,N_9205);
nor U10187 (N_10187,N_9240,N_9179);
xor U10188 (N_10188,N_9783,N_9801);
nand U10189 (N_10189,N_9768,N_9334);
or U10190 (N_10190,N_9689,N_9370);
or U10191 (N_10191,N_9720,N_9136);
and U10192 (N_10192,N_9861,N_9259);
or U10193 (N_10193,N_9554,N_9329);
nor U10194 (N_10194,N_9053,N_9959);
nor U10195 (N_10195,N_9252,N_9439);
xnor U10196 (N_10196,N_9086,N_9321);
nand U10197 (N_10197,N_9443,N_9815);
xnor U10198 (N_10198,N_9827,N_9675);
or U10199 (N_10199,N_9992,N_9607);
nor U10200 (N_10200,N_9767,N_9512);
and U10201 (N_10201,N_9867,N_9111);
or U10202 (N_10202,N_9883,N_9929);
or U10203 (N_10203,N_9264,N_9547);
xnor U10204 (N_10204,N_9165,N_9275);
or U10205 (N_10205,N_9593,N_9061);
nor U10206 (N_10206,N_9127,N_9095);
nand U10207 (N_10207,N_9517,N_9871);
xor U10208 (N_10208,N_9918,N_9977);
nor U10209 (N_10209,N_9401,N_9049);
nor U10210 (N_10210,N_9010,N_9182);
and U10211 (N_10211,N_9924,N_9407);
nor U10212 (N_10212,N_9725,N_9999);
and U10213 (N_10213,N_9327,N_9983);
or U10214 (N_10214,N_9212,N_9551);
and U10215 (N_10215,N_9335,N_9006);
nand U10216 (N_10216,N_9352,N_9655);
and U10217 (N_10217,N_9402,N_9686);
nand U10218 (N_10218,N_9691,N_9591);
and U10219 (N_10219,N_9036,N_9952);
or U10220 (N_10220,N_9800,N_9715);
and U10221 (N_10221,N_9027,N_9972);
or U10222 (N_10222,N_9814,N_9760);
nand U10223 (N_10223,N_9143,N_9234);
nor U10224 (N_10224,N_9041,N_9565);
nand U10225 (N_10225,N_9261,N_9292);
nand U10226 (N_10226,N_9176,N_9332);
and U10227 (N_10227,N_9258,N_9074);
and U10228 (N_10228,N_9834,N_9262);
and U10229 (N_10229,N_9755,N_9355);
nor U10230 (N_10230,N_9076,N_9650);
or U10231 (N_10231,N_9295,N_9612);
nor U10232 (N_10232,N_9958,N_9024);
and U10233 (N_10233,N_9395,N_9263);
or U10234 (N_10234,N_9863,N_9048);
xor U10235 (N_10235,N_9906,N_9605);
nand U10236 (N_10236,N_9927,N_9774);
nor U10237 (N_10237,N_9853,N_9680);
or U10238 (N_10238,N_9423,N_9789);
or U10239 (N_10239,N_9842,N_9246);
xor U10240 (N_10240,N_9525,N_9564);
nor U10241 (N_10241,N_9196,N_9481);
and U10242 (N_10242,N_9409,N_9658);
nor U10243 (N_10243,N_9540,N_9207);
nand U10244 (N_10244,N_9124,N_9682);
nand U10245 (N_10245,N_9550,N_9324);
nor U10246 (N_10246,N_9158,N_9529);
and U10247 (N_10247,N_9160,N_9928);
xnor U10248 (N_10248,N_9652,N_9634);
nand U10249 (N_10249,N_9139,N_9797);
or U10250 (N_10250,N_9129,N_9478);
nand U10251 (N_10251,N_9810,N_9955);
nand U10252 (N_10252,N_9096,N_9708);
nor U10253 (N_10253,N_9803,N_9062);
nor U10254 (N_10254,N_9943,N_9946);
or U10255 (N_10255,N_9847,N_9966);
nand U10256 (N_10256,N_9514,N_9986);
nand U10257 (N_10257,N_9695,N_9488);
nor U10258 (N_10258,N_9229,N_9897);
and U10259 (N_10259,N_9322,N_9294);
and U10260 (N_10260,N_9651,N_9622);
nand U10261 (N_10261,N_9723,N_9161);
nor U10262 (N_10262,N_9621,N_9328);
nor U10263 (N_10263,N_9185,N_9681);
nor U10264 (N_10264,N_9982,N_9843);
nor U10265 (N_10265,N_9942,N_9241);
and U10266 (N_10266,N_9441,N_9042);
nand U10267 (N_10267,N_9548,N_9391);
nand U10268 (N_10268,N_9138,N_9510);
or U10269 (N_10269,N_9425,N_9542);
xnor U10270 (N_10270,N_9519,N_9792);
or U10271 (N_10271,N_9702,N_9417);
nand U10272 (N_10272,N_9109,N_9175);
xor U10273 (N_10273,N_9440,N_9368);
nor U10274 (N_10274,N_9385,N_9846);
nand U10275 (N_10275,N_9854,N_9870);
and U10276 (N_10276,N_9889,N_9080);
nor U10277 (N_10277,N_9219,N_9008);
and U10278 (N_10278,N_9751,N_9394);
or U10279 (N_10279,N_9886,N_9762);
or U10280 (N_10280,N_9830,N_9832);
nor U10281 (N_10281,N_9154,N_9100);
or U10282 (N_10282,N_9936,N_9426);
and U10283 (N_10283,N_9277,N_9811);
or U10284 (N_10284,N_9376,N_9031);
nand U10285 (N_10285,N_9567,N_9224);
nor U10286 (N_10286,N_9892,N_9311);
or U10287 (N_10287,N_9984,N_9805);
nand U10288 (N_10288,N_9993,N_9306);
nor U10289 (N_10289,N_9947,N_9582);
nand U10290 (N_10290,N_9588,N_9911);
nor U10291 (N_10291,N_9415,N_9638);
and U10292 (N_10292,N_9666,N_9899);
and U10293 (N_10293,N_9173,N_9613);
or U10294 (N_10294,N_9849,N_9383);
and U10295 (N_10295,N_9044,N_9269);
nand U10296 (N_10296,N_9004,N_9422);
nand U10297 (N_10297,N_9528,N_9765);
xnor U10298 (N_10298,N_9177,N_9186);
nand U10299 (N_10299,N_9938,N_9719);
nand U10300 (N_10300,N_9630,N_9116);
and U10301 (N_10301,N_9836,N_9839);
nor U10302 (N_10302,N_9393,N_9464);
and U10303 (N_10303,N_9736,N_9756);
nor U10304 (N_10304,N_9192,N_9472);
nor U10305 (N_10305,N_9437,N_9898);
or U10306 (N_10306,N_9880,N_9688);
nand U10307 (N_10307,N_9097,N_9507);
or U10308 (N_10308,N_9971,N_9887);
nand U10309 (N_10309,N_9844,N_9973);
or U10310 (N_10310,N_9590,N_9692);
nand U10311 (N_10311,N_9597,N_9360);
or U10312 (N_10312,N_9799,N_9601);
and U10313 (N_10313,N_9380,N_9087);
nor U10314 (N_10314,N_9141,N_9562);
nor U10315 (N_10315,N_9553,N_9572);
nor U10316 (N_10316,N_9183,N_9001);
nand U10317 (N_10317,N_9137,N_9364);
nor U10318 (N_10318,N_9028,N_9965);
nor U10319 (N_10319,N_9466,N_9901);
nor U10320 (N_10320,N_9305,N_9669);
and U10321 (N_10321,N_9824,N_9989);
nor U10322 (N_10322,N_9737,N_9521);
nor U10323 (N_10323,N_9115,N_9665);
nor U10324 (N_10324,N_9931,N_9611);
nand U10325 (N_10325,N_9194,N_9996);
and U10326 (N_10326,N_9343,N_9840);
nand U10327 (N_10327,N_9301,N_9818);
and U10328 (N_10328,N_9122,N_9769);
or U10329 (N_10329,N_9079,N_9410);
nand U10330 (N_10330,N_9808,N_9297);
or U10331 (N_10331,N_9802,N_9627);
nor U10332 (N_10332,N_9804,N_9881);
or U10333 (N_10333,N_9628,N_9435);
xor U10334 (N_10334,N_9595,N_9704);
or U10335 (N_10335,N_9220,N_9576);
nor U10336 (N_10336,N_9315,N_9083);
and U10337 (N_10337,N_9467,N_9858);
nand U10338 (N_10338,N_9427,N_9000);
or U10339 (N_10339,N_9974,N_9108);
nor U10340 (N_10340,N_9150,N_9531);
nor U10341 (N_10341,N_9250,N_9130);
and U10342 (N_10342,N_9895,N_9491);
and U10343 (N_10343,N_9416,N_9142);
nand U10344 (N_10344,N_9032,N_9208);
nand U10345 (N_10345,N_9499,N_9398);
nand U10346 (N_10346,N_9089,N_9648);
nand U10347 (N_10347,N_9077,N_9412);
or U10348 (N_10348,N_9436,N_9468);
or U10349 (N_10349,N_9304,N_9845);
nor U10350 (N_10350,N_9980,N_9949);
nand U10351 (N_10351,N_9752,N_9251);
or U10352 (N_10352,N_9874,N_9477);
nor U10353 (N_10353,N_9121,N_9922);
xor U10354 (N_10354,N_9825,N_9937);
xnor U10355 (N_10355,N_9102,N_9047);
and U10356 (N_10356,N_9618,N_9790);
nor U10357 (N_10357,N_9163,N_9023);
nor U10358 (N_10358,N_9994,N_9709);
nor U10359 (N_10359,N_9614,N_9493);
or U10360 (N_10360,N_9405,N_9904);
nor U10361 (N_10361,N_9134,N_9850);
and U10362 (N_10362,N_9473,N_9396);
or U10363 (N_10363,N_9759,N_9288);
or U10364 (N_10364,N_9293,N_9345);
nor U10365 (N_10365,N_9910,N_9821);
and U10366 (N_10366,N_9432,N_9090);
or U10367 (N_10367,N_9730,N_9448);
nor U10368 (N_10368,N_9855,N_9660);
nor U10369 (N_10369,N_9050,N_9594);
or U10370 (N_10370,N_9495,N_9103);
nor U10371 (N_10371,N_9156,N_9642);
or U10372 (N_10372,N_9446,N_9453);
and U10373 (N_10373,N_9747,N_9530);
and U10374 (N_10374,N_9505,N_9728);
xor U10375 (N_10375,N_9596,N_9017);
nand U10376 (N_10376,N_9081,N_9888);
xor U10377 (N_10377,N_9951,N_9411);
or U10378 (N_10378,N_9629,N_9930);
and U10379 (N_10379,N_9644,N_9056);
and U10380 (N_10380,N_9738,N_9377);
or U10381 (N_10381,N_9772,N_9366);
xor U10382 (N_10382,N_9424,N_9286);
or U10383 (N_10383,N_9990,N_9731);
and U10384 (N_10384,N_9533,N_9168);
or U10385 (N_10385,N_9833,N_9420);
nor U10386 (N_10386,N_9552,N_9776);
or U10387 (N_10387,N_9794,N_9178);
nor U10388 (N_10388,N_9641,N_9513);
and U10389 (N_10389,N_9012,N_9826);
nand U10390 (N_10390,N_9745,N_9851);
xor U10391 (N_10391,N_9592,N_9461);
and U10392 (N_10392,N_9604,N_9492);
xor U10393 (N_10393,N_9643,N_9893);
or U10394 (N_10394,N_9354,N_9940);
nand U10395 (N_10395,N_9438,N_9782);
or U10396 (N_10396,N_9693,N_9456);
nand U10397 (N_10397,N_9908,N_9228);
or U10398 (N_10398,N_9272,N_9147);
nor U10399 (N_10399,N_9484,N_9033);
xor U10400 (N_10400,N_9055,N_9233);
and U10401 (N_10401,N_9002,N_9195);
nor U10402 (N_10402,N_9326,N_9085);
or U10403 (N_10403,N_9353,N_9781);
and U10404 (N_10404,N_9356,N_9896);
and U10405 (N_10405,N_9218,N_9279);
xnor U10406 (N_10406,N_9933,N_9667);
or U10407 (N_10407,N_9067,N_9891);
nor U10408 (N_10408,N_9970,N_9479);
and U10409 (N_10409,N_9511,N_9217);
and U10410 (N_10410,N_9257,N_9640);
nor U10411 (N_10411,N_9159,N_9549);
or U10412 (N_10412,N_9287,N_9403);
and U10413 (N_10413,N_9431,N_9835);
nor U10414 (N_10414,N_9829,N_9502);
or U10415 (N_10415,N_9333,N_9128);
nor U10416 (N_10416,N_9706,N_9953);
nand U10417 (N_10417,N_9221,N_9166);
nand U10418 (N_10418,N_9671,N_9365);
or U10419 (N_10419,N_9348,N_9579);
or U10420 (N_10420,N_9457,N_9389);
or U10421 (N_10421,N_9362,N_9524);
nor U10422 (N_10422,N_9092,N_9057);
or U10423 (N_10423,N_9347,N_9603);
and U10424 (N_10424,N_9761,N_9162);
or U10425 (N_10425,N_9126,N_9152);
nand U10426 (N_10426,N_9981,N_9112);
nor U10427 (N_10427,N_9791,N_9961);
nor U10428 (N_10428,N_9575,N_9589);
nor U10429 (N_10429,N_9677,N_9151);
xor U10430 (N_10430,N_9764,N_9203);
and U10431 (N_10431,N_9266,N_9878);
xnor U10432 (N_10432,N_9506,N_9664);
or U10433 (N_10433,N_9199,N_9174);
or U10434 (N_10434,N_9382,N_9274);
nor U10435 (N_10435,N_9238,N_9302);
nor U10436 (N_10436,N_9561,N_9054);
or U10437 (N_10437,N_9167,N_9920);
or U10438 (N_10438,N_9773,N_9058);
nor U10439 (N_10439,N_9654,N_9766);
nand U10440 (N_10440,N_9260,N_9979);
nand U10441 (N_10441,N_9214,N_9917);
xnor U10442 (N_10442,N_9668,N_9872);
or U10443 (N_10443,N_9068,N_9098);
xnor U10444 (N_10444,N_9950,N_9632);
xor U10445 (N_10445,N_9932,N_9476);
nor U10446 (N_10446,N_9771,N_9964);
nor U10447 (N_10447,N_9763,N_9976);
or U10448 (N_10448,N_9191,N_9570);
or U10449 (N_10449,N_9338,N_9060);
xor U10450 (N_10450,N_9021,N_9387);
and U10451 (N_10451,N_9013,N_9188);
nor U10452 (N_10452,N_9975,N_9848);
nand U10453 (N_10453,N_9857,N_9104);
and U10454 (N_10454,N_9132,N_9687);
or U10455 (N_10455,N_9712,N_9157);
nor U10456 (N_10456,N_9284,N_9118);
nand U10457 (N_10457,N_9072,N_9573);
nor U10458 (N_10458,N_9135,N_9066);
nand U10459 (N_10459,N_9172,N_9823);
nor U10460 (N_10460,N_9879,N_9574);
or U10461 (N_10461,N_9323,N_9201);
nor U10462 (N_10462,N_9131,N_9019);
or U10463 (N_10463,N_9430,N_9657);
xor U10464 (N_10464,N_9237,N_9419);
xor U10465 (N_10465,N_9390,N_9123);
and U10466 (N_10466,N_9819,N_9039);
and U10467 (N_10467,N_9508,N_9035);
or U10468 (N_10468,N_9678,N_9537);
nor U10469 (N_10469,N_9392,N_9788);
or U10470 (N_10470,N_9344,N_9625);
nor U10471 (N_10471,N_9718,N_9796);
nor U10472 (N_10472,N_9740,N_9434);
nand U10473 (N_10473,N_9914,N_9303);
nand U10474 (N_10474,N_9923,N_9190);
and U10475 (N_10475,N_9236,N_9750);
and U10476 (N_10476,N_9963,N_9270);
and U10477 (N_10477,N_9987,N_9882);
nand U10478 (N_10478,N_9300,N_9890);
or U10479 (N_10479,N_9907,N_9721);
and U10480 (N_10480,N_9516,N_9988);
nor U10481 (N_10481,N_9357,N_9598);
nand U10482 (N_10482,N_9308,N_9117);
nand U10483 (N_10483,N_9779,N_9916);
and U10484 (N_10484,N_9487,N_9884);
nand U10485 (N_10485,N_9065,N_9873);
or U10486 (N_10486,N_9902,N_9189);
and U10487 (N_10487,N_9119,N_9227);
nor U10488 (N_10488,N_9515,N_9462);
nand U10489 (N_10489,N_9280,N_9586);
and U10490 (N_10490,N_9813,N_9684);
xnor U10491 (N_10491,N_9414,N_9536);
and U10492 (N_10492,N_9340,N_9400);
nand U10493 (N_10493,N_9710,N_9558);
nand U10494 (N_10494,N_9822,N_9445);
nand U10495 (N_10495,N_9919,N_9617);
nor U10496 (N_10496,N_9107,N_9206);
and U10497 (N_10497,N_9793,N_9741);
nand U10498 (N_10498,N_9273,N_9342);
nor U10499 (N_10499,N_9518,N_9091);
nor U10500 (N_10500,N_9847,N_9414);
or U10501 (N_10501,N_9979,N_9675);
nand U10502 (N_10502,N_9888,N_9322);
or U10503 (N_10503,N_9737,N_9018);
nor U10504 (N_10504,N_9204,N_9635);
and U10505 (N_10505,N_9430,N_9832);
or U10506 (N_10506,N_9657,N_9251);
and U10507 (N_10507,N_9666,N_9589);
nand U10508 (N_10508,N_9718,N_9897);
or U10509 (N_10509,N_9096,N_9638);
or U10510 (N_10510,N_9584,N_9956);
and U10511 (N_10511,N_9560,N_9344);
nor U10512 (N_10512,N_9282,N_9856);
nand U10513 (N_10513,N_9070,N_9909);
and U10514 (N_10514,N_9598,N_9786);
and U10515 (N_10515,N_9609,N_9902);
or U10516 (N_10516,N_9624,N_9319);
nor U10517 (N_10517,N_9752,N_9609);
and U10518 (N_10518,N_9245,N_9015);
nand U10519 (N_10519,N_9124,N_9129);
nand U10520 (N_10520,N_9730,N_9244);
nand U10521 (N_10521,N_9413,N_9229);
xnor U10522 (N_10522,N_9175,N_9816);
nand U10523 (N_10523,N_9956,N_9452);
or U10524 (N_10524,N_9187,N_9634);
nand U10525 (N_10525,N_9893,N_9651);
nor U10526 (N_10526,N_9575,N_9935);
xnor U10527 (N_10527,N_9783,N_9150);
and U10528 (N_10528,N_9904,N_9004);
or U10529 (N_10529,N_9350,N_9207);
and U10530 (N_10530,N_9444,N_9478);
and U10531 (N_10531,N_9336,N_9052);
nor U10532 (N_10532,N_9158,N_9930);
and U10533 (N_10533,N_9064,N_9042);
or U10534 (N_10534,N_9350,N_9485);
or U10535 (N_10535,N_9570,N_9513);
and U10536 (N_10536,N_9879,N_9820);
nand U10537 (N_10537,N_9656,N_9808);
nand U10538 (N_10538,N_9887,N_9275);
nand U10539 (N_10539,N_9825,N_9061);
xor U10540 (N_10540,N_9198,N_9750);
nor U10541 (N_10541,N_9830,N_9172);
nand U10542 (N_10542,N_9099,N_9135);
and U10543 (N_10543,N_9237,N_9378);
nand U10544 (N_10544,N_9296,N_9601);
nand U10545 (N_10545,N_9236,N_9880);
or U10546 (N_10546,N_9081,N_9569);
or U10547 (N_10547,N_9945,N_9075);
and U10548 (N_10548,N_9453,N_9217);
and U10549 (N_10549,N_9004,N_9826);
and U10550 (N_10550,N_9852,N_9717);
or U10551 (N_10551,N_9815,N_9113);
or U10552 (N_10552,N_9299,N_9079);
and U10553 (N_10553,N_9848,N_9850);
nand U10554 (N_10554,N_9962,N_9425);
or U10555 (N_10555,N_9757,N_9323);
and U10556 (N_10556,N_9422,N_9270);
and U10557 (N_10557,N_9790,N_9920);
nor U10558 (N_10558,N_9126,N_9399);
or U10559 (N_10559,N_9523,N_9648);
or U10560 (N_10560,N_9249,N_9322);
or U10561 (N_10561,N_9530,N_9717);
nand U10562 (N_10562,N_9737,N_9854);
or U10563 (N_10563,N_9965,N_9356);
or U10564 (N_10564,N_9937,N_9820);
nand U10565 (N_10565,N_9279,N_9358);
nand U10566 (N_10566,N_9688,N_9329);
and U10567 (N_10567,N_9771,N_9445);
nor U10568 (N_10568,N_9169,N_9401);
nor U10569 (N_10569,N_9341,N_9332);
and U10570 (N_10570,N_9982,N_9176);
nand U10571 (N_10571,N_9484,N_9739);
and U10572 (N_10572,N_9111,N_9460);
and U10573 (N_10573,N_9459,N_9000);
nor U10574 (N_10574,N_9615,N_9786);
or U10575 (N_10575,N_9015,N_9194);
nand U10576 (N_10576,N_9933,N_9186);
and U10577 (N_10577,N_9091,N_9319);
nor U10578 (N_10578,N_9526,N_9846);
nand U10579 (N_10579,N_9751,N_9670);
xor U10580 (N_10580,N_9743,N_9631);
nor U10581 (N_10581,N_9086,N_9079);
nor U10582 (N_10582,N_9177,N_9922);
or U10583 (N_10583,N_9169,N_9554);
and U10584 (N_10584,N_9024,N_9496);
nor U10585 (N_10585,N_9577,N_9188);
nor U10586 (N_10586,N_9397,N_9839);
and U10587 (N_10587,N_9543,N_9423);
nor U10588 (N_10588,N_9536,N_9212);
or U10589 (N_10589,N_9351,N_9529);
or U10590 (N_10590,N_9858,N_9501);
nor U10591 (N_10591,N_9040,N_9306);
nand U10592 (N_10592,N_9590,N_9659);
or U10593 (N_10593,N_9016,N_9971);
xor U10594 (N_10594,N_9272,N_9774);
and U10595 (N_10595,N_9832,N_9696);
xor U10596 (N_10596,N_9288,N_9597);
nand U10597 (N_10597,N_9232,N_9450);
or U10598 (N_10598,N_9887,N_9157);
and U10599 (N_10599,N_9603,N_9856);
and U10600 (N_10600,N_9065,N_9281);
or U10601 (N_10601,N_9621,N_9354);
nor U10602 (N_10602,N_9994,N_9265);
xor U10603 (N_10603,N_9619,N_9773);
nand U10604 (N_10604,N_9511,N_9926);
nor U10605 (N_10605,N_9778,N_9043);
and U10606 (N_10606,N_9792,N_9836);
nor U10607 (N_10607,N_9032,N_9005);
nand U10608 (N_10608,N_9949,N_9379);
nand U10609 (N_10609,N_9991,N_9531);
nor U10610 (N_10610,N_9097,N_9856);
and U10611 (N_10611,N_9674,N_9913);
nand U10612 (N_10612,N_9087,N_9164);
nand U10613 (N_10613,N_9169,N_9012);
or U10614 (N_10614,N_9859,N_9450);
or U10615 (N_10615,N_9569,N_9969);
nand U10616 (N_10616,N_9029,N_9278);
xor U10617 (N_10617,N_9025,N_9976);
xor U10618 (N_10618,N_9398,N_9551);
or U10619 (N_10619,N_9019,N_9490);
nand U10620 (N_10620,N_9988,N_9396);
xor U10621 (N_10621,N_9819,N_9779);
or U10622 (N_10622,N_9352,N_9252);
or U10623 (N_10623,N_9888,N_9449);
nor U10624 (N_10624,N_9768,N_9184);
and U10625 (N_10625,N_9811,N_9470);
and U10626 (N_10626,N_9895,N_9561);
nand U10627 (N_10627,N_9533,N_9284);
nor U10628 (N_10628,N_9529,N_9645);
nor U10629 (N_10629,N_9399,N_9667);
and U10630 (N_10630,N_9666,N_9430);
or U10631 (N_10631,N_9990,N_9170);
nor U10632 (N_10632,N_9049,N_9505);
nor U10633 (N_10633,N_9343,N_9114);
and U10634 (N_10634,N_9969,N_9076);
xor U10635 (N_10635,N_9029,N_9381);
nand U10636 (N_10636,N_9522,N_9788);
or U10637 (N_10637,N_9520,N_9769);
nor U10638 (N_10638,N_9800,N_9378);
xnor U10639 (N_10639,N_9155,N_9038);
xor U10640 (N_10640,N_9864,N_9120);
and U10641 (N_10641,N_9143,N_9885);
nand U10642 (N_10642,N_9052,N_9642);
nand U10643 (N_10643,N_9522,N_9980);
nand U10644 (N_10644,N_9430,N_9715);
and U10645 (N_10645,N_9882,N_9572);
and U10646 (N_10646,N_9666,N_9002);
and U10647 (N_10647,N_9281,N_9248);
xnor U10648 (N_10648,N_9252,N_9317);
nand U10649 (N_10649,N_9422,N_9773);
nor U10650 (N_10650,N_9344,N_9733);
and U10651 (N_10651,N_9432,N_9844);
nor U10652 (N_10652,N_9093,N_9015);
and U10653 (N_10653,N_9649,N_9042);
xor U10654 (N_10654,N_9623,N_9024);
or U10655 (N_10655,N_9112,N_9631);
nor U10656 (N_10656,N_9476,N_9709);
nor U10657 (N_10657,N_9370,N_9259);
nand U10658 (N_10658,N_9209,N_9846);
nor U10659 (N_10659,N_9229,N_9377);
or U10660 (N_10660,N_9136,N_9265);
and U10661 (N_10661,N_9732,N_9591);
nand U10662 (N_10662,N_9473,N_9597);
xnor U10663 (N_10663,N_9808,N_9956);
nand U10664 (N_10664,N_9226,N_9645);
nor U10665 (N_10665,N_9573,N_9901);
nand U10666 (N_10666,N_9848,N_9188);
or U10667 (N_10667,N_9604,N_9608);
nand U10668 (N_10668,N_9731,N_9695);
nand U10669 (N_10669,N_9262,N_9290);
or U10670 (N_10670,N_9711,N_9960);
and U10671 (N_10671,N_9792,N_9966);
and U10672 (N_10672,N_9818,N_9692);
xnor U10673 (N_10673,N_9927,N_9072);
nor U10674 (N_10674,N_9671,N_9080);
nor U10675 (N_10675,N_9795,N_9463);
or U10676 (N_10676,N_9650,N_9791);
or U10677 (N_10677,N_9481,N_9230);
or U10678 (N_10678,N_9139,N_9028);
and U10679 (N_10679,N_9677,N_9011);
or U10680 (N_10680,N_9166,N_9061);
xnor U10681 (N_10681,N_9978,N_9416);
nand U10682 (N_10682,N_9215,N_9217);
and U10683 (N_10683,N_9178,N_9428);
and U10684 (N_10684,N_9857,N_9849);
and U10685 (N_10685,N_9602,N_9267);
and U10686 (N_10686,N_9857,N_9379);
or U10687 (N_10687,N_9442,N_9208);
nand U10688 (N_10688,N_9867,N_9727);
xnor U10689 (N_10689,N_9057,N_9566);
and U10690 (N_10690,N_9584,N_9293);
and U10691 (N_10691,N_9592,N_9300);
or U10692 (N_10692,N_9154,N_9388);
and U10693 (N_10693,N_9785,N_9810);
nor U10694 (N_10694,N_9590,N_9172);
and U10695 (N_10695,N_9835,N_9998);
or U10696 (N_10696,N_9831,N_9150);
nor U10697 (N_10697,N_9772,N_9559);
nand U10698 (N_10698,N_9262,N_9629);
nor U10699 (N_10699,N_9055,N_9157);
nand U10700 (N_10700,N_9666,N_9266);
and U10701 (N_10701,N_9326,N_9458);
nand U10702 (N_10702,N_9411,N_9237);
and U10703 (N_10703,N_9686,N_9404);
and U10704 (N_10704,N_9697,N_9320);
nand U10705 (N_10705,N_9441,N_9865);
nor U10706 (N_10706,N_9347,N_9039);
or U10707 (N_10707,N_9026,N_9105);
nor U10708 (N_10708,N_9526,N_9383);
nor U10709 (N_10709,N_9646,N_9388);
or U10710 (N_10710,N_9370,N_9252);
or U10711 (N_10711,N_9449,N_9257);
nor U10712 (N_10712,N_9599,N_9196);
xor U10713 (N_10713,N_9011,N_9984);
or U10714 (N_10714,N_9762,N_9304);
and U10715 (N_10715,N_9239,N_9877);
xor U10716 (N_10716,N_9080,N_9844);
and U10717 (N_10717,N_9072,N_9374);
nor U10718 (N_10718,N_9279,N_9471);
or U10719 (N_10719,N_9391,N_9912);
nand U10720 (N_10720,N_9983,N_9244);
nand U10721 (N_10721,N_9051,N_9434);
xor U10722 (N_10722,N_9385,N_9029);
or U10723 (N_10723,N_9274,N_9612);
and U10724 (N_10724,N_9958,N_9453);
nor U10725 (N_10725,N_9658,N_9914);
nand U10726 (N_10726,N_9747,N_9948);
or U10727 (N_10727,N_9094,N_9902);
nand U10728 (N_10728,N_9539,N_9542);
and U10729 (N_10729,N_9778,N_9724);
or U10730 (N_10730,N_9763,N_9156);
and U10731 (N_10731,N_9928,N_9686);
or U10732 (N_10732,N_9111,N_9284);
nand U10733 (N_10733,N_9255,N_9396);
nor U10734 (N_10734,N_9781,N_9568);
and U10735 (N_10735,N_9465,N_9961);
nand U10736 (N_10736,N_9695,N_9739);
nand U10737 (N_10737,N_9937,N_9562);
and U10738 (N_10738,N_9963,N_9889);
or U10739 (N_10739,N_9199,N_9902);
nor U10740 (N_10740,N_9041,N_9140);
nand U10741 (N_10741,N_9352,N_9371);
and U10742 (N_10742,N_9922,N_9938);
or U10743 (N_10743,N_9052,N_9329);
and U10744 (N_10744,N_9039,N_9895);
nor U10745 (N_10745,N_9792,N_9638);
xor U10746 (N_10746,N_9951,N_9812);
nor U10747 (N_10747,N_9137,N_9330);
nor U10748 (N_10748,N_9629,N_9257);
xor U10749 (N_10749,N_9515,N_9987);
and U10750 (N_10750,N_9614,N_9796);
nor U10751 (N_10751,N_9245,N_9294);
xnor U10752 (N_10752,N_9207,N_9566);
nand U10753 (N_10753,N_9404,N_9619);
xnor U10754 (N_10754,N_9593,N_9291);
nand U10755 (N_10755,N_9032,N_9613);
and U10756 (N_10756,N_9589,N_9379);
or U10757 (N_10757,N_9439,N_9115);
or U10758 (N_10758,N_9776,N_9753);
and U10759 (N_10759,N_9805,N_9236);
and U10760 (N_10760,N_9570,N_9995);
nand U10761 (N_10761,N_9849,N_9725);
or U10762 (N_10762,N_9818,N_9495);
or U10763 (N_10763,N_9567,N_9705);
xor U10764 (N_10764,N_9402,N_9532);
or U10765 (N_10765,N_9001,N_9122);
or U10766 (N_10766,N_9061,N_9094);
nand U10767 (N_10767,N_9529,N_9572);
or U10768 (N_10768,N_9208,N_9884);
nor U10769 (N_10769,N_9296,N_9288);
or U10770 (N_10770,N_9128,N_9279);
nand U10771 (N_10771,N_9293,N_9499);
nand U10772 (N_10772,N_9252,N_9886);
or U10773 (N_10773,N_9641,N_9956);
or U10774 (N_10774,N_9932,N_9767);
nor U10775 (N_10775,N_9992,N_9061);
nor U10776 (N_10776,N_9042,N_9873);
nor U10777 (N_10777,N_9480,N_9121);
xnor U10778 (N_10778,N_9164,N_9982);
nand U10779 (N_10779,N_9708,N_9693);
nand U10780 (N_10780,N_9075,N_9390);
and U10781 (N_10781,N_9931,N_9232);
nor U10782 (N_10782,N_9628,N_9881);
or U10783 (N_10783,N_9002,N_9180);
and U10784 (N_10784,N_9127,N_9819);
nor U10785 (N_10785,N_9654,N_9635);
xnor U10786 (N_10786,N_9117,N_9968);
or U10787 (N_10787,N_9202,N_9389);
nand U10788 (N_10788,N_9923,N_9527);
nand U10789 (N_10789,N_9738,N_9000);
xnor U10790 (N_10790,N_9503,N_9191);
nor U10791 (N_10791,N_9909,N_9311);
nand U10792 (N_10792,N_9184,N_9487);
nor U10793 (N_10793,N_9950,N_9716);
and U10794 (N_10794,N_9509,N_9457);
or U10795 (N_10795,N_9011,N_9711);
nor U10796 (N_10796,N_9638,N_9100);
xor U10797 (N_10797,N_9072,N_9172);
and U10798 (N_10798,N_9973,N_9359);
nand U10799 (N_10799,N_9389,N_9608);
and U10800 (N_10800,N_9231,N_9123);
or U10801 (N_10801,N_9094,N_9277);
or U10802 (N_10802,N_9924,N_9442);
or U10803 (N_10803,N_9512,N_9069);
nor U10804 (N_10804,N_9077,N_9966);
or U10805 (N_10805,N_9345,N_9889);
nor U10806 (N_10806,N_9212,N_9929);
or U10807 (N_10807,N_9864,N_9087);
or U10808 (N_10808,N_9211,N_9509);
xor U10809 (N_10809,N_9884,N_9101);
or U10810 (N_10810,N_9794,N_9710);
nand U10811 (N_10811,N_9209,N_9001);
xor U10812 (N_10812,N_9903,N_9475);
or U10813 (N_10813,N_9531,N_9253);
or U10814 (N_10814,N_9571,N_9695);
and U10815 (N_10815,N_9844,N_9366);
nor U10816 (N_10816,N_9451,N_9239);
and U10817 (N_10817,N_9609,N_9807);
and U10818 (N_10818,N_9390,N_9485);
and U10819 (N_10819,N_9535,N_9866);
and U10820 (N_10820,N_9225,N_9227);
nand U10821 (N_10821,N_9248,N_9594);
or U10822 (N_10822,N_9418,N_9927);
nand U10823 (N_10823,N_9927,N_9795);
nand U10824 (N_10824,N_9054,N_9379);
nand U10825 (N_10825,N_9200,N_9031);
or U10826 (N_10826,N_9162,N_9913);
nor U10827 (N_10827,N_9234,N_9954);
nor U10828 (N_10828,N_9601,N_9260);
and U10829 (N_10829,N_9234,N_9506);
or U10830 (N_10830,N_9852,N_9913);
and U10831 (N_10831,N_9858,N_9520);
nand U10832 (N_10832,N_9800,N_9272);
or U10833 (N_10833,N_9971,N_9837);
or U10834 (N_10834,N_9050,N_9118);
and U10835 (N_10835,N_9166,N_9483);
nand U10836 (N_10836,N_9227,N_9545);
nand U10837 (N_10837,N_9154,N_9613);
and U10838 (N_10838,N_9961,N_9964);
nor U10839 (N_10839,N_9002,N_9314);
or U10840 (N_10840,N_9811,N_9252);
xor U10841 (N_10841,N_9774,N_9373);
nor U10842 (N_10842,N_9812,N_9328);
nand U10843 (N_10843,N_9695,N_9831);
and U10844 (N_10844,N_9869,N_9905);
nor U10845 (N_10845,N_9755,N_9711);
or U10846 (N_10846,N_9582,N_9111);
or U10847 (N_10847,N_9457,N_9997);
nand U10848 (N_10848,N_9447,N_9017);
nor U10849 (N_10849,N_9559,N_9064);
nand U10850 (N_10850,N_9443,N_9827);
nand U10851 (N_10851,N_9551,N_9854);
or U10852 (N_10852,N_9197,N_9644);
nand U10853 (N_10853,N_9872,N_9975);
and U10854 (N_10854,N_9459,N_9892);
xor U10855 (N_10855,N_9530,N_9901);
and U10856 (N_10856,N_9704,N_9493);
or U10857 (N_10857,N_9011,N_9374);
nand U10858 (N_10858,N_9362,N_9854);
and U10859 (N_10859,N_9053,N_9399);
nor U10860 (N_10860,N_9573,N_9078);
and U10861 (N_10861,N_9845,N_9287);
nand U10862 (N_10862,N_9524,N_9983);
and U10863 (N_10863,N_9407,N_9166);
nor U10864 (N_10864,N_9652,N_9399);
xor U10865 (N_10865,N_9854,N_9063);
and U10866 (N_10866,N_9560,N_9561);
and U10867 (N_10867,N_9006,N_9084);
nand U10868 (N_10868,N_9437,N_9997);
nor U10869 (N_10869,N_9503,N_9687);
nand U10870 (N_10870,N_9906,N_9451);
nor U10871 (N_10871,N_9362,N_9578);
nor U10872 (N_10872,N_9817,N_9226);
or U10873 (N_10873,N_9000,N_9791);
or U10874 (N_10874,N_9892,N_9275);
and U10875 (N_10875,N_9200,N_9443);
nor U10876 (N_10876,N_9882,N_9573);
and U10877 (N_10877,N_9112,N_9253);
and U10878 (N_10878,N_9594,N_9245);
and U10879 (N_10879,N_9785,N_9847);
or U10880 (N_10880,N_9145,N_9203);
nor U10881 (N_10881,N_9460,N_9475);
nand U10882 (N_10882,N_9222,N_9480);
and U10883 (N_10883,N_9000,N_9909);
and U10884 (N_10884,N_9071,N_9472);
xnor U10885 (N_10885,N_9859,N_9298);
and U10886 (N_10886,N_9389,N_9656);
nand U10887 (N_10887,N_9661,N_9382);
nor U10888 (N_10888,N_9033,N_9768);
and U10889 (N_10889,N_9773,N_9544);
nand U10890 (N_10890,N_9877,N_9726);
nand U10891 (N_10891,N_9852,N_9671);
nand U10892 (N_10892,N_9744,N_9691);
and U10893 (N_10893,N_9330,N_9566);
nor U10894 (N_10894,N_9786,N_9346);
nor U10895 (N_10895,N_9306,N_9749);
xnor U10896 (N_10896,N_9456,N_9496);
nand U10897 (N_10897,N_9313,N_9343);
or U10898 (N_10898,N_9471,N_9966);
nor U10899 (N_10899,N_9471,N_9867);
and U10900 (N_10900,N_9463,N_9666);
and U10901 (N_10901,N_9774,N_9763);
nor U10902 (N_10902,N_9299,N_9563);
or U10903 (N_10903,N_9750,N_9502);
nor U10904 (N_10904,N_9710,N_9610);
and U10905 (N_10905,N_9014,N_9770);
nor U10906 (N_10906,N_9124,N_9558);
or U10907 (N_10907,N_9375,N_9325);
nor U10908 (N_10908,N_9285,N_9736);
xnor U10909 (N_10909,N_9397,N_9114);
nor U10910 (N_10910,N_9184,N_9821);
xnor U10911 (N_10911,N_9026,N_9963);
or U10912 (N_10912,N_9198,N_9473);
xnor U10913 (N_10913,N_9992,N_9090);
xor U10914 (N_10914,N_9099,N_9873);
nor U10915 (N_10915,N_9000,N_9602);
nor U10916 (N_10916,N_9733,N_9543);
nor U10917 (N_10917,N_9096,N_9830);
nand U10918 (N_10918,N_9557,N_9105);
xor U10919 (N_10919,N_9383,N_9919);
and U10920 (N_10920,N_9520,N_9819);
and U10921 (N_10921,N_9922,N_9249);
nand U10922 (N_10922,N_9837,N_9702);
and U10923 (N_10923,N_9177,N_9999);
xnor U10924 (N_10924,N_9521,N_9574);
and U10925 (N_10925,N_9647,N_9555);
or U10926 (N_10926,N_9439,N_9138);
or U10927 (N_10927,N_9129,N_9981);
and U10928 (N_10928,N_9382,N_9259);
and U10929 (N_10929,N_9283,N_9565);
and U10930 (N_10930,N_9561,N_9847);
and U10931 (N_10931,N_9772,N_9073);
or U10932 (N_10932,N_9456,N_9550);
nor U10933 (N_10933,N_9302,N_9827);
nor U10934 (N_10934,N_9316,N_9560);
or U10935 (N_10935,N_9456,N_9011);
nor U10936 (N_10936,N_9131,N_9008);
nand U10937 (N_10937,N_9705,N_9904);
and U10938 (N_10938,N_9021,N_9150);
and U10939 (N_10939,N_9942,N_9582);
and U10940 (N_10940,N_9720,N_9332);
nand U10941 (N_10941,N_9204,N_9786);
and U10942 (N_10942,N_9350,N_9088);
nand U10943 (N_10943,N_9472,N_9497);
and U10944 (N_10944,N_9307,N_9889);
or U10945 (N_10945,N_9591,N_9169);
nand U10946 (N_10946,N_9078,N_9741);
nor U10947 (N_10947,N_9141,N_9748);
nand U10948 (N_10948,N_9142,N_9605);
or U10949 (N_10949,N_9756,N_9297);
nand U10950 (N_10950,N_9496,N_9860);
nor U10951 (N_10951,N_9281,N_9854);
or U10952 (N_10952,N_9265,N_9551);
nor U10953 (N_10953,N_9801,N_9122);
or U10954 (N_10954,N_9592,N_9798);
nand U10955 (N_10955,N_9666,N_9334);
nor U10956 (N_10956,N_9090,N_9813);
and U10957 (N_10957,N_9803,N_9499);
or U10958 (N_10958,N_9539,N_9313);
nand U10959 (N_10959,N_9691,N_9294);
or U10960 (N_10960,N_9116,N_9298);
xnor U10961 (N_10961,N_9055,N_9512);
nor U10962 (N_10962,N_9261,N_9723);
xnor U10963 (N_10963,N_9490,N_9586);
nand U10964 (N_10964,N_9662,N_9320);
or U10965 (N_10965,N_9720,N_9988);
xnor U10966 (N_10966,N_9376,N_9074);
and U10967 (N_10967,N_9543,N_9372);
and U10968 (N_10968,N_9909,N_9201);
xnor U10969 (N_10969,N_9358,N_9501);
and U10970 (N_10970,N_9246,N_9399);
nand U10971 (N_10971,N_9008,N_9671);
nand U10972 (N_10972,N_9768,N_9734);
and U10973 (N_10973,N_9138,N_9355);
and U10974 (N_10974,N_9423,N_9573);
and U10975 (N_10975,N_9185,N_9214);
and U10976 (N_10976,N_9243,N_9545);
nor U10977 (N_10977,N_9894,N_9239);
and U10978 (N_10978,N_9066,N_9628);
nand U10979 (N_10979,N_9383,N_9877);
nand U10980 (N_10980,N_9148,N_9199);
or U10981 (N_10981,N_9187,N_9570);
and U10982 (N_10982,N_9195,N_9396);
nor U10983 (N_10983,N_9928,N_9204);
and U10984 (N_10984,N_9265,N_9739);
and U10985 (N_10985,N_9003,N_9099);
nor U10986 (N_10986,N_9297,N_9543);
nor U10987 (N_10987,N_9468,N_9095);
and U10988 (N_10988,N_9936,N_9131);
and U10989 (N_10989,N_9168,N_9064);
nand U10990 (N_10990,N_9002,N_9053);
and U10991 (N_10991,N_9529,N_9396);
or U10992 (N_10992,N_9685,N_9244);
nor U10993 (N_10993,N_9939,N_9735);
and U10994 (N_10994,N_9061,N_9843);
nand U10995 (N_10995,N_9730,N_9641);
nand U10996 (N_10996,N_9846,N_9670);
and U10997 (N_10997,N_9370,N_9430);
or U10998 (N_10998,N_9612,N_9563);
nand U10999 (N_10999,N_9521,N_9798);
and U11000 (N_11000,N_10470,N_10970);
nor U11001 (N_11001,N_10843,N_10395);
and U11002 (N_11002,N_10789,N_10528);
nand U11003 (N_11003,N_10040,N_10839);
nand U11004 (N_11004,N_10707,N_10036);
nor U11005 (N_11005,N_10238,N_10142);
and U11006 (N_11006,N_10950,N_10364);
and U11007 (N_11007,N_10847,N_10675);
nor U11008 (N_11008,N_10210,N_10713);
nand U11009 (N_11009,N_10367,N_10887);
nand U11010 (N_11010,N_10029,N_10923);
nor U11011 (N_11011,N_10648,N_10737);
nand U11012 (N_11012,N_10141,N_10506);
and U11013 (N_11013,N_10568,N_10001);
and U11014 (N_11014,N_10867,N_10914);
nand U11015 (N_11015,N_10747,N_10077);
nand U11016 (N_11016,N_10301,N_10408);
nand U11017 (N_11017,N_10602,N_10615);
nor U11018 (N_11018,N_10584,N_10700);
or U11019 (N_11019,N_10582,N_10290);
or U11020 (N_11020,N_10668,N_10986);
xnor U11021 (N_11021,N_10913,N_10921);
nand U11022 (N_11022,N_10006,N_10929);
nand U11023 (N_11023,N_10566,N_10828);
or U11024 (N_11024,N_10033,N_10456);
or U11025 (N_11025,N_10162,N_10698);
or U11026 (N_11026,N_10529,N_10341);
or U11027 (N_11027,N_10386,N_10772);
or U11028 (N_11028,N_10540,N_10565);
nor U11029 (N_11029,N_10037,N_10235);
and U11030 (N_11030,N_10373,N_10837);
xnor U11031 (N_11031,N_10908,N_10236);
xor U11032 (N_11032,N_10024,N_10255);
and U11033 (N_11033,N_10628,N_10857);
nor U11034 (N_11034,N_10343,N_10361);
nand U11035 (N_11035,N_10625,N_10308);
and U11036 (N_11036,N_10518,N_10274);
and U11037 (N_11037,N_10441,N_10834);
and U11038 (N_11038,N_10999,N_10905);
or U11039 (N_11039,N_10375,N_10579);
nand U11040 (N_11040,N_10475,N_10760);
xor U11041 (N_11041,N_10152,N_10878);
nand U11042 (N_11042,N_10803,N_10880);
and U11043 (N_11043,N_10727,N_10903);
and U11044 (N_11044,N_10734,N_10153);
nor U11045 (N_11045,N_10937,N_10320);
or U11046 (N_11046,N_10028,N_10632);
nor U11047 (N_11047,N_10273,N_10511);
and U11048 (N_11048,N_10841,N_10881);
nor U11049 (N_11049,N_10168,N_10699);
xor U11050 (N_11050,N_10995,N_10149);
nor U11051 (N_11051,N_10313,N_10716);
nand U11052 (N_11052,N_10773,N_10335);
and U11053 (N_11053,N_10337,N_10187);
or U11054 (N_11054,N_10346,N_10144);
nor U11055 (N_11055,N_10398,N_10665);
xor U11056 (N_11056,N_10497,N_10626);
and U11057 (N_11057,N_10939,N_10151);
and U11058 (N_11058,N_10550,N_10260);
and U11059 (N_11059,N_10073,N_10424);
and U11060 (N_11060,N_10882,N_10865);
or U11061 (N_11061,N_10790,N_10598);
and U11062 (N_11062,N_10534,N_10808);
nand U11063 (N_11063,N_10163,N_10230);
and U11064 (N_11064,N_10557,N_10358);
nand U11065 (N_11065,N_10562,N_10336);
nor U11066 (N_11066,N_10440,N_10067);
and U11067 (N_11067,N_10084,N_10026);
nand U11068 (N_11068,N_10780,N_10183);
nand U11069 (N_11069,N_10059,N_10622);
nand U11070 (N_11070,N_10610,N_10300);
nand U11071 (N_11071,N_10546,N_10436);
xor U11072 (N_11072,N_10606,N_10262);
or U11073 (N_11073,N_10692,N_10414);
and U11074 (N_11074,N_10357,N_10697);
nor U11075 (N_11075,N_10179,N_10081);
and U11076 (N_11076,N_10781,N_10046);
nand U11077 (N_11077,N_10705,N_10286);
or U11078 (N_11078,N_10891,N_10442);
nand U11079 (N_11079,N_10353,N_10463);
and U11080 (N_11080,N_10292,N_10725);
nor U11081 (N_11081,N_10114,N_10186);
xnor U11082 (N_11082,N_10322,N_10647);
nand U11083 (N_11083,N_10748,N_10087);
or U11084 (N_11084,N_10541,N_10879);
nand U11085 (N_11085,N_10056,N_10121);
or U11086 (N_11086,N_10943,N_10108);
nand U11087 (N_11087,N_10985,N_10178);
and U11088 (N_11088,N_10852,N_10385);
nor U11089 (N_11089,N_10821,N_10275);
or U11090 (N_11090,N_10074,N_10011);
nand U11091 (N_11091,N_10493,N_10832);
nor U11092 (N_11092,N_10526,N_10448);
or U11093 (N_11093,N_10502,N_10793);
xnor U11094 (N_11094,N_10754,N_10287);
and U11095 (N_11095,N_10302,N_10979);
nor U11096 (N_11096,N_10244,N_10093);
or U11097 (N_11097,N_10679,N_10406);
nand U11098 (N_11098,N_10912,N_10888);
or U11099 (N_11099,N_10663,N_10989);
xor U11100 (N_11100,N_10718,N_10092);
and U11101 (N_11101,N_10954,N_10237);
or U11102 (N_11102,N_10992,N_10655);
or U11103 (N_11103,N_10927,N_10213);
nand U11104 (N_11104,N_10677,N_10809);
nor U11105 (N_11105,N_10884,N_10597);
and U11106 (N_11106,N_10297,N_10614);
or U11107 (N_11107,N_10695,N_10538);
and U11108 (N_11108,N_10846,N_10942);
and U11109 (N_11109,N_10599,N_10791);
xnor U11110 (N_11110,N_10785,N_10787);
or U11111 (N_11111,N_10418,N_10501);
xnor U11112 (N_11112,N_10629,N_10376);
and U11113 (N_11113,N_10778,N_10473);
nand U11114 (N_11114,N_10279,N_10531);
nand U11115 (N_11115,N_10083,N_10953);
or U11116 (N_11116,N_10131,N_10064);
and U11117 (N_11117,N_10225,N_10390);
nor U11118 (N_11118,N_10160,N_10161);
and U11119 (N_11119,N_10799,N_10082);
xor U11120 (N_11120,N_10769,N_10685);
nand U11121 (N_11121,N_10045,N_10269);
nor U11122 (N_11122,N_10305,N_10894);
or U11123 (N_11123,N_10066,N_10044);
nand U11124 (N_11124,N_10447,N_10527);
nand U11125 (N_11125,N_10415,N_10451);
or U11126 (N_11126,N_10014,N_10472);
nand U11127 (N_11127,N_10673,N_10840);
nor U11128 (N_11128,N_10360,N_10859);
and U11129 (N_11129,N_10078,N_10392);
nand U11130 (N_11130,N_10691,N_10423);
xnor U11131 (N_11131,N_10462,N_10379);
or U11132 (N_11132,N_10570,N_10198);
or U11133 (N_11133,N_10554,N_10958);
nand U11134 (N_11134,N_10826,N_10053);
nand U11135 (N_11135,N_10553,N_10318);
and U11136 (N_11136,N_10963,N_10195);
xor U11137 (N_11137,N_10063,N_10783);
nand U11138 (N_11138,N_10637,N_10898);
nand U11139 (N_11139,N_10136,N_10166);
nand U11140 (N_11140,N_10577,N_10215);
nor U11141 (N_11141,N_10330,N_10978);
nand U11142 (N_11142,N_10129,N_10544);
nor U11143 (N_11143,N_10515,N_10766);
nor U11144 (N_11144,N_10477,N_10890);
and U11145 (N_11145,N_10720,N_10805);
and U11146 (N_11146,N_10116,N_10758);
nor U11147 (N_11147,N_10319,N_10259);
and U11148 (N_11148,N_10678,N_10601);
nand U11149 (N_11149,N_10587,N_10701);
xnor U11150 (N_11150,N_10150,N_10249);
or U11151 (N_11151,N_10214,N_10944);
nor U11152 (N_11152,N_10167,N_10689);
or U11153 (N_11153,N_10118,N_10248);
xnor U11154 (N_11154,N_10315,N_10621);
nand U11155 (N_11155,N_10219,N_10911);
nor U11156 (N_11156,N_10771,N_10323);
or U11157 (N_11157,N_10654,N_10571);
nand U11158 (N_11158,N_10982,N_10619);
and U11159 (N_11159,N_10245,N_10512);
and U11160 (N_11160,N_10062,N_10813);
nand U11161 (N_11161,N_10591,N_10217);
and U11162 (N_11162,N_10103,N_10350);
nand U11163 (N_11163,N_10551,N_10316);
and U11164 (N_11164,N_10674,N_10430);
and U11165 (N_11165,N_10997,N_10095);
or U11166 (N_11166,N_10384,N_10391);
and U11167 (N_11167,N_10946,N_10817);
xor U11168 (N_11168,N_10331,N_10388);
nor U11169 (N_11169,N_10653,N_10508);
xnor U11170 (N_11170,N_10090,N_10712);
nor U11171 (N_11171,N_10422,N_10833);
nand U11172 (N_11172,N_10972,N_10293);
nand U11173 (N_11173,N_10586,N_10509);
or U11174 (N_11174,N_10850,N_10058);
and U11175 (N_11175,N_10750,N_10104);
nand U11176 (N_11176,N_10812,N_10635);
nand U11177 (N_11177,N_10684,N_10844);
and U11178 (N_11178,N_10208,N_10101);
and U11179 (N_11179,N_10362,N_10296);
or U11180 (N_11180,N_10552,N_10450);
xnor U11181 (N_11181,N_10251,N_10572);
and U11182 (N_11182,N_10175,N_10055);
nand U11183 (N_11183,N_10306,N_10875);
and U11184 (N_11184,N_10212,N_10339);
or U11185 (N_11185,N_10542,N_10814);
and U11186 (N_11186,N_10547,N_10688);
nor U11187 (N_11187,N_10389,N_10856);
nand U11188 (N_11188,N_10003,N_10027);
nor U11189 (N_11189,N_10936,N_10457);
nor U11190 (N_11190,N_10170,N_10756);
xnor U11191 (N_11191,N_10644,N_10764);
or U11192 (N_11192,N_10054,N_10981);
nor U11193 (N_11193,N_10495,N_10794);
or U11194 (N_11194,N_10489,N_10966);
nand U11195 (N_11195,N_10471,N_10592);
nand U11196 (N_11196,N_10304,N_10706);
nand U11197 (N_11197,N_10971,N_10117);
or U11198 (N_11198,N_10349,N_10662);
nand U11199 (N_11199,N_10266,N_10123);
xnor U11200 (N_11200,N_10257,N_10798);
nor U11201 (N_11201,N_10897,N_10545);
nor U11202 (N_11202,N_10374,N_10252);
and U11203 (N_11203,N_10576,N_10480);
nand U11204 (N_11204,N_10634,N_10749);
or U11205 (N_11205,N_10231,N_10159);
or U11206 (N_11206,N_10025,N_10034);
nand U11207 (N_11207,N_10413,N_10446);
or U11208 (N_11208,N_10977,N_10835);
and U11209 (N_11209,N_10076,N_10071);
or U11210 (N_11210,N_10061,N_10474);
nor U11211 (N_11211,N_10299,N_10354);
nand U11212 (N_11212,N_10609,N_10145);
nand U11213 (N_11213,N_10445,N_10792);
or U11214 (N_11214,N_10291,N_10605);
nor U11215 (N_11215,N_10731,N_10770);
or U11216 (N_11216,N_10974,N_10928);
or U11217 (N_11217,N_10774,N_10855);
nand U11218 (N_11218,N_10962,N_10365);
nor U11219 (N_11219,N_10735,N_10294);
and U11220 (N_11220,N_10922,N_10940);
and U11221 (N_11221,N_10193,N_10021);
xnor U11222 (N_11222,N_10845,N_10321);
or U11223 (N_11223,N_10952,N_10746);
and U11224 (N_11224,N_10465,N_10079);
nand U11225 (N_11225,N_10065,N_10902);
nand U11226 (N_11226,N_10484,N_10184);
nor U11227 (N_11227,N_10889,N_10642);
nor U11228 (N_11228,N_10454,N_10519);
nor U11229 (N_11229,N_10608,N_10122);
or U11230 (N_11230,N_10106,N_10759);
nor U11231 (N_11231,N_10052,N_10372);
nor U11232 (N_11232,N_10500,N_10652);
xnor U11233 (N_11233,N_10851,N_10125);
nor U11234 (N_11234,N_10172,N_10830);
xor U11235 (N_11235,N_10824,N_10827);
nor U11236 (N_11236,N_10334,N_10466);
nand U11237 (N_11237,N_10307,N_10048);
nand U11238 (N_11238,N_10250,N_10868);
and U11239 (N_11239,N_10990,N_10281);
or U11240 (N_11240,N_10969,N_10504);
nand U11241 (N_11241,N_10567,N_10589);
nand U11242 (N_11242,N_10968,N_10539);
nor U11243 (N_11243,N_10008,N_10267);
nand U11244 (N_11244,N_10514,N_10091);
nor U11245 (N_11245,N_10893,N_10209);
nand U11246 (N_11246,N_10672,N_10325);
and U11247 (N_11247,N_10478,N_10869);
and U11248 (N_11248,N_10831,N_10128);
and U11249 (N_11249,N_10173,N_10516);
nand U11250 (N_11250,N_10853,N_10696);
and U11251 (N_11251,N_10595,N_10917);
or U11252 (N_11252,N_10800,N_10070);
and U11253 (N_11253,N_10871,N_10961);
nor U11254 (N_11254,N_10113,N_10181);
and U11255 (N_11255,N_10263,N_10752);
and U11256 (N_11256,N_10736,N_10924);
nand U11257 (N_11257,N_10607,N_10646);
or U11258 (N_11258,N_10656,N_10892);
or U11259 (N_11259,N_10031,N_10765);
nor U11260 (N_11260,N_10594,N_10485);
xor U11261 (N_11261,N_10254,N_10904);
or U11262 (N_11262,N_10492,N_10521);
and U11263 (N_11263,N_10704,N_10176);
nor U11264 (N_11264,N_10671,N_10657);
nor U11265 (N_11265,N_10435,N_10624);
or U11266 (N_11266,N_10233,N_10741);
or U11267 (N_11267,N_10767,N_10280);
or U11268 (N_11268,N_10177,N_10938);
xor U11269 (N_11269,N_10314,N_10666);
nand U11270 (N_11270,N_10667,N_10755);
and U11271 (N_11271,N_10549,N_10630);
and U11272 (N_11272,N_10548,N_10739);
or U11273 (N_11273,N_10693,N_10427);
nor U11274 (N_11274,N_10745,N_10920);
or U11275 (N_11275,N_10555,N_10140);
nand U11276 (N_11276,N_10007,N_10872);
or U11277 (N_11277,N_10866,N_10107);
nand U11278 (N_11278,N_10721,N_10110);
xor U11279 (N_11279,N_10370,N_10561);
xor U11280 (N_11280,N_10405,N_10197);
and U11281 (N_11281,N_10443,N_10295);
and U11282 (N_11282,N_10503,N_10951);
nand U11283 (N_11283,N_10639,N_10133);
or U11284 (N_11284,N_10910,N_10596);
nand U11285 (N_11285,N_10569,N_10206);
or U11286 (N_11286,N_10222,N_10359);
or U11287 (N_11287,N_10366,N_10660);
nand U11288 (N_11288,N_10333,N_10165);
and U11289 (N_11289,N_10682,N_10156);
and U11290 (N_11290,N_10680,N_10042);
or U11291 (N_11291,N_10728,N_10991);
nor U11292 (N_11292,N_10348,N_10180);
nand U11293 (N_11293,N_10015,N_10967);
nand U11294 (N_11294,N_10883,N_10710);
nand U11295 (N_11295,N_10810,N_10564);
or U11296 (N_11296,N_10310,N_10543);
and U11297 (N_11297,N_10396,N_10139);
nand U11298 (N_11298,N_10253,N_10038);
nor U11299 (N_11299,N_10239,N_10075);
nand U11300 (N_11300,N_10438,N_10873);
nand U11301 (N_11301,N_10203,N_10876);
and U11302 (N_11302,N_10931,N_10957);
or U11303 (N_11303,N_10714,N_10513);
nor U11304 (N_11304,N_10616,N_10407);
and U11305 (N_11305,N_10988,N_10948);
nor U11306 (N_11306,N_10930,N_10722);
and U11307 (N_11307,N_10051,N_10670);
and U11308 (N_11308,N_10815,N_10368);
and U11309 (N_11309,N_10459,N_10494);
nor U11310 (N_11310,N_10686,N_10115);
nand U11311 (N_11311,N_10633,N_10520);
and U11312 (N_11312,N_10009,N_10761);
or U11313 (N_11313,N_10575,N_10804);
and U11314 (N_11314,N_10345,N_10229);
and U11315 (N_11315,N_10189,N_10425);
nor U11316 (N_11316,N_10532,N_10363);
nor U11317 (N_11317,N_10535,N_10285);
and U11318 (N_11318,N_10102,N_10387);
nand U11319 (N_11319,N_10433,N_10017);
xor U11320 (N_11320,N_10949,N_10050);
nand U11321 (N_11321,N_10099,N_10243);
or U11322 (N_11322,N_10687,N_10196);
nand U11323 (N_11323,N_10256,N_10870);
nor U11324 (N_11324,N_10211,N_10041);
or U11325 (N_11325,N_10199,N_10383);
and U11326 (N_11326,N_10732,N_10730);
and U11327 (N_11327,N_10278,N_10094);
nor U11328 (N_11328,N_10811,N_10411);
and U11329 (N_11329,N_10858,N_10127);
and U11330 (N_11330,N_10536,N_10138);
nor U11331 (N_11331,N_10818,N_10220);
or U11332 (N_11332,N_10119,N_10039);
xnor U11333 (N_11333,N_10763,N_10100);
nor U11334 (N_11334,N_10143,N_10378);
nand U11335 (N_11335,N_10482,N_10499);
or U11336 (N_11336,N_10643,N_10158);
nand U11337 (N_11337,N_10973,N_10537);
nand U11338 (N_11338,N_10715,N_10885);
nand U11339 (N_11339,N_10468,N_10915);
or U11340 (N_11340,N_10965,N_10488);
nor U11341 (N_11341,N_10510,N_10620);
and U11342 (N_11342,N_10934,N_10861);
xor U11343 (N_11343,N_10420,N_10207);
xnor U11344 (N_11344,N_10018,N_10795);
nor U11345 (N_11345,N_10347,N_10155);
and U11346 (N_11346,N_10483,N_10702);
xor U11347 (N_11347,N_10505,N_10298);
or U11348 (N_11348,N_10807,N_10218);
or U11349 (N_11349,N_10264,N_10724);
nor U11350 (N_11350,N_10676,N_10221);
and U11351 (N_11351,N_10583,N_10194);
nor U11352 (N_11352,N_10976,N_10690);
or U11353 (N_11353,N_10842,N_10517);
xnor U11354 (N_11354,N_10964,N_10659);
or U11355 (N_11355,N_10088,N_10188);
nand U11356 (N_11356,N_10533,N_10444);
nand U11357 (N_11357,N_10068,N_10733);
and U11358 (N_11358,N_10080,N_10980);
or U11359 (N_11359,N_10010,N_10801);
nand U11360 (N_11360,N_10788,N_10174);
xor U11361 (N_11361,N_10664,N_10895);
nor U11362 (N_11362,N_10192,N_10556);
nand U11363 (N_11363,N_10246,N_10240);
nand U11364 (N_11364,N_10525,N_10578);
nand U11365 (N_11365,N_10288,N_10342);
nand U11366 (N_11366,N_10822,N_10202);
or U11367 (N_11367,N_10854,N_10410);
nand U11368 (N_11368,N_10270,N_10651);
nor U11369 (N_11369,N_10402,N_10004);
nand U11370 (N_11370,N_10340,N_10111);
or U11371 (N_11371,N_10130,N_10224);
xnor U11372 (N_11372,N_10896,N_10434);
nor U11373 (N_11373,N_10559,N_10169);
xnor U11374 (N_11374,N_10057,N_10429);
xnor U11375 (N_11375,N_10581,N_10907);
xnor U11376 (N_11376,N_10439,N_10849);
nor U11377 (N_11377,N_10137,N_10317);
and U11378 (N_11378,N_10190,N_10975);
or U11379 (N_11379,N_10132,N_10098);
and U11380 (N_11380,N_10820,N_10558);
nor U11381 (N_11381,N_10522,N_10779);
xnor U11382 (N_11382,N_10428,N_10636);
nor U11383 (N_11383,N_10185,N_10157);
xor U11384 (N_11384,N_10394,N_10600);
or U11385 (N_11385,N_10000,N_10309);
nor U11386 (N_11386,N_10711,N_10909);
nor U11387 (N_11387,N_10171,N_10352);
or U11388 (N_11388,N_10458,N_10743);
and U11389 (N_11389,N_10983,N_10393);
nand U11390 (N_11390,N_10574,N_10089);
and U11391 (N_11391,N_10344,N_10738);
nor U11392 (N_11392,N_10487,N_10640);
nor U11393 (N_11393,N_10862,N_10901);
and U11394 (N_11394,N_10303,N_10918);
nand U11395 (N_11395,N_10328,N_10311);
and U11396 (N_11396,N_10096,N_10242);
nand U11397 (N_11397,N_10023,N_10658);
nor U11398 (N_11398,N_10836,N_10593);
nor U11399 (N_11399,N_10481,N_10412);
nor U11400 (N_11400,N_10588,N_10984);
nor U11401 (N_11401,N_10782,N_10329);
and U11402 (N_11402,N_10226,N_10530);
and U11403 (N_11403,N_10105,N_10573);
or U11404 (N_11404,N_10825,N_10277);
nor U11405 (N_11405,N_10786,N_10449);
nor U11406 (N_11406,N_10191,N_10708);
nor U11407 (N_11407,N_10627,N_10421);
or U11408 (N_11408,N_10806,N_10204);
or U11409 (N_11409,N_10563,N_10816);
or U11410 (N_11410,N_10613,N_10327);
or U11411 (N_11411,N_10135,N_10703);
xor U11412 (N_11412,N_10523,N_10013);
nor U11413 (N_11413,N_10899,N_10426);
nand U11414 (N_11414,N_10416,N_10284);
or U11415 (N_11415,N_10560,N_10524);
xor U11416 (N_11416,N_10247,N_10241);
and U11417 (N_11417,N_10332,N_10460);
nand U11418 (N_11418,N_10960,N_10124);
nand U11419 (N_11419,N_10400,N_10823);
nor U11420 (N_11420,N_10603,N_10476);
or U11421 (N_11421,N_10604,N_10437);
and U11422 (N_11422,N_10941,N_10906);
nor U11423 (N_11423,N_10399,N_10002);
nand U11424 (N_11424,N_10618,N_10043);
nand U11425 (N_11425,N_10987,N_10694);
nor U11426 (N_11426,N_10631,N_10380);
nor U11427 (N_11427,N_10265,N_10819);
nand U11428 (N_11428,N_10261,N_10258);
or U11429 (N_11429,N_10030,N_10369);
nor U11430 (N_11430,N_10276,N_10461);
nand U11431 (N_11431,N_10020,N_10926);
nor U11432 (N_11432,N_10355,N_10864);
and U11433 (N_11433,N_10469,N_10955);
nor U11434 (N_11434,N_10757,N_10996);
nor U11435 (N_11435,N_10289,N_10019);
nor U11436 (N_11436,N_10200,N_10126);
or U11437 (N_11437,N_10409,N_10498);
or U11438 (N_11438,N_10611,N_10356);
nor U11439 (N_11439,N_10382,N_10998);
xnor U11440 (N_11440,N_10863,N_10060);
xnor U11441 (N_11441,N_10326,N_10232);
nor U11442 (N_11442,N_10147,N_10086);
and U11443 (N_11443,N_10829,N_10935);
nor U11444 (N_11444,N_10669,N_10377);
or U11445 (N_11445,N_10947,N_10886);
and U11446 (N_11446,N_10455,N_10507);
nand U11447 (N_11447,N_10638,N_10993);
nand U11448 (N_11448,N_10762,N_10069);
xnor U11449 (N_11449,N_10617,N_10403);
nand U11450 (N_11450,N_10959,N_10479);
nor U11451 (N_11451,N_10201,N_10109);
and U11452 (N_11452,N_10032,N_10838);
nand U11453 (N_11453,N_10623,N_10216);
and U11454 (N_11454,N_10723,N_10223);
and U11455 (N_11455,N_10612,N_10775);
xor U11456 (N_11456,N_10035,N_10282);
xnor U11457 (N_11457,N_10228,N_10148);
and U11458 (N_11458,N_10681,N_10419);
and U11459 (N_11459,N_10283,N_10154);
xor U11460 (N_11460,N_10351,N_10085);
xnor U11461 (N_11461,N_10994,N_10072);
or U11462 (N_11462,N_10047,N_10709);
xor U11463 (N_11463,N_10397,N_10312);
nand U11464 (N_11464,N_10401,N_10134);
or U11465 (N_11465,N_10683,N_10112);
nor U11466 (N_11466,N_10661,N_10784);
or U11467 (N_11467,N_10005,N_10585);
or U11468 (N_11468,N_10467,N_10120);
nor U11469 (N_11469,N_10182,N_10146);
and U11470 (N_11470,N_10645,N_10726);
nand U11471 (N_11471,N_10848,N_10381);
or U11472 (N_11472,N_10945,N_10486);
or U11473 (N_11473,N_10268,N_10205);
nor U11474 (N_11474,N_10900,N_10742);
nor U11475 (N_11475,N_10227,N_10590);
nor U11476 (N_11476,N_10496,N_10464);
or U11477 (N_11477,N_10860,N_10404);
and U11478 (N_11478,N_10768,N_10491);
nor U11479 (N_11479,N_10796,N_10338);
and U11480 (N_11480,N_10012,N_10164);
nand U11481 (N_11481,N_10371,N_10431);
nand U11482 (N_11482,N_10049,N_10933);
or U11483 (N_11483,N_10932,N_10417);
nor U11484 (N_11484,N_10751,N_10919);
xor U11485 (N_11485,N_10753,N_10777);
nand U11486 (N_11486,N_10916,N_10797);
and U11487 (N_11487,N_10272,N_10925);
nand U11488 (N_11488,N_10490,N_10719);
and U11489 (N_11489,N_10776,N_10744);
nand U11490 (N_11490,N_10271,N_10877);
or U11491 (N_11491,N_10649,N_10016);
or U11492 (N_11492,N_10650,N_10729);
nor U11493 (N_11493,N_10452,N_10641);
nor U11494 (N_11494,N_10874,N_10802);
and U11495 (N_11495,N_10432,N_10022);
and U11496 (N_11496,N_10580,N_10097);
and U11497 (N_11497,N_10717,N_10956);
or U11498 (N_11498,N_10234,N_10453);
and U11499 (N_11499,N_10740,N_10324);
and U11500 (N_11500,N_10228,N_10354);
nand U11501 (N_11501,N_10752,N_10445);
or U11502 (N_11502,N_10968,N_10075);
and U11503 (N_11503,N_10031,N_10741);
or U11504 (N_11504,N_10589,N_10127);
or U11505 (N_11505,N_10578,N_10686);
and U11506 (N_11506,N_10799,N_10119);
nor U11507 (N_11507,N_10450,N_10010);
xor U11508 (N_11508,N_10254,N_10029);
nor U11509 (N_11509,N_10262,N_10783);
xor U11510 (N_11510,N_10553,N_10703);
or U11511 (N_11511,N_10097,N_10540);
xnor U11512 (N_11512,N_10089,N_10485);
nand U11513 (N_11513,N_10855,N_10436);
and U11514 (N_11514,N_10604,N_10518);
nor U11515 (N_11515,N_10070,N_10254);
or U11516 (N_11516,N_10609,N_10104);
or U11517 (N_11517,N_10563,N_10604);
or U11518 (N_11518,N_10101,N_10699);
or U11519 (N_11519,N_10517,N_10782);
and U11520 (N_11520,N_10486,N_10213);
nand U11521 (N_11521,N_10009,N_10089);
nand U11522 (N_11522,N_10957,N_10093);
nand U11523 (N_11523,N_10485,N_10894);
and U11524 (N_11524,N_10873,N_10526);
nor U11525 (N_11525,N_10398,N_10178);
or U11526 (N_11526,N_10795,N_10381);
nand U11527 (N_11527,N_10694,N_10441);
nor U11528 (N_11528,N_10882,N_10361);
or U11529 (N_11529,N_10919,N_10975);
xor U11530 (N_11530,N_10399,N_10306);
nor U11531 (N_11531,N_10513,N_10732);
nor U11532 (N_11532,N_10269,N_10727);
nor U11533 (N_11533,N_10566,N_10255);
and U11534 (N_11534,N_10987,N_10323);
and U11535 (N_11535,N_10622,N_10377);
nor U11536 (N_11536,N_10428,N_10169);
or U11537 (N_11537,N_10356,N_10864);
or U11538 (N_11538,N_10160,N_10131);
and U11539 (N_11539,N_10082,N_10451);
or U11540 (N_11540,N_10745,N_10018);
and U11541 (N_11541,N_10441,N_10942);
nor U11542 (N_11542,N_10539,N_10459);
nand U11543 (N_11543,N_10243,N_10064);
nand U11544 (N_11544,N_10992,N_10463);
nand U11545 (N_11545,N_10820,N_10062);
and U11546 (N_11546,N_10789,N_10862);
xor U11547 (N_11547,N_10219,N_10075);
nor U11548 (N_11548,N_10314,N_10877);
and U11549 (N_11549,N_10605,N_10062);
or U11550 (N_11550,N_10138,N_10938);
nand U11551 (N_11551,N_10367,N_10279);
or U11552 (N_11552,N_10423,N_10375);
xnor U11553 (N_11553,N_10132,N_10797);
xnor U11554 (N_11554,N_10709,N_10586);
and U11555 (N_11555,N_10266,N_10501);
or U11556 (N_11556,N_10931,N_10418);
nand U11557 (N_11557,N_10395,N_10838);
and U11558 (N_11558,N_10410,N_10328);
or U11559 (N_11559,N_10993,N_10588);
nor U11560 (N_11560,N_10257,N_10306);
nand U11561 (N_11561,N_10317,N_10419);
or U11562 (N_11562,N_10988,N_10493);
or U11563 (N_11563,N_10208,N_10275);
and U11564 (N_11564,N_10227,N_10136);
and U11565 (N_11565,N_10024,N_10917);
nor U11566 (N_11566,N_10925,N_10118);
or U11567 (N_11567,N_10395,N_10592);
and U11568 (N_11568,N_10712,N_10041);
or U11569 (N_11569,N_10954,N_10558);
and U11570 (N_11570,N_10992,N_10475);
or U11571 (N_11571,N_10987,N_10434);
and U11572 (N_11572,N_10564,N_10801);
or U11573 (N_11573,N_10186,N_10296);
nor U11574 (N_11574,N_10514,N_10066);
or U11575 (N_11575,N_10191,N_10950);
and U11576 (N_11576,N_10096,N_10080);
nand U11577 (N_11577,N_10084,N_10979);
or U11578 (N_11578,N_10665,N_10174);
and U11579 (N_11579,N_10622,N_10324);
or U11580 (N_11580,N_10913,N_10437);
nand U11581 (N_11581,N_10663,N_10818);
nor U11582 (N_11582,N_10296,N_10786);
and U11583 (N_11583,N_10414,N_10208);
nand U11584 (N_11584,N_10273,N_10070);
or U11585 (N_11585,N_10844,N_10425);
nor U11586 (N_11586,N_10310,N_10224);
or U11587 (N_11587,N_10930,N_10439);
or U11588 (N_11588,N_10222,N_10447);
nor U11589 (N_11589,N_10866,N_10125);
nand U11590 (N_11590,N_10985,N_10885);
or U11591 (N_11591,N_10381,N_10559);
and U11592 (N_11592,N_10686,N_10801);
or U11593 (N_11593,N_10162,N_10367);
nor U11594 (N_11594,N_10149,N_10837);
or U11595 (N_11595,N_10713,N_10414);
or U11596 (N_11596,N_10316,N_10712);
nor U11597 (N_11597,N_10390,N_10903);
and U11598 (N_11598,N_10927,N_10823);
nand U11599 (N_11599,N_10908,N_10497);
or U11600 (N_11600,N_10208,N_10042);
nand U11601 (N_11601,N_10607,N_10101);
nand U11602 (N_11602,N_10638,N_10691);
and U11603 (N_11603,N_10015,N_10589);
nand U11604 (N_11604,N_10825,N_10955);
nor U11605 (N_11605,N_10522,N_10432);
nor U11606 (N_11606,N_10411,N_10395);
xnor U11607 (N_11607,N_10401,N_10444);
nor U11608 (N_11608,N_10734,N_10944);
nor U11609 (N_11609,N_10801,N_10039);
nor U11610 (N_11610,N_10650,N_10331);
nand U11611 (N_11611,N_10379,N_10127);
and U11612 (N_11612,N_10489,N_10843);
xnor U11613 (N_11613,N_10788,N_10008);
nand U11614 (N_11614,N_10546,N_10442);
nor U11615 (N_11615,N_10939,N_10395);
xnor U11616 (N_11616,N_10622,N_10055);
nor U11617 (N_11617,N_10485,N_10806);
nor U11618 (N_11618,N_10064,N_10306);
and U11619 (N_11619,N_10780,N_10173);
and U11620 (N_11620,N_10070,N_10940);
nor U11621 (N_11621,N_10697,N_10826);
or U11622 (N_11622,N_10249,N_10246);
nor U11623 (N_11623,N_10737,N_10226);
nor U11624 (N_11624,N_10640,N_10094);
nand U11625 (N_11625,N_10699,N_10766);
xnor U11626 (N_11626,N_10641,N_10790);
or U11627 (N_11627,N_10615,N_10541);
nor U11628 (N_11628,N_10588,N_10955);
nand U11629 (N_11629,N_10558,N_10114);
or U11630 (N_11630,N_10828,N_10996);
nor U11631 (N_11631,N_10758,N_10078);
nor U11632 (N_11632,N_10009,N_10034);
or U11633 (N_11633,N_10022,N_10903);
and U11634 (N_11634,N_10359,N_10943);
and U11635 (N_11635,N_10361,N_10417);
or U11636 (N_11636,N_10515,N_10998);
nor U11637 (N_11637,N_10922,N_10532);
xor U11638 (N_11638,N_10656,N_10625);
or U11639 (N_11639,N_10011,N_10086);
or U11640 (N_11640,N_10114,N_10135);
and U11641 (N_11641,N_10246,N_10447);
nand U11642 (N_11642,N_10056,N_10022);
or U11643 (N_11643,N_10730,N_10623);
and U11644 (N_11644,N_10267,N_10849);
and U11645 (N_11645,N_10600,N_10341);
or U11646 (N_11646,N_10671,N_10368);
or U11647 (N_11647,N_10366,N_10782);
nand U11648 (N_11648,N_10674,N_10118);
nor U11649 (N_11649,N_10712,N_10667);
and U11650 (N_11650,N_10844,N_10430);
and U11651 (N_11651,N_10177,N_10646);
and U11652 (N_11652,N_10902,N_10179);
xor U11653 (N_11653,N_10247,N_10840);
nor U11654 (N_11654,N_10335,N_10895);
xnor U11655 (N_11655,N_10485,N_10851);
nor U11656 (N_11656,N_10525,N_10737);
or U11657 (N_11657,N_10368,N_10548);
nand U11658 (N_11658,N_10955,N_10247);
and U11659 (N_11659,N_10564,N_10144);
nor U11660 (N_11660,N_10211,N_10155);
and U11661 (N_11661,N_10767,N_10906);
or U11662 (N_11662,N_10889,N_10016);
or U11663 (N_11663,N_10369,N_10125);
nand U11664 (N_11664,N_10022,N_10546);
or U11665 (N_11665,N_10905,N_10964);
nor U11666 (N_11666,N_10264,N_10815);
nor U11667 (N_11667,N_10341,N_10644);
and U11668 (N_11668,N_10870,N_10808);
nand U11669 (N_11669,N_10458,N_10868);
nor U11670 (N_11670,N_10879,N_10790);
nor U11671 (N_11671,N_10045,N_10021);
and U11672 (N_11672,N_10639,N_10143);
nor U11673 (N_11673,N_10754,N_10521);
or U11674 (N_11674,N_10968,N_10961);
nand U11675 (N_11675,N_10905,N_10358);
or U11676 (N_11676,N_10224,N_10783);
nand U11677 (N_11677,N_10115,N_10650);
nor U11678 (N_11678,N_10445,N_10351);
nand U11679 (N_11679,N_10403,N_10729);
xnor U11680 (N_11680,N_10268,N_10925);
nand U11681 (N_11681,N_10781,N_10771);
xor U11682 (N_11682,N_10817,N_10300);
nand U11683 (N_11683,N_10040,N_10967);
or U11684 (N_11684,N_10746,N_10595);
or U11685 (N_11685,N_10563,N_10873);
nand U11686 (N_11686,N_10281,N_10091);
or U11687 (N_11687,N_10099,N_10268);
or U11688 (N_11688,N_10910,N_10829);
nand U11689 (N_11689,N_10162,N_10133);
nand U11690 (N_11690,N_10691,N_10404);
or U11691 (N_11691,N_10810,N_10344);
and U11692 (N_11692,N_10193,N_10660);
nand U11693 (N_11693,N_10753,N_10950);
or U11694 (N_11694,N_10436,N_10011);
or U11695 (N_11695,N_10628,N_10552);
nor U11696 (N_11696,N_10316,N_10773);
nor U11697 (N_11697,N_10413,N_10433);
nor U11698 (N_11698,N_10472,N_10302);
and U11699 (N_11699,N_10173,N_10324);
and U11700 (N_11700,N_10863,N_10965);
nand U11701 (N_11701,N_10910,N_10261);
or U11702 (N_11702,N_10293,N_10298);
nand U11703 (N_11703,N_10929,N_10831);
nor U11704 (N_11704,N_10532,N_10571);
or U11705 (N_11705,N_10302,N_10103);
or U11706 (N_11706,N_10631,N_10796);
or U11707 (N_11707,N_10802,N_10804);
and U11708 (N_11708,N_10984,N_10992);
or U11709 (N_11709,N_10875,N_10486);
and U11710 (N_11710,N_10179,N_10526);
nor U11711 (N_11711,N_10585,N_10197);
or U11712 (N_11712,N_10370,N_10522);
and U11713 (N_11713,N_10248,N_10582);
nor U11714 (N_11714,N_10217,N_10978);
nand U11715 (N_11715,N_10156,N_10989);
or U11716 (N_11716,N_10864,N_10684);
and U11717 (N_11717,N_10549,N_10205);
and U11718 (N_11718,N_10316,N_10209);
nor U11719 (N_11719,N_10811,N_10611);
and U11720 (N_11720,N_10649,N_10442);
nand U11721 (N_11721,N_10341,N_10722);
and U11722 (N_11722,N_10406,N_10258);
or U11723 (N_11723,N_10971,N_10593);
nor U11724 (N_11724,N_10975,N_10950);
and U11725 (N_11725,N_10754,N_10042);
nor U11726 (N_11726,N_10568,N_10493);
nor U11727 (N_11727,N_10889,N_10267);
nand U11728 (N_11728,N_10645,N_10716);
xnor U11729 (N_11729,N_10628,N_10391);
or U11730 (N_11730,N_10433,N_10681);
nand U11731 (N_11731,N_10348,N_10882);
nand U11732 (N_11732,N_10342,N_10685);
xnor U11733 (N_11733,N_10606,N_10571);
xor U11734 (N_11734,N_10014,N_10531);
and U11735 (N_11735,N_10162,N_10079);
and U11736 (N_11736,N_10329,N_10536);
or U11737 (N_11737,N_10242,N_10243);
and U11738 (N_11738,N_10672,N_10298);
and U11739 (N_11739,N_10814,N_10338);
and U11740 (N_11740,N_10821,N_10005);
xnor U11741 (N_11741,N_10370,N_10980);
and U11742 (N_11742,N_10822,N_10116);
xor U11743 (N_11743,N_10459,N_10067);
nor U11744 (N_11744,N_10356,N_10571);
and U11745 (N_11745,N_10744,N_10895);
nand U11746 (N_11746,N_10713,N_10659);
or U11747 (N_11747,N_10816,N_10039);
nor U11748 (N_11748,N_10009,N_10196);
xor U11749 (N_11749,N_10456,N_10988);
nand U11750 (N_11750,N_10768,N_10481);
or U11751 (N_11751,N_10108,N_10381);
nor U11752 (N_11752,N_10648,N_10367);
or U11753 (N_11753,N_10743,N_10169);
nand U11754 (N_11754,N_10597,N_10937);
and U11755 (N_11755,N_10441,N_10193);
nor U11756 (N_11756,N_10274,N_10439);
and U11757 (N_11757,N_10399,N_10383);
and U11758 (N_11758,N_10533,N_10641);
nand U11759 (N_11759,N_10441,N_10635);
nand U11760 (N_11760,N_10748,N_10450);
and U11761 (N_11761,N_10091,N_10791);
nand U11762 (N_11762,N_10646,N_10123);
xnor U11763 (N_11763,N_10433,N_10730);
or U11764 (N_11764,N_10179,N_10167);
nor U11765 (N_11765,N_10332,N_10645);
nand U11766 (N_11766,N_10128,N_10384);
nor U11767 (N_11767,N_10408,N_10684);
nand U11768 (N_11768,N_10338,N_10210);
nand U11769 (N_11769,N_10485,N_10183);
nand U11770 (N_11770,N_10391,N_10907);
nand U11771 (N_11771,N_10024,N_10521);
or U11772 (N_11772,N_10439,N_10925);
nand U11773 (N_11773,N_10246,N_10672);
and U11774 (N_11774,N_10514,N_10871);
xnor U11775 (N_11775,N_10968,N_10869);
and U11776 (N_11776,N_10777,N_10703);
nand U11777 (N_11777,N_10743,N_10412);
xnor U11778 (N_11778,N_10036,N_10140);
xnor U11779 (N_11779,N_10297,N_10195);
nand U11780 (N_11780,N_10201,N_10486);
or U11781 (N_11781,N_10596,N_10601);
and U11782 (N_11782,N_10889,N_10513);
xnor U11783 (N_11783,N_10775,N_10863);
nor U11784 (N_11784,N_10961,N_10028);
xnor U11785 (N_11785,N_10985,N_10424);
nor U11786 (N_11786,N_10294,N_10261);
or U11787 (N_11787,N_10368,N_10924);
and U11788 (N_11788,N_10968,N_10245);
xor U11789 (N_11789,N_10273,N_10174);
and U11790 (N_11790,N_10087,N_10081);
or U11791 (N_11791,N_10704,N_10078);
or U11792 (N_11792,N_10522,N_10245);
and U11793 (N_11793,N_10452,N_10736);
nand U11794 (N_11794,N_10330,N_10300);
or U11795 (N_11795,N_10781,N_10607);
or U11796 (N_11796,N_10413,N_10254);
nor U11797 (N_11797,N_10957,N_10741);
and U11798 (N_11798,N_10284,N_10186);
nand U11799 (N_11799,N_10166,N_10340);
and U11800 (N_11800,N_10949,N_10200);
nand U11801 (N_11801,N_10598,N_10170);
and U11802 (N_11802,N_10114,N_10567);
nand U11803 (N_11803,N_10986,N_10769);
nand U11804 (N_11804,N_10198,N_10515);
nor U11805 (N_11805,N_10822,N_10417);
or U11806 (N_11806,N_10433,N_10412);
and U11807 (N_11807,N_10254,N_10052);
or U11808 (N_11808,N_10446,N_10326);
and U11809 (N_11809,N_10892,N_10342);
nand U11810 (N_11810,N_10239,N_10698);
nor U11811 (N_11811,N_10080,N_10537);
nor U11812 (N_11812,N_10782,N_10682);
nand U11813 (N_11813,N_10463,N_10579);
and U11814 (N_11814,N_10613,N_10129);
and U11815 (N_11815,N_10580,N_10718);
and U11816 (N_11816,N_10269,N_10553);
and U11817 (N_11817,N_10329,N_10961);
or U11818 (N_11818,N_10409,N_10462);
and U11819 (N_11819,N_10694,N_10831);
and U11820 (N_11820,N_10306,N_10890);
xnor U11821 (N_11821,N_10927,N_10430);
nor U11822 (N_11822,N_10523,N_10945);
and U11823 (N_11823,N_10982,N_10480);
nand U11824 (N_11824,N_10964,N_10514);
xnor U11825 (N_11825,N_10547,N_10734);
or U11826 (N_11826,N_10897,N_10501);
and U11827 (N_11827,N_10565,N_10290);
and U11828 (N_11828,N_10344,N_10380);
nand U11829 (N_11829,N_10477,N_10765);
xor U11830 (N_11830,N_10758,N_10544);
or U11831 (N_11831,N_10347,N_10897);
nand U11832 (N_11832,N_10130,N_10020);
nor U11833 (N_11833,N_10205,N_10084);
nor U11834 (N_11834,N_10300,N_10849);
or U11835 (N_11835,N_10143,N_10956);
nor U11836 (N_11836,N_10569,N_10266);
or U11837 (N_11837,N_10502,N_10471);
nor U11838 (N_11838,N_10248,N_10780);
and U11839 (N_11839,N_10839,N_10897);
nand U11840 (N_11840,N_10787,N_10363);
and U11841 (N_11841,N_10077,N_10624);
nor U11842 (N_11842,N_10944,N_10875);
nor U11843 (N_11843,N_10946,N_10628);
nand U11844 (N_11844,N_10731,N_10171);
nor U11845 (N_11845,N_10701,N_10240);
and U11846 (N_11846,N_10309,N_10179);
nor U11847 (N_11847,N_10180,N_10276);
nor U11848 (N_11848,N_10742,N_10234);
and U11849 (N_11849,N_10658,N_10041);
nand U11850 (N_11850,N_10829,N_10061);
and U11851 (N_11851,N_10506,N_10792);
or U11852 (N_11852,N_10764,N_10892);
or U11853 (N_11853,N_10368,N_10162);
or U11854 (N_11854,N_10785,N_10293);
nand U11855 (N_11855,N_10824,N_10260);
nor U11856 (N_11856,N_10533,N_10981);
or U11857 (N_11857,N_10935,N_10400);
or U11858 (N_11858,N_10635,N_10817);
nand U11859 (N_11859,N_10046,N_10017);
or U11860 (N_11860,N_10132,N_10970);
or U11861 (N_11861,N_10202,N_10650);
nor U11862 (N_11862,N_10528,N_10794);
or U11863 (N_11863,N_10892,N_10876);
xor U11864 (N_11864,N_10676,N_10574);
and U11865 (N_11865,N_10866,N_10393);
nand U11866 (N_11866,N_10691,N_10388);
or U11867 (N_11867,N_10970,N_10701);
and U11868 (N_11868,N_10135,N_10656);
nor U11869 (N_11869,N_10795,N_10975);
nand U11870 (N_11870,N_10044,N_10035);
nor U11871 (N_11871,N_10290,N_10431);
nand U11872 (N_11872,N_10044,N_10632);
or U11873 (N_11873,N_10416,N_10768);
nor U11874 (N_11874,N_10543,N_10355);
nor U11875 (N_11875,N_10994,N_10028);
nand U11876 (N_11876,N_10575,N_10642);
or U11877 (N_11877,N_10009,N_10890);
or U11878 (N_11878,N_10458,N_10278);
nand U11879 (N_11879,N_10678,N_10914);
or U11880 (N_11880,N_10924,N_10282);
nor U11881 (N_11881,N_10106,N_10344);
nand U11882 (N_11882,N_10633,N_10942);
nor U11883 (N_11883,N_10247,N_10611);
nor U11884 (N_11884,N_10279,N_10631);
nand U11885 (N_11885,N_10027,N_10881);
nand U11886 (N_11886,N_10323,N_10233);
nand U11887 (N_11887,N_10087,N_10764);
or U11888 (N_11888,N_10801,N_10017);
or U11889 (N_11889,N_10029,N_10176);
and U11890 (N_11890,N_10898,N_10023);
and U11891 (N_11891,N_10617,N_10929);
nor U11892 (N_11892,N_10731,N_10684);
and U11893 (N_11893,N_10075,N_10920);
nor U11894 (N_11894,N_10643,N_10949);
nor U11895 (N_11895,N_10772,N_10505);
nand U11896 (N_11896,N_10635,N_10115);
or U11897 (N_11897,N_10814,N_10053);
and U11898 (N_11898,N_10974,N_10010);
or U11899 (N_11899,N_10086,N_10506);
and U11900 (N_11900,N_10760,N_10015);
nor U11901 (N_11901,N_10883,N_10706);
nor U11902 (N_11902,N_10680,N_10708);
or U11903 (N_11903,N_10524,N_10979);
xnor U11904 (N_11904,N_10753,N_10052);
nand U11905 (N_11905,N_10662,N_10177);
or U11906 (N_11906,N_10908,N_10468);
or U11907 (N_11907,N_10433,N_10411);
or U11908 (N_11908,N_10654,N_10456);
nor U11909 (N_11909,N_10879,N_10225);
nor U11910 (N_11910,N_10236,N_10665);
nor U11911 (N_11911,N_10967,N_10497);
or U11912 (N_11912,N_10606,N_10633);
or U11913 (N_11913,N_10256,N_10875);
nor U11914 (N_11914,N_10218,N_10777);
and U11915 (N_11915,N_10299,N_10431);
or U11916 (N_11916,N_10567,N_10499);
nor U11917 (N_11917,N_10376,N_10386);
or U11918 (N_11918,N_10732,N_10332);
or U11919 (N_11919,N_10411,N_10324);
and U11920 (N_11920,N_10764,N_10682);
or U11921 (N_11921,N_10010,N_10868);
or U11922 (N_11922,N_10652,N_10212);
and U11923 (N_11923,N_10782,N_10343);
xor U11924 (N_11924,N_10230,N_10178);
or U11925 (N_11925,N_10206,N_10242);
or U11926 (N_11926,N_10980,N_10649);
xnor U11927 (N_11927,N_10493,N_10787);
nor U11928 (N_11928,N_10221,N_10739);
nor U11929 (N_11929,N_10737,N_10095);
nor U11930 (N_11930,N_10136,N_10044);
nor U11931 (N_11931,N_10197,N_10635);
nand U11932 (N_11932,N_10768,N_10494);
xnor U11933 (N_11933,N_10202,N_10468);
nor U11934 (N_11934,N_10011,N_10191);
nor U11935 (N_11935,N_10090,N_10606);
or U11936 (N_11936,N_10793,N_10371);
nand U11937 (N_11937,N_10252,N_10403);
and U11938 (N_11938,N_10084,N_10208);
and U11939 (N_11939,N_10392,N_10252);
nor U11940 (N_11940,N_10496,N_10192);
and U11941 (N_11941,N_10494,N_10277);
nor U11942 (N_11942,N_10033,N_10979);
nand U11943 (N_11943,N_10345,N_10325);
nand U11944 (N_11944,N_10993,N_10270);
nand U11945 (N_11945,N_10409,N_10807);
and U11946 (N_11946,N_10235,N_10892);
or U11947 (N_11947,N_10472,N_10951);
xor U11948 (N_11948,N_10595,N_10536);
nor U11949 (N_11949,N_10462,N_10546);
xnor U11950 (N_11950,N_10382,N_10120);
and U11951 (N_11951,N_10109,N_10470);
nor U11952 (N_11952,N_10262,N_10927);
nor U11953 (N_11953,N_10178,N_10602);
nand U11954 (N_11954,N_10085,N_10510);
nor U11955 (N_11955,N_10395,N_10591);
and U11956 (N_11956,N_10616,N_10406);
or U11957 (N_11957,N_10283,N_10052);
nor U11958 (N_11958,N_10642,N_10198);
or U11959 (N_11959,N_10645,N_10125);
and U11960 (N_11960,N_10929,N_10829);
or U11961 (N_11961,N_10295,N_10721);
nand U11962 (N_11962,N_10169,N_10232);
and U11963 (N_11963,N_10449,N_10217);
nand U11964 (N_11964,N_10870,N_10698);
xnor U11965 (N_11965,N_10711,N_10266);
or U11966 (N_11966,N_10399,N_10855);
nor U11967 (N_11967,N_10306,N_10196);
and U11968 (N_11968,N_10819,N_10467);
and U11969 (N_11969,N_10425,N_10071);
or U11970 (N_11970,N_10051,N_10072);
or U11971 (N_11971,N_10310,N_10920);
nor U11972 (N_11972,N_10303,N_10179);
xor U11973 (N_11973,N_10693,N_10762);
nor U11974 (N_11974,N_10425,N_10210);
nor U11975 (N_11975,N_10076,N_10450);
or U11976 (N_11976,N_10356,N_10911);
nor U11977 (N_11977,N_10844,N_10479);
and U11978 (N_11978,N_10775,N_10014);
and U11979 (N_11979,N_10073,N_10113);
and U11980 (N_11980,N_10749,N_10491);
nor U11981 (N_11981,N_10460,N_10687);
nor U11982 (N_11982,N_10163,N_10219);
nor U11983 (N_11983,N_10854,N_10592);
or U11984 (N_11984,N_10456,N_10816);
and U11985 (N_11985,N_10098,N_10991);
or U11986 (N_11986,N_10987,N_10689);
xor U11987 (N_11987,N_10506,N_10269);
nor U11988 (N_11988,N_10254,N_10601);
nand U11989 (N_11989,N_10258,N_10982);
nand U11990 (N_11990,N_10719,N_10371);
and U11991 (N_11991,N_10347,N_10569);
nand U11992 (N_11992,N_10421,N_10408);
nor U11993 (N_11993,N_10289,N_10682);
or U11994 (N_11994,N_10566,N_10812);
and U11995 (N_11995,N_10565,N_10605);
or U11996 (N_11996,N_10514,N_10838);
or U11997 (N_11997,N_10011,N_10942);
nand U11998 (N_11998,N_10081,N_10473);
or U11999 (N_11999,N_10251,N_10561);
nand U12000 (N_12000,N_11913,N_11458);
and U12001 (N_12001,N_11055,N_11481);
nand U12002 (N_12002,N_11485,N_11126);
nand U12003 (N_12003,N_11045,N_11155);
or U12004 (N_12004,N_11486,N_11016);
and U12005 (N_12005,N_11651,N_11991);
and U12006 (N_12006,N_11551,N_11043);
and U12007 (N_12007,N_11897,N_11544);
or U12008 (N_12008,N_11097,N_11877);
and U12009 (N_12009,N_11215,N_11953);
nand U12010 (N_12010,N_11052,N_11150);
and U12011 (N_12011,N_11316,N_11313);
and U12012 (N_12012,N_11800,N_11391);
nand U12013 (N_12013,N_11618,N_11034);
or U12014 (N_12014,N_11219,N_11275);
nand U12015 (N_12015,N_11955,N_11373);
nor U12016 (N_12016,N_11254,N_11195);
or U12017 (N_12017,N_11904,N_11790);
nor U12018 (N_12018,N_11082,N_11850);
and U12019 (N_12019,N_11437,N_11410);
and U12020 (N_12020,N_11846,N_11228);
and U12021 (N_12021,N_11687,N_11030);
or U12022 (N_12022,N_11114,N_11958);
or U12023 (N_12023,N_11723,N_11200);
and U12024 (N_12024,N_11883,N_11835);
xor U12025 (N_12025,N_11546,N_11435);
nand U12026 (N_12026,N_11364,N_11803);
nor U12027 (N_12027,N_11103,N_11164);
or U12028 (N_12028,N_11068,N_11880);
or U12029 (N_12029,N_11054,N_11425);
and U12030 (N_12030,N_11918,N_11564);
nand U12031 (N_12031,N_11325,N_11035);
and U12032 (N_12032,N_11999,N_11939);
or U12033 (N_12033,N_11205,N_11444);
or U12034 (N_12034,N_11845,N_11375);
nand U12035 (N_12035,N_11297,N_11242);
and U12036 (N_12036,N_11156,N_11744);
nand U12037 (N_12037,N_11345,N_11754);
nor U12038 (N_12038,N_11025,N_11426);
or U12039 (N_12039,N_11004,N_11111);
nand U12040 (N_12040,N_11370,N_11158);
nand U12041 (N_12041,N_11884,N_11533);
nor U12042 (N_12042,N_11995,N_11066);
xnor U12043 (N_12043,N_11636,N_11921);
nand U12044 (N_12044,N_11616,N_11132);
nand U12045 (N_12045,N_11630,N_11062);
nand U12046 (N_12046,N_11051,N_11312);
and U12047 (N_12047,N_11733,N_11732);
nor U12048 (N_12048,N_11702,N_11949);
and U12049 (N_12049,N_11760,N_11181);
and U12050 (N_12050,N_11730,N_11241);
nor U12051 (N_12051,N_11377,N_11168);
xor U12052 (N_12052,N_11827,N_11130);
xor U12053 (N_12053,N_11087,N_11549);
nand U12054 (N_12054,N_11898,N_11173);
nor U12055 (N_12055,N_11890,N_11886);
nand U12056 (N_12056,N_11547,N_11000);
and U12057 (N_12057,N_11960,N_11617);
or U12058 (N_12058,N_11752,N_11133);
and U12059 (N_12059,N_11053,N_11865);
and U12060 (N_12060,N_11633,N_11488);
nor U12061 (N_12061,N_11327,N_11820);
nor U12062 (N_12062,N_11771,N_11994);
or U12063 (N_12063,N_11008,N_11143);
xor U12064 (N_12064,N_11829,N_11614);
nor U12065 (N_12065,N_11397,N_11296);
xor U12066 (N_12066,N_11235,N_11073);
nor U12067 (N_12067,N_11930,N_11644);
nand U12068 (N_12068,N_11922,N_11094);
and U12069 (N_12069,N_11905,N_11106);
and U12070 (N_12070,N_11575,N_11659);
nand U12071 (N_12071,N_11154,N_11794);
nor U12072 (N_12072,N_11677,N_11531);
or U12073 (N_12073,N_11772,N_11302);
or U12074 (N_12074,N_11650,N_11973);
and U12075 (N_12075,N_11116,N_11590);
nor U12076 (N_12076,N_11576,N_11487);
and U12077 (N_12077,N_11141,N_11037);
nand U12078 (N_12078,N_11322,N_11121);
or U12079 (N_12079,N_11482,N_11331);
nand U12080 (N_12080,N_11613,N_11263);
nor U12081 (N_12081,N_11204,N_11882);
nand U12082 (N_12082,N_11117,N_11822);
and U12083 (N_12083,N_11212,N_11246);
nand U12084 (N_12084,N_11323,N_11202);
nor U12085 (N_12085,N_11854,N_11520);
or U12086 (N_12086,N_11681,N_11027);
or U12087 (N_12087,N_11697,N_11372);
nand U12088 (N_12088,N_11041,N_11095);
nor U12089 (N_12089,N_11099,N_11556);
nor U12090 (N_12090,N_11285,N_11050);
or U12091 (N_12091,N_11226,N_11802);
nor U12092 (N_12092,N_11784,N_11236);
or U12093 (N_12093,N_11413,N_11291);
and U12094 (N_12094,N_11338,N_11321);
or U12095 (N_12095,N_11701,N_11249);
or U12096 (N_12096,N_11398,N_11852);
and U12097 (N_12097,N_11574,N_11180);
xnor U12098 (N_12098,N_11257,N_11265);
nand U12099 (N_12099,N_11596,N_11699);
or U12100 (N_12100,N_11163,N_11252);
nand U12101 (N_12101,N_11347,N_11288);
nor U12102 (N_12102,N_11567,N_11530);
or U12103 (N_12103,N_11023,N_11587);
nand U12104 (N_12104,N_11559,N_11553);
or U12105 (N_12105,N_11303,N_11378);
nor U12106 (N_12106,N_11183,N_11147);
or U12107 (N_12107,N_11198,N_11229);
xnor U12108 (N_12108,N_11072,N_11795);
nor U12109 (N_12109,N_11174,N_11920);
nand U12110 (N_12110,N_11625,N_11390);
or U12111 (N_12111,N_11770,N_11662);
or U12112 (N_12112,N_11766,N_11764);
xor U12113 (N_12113,N_11048,N_11934);
xnor U12114 (N_12114,N_11479,N_11237);
and U12115 (N_12115,N_11527,N_11078);
or U12116 (N_12116,N_11786,N_11534);
and U12117 (N_12117,N_11859,N_11814);
nor U12118 (N_12118,N_11509,N_11821);
xnor U12119 (N_12119,N_11495,N_11649);
and U12120 (N_12120,N_11695,N_11661);
nand U12121 (N_12121,N_11255,N_11127);
nand U12122 (N_12122,N_11669,N_11361);
or U12123 (N_12123,N_11340,N_11476);
or U12124 (N_12124,N_11192,N_11137);
nand U12125 (N_12125,N_11716,N_11935);
nand U12126 (N_12126,N_11963,N_11088);
nand U12127 (N_12127,N_11804,N_11477);
nand U12128 (N_12128,N_11997,N_11196);
or U12129 (N_12129,N_11243,N_11315);
and U12130 (N_12130,N_11683,N_11317);
or U12131 (N_12131,N_11157,N_11401);
nand U12132 (N_12132,N_11857,N_11956);
and U12133 (N_12133,N_11344,N_11735);
xnor U12134 (N_12134,N_11282,N_11416);
and U12135 (N_12135,N_11694,N_11684);
nor U12136 (N_12136,N_11581,N_11739);
xnor U12137 (N_12137,N_11670,N_11194);
nand U12138 (N_12138,N_11091,N_11266);
or U12139 (N_12139,N_11366,N_11188);
nor U12140 (N_12140,N_11562,N_11367);
nor U12141 (N_12141,N_11672,N_11319);
nand U12142 (N_12142,N_11887,N_11337);
xor U12143 (N_12143,N_11436,N_11809);
nand U12144 (N_12144,N_11463,N_11199);
nor U12145 (N_12145,N_11492,N_11467);
nor U12146 (N_12146,N_11295,N_11743);
nand U12147 (N_12147,N_11261,N_11863);
and U12148 (N_12148,N_11368,N_11902);
nand U12149 (N_12149,N_11641,N_11640);
nor U12150 (N_12150,N_11819,N_11706);
or U12151 (N_12151,N_11334,N_11060);
nor U12152 (N_12152,N_11069,N_11594);
nand U12153 (N_12153,N_11365,N_11404);
xor U12154 (N_12154,N_11805,N_11832);
nand U12155 (N_12155,N_11992,N_11500);
nand U12156 (N_12156,N_11548,N_11271);
or U12157 (N_12157,N_11592,N_11565);
nand U12158 (N_12158,N_11421,N_11234);
xnor U12159 (N_12159,N_11287,N_11167);
or U12160 (N_12160,N_11359,N_11191);
nor U12161 (N_12161,N_11042,N_11799);
xnor U12162 (N_12162,N_11729,N_11248);
and U12163 (N_12163,N_11273,N_11688);
nor U12164 (N_12164,N_11864,N_11709);
nand U12165 (N_12165,N_11171,N_11775);
or U12166 (N_12166,N_11776,N_11823);
or U12167 (N_12167,N_11708,N_11244);
xor U12168 (N_12168,N_11270,N_11653);
and U12169 (N_12169,N_11406,N_11923);
or U12170 (N_12170,N_11810,N_11536);
or U12171 (N_12171,N_11676,N_11742);
xnor U12172 (N_12172,N_11703,N_11705);
nor U12173 (N_12173,N_11057,N_11018);
xor U12174 (N_12174,N_11113,N_11120);
nor U12175 (N_12175,N_11988,N_11203);
or U12176 (N_12176,N_11635,N_11873);
or U12177 (N_12177,N_11431,N_11881);
nand U12178 (N_12178,N_11101,N_11901);
nor U12179 (N_12179,N_11746,N_11400);
and U12180 (N_12180,N_11507,N_11895);
nand U12181 (N_12181,N_11335,N_11726);
and U12182 (N_12182,N_11542,N_11622);
or U12183 (N_12183,N_11712,N_11686);
nor U12184 (N_12184,N_11588,N_11351);
nand U12185 (N_12185,N_11429,N_11318);
nor U12186 (N_12186,N_11478,N_11142);
and U12187 (N_12187,N_11409,N_11301);
nor U12188 (N_12188,N_11720,N_11842);
and U12189 (N_12189,N_11017,N_11457);
nand U12190 (N_12190,N_11358,N_11233);
or U12191 (N_12191,N_11501,N_11666);
and U12192 (N_12192,N_11721,N_11658);
xor U12193 (N_12193,N_11209,N_11981);
and U12194 (N_12194,N_11806,N_11001);
nor U12195 (N_12195,N_11755,N_11352);
nor U12196 (N_12196,N_11355,N_11719);
xor U12197 (N_12197,N_11830,N_11418);
or U12198 (N_12198,N_11014,N_11208);
or U12199 (N_12199,N_11029,N_11153);
and U12200 (N_12200,N_11262,N_11349);
nor U12201 (N_12201,N_11521,N_11971);
and U12202 (N_12202,N_11947,N_11129);
or U12203 (N_12203,N_11399,N_11184);
nor U12204 (N_12204,N_11936,N_11395);
and U12205 (N_12205,N_11668,N_11128);
xnor U12206 (N_12206,N_11454,N_11433);
xor U12207 (N_12207,N_11460,N_11535);
nor U12208 (N_12208,N_11189,N_11748);
nand U12209 (N_12209,N_11554,N_11675);
nor U12210 (N_12210,N_11987,N_11928);
and U12211 (N_12211,N_11186,N_11269);
nand U12212 (N_12212,N_11778,N_11290);
nand U12213 (N_12213,N_11734,N_11580);
or U12214 (N_12214,N_11959,N_11462);
and U12215 (N_12215,N_11278,N_11505);
or U12216 (N_12216,N_11837,N_11655);
and U12217 (N_12217,N_11889,N_11240);
nor U12218 (N_12218,N_11443,N_11245);
or U12219 (N_12219,N_11591,N_11996);
and U12220 (N_12220,N_11508,N_11678);
nand U12221 (N_12221,N_11532,N_11063);
nor U12222 (N_12222,N_11552,N_11516);
or U12223 (N_12223,N_11761,N_11038);
nor U12224 (N_12224,N_11777,N_11951);
and U12225 (N_12225,N_11298,N_11356);
or U12226 (N_12226,N_11757,N_11558);
xor U12227 (N_12227,N_11439,N_11131);
and U12228 (N_12228,N_11931,N_11305);
nand U12229 (N_12229,N_11145,N_11251);
or U12230 (N_12230,N_11159,N_11108);
nand U12231 (N_12231,N_11496,N_11354);
nor U12232 (N_12232,N_11888,N_11224);
xor U12233 (N_12233,N_11660,N_11470);
xnor U12234 (N_12234,N_11780,N_11568);
and U12235 (N_12235,N_11115,N_11059);
or U12236 (N_12236,N_11774,N_11138);
nor U12237 (N_12237,N_11689,N_11392);
or U12238 (N_12238,N_11541,N_11862);
nor U12239 (N_12239,N_11911,N_11982);
xnor U12240 (N_12240,N_11007,N_11910);
and U12241 (N_12241,N_11172,N_11148);
nand U12242 (N_12242,N_11450,N_11028);
nand U12243 (N_12243,N_11071,N_11459);
nor U12244 (N_12244,N_11441,N_11779);
nor U12245 (N_12245,N_11637,N_11950);
nand U12246 (N_12246,N_11006,N_11308);
nor U12247 (N_12247,N_11741,N_11872);
or U12248 (N_12248,N_11220,N_11110);
or U12249 (N_12249,N_11214,N_11283);
or U12250 (N_12250,N_11903,N_11207);
or U12251 (N_12251,N_11933,N_11586);
and U12252 (N_12252,N_11976,N_11628);
and U12253 (N_12253,N_11798,N_11092);
and U12254 (N_12254,N_11573,N_11506);
or U12255 (N_12255,N_11634,N_11304);
and U12256 (N_12256,N_11948,N_11942);
nor U12257 (N_12257,N_11696,N_11396);
or U12258 (N_12258,N_11466,N_11908);
nand U12259 (N_12259,N_11891,N_11281);
nand U12260 (N_12260,N_11750,N_11497);
nor U12261 (N_12261,N_11169,N_11685);
nor U12262 (N_12262,N_11753,N_11624);
nor U12263 (N_12263,N_11449,N_11494);
nor U12264 (N_12264,N_11844,N_11333);
and U12265 (N_12265,N_11387,N_11510);
nor U12266 (N_12266,N_11084,N_11190);
nand U12267 (N_12267,N_11118,N_11577);
or U12268 (N_12268,N_11728,N_11700);
nor U12269 (N_12269,N_11022,N_11216);
or U12270 (N_12270,N_11136,N_11858);
or U12271 (N_12271,N_11807,N_11943);
nand U12272 (N_12272,N_11098,N_11277);
nor U12273 (N_12273,N_11484,N_11816);
or U12274 (N_12274,N_11749,N_11112);
or U12275 (N_12275,N_11299,N_11967);
nand U12276 (N_12276,N_11906,N_11074);
and U12277 (N_12277,N_11374,N_11927);
nand U12278 (N_12278,N_11289,N_11346);
nor U12279 (N_12279,N_11773,N_11348);
nor U12280 (N_12280,N_11768,N_11093);
nand U12281 (N_12281,N_11990,N_11268);
and U12282 (N_12282,N_11013,N_11851);
or U12283 (N_12283,N_11639,N_11589);
xnor U12284 (N_12284,N_11643,N_11671);
and U12285 (N_12285,N_11715,N_11808);
or U12286 (N_12286,N_11343,N_11342);
and U12287 (N_12287,N_11293,N_11940);
or U12288 (N_12288,N_11040,N_11945);
or U12289 (N_12289,N_11306,N_11124);
xor U12290 (N_12290,N_11498,N_11061);
nand U12291 (N_12291,N_11788,N_11974);
xor U12292 (N_12292,N_11598,N_11430);
or U12293 (N_12293,N_11079,N_11543);
or U12294 (N_12294,N_11440,N_11718);
nor U12295 (N_12295,N_11915,N_11525);
or U12296 (N_12296,N_11893,N_11020);
xor U12297 (N_12297,N_11885,N_11123);
nor U12298 (N_12298,N_11892,N_11201);
and U12299 (N_12299,N_11691,N_11612);
and U12300 (N_12300,N_11875,N_11966);
nor U12301 (N_12301,N_11026,N_11272);
nand U12302 (N_12302,N_11503,N_11919);
nand U12303 (N_12303,N_11916,N_11731);
or U12304 (N_12304,N_11824,N_11593);
nand U12305 (N_12305,N_11899,N_11941);
or U12306 (N_12306,N_11605,N_11572);
or U12307 (N_12307,N_11968,N_11031);
or U12308 (N_12308,N_11944,N_11274);
or U12309 (N_12309,N_11693,N_11360);
nand U12310 (N_12310,N_11504,N_11314);
or U12311 (N_12311,N_11489,N_11002);
nand U12312 (N_12312,N_11597,N_11738);
and U12313 (N_12313,N_11329,N_11292);
nand U12314 (N_12314,N_11557,N_11239);
nor U12315 (N_12315,N_11871,N_11818);
nand U12316 (N_12316,N_11664,N_11538);
nor U12317 (N_12317,N_11332,N_11600);
nand U12318 (N_12318,N_11511,N_11985);
or U12319 (N_12319,N_11284,N_11067);
or U12320 (N_12320,N_11044,N_11896);
nor U12321 (N_12321,N_11610,N_11096);
or U12322 (N_12322,N_11213,N_11330);
or U12323 (N_12323,N_11386,N_11369);
nand U12324 (N_12324,N_11642,N_11980);
nor U12325 (N_12325,N_11075,N_11599);
and U12326 (N_12326,N_11646,N_11009);
nor U12327 (N_12327,N_11583,N_11256);
nor U12328 (N_12328,N_11468,N_11870);
nor U12329 (N_12329,N_11162,N_11550);
or U12330 (N_12330,N_11841,N_11490);
nor U12331 (N_12331,N_11371,N_11964);
and U12332 (N_12332,N_11221,N_11912);
nor U12333 (N_12333,N_11144,N_11657);
or U12334 (N_12334,N_11579,N_11638);
or U12335 (N_12335,N_11187,N_11894);
or U12336 (N_12336,N_11182,N_11403);
and U12337 (N_12337,N_11682,N_11667);
and U12338 (N_12338,N_11914,N_11611);
and U12339 (N_12339,N_11647,N_11193);
nand U12340 (N_12340,N_11326,N_11725);
and U12341 (N_12341,N_11517,N_11817);
or U12342 (N_12342,N_11247,N_11623);
and U12343 (N_12343,N_11789,N_11310);
and U12344 (N_12344,N_11019,N_11876);
nand U12345 (N_12345,N_11179,N_11979);
nand U12346 (N_12346,N_11801,N_11765);
or U12347 (N_12347,N_11522,N_11077);
and U12348 (N_12348,N_11279,N_11227);
and U12349 (N_12349,N_11453,N_11139);
nand U12350 (N_12350,N_11491,N_11472);
nor U12351 (N_12351,N_11710,N_11926);
or U12352 (N_12352,N_11843,N_11336);
nor U12353 (N_12353,N_11197,N_11714);
and U12354 (N_12354,N_11740,N_11631);
or U12355 (N_12355,N_11151,N_11632);
nand U12356 (N_12356,N_11724,N_11796);
nor U12357 (N_12357,N_11140,N_11217);
and U12358 (N_12358,N_11146,N_11977);
nor U12359 (N_12359,N_11698,N_11465);
nor U12360 (N_12360,N_11620,N_11972);
nor U12361 (N_12361,N_11962,N_11656);
and U12362 (N_12362,N_11428,N_11253);
nand U12363 (N_12363,N_11086,N_11736);
nand U12364 (N_12364,N_11104,N_11280);
and U12365 (N_12365,N_11480,N_11388);
nor U12366 (N_12366,N_11380,N_11161);
nor U12367 (N_12367,N_11381,N_11602);
xnor U12368 (N_12368,N_11135,N_11058);
nor U12369 (N_12369,N_11834,N_11383);
nor U12370 (N_12370,N_11989,N_11411);
or U12371 (N_12371,N_11907,N_11405);
and U12372 (N_12372,N_11518,N_11003);
xnor U12373 (N_12373,N_11606,N_11607);
xor U12374 (N_12374,N_11645,N_11230);
and U12375 (N_12375,N_11540,N_11566);
nand U12376 (N_12376,N_11866,N_11563);
or U12377 (N_12377,N_11011,N_11601);
nor U12378 (N_12378,N_11102,N_11047);
or U12379 (N_12379,N_11176,N_11555);
nand U12380 (N_12380,N_11578,N_11869);
nand U12381 (N_12381,N_11357,N_11582);
nand U12382 (N_12382,N_11957,N_11673);
nor U12383 (N_12383,N_11847,N_11758);
nor U12384 (N_12384,N_11762,N_11978);
and U12385 (N_12385,N_11690,N_11065);
xor U12386 (N_12386,N_11438,N_11134);
nand U12387 (N_12387,N_11122,N_11791);
or U12388 (N_12388,N_11692,N_11185);
and U12389 (N_12389,N_11983,N_11385);
or U12390 (N_12390,N_11473,N_11276);
or U12391 (N_12391,N_11417,N_11456);
xor U12392 (N_12392,N_11603,N_11998);
nand U12393 (N_12393,N_11464,N_11455);
nand U12394 (N_12394,N_11993,N_11604);
nor U12395 (N_12395,N_11674,N_11946);
nor U12396 (N_12396,N_11727,N_11561);
nor U12397 (N_12397,N_11502,N_11307);
nand U12398 (N_12398,N_11419,N_11149);
and U12399 (N_12399,N_11427,N_11056);
nand U12400 (N_12400,N_11868,N_11961);
nor U12401 (N_12401,N_11382,N_11422);
and U12402 (N_12402,N_11379,N_11840);
and U12403 (N_12403,N_11394,N_11415);
or U12404 (N_12404,N_11223,N_11737);
or U12405 (N_12405,N_11448,N_11469);
and U12406 (N_12406,N_11036,N_11759);
nand U12407 (N_12407,N_11175,N_11238);
and U12408 (N_12408,N_11783,N_11909);
or U12409 (N_12409,N_11015,N_11984);
or U12410 (N_12410,N_11585,N_11309);
nor U12411 (N_12411,N_11717,N_11679);
xor U12412 (N_12412,N_11654,N_11619);
or U12413 (N_12413,N_11178,N_11320);
nor U12414 (N_12414,N_11537,N_11166);
nor U12415 (N_12415,N_11813,N_11849);
and U12416 (N_12416,N_11648,N_11107);
or U12417 (N_12417,N_11049,N_11855);
and U12418 (N_12418,N_11021,N_11751);
or U12419 (N_12419,N_11211,N_11826);
nor U12420 (N_12420,N_11514,N_11076);
or U12421 (N_12421,N_11493,N_11811);
xor U12422 (N_12422,N_11210,N_11033);
nor U12423 (N_12423,N_11408,N_11445);
and U12424 (N_12424,N_11471,N_11609);
xnor U12425 (N_12425,N_11225,N_11932);
nor U12426 (N_12426,N_11867,N_11259);
and U12427 (N_12427,N_11782,N_11797);
nor U12428 (N_12428,N_11781,N_11787);
nand U12429 (N_12429,N_11165,N_11680);
nand U12430 (N_12430,N_11170,N_11446);
nor U12431 (N_12431,N_11707,N_11952);
or U12432 (N_12432,N_11384,N_11039);
nor U12433 (N_12433,N_11010,N_11584);
nand U12434 (N_12434,N_11570,N_11085);
xnor U12435 (N_12435,N_11767,N_11621);
nand U12436 (N_12436,N_11081,N_11005);
or U12437 (N_12437,N_11860,N_11515);
nor U12438 (N_12438,N_11970,N_11713);
and U12439 (N_12439,N_11747,N_11711);
nand U12440 (N_12440,N_11792,N_11831);
or U12441 (N_12441,N_11451,N_11434);
and U12442 (N_12442,N_11177,N_11499);
nand U12443 (N_12443,N_11090,N_11420);
nand U12444 (N_12444,N_11745,N_11363);
and U12445 (N_12445,N_11032,N_11763);
and U12446 (N_12446,N_11339,N_11070);
nand U12447 (N_12447,N_11447,N_11975);
nor U12448 (N_12448,N_11722,N_11793);
or U12449 (N_12449,N_11545,N_11424);
or U12450 (N_12450,N_11704,N_11353);
and U12451 (N_12451,N_11652,N_11350);
nand U12452 (N_12452,N_11152,N_11475);
or U12453 (N_12453,N_11560,N_11595);
or U12454 (N_12454,N_11848,N_11608);
nor U12455 (N_12455,N_11519,N_11756);
or U12456 (N_12456,N_11615,N_11206);
nand U12457 (N_12457,N_11105,N_11218);
nand U12458 (N_12458,N_11815,N_11407);
nand U12459 (N_12459,N_11089,N_11929);
or U12460 (N_12460,N_11569,N_11924);
and U12461 (N_12461,N_11529,N_11986);
nor U12462 (N_12462,N_11769,N_11119);
nor U12463 (N_12463,N_11046,N_11432);
and U12464 (N_12464,N_11264,N_11812);
and U12465 (N_12465,N_11232,N_11954);
and U12466 (N_12466,N_11833,N_11402);
nand U12467 (N_12467,N_11938,N_11024);
nor U12468 (N_12468,N_11512,N_11412);
nand U12469 (N_12469,N_11080,N_11286);
or U12470 (N_12470,N_11626,N_11523);
nor U12471 (N_12471,N_11012,N_11900);
nand U12472 (N_12472,N_11389,N_11267);
nand U12473 (N_12473,N_11442,N_11629);
nand U12474 (N_12474,N_11663,N_11836);
or U12475 (N_12475,N_11539,N_11925);
nand U12476 (N_12476,N_11627,N_11878);
nand U12477 (N_12477,N_11125,N_11879);
nor U12478 (N_12478,N_11785,N_11917);
nor U12479 (N_12479,N_11294,N_11825);
or U12480 (N_12480,N_11528,N_11474);
and U12481 (N_12481,N_11393,N_11109);
and U12482 (N_12482,N_11965,N_11100);
nand U12483 (N_12483,N_11874,N_11414);
or U12484 (N_12484,N_11571,N_11937);
or U12485 (N_12485,N_11258,N_11461);
or U12486 (N_12486,N_11526,N_11160);
nand U12487 (N_12487,N_11861,N_11376);
nor U12488 (N_12488,N_11362,N_11483);
or U12489 (N_12489,N_11328,N_11260);
or U12490 (N_12490,N_11341,N_11665);
or U12491 (N_12491,N_11828,N_11853);
and U12492 (N_12492,N_11513,N_11300);
nor U12493 (N_12493,N_11064,N_11524);
and U12494 (N_12494,N_11222,N_11856);
xnor U12495 (N_12495,N_11423,N_11311);
and U12496 (N_12496,N_11969,N_11838);
and U12497 (N_12497,N_11083,N_11324);
and U12498 (N_12498,N_11231,N_11839);
and U12499 (N_12499,N_11250,N_11452);
xor U12500 (N_12500,N_11214,N_11554);
xor U12501 (N_12501,N_11139,N_11192);
and U12502 (N_12502,N_11346,N_11524);
nor U12503 (N_12503,N_11792,N_11038);
or U12504 (N_12504,N_11728,N_11759);
and U12505 (N_12505,N_11220,N_11786);
and U12506 (N_12506,N_11372,N_11063);
nand U12507 (N_12507,N_11006,N_11863);
and U12508 (N_12508,N_11205,N_11437);
xor U12509 (N_12509,N_11133,N_11955);
and U12510 (N_12510,N_11544,N_11094);
nor U12511 (N_12511,N_11377,N_11539);
nand U12512 (N_12512,N_11242,N_11665);
and U12513 (N_12513,N_11303,N_11400);
nand U12514 (N_12514,N_11308,N_11658);
and U12515 (N_12515,N_11250,N_11086);
nor U12516 (N_12516,N_11510,N_11826);
nand U12517 (N_12517,N_11557,N_11984);
nor U12518 (N_12518,N_11477,N_11613);
nand U12519 (N_12519,N_11037,N_11845);
nor U12520 (N_12520,N_11940,N_11263);
and U12521 (N_12521,N_11144,N_11264);
and U12522 (N_12522,N_11424,N_11951);
or U12523 (N_12523,N_11950,N_11917);
nor U12524 (N_12524,N_11726,N_11076);
or U12525 (N_12525,N_11537,N_11618);
nand U12526 (N_12526,N_11664,N_11871);
nor U12527 (N_12527,N_11276,N_11751);
nand U12528 (N_12528,N_11644,N_11420);
nand U12529 (N_12529,N_11008,N_11022);
or U12530 (N_12530,N_11913,N_11851);
nor U12531 (N_12531,N_11879,N_11200);
or U12532 (N_12532,N_11471,N_11213);
nor U12533 (N_12533,N_11633,N_11788);
and U12534 (N_12534,N_11588,N_11183);
nor U12535 (N_12535,N_11083,N_11817);
or U12536 (N_12536,N_11331,N_11534);
nand U12537 (N_12537,N_11789,N_11203);
and U12538 (N_12538,N_11022,N_11838);
xnor U12539 (N_12539,N_11783,N_11646);
and U12540 (N_12540,N_11079,N_11516);
and U12541 (N_12541,N_11153,N_11134);
and U12542 (N_12542,N_11628,N_11824);
nor U12543 (N_12543,N_11055,N_11933);
and U12544 (N_12544,N_11960,N_11505);
and U12545 (N_12545,N_11195,N_11249);
nor U12546 (N_12546,N_11362,N_11122);
and U12547 (N_12547,N_11942,N_11826);
or U12548 (N_12548,N_11939,N_11769);
and U12549 (N_12549,N_11132,N_11746);
or U12550 (N_12550,N_11571,N_11995);
and U12551 (N_12551,N_11488,N_11413);
and U12552 (N_12552,N_11903,N_11746);
xnor U12553 (N_12553,N_11482,N_11081);
nand U12554 (N_12554,N_11777,N_11812);
and U12555 (N_12555,N_11765,N_11615);
nor U12556 (N_12556,N_11253,N_11487);
nor U12557 (N_12557,N_11577,N_11673);
nand U12558 (N_12558,N_11848,N_11793);
nand U12559 (N_12559,N_11986,N_11465);
nand U12560 (N_12560,N_11643,N_11982);
or U12561 (N_12561,N_11474,N_11499);
xnor U12562 (N_12562,N_11680,N_11403);
nor U12563 (N_12563,N_11408,N_11102);
or U12564 (N_12564,N_11398,N_11249);
nand U12565 (N_12565,N_11087,N_11018);
or U12566 (N_12566,N_11689,N_11342);
nand U12567 (N_12567,N_11345,N_11455);
and U12568 (N_12568,N_11947,N_11510);
or U12569 (N_12569,N_11661,N_11584);
nand U12570 (N_12570,N_11748,N_11347);
or U12571 (N_12571,N_11255,N_11418);
nor U12572 (N_12572,N_11373,N_11290);
xnor U12573 (N_12573,N_11293,N_11342);
or U12574 (N_12574,N_11711,N_11254);
nand U12575 (N_12575,N_11443,N_11622);
nor U12576 (N_12576,N_11680,N_11850);
nor U12577 (N_12577,N_11693,N_11802);
nand U12578 (N_12578,N_11099,N_11203);
nand U12579 (N_12579,N_11885,N_11245);
nor U12580 (N_12580,N_11142,N_11362);
nor U12581 (N_12581,N_11704,N_11364);
or U12582 (N_12582,N_11726,N_11245);
and U12583 (N_12583,N_11958,N_11065);
nor U12584 (N_12584,N_11187,N_11107);
and U12585 (N_12585,N_11283,N_11220);
xor U12586 (N_12586,N_11110,N_11107);
and U12587 (N_12587,N_11450,N_11792);
nand U12588 (N_12588,N_11106,N_11767);
xnor U12589 (N_12589,N_11543,N_11039);
xnor U12590 (N_12590,N_11872,N_11415);
nor U12591 (N_12591,N_11925,N_11082);
nor U12592 (N_12592,N_11297,N_11809);
and U12593 (N_12593,N_11399,N_11332);
nand U12594 (N_12594,N_11483,N_11897);
nor U12595 (N_12595,N_11348,N_11137);
nand U12596 (N_12596,N_11254,N_11707);
nor U12597 (N_12597,N_11546,N_11095);
nand U12598 (N_12598,N_11040,N_11809);
xnor U12599 (N_12599,N_11417,N_11735);
nand U12600 (N_12600,N_11085,N_11996);
nand U12601 (N_12601,N_11117,N_11724);
or U12602 (N_12602,N_11842,N_11237);
nor U12603 (N_12603,N_11419,N_11389);
nor U12604 (N_12604,N_11110,N_11137);
and U12605 (N_12605,N_11157,N_11920);
nand U12606 (N_12606,N_11302,N_11154);
nand U12607 (N_12607,N_11276,N_11971);
or U12608 (N_12608,N_11652,N_11588);
nor U12609 (N_12609,N_11957,N_11305);
nor U12610 (N_12610,N_11220,N_11572);
or U12611 (N_12611,N_11498,N_11664);
or U12612 (N_12612,N_11053,N_11597);
and U12613 (N_12613,N_11674,N_11168);
xnor U12614 (N_12614,N_11719,N_11361);
and U12615 (N_12615,N_11573,N_11625);
and U12616 (N_12616,N_11966,N_11558);
xor U12617 (N_12617,N_11866,N_11755);
or U12618 (N_12618,N_11584,N_11518);
nor U12619 (N_12619,N_11317,N_11549);
nor U12620 (N_12620,N_11903,N_11537);
and U12621 (N_12621,N_11354,N_11261);
nand U12622 (N_12622,N_11743,N_11368);
or U12623 (N_12623,N_11648,N_11099);
nand U12624 (N_12624,N_11679,N_11554);
nor U12625 (N_12625,N_11801,N_11193);
or U12626 (N_12626,N_11496,N_11337);
and U12627 (N_12627,N_11677,N_11105);
xnor U12628 (N_12628,N_11027,N_11581);
nor U12629 (N_12629,N_11882,N_11847);
and U12630 (N_12630,N_11313,N_11707);
nand U12631 (N_12631,N_11182,N_11015);
or U12632 (N_12632,N_11608,N_11722);
nor U12633 (N_12633,N_11585,N_11936);
xor U12634 (N_12634,N_11193,N_11913);
nor U12635 (N_12635,N_11603,N_11449);
nor U12636 (N_12636,N_11038,N_11646);
xnor U12637 (N_12637,N_11723,N_11400);
and U12638 (N_12638,N_11011,N_11562);
nor U12639 (N_12639,N_11666,N_11650);
xor U12640 (N_12640,N_11778,N_11246);
nor U12641 (N_12641,N_11330,N_11491);
or U12642 (N_12642,N_11598,N_11440);
xor U12643 (N_12643,N_11431,N_11140);
and U12644 (N_12644,N_11131,N_11782);
and U12645 (N_12645,N_11049,N_11668);
nor U12646 (N_12646,N_11086,N_11585);
and U12647 (N_12647,N_11200,N_11824);
xor U12648 (N_12648,N_11476,N_11096);
and U12649 (N_12649,N_11281,N_11945);
nand U12650 (N_12650,N_11393,N_11265);
or U12651 (N_12651,N_11886,N_11327);
xnor U12652 (N_12652,N_11042,N_11205);
nand U12653 (N_12653,N_11545,N_11266);
xor U12654 (N_12654,N_11005,N_11746);
or U12655 (N_12655,N_11741,N_11873);
and U12656 (N_12656,N_11354,N_11716);
nand U12657 (N_12657,N_11141,N_11460);
or U12658 (N_12658,N_11299,N_11525);
nor U12659 (N_12659,N_11136,N_11333);
nand U12660 (N_12660,N_11478,N_11905);
nor U12661 (N_12661,N_11911,N_11545);
nor U12662 (N_12662,N_11759,N_11977);
nor U12663 (N_12663,N_11250,N_11606);
or U12664 (N_12664,N_11277,N_11804);
and U12665 (N_12665,N_11059,N_11140);
and U12666 (N_12666,N_11335,N_11975);
nor U12667 (N_12667,N_11596,N_11044);
nor U12668 (N_12668,N_11632,N_11295);
nor U12669 (N_12669,N_11850,N_11408);
and U12670 (N_12670,N_11519,N_11508);
or U12671 (N_12671,N_11976,N_11179);
or U12672 (N_12672,N_11705,N_11026);
and U12673 (N_12673,N_11003,N_11517);
nor U12674 (N_12674,N_11699,N_11886);
nor U12675 (N_12675,N_11045,N_11326);
nand U12676 (N_12676,N_11479,N_11332);
xnor U12677 (N_12677,N_11816,N_11048);
and U12678 (N_12678,N_11263,N_11638);
or U12679 (N_12679,N_11643,N_11171);
nor U12680 (N_12680,N_11051,N_11943);
or U12681 (N_12681,N_11500,N_11815);
and U12682 (N_12682,N_11619,N_11055);
nand U12683 (N_12683,N_11633,N_11174);
nor U12684 (N_12684,N_11944,N_11540);
xor U12685 (N_12685,N_11895,N_11334);
nor U12686 (N_12686,N_11395,N_11459);
and U12687 (N_12687,N_11284,N_11717);
nor U12688 (N_12688,N_11246,N_11621);
and U12689 (N_12689,N_11122,N_11871);
nor U12690 (N_12690,N_11692,N_11913);
or U12691 (N_12691,N_11351,N_11485);
nor U12692 (N_12692,N_11460,N_11099);
xnor U12693 (N_12693,N_11224,N_11469);
nand U12694 (N_12694,N_11002,N_11150);
nand U12695 (N_12695,N_11345,N_11923);
nand U12696 (N_12696,N_11133,N_11390);
nor U12697 (N_12697,N_11377,N_11892);
nor U12698 (N_12698,N_11631,N_11557);
nand U12699 (N_12699,N_11285,N_11199);
and U12700 (N_12700,N_11480,N_11927);
nand U12701 (N_12701,N_11681,N_11320);
nor U12702 (N_12702,N_11377,N_11870);
or U12703 (N_12703,N_11818,N_11974);
and U12704 (N_12704,N_11112,N_11791);
nand U12705 (N_12705,N_11084,N_11928);
xnor U12706 (N_12706,N_11244,N_11028);
nor U12707 (N_12707,N_11553,N_11645);
or U12708 (N_12708,N_11796,N_11101);
or U12709 (N_12709,N_11300,N_11524);
nor U12710 (N_12710,N_11220,N_11350);
or U12711 (N_12711,N_11612,N_11083);
and U12712 (N_12712,N_11832,N_11347);
nand U12713 (N_12713,N_11888,N_11194);
or U12714 (N_12714,N_11852,N_11858);
nand U12715 (N_12715,N_11985,N_11907);
nor U12716 (N_12716,N_11559,N_11992);
and U12717 (N_12717,N_11630,N_11524);
nand U12718 (N_12718,N_11619,N_11865);
nor U12719 (N_12719,N_11280,N_11915);
or U12720 (N_12720,N_11903,N_11529);
and U12721 (N_12721,N_11773,N_11583);
xor U12722 (N_12722,N_11672,N_11225);
or U12723 (N_12723,N_11041,N_11911);
nand U12724 (N_12724,N_11071,N_11584);
or U12725 (N_12725,N_11101,N_11370);
nor U12726 (N_12726,N_11536,N_11306);
nor U12727 (N_12727,N_11839,N_11613);
or U12728 (N_12728,N_11709,N_11648);
nor U12729 (N_12729,N_11733,N_11241);
and U12730 (N_12730,N_11417,N_11991);
and U12731 (N_12731,N_11881,N_11290);
nand U12732 (N_12732,N_11356,N_11434);
and U12733 (N_12733,N_11973,N_11166);
nor U12734 (N_12734,N_11999,N_11175);
and U12735 (N_12735,N_11170,N_11335);
xnor U12736 (N_12736,N_11796,N_11006);
and U12737 (N_12737,N_11732,N_11076);
xnor U12738 (N_12738,N_11502,N_11412);
nor U12739 (N_12739,N_11781,N_11914);
nor U12740 (N_12740,N_11227,N_11904);
nor U12741 (N_12741,N_11992,N_11083);
nand U12742 (N_12742,N_11490,N_11007);
nor U12743 (N_12743,N_11058,N_11475);
nand U12744 (N_12744,N_11964,N_11451);
nor U12745 (N_12745,N_11963,N_11789);
and U12746 (N_12746,N_11636,N_11403);
and U12747 (N_12747,N_11088,N_11821);
or U12748 (N_12748,N_11117,N_11180);
xnor U12749 (N_12749,N_11299,N_11759);
nand U12750 (N_12750,N_11407,N_11277);
nor U12751 (N_12751,N_11803,N_11494);
or U12752 (N_12752,N_11236,N_11057);
nor U12753 (N_12753,N_11631,N_11533);
and U12754 (N_12754,N_11296,N_11399);
or U12755 (N_12755,N_11010,N_11479);
nand U12756 (N_12756,N_11361,N_11390);
nor U12757 (N_12757,N_11371,N_11412);
and U12758 (N_12758,N_11101,N_11728);
or U12759 (N_12759,N_11903,N_11390);
nor U12760 (N_12760,N_11438,N_11573);
nand U12761 (N_12761,N_11687,N_11385);
nor U12762 (N_12762,N_11450,N_11262);
nor U12763 (N_12763,N_11770,N_11629);
nor U12764 (N_12764,N_11939,N_11269);
and U12765 (N_12765,N_11521,N_11082);
nand U12766 (N_12766,N_11360,N_11774);
nor U12767 (N_12767,N_11500,N_11238);
and U12768 (N_12768,N_11046,N_11874);
nand U12769 (N_12769,N_11108,N_11254);
nand U12770 (N_12770,N_11570,N_11494);
and U12771 (N_12771,N_11728,N_11182);
xnor U12772 (N_12772,N_11504,N_11693);
or U12773 (N_12773,N_11619,N_11264);
and U12774 (N_12774,N_11841,N_11224);
nor U12775 (N_12775,N_11832,N_11432);
or U12776 (N_12776,N_11731,N_11027);
nor U12777 (N_12777,N_11565,N_11726);
nand U12778 (N_12778,N_11828,N_11793);
or U12779 (N_12779,N_11190,N_11865);
or U12780 (N_12780,N_11991,N_11332);
nor U12781 (N_12781,N_11889,N_11276);
or U12782 (N_12782,N_11838,N_11057);
or U12783 (N_12783,N_11345,N_11049);
or U12784 (N_12784,N_11515,N_11867);
or U12785 (N_12785,N_11068,N_11628);
or U12786 (N_12786,N_11410,N_11950);
and U12787 (N_12787,N_11271,N_11072);
and U12788 (N_12788,N_11092,N_11702);
or U12789 (N_12789,N_11228,N_11591);
xnor U12790 (N_12790,N_11244,N_11410);
nor U12791 (N_12791,N_11345,N_11949);
nand U12792 (N_12792,N_11993,N_11836);
or U12793 (N_12793,N_11986,N_11460);
or U12794 (N_12794,N_11606,N_11729);
nand U12795 (N_12795,N_11548,N_11340);
and U12796 (N_12796,N_11833,N_11071);
nand U12797 (N_12797,N_11330,N_11322);
nor U12798 (N_12798,N_11213,N_11546);
and U12799 (N_12799,N_11575,N_11217);
nand U12800 (N_12800,N_11137,N_11638);
or U12801 (N_12801,N_11283,N_11535);
nor U12802 (N_12802,N_11002,N_11263);
and U12803 (N_12803,N_11222,N_11718);
or U12804 (N_12804,N_11590,N_11324);
nor U12805 (N_12805,N_11585,N_11921);
nor U12806 (N_12806,N_11867,N_11740);
nand U12807 (N_12807,N_11145,N_11545);
nand U12808 (N_12808,N_11761,N_11758);
and U12809 (N_12809,N_11550,N_11873);
nor U12810 (N_12810,N_11425,N_11169);
or U12811 (N_12811,N_11177,N_11878);
nor U12812 (N_12812,N_11371,N_11402);
nor U12813 (N_12813,N_11218,N_11804);
and U12814 (N_12814,N_11335,N_11077);
and U12815 (N_12815,N_11257,N_11281);
nand U12816 (N_12816,N_11054,N_11846);
or U12817 (N_12817,N_11099,N_11036);
or U12818 (N_12818,N_11098,N_11535);
nor U12819 (N_12819,N_11941,N_11393);
nand U12820 (N_12820,N_11325,N_11227);
nand U12821 (N_12821,N_11827,N_11276);
nor U12822 (N_12822,N_11443,N_11441);
xnor U12823 (N_12823,N_11050,N_11735);
nand U12824 (N_12824,N_11960,N_11893);
nor U12825 (N_12825,N_11784,N_11047);
nand U12826 (N_12826,N_11036,N_11383);
and U12827 (N_12827,N_11387,N_11350);
xor U12828 (N_12828,N_11344,N_11414);
and U12829 (N_12829,N_11636,N_11081);
nor U12830 (N_12830,N_11301,N_11709);
nand U12831 (N_12831,N_11605,N_11464);
or U12832 (N_12832,N_11026,N_11962);
nor U12833 (N_12833,N_11805,N_11710);
nor U12834 (N_12834,N_11338,N_11363);
xnor U12835 (N_12835,N_11672,N_11413);
xnor U12836 (N_12836,N_11116,N_11859);
and U12837 (N_12837,N_11637,N_11818);
nand U12838 (N_12838,N_11641,N_11059);
nor U12839 (N_12839,N_11992,N_11908);
and U12840 (N_12840,N_11350,N_11879);
and U12841 (N_12841,N_11782,N_11529);
or U12842 (N_12842,N_11899,N_11871);
or U12843 (N_12843,N_11559,N_11582);
and U12844 (N_12844,N_11083,N_11302);
nor U12845 (N_12845,N_11745,N_11148);
xor U12846 (N_12846,N_11577,N_11319);
nand U12847 (N_12847,N_11936,N_11192);
xor U12848 (N_12848,N_11468,N_11830);
nor U12849 (N_12849,N_11886,N_11817);
and U12850 (N_12850,N_11016,N_11259);
nand U12851 (N_12851,N_11066,N_11432);
nor U12852 (N_12852,N_11034,N_11476);
nor U12853 (N_12853,N_11886,N_11380);
nor U12854 (N_12854,N_11365,N_11038);
xor U12855 (N_12855,N_11255,N_11906);
and U12856 (N_12856,N_11821,N_11657);
nor U12857 (N_12857,N_11733,N_11014);
and U12858 (N_12858,N_11263,N_11791);
and U12859 (N_12859,N_11563,N_11262);
nor U12860 (N_12860,N_11568,N_11075);
or U12861 (N_12861,N_11820,N_11152);
nand U12862 (N_12862,N_11989,N_11902);
nor U12863 (N_12863,N_11254,N_11917);
nand U12864 (N_12864,N_11948,N_11433);
and U12865 (N_12865,N_11632,N_11541);
or U12866 (N_12866,N_11309,N_11419);
nor U12867 (N_12867,N_11527,N_11882);
nand U12868 (N_12868,N_11359,N_11199);
xor U12869 (N_12869,N_11926,N_11259);
nand U12870 (N_12870,N_11794,N_11338);
and U12871 (N_12871,N_11239,N_11208);
or U12872 (N_12872,N_11290,N_11439);
nor U12873 (N_12873,N_11427,N_11486);
nor U12874 (N_12874,N_11550,N_11338);
or U12875 (N_12875,N_11659,N_11851);
and U12876 (N_12876,N_11908,N_11716);
xnor U12877 (N_12877,N_11186,N_11965);
xor U12878 (N_12878,N_11885,N_11796);
and U12879 (N_12879,N_11638,N_11694);
nor U12880 (N_12880,N_11042,N_11660);
nand U12881 (N_12881,N_11998,N_11154);
or U12882 (N_12882,N_11092,N_11423);
or U12883 (N_12883,N_11175,N_11337);
nor U12884 (N_12884,N_11690,N_11391);
and U12885 (N_12885,N_11841,N_11748);
nand U12886 (N_12886,N_11370,N_11904);
nor U12887 (N_12887,N_11002,N_11987);
xnor U12888 (N_12888,N_11507,N_11600);
nand U12889 (N_12889,N_11359,N_11858);
and U12890 (N_12890,N_11829,N_11654);
xnor U12891 (N_12891,N_11857,N_11949);
and U12892 (N_12892,N_11748,N_11183);
xor U12893 (N_12893,N_11883,N_11739);
xnor U12894 (N_12894,N_11993,N_11282);
nor U12895 (N_12895,N_11497,N_11822);
or U12896 (N_12896,N_11070,N_11285);
and U12897 (N_12897,N_11648,N_11130);
or U12898 (N_12898,N_11460,N_11663);
xor U12899 (N_12899,N_11622,N_11835);
nor U12900 (N_12900,N_11652,N_11434);
nor U12901 (N_12901,N_11197,N_11261);
or U12902 (N_12902,N_11199,N_11196);
nor U12903 (N_12903,N_11076,N_11733);
or U12904 (N_12904,N_11083,N_11941);
or U12905 (N_12905,N_11961,N_11523);
and U12906 (N_12906,N_11222,N_11802);
nor U12907 (N_12907,N_11976,N_11509);
nor U12908 (N_12908,N_11316,N_11656);
nor U12909 (N_12909,N_11407,N_11086);
or U12910 (N_12910,N_11776,N_11337);
and U12911 (N_12911,N_11657,N_11386);
nor U12912 (N_12912,N_11883,N_11743);
xnor U12913 (N_12913,N_11033,N_11679);
and U12914 (N_12914,N_11763,N_11292);
nor U12915 (N_12915,N_11677,N_11806);
and U12916 (N_12916,N_11489,N_11536);
nand U12917 (N_12917,N_11370,N_11389);
nand U12918 (N_12918,N_11977,N_11373);
nand U12919 (N_12919,N_11725,N_11129);
or U12920 (N_12920,N_11835,N_11947);
nor U12921 (N_12921,N_11451,N_11521);
nand U12922 (N_12922,N_11690,N_11856);
nand U12923 (N_12923,N_11058,N_11018);
nand U12924 (N_12924,N_11369,N_11977);
or U12925 (N_12925,N_11611,N_11187);
nor U12926 (N_12926,N_11591,N_11440);
or U12927 (N_12927,N_11253,N_11992);
and U12928 (N_12928,N_11621,N_11036);
nand U12929 (N_12929,N_11454,N_11015);
or U12930 (N_12930,N_11912,N_11892);
nor U12931 (N_12931,N_11737,N_11598);
and U12932 (N_12932,N_11628,N_11777);
xnor U12933 (N_12933,N_11773,N_11438);
or U12934 (N_12934,N_11191,N_11509);
or U12935 (N_12935,N_11696,N_11373);
or U12936 (N_12936,N_11681,N_11246);
and U12937 (N_12937,N_11020,N_11897);
or U12938 (N_12938,N_11513,N_11361);
xor U12939 (N_12939,N_11881,N_11673);
nand U12940 (N_12940,N_11469,N_11005);
and U12941 (N_12941,N_11480,N_11262);
and U12942 (N_12942,N_11032,N_11754);
xor U12943 (N_12943,N_11094,N_11542);
nor U12944 (N_12944,N_11341,N_11748);
nand U12945 (N_12945,N_11698,N_11602);
xor U12946 (N_12946,N_11445,N_11798);
or U12947 (N_12947,N_11384,N_11541);
and U12948 (N_12948,N_11594,N_11191);
nor U12949 (N_12949,N_11971,N_11041);
or U12950 (N_12950,N_11613,N_11032);
or U12951 (N_12951,N_11951,N_11187);
nor U12952 (N_12952,N_11579,N_11646);
or U12953 (N_12953,N_11207,N_11510);
or U12954 (N_12954,N_11625,N_11394);
xor U12955 (N_12955,N_11329,N_11381);
or U12956 (N_12956,N_11502,N_11595);
xnor U12957 (N_12957,N_11921,N_11887);
nand U12958 (N_12958,N_11483,N_11938);
or U12959 (N_12959,N_11292,N_11798);
or U12960 (N_12960,N_11460,N_11914);
xor U12961 (N_12961,N_11238,N_11631);
and U12962 (N_12962,N_11629,N_11365);
and U12963 (N_12963,N_11948,N_11307);
nor U12964 (N_12964,N_11579,N_11152);
or U12965 (N_12965,N_11144,N_11432);
nand U12966 (N_12966,N_11436,N_11791);
nand U12967 (N_12967,N_11542,N_11004);
nand U12968 (N_12968,N_11616,N_11471);
nand U12969 (N_12969,N_11179,N_11728);
nand U12970 (N_12970,N_11926,N_11552);
nor U12971 (N_12971,N_11470,N_11391);
or U12972 (N_12972,N_11279,N_11314);
nor U12973 (N_12973,N_11854,N_11327);
xor U12974 (N_12974,N_11557,N_11620);
and U12975 (N_12975,N_11557,N_11806);
nor U12976 (N_12976,N_11791,N_11163);
or U12977 (N_12977,N_11396,N_11082);
or U12978 (N_12978,N_11534,N_11656);
and U12979 (N_12979,N_11524,N_11442);
and U12980 (N_12980,N_11049,N_11656);
nor U12981 (N_12981,N_11734,N_11226);
xnor U12982 (N_12982,N_11742,N_11581);
nand U12983 (N_12983,N_11678,N_11298);
nand U12984 (N_12984,N_11990,N_11840);
xnor U12985 (N_12985,N_11559,N_11394);
or U12986 (N_12986,N_11822,N_11538);
nand U12987 (N_12987,N_11043,N_11471);
nand U12988 (N_12988,N_11451,N_11943);
nand U12989 (N_12989,N_11270,N_11351);
or U12990 (N_12990,N_11278,N_11243);
or U12991 (N_12991,N_11623,N_11406);
nor U12992 (N_12992,N_11011,N_11047);
and U12993 (N_12993,N_11933,N_11626);
xnor U12994 (N_12994,N_11340,N_11195);
and U12995 (N_12995,N_11239,N_11575);
nor U12996 (N_12996,N_11134,N_11960);
nand U12997 (N_12997,N_11792,N_11698);
or U12998 (N_12998,N_11269,N_11689);
nand U12999 (N_12999,N_11819,N_11021);
nor U13000 (N_13000,N_12719,N_12699);
and U13001 (N_13001,N_12825,N_12709);
or U13002 (N_13002,N_12624,N_12094);
nor U13003 (N_13003,N_12451,N_12492);
or U13004 (N_13004,N_12490,N_12707);
nor U13005 (N_13005,N_12248,N_12395);
nand U13006 (N_13006,N_12364,N_12590);
xnor U13007 (N_13007,N_12425,N_12276);
or U13008 (N_13008,N_12156,N_12204);
or U13009 (N_13009,N_12401,N_12378);
nor U13010 (N_13010,N_12754,N_12135);
nor U13011 (N_13011,N_12381,N_12999);
or U13012 (N_13012,N_12234,N_12374);
xnor U13013 (N_13013,N_12314,N_12457);
and U13014 (N_13014,N_12211,N_12169);
nand U13015 (N_13015,N_12918,N_12201);
or U13016 (N_13016,N_12546,N_12812);
and U13017 (N_13017,N_12220,N_12046);
xor U13018 (N_13018,N_12871,N_12938);
or U13019 (N_13019,N_12838,N_12856);
or U13020 (N_13020,N_12223,N_12003);
nand U13021 (N_13021,N_12500,N_12720);
and U13022 (N_13022,N_12133,N_12956);
xor U13023 (N_13023,N_12961,N_12322);
nand U13024 (N_13024,N_12847,N_12319);
and U13025 (N_13025,N_12281,N_12298);
xor U13026 (N_13026,N_12170,N_12723);
nor U13027 (N_13027,N_12888,N_12743);
nor U13028 (N_13028,N_12066,N_12829);
nor U13029 (N_13029,N_12379,N_12869);
and U13030 (N_13030,N_12540,N_12670);
or U13031 (N_13031,N_12102,N_12832);
nor U13032 (N_13032,N_12702,N_12266);
xor U13033 (N_13033,N_12041,N_12718);
xnor U13034 (N_13034,N_12311,N_12712);
nand U13035 (N_13035,N_12076,N_12556);
and U13036 (N_13036,N_12687,N_12142);
nand U13037 (N_13037,N_12932,N_12139);
and U13038 (N_13038,N_12384,N_12031);
or U13039 (N_13039,N_12431,N_12749);
or U13040 (N_13040,N_12108,N_12496);
nor U13041 (N_13041,N_12997,N_12423);
nor U13042 (N_13042,N_12522,N_12755);
or U13043 (N_13043,N_12441,N_12786);
nand U13044 (N_13044,N_12734,N_12567);
nor U13045 (N_13045,N_12766,N_12898);
and U13046 (N_13046,N_12148,N_12853);
nand U13047 (N_13047,N_12525,N_12370);
nand U13048 (N_13048,N_12554,N_12769);
and U13049 (N_13049,N_12030,N_12412);
nor U13050 (N_13050,N_12273,N_12666);
or U13051 (N_13051,N_12153,N_12328);
nand U13052 (N_13052,N_12009,N_12551);
or U13053 (N_13053,N_12122,N_12351);
or U13054 (N_13054,N_12713,N_12845);
nor U13055 (N_13055,N_12627,N_12430);
and U13056 (N_13056,N_12916,N_12239);
xnor U13057 (N_13057,N_12919,N_12501);
xor U13058 (N_13058,N_12930,N_12538);
and U13059 (N_13059,N_12461,N_12692);
and U13060 (N_13060,N_12489,N_12329);
nor U13061 (N_13061,N_12249,N_12576);
nor U13062 (N_13062,N_12990,N_12811);
nand U13063 (N_13063,N_12025,N_12776);
or U13064 (N_13064,N_12126,N_12427);
nor U13065 (N_13065,N_12198,N_12965);
and U13066 (N_13066,N_12032,N_12879);
or U13067 (N_13067,N_12323,N_12992);
nand U13068 (N_13068,N_12438,N_12778);
nor U13069 (N_13069,N_12969,N_12596);
xnor U13070 (N_13070,N_12691,N_12482);
nor U13071 (N_13071,N_12034,N_12343);
nand U13072 (N_13072,N_12040,N_12964);
or U13073 (N_13073,N_12012,N_12217);
nor U13074 (N_13074,N_12453,N_12528);
or U13075 (N_13075,N_12388,N_12664);
xnor U13076 (N_13076,N_12909,N_12305);
nor U13077 (N_13077,N_12111,N_12793);
xnor U13078 (N_13078,N_12268,N_12112);
nand U13079 (N_13079,N_12420,N_12468);
nand U13080 (N_13080,N_12353,N_12020);
nor U13081 (N_13081,N_12448,N_12405);
and U13082 (N_13082,N_12459,N_12739);
nand U13083 (N_13083,N_12195,N_12503);
nand U13084 (N_13084,N_12746,N_12458);
xor U13085 (N_13085,N_12147,N_12418);
and U13086 (N_13086,N_12790,N_12107);
nand U13087 (N_13087,N_12649,N_12098);
and U13088 (N_13088,N_12610,N_12494);
nand U13089 (N_13089,N_12611,N_12715);
nand U13090 (N_13090,N_12660,N_12868);
nor U13091 (N_13091,N_12658,N_12072);
or U13092 (N_13092,N_12117,N_12228);
nand U13093 (N_13093,N_12760,N_12493);
nand U13094 (N_13094,N_12599,N_12140);
nor U13095 (N_13095,N_12327,N_12800);
and U13096 (N_13096,N_12928,N_12529);
xnor U13097 (N_13097,N_12758,N_12864);
xor U13098 (N_13098,N_12113,N_12360);
nor U13099 (N_13099,N_12238,N_12345);
nand U13100 (N_13100,N_12836,N_12733);
nor U13101 (N_13101,N_12834,N_12306);
and U13102 (N_13102,N_12612,N_12792);
and U13103 (N_13103,N_12550,N_12245);
and U13104 (N_13104,N_12725,N_12741);
nand U13105 (N_13105,N_12049,N_12481);
or U13106 (N_13106,N_12545,N_12044);
nor U13107 (N_13107,N_12697,N_12943);
or U13108 (N_13108,N_12075,N_12752);
nor U13109 (N_13109,N_12149,N_12972);
or U13110 (N_13110,N_12318,N_12613);
nand U13111 (N_13111,N_12277,N_12059);
and U13112 (N_13112,N_12183,N_12189);
nor U13113 (N_13113,N_12410,N_12101);
nor U13114 (N_13114,N_12645,N_12141);
nor U13115 (N_13115,N_12167,N_12827);
nor U13116 (N_13116,N_12700,N_12794);
nand U13117 (N_13117,N_12465,N_12215);
xor U13118 (N_13118,N_12502,N_12002);
and U13119 (N_13119,N_12386,N_12770);
nand U13120 (N_13120,N_12678,N_12882);
and U13121 (N_13121,N_12051,N_12574);
or U13122 (N_13122,N_12548,N_12250);
xor U13123 (N_13123,N_12667,N_12475);
xor U13124 (N_13124,N_12162,N_12432);
nand U13125 (N_13125,N_12115,N_12783);
and U13126 (N_13126,N_12192,N_12352);
nand U13127 (N_13127,N_12143,N_12464);
nor U13128 (N_13128,N_12454,N_12690);
nor U13129 (N_13129,N_12945,N_12279);
nand U13130 (N_13130,N_12299,N_12340);
or U13131 (N_13131,N_12206,N_12802);
or U13132 (N_13132,N_12698,N_12000);
or U13133 (N_13133,N_12067,N_12337);
or U13134 (N_13134,N_12443,N_12643);
and U13135 (N_13135,N_12803,N_12638);
xor U13136 (N_13136,N_12841,N_12214);
xor U13137 (N_13137,N_12495,N_12607);
xnor U13138 (N_13138,N_12578,N_12870);
and U13139 (N_13139,N_12436,N_12620);
nand U13140 (N_13140,N_12657,N_12161);
and U13141 (N_13141,N_12924,N_12132);
or U13142 (N_13142,N_12282,N_12773);
and U13143 (N_13143,N_12477,N_12842);
xor U13144 (N_13144,N_12929,N_12602);
or U13145 (N_13145,N_12287,N_12199);
nand U13146 (N_13146,N_12512,N_12335);
nor U13147 (N_13147,N_12855,N_12526);
and U13148 (N_13148,N_12908,N_12336);
or U13149 (N_13149,N_12226,N_12190);
and U13150 (N_13150,N_12019,N_12534);
or U13151 (N_13151,N_12285,N_12603);
or U13152 (N_13152,N_12594,N_12124);
nand U13153 (N_13153,N_12208,N_12301);
nor U13154 (N_13154,N_12609,N_12200);
or U13155 (N_13155,N_12744,N_12768);
or U13156 (N_13156,N_12110,N_12974);
and U13157 (N_13157,N_12038,N_12524);
or U13158 (N_13158,N_12780,N_12865);
nand U13159 (N_13159,N_12785,N_12806);
or U13160 (N_13160,N_12325,N_12530);
xnor U13161 (N_13161,N_12092,N_12136);
or U13162 (N_13162,N_12194,N_12380);
xor U13163 (N_13163,N_12202,N_12315);
or U13164 (N_13164,N_12821,N_12073);
or U13165 (N_13165,N_12417,N_12696);
or U13166 (N_13166,N_12058,N_12523);
nor U13167 (N_13167,N_12042,N_12818);
xor U13168 (N_13168,N_12949,N_12767);
or U13169 (N_13169,N_12456,N_12617);
and U13170 (N_13170,N_12463,N_12580);
nand U13171 (N_13171,N_12317,N_12584);
and U13172 (N_13172,N_12497,N_12860);
and U13173 (N_13173,N_12573,N_12986);
or U13174 (N_13174,N_12669,N_12283);
nand U13175 (N_13175,N_12056,N_12396);
and U13176 (N_13176,N_12414,N_12679);
nor U13177 (N_13177,N_12555,N_12158);
or U13178 (N_13178,N_12680,N_12119);
xnor U13179 (N_13179,N_12730,N_12553);
nor U13180 (N_13180,N_12398,N_12907);
and U13181 (N_13181,N_12007,N_12387);
nor U13182 (N_13182,N_12586,N_12389);
nor U13183 (N_13183,N_12488,N_12369);
nor U13184 (N_13184,N_12628,N_12373);
nor U13185 (N_13185,N_12207,N_12349);
or U13186 (N_13186,N_12368,N_12906);
nand U13187 (N_13187,N_12506,N_12127);
xnor U13188 (N_13188,N_12491,N_12994);
and U13189 (N_13189,N_12963,N_12925);
or U13190 (N_13190,N_12828,N_12896);
or U13191 (N_13191,N_12371,N_12948);
or U13192 (N_13192,N_12814,N_12630);
nor U13193 (N_13193,N_12951,N_12191);
nand U13194 (N_13194,N_12471,N_12772);
and U13195 (N_13195,N_12247,N_12023);
nand U13196 (N_13196,N_12593,N_12840);
nor U13197 (N_13197,N_12426,N_12236);
nor U13198 (N_13198,N_12577,N_12676);
and U13199 (N_13199,N_12510,N_12015);
nand U13200 (N_13200,N_12960,N_12375);
xor U13201 (N_13201,N_12656,N_12174);
or U13202 (N_13202,N_12077,N_12957);
or U13203 (N_13203,N_12237,N_12606);
nor U13204 (N_13204,N_12258,N_12672);
and U13205 (N_13205,N_12784,N_12138);
and U13206 (N_13206,N_12449,N_12120);
and U13207 (N_13207,N_12260,N_12937);
and U13208 (N_13208,N_12027,N_12867);
nand U13209 (N_13209,N_12099,N_12762);
nand U13210 (N_13210,N_12232,N_12419);
nand U13211 (N_13211,N_12947,N_12716);
nand U13212 (N_13212,N_12674,N_12022);
nand U13213 (N_13213,N_12857,N_12295);
and U13214 (N_13214,N_12682,N_12382);
nor U13215 (N_13215,N_12976,N_12823);
nand U13216 (N_13216,N_12757,N_12332);
or U13217 (N_13217,N_12155,N_12533);
nor U13218 (N_13218,N_12984,N_12354);
nor U13219 (N_13219,N_12391,N_12695);
nand U13220 (N_13220,N_12362,N_12243);
and U13221 (N_13221,N_12474,N_12995);
or U13222 (N_13222,N_12587,N_12350);
and U13223 (N_13223,N_12642,N_12128);
and U13224 (N_13224,N_12004,N_12383);
or U13225 (N_13225,N_12307,N_12789);
or U13226 (N_13226,N_12891,N_12618);
nor U13227 (N_13227,N_12303,N_12899);
and U13228 (N_13228,N_12193,N_12404);
nor U13229 (N_13229,N_12447,N_12728);
nand U13230 (N_13230,N_12854,N_12996);
or U13231 (N_13231,N_12230,N_12511);
nor U13232 (N_13232,N_12269,N_12748);
xnor U13233 (N_13233,N_12045,N_12097);
and U13234 (N_13234,N_12621,N_12498);
and U13235 (N_13235,N_12588,N_12326);
or U13236 (N_13236,N_12321,N_12035);
and U13237 (N_13237,N_12881,N_12085);
and U13238 (N_13238,N_12087,N_12255);
or U13239 (N_13239,N_12235,N_12017);
and U13240 (N_13240,N_12704,N_12859);
or U13241 (N_13241,N_12377,N_12437);
nor U13242 (N_13242,N_12982,N_12581);
nor U13243 (N_13243,N_12356,N_12765);
nand U13244 (N_13244,N_12654,N_12082);
or U13245 (N_13245,N_12872,N_12262);
and U13246 (N_13246,N_12355,N_12668);
and U13247 (N_13247,N_12822,N_12625);
nor U13248 (N_13248,N_12145,N_12900);
nand U13249 (N_13249,N_12125,N_12415);
and U13250 (N_13250,N_12653,N_12413);
nand U13251 (N_13251,N_12320,N_12705);
nor U13252 (N_13252,N_12114,N_12913);
nand U13253 (N_13253,N_12886,N_12069);
or U13254 (N_13254,N_12851,N_12950);
nor U13255 (N_13255,N_12646,N_12884);
and U13256 (N_13256,N_12626,N_12689);
nand U13257 (N_13257,N_12892,N_12589);
and U13258 (N_13258,N_12717,N_12751);
nand U13259 (N_13259,N_12629,N_12168);
nand U13260 (N_13260,N_12923,N_12693);
and U13261 (N_13261,N_12499,N_12100);
nor U13262 (N_13262,N_12361,N_12104);
nand U13263 (N_13263,N_12544,N_12348);
or U13264 (N_13264,N_12134,N_12181);
nor U13265 (N_13265,N_12406,N_12172);
and U13266 (N_13266,N_12917,N_12016);
or U13267 (N_13267,N_12053,N_12542);
nand U13268 (N_13268,N_12256,N_12787);
nand U13269 (N_13269,N_12402,N_12846);
and U13270 (N_13270,N_12835,N_12446);
or U13271 (N_13271,N_12559,N_12060);
and U13272 (N_13272,N_12105,N_12991);
nand U13273 (N_13273,N_12026,N_12397);
nor U13274 (N_13274,N_12547,N_12472);
nor U13275 (N_13275,N_12946,N_12342);
nor U13276 (N_13276,N_12952,N_12777);
nand U13277 (N_13277,N_12731,N_12054);
and U13278 (N_13278,N_12090,N_12601);
or U13279 (N_13279,N_12635,N_12647);
or U13280 (N_13280,N_12088,N_12324);
nand U13281 (N_13281,N_12347,N_12637);
nand U13282 (N_13282,N_12165,N_12175);
and U13283 (N_13283,N_12557,N_12759);
nand U13284 (N_13284,N_12592,N_12850);
and U13285 (N_13285,N_12808,N_12675);
nand U13286 (N_13286,N_12953,N_12640);
and U13287 (N_13287,N_12971,N_12517);
or U13288 (N_13288,N_12313,N_12876);
and U13289 (N_13289,N_12484,N_12543);
nor U13290 (N_13290,N_12959,N_12595);
nor U13291 (N_13291,N_12745,N_12344);
xor U13292 (N_13292,N_12409,N_12569);
nor U13293 (N_13293,N_12052,N_12970);
xnor U13294 (N_13294,N_12644,N_12706);
or U13295 (N_13295,N_12316,N_12967);
or U13296 (N_13296,N_12291,N_12966);
nand U13297 (N_13297,N_12979,N_12166);
xnor U13298 (N_13298,N_12819,N_12962);
nand U13299 (N_13299,N_12341,N_12508);
and U13300 (N_13300,N_12244,N_12209);
nand U13301 (N_13301,N_12936,N_12467);
nand U13302 (N_13302,N_12180,N_12150);
nand U13303 (N_13303,N_12205,N_12008);
nor U13304 (N_13304,N_12251,N_12159);
nor U13305 (N_13305,N_12095,N_12686);
and U13306 (N_13306,N_12179,N_12460);
nand U13307 (N_13307,N_12583,N_12103);
and U13308 (N_13308,N_12338,N_12615);
or U13309 (N_13309,N_12895,N_12036);
and U13310 (N_13310,N_12981,N_12428);
or U13311 (N_13311,N_12761,N_12805);
or U13312 (N_13312,N_12253,N_12521);
nor U13313 (N_13313,N_12504,N_12057);
and U13314 (N_13314,N_12037,N_12271);
nand U13315 (N_13315,N_12470,N_12650);
nor U13316 (N_13316,N_12176,N_12993);
nand U13317 (N_13317,N_12080,N_12849);
nor U13318 (N_13318,N_12597,N_12655);
xor U13319 (N_13319,N_12632,N_12272);
nand U13320 (N_13320,N_12429,N_12782);
nand U13321 (N_13321,N_12302,N_12722);
nor U13322 (N_13322,N_12921,N_12639);
xor U13323 (N_13323,N_12861,N_12659);
or U13324 (N_13324,N_12346,N_12310);
xor U13325 (N_13325,N_12435,N_12188);
or U13326 (N_13326,N_12393,N_12222);
nand U13327 (N_13327,N_12652,N_12096);
nand U13328 (N_13328,N_12330,N_12939);
nand U13329 (N_13329,N_12889,N_12357);
or U13330 (N_13330,N_12083,N_12411);
nor U13331 (N_13331,N_12527,N_12309);
nand U13332 (N_13332,N_12688,N_12940);
nor U13333 (N_13333,N_12050,N_12422);
or U13334 (N_13334,N_12958,N_12157);
and U13335 (N_13335,N_12146,N_12263);
or U13336 (N_13336,N_12478,N_12797);
or U13337 (N_13337,N_12365,N_12312);
and U13338 (N_13338,N_12252,N_12186);
or U13339 (N_13339,N_12756,N_12182);
or U13340 (N_13340,N_12614,N_12163);
nor U13341 (N_13341,N_12651,N_12973);
xor U13342 (N_13342,N_12485,N_12575);
xnor U13343 (N_13343,N_12296,N_12359);
or U13344 (N_13344,N_12562,N_12018);
and U13345 (N_13345,N_12505,N_12863);
or U13346 (N_13346,N_12385,N_12753);
or U13347 (N_13347,N_12781,N_12536);
nand U13348 (N_13348,N_12837,N_12093);
nand U13349 (N_13349,N_12985,N_12893);
nand U13350 (N_13350,N_12552,N_12604);
nand U13351 (N_13351,N_12297,N_12742);
and U13352 (N_13352,N_12775,N_12619);
and U13353 (N_13353,N_12570,N_12513);
or U13354 (N_13354,N_12983,N_12440);
or U13355 (N_13355,N_12844,N_12874);
nand U13356 (N_13356,N_12641,N_12915);
nor U13357 (N_13357,N_12541,N_12469);
nand U13358 (N_13358,N_12537,N_12520);
nor U13359 (N_13359,N_12998,N_12633);
and U13360 (N_13360,N_12065,N_12729);
nand U13361 (N_13361,N_12815,N_12333);
nand U13362 (N_13362,N_12278,N_12518);
nor U13363 (N_13363,N_12394,N_12931);
or U13364 (N_13364,N_12434,N_12028);
nand U13365 (N_13365,N_12852,N_12259);
nor U13366 (N_13366,N_12339,N_12064);
or U13367 (N_13367,N_12600,N_12839);
nor U13368 (N_13368,N_12400,N_12416);
and U13369 (N_13369,N_12796,N_12363);
xnor U13370 (N_13370,N_12684,N_12462);
xnor U13371 (N_13371,N_12880,N_12079);
or U13372 (N_13372,N_12582,N_12331);
nand U13373 (N_13373,N_12816,N_12476);
nor U13374 (N_13374,N_12144,N_12203);
nor U13375 (N_13375,N_12479,N_12694);
and U13376 (N_13376,N_12568,N_12450);
nor U13377 (N_13377,N_12480,N_12300);
or U13378 (N_13378,N_12560,N_12171);
or U13379 (N_13379,N_12735,N_12151);
or U13380 (N_13380,N_12137,N_12063);
and U13381 (N_13381,N_12442,N_12514);
nand U13382 (N_13382,N_12809,N_12010);
or U13383 (N_13383,N_12662,N_12293);
nand U13384 (N_13384,N_12914,N_12902);
and U13385 (N_13385,N_12944,N_12225);
or U13386 (N_13386,N_12288,N_12224);
or U13387 (N_13387,N_12121,N_12231);
xor U13388 (N_13388,N_12831,N_12873);
or U13389 (N_13389,N_12933,N_12084);
nor U13390 (N_13390,N_12390,N_12774);
nand U13391 (N_13391,N_12216,N_12875);
nand U13392 (N_13392,N_12622,N_12671);
or U13393 (N_13393,N_12903,N_12631);
nor U13394 (N_13394,N_12274,N_12877);
or U13395 (N_13395,N_12636,N_12024);
nand U13396 (N_13396,N_12106,N_12565);
or U13397 (N_13397,N_12061,N_12118);
xnor U13398 (N_13398,N_12033,N_12519);
nand U13399 (N_13399,N_12487,N_12021);
nor U13400 (N_13400,N_12732,N_12791);
and U13401 (N_13401,N_12261,N_12358);
and U13402 (N_13402,N_12724,N_12011);
xor U13403 (N_13403,N_12532,N_12885);
and U13404 (N_13404,N_12623,N_12935);
or U13405 (N_13405,N_12771,N_12566);
xnor U13406 (N_13406,N_12424,N_12164);
or U13407 (N_13407,N_12509,N_12710);
nor U13408 (N_13408,N_12708,N_12196);
and U13409 (N_13409,N_12116,N_12920);
and U13410 (N_13410,N_12071,N_12862);
or U13411 (N_13411,N_12403,N_12813);
nand U13412 (N_13412,N_12934,N_12091);
and U13413 (N_13413,N_12241,N_12910);
nand U13414 (N_13414,N_12798,N_12286);
nand U13415 (N_13415,N_12598,N_12294);
nor U13416 (N_13416,N_12372,N_12507);
nor U13417 (N_13417,N_12154,N_12740);
and U13418 (N_13418,N_12047,N_12807);
or U13419 (N_13419,N_12820,N_12685);
nand U13420 (N_13420,N_12616,N_12013);
nor U13421 (N_13421,N_12824,N_12421);
nand U13422 (N_13422,N_12591,N_12376);
or U13423 (N_13423,N_12055,N_12086);
nand U13424 (N_13424,N_12264,N_12683);
nor U13425 (N_13425,N_12585,N_12152);
or U13426 (N_13426,N_12246,N_12289);
nand U13427 (N_13427,N_12954,N_12178);
nor U13428 (N_13428,N_12292,N_12779);
nor U13429 (N_13429,N_12788,N_12212);
nand U13430 (N_13430,N_12801,N_12197);
and U13431 (N_13431,N_12160,N_12737);
and U13432 (N_13432,N_12081,N_12905);
or U13433 (N_13433,N_12515,N_12539);
nor U13434 (N_13434,N_12455,N_12270);
nand U13435 (N_13435,N_12433,N_12187);
nor U13436 (N_13436,N_12564,N_12227);
or U13437 (N_13437,N_12014,N_12736);
and U13438 (N_13438,N_12810,N_12608);
xnor U13439 (N_13439,N_12763,N_12681);
and U13440 (N_13440,N_12275,N_12795);
or U13441 (N_13441,N_12109,N_12473);
nand U13442 (N_13442,N_12219,N_12392);
or U13443 (N_13443,N_12334,N_12848);
and U13444 (N_13444,N_12367,N_12701);
and U13445 (N_13445,N_12130,N_12901);
or U13446 (N_13446,N_12254,N_12665);
or U13447 (N_13447,N_12308,N_12673);
nor U13448 (N_13448,N_12131,N_12267);
or U13449 (N_13449,N_12843,N_12579);
or U13450 (N_13450,N_12452,N_12922);
or U13451 (N_13451,N_12516,N_12048);
and U13452 (N_13452,N_12764,N_12408);
and U13453 (N_13453,N_12185,N_12663);
and U13454 (N_13454,N_12941,N_12444);
and U13455 (N_13455,N_12927,N_12561);
and U13456 (N_13456,N_12445,N_12304);
or U13457 (N_13457,N_12486,N_12980);
nand U13458 (N_13458,N_12830,N_12866);
nand U13459 (N_13459,N_12290,N_12070);
nand U13460 (N_13460,N_12799,N_12721);
and U13461 (N_13461,N_12265,N_12883);
and U13462 (N_13462,N_12043,N_12988);
nor U13463 (N_13463,N_12284,N_12177);
and U13464 (N_13464,N_12738,N_12750);
or U13465 (N_13465,N_12005,N_12711);
or U13466 (N_13466,N_12242,N_12897);
and U13467 (N_13467,N_12677,N_12926);
nor U13468 (N_13468,N_12240,N_12605);
and U13469 (N_13469,N_12878,N_12218);
nand U13470 (N_13470,N_12280,N_12942);
or U13471 (N_13471,N_12233,N_12977);
and U13472 (N_13472,N_12634,N_12858);
xnor U13473 (N_13473,N_12890,N_12123);
nor U13474 (N_13474,N_12213,N_12229);
nand U13475 (N_13475,N_12257,N_12703);
nand U13476 (N_13476,N_12572,N_12989);
nor U13477 (N_13477,N_12466,N_12726);
or U13478 (N_13478,N_12978,N_12439);
or U13479 (N_13479,N_12089,N_12074);
and U13480 (N_13480,N_12184,N_12648);
or U13481 (N_13481,N_12549,N_12804);
nor U13482 (N_13482,N_12975,N_12535);
and U13483 (N_13483,N_12366,N_12571);
and U13484 (N_13484,N_12531,N_12006);
or U13485 (N_13485,N_12894,N_12407);
or U13486 (N_13486,N_12987,N_12904);
and U13487 (N_13487,N_12399,N_12563);
or U13488 (N_13488,N_12129,N_12887);
and U13489 (N_13489,N_12001,N_12062);
and U13490 (N_13490,N_12826,N_12817);
nor U13491 (N_13491,N_12955,N_12039);
nor U13492 (N_13492,N_12912,N_12029);
and U13493 (N_13493,N_12483,N_12078);
or U13494 (N_13494,N_12747,N_12968);
or U13495 (N_13495,N_12661,N_12833);
nor U13496 (N_13496,N_12221,N_12173);
and U13497 (N_13497,N_12727,N_12210);
nand U13498 (N_13498,N_12714,N_12068);
or U13499 (N_13499,N_12558,N_12911);
or U13500 (N_13500,N_12478,N_12132);
or U13501 (N_13501,N_12870,N_12233);
nand U13502 (N_13502,N_12533,N_12283);
and U13503 (N_13503,N_12162,N_12640);
xnor U13504 (N_13504,N_12300,N_12122);
nand U13505 (N_13505,N_12251,N_12333);
xor U13506 (N_13506,N_12420,N_12304);
nand U13507 (N_13507,N_12186,N_12714);
nor U13508 (N_13508,N_12711,N_12762);
xnor U13509 (N_13509,N_12486,N_12779);
or U13510 (N_13510,N_12549,N_12446);
or U13511 (N_13511,N_12621,N_12723);
nand U13512 (N_13512,N_12081,N_12254);
or U13513 (N_13513,N_12959,N_12862);
nor U13514 (N_13514,N_12140,N_12035);
nor U13515 (N_13515,N_12184,N_12172);
and U13516 (N_13516,N_12218,N_12389);
xor U13517 (N_13517,N_12823,N_12148);
or U13518 (N_13518,N_12178,N_12799);
or U13519 (N_13519,N_12895,N_12553);
nand U13520 (N_13520,N_12241,N_12778);
xor U13521 (N_13521,N_12178,N_12568);
nand U13522 (N_13522,N_12223,N_12418);
nor U13523 (N_13523,N_12839,N_12311);
xnor U13524 (N_13524,N_12198,N_12686);
nor U13525 (N_13525,N_12715,N_12630);
xor U13526 (N_13526,N_12533,N_12016);
nand U13527 (N_13527,N_12081,N_12208);
and U13528 (N_13528,N_12860,N_12768);
and U13529 (N_13529,N_12460,N_12191);
xnor U13530 (N_13530,N_12557,N_12146);
and U13531 (N_13531,N_12926,N_12688);
or U13532 (N_13532,N_12240,N_12720);
nand U13533 (N_13533,N_12386,N_12538);
nand U13534 (N_13534,N_12140,N_12668);
and U13535 (N_13535,N_12343,N_12018);
xor U13536 (N_13536,N_12569,N_12034);
and U13537 (N_13537,N_12926,N_12520);
nor U13538 (N_13538,N_12649,N_12055);
nand U13539 (N_13539,N_12665,N_12780);
or U13540 (N_13540,N_12916,N_12133);
or U13541 (N_13541,N_12299,N_12359);
nand U13542 (N_13542,N_12804,N_12207);
xor U13543 (N_13543,N_12279,N_12869);
and U13544 (N_13544,N_12648,N_12093);
nor U13545 (N_13545,N_12669,N_12572);
and U13546 (N_13546,N_12592,N_12989);
and U13547 (N_13547,N_12528,N_12679);
nor U13548 (N_13548,N_12002,N_12519);
nand U13549 (N_13549,N_12720,N_12605);
nor U13550 (N_13550,N_12646,N_12973);
and U13551 (N_13551,N_12876,N_12399);
nand U13552 (N_13552,N_12015,N_12854);
or U13553 (N_13553,N_12979,N_12864);
nand U13554 (N_13554,N_12627,N_12863);
and U13555 (N_13555,N_12496,N_12294);
nor U13556 (N_13556,N_12072,N_12232);
nand U13557 (N_13557,N_12322,N_12776);
nand U13558 (N_13558,N_12932,N_12963);
nor U13559 (N_13559,N_12135,N_12206);
nor U13560 (N_13560,N_12259,N_12694);
and U13561 (N_13561,N_12243,N_12915);
or U13562 (N_13562,N_12560,N_12221);
nor U13563 (N_13563,N_12999,N_12630);
and U13564 (N_13564,N_12486,N_12916);
xnor U13565 (N_13565,N_12152,N_12912);
nand U13566 (N_13566,N_12967,N_12345);
and U13567 (N_13567,N_12494,N_12611);
nor U13568 (N_13568,N_12398,N_12591);
and U13569 (N_13569,N_12795,N_12969);
nor U13570 (N_13570,N_12530,N_12038);
nor U13571 (N_13571,N_12377,N_12797);
nand U13572 (N_13572,N_12330,N_12794);
xnor U13573 (N_13573,N_12265,N_12434);
and U13574 (N_13574,N_12255,N_12670);
or U13575 (N_13575,N_12228,N_12149);
nand U13576 (N_13576,N_12930,N_12752);
nor U13577 (N_13577,N_12244,N_12658);
or U13578 (N_13578,N_12395,N_12446);
nand U13579 (N_13579,N_12097,N_12519);
and U13580 (N_13580,N_12618,N_12782);
nand U13581 (N_13581,N_12783,N_12010);
or U13582 (N_13582,N_12584,N_12665);
xor U13583 (N_13583,N_12032,N_12804);
and U13584 (N_13584,N_12414,N_12743);
nand U13585 (N_13585,N_12438,N_12257);
nor U13586 (N_13586,N_12941,N_12528);
nand U13587 (N_13587,N_12927,N_12968);
nand U13588 (N_13588,N_12178,N_12145);
nand U13589 (N_13589,N_12836,N_12415);
and U13590 (N_13590,N_12360,N_12791);
nor U13591 (N_13591,N_12694,N_12018);
or U13592 (N_13592,N_12864,N_12594);
or U13593 (N_13593,N_12717,N_12761);
nand U13594 (N_13594,N_12662,N_12986);
and U13595 (N_13595,N_12125,N_12614);
or U13596 (N_13596,N_12666,N_12835);
xnor U13597 (N_13597,N_12167,N_12058);
or U13598 (N_13598,N_12088,N_12191);
and U13599 (N_13599,N_12139,N_12256);
and U13600 (N_13600,N_12969,N_12112);
or U13601 (N_13601,N_12245,N_12593);
nand U13602 (N_13602,N_12606,N_12378);
xor U13603 (N_13603,N_12999,N_12247);
and U13604 (N_13604,N_12254,N_12100);
or U13605 (N_13605,N_12128,N_12951);
or U13606 (N_13606,N_12477,N_12434);
nor U13607 (N_13607,N_12201,N_12915);
nor U13608 (N_13608,N_12243,N_12530);
and U13609 (N_13609,N_12984,N_12326);
xor U13610 (N_13610,N_12896,N_12643);
nand U13611 (N_13611,N_12386,N_12422);
nand U13612 (N_13612,N_12500,N_12477);
or U13613 (N_13613,N_12913,N_12605);
nand U13614 (N_13614,N_12589,N_12703);
and U13615 (N_13615,N_12681,N_12894);
nand U13616 (N_13616,N_12428,N_12653);
nand U13617 (N_13617,N_12129,N_12002);
nand U13618 (N_13618,N_12886,N_12361);
or U13619 (N_13619,N_12695,N_12975);
and U13620 (N_13620,N_12435,N_12635);
and U13621 (N_13621,N_12530,N_12581);
nand U13622 (N_13622,N_12264,N_12593);
nor U13623 (N_13623,N_12856,N_12417);
and U13624 (N_13624,N_12124,N_12553);
nand U13625 (N_13625,N_12224,N_12025);
nand U13626 (N_13626,N_12995,N_12819);
or U13627 (N_13627,N_12336,N_12259);
nor U13628 (N_13628,N_12080,N_12013);
and U13629 (N_13629,N_12568,N_12322);
nor U13630 (N_13630,N_12721,N_12452);
nor U13631 (N_13631,N_12612,N_12836);
and U13632 (N_13632,N_12572,N_12428);
and U13633 (N_13633,N_12651,N_12347);
or U13634 (N_13634,N_12613,N_12572);
nor U13635 (N_13635,N_12533,N_12268);
xnor U13636 (N_13636,N_12633,N_12671);
or U13637 (N_13637,N_12594,N_12835);
nor U13638 (N_13638,N_12222,N_12374);
nor U13639 (N_13639,N_12715,N_12176);
or U13640 (N_13640,N_12100,N_12726);
nor U13641 (N_13641,N_12570,N_12047);
nor U13642 (N_13642,N_12714,N_12373);
and U13643 (N_13643,N_12121,N_12111);
nand U13644 (N_13644,N_12858,N_12820);
nor U13645 (N_13645,N_12644,N_12675);
and U13646 (N_13646,N_12988,N_12177);
nor U13647 (N_13647,N_12941,N_12311);
and U13648 (N_13648,N_12378,N_12071);
or U13649 (N_13649,N_12155,N_12292);
nor U13650 (N_13650,N_12047,N_12408);
or U13651 (N_13651,N_12944,N_12837);
nor U13652 (N_13652,N_12542,N_12775);
or U13653 (N_13653,N_12159,N_12717);
nor U13654 (N_13654,N_12895,N_12833);
and U13655 (N_13655,N_12143,N_12815);
or U13656 (N_13656,N_12731,N_12486);
and U13657 (N_13657,N_12907,N_12585);
nor U13658 (N_13658,N_12216,N_12468);
and U13659 (N_13659,N_12342,N_12870);
nor U13660 (N_13660,N_12852,N_12514);
and U13661 (N_13661,N_12571,N_12804);
xor U13662 (N_13662,N_12499,N_12563);
xor U13663 (N_13663,N_12063,N_12992);
and U13664 (N_13664,N_12443,N_12012);
and U13665 (N_13665,N_12807,N_12751);
nand U13666 (N_13666,N_12377,N_12663);
xnor U13667 (N_13667,N_12903,N_12568);
xnor U13668 (N_13668,N_12209,N_12991);
nand U13669 (N_13669,N_12332,N_12942);
and U13670 (N_13670,N_12011,N_12075);
nand U13671 (N_13671,N_12763,N_12700);
nor U13672 (N_13672,N_12091,N_12064);
and U13673 (N_13673,N_12493,N_12942);
or U13674 (N_13674,N_12697,N_12668);
and U13675 (N_13675,N_12805,N_12287);
xnor U13676 (N_13676,N_12950,N_12710);
nor U13677 (N_13677,N_12058,N_12154);
nand U13678 (N_13678,N_12524,N_12055);
and U13679 (N_13679,N_12816,N_12646);
nor U13680 (N_13680,N_12246,N_12134);
nor U13681 (N_13681,N_12852,N_12885);
xnor U13682 (N_13682,N_12311,N_12435);
nor U13683 (N_13683,N_12830,N_12928);
or U13684 (N_13684,N_12681,N_12347);
nor U13685 (N_13685,N_12033,N_12607);
or U13686 (N_13686,N_12123,N_12186);
xnor U13687 (N_13687,N_12251,N_12398);
or U13688 (N_13688,N_12857,N_12639);
nor U13689 (N_13689,N_12391,N_12609);
and U13690 (N_13690,N_12138,N_12630);
xnor U13691 (N_13691,N_12197,N_12608);
xnor U13692 (N_13692,N_12495,N_12246);
and U13693 (N_13693,N_12641,N_12638);
nor U13694 (N_13694,N_12077,N_12596);
or U13695 (N_13695,N_12379,N_12668);
nor U13696 (N_13696,N_12522,N_12405);
or U13697 (N_13697,N_12081,N_12601);
nand U13698 (N_13698,N_12305,N_12618);
and U13699 (N_13699,N_12412,N_12074);
nand U13700 (N_13700,N_12562,N_12952);
nand U13701 (N_13701,N_12796,N_12093);
or U13702 (N_13702,N_12623,N_12603);
nor U13703 (N_13703,N_12270,N_12876);
nor U13704 (N_13704,N_12636,N_12741);
and U13705 (N_13705,N_12168,N_12223);
xnor U13706 (N_13706,N_12707,N_12144);
and U13707 (N_13707,N_12232,N_12917);
or U13708 (N_13708,N_12416,N_12135);
or U13709 (N_13709,N_12846,N_12884);
nor U13710 (N_13710,N_12789,N_12157);
or U13711 (N_13711,N_12022,N_12948);
xnor U13712 (N_13712,N_12992,N_12037);
and U13713 (N_13713,N_12475,N_12736);
nor U13714 (N_13714,N_12136,N_12603);
and U13715 (N_13715,N_12406,N_12733);
and U13716 (N_13716,N_12852,N_12358);
nand U13717 (N_13717,N_12478,N_12592);
or U13718 (N_13718,N_12595,N_12346);
nor U13719 (N_13719,N_12489,N_12948);
or U13720 (N_13720,N_12000,N_12928);
nor U13721 (N_13721,N_12785,N_12521);
and U13722 (N_13722,N_12988,N_12375);
and U13723 (N_13723,N_12556,N_12079);
and U13724 (N_13724,N_12657,N_12297);
and U13725 (N_13725,N_12058,N_12357);
or U13726 (N_13726,N_12832,N_12764);
nor U13727 (N_13727,N_12846,N_12765);
or U13728 (N_13728,N_12948,N_12965);
nor U13729 (N_13729,N_12477,N_12852);
and U13730 (N_13730,N_12283,N_12518);
or U13731 (N_13731,N_12216,N_12923);
or U13732 (N_13732,N_12221,N_12079);
nand U13733 (N_13733,N_12570,N_12514);
nand U13734 (N_13734,N_12191,N_12677);
nor U13735 (N_13735,N_12839,N_12617);
nand U13736 (N_13736,N_12939,N_12985);
nand U13737 (N_13737,N_12720,N_12990);
nor U13738 (N_13738,N_12648,N_12394);
or U13739 (N_13739,N_12812,N_12506);
nand U13740 (N_13740,N_12403,N_12348);
and U13741 (N_13741,N_12206,N_12290);
or U13742 (N_13742,N_12125,N_12540);
nor U13743 (N_13743,N_12606,N_12187);
nor U13744 (N_13744,N_12175,N_12400);
nand U13745 (N_13745,N_12306,N_12101);
or U13746 (N_13746,N_12818,N_12799);
nand U13747 (N_13747,N_12066,N_12396);
or U13748 (N_13748,N_12097,N_12448);
nor U13749 (N_13749,N_12088,N_12960);
and U13750 (N_13750,N_12886,N_12512);
or U13751 (N_13751,N_12657,N_12192);
nor U13752 (N_13752,N_12391,N_12406);
and U13753 (N_13753,N_12457,N_12998);
nand U13754 (N_13754,N_12751,N_12486);
or U13755 (N_13755,N_12963,N_12066);
or U13756 (N_13756,N_12415,N_12431);
nand U13757 (N_13757,N_12505,N_12915);
nor U13758 (N_13758,N_12773,N_12273);
nor U13759 (N_13759,N_12740,N_12829);
xor U13760 (N_13760,N_12463,N_12988);
nor U13761 (N_13761,N_12334,N_12496);
nand U13762 (N_13762,N_12530,N_12576);
nand U13763 (N_13763,N_12432,N_12102);
nand U13764 (N_13764,N_12930,N_12371);
nor U13765 (N_13765,N_12713,N_12711);
nand U13766 (N_13766,N_12905,N_12706);
or U13767 (N_13767,N_12977,N_12580);
nand U13768 (N_13768,N_12376,N_12612);
or U13769 (N_13769,N_12620,N_12749);
nor U13770 (N_13770,N_12030,N_12876);
nand U13771 (N_13771,N_12370,N_12496);
nand U13772 (N_13772,N_12922,N_12271);
nor U13773 (N_13773,N_12609,N_12860);
or U13774 (N_13774,N_12112,N_12079);
nor U13775 (N_13775,N_12807,N_12711);
and U13776 (N_13776,N_12268,N_12147);
nor U13777 (N_13777,N_12323,N_12407);
or U13778 (N_13778,N_12685,N_12459);
nor U13779 (N_13779,N_12998,N_12916);
nand U13780 (N_13780,N_12374,N_12700);
nor U13781 (N_13781,N_12847,N_12982);
or U13782 (N_13782,N_12474,N_12510);
nand U13783 (N_13783,N_12634,N_12703);
and U13784 (N_13784,N_12569,N_12731);
and U13785 (N_13785,N_12623,N_12663);
xnor U13786 (N_13786,N_12963,N_12991);
nand U13787 (N_13787,N_12243,N_12553);
nand U13788 (N_13788,N_12867,N_12626);
nor U13789 (N_13789,N_12302,N_12019);
or U13790 (N_13790,N_12306,N_12635);
and U13791 (N_13791,N_12909,N_12759);
and U13792 (N_13792,N_12300,N_12965);
or U13793 (N_13793,N_12989,N_12497);
and U13794 (N_13794,N_12099,N_12787);
or U13795 (N_13795,N_12979,N_12543);
nand U13796 (N_13796,N_12723,N_12733);
nor U13797 (N_13797,N_12528,N_12513);
and U13798 (N_13798,N_12635,N_12341);
and U13799 (N_13799,N_12297,N_12030);
nor U13800 (N_13800,N_12763,N_12958);
or U13801 (N_13801,N_12880,N_12943);
and U13802 (N_13802,N_12818,N_12696);
and U13803 (N_13803,N_12136,N_12286);
nand U13804 (N_13804,N_12340,N_12042);
nand U13805 (N_13805,N_12297,N_12314);
nor U13806 (N_13806,N_12839,N_12419);
or U13807 (N_13807,N_12902,N_12429);
nand U13808 (N_13808,N_12864,N_12357);
or U13809 (N_13809,N_12567,N_12715);
and U13810 (N_13810,N_12155,N_12048);
and U13811 (N_13811,N_12113,N_12742);
and U13812 (N_13812,N_12616,N_12442);
nor U13813 (N_13813,N_12881,N_12782);
nor U13814 (N_13814,N_12167,N_12728);
xor U13815 (N_13815,N_12829,N_12617);
and U13816 (N_13816,N_12152,N_12741);
and U13817 (N_13817,N_12812,N_12985);
xor U13818 (N_13818,N_12895,N_12391);
or U13819 (N_13819,N_12459,N_12201);
nand U13820 (N_13820,N_12480,N_12456);
nand U13821 (N_13821,N_12439,N_12815);
xnor U13822 (N_13822,N_12060,N_12669);
nor U13823 (N_13823,N_12672,N_12234);
or U13824 (N_13824,N_12175,N_12620);
and U13825 (N_13825,N_12246,N_12424);
or U13826 (N_13826,N_12276,N_12297);
and U13827 (N_13827,N_12835,N_12699);
xnor U13828 (N_13828,N_12489,N_12740);
and U13829 (N_13829,N_12733,N_12475);
xnor U13830 (N_13830,N_12545,N_12775);
or U13831 (N_13831,N_12458,N_12119);
nor U13832 (N_13832,N_12072,N_12088);
nor U13833 (N_13833,N_12740,N_12973);
xnor U13834 (N_13834,N_12239,N_12029);
nand U13835 (N_13835,N_12421,N_12188);
nor U13836 (N_13836,N_12359,N_12723);
nor U13837 (N_13837,N_12009,N_12489);
nor U13838 (N_13838,N_12440,N_12956);
xor U13839 (N_13839,N_12205,N_12520);
or U13840 (N_13840,N_12917,N_12392);
nand U13841 (N_13841,N_12147,N_12009);
and U13842 (N_13842,N_12865,N_12856);
nor U13843 (N_13843,N_12576,N_12344);
or U13844 (N_13844,N_12231,N_12598);
xnor U13845 (N_13845,N_12994,N_12474);
xor U13846 (N_13846,N_12096,N_12317);
nor U13847 (N_13847,N_12083,N_12610);
and U13848 (N_13848,N_12883,N_12216);
nor U13849 (N_13849,N_12506,N_12492);
or U13850 (N_13850,N_12286,N_12568);
nand U13851 (N_13851,N_12926,N_12533);
nand U13852 (N_13852,N_12336,N_12380);
or U13853 (N_13853,N_12376,N_12285);
or U13854 (N_13854,N_12484,N_12927);
or U13855 (N_13855,N_12208,N_12586);
or U13856 (N_13856,N_12592,N_12731);
and U13857 (N_13857,N_12789,N_12912);
xor U13858 (N_13858,N_12190,N_12670);
nand U13859 (N_13859,N_12367,N_12436);
nor U13860 (N_13860,N_12634,N_12974);
nand U13861 (N_13861,N_12989,N_12255);
nor U13862 (N_13862,N_12892,N_12323);
nor U13863 (N_13863,N_12713,N_12605);
nand U13864 (N_13864,N_12138,N_12376);
nand U13865 (N_13865,N_12127,N_12297);
nand U13866 (N_13866,N_12921,N_12907);
nor U13867 (N_13867,N_12500,N_12412);
nor U13868 (N_13868,N_12972,N_12376);
nor U13869 (N_13869,N_12283,N_12393);
nand U13870 (N_13870,N_12303,N_12092);
or U13871 (N_13871,N_12827,N_12348);
nor U13872 (N_13872,N_12763,N_12136);
and U13873 (N_13873,N_12082,N_12451);
nor U13874 (N_13874,N_12243,N_12640);
and U13875 (N_13875,N_12453,N_12393);
and U13876 (N_13876,N_12931,N_12526);
nor U13877 (N_13877,N_12667,N_12857);
nand U13878 (N_13878,N_12767,N_12469);
nor U13879 (N_13879,N_12778,N_12247);
nor U13880 (N_13880,N_12079,N_12085);
nand U13881 (N_13881,N_12354,N_12446);
and U13882 (N_13882,N_12741,N_12201);
nand U13883 (N_13883,N_12500,N_12618);
nor U13884 (N_13884,N_12941,N_12654);
or U13885 (N_13885,N_12806,N_12240);
or U13886 (N_13886,N_12385,N_12617);
nor U13887 (N_13887,N_12951,N_12824);
nor U13888 (N_13888,N_12132,N_12507);
and U13889 (N_13889,N_12579,N_12091);
nand U13890 (N_13890,N_12917,N_12957);
nand U13891 (N_13891,N_12607,N_12662);
and U13892 (N_13892,N_12381,N_12281);
nand U13893 (N_13893,N_12368,N_12568);
or U13894 (N_13894,N_12327,N_12420);
or U13895 (N_13895,N_12579,N_12358);
nand U13896 (N_13896,N_12179,N_12094);
or U13897 (N_13897,N_12562,N_12281);
nand U13898 (N_13898,N_12039,N_12383);
or U13899 (N_13899,N_12130,N_12808);
nand U13900 (N_13900,N_12908,N_12371);
or U13901 (N_13901,N_12568,N_12271);
xor U13902 (N_13902,N_12862,N_12750);
and U13903 (N_13903,N_12147,N_12399);
or U13904 (N_13904,N_12934,N_12536);
xor U13905 (N_13905,N_12135,N_12837);
nor U13906 (N_13906,N_12190,N_12678);
or U13907 (N_13907,N_12840,N_12366);
or U13908 (N_13908,N_12271,N_12460);
nand U13909 (N_13909,N_12804,N_12807);
xnor U13910 (N_13910,N_12865,N_12763);
nand U13911 (N_13911,N_12358,N_12966);
nor U13912 (N_13912,N_12025,N_12101);
and U13913 (N_13913,N_12600,N_12667);
and U13914 (N_13914,N_12503,N_12402);
nand U13915 (N_13915,N_12909,N_12622);
and U13916 (N_13916,N_12765,N_12961);
xor U13917 (N_13917,N_12675,N_12798);
nor U13918 (N_13918,N_12632,N_12634);
nand U13919 (N_13919,N_12710,N_12204);
nor U13920 (N_13920,N_12927,N_12378);
and U13921 (N_13921,N_12336,N_12998);
and U13922 (N_13922,N_12619,N_12540);
or U13923 (N_13923,N_12396,N_12993);
or U13924 (N_13924,N_12058,N_12363);
nand U13925 (N_13925,N_12816,N_12223);
nand U13926 (N_13926,N_12458,N_12662);
nand U13927 (N_13927,N_12746,N_12261);
nand U13928 (N_13928,N_12933,N_12643);
and U13929 (N_13929,N_12140,N_12948);
or U13930 (N_13930,N_12256,N_12318);
xnor U13931 (N_13931,N_12725,N_12370);
and U13932 (N_13932,N_12272,N_12836);
nor U13933 (N_13933,N_12073,N_12734);
and U13934 (N_13934,N_12270,N_12563);
nand U13935 (N_13935,N_12562,N_12546);
or U13936 (N_13936,N_12585,N_12434);
nand U13937 (N_13937,N_12639,N_12868);
and U13938 (N_13938,N_12970,N_12631);
or U13939 (N_13939,N_12800,N_12530);
nor U13940 (N_13940,N_12980,N_12586);
and U13941 (N_13941,N_12514,N_12946);
or U13942 (N_13942,N_12050,N_12399);
or U13943 (N_13943,N_12273,N_12373);
nor U13944 (N_13944,N_12079,N_12168);
nor U13945 (N_13945,N_12873,N_12054);
nor U13946 (N_13946,N_12697,N_12412);
xor U13947 (N_13947,N_12979,N_12020);
and U13948 (N_13948,N_12987,N_12112);
nand U13949 (N_13949,N_12318,N_12166);
and U13950 (N_13950,N_12405,N_12268);
nand U13951 (N_13951,N_12720,N_12777);
and U13952 (N_13952,N_12605,N_12163);
nor U13953 (N_13953,N_12304,N_12206);
and U13954 (N_13954,N_12267,N_12118);
nand U13955 (N_13955,N_12915,N_12916);
and U13956 (N_13956,N_12210,N_12477);
and U13957 (N_13957,N_12818,N_12421);
and U13958 (N_13958,N_12031,N_12881);
or U13959 (N_13959,N_12045,N_12658);
or U13960 (N_13960,N_12553,N_12722);
nand U13961 (N_13961,N_12563,N_12908);
and U13962 (N_13962,N_12145,N_12477);
or U13963 (N_13963,N_12983,N_12623);
or U13964 (N_13964,N_12576,N_12731);
and U13965 (N_13965,N_12435,N_12935);
or U13966 (N_13966,N_12317,N_12840);
nor U13967 (N_13967,N_12015,N_12016);
and U13968 (N_13968,N_12254,N_12531);
nor U13969 (N_13969,N_12234,N_12604);
nor U13970 (N_13970,N_12476,N_12929);
and U13971 (N_13971,N_12730,N_12643);
nand U13972 (N_13972,N_12125,N_12479);
or U13973 (N_13973,N_12401,N_12840);
xnor U13974 (N_13974,N_12117,N_12472);
or U13975 (N_13975,N_12186,N_12934);
and U13976 (N_13976,N_12601,N_12333);
or U13977 (N_13977,N_12655,N_12333);
nor U13978 (N_13978,N_12425,N_12893);
nor U13979 (N_13979,N_12141,N_12638);
and U13980 (N_13980,N_12728,N_12583);
nor U13981 (N_13981,N_12153,N_12651);
nor U13982 (N_13982,N_12438,N_12898);
nor U13983 (N_13983,N_12238,N_12406);
and U13984 (N_13984,N_12805,N_12571);
nand U13985 (N_13985,N_12675,N_12322);
xnor U13986 (N_13986,N_12096,N_12770);
and U13987 (N_13987,N_12518,N_12338);
nor U13988 (N_13988,N_12580,N_12362);
or U13989 (N_13989,N_12674,N_12032);
and U13990 (N_13990,N_12443,N_12214);
nor U13991 (N_13991,N_12011,N_12302);
nand U13992 (N_13992,N_12856,N_12679);
xnor U13993 (N_13993,N_12719,N_12874);
nor U13994 (N_13994,N_12767,N_12380);
xnor U13995 (N_13995,N_12369,N_12948);
and U13996 (N_13996,N_12495,N_12119);
nor U13997 (N_13997,N_12266,N_12202);
and U13998 (N_13998,N_12852,N_12438);
nand U13999 (N_13999,N_12426,N_12461);
and U14000 (N_14000,N_13856,N_13932);
nor U14001 (N_14001,N_13652,N_13472);
or U14002 (N_14002,N_13200,N_13124);
xor U14003 (N_14003,N_13260,N_13496);
xor U14004 (N_14004,N_13017,N_13855);
nand U14005 (N_14005,N_13187,N_13356);
nand U14006 (N_14006,N_13543,N_13815);
nor U14007 (N_14007,N_13629,N_13372);
and U14008 (N_14008,N_13140,N_13046);
nand U14009 (N_14009,N_13387,N_13926);
or U14010 (N_14010,N_13686,N_13096);
or U14011 (N_14011,N_13203,N_13661);
nand U14012 (N_14012,N_13454,N_13117);
nand U14013 (N_14013,N_13938,N_13732);
nand U14014 (N_14014,N_13004,N_13347);
or U14015 (N_14015,N_13104,N_13675);
and U14016 (N_14016,N_13476,N_13982);
xnor U14017 (N_14017,N_13175,N_13388);
and U14018 (N_14018,N_13863,N_13739);
or U14019 (N_14019,N_13719,N_13824);
nor U14020 (N_14020,N_13792,N_13624);
or U14021 (N_14021,N_13530,N_13746);
nand U14022 (N_14022,N_13781,N_13394);
and U14023 (N_14023,N_13945,N_13861);
nand U14024 (N_14024,N_13744,N_13099);
or U14025 (N_14025,N_13042,N_13509);
nand U14026 (N_14026,N_13079,N_13326);
nor U14027 (N_14027,N_13868,N_13314);
nand U14028 (N_14028,N_13890,N_13223);
nor U14029 (N_14029,N_13374,N_13603);
nand U14030 (N_14030,N_13378,N_13122);
and U14031 (N_14031,N_13438,N_13473);
and U14032 (N_14032,N_13163,N_13487);
or U14033 (N_14033,N_13297,N_13333);
nand U14034 (N_14034,N_13450,N_13261);
and U14035 (N_14035,N_13909,N_13900);
and U14036 (N_14036,N_13044,N_13155);
nor U14037 (N_14037,N_13797,N_13832);
nor U14038 (N_14038,N_13523,N_13330);
or U14039 (N_14039,N_13666,N_13174);
nand U14040 (N_14040,N_13960,N_13622);
or U14041 (N_14041,N_13384,N_13107);
or U14042 (N_14042,N_13741,N_13870);
and U14043 (N_14043,N_13048,N_13788);
xnor U14044 (N_14044,N_13625,N_13687);
nor U14045 (N_14045,N_13541,N_13241);
or U14046 (N_14046,N_13296,N_13136);
or U14047 (N_14047,N_13951,N_13897);
or U14048 (N_14048,N_13243,N_13440);
nor U14049 (N_14049,N_13114,N_13840);
xnor U14050 (N_14050,N_13071,N_13611);
and U14051 (N_14051,N_13933,N_13923);
or U14052 (N_14052,N_13838,N_13153);
xnor U14053 (N_14053,N_13289,N_13710);
and U14054 (N_14054,N_13720,N_13025);
xor U14055 (N_14055,N_13045,N_13874);
nand U14056 (N_14056,N_13468,N_13285);
nand U14057 (N_14057,N_13430,N_13845);
and U14058 (N_14058,N_13217,N_13366);
nor U14059 (N_14059,N_13711,N_13808);
and U14060 (N_14060,N_13783,N_13574);
and U14061 (N_14061,N_13278,N_13251);
nand U14062 (N_14062,N_13070,N_13764);
nand U14063 (N_14063,N_13427,N_13787);
nor U14064 (N_14064,N_13369,N_13007);
or U14065 (N_14065,N_13912,N_13602);
nand U14066 (N_14066,N_13731,N_13442);
xor U14067 (N_14067,N_13247,N_13995);
nand U14068 (N_14068,N_13585,N_13049);
xor U14069 (N_14069,N_13090,N_13804);
or U14070 (N_14070,N_13579,N_13225);
nand U14071 (N_14071,N_13906,N_13368);
or U14072 (N_14072,N_13228,N_13059);
and U14073 (N_14073,N_13133,N_13963);
nor U14074 (N_14074,N_13435,N_13955);
and U14075 (N_14075,N_13293,N_13650);
and U14076 (N_14076,N_13425,N_13307);
xor U14077 (N_14077,N_13696,N_13418);
and U14078 (N_14078,N_13498,N_13620);
and U14079 (N_14079,N_13789,N_13795);
and U14080 (N_14080,N_13121,N_13379);
and U14081 (N_14081,N_13000,N_13616);
nor U14082 (N_14082,N_13967,N_13670);
nand U14083 (N_14083,N_13779,N_13373);
nand U14084 (N_14084,N_13749,N_13705);
xor U14085 (N_14085,N_13306,N_13299);
or U14086 (N_14086,N_13984,N_13939);
nor U14087 (N_14087,N_13769,N_13263);
nand U14088 (N_14088,N_13847,N_13821);
and U14089 (N_14089,N_13648,N_13695);
nor U14090 (N_14090,N_13910,N_13619);
or U14091 (N_14091,N_13922,N_13202);
nor U14092 (N_14092,N_13817,N_13962);
nor U14093 (N_14093,N_13001,N_13645);
or U14094 (N_14094,N_13294,N_13097);
nand U14095 (N_14095,N_13814,N_13974);
nand U14096 (N_14096,N_13752,N_13807);
nor U14097 (N_14097,N_13084,N_13050);
nand U14098 (N_14098,N_13103,N_13823);
xor U14099 (N_14099,N_13295,N_13937);
and U14100 (N_14100,N_13165,N_13707);
and U14101 (N_14101,N_13522,N_13786);
and U14102 (N_14102,N_13891,N_13632);
nor U14103 (N_14103,N_13259,N_13382);
nor U14104 (N_14104,N_13902,N_13304);
nand U14105 (N_14105,N_13849,N_13030);
xor U14106 (N_14106,N_13637,N_13997);
and U14107 (N_14107,N_13189,N_13865);
or U14108 (N_14108,N_13751,N_13375);
and U14109 (N_14109,N_13069,N_13886);
nand U14110 (N_14110,N_13231,N_13181);
nor U14111 (N_14111,N_13180,N_13053);
nor U14112 (N_14112,N_13676,N_13342);
nor U14113 (N_14113,N_13564,N_13419);
nor U14114 (N_14114,N_13846,N_13542);
nand U14115 (N_14115,N_13584,N_13459);
nor U14116 (N_14116,N_13460,N_13486);
or U14117 (N_14117,N_13074,N_13322);
nor U14118 (N_14118,N_13346,N_13527);
nor U14119 (N_14119,N_13753,N_13396);
and U14120 (N_14120,N_13991,N_13286);
nor U14121 (N_14121,N_13420,N_13086);
nor U14122 (N_14122,N_13575,N_13463);
or U14123 (N_14123,N_13975,N_13218);
nand U14124 (N_14124,N_13742,N_13614);
nand U14125 (N_14125,N_13596,N_13727);
and U14126 (N_14126,N_13514,N_13833);
or U14127 (N_14127,N_13690,N_13483);
xnor U14128 (N_14128,N_13842,N_13467);
nand U14129 (N_14129,N_13935,N_13524);
nor U14130 (N_14130,N_13207,N_13106);
or U14131 (N_14131,N_13757,N_13580);
or U14132 (N_14132,N_13577,N_13201);
or U14133 (N_14133,N_13839,N_13777);
nor U14134 (N_14134,N_13465,N_13078);
nand U14135 (N_14135,N_13561,N_13367);
and U14136 (N_14136,N_13221,N_13703);
nand U14137 (N_14137,N_13308,N_13392);
xnor U14138 (N_14138,N_13248,N_13101);
and U14139 (N_14139,N_13398,N_13641);
nor U14140 (N_14140,N_13623,N_13344);
nand U14141 (N_14141,N_13733,N_13421);
and U14142 (N_14142,N_13879,N_13488);
nor U14143 (N_14143,N_13351,N_13162);
and U14144 (N_14144,N_13966,N_13607);
or U14145 (N_14145,N_13037,N_13386);
xor U14146 (N_14146,N_13417,N_13680);
or U14147 (N_14147,N_13844,N_13581);
or U14148 (N_14148,N_13829,N_13875);
nand U14149 (N_14149,N_13736,N_13455);
and U14150 (N_14150,N_13681,N_13776);
and U14151 (N_14151,N_13659,N_13631);
nand U14152 (N_14152,N_13635,N_13083);
or U14153 (N_14153,N_13002,N_13745);
nor U14154 (N_14154,N_13993,N_13920);
and U14155 (N_14155,N_13547,N_13529);
and U14156 (N_14156,N_13323,N_13925);
nand U14157 (N_14157,N_13885,N_13210);
nor U14158 (N_14158,N_13663,N_13766);
or U14159 (N_14159,N_13737,N_13456);
nand U14160 (N_14160,N_13972,N_13985);
nand U14161 (N_14161,N_13860,N_13432);
or U14162 (N_14162,N_13208,N_13971);
and U14163 (N_14163,N_13904,N_13519);
or U14164 (N_14164,N_13157,N_13994);
xor U14165 (N_14165,N_13056,N_13837);
nor U14166 (N_14166,N_13682,N_13081);
nor U14167 (N_14167,N_13812,N_13428);
nand U14168 (N_14168,N_13697,N_13612);
nand U14169 (N_14169,N_13944,N_13989);
nor U14170 (N_14170,N_13469,N_13088);
nand U14171 (N_14171,N_13149,N_13583);
nor U14172 (N_14172,N_13371,N_13717);
or U14173 (N_14173,N_13538,N_13598);
and U14174 (N_14174,N_13565,N_13771);
or U14175 (N_14175,N_13234,N_13878);
nand U14176 (N_14176,N_13021,N_13843);
and U14177 (N_14177,N_13446,N_13907);
nor U14178 (N_14178,N_13331,N_13305);
and U14179 (N_14179,N_13708,N_13236);
nand U14180 (N_14180,N_13076,N_13087);
nor U14181 (N_14181,N_13453,N_13759);
or U14182 (N_14182,N_13313,N_13826);
nor U14183 (N_14183,N_13132,N_13434);
and U14184 (N_14184,N_13630,N_13871);
and U14185 (N_14185,N_13146,N_13118);
nor U14186 (N_14186,N_13254,N_13532);
nand U14187 (N_14187,N_13319,N_13010);
nand U14188 (N_14188,N_13747,N_13409);
nand U14189 (N_14189,N_13743,N_13287);
and U14190 (N_14190,N_13031,N_13665);
nand U14191 (N_14191,N_13038,N_13570);
nor U14192 (N_14192,N_13292,N_13258);
and U14193 (N_14193,N_13600,N_13277);
and U14194 (N_14194,N_13204,N_13437);
and U14195 (N_14195,N_13300,N_13721);
nor U14196 (N_14196,N_13672,N_13230);
nand U14197 (N_14197,N_13397,N_13640);
or U14198 (N_14198,N_13917,N_13485);
nand U14199 (N_14199,N_13599,N_13197);
or U14200 (N_14200,N_13558,N_13706);
and U14201 (N_14201,N_13836,N_13478);
or U14202 (N_14202,N_13164,N_13948);
xnor U14203 (N_14203,N_13726,N_13255);
nor U14204 (N_14204,N_13798,N_13018);
xnor U14205 (N_14205,N_13229,N_13507);
and U14206 (N_14206,N_13237,N_13232);
nand U14207 (N_14207,N_13338,N_13859);
and U14208 (N_14208,N_13592,N_13271);
and U14209 (N_14209,N_13537,N_13634);
nor U14210 (N_14210,N_13395,N_13883);
and U14211 (N_14211,N_13257,N_13756);
nand U14212 (N_14212,N_13872,N_13867);
nand U14213 (N_14213,N_13284,N_13345);
and U14214 (N_14214,N_13533,N_13740);
nor U14215 (N_14215,N_13327,N_13760);
nor U14216 (N_14216,N_13723,N_13679);
nor U14217 (N_14217,N_13172,N_13281);
nor U14218 (N_14218,N_13589,N_13361);
and U14219 (N_14219,N_13276,N_13416);
or U14220 (N_14220,N_13851,N_13990);
and U14221 (N_14221,N_13317,N_13449);
or U14222 (N_14222,N_13638,N_13128);
or U14223 (N_14223,N_13439,N_13947);
nand U14224 (N_14224,N_13220,N_13301);
and U14225 (N_14225,N_13458,N_13154);
and U14226 (N_14226,N_13969,N_13063);
nor U14227 (N_14227,N_13095,N_13350);
and U14228 (N_14228,N_13072,N_13012);
nand U14229 (N_14229,N_13098,N_13692);
or U14230 (N_14230,N_13588,N_13853);
nor U14231 (N_14231,N_13363,N_13340);
nor U14232 (N_14232,N_13275,N_13793);
nand U14233 (N_14233,N_13192,N_13075);
or U14234 (N_14234,N_13073,N_13942);
and U14235 (N_14235,N_13791,N_13365);
or U14236 (N_14236,N_13080,N_13239);
nand U14237 (N_14237,N_13864,N_13362);
nand U14238 (N_14238,N_13482,N_13481);
or U14239 (N_14239,N_13977,N_13318);
or U14240 (N_14240,N_13660,N_13125);
nor U14241 (N_14241,N_13116,N_13490);
and U14242 (N_14242,N_13573,N_13688);
and U14243 (N_14243,N_13884,N_13671);
nor U14244 (N_14244,N_13763,N_13452);
nor U14245 (N_14245,N_13544,N_13968);
xnor U14246 (N_14246,N_13805,N_13518);
or U14247 (N_14247,N_13889,N_13120);
and U14248 (N_14248,N_13782,N_13170);
or U14249 (N_14249,N_13735,N_13712);
nand U14250 (N_14250,N_13502,N_13320);
or U14251 (N_14251,N_13662,N_13269);
and U14252 (N_14252,N_13267,N_13402);
xnor U14253 (N_14253,N_13950,N_13615);
and U14254 (N_14254,N_13609,N_13664);
or U14255 (N_14255,N_13178,N_13283);
or U14256 (N_14256,N_13822,N_13131);
xor U14257 (N_14257,N_13961,N_13550);
xor U14258 (N_14258,N_13159,N_13415);
or U14259 (N_14259,N_13321,N_13773);
xnor U14260 (N_14260,N_13355,N_13214);
xnor U14261 (N_14261,N_13272,N_13656);
and U14262 (N_14262,N_13068,N_13359);
or U14263 (N_14263,N_13184,N_13385);
nor U14264 (N_14264,N_13470,N_13852);
and U14265 (N_14265,N_13667,N_13970);
nand U14266 (N_14266,N_13414,N_13953);
or U14267 (N_14267,N_13256,N_13601);
xor U14268 (N_14268,N_13905,N_13504);
nor U14269 (N_14269,N_13457,N_13495);
xnor U14270 (N_14270,N_13934,N_13552);
or U14271 (N_14271,N_13730,N_13651);
or U14272 (N_14272,N_13092,N_13213);
nor U14273 (N_14273,N_13894,N_13156);
nor U14274 (N_14274,N_13576,N_13176);
xnor U14275 (N_14275,N_13043,N_13193);
xnor U14276 (N_14276,N_13593,N_13058);
nand U14277 (N_14277,N_13123,N_13578);
nor U14278 (N_14278,N_13709,N_13041);
or U14279 (N_14279,N_13475,N_13102);
xor U14280 (N_14280,N_13246,N_13525);
nand U14281 (N_14281,N_13893,N_13591);
and U14282 (N_14282,N_13358,N_13339);
xor U14283 (N_14283,N_13381,N_13899);
and U14284 (N_14284,N_13262,N_13540);
nand U14285 (N_14285,N_13834,N_13110);
or U14286 (N_14286,N_13226,N_13536);
nor U14287 (N_14287,N_13151,N_13901);
xor U14288 (N_14288,N_13186,N_13981);
nor U14289 (N_14289,N_13160,N_13940);
nand U14290 (N_14290,N_13198,N_13288);
and U14291 (N_14291,N_13590,N_13082);
and U14292 (N_14292,N_13813,N_13195);
nor U14293 (N_14293,N_13605,N_13216);
nand U14294 (N_14294,N_13657,N_13921);
nand U14295 (N_14295,N_13093,N_13423);
nand U14296 (N_14296,N_13597,N_13979);
nand U14297 (N_14297,N_13772,N_13765);
nor U14298 (N_14298,N_13335,N_13572);
nand U14299 (N_14299,N_13857,N_13413);
and U14300 (N_14300,N_13206,N_13965);
and U14301 (N_14301,N_13280,N_13222);
nand U14302 (N_14302,N_13761,N_13827);
or U14303 (N_14303,N_13790,N_13461);
or U14304 (N_14304,N_13728,N_13380);
and U14305 (N_14305,N_13245,N_13556);
and U14306 (N_14306,N_13956,N_13065);
xnor U14307 (N_14307,N_13535,N_13903);
nor U14308 (N_14308,N_13199,N_13100);
xor U14309 (N_14309,N_13515,N_13555);
nor U14310 (N_14310,N_13545,N_13913);
or U14311 (N_14311,N_13560,N_13499);
xnor U14312 (N_14312,N_13768,N_13862);
nor U14313 (N_14313,N_13253,N_13235);
or U14314 (N_14314,N_13762,N_13887);
nor U14315 (N_14315,N_13528,N_13562);
and U14316 (N_14316,N_13242,N_13479);
nand U14317 (N_14317,N_13051,N_13168);
and U14318 (N_14318,N_13064,N_13024);
or U14319 (N_14319,N_13400,N_13268);
nor U14320 (N_14320,N_13626,N_13119);
nand U14321 (N_14321,N_13215,N_13848);
or U14322 (N_14322,N_13546,N_13767);
nor U14323 (N_14323,N_13150,N_13850);
or U14324 (N_14324,N_13316,N_13784);
nand U14325 (N_14325,N_13606,N_13006);
or U14326 (N_14326,N_13698,N_13582);
and U14327 (N_14327,N_13061,N_13608);
nor U14328 (N_14328,N_13244,N_13066);
and U14329 (N_14329,N_13931,N_13055);
nor U14330 (N_14330,N_13594,N_13028);
nand U14331 (N_14331,N_13526,N_13022);
and U14332 (N_14332,N_13818,N_13587);
and U14333 (N_14333,N_13034,N_13513);
or U14334 (N_14334,N_13445,N_13112);
nor U14335 (N_14335,N_13801,N_13399);
nor U14336 (N_14336,N_13551,N_13447);
or U14337 (N_14337,N_13135,N_13655);
nand U14338 (N_14338,N_13334,N_13724);
nor U14339 (N_14339,N_13312,N_13754);
nor U14340 (N_14340,N_13952,N_13182);
nor U14341 (N_14341,N_13127,N_13716);
or U14342 (N_14342,N_13166,N_13143);
and U14343 (N_14343,N_13673,N_13183);
xor U14344 (N_14344,N_13512,N_13877);
nor U14345 (N_14345,N_13298,N_13406);
nor U14346 (N_14346,N_13976,N_13169);
or U14347 (N_14347,N_13554,N_13866);
nor U14348 (N_14348,N_13403,N_13161);
or U14349 (N_14349,N_13130,N_13310);
nand U14350 (N_14350,N_13704,N_13531);
nand U14351 (N_14351,N_13354,N_13353);
and U14352 (N_14352,N_13806,N_13964);
nand U14353 (N_14353,N_13383,N_13196);
and U14354 (N_14354,N_13139,N_13410);
or U14355 (N_14355,N_13085,N_13503);
or U14356 (N_14356,N_13389,N_13040);
nand U14357 (N_14357,N_13451,N_13290);
nand U14358 (N_14358,N_13986,N_13111);
or U14359 (N_14359,N_13954,N_13998);
nor U14360 (N_14360,N_13811,N_13658);
or U14361 (N_14361,N_13302,N_13802);
nand U14362 (N_14362,N_13138,N_13915);
nand U14363 (N_14363,N_13566,N_13559);
or U14364 (N_14364,N_13816,N_13194);
and U14365 (N_14365,N_13108,N_13343);
xnor U14366 (N_14366,N_13835,N_13500);
nand U14367 (N_14367,N_13026,N_13489);
and U14368 (N_14368,N_13315,N_13983);
nor U14369 (N_14369,N_13534,N_13273);
and U14370 (N_14370,N_13595,N_13003);
nand U14371 (N_14371,N_13027,N_13854);
nand U14372 (N_14372,N_13809,N_13474);
or U14373 (N_14373,N_13685,N_13426);
and U14374 (N_14374,N_13888,N_13785);
and U14375 (N_14375,N_13729,N_13799);
or U14376 (N_14376,N_13360,N_13443);
nor U14377 (N_14377,N_13882,N_13142);
or U14378 (N_14378,N_13508,N_13959);
and U14379 (N_14379,N_13390,N_13491);
or U14380 (N_14380,N_13190,N_13014);
or U14381 (N_14381,N_13946,N_13873);
nor U14382 (N_14382,N_13336,N_13571);
nand U14383 (N_14383,N_13444,N_13794);
or U14384 (N_14384,N_13497,N_13405);
nand U14385 (N_14385,N_13668,N_13325);
nand U14386 (N_14386,N_13352,N_13349);
nor U14387 (N_14387,N_13249,N_13678);
nand U14388 (N_14388,N_13091,N_13039);
nand U14389 (N_14389,N_13089,N_13683);
xnor U14390 (N_14390,N_13618,N_13436);
nand U14391 (N_14391,N_13477,N_13370);
nor U14392 (N_14392,N_13462,N_13191);
or U14393 (N_14393,N_13265,N_13148);
nor U14394 (N_14394,N_13211,N_13738);
nand U14395 (N_14395,N_13924,N_13778);
and U14396 (N_14396,N_13376,N_13109);
xor U14397 (N_14397,N_13930,N_13617);
and U14398 (N_14398,N_13011,N_13015);
or U14399 (N_14399,N_13173,N_13433);
nor U14400 (N_14400,N_13553,N_13147);
and U14401 (N_14401,N_13501,N_13141);
nand U14402 (N_14402,N_13005,N_13105);
or U14403 (N_14403,N_13684,N_13377);
and U14404 (N_14404,N_13699,N_13016);
and U14405 (N_14405,N_13047,N_13702);
nand U14406 (N_14406,N_13548,N_13480);
and U14407 (N_14407,N_13693,N_13219);
or U14408 (N_14408,N_13209,N_13803);
nand U14409 (N_14409,N_13918,N_13060);
and U14410 (N_14410,N_13401,N_13224);
or U14411 (N_14411,N_13694,N_13691);
nand U14412 (N_14412,N_13639,N_13610);
and U14413 (N_14413,N_13780,N_13291);
nor U14414 (N_14414,N_13404,N_13493);
xnor U14415 (N_14415,N_13145,N_13567);
nand U14416 (N_14416,N_13033,N_13422);
and U14417 (N_14417,N_13324,N_13113);
nor U14418 (N_14418,N_13510,N_13563);
nor U14419 (N_14419,N_13569,N_13700);
and U14420 (N_14420,N_13185,N_13825);
and U14421 (N_14421,N_13407,N_13332);
and U14422 (N_14422,N_13054,N_13627);
and U14423 (N_14423,N_13252,N_13188);
nor U14424 (N_14424,N_13516,N_13035);
and U14425 (N_14425,N_13032,N_13052);
and U14426 (N_14426,N_13715,N_13233);
or U14427 (N_14427,N_13770,N_13282);
nand U14428 (N_14428,N_13568,N_13929);
or U14429 (N_14429,N_13869,N_13303);
nand U14430 (N_14430,N_13820,N_13205);
or U14431 (N_14431,N_13774,N_13412);
nand U14432 (N_14432,N_13895,N_13828);
or U14433 (N_14433,N_13750,N_13713);
nand U14434 (N_14434,N_13628,N_13521);
or U14435 (N_14435,N_13941,N_13429);
xnor U14436 (N_14436,N_13876,N_13755);
or U14437 (N_14437,N_13701,N_13549);
nand U14438 (N_14438,N_13800,N_13464);
or U14439 (N_14439,N_13448,N_13466);
xnor U14440 (N_14440,N_13391,N_13357);
nor U14441 (N_14441,N_13238,N_13621);
xor U14442 (N_14442,N_13943,N_13831);
nor U14443 (N_14443,N_13654,N_13919);
nand U14444 (N_14444,N_13936,N_13311);
nor U14445 (N_14445,N_13393,N_13494);
xnor U14446 (N_14446,N_13009,N_13689);
nor U14447 (N_14447,N_13604,N_13179);
nand U14448 (N_14448,N_13408,N_13908);
xnor U14449 (N_14449,N_13279,N_13987);
and U14450 (N_14450,N_13013,N_13674);
or U14451 (N_14451,N_13329,N_13722);
or U14452 (N_14452,N_13748,N_13988);
and U14453 (N_14453,N_13227,N_13819);
nand U14454 (N_14454,N_13240,N_13928);
nor U14455 (N_14455,N_13796,N_13471);
nand U14456 (N_14456,N_13646,N_13029);
nor U14457 (N_14457,N_13266,N_13914);
xnor U14458 (N_14458,N_13177,N_13484);
nor U14459 (N_14459,N_13441,N_13898);
xor U14460 (N_14460,N_13999,N_13036);
xnor U14461 (N_14461,N_13810,N_13911);
and U14462 (N_14462,N_13057,N_13328);
nand U14463 (N_14463,N_13337,N_13949);
nor U14464 (N_14464,N_13094,N_13649);
nand U14465 (N_14465,N_13309,N_13019);
and U14466 (N_14466,N_13647,N_13008);
nand U14467 (N_14467,N_13411,N_13511);
nor U14468 (N_14468,N_13669,N_13152);
nand U14469 (N_14469,N_13725,N_13062);
and U14470 (N_14470,N_13144,N_13364);
nor U14471 (N_14471,N_13158,N_13539);
or U14472 (N_14472,N_13505,N_13958);
and U14473 (N_14473,N_13858,N_13520);
xor U14474 (N_14474,N_13020,N_13250);
nor U14475 (N_14475,N_13927,N_13644);
nor U14476 (N_14476,N_13978,N_13137);
or U14477 (N_14477,N_13586,N_13067);
nand U14478 (N_14478,N_13775,N_13270);
or U14479 (N_14479,N_13126,N_13212);
xnor U14480 (N_14480,N_13424,N_13677);
nor U14481 (N_14481,N_13980,N_13115);
and U14482 (N_14482,N_13643,N_13129);
xor U14483 (N_14483,N_13880,N_13992);
and U14484 (N_14484,N_13896,N_13642);
nand U14485 (N_14485,N_13881,N_13341);
and U14486 (N_14486,N_13167,N_13633);
nand U14487 (N_14487,N_13506,N_13714);
nand U14488 (N_14488,N_13653,N_13492);
or U14489 (N_14489,N_13636,N_13718);
xnor U14490 (N_14490,N_13758,N_13348);
nand U14491 (N_14491,N_13892,N_13431);
nor U14492 (N_14492,N_13171,N_13134);
and U14493 (N_14493,N_13830,N_13957);
and U14494 (N_14494,N_13916,N_13517);
nor U14495 (N_14495,N_13274,N_13557);
and U14496 (N_14496,N_13264,N_13734);
nand U14497 (N_14497,N_13996,N_13613);
or U14498 (N_14498,N_13973,N_13841);
or U14499 (N_14499,N_13023,N_13077);
or U14500 (N_14500,N_13124,N_13479);
or U14501 (N_14501,N_13129,N_13389);
or U14502 (N_14502,N_13909,N_13863);
or U14503 (N_14503,N_13235,N_13206);
nor U14504 (N_14504,N_13278,N_13858);
nand U14505 (N_14505,N_13388,N_13246);
and U14506 (N_14506,N_13167,N_13746);
or U14507 (N_14507,N_13930,N_13376);
nor U14508 (N_14508,N_13970,N_13284);
and U14509 (N_14509,N_13483,N_13933);
xnor U14510 (N_14510,N_13090,N_13880);
and U14511 (N_14511,N_13295,N_13309);
nor U14512 (N_14512,N_13811,N_13874);
nand U14513 (N_14513,N_13481,N_13439);
nor U14514 (N_14514,N_13680,N_13453);
xor U14515 (N_14515,N_13903,N_13160);
nand U14516 (N_14516,N_13006,N_13187);
or U14517 (N_14517,N_13021,N_13101);
and U14518 (N_14518,N_13849,N_13025);
nand U14519 (N_14519,N_13871,N_13142);
nor U14520 (N_14520,N_13371,N_13671);
and U14521 (N_14521,N_13320,N_13520);
nor U14522 (N_14522,N_13281,N_13065);
and U14523 (N_14523,N_13701,N_13856);
xor U14524 (N_14524,N_13451,N_13406);
xnor U14525 (N_14525,N_13374,N_13281);
and U14526 (N_14526,N_13273,N_13987);
or U14527 (N_14527,N_13395,N_13934);
xor U14528 (N_14528,N_13722,N_13944);
nand U14529 (N_14529,N_13987,N_13956);
or U14530 (N_14530,N_13275,N_13412);
nor U14531 (N_14531,N_13041,N_13738);
or U14532 (N_14532,N_13674,N_13401);
nor U14533 (N_14533,N_13195,N_13659);
or U14534 (N_14534,N_13052,N_13792);
and U14535 (N_14535,N_13065,N_13035);
or U14536 (N_14536,N_13854,N_13409);
nor U14537 (N_14537,N_13055,N_13764);
and U14538 (N_14538,N_13893,N_13853);
nand U14539 (N_14539,N_13030,N_13260);
or U14540 (N_14540,N_13494,N_13240);
nor U14541 (N_14541,N_13247,N_13607);
xnor U14542 (N_14542,N_13030,N_13871);
or U14543 (N_14543,N_13009,N_13304);
nand U14544 (N_14544,N_13708,N_13578);
xnor U14545 (N_14545,N_13869,N_13488);
nand U14546 (N_14546,N_13645,N_13944);
nand U14547 (N_14547,N_13325,N_13885);
nor U14548 (N_14548,N_13175,N_13365);
xor U14549 (N_14549,N_13309,N_13072);
or U14550 (N_14550,N_13285,N_13862);
nor U14551 (N_14551,N_13802,N_13896);
and U14552 (N_14552,N_13939,N_13625);
xor U14553 (N_14553,N_13883,N_13155);
nand U14554 (N_14554,N_13778,N_13328);
or U14555 (N_14555,N_13033,N_13478);
nor U14556 (N_14556,N_13567,N_13168);
and U14557 (N_14557,N_13859,N_13531);
nand U14558 (N_14558,N_13157,N_13692);
nand U14559 (N_14559,N_13460,N_13320);
or U14560 (N_14560,N_13166,N_13465);
or U14561 (N_14561,N_13352,N_13511);
and U14562 (N_14562,N_13685,N_13909);
nand U14563 (N_14563,N_13017,N_13953);
and U14564 (N_14564,N_13058,N_13186);
xnor U14565 (N_14565,N_13798,N_13717);
nor U14566 (N_14566,N_13486,N_13957);
nand U14567 (N_14567,N_13104,N_13676);
and U14568 (N_14568,N_13766,N_13067);
nand U14569 (N_14569,N_13934,N_13220);
and U14570 (N_14570,N_13492,N_13812);
or U14571 (N_14571,N_13718,N_13472);
xor U14572 (N_14572,N_13222,N_13229);
nor U14573 (N_14573,N_13668,N_13476);
nor U14574 (N_14574,N_13093,N_13075);
or U14575 (N_14575,N_13850,N_13062);
and U14576 (N_14576,N_13460,N_13404);
nor U14577 (N_14577,N_13831,N_13535);
or U14578 (N_14578,N_13197,N_13688);
nor U14579 (N_14579,N_13540,N_13995);
nand U14580 (N_14580,N_13439,N_13891);
nor U14581 (N_14581,N_13718,N_13823);
and U14582 (N_14582,N_13403,N_13828);
nor U14583 (N_14583,N_13594,N_13781);
nand U14584 (N_14584,N_13764,N_13744);
or U14585 (N_14585,N_13615,N_13143);
and U14586 (N_14586,N_13392,N_13479);
or U14587 (N_14587,N_13905,N_13765);
xor U14588 (N_14588,N_13099,N_13920);
or U14589 (N_14589,N_13391,N_13938);
nor U14590 (N_14590,N_13252,N_13362);
nand U14591 (N_14591,N_13563,N_13864);
xor U14592 (N_14592,N_13557,N_13395);
nand U14593 (N_14593,N_13451,N_13506);
nor U14594 (N_14594,N_13951,N_13319);
nor U14595 (N_14595,N_13917,N_13278);
nand U14596 (N_14596,N_13023,N_13375);
xnor U14597 (N_14597,N_13739,N_13134);
nand U14598 (N_14598,N_13872,N_13182);
and U14599 (N_14599,N_13415,N_13180);
xnor U14600 (N_14600,N_13944,N_13409);
nor U14601 (N_14601,N_13316,N_13991);
and U14602 (N_14602,N_13669,N_13418);
nand U14603 (N_14603,N_13680,N_13438);
nand U14604 (N_14604,N_13511,N_13306);
nand U14605 (N_14605,N_13454,N_13699);
nand U14606 (N_14606,N_13813,N_13433);
or U14607 (N_14607,N_13398,N_13985);
nand U14608 (N_14608,N_13653,N_13488);
and U14609 (N_14609,N_13683,N_13674);
and U14610 (N_14610,N_13398,N_13120);
nor U14611 (N_14611,N_13216,N_13692);
and U14612 (N_14612,N_13530,N_13747);
or U14613 (N_14613,N_13925,N_13793);
or U14614 (N_14614,N_13943,N_13527);
or U14615 (N_14615,N_13815,N_13710);
or U14616 (N_14616,N_13779,N_13197);
or U14617 (N_14617,N_13137,N_13427);
nand U14618 (N_14618,N_13847,N_13335);
and U14619 (N_14619,N_13237,N_13823);
nor U14620 (N_14620,N_13098,N_13651);
nor U14621 (N_14621,N_13754,N_13007);
and U14622 (N_14622,N_13810,N_13715);
and U14623 (N_14623,N_13217,N_13640);
or U14624 (N_14624,N_13290,N_13363);
or U14625 (N_14625,N_13289,N_13785);
nand U14626 (N_14626,N_13273,N_13766);
nor U14627 (N_14627,N_13010,N_13560);
and U14628 (N_14628,N_13845,N_13816);
nor U14629 (N_14629,N_13587,N_13262);
or U14630 (N_14630,N_13674,N_13601);
xor U14631 (N_14631,N_13114,N_13597);
nand U14632 (N_14632,N_13942,N_13500);
or U14633 (N_14633,N_13042,N_13539);
nand U14634 (N_14634,N_13468,N_13896);
nor U14635 (N_14635,N_13408,N_13504);
nor U14636 (N_14636,N_13829,N_13747);
or U14637 (N_14637,N_13692,N_13977);
nor U14638 (N_14638,N_13225,N_13053);
nor U14639 (N_14639,N_13354,N_13778);
and U14640 (N_14640,N_13187,N_13488);
and U14641 (N_14641,N_13395,N_13702);
nor U14642 (N_14642,N_13624,N_13029);
and U14643 (N_14643,N_13030,N_13075);
nor U14644 (N_14644,N_13885,N_13894);
nor U14645 (N_14645,N_13228,N_13906);
nand U14646 (N_14646,N_13519,N_13304);
nand U14647 (N_14647,N_13633,N_13547);
xnor U14648 (N_14648,N_13338,N_13558);
xor U14649 (N_14649,N_13626,N_13873);
nand U14650 (N_14650,N_13278,N_13993);
and U14651 (N_14651,N_13694,N_13001);
nor U14652 (N_14652,N_13973,N_13446);
nand U14653 (N_14653,N_13651,N_13617);
xor U14654 (N_14654,N_13528,N_13863);
or U14655 (N_14655,N_13956,N_13153);
and U14656 (N_14656,N_13300,N_13769);
nand U14657 (N_14657,N_13231,N_13799);
nand U14658 (N_14658,N_13538,N_13272);
xnor U14659 (N_14659,N_13389,N_13727);
or U14660 (N_14660,N_13272,N_13733);
nor U14661 (N_14661,N_13127,N_13478);
or U14662 (N_14662,N_13766,N_13431);
and U14663 (N_14663,N_13887,N_13690);
and U14664 (N_14664,N_13800,N_13466);
nand U14665 (N_14665,N_13785,N_13093);
nand U14666 (N_14666,N_13374,N_13774);
nand U14667 (N_14667,N_13207,N_13448);
nand U14668 (N_14668,N_13812,N_13589);
and U14669 (N_14669,N_13421,N_13389);
nand U14670 (N_14670,N_13809,N_13180);
nor U14671 (N_14671,N_13812,N_13787);
or U14672 (N_14672,N_13640,N_13645);
nand U14673 (N_14673,N_13288,N_13582);
nand U14674 (N_14674,N_13662,N_13737);
and U14675 (N_14675,N_13762,N_13578);
and U14676 (N_14676,N_13547,N_13376);
nand U14677 (N_14677,N_13970,N_13884);
or U14678 (N_14678,N_13581,N_13221);
and U14679 (N_14679,N_13138,N_13648);
or U14680 (N_14680,N_13419,N_13443);
and U14681 (N_14681,N_13017,N_13155);
and U14682 (N_14682,N_13846,N_13459);
xor U14683 (N_14683,N_13548,N_13782);
nor U14684 (N_14684,N_13049,N_13365);
or U14685 (N_14685,N_13199,N_13334);
xnor U14686 (N_14686,N_13188,N_13987);
nor U14687 (N_14687,N_13729,N_13333);
and U14688 (N_14688,N_13987,N_13432);
nor U14689 (N_14689,N_13461,N_13614);
or U14690 (N_14690,N_13702,N_13555);
nor U14691 (N_14691,N_13704,N_13856);
nor U14692 (N_14692,N_13023,N_13646);
nor U14693 (N_14693,N_13661,N_13950);
or U14694 (N_14694,N_13708,N_13143);
xnor U14695 (N_14695,N_13588,N_13460);
xor U14696 (N_14696,N_13518,N_13049);
xnor U14697 (N_14697,N_13538,N_13482);
nand U14698 (N_14698,N_13134,N_13537);
or U14699 (N_14699,N_13930,N_13584);
nand U14700 (N_14700,N_13359,N_13942);
nor U14701 (N_14701,N_13598,N_13046);
and U14702 (N_14702,N_13027,N_13878);
or U14703 (N_14703,N_13667,N_13193);
nor U14704 (N_14704,N_13924,N_13161);
nand U14705 (N_14705,N_13071,N_13549);
nor U14706 (N_14706,N_13971,N_13407);
or U14707 (N_14707,N_13112,N_13942);
nand U14708 (N_14708,N_13565,N_13473);
and U14709 (N_14709,N_13610,N_13586);
nand U14710 (N_14710,N_13715,N_13246);
nand U14711 (N_14711,N_13264,N_13134);
and U14712 (N_14712,N_13119,N_13137);
nand U14713 (N_14713,N_13881,N_13159);
nand U14714 (N_14714,N_13058,N_13723);
nand U14715 (N_14715,N_13847,N_13113);
and U14716 (N_14716,N_13403,N_13841);
or U14717 (N_14717,N_13467,N_13311);
and U14718 (N_14718,N_13809,N_13105);
or U14719 (N_14719,N_13856,N_13613);
xor U14720 (N_14720,N_13920,N_13310);
nor U14721 (N_14721,N_13438,N_13655);
nor U14722 (N_14722,N_13492,N_13742);
nor U14723 (N_14723,N_13188,N_13094);
nand U14724 (N_14724,N_13450,N_13367);
or U14725 (N_14725,N_13976,N_13094);
and U14726 (N_14726,N_13563,N_13743);
xnor U14727 (N_14727,N_13905,N_13809);
xnor U14728 (N_14728,N_13620,N_13236);
and U14729 (N_14729,N_13654,N_13184);
nand U14730 (N_14730,N_13470,N_13266);
and U14731 (N_14731,N_13442,N_13739);
or U14732 (N_14732,N_13914,N_13410);
nor U14733 (N_14733,N_13394,N_13860);
or U14734 (N_14734,N_13139,N_13038);
nor U14735 (N_14735,N_13414,N_13652);
nor U14736 (N_14736,N_13492,N_13060);
and U14737 (N_14737,N_13702,N_13775);
nand U14738 (N_14738,N_13018,N_13066);
nor U14739 (N_14739,N_13510,N_13583);
or U14740 (N_14740,N_13953,N_13322);
and U14741 (N_14741,N_13122,N_13354);
or U14742 (N_14742,N_13754,N_13468);
nand U14743 (N_14743,N_13394,N_13536);
and U14744 (N_14744,N_13437,N_13100);
or U14745 (N_14745,N_13416,N_13842);
nor U14746 (N_14746,N_13601,N_13412);
nor U14747 (N_14747,N_13990,N_13945);
xor U14748 (N_14748,N_13799,N_13069);
or U14749 (N_14749,N_13458,N_13142);
nand U14750 (N_14750,N_13724,N_13821);
nor U14751 (N_14751,N_13717,N_13930);
nand U14752 (N_14752,N_13229,N_13477);
nand U14753 (N_14753,N_13975,N_13436);
nor U14754 (N_14754,N_13336,N_13325);
nand U14755 (N_14755,N_13545,N_13512);
or U14756 (N_14756,N_13802,N_13764);
nand U14757 (N_14757,N_13018,N_13295);
nor U14758 (N_14758,N_13940,N_13509);
or U14759 (N_14759,N_13410,N_13676);
or U14760 (N_14760,N_13172,N_13009);
and U14761 (N_14761,N_13489,N_13629);
or U14762 (N_14762,N_13375,N_13302);
or U14763 (N_14763,N_13312,N_13213);
and U14764 (N_14764,N_13193,N_13385);
and U14765 (N_14765,N_13922,N_13741);
nand U14766 (N_14766,N_13328,N_13952);
xor U14767 (N_14767,N_13873,N_13433);
and U14768 (N_14768,N_13855,N_13500);
nor U14769 (N_14769,N_13290,N_13586);
nor U14770 (N_14770,N_13948,N_13517);
nor U14771 (N_14771,N_13507,N_13030);
or U14772 (N_14772,N_13810,N_13296);
or U14773 (N_14773,N_13509,N_13022);
nand U14774 (N_14774,N_13208,N_13535);
or U14775 (N_14775,N_13477,N_13790);
nand U14776 (N_14776,N_13600,N_13183);
or U14777 (N_14777,N_13674,N_13476);
nand U14778 (N_14778,N_13978,N_13690);
xnor U14779 (N_14779,N_13320,N_13617);
nor U14780 (N_14780,N_13559,N_13622);
nor U14781 (N_14781,N_13045,N_13456);
or U14782 (N_14782,N_13022,N_13913);
and U14783 (N_14783,N_13508,N_13776);
nor U14784 (N_14784,N_13889,N_13210);
nand U14785 (N_14785,N_13984,N_13173);
nand U14786 (N_14786,N_13107,N_13301);
nand U14787 (N_14787,N_13875,N_13579);
xor U14788 (N_14788,N_13387,N_13490);
nor U14789 (N_14789,N_13290,N_13708);
nor U14790 (N_14790,N_13982,N_13472);
and U14791 (N_14791,N_13444,N_13851);
or U14792 (N_14792,N_13882,N_13643);
or U14793 (N_14793,N_13943,N_13654);
xnor U14794 (N_14794,N_13569,N_13164);
nor U14795 (N_14795,N_13864,N_13423);
nand U14796 (N_14796,N_13486,N_13242);
and U14797 (N_14797,N_13444,N_13947);
and U14798 (N_14798,N_13052,N_13865);
and U14799 (N_14799,N_13272,N_13971);
and U14800 (N_14800,N_13896,N_13204);
nand U14801 (N_14801,N_13063,N_13684);
or U14802 (N_14802,N_13730,N_13536);
nor U14803 (N_14803,N_13594,N_13158);
nor U14804 (N_14804,N_13754,N_13356);
and U14805 (N_14805,N_13924,N_13154);
or U14806 (N_14806,N_13411,N_13212);
nand U14807 (N_14807,N_13533,N_13771);
nor U14808 (N_14808,N_13762,N_13638);
and U14809 (N_14809,N_13592,N_13834);
nor U14810 (N_14810,N_13072,N_13916);
and U14811 (N_14811,N_13336,N_13885);
and U14812 (N_14812,N_13159,N_13131);
or U14813 (N_14813,N_13679,N_13217);
or U14814 (N_14814,N_13842,N_13562);
and U14815 (N_14815,N_13966,N_13990);
and U14816 (N_14816,N_13150,N_13340);
nand U14817 (N_14817,N_13626,N_13812);
nand U14818 (N_14818,N_13421,N_13099);
or U14819 (N_14819,N_13207,N_13125);
and U14820 (N_14820,N_13755,N_13495);
xor U14821 (N_14821,N_13121,N_13122);
and U14822 (N_14822,N_13668,N_13542);
nor U14823 (N_14823,N_13422,N_13957);
nand U14824 (N_14824,N_13582,N_13454);
nor U14825 (N_14825,N_13574,N_13492);
or U14826 (N_14826,N_13270,N_13646);
nor U14827 (N_14827,N_13305,N_13971);
or U14828 (N_14828,N_13106,N_13167);
nand U14829 (N_14829,N_13611,N_13168);
xor U14830 (N_14830,N_13904,N_13960);
or U14831 (N_14831,N_13752,N_13690);
xor U14832 (N_14832,N_13912,N_13802);
nand U14833 (N_14833,N_13984,N_13460);
and U14834 (N_14834,N_13508,N_13799);
nand U14835 (N_14835,N_13007,N_13752);
nand U14836 (N_14836,N_13741,N_13776);
nor U14837 (N_14837,N_13098,N_13003);
or U14838 (N_14838,N_13559,N_13061);
nor U14839 (N_14839,N_13559,N_13511);
nand U14840 (N_14840,N_13840,N_13227);
or U14841 (N_14841,N_13245,N_13005);
or U14842 (N_14842,N_13096,N_13867);
and U14843 (N_14843,N_13460,N_13061);
or U14844 (N_14844,N_13772,N_13864);
nor U14845 (N_14845,N_13855,N_13672);
or U14846 (N_14846,N_13685,N_13856);
nor U14847 (N_14847,N_13003,N_13562);
or U14848 (N_14848,N_13629,N_13502);
nor U14849 (N_14849,N_13913,N_13794);
nor U14850 (N_14850,N_13712,N_13993);
nand U14851 (N_14851,N_13836,N_13654);
nand U14852 (N_14852,N_13063,N_13925);
nor U14853 (N_14853,N_13400,N_13207);
or U14854 (N_14854,N_13649,N_13905);
or U14855 (N_14855,N_13274,N_13533);
nor U14856 (N_14856,N_13098,N_13761);
nor U14857 (N_14857,N_13875,N_13190);
xor U14858 (N_14858,N_13482,N_13673);
nand U14859 (N_14859,N_13052,N_13204);
nand U14860 (N_14860,N_13405,N_13874);
or U14861 (N_14861,N_13109,N_13365);
nand U14862 (N_14862,N_13283,N_13478);
nand U14863 (N_14863,N_13228,N_13400);
and U14864 (N_14864,N_13897,N_13065);
or U14865 (N_14865,N_13019,N_13337);
nor U14866 (N_14866,N_13896,N_13645);
xor U14867 (N_14867,N_13628,N_13686);
nand U14868 (N_14868,N_13753,N_13687);
and U14869 (N_14869,N_13308,N_13343);
nor U14870 (N_14870,N_13610,N_13449);
nand U14871 (N_14871,N_13534,N_13416);
or U14872 (N_14872,N_13760,N_13812);
or U14873 (N_14873,N_13148,N_13716);
and U14874 (N_14874,N_13869,N_13383);
nor U14875 (N_14875,N_13953,N_13505);
xnor U14876 (N_14876,N_13266,N_13541);
or U14877 (N_14877,N_13112,N_13962);
and U14878 (N_14878,N_13078,N_13476);
nor U14879 (N_14879,N_13115,N_13725);
nor U14880 (N_14880,N_13712,N_13677);
nor U14881 (N_14881,N_13655,N_13396);
xor U14882 (N_14882,N_13052,N_13505);
nor U14883 (N_14883,N_13521,N_13369);
nand U14884 (N_14884,N_13680,N_13341);
and U14885 (N_14885,N_13140,N_13044);
nand U14886 (N_14886,N_13909,N_13214);
and U14887 (N_14887,N_13841,N_13491);
xor U14888 (N_14888,N_13668,N_13108);
and U14889 (N_14889,N_13007,N_13657);
or U14890 (N_14890,N_13231,N_13668);
or U14891 (N_14891,N_13794,N_13118);
and U14892 (N_14892,N_13707,N_13225);
or U14893 (N_14893,N_13631,N_13308);
or U14894 (N_14894,N_13415,N_13703);
xor U14895 (N_14895,N_13798,N_13260);
xor U14896 (N_14896,N_13031,N_13635);
or U14897 (N_14897,N_13809,N_13781);
or U14898 (N_14898,N_13005,N_13101);
nor U14899 (N_14899,N_13630,N_13484);
xor U14900 (N_14900,N_13159,N_13351);
nor U14901 (N_14901,N_13788,N_13556);
or U14902 (N_14902,N_13958,N_13046);
nand U14903 (N_14903,N_13141,N_13942);
and U14904 (N_14904,N_13507,N_13736);
xnor U14905 (N_14905,N_13555,N_13179);
xnor U14906 (N_14906,N_13971,N_13400);
nand U14907 (N_14907,N_13860,N_13810);
nor U14908 (N_14908,N_13413,N_13146);
and U14909 (N_14909,N_13980,N_13173);
nand U14910 (N_14910,N_13055,N_13031);
nand U14911 (N_14911,N_13331,N_13026);
nand U14912 (N_14912,N_13788,N_13619);
nand U14913 (N_14913,N_13202,N_13366);
nor U14914 (N_14914,N_13137,N_13574);
and U14915 (N_14915,N_13658,N_13970);
or U14916 (N_14916,N_13141,N_13265);
xor U14917 (N_14917,N_13356,N_13974);
or U14918 (N_14918,N_13816,N_13775);
nand U14919 (N_14919,N_13076,N_13985);
nand U14920 (N_14920,N_13162,N_13310);
or U14921 (N_14921,N_13192,N_13057);
or U14922 (N_14922,N_13085,N_13635);
nor U14923 (N_14923,N_13191,N_13260);
nand U14924 (N_14924,N_13537,N_13794);
nor U14925 (N_14925,N_13964,N_13133);
and U14926 (N_14926,N_13100,N_13393);
nand U14927 (N_14927,N_13419,N_13848);
xor U14928 (N_14928,N_13384,N_13844);
nand U14929 (N_14929,N_13303,N_13404);
nand U14930 (N_14930,N_13582,N_13895);
nand U14931 (N_14931,N_13888,N_13580);
and U14932 (N_14932,N_13345,N_13710);
and U14933 (N_14933,N_13234,N_13801);
or U14934 (N_14934,N_13617,N_13778);
xnor U14935 (N_14935,N_13339,N_13562);
nand U14936 (N_14936,N_13481,N_13388);
nor U14937 (N_14937,N_13933,N_13278);
and U14938 (N_14938,N_13565,N_13945);
nor U14939 (N_14939,N_13711,N_13932);
and U14940 (N_14940,N_13176,N_13045);
nor U14941 (N_14941,N_13536,N_13307);
and U14942 (N_14942,N_13664,N_13100);
nand U14943 (N_14943,N_13017,N_13866);
nor U14944 (N_14944,N_13931,N_13319);
and U14945 (N_14945,N_13263,N_13958);
or U14946 (N_14946,N_13342,N_13071);
nor U14947 (N_14947,N_13646,N_13685);
and U14948 (N_14948,N_13656,N_13930);
nor U14949 (N_14949,N_13202,N_13489);
and U14950 (N_14950,N_13276,N_13261);
and U14951 (N_14951,N_13484,N_13361);
xor U14952 (N_14952,N_13995,N_13318);
xnor U14953 (N_14953,N_13245,N_13353);
and U14954 (N_14954,N_13906,N_13059);
nor U14955 (N_14955,N_13137,N_13722);
and U14956 (N_14956,N_13279,N_13573);
or U14957 (N_14957,N_13587,N_13249);
and U14958 (N_14958,N_13558,N_13531);
xnor U14959 (N_14959,N_13244,N_13333);
nor U14960 (N_14960,N_13889,N_13097);
or U14961 (N_14961,N_13376,N_13083);
nor U14962 (N_14962,N_13577,N_13502);
and U14963 (N_14963,N_13930,N_13989);
xnor U14964 (N_14964,N_13390,N_13627);
or U14965 (N_14965,N_13212,N_13884);
nor U14966 (N_14966,N_13624,N_13132);
nor U14967 (N_14967,N_13118,N_13595);
xor U14968 (N_14968,N_13514,N_13702);
xnor U14969 (N_14969,N_13693,N_13157);
nor U14970 (N_14970,N_13680,N_13088);
and U14971 (N_14971,N_13968,N_13597);
and U14972 (N_14972,N_13441,N_13310);
or U14973 (N_14973,N_13228,N_13558);
and U14974 (N_14974,N_13571,N_13487);
and U14975 (N_14975,N_13214,N_13613);
or U14976 (N_14976,N_13997,N_13857);
xor U14977 (N_14977,N_13734,N_13951);
nand U14978 (N_14978,N_13912,N_13779);
and U14979 (N_14979,N_13536,N_13762);
and U14980 (N_14980,N_13194,N_13449);
nand U14981 (N_14981,N_13945,N_13146);
and U14982 (N_14982,N_13836,N_13323);
xnor U14983 (N_14983,N_13268,N_13914);
nand U14984 (N_14984,N_13308,N_13990);
nor U14985 (N_14985,N_13767,N_13751);
nor U14986 (N_14986,N_13099,N_13227);
or U14987 (N_14987,N_13396,N_13386);
and U14988 (N_14988,N_13379,N_13232);
xor U14989 (N_14989,N_13019,N_13626);
nand U14990 (N_14990,N_13211,N_13929);
or U14991 (N_14991,N_13907,N_13785);
nor U14992 (N_14992,N_13153,N_13665);
or U14993 (N_14993,N_13821,N_13852);
nor U14994 (N_14994,N_13081,N_13693);
nor U14995 (N_14995,N_13943,N_13055);
and U14996 (N_14996,N_13904,N_13648);
or U14997 (N_14997,N_13898,N_13930);
and U14998 (N_14998,N_13404,N_13487);
or U14999 (N_14999,N_13190,N_13638);
and UO_0 (O_0,N_14584,N_14347);
nand UO_1 (O_1,N_14383,N_14412);
or UO_2 (O_2,N_14311,N_14614);
nor UO_3 (O_3,N_14610,N_14053);
or UO_4 (O_4,N_14446,N_14884);
nand UO_5 (O_5,N_14439,N_14451);
nor UO_6 (O_6,N_14397,N_14068);
or UO_7 (O_7,N_14281,N_14806);
and UO_8 (O_8,N_14323,N_14407);
or UO_9 (O_9,N_14164,N_14623);
nor UO_10 (O_10,N_14106,N_14284);
and UO_11 (O_11,N_14608,N_14982);
nand UO_12 (O_12,N_14585,N_14219);
and UO_13 (O_13,N_14770,N_14073);
and UO_14 (O_14,N_14315,N_14196);
nor UO_15 (O_15,N_14405,N_14440);
nor UO_16 (O_16,N_14750,N_14067);
xnor UO_17 (O_17,N_14709,N_14208);
or UO_18 (O_18,N_14015,N_14892);
and UO_19 (O_19,N_14080,N_14613);
and UO_20 (O_20,N_14824,N_14466);
and UO_21 (O_21,N_14988,N_14695);
xor UO_22 (O_22,N_14426,N_14151);
nand UO_23 (O_23,N_14571,N_14897);
nor UO_24 (O_24,N_14257,N_14913);
or UO_25 (O_25,N_14510,N_14183);
and UO_26 (O_26,N_14538,N_14772);
nand UO_27 (O_27,N_14237,N_14098);
xnor UO_28 (O_28,N_14829,N_14222);
nor UO_29 (O_29,N_14187,N_14743);
or UO_30 (O_30,N_14018,N_14138);
xnor UO_31 (O_31,N_14767,N_14574);
or UO_32 (O_32,N_14305,N_14153);
or UO_33 (O_33,N_14903,N_14842);
xnor UO_34 (O_34,N_14508,N_14643);
and UO_35 (O_35,N_14720,N_14065);
and UO_36 (O_36,N_14373,N_14417);
or UO_37 (O_37,N_14423,N_14539);
nor UO_38 (O_38,N_14428,N_14130);
and UO_39 (O_39,N_14007,N_14447);
or UO_40 (O_40,N_14485,N_14231);
nor UO_41 (O_41,N_14513,N_14194);
nor UO_42 (O_42,N_14966,N_14169);
nand UO_43 (O_43,N_14274,N_14042);
or UO_44 (O_44,N_14896,N_14483);
nor UO_45 (O_45,N_14785,N_14490);
or UO_46 (O_46,N_14283,N_14351);
nand UO_47 (O_47,N_14109,N_14902);
xnor UO_48 (O_48,N_14798,N_14552);
nor UO_49 (O_49,N_14983,N_14502);
nor UO_50 (O_50,N_14167,N_14678);
and UO_51 (O_51,N_14604,N_14264);
nor UO_52 (O_52,N_14813,N_14648);
or UO_53 (O_53,N_14577,N_14127);
nand UO_54 (O_54,N_14946,N_14774);
nand UO_55 (O_55,N_14409,N_14805);
and UO_56 (O_56,N_14267,N_14043);
xnor UO_57 (O_57,N_14905,N_14396);
nand UO_58 (O_58,N_14273,N_14780);
or UO_59 (O_59,N_14697,N_14551);
nand UO_60 (O_60,N_14557,N_14924);
or UO_61 (O_61,N_14779,N_14074);
nand UO_62 (O_62,N_14736,N_14880);
and UO_63 (O_63,N_14083,N_14209);
and UO_64 (O_64,N_14023,N_14265);
and UO_65 (O_65,N_14576,N_14233);
nand UO_66 (O_66,N_14521,N_14995);
nor UO_67 (O_67,N_14454,N_14091);
nor UO_68 (O_68,N_14480,N_14854);
nand UO_69 (O_69,N_14642,N_14227);
nor UO_70 (O_70,N_14699,N_14645);
xor UO_71 (O_71,N_14596,N_14803);
and UO_72 (O_72,N_14246,N_14484);
xor UO_73 (O_73,N_14181,N_14816);
nor UO_74 (O_74,N_14634,N_14932);
and UO_75 (O_75,N_14994,N_14625);
nand UO_76 (O_76,N_14639,N_14890);
nor UO_77 (O_77,N_14408,N_14541);
nand UO_78 (O_78,N_14741,N_14319);
or UO_79 (O_79,N_14630,N_14954);
and UO_80 (O_80,N_14386,N_14911);
xor UO_81 (O_81,N_14533,N_14711);
or UO_82 (O_82,N_14518,N_14449);
and UO_83 (O_83,N_14673,N_14692);
or UO_84 (O_84,N_14685,N_14163);
xor UO_85 (O_85,N_14026,N_14955);
or UO_86 (O_86,N_14325,N_14293);
or UO_87 (O_87,N_14118,N_14089);
and UO_88 (O_88,N_14148,N_14135);
nand UO_89 (O_89,N_14182,N_14839);
nor UO_90 (O_90,N_14650,N_14885);
and UO_91 (O_91,N_14251,N_14989);
xnor UO_92 (O_92,N_14477,N_14342);
or UO_93 (O_93,N_14964,N_14154);
nand UO_94 (O_94,N_14618,N_14441);
and UO_95 (O_95,N_14509,N_14870);
nor UO_96 (O_96,N_14456,N_14934);
or UO_97 (O_97,N_14561,N_14256);
nor UO_98 (O_98,N_14278,N_14769);
nand UO_99 (O_99,N_14638,N_14554);
and UO_100 (O_100,N_14708,N_14835);
xor UO_101 (O_101,N_14531,N_14981);
nor UO_102 (O_102,N_14272,N_14811);
nand UO_103 (O_103,N_14092,N_14318);
and UO_104 (O_104,N_14263,N_14560);
nand UO_105 (O_105,N_14782,N_14668);
or UO_106 (O_106,N_14810,N_14374);
or UO_107 (O_107,N_14430,N_14609);
nand UO_108 (O_108,N_14476,N_14195);
xor UO_109 (O_109,N_14308,N_14629);
nor UO_110 (O_110,N_14165,N_14081);
or UO_111 (O_111,N_14355,N_14482);
or UO_112 (O_112,N_14635,N_14243);
and UO_113 (O_113,N_14545,N_14591);
and UO_114 (O_114,N_14716,N_14918);
nor UO_115 (O_115,N_14357,N_14158);
nand UO_116 (O_116,N_14666,N_14301);
nand UO_117 (O_117,N_14529,N_14881);
or UO_118 (O_118,N_14783,N_14559);
xnor UO_119 (O_119,N_14809,N_14052);
nor UO_120 (O_120,N_14605,N_14398);
nand UO_121 (O_121,N_14090,N_14300);
and UO_122 (O_122,N_14242,N_14268);
nand UO_123 (O_123,N_14786,N_14376);
xor UO_124 (O_124,N_14058,N_14689);
or UO_125 (O_125,N_14710,N_14204);
xnor UO_126 (O_126,N_14760,N_14620);
nand UO_127 (O_127,N_14794,N_14136);
xnor UO_128 (O_128,N_14461,N_14329);
or UO_129 (O_129,N_14768,N_14724);
and UO_130 (O_130,N_14122,N_14380);
nor UO_131 (O_131,N_14929,N_14086);
or UO_132 (O_132,N_14140,N_14927);
xor UO_133 (O_133,N_14907,N_14356);
nand UO_134 (O_134,N_14358,N_14110);
nor UO_135 (O_135,N_14910,N_14202);
or UO_136 (O_136,N_14453,N_14761);
and UO_137 (O_137,N_14402,N_14201);
nor UO_138 (O_138,N_14354,N_14048);
xor UO_139 (O_139,N_14746,N_14258);
xor UO_140 (O_140,N_14393,N_14737);
and UO_141 (O_141,N_14463,N_14850);
nand UO_142 (O_142,N_14403,N_14221);
nor UO_143 (O_143,N_14525,N_14079);
and UO_144 (O_144,N_14500,N_14544);
and UO_145 (O_145,N_14705,N_14640);
nor UO_146 (O_146,N_14146,N_14965);
nand UO_147 (O_147,N_14787,N_14011);
xnor UO_148 (O_148,N_14844,N_14649);
and UO_149 (O_149,N_14797,N_14096);
or UO_150 (O_150,N_14861,N_14427);
nor UO_151 (O_151,N_14660,N_14587);
nand UO_152 (O_152,N_14132,N_14998);
nand UO_153 (O_153,N_14271,N_14900);
nand UO_154 (O_154,N_14877,N_14588);
and UO_155 (O_155,N_14951,N_14947);
or UO_156 (O_156,N_14626,N_14771);
nand UO_157 (O_157,N_14419,N_14343);
and UO_158 (O_158,N_14831,N_14808);
nand UO_159 (O_159,N_14247,N_14945);
nand UO_160 (O_160,N_14681,N_14107);
or UO_161 (O_161,N_14178,N_14622);
nor UO_162 (O_162,N_14933,N_14693);
nand UO_163 (O_163,N_14050,N_14475);
nor UO_164 (O_164,N_14312,N_14690);
xor UO_165 (O_165,N_14624,N_14987);
nor UO_166 (O_166,N_14899,N_14759);
nor UO_167 (O_167,N_14856,N_14168);
nor UO_168 (O_168,N_14742,N_14205);
nor UO_169 (O_169,N_14166,N_14150);
xor UO_170 (O_170,N_14159,N_14156);
nand UO_171 (O_171,N_14286,N_14336);
nor UO_172 (O_172,N_14418,N_14059);
and UO_173 (O_173,N_14647,N_14180);
and UO_174 (O_174,N_14249,N_14395);
xor UO_175 (O_175,N_14002,N_14119);
or UO_176 (O_176,N_14321,N_14819);
nand UO_177 (O_177,N_14784,N_14843);
xnor UO_178 (O_178,N_14491,N_14940);
nand UO_179 (O_179,N_14788,N_14662);
or UO_180 (O_180,N_14719,N_14290);
nor UO_181 (O_181,N_14879,N_14443);
nor UO_182 (O_182,N_14269,N_14641);
xor UO_183 (O_183,N_14517,N_14006);
and UO_184 (O_184,N_14145,N_14467);
or UO_185 (O_185,N_14543,N_14377);
or UO_186 (O_186,N_14516,N_14339);
and UO_187 (O_187,N_14962,N_14344);
nand UO_188 (O_188,N_14225,N_14341);
nor UO_189 (O_189,N_14241,N_14005);
nand UO_190 (O_190,N_14667,N_14324);
nor UO_191 (O_191,N_14128,N_14676);
and UO_192 (O_192,N_14238,N_14175);
xor UO_193 (O_193,N_14367,N_14149);
and UO_194 (O_194,N_14390,N_14572);
nor UO_195 (O_195,N_14188,N_14586);
and UO_196 (O_196,N_14970,N_14712);
nor UO_197 (O_197,N_14921,N_14817);
or UO_198 (O_198,N_14828,N_14665);
nand UO_199 (O_199,N_14536,N_14555);
nor UO_200 (O_200,N_14908,N_14976);
and UO_201 (O_201,N_14827,N_14352);
nand UO_202 (O_202,N_14567,N_14051);
nor UO_203 (O_203,N_14022,N_14914);
or UO_204 (O_204,N_14563,N_14392);
and UO_205 (O_205,N_14313,N_14171);
nand UO_206 (O_206,N_14060,N_14867);
xnor UO_207 (O_207,N_14046,N_14777);
and UO_208 (O_208,N_14024,N_14949);
nor UO_209 (O_209,N_14621,N_14706);
nor UO_210 (O_210,N_14112,N_14534);
or UO_211 (O_211,N_14391,N_14744);
nor UO_212 (O_212,N_14790,N_14943);
and UO_213 (O_213,N_14287,N_14549);
and UO_214 (O_214,N_14459,N_14592);
or UO_215 (O_215,N_14299,N_14972);
nand UO_216 (O_216,N_14414,N_14384);
or UO_217 (O_217,N_14142,N_14826);
or UO_218 (O_218,N_14923,N_14580);
or UO_219 (O_219,N_14566,N_14270);
or UO_220 (O_220,N_14298,N_14564);
or UO_221 (O_221,N_14192,N_14117);
xor UO_222 (O_222,N_14766,N_14996);
and UO_223 (O_223,N_14422,N_14226);
and UO_224 (O_224,N_14199,N_14114);
and UO_225 (O_225,N_14100,N_14959);
xor UO_226 (O_226,N_14916,N_14245);
nand UO_227 (O_227,N_14830,N_14364);
nand UO_228 (O_228,N_14922,N_14594);
nor UO_229 (O_229,N_14872,N_14825);
or UO_230 (O_230,N_14472,N_14986);
nand UO_231 (O_231,N_14595,N_14203);
and UO_232 (O_232,N_14152,N_14528);
nand UO_233 (O_233,N_14064,N_14277);
nor UO_234 (O_234,N_14631,N_14573);
or UO_235 (O_235,N_14993,N_14413);
and UO_236 (O_236,N_14677,N_14675);
nand UO_237 (O_237,N_14953,N_14057);
nand UO_238 (O_238,N_14530,N_14223);
and UO_239 (O_239,N_14473,N_14958);
or UO_240 (O_240,N_14433,N_14520);
xnor UO_241 (O_241,N_14756,N_14017);
or UO_242 (O_242,N_14411,N_14597);
or UO_243 (O_243,N_14088,N_14714);
and UO_244 (O_244,N_14436,N_14310);
nand UO_245 (O_245,N_14542,N_14230);
nor UO_246 (O_246,N_14029,N_14778);
nor UO_247 (O_247,N_14939,N_14044);
and UO_248 (O_248,N_14715,N_14800);
nor UO_249 (O_249,N_14296,N_14963);
nand UO_250 (O_250,N_14049,N_14859);
nor UO_251 (O_251,N_14537,N_14031);
and UO_252 (O_252,N_14570,N_14361);
or UO_253 (O_253,N_14801,N_14590);
or UO_254 (O_254,N_14886,N_14721);
nor UO_255 (O_255,N_14493,N_14812);
or UO_256 (O_256,N_14734,N_14087);
xnor UO_257 (O_257,N_14499,N_14193);
xor UO_258 (O_258,N_14304,N_14713);
or UO_259 (O_259,N_14314,N_14926);
or UO_260 (O_260,N_14838,N_14108);
or UO_261 (O_261,N_14878,N_14346);
or UO_262 (O_262,N_14874,N_14008);
nand UO_263 (O_263,N_14496,N_14462);
nor UO_264 (O_264,N_14589,N_14823);
nand UO_265 (O_265,N_14920,N_14655);
and UO_266 (O_266,N_14198,N_14335);
nand UO_267 (O_267,N_14445,N_14061);
nor UO_268 (O_268,N_14047,N_14847);
nor UO_269 (O_269,N_14206,N_14731);
and UO_270 (O_270,N_14745,N_14186);
nor UO_271 (O_271,N_14470,N_14925);
or UO_272 (O_272,N_14099,N_14285);
and UO_273 (O_273,N_14519,N_14228);
nor UO_274 (O_274,N_14240,N_14568);
nand UO_275 (O_275,N_14703,N_14253);
and UO_276 (O_276,N_14309,N_14973);
nor UO_277 (O_277,N_14001,N_14292);
nand UO_278 (O_278,N_14252,N_14365);
or UO_279 (O_279,N_14094,N_14653);
xnor UO_280 (O_280,N_14210,N_14035);
or UO_281 (O_281,N_14532,N_14468);
and UO_282 (O_282,N_14303,N_14575);
xnor UO_283 (O_283,N_14799,N_14214);
and UO_284 (O_284,N_14276,N_14616);
or UO_285 (O_285,N_14763,N_14294);
and UO_286 (O_286,N_14818,N_14753);
nand UO_287 (O_287,N_14935,N_14372);
nand UO_288 (O_288,N_14232,N_14184);
and UO_289 (O_289,N_14984,N_14974);
or UO_290 (O_290,N_14762,N_14124);
nor UO_291 (O_291,N_14707,N_14471);
or UO_292 (O_292,N_14280,N_14891);
nand UO_293 (O_293,N_14637,N_14038);
and UO_294 (O_294,N_14291,N_14322);
nor UO_295 (O_295,N_14833,N_14045);
or UO_296 (O_296,N_14056,N_14478);
or UO_297 (O_297,N_14895,N_14434);
nor UO_298 (O_298,N_14489,N_14220);
xor UO_299 (O_299,N_14978,N_14378);
nor UO_300 (O_300,N_14917,N_14550);
nand UO_301 (O_301,N_14021,N_14388);
nand UO_302 (O_302,N_14535,N_14952);
xnor UO_303 (O_303,N_14404,N_14350);
nor UO_304 (O_304,N_14144,N_14524);
or UO_305 (O_305,N_14956,N_14170);
xnor UO_306 (O_306,N_14834,N_14070);
and UO_307 (O_307,N_14619,N_14841);
and UO_308 (O_308,N_14328,N_14327);
or UO_309 (O_309,N_14999,N_14765);
nor UO_310 (O_310,N_14362,N_14793);
and UO_311 (O_311,N_14961,N_14944);
xnor UO_312 (O_312,N_14873,N_14345);
nand UO_313 (O_313,N_14928,N_14075);
nor UO_314 (O_314,N_14652,N_14837);
nand UO_315 (O_315,N_14093,N_14041);
nand UO_316 (O_316,N_14494,N_14368);
nand UO_317 (O_317,N_14275,N_14382);
or UO_318 (O_318,N_14656,N_14359);
or UO_319 (O_319,N_14431,N_14582);
and UO_320 (O_320,N_14254,N_14424);
and UO_321 (O_321,N_14694,N_14033);
and UO_322 (O_322,N_14452,N_14612);
nor UO_323 (O_323,N_14600,N_14248);
nor UO_324 (O_324,N_14120,N_14229);
nand UO_325 (O_325,N_14729,N_14333);
or UO_326 (O_326,N_14034,N_14234);
or UO_327 (O_327,N_14858,N_14740);
and UO_328 (O_328,N_14084,N_14749);
nand UO_329 (O_329,N_14791,N_14680);
and UO_330 (O_330,N_14822,N_14894);
or UO_331 (O_331,N_14394,N_14775);
nor UO_332 (O_332,N_14379,N_14448);
nor UO_333 (O_333,N_14215,N_14569);
or UO_334 (O_334,N_14071,N_14212);
nand UO_335 (O_335,N_14211,N_14565);
or UO_336 (O_336,N_14218,N_14004);
or UO_337 (O_337,N_14429,N_14032);
nand UO_338 (O_338,N_14028,N_14599);
nand UO_339 (O_339,N_14628,N_14919);
nor UO_340 (O_340,N_14698,N_14848);
and UO_341 (O_341,N_14863,N_14217);
or UO_342 (O_342,N_14754,N_14191);
or UO_343 (O_343,N_14686,N_14971);
nand UO_344 (O_344,N_14190,N_14522);
nor UO_345 (O_345,N_14134,N_14887);
nand UO_346 (O_346,N_14330,N_14792);
nand UO_347 (O_347,N_14882,N_14009);
and UO_348 (O_348,N_14039,N_14331);
nor UO_349 (O_349,N_14349,N_14735);
nand UO_350 (O_350,N_14723,N_14207);
nand UO_351 (O_351,N_14465,N_14845);
and UO_352 (O_352,N_14898,N_14072);
or UO_353 (O_353,N_14381,N_14279);
nand UO_354 (O_354,N_14661,N_14670);
or UO_355 (O_355,N_14871,N_14326);
or UO_356 (O_356,N_14450,N_14738);
or UO_357 (O_357,N_14438,N_14948);
nand UO_358 (O_358,N_14980,N_14025);
nor UO_359 (O_359,N_14224,N_14511);
and UO_360 (O_360,N_14406,N_14865);
nor UO_361 (O_361,N_14730,N_14486);
and UO_362 (O_362,N_14101,N_14912);
nor UO_363 (O_363,N_14627,N_14755);
or UO_364 (O_364,N_14869,N_14337);
or UO_365 (O_365,N_14646,N_14506);
or UO_366 (O_366,N_14722,N_14479);
nor UO_367 (O_367,N_14307,N_14636);
or UO_368 (O_368,N_14157,N_14930);
or UO_369 (O_369,N_14846,N_14733);
or UO_370 (O_370,N_14968,N_14679);
nand UO_371 (O_371,N_14155,N_14702);
and UO_372 (O_372,N_14505,N_14316);
or UO_373 (O_373,N_14030,N_14888);
nand UO_374 (O_374,N_14000,N_14657);
nor UO_375 (O_375,N_14547,N_14937);
or UO_376 (O_376,N_14503,N_14261);
xor UO_377 (O_377,N_14860,N_14901);
or UO_378 (O_378,N_14062,N_14410);
or UO_379 (O_379,N_14815,N_14764);
nor UO_380 (O_380,N_14868,N_14104);
or UO_381 (O_381,N_14370,N_14663);
nor UO_382 (O_382,N_14115,N_14758);
nand UO_383 (O_383,N_14526,N_14751);
and UO_384 (O_384,N_14684,N_14598);
and UO_385 (O_385,N_14085,N_14701);
or UO_386 (O_386,N_14338,N_14421);
nand UO_387 (O_387,N_14495,N_14967);
nor UO_388 (O_388,N_14054,N_14137);
or UO_389 (O_389,N_14603,N_14010);
and UO_390 (O_390,N_14683,N_14360);
nand UO_391 (O_391,N_14082,N_14727);
nand UO_392 (O_392,N_14583,N_14348);
or UO_393 (O_393,N_14804,N_14162);
or UO_394 (O_394,N_14027,N_14259);
or UO_395 (O_395,N_14936,N_14950);
nand UO_396 (O_396,N_14696,N_14832);
and UO_397 (O_397,N_14985,N_14415);
nor UO_398 (O_398,N_14632,N_14317);
or UO_399 (O_399,N_14197,N_14669);
nor UO_400 (O_400,N_14579,N_14401);
and UO_401 (O_401,N_14295,N_14400);
nor UO_402 (O_402,N_14385,N_14747);
xnor UO_403 (O_403,N_14332,N_14113);
xnor UO_404 (O_404,N_14302,N_14606);
nand UO_405 (O_405,N_14553,N_14003);
nor UO_406 (O_406,N_14013,N_14836);
xnor UO_407 (O_407,N_14236,N_14160);
and UO_408 (O_408,N_14416,N_14802);
nor UO_409 (O_409,N_14909,N_14375);
nor UO_410 (O_410,N_14726,N_14991);
and UO_411 (O_411,N_14282,N_14725);
or UO_412 (O_412,N_14617,N_14960);
nand UO_413 (O_413,N_14063,N_14717);
or UO_414 (O_414,N_14444,N_14975);
xor UO_415 (O_415,N_14931,N_14658);
nand UO_416 (O_416,N_14250,N_14123);
nand UO_417 (O_417,N_14432,N_14781);
nand UO_418 (O_418,N_14562,N_14387);
or UO_419 (O_419,N_14177,N_14789);
or UO_420 (O_420,N_14425,N_14523);
or UO_421 (O_421,N_14014,N_14688);
nand UO_422 (O_422,N_14992,N_14938);
and UO_423 (O_423,N_14040,N_14172);
or UO_424 (O_424,N_14548,N_14507);
or UO_425 (O_425,N_14851,N_14997);
nand UO_426 (O_426,N_14682,N_14102);
nand UO_427 (O_427,N_14469,N_14097);
nor UO_428 (O_428,N_14820,N_14875);
nor UO_429 (O_429,N_14514,N_14906);
nor UO_430 (O_430,N_14216,N_14176);
and UO_431 (O_431,N_14889,N_14353);
and UO_432 (O_432,N_14179,N_14457);
nor UO_433 (O_433,N_14795,N_14977);
or UO_434 (O_434,N_14289,N_14578);
nand UO_435 (O_435,N_14849,N_14139);
nand UO_436 (O_436,N_14644,N_14672);
nor UO_437 (O_437,N_14488,N_14855);
and UO_438 (O_438,N_14334,N_14244);
and UO_439 (O_439,N_14185,N_14674);
nand UO_440 (O_440,N_14147,N_14213);
xnor UO_441 (O_441,N_14807,N_14340);
xnor UO_442 (O_442,N_14288,N_14664);
xnor UO_443 (O_443,N_14055,N_14037);
nand UO_444 (O_444,N_14442,N_14990);
nor UO_445 (O_445,N_14602,N_14718);
xor UO_446 (O_446,N_14915,N_14077);
nand UO_447 (O_447,N_14369,N_14659);
or UO_448 (O_448,N_14601,N_14633);
nor UO_449 (O_449,N_14235,N_14857);
or UO_450 (O_450,N_14941,N_14487);
xnor UO_451 (O_451,N_14095,N_14474);
xnor UO_452 (O_452,N_14757,N_14739);
or UO_453 (O_453,N_14020,N_14687);
or UO_454 (O_454,N_14752,N_14512);
nor UO_455 (O_455,N_14066,N_14129);
nand UO_456 (O_456,N_14969,N_14076);
nand UO_457 (O_457,N_14455,N_14691);
and UO_458 (O_458,N_14069,N_14558);
nand UO_459 (O_459,N_14864,N_14671);
or UO_460 (O_460,N_14501,N_14111);
and UO_461 (O_461,N_14942,N_14796);
nor UO_462 (O_462,N_14019,N_14141);
or UO_463 (O_463,N_14420,N_14200);
nand UO_464 (O_464,N_14016,N_14540);
xor UO_465 (O_465,N_14497,N_14126);
nand UO_466 (O_466,N_14320,N_14876);
or UO_467 (O_467,N_14189,N_14078);
xnor UO_468 (O_468,N_14773,N_14399);
or UO_469 (O_469,N_14776,N_14121);
and UO_470 (O_470,N_14435,N_14748);
or UO_471 (O_471,N_14498,N_14389);
xor UO_472 (O_472,N_14704,N_14458);
nand UO_473 (O_473,N_14125,N_14814);
or UO_474 (O_474,N_14161,N_14979);
nand UO_475 (O_475,N_14904,N_14012);
xor UO_476 (O_476,N_14437,N_14239);
nand UO_477 (O_477,N_14460,N_14297);
and UO_478 (O_478,N_14957,N_14492);
nor UO_479 (O_479,N_14266,N_14174);
nor UO_480 (O_480,N_14654,N_14105);
or UO_481 (O_481,N_14700,N_14862);
nand UO_482 (O_482,N_14527,N_14116);
or UO_483 (O_483,N_14262,N_14371);
or UO_484 (O_484,N_14556,N_14853);
or UO_485 (O_485,N_14866,N_14103);
xnor UO_486 (O_486,N_14363,N_14515);
and UO_487 (O_487,N_14366,N_14143);
nand UO_488 (O_488,N_14883,N_14651);
nor UO_489 (O_489,N_14893,N_14611);
nand UO_490 (O_490,N_14504,N_14728);
nor UO_491 (O_491,N_14732,N_14581);
nand UO_492 (O_492,N_14852,N_14255);
nand UO_493 (O_493,N_14464,N_14306);
and UO_494 (O_494,N_14173,N_14133);
xor UO_495 (O_495,N_14821,N_14481);
or UO_496 (O_496,N_14607,N_14593);
nor UO_497 (O_497,N_14036,N_14546);
and UO_498 (O_498,N_14615,N_14840);
nand UO_499 (O_499,N_14260,N_14131);
nor UO_500 (O_500,N_14956,N_14596);
or UO_501 (O_501,N_14057,N_14296);
nor UO_502 (O_502,N_14191,N_14550);
or UO_503 (O_503,N_14207,N_14078);
nand UO_504 (O_504,N_14179,N_14639);
nor UO_505 (O_505,N_14698,N_14624);
xnor UO_506 (O_506,N_14392,N_14373);
or UO_507 (O_507,N_14189,N_14697);
and UO_508 (O_508,N_14896,N_14476);
and UO_509 (O_509,N_14124,N_14240);
xnor UO_510 (O_510,N_14400,N_14495);
or UO_511 (O_511,N_14116,N_14242);
nand UO_512 (O_512,N_14408,N_14687);
or UO_513 (O_513,N_14169,N_14682);
and UO_514 (O_514,N_14575,N_14982);
nand UO_515 (O_515,N_14612,N_14804);
nand UO_516 (O_516,N_14020,N_14548);
xor UO_517 (O_517,N_14821,N_14208);
xor UO_518 (O_518,N_14023,N_14059);
xor UO_519 (O_519,N_14942,N_14522);
nor UO_520 (O_520,N_14331,N_14718);
or UO_521 (O_521,N_14797,N_14069);
xnor UO_522 (O_522,N_14834,N_14199);
or UO_523 (O_523,N_14196,N_14929);
and UO_524 (O_524,N_14541,N_14618);
nand UO_525 (O_525,N_14504,N_14191);
and UO_526 (O_526,N_14812,N_14794);
nor UO_527 (O_527,N_14696,N_14321);
nand UO_528 (O_528,N_14342,N_14235);
xnor UO_529 (O_529,N_14497,N_14635);
or UO_530 (O_530,N_14827,N_14847);
xnor UO_531 (O_531,N_14416,N_14239);
nand UO_532 (O_532,N_14361,N_14013);
or UO_533 (O_533,N_14731,N_14185);
nand UO_534 (O_534,N_14921,N_14337);
and UO_535 (O_535,N_14738,N_14929);
or UO_536 (O_536,N_14141,N_14702);
nand UO_537 (O_537,N_14585,N_14505);
nor UO_538 (O_538,N_14188,N_14378);
nand UO_539 (O_539,N_14267,N_14897);
xnor UO_540 (O_540,N_14517,N_14124);
xnor UO_541 (O_541,N_14660,N_14292);
or UO_542 (O_542,N_14291,N_14396);
nand UO_543 (O_543,N_14696,N_14145);
and UO_544 (O_544,N_14937,N_14072);
or UO_545 (O_545,N_14339,N_14093);
and UO_546 (O_546,N_14636,N_14175);
and UO_547 (O_547,N_14189,N_14048);
nor UO_548 (O_548,N_14014,N_14146);
and UO_549 (O_549,N_14971,N_14566);
and UO_550 (O_550,N_14697,N_14448);
and UO_551 (O_551,N_14146,N_14642);
or UO_552 (O_552,N_14559,N_14515);
and UO_553 (O_553,N_14295,N_14362);
nand UO_554 (O_554,N_14482,N_14934);
nand UO_555 (O_555,N_14415,N_14297);
nor UO_556 (O_556,N_14025,N_14605);
or UO_557 (O_557,N_14295,N_14911);
and UO_558 (O_558,N_14381,N_14708);
or UO_559 (O_559,N_14261,N_14521);
and UO_560 (O_560,N_14864,N_14596);
and UO_561 (O_561,N_14937,N_14239);
and UO_562 (O_562,N_14612,N_14327);
nor UO_563 (O_563,N_14144,N_14566);
and UO_564 (O_564,N_14791,N_14723);
nand UO_565 (O_565,N_14019,N_14201);
xor UO_566 (O_566,N_14420,N_14433);
nand UO_567 (O_567,N_14805,N_14491);
and UO_568 (O_568,N_14245,N_14415);
nand UO_569 (O_569,N_14775,N_14118);
and UO_570 (O_570,N_14476,N_14976);
xnor UO_571 (O_571,N_14372,N_14514);
and UO_572 (O_572,N_14294,N_14440);
xor UO_573 (O_573,N_14470,N_14145);
nor UO_574 (O_574,N_14663,N_14096);
nor UO_575 (O_575,N_14647,N_14671);
and UO_576 (O_576,N_14437,N_14561);
and UO_577 (O_577,N_14003,N_14944);
xor UO_578 (O_578,N_14249,N_14922);
nand UO_579 (O_579,N_14601,N_14278);
and UO_580 (O_580,N_14687,N_14989);
nor UO_581 (O_581,N_14982,N_14878);
or UO_582 (O_582,N_14125,N_14445);
xor UO_583 (O_583,N_14257,N_14992);
nor UO_584 (O_584,N_14892,N_14778);
and UO_585 (O_585,N_14490,N_14012);
nand UO_586 (O_586,N_14315,N_14109);
or UO_587 (O_587,N_14423,N_14255);
nand UO_588 (O_588,N_14827,N_14452);
or UO_589 (O_589,N_14420,N_14252);
or UO_590 (O_590,N_14989,N_14953);
or UO_591 (O_591,N_14729,N_14536);
xnor UO_592 (O_592,N_14356,N_14454);
nand UO_593 (O_593,N_14458,N_14299);
nand UO_594 (O_594,N_14417,N_14443);
nor UO_595 (O_595,N_14731,N_14643);
xor UO_596 (O_596,N_14401,N_14396);
nor UO_597 (O_597,N_14546,N_14191);
nand UO_598 (O_598,N_14288,N_14477);
nand UO_599 (O_599,N_14886,N_14023);
xnor UO_600 (O_600,N_14122,N_14517);
nand UO_601 (O_601,N_14797,N_14316);
xor UO_602 (O_602,N_14504,N_14763);
or UO_603 (O_603,N_14202,N_14356);
nand UO_604 (O_604,N_14282,N_14378);
xor UO_605 (O_605,N_14138,N_14828);
or UO_606 (O_606,N_14408,N_14224);
nand UO_607 (O_607,N_14261,N_14945);
and UO_608 (O_608,N_14300,N_14081);
or UO_609 (O_609,N_14423,N_14156);
or UO_610 (O_610,N_14487,N_14137);
nor UO_611 (O_611,N_14293,N_14894);
nand UO_612 (O_612,N_14893,N_14771);
and UO_613 (O_613,N_14003,N_14242);
xor UO_614 (O_614,N_14699,N_14332);
nor UO_615 (O_615,N_14418,N_14415);
nand UO_616 (O_616,N_14846,N_14495);
nand UO_617 (O_617,N_14918,N_14398);
nand UO_618 (O_618,N_14869,N_14072);
and UO_619 (O_619,N_14110,N_14295);
xor UO_620 (O_620,N_14082,N_14946);
or UO_621 (O_621,N_14811,N_14757);
nor UO_622 (O_622,N_14158,N_14379);
or UO_623 (O_623,N_14534,N_14793);
or UO_624 (O_624,N_14021,N_14183);
and UO_625 (O_625,N_14444,N_14633);
nor UO_626 (O_626,N_14402,N_14944);
or UO_627 (O_627,N_14418,N_14867);
and UO_628 (O_628,N_14980,N_14411);
nand UO_629 (O_629,N_14826,N_14371);
nor UO_630 (O_630,N_14704,N_14624);
or UO_631 (O_631,N_14591,N_14259);
nand UO_632 (O_632,N_14231,N_14571);
and UO_633 (O_633,N_14056,N_14400);
nand UO_634 (O_634,N_14317,N_14966);
and UO_635 (O_635,N_14141,N_14115);
xor UO_636 (O_636,N_14082,N_14706);
and UO_637 (O_637,N_14057,N_14014);
or UO_638 (O_638,N_14163,N_14329);
and UO_639 (O_639,N_14120,N_14965);
and UO_640 (O_640,N_14640,N_14540);
nor UO_641 (O_641,N_14292,N_14464);
nand UO_642 (O_642,N_14378,N_14063);
nor UO_643 (O_643,N_14388,N_14082);
and UO_644 (O_644,N_14125,N_14863);
nand UO_645 (O_645,N_14228,N_14685);
or UO_646 (O_646,N_14242,N_14394);
and UO_647 (O_647,N_14624,N_14026);
nand UO_648 (O_648,N_14085,N_14714);
nor UO_649 (O_649,N_14243,N_14264);
nor UO_650 (O_650,N_14975,N_14764);
and UO_651 (O_651,N_14203,N_14132);
nor UO_652 (O_652,N_14318,N_14878);
nand UO_653 (O_653,N_14890,N_14731);
nor UO_654 (O_654,N_14470,N_14630);
or UO_655 (O_655,N_14976,N_14004);
or UO_656 (O_656,N_14737,N_14150);
or UO_657 (O_657,N_14329,N_14911);
nand UO_658 (O_658,N_14670,N_14956);
xor UO_659 (O_659,N_14443,N_14231);
xor UO_660 (O_660,N_14686,N_14967);
nor UO_661 (O_661,N_14861,N_14856);
and UO_662 (O_662,N_14136,N_14647);
and UO_663 (O_663,N_14496,N_14134);
nand UO_664 (O_664,N_14396,N_14831);
nor UO_665 (O_665,N_14948,N_14350);
nand UO_666 (O_666,N_14560,N_14565);
nor UO_667 (O_667,N_14116,N_14871);
or UO_668 (O_668,N_14350,N_14601);
nor UO_669 (O_669,N_14650,N_14546);
and UO_670 (O_670,N_14282,N_14177);
xnor UO_671 (O_671,N_14803,N_14804);
nor UO_672 (O_672,N_14232,N_14621);
nand UO_673 (O_673,N_14240,N_14005);
xnor UO_674 (O_674,N_14443,N_14809);
nor UO_675 (O_675,N_14471,N_14509);
nand UO_676 (O_676,N_14278,N_14202);
nor UO_677 (O_677,N_14817,N_14912);
and UO_678 (O_678,N_14947,N_14797);
nor UO_679 (O_679,N_14786,N_14128);
or UO_680 (O_680,N_14373,N_14707);
xor UO_681 (O_681,N_14851,N_14176);
or UO_682 (O_682,N_14472,N_14529);
or UO_683 (O_683,N_14438,N_14257);
and UO_684 (O_684,N_14376,N_14212);
and UO_685 (O_685,N_14783,N_14056);
nand UO_686 (O_686,N_14795,N_14218);
nor UO_687 (O_687,N_14746,N_14127);
or UO_688 (O_688,N_14595,N_14673);
nor UO_689 (O_689,N_14407,N_14606);
or UO_690 (O_690,N_14833,N_14948);
nand UO_691 (O_691,N_14689,N_14961);
and UO_692 (O_692,N_14953,N_14858);
and UO_693 (O_693,N_14385,N_14167);
or UO_694 (O_694,N_14059,N_14511);
nor UO_695 (O_695,N_14982,N_14870);
nor UO_696 (O_696,N_14414,N_14631);
nand UO_697 (O_697,N_14944,N_14780);
and UO_698 (O_698,N_14897,N_14844);
or UO_699 (O_699,N_14110,N_14562);
nor UO_700 (O_700,N_14661,N_14872);
and UO_701 (O_701,N_14865,N_14811);
or UO_702 (O_702,N_14438,N_14753);
and UO_703 (O_703,N_14670,N_14304);
or UO_704 (O_704,N_14046,N_14827);
or UO_705 (O_705,N_14042,N_14205);
and UO_706 (O_706,N_14310,N_14111);
nor UO_707 (O_707,N_14203,N_14274);
nand UO_708 (O_708,N_14470,N_14207);
nor UO_709 (O_709,N_14239,N_14658);
and UO_710 (O_710,N_14118,N_14631);
nor UO_711 (O_711,N_14704,N_14488);
and UO_712 (O_712,N_14578,N_14434);
and UO_713 (O_713,N_14379,N_14639);
nor UO_714 (O_714,N_14878,N_14187);
or UO_715 (O_715,N_14209,N_14268);
nand UO_716 (O_716,N_14233,N_14649);
or UO_717 (O_717,N_14309,N_14979);
nand UO_718 (O_718,N_14926,N_14900);
nor UO_719 (O_719,N_14040,N_14455);
nor UO_720 (O_720,N_14794,N_14018);
and UO_721 (O_721,N_14101,N_14580);
or UO_722 (O_722,N_14056,N_14457);
or UO_723 (O_723,N_14486,N_14206);
or UO_724 (O_724,N_14696,N_14736);
nor UO_725 (O_725,N_14697,N_14684);
nand UO_726 (O_726,N_14221,N_14534);
and UO_727 (O_727,N_14475,N_14304);
nand UO_728 (O_728,N_14426,N_14611);
xor UO_729 (O_729,N_14739,N_14894);
or UO_730 (O_730,N_14002,N_14742);
xnor UO_731 (O_731,N_14704,N_14523);
or UO_732 (O_732,N_14947,N_14179);
and UO_733 (O_733,N_14754,N_14019);
nor UO_734 (O_734,N_14565,N_14347);
nand UO_735 (O_735,N_14787,N_14535);
and UO_736 (O_736,N_14396,N_14841);
and UO_737 (O_737,N_14865,N_14852);
or UO_738 (O_738,N_14138,N_14983);
and UO_739 (O_739,N_14472,N_14000);
nor UO_740 (O_740,N_14553,N_14335);
or UO_741 (O_741,N_14900,N_14852);
nor UO_742 (O_742,N_14506,N_14834);
nand UO_743 (O_743,N_14351,N_14903);
nor UO_744 (O_744,N_14733,N_14848);
nand UO_745 (O_745,N_14502,N_14051);
nand UO_746 (O_746,N_14110,N_14173);
or UO_747 (O_747,N_14948,N_14233);
xor UO_748 (O_748,N_14013,N_14051);
or UO_749 (O_749,N_14817,N_14014);
or UO_750 (O_750,N_14671,N_14558);
nor UO_751 (O_751,N_14657,N_14138);
nor UO_752 (O_752,N_14380,N_14423);
nand UO_753 (O_753,N_14891,N_14366);
xor UO_754 (O_754,N_14656,N_14176);
nand UO_755 (O_755,N_14585,N_14679);
nor UO_756 (O_756,N_14498,N_14456);
or UO_757 (O_757,N_14579,N_14980);
nand UO_758 (O_758,N_14421,N_14482);
nor UO_759 (O_759,N_14049,N_14336);
nand UO_760 (O_760,N_14462,N_14545);
nor UO_761 (O_761,N_14356,N_14668);
nor UO_762 (O_762,N_14453,N_14389);
nand UO_763 (O_763,N_14852,N_14572);
nand UO_764 (O_764,N_14354,N_14239);
and UO_765 (O_765,N_14237,N_14536);
and UO_766 (O_766,N_14937,N_14226);
or UO_767 (O_767,N_14411,N_14601);
or UO_768 (O_768,N_14624,N_14554);
or UO_769 (O_769,N_14419,N_14858);
and UO_770 (O_770,N_14858,N_14732);
nand UO_771 (O_771,N_14124,N_14322);
and UO_772 (O_772,N_14788,N_14065);
xnor UO_773 (O_773,N_14631,N_14317);
or UO_774 (O_774,N_14501,N_14598);
nor UO_775 (O_775,N_14072,N_14475);
nand UO_776 (O_776,N_14877,N_14819);
and UO_777 (O_777,N_14840,N_14366);
and UO_778 (O_778,N_14931,N_14874);
nand UO_779 (O_779,N_14335,N_14000);
or UO_780 (O_780,N_14430,N_14304);
and UO_781 (O_781,N_14533,N_14159);
nor UO_782 (O_782,N_14939,N_14996);
nor UO_783 (O_783,N_14261,N_14975);
or UO_784 (O_784,N_14938,N_14530);
nor UO_785 (O_785,N_14949,N_14063);
and UO_786 (O_786,N_14777,N_14210);
xnor UO_787 (O_787,N_14968,N_14672);
nand UO_788 (O_788,N_14931,N_14939);
xor UO_789 (O_789,N_14895,N_14448);
nor UO_790 (O_790,N_14636,N_14329);
nand UO_791 (O_791,N_14989,N_14054);
nand UO_792 (O_792,N_14879,N_14911);
nor UO_793 (O_793,N_14247,N_14408);
nand UO_794 (O_794,N_14917,N_14710);
nand UO_795 (O_795,N_14713,N_14541);
nand UO_796 (O_796,N_14667,N_14719);
and UO_797 (O_797,N_14820,N_14269);
or UO_798 (O_798,N_14175,N_14026);
or UO_799 (O_799,N_14570,N_14822);
nor UO_800 (O_800,N_14242,N_14206);
and UO_801 (O_801,N_14721,N_14356);
nand UO_802 (O_802,N_14899,N_14770);
and UO_803 (O_803,N_14403,N_14657);
nand UO_804 (O_804,N_14936,N_14128);
nor UO_805 (O_805,N_14801,N_14481);
and UO_806 (O_806,N_14347,N_14863);
or UO_807 (O_807,N_14118,N_14504);
nor UO_808 (O_808,N_14484,N_14615);
nor UO_809 (O_809,N_14758,N_14306);
or UO_810 (O_810,N_14765,N_14858);
and UO_811 (O_811,N_14681,N_14370);
and UO_812 (O_812,N_14270,N_14622);
nor UO_813 (O_813,N_14451,N_14063);
or UO_814 (O_814,N_14300,N_14221);
or UO_815 (O_815,N_14820,N_14765);
nor UO_816 (O_816,N_14920,N_14047);
xnor UO_817 (O_817,N_14181,N_14337);
and UO_818 (O_818,N_14470,N_14536);
or UO_819 (O_819,N_14497,N_14364);
or UO_820 (O_820,N_14659,N_14647);
nor UO_821 (O_821,N_14850,N_14053);
nor UO_822 (O_822,N_14913,N_14344);
nor UO_823 (O_823,N_14677,N_14861);
nor UO_824 (O_824,N_14942,N_14556);
and UO_825 (O_825,N_14024,N_14742);
nand UO_826 (O_826,N_14340,N_14424);
xnor UO_827 (O_827,N_14016,N_14372);
and UO_828 (O_828,N_14823,N_14130);
nor UO_829 (O_829,N_14906,N_14708);
nand UO_830 (O_830,N_14178,N_14668);
nor UO_831 (O_831,N_14887,N_14526);
and UO_832 (O_832,N_14937,N_14733);
nor UO_833 (O_833,N_14696,N_14763);
nand UO_834 (O_834,N_14217,N_14416);
or UO_835 (O_835,N_14024,N_14436);
nor UO_836 (O_836,N_14964,N_14473);
nor UO_837 (O_837,N_14524,N_14339);
nand UO_838 (O_838,N_14496,N_14533);
nor UO_839 (O_839,N_14435,N_14804);
or UO_840 (O_840,N_14072,N_14667);
nor UO_841 (O_841,N_14250,N_14168);
nor UO_842 (O_842,N_14533,N_14967);
nor UO_843 (O_843,N_14467,N_14230);
nand UO_844 (O_844,N_14493,N_14470);
and UO_845 (O_845,N_14788,N_14038);
nand UO_846 (O_846,N_14006,N_14424);
and UO_847 (O_847,N_14111,N_14429);
and UO_848 (O_848,N_14460,N_14695);
nand UO_849 (O_849,N_14685,N_14528);
nor UO_850 (O_850,N_14182,N_14294);
nor UO_851 (O_851,N_14768,N_14195);
or UO_852 (O_852,N_14093,N_14883);
nor UO_853 (O_853,N_14297,N_14480);
xnor UO_854 (O_854,N_14634,N_14540);
and UO_855 (O_855,N_14250,N_14993);
and UO_856 (O_856,N_14708,N_14705);
or UO_857 (O_857,N_14218,N_14738);
xnor UO_858 (O_858,N_14191,N_14442);
and UO_859 (O_859,N_14759,N_14524);
xnor UO_860 (O_860,N_14228,N_14283);
xor UO_861 (O_861,N_14589,N_14886);
and UO_862 (O_862,N_14795,N_14045);
or UO_863 (O_863,N_14717,N_14880);
and UO_864 (O_864,N_14900,N_14425);
and UO_865 (O_865,N_14687,N_14361);
or UO_866 (O_866,N_14027,N_14450);
nor UO_867 (O_867,N_14924,N_14572);
nand UO_868 (O_868,N_14122,N_14240);
or UO_869 (O_869,N_14308,N_14861);
and UO_870 (O_870,N_14435,N_14927);
and UO_871 (O_871,N_14041,N_14469);
nand UO_872 (O_872,N_14199,N_14288);
and UO_873 (O_873,N_14044,N_14865);
or UO_874 (O_874,N_14322,N_14305);
or UO_875 (O_875,N_14711,N_14830);
xor UO_876 (O_876,N_14140,N_14202);
and UO_877 (O_877,N_14193,N_14173);
nor UO_878 (O_878,N_14496,N_14082);
or UO_879 (O_879,N_14201,N_14948);
xor UO_880 (O_880,N_14812,N_14574);
nand UO_881 (O_881,N_14533,N_14477);
nor UO_882 (O_882,N_14249,N_14349);
and UO_883 (O_883,N_14940,N_14661);
or UO_884 (O_884,N_14870,N_14696);
or UO_885 (O_885,N_14647,N_14395);
or UO_886 (O_886,N_14509,N_14782);
and UO_887 (O_887,N_14774,N_14037);
xor UO_888 (O_888,N_14377,N_14972);
nor UO_889 (O_889,N_14779,N_14605);
nand UO_890 (O_890,N_14790,N_14353);
and UO_891 (O_891,N_14375,N_14379);
nand UO_892 (O_892,N_14165,N_14781);
or UO_893 (O_893,N_14815,N_14138);
nand UO_894 (O_894,N_14092,N_14366);
nor UO_895 (O_895,N_14598,N_14369);
nand UO_896 (O_896,N_14963,N_14096);
xnor UO_897 (O_897,N_14104,N_14871);
or UO_898 (O_898,N_14890,N_14960);
and UO_899 (O_899,N_14181,N_14674);
nand UO_900 (O_900,N_14116,N_14341);
or UO_901 (O_901,N_14655,N_14307);
or UO_902 (O_902,N_14881,N_14777);
nor UO_903 (O_903,N_14309,N_14465);
nand UO_904 (O_904,N_14279,N_14402);
nand UO_905 (O_905,N_14123,N_14708);
nor UO_906 (O_906,N_14753,N_14218);
and UO_907 (O_907,N_14630,N_14506);
nor UO_908 (O_908,N_14891,N_14597);
nand UO_909 (O_909,N_14987,N_14826);
nand UO_910 (O_910,N_14876,N_14808);
or UO_911 (O_911,N_14803,N_14517);
and UO_912 (O_912,N_14940,N_14480);
nor UO_913 (O_913,N_14509,N_14034);
nor UO_914 (O_914,N_14753,N_14555);
xnor UO_915 (O_915,N_14748,N_14787);
nand UO_916 (O_916,N_14633,N_14173);
or UO_917 (O_917,N_14459,N_14359);
nand UO_918 (O_918,N_14294,N_14583);
nor UO_919 (O_919,N_14092,N_14442);
and UO_920 (O_920,N_14889,N_14328);
nor UO_921 (O_921,N_14969,N_14238);
and UO_922 (O_922,N_14245,N_14149);
nand UO_923 (O_923,N_14339,N_14520);
and UO_924 (O_924,N_14370,N_14640);
nand UO_925 (O_925,N_14953,N_14567);
or UO_926 (O_926,N_14395,N_14132);
nor UO_927 (O_927,N_14540,N_14129);
and UO_928 (O_928,N_14657,N_14964);
or UO_929 (O_929,N_14248,N_14167);
nand UO_930 (O_930,N_14702,N_14534);
nor UO_931 (O_931,N_14173,N_14592);
xnor UO_932 (O_932,N_14552,N_14522);
xor UO_933 (O_933,N_14625,N_14182);
or UO_934 (O_934,N_14223,N_14904);
nand UO_935 (O_935,N_14929,N_14494);
nor UO_936 (O_936,N_14751,N_14443);
or UO_937 (O_937,N_14641,N_14954);
nand UO_938 (O_938,N_14529,N_14364);
and UO_939 (O_939,N_14916,N_14316);
nand UO_940 (O_940,N_14899,N_14702);
and UO_941 (O_941,N_14805,N_14110);
and UO_942 (O_942,N_14851,N_14192);
xnor UO_943 (O_943,N_14195,N_14133);
and UO_944 (O_944,N_14119,N_14652);
xor UO_945 (O_945,N_14428,N_14088);
nand UO_946 (O_946,N_14208,N_14427);
and UO_947 (O_947,N_14901,N_14182);
nand UO_948 (O_948,N_14972,N_14472);
or UO_949 (O_949,N_14656,N_14803);
and UO_950 (O_950,N_14440,N_14199);
nor UO_951 (O_951,N_14195,N_14367);
and UO_952 (O_952,N_14761,N_14971);
or UO_953 (O_953,N_14117,N_14619);
and UO_954 (O_954,N_14281,N_14081);
and UO_955 (O_955,N_14837,N_14792);
nand UO_956 (O_956,N_14652,N_14774);
nand UO_957 (O_957,N_14003,N_14315);
nor UO_958 (O_958,N_14624,N_14369);
nand UO_959 (O_959,N_14134,N_14004);
and UO_960 (O_960,N_14925,N_14757);
xnor UO_961 (O_961,N_14729,N_14906);
and UO_962 (O_962,N_14998,N_14899);
nor UO_963 (O_963,N_14687,N_14695);
or UO_964 (O_964,N_14369,N_14552);
and UO_965 (O_965,N_14483,N_14015);
nor UO_966 (O_966,N_14539,N_14323);
nand UO_967 (O_967,N_14472,N_14539);
or UO_968 (O_968,N_14292,N_14809);
nor UO_969 (O_969,N_14209,N_14854);
xnor UO_970 (O_970,N_14315,N_14378);
nand UO_971 (O_971,N_14732,N_14282);
or UO_972 (O_972,N_14700,N_14624);
nor UO_973 (O_973,N_14512,N_14649);
nor UO_974 (O_974,N_14222,N_14324);
nor UO_975 (O_975,N_14779,N_14765);
and UO_976 (O_976,N_14781,N_14548);
xor UO_977 (O_977,N_14315,N_14609);
and UO_978 (O_978,N_14025,N_14594);
nor UO_979 (O_979,N_14842,N_14360);
and UO_980 (O_980,N_14548,N_14766);
nor UO_981 (O_981,N_14311,N_14714);
nand UO_982 (O_982,N_14106,N_14165);
or UO_983 (O_983,N_14069,N_14431);
nor UO_984 (O_984,N_14999,N_14397);
or UO_985 (O_985,N_14776,N_14822);
or UO_986 (O_986,N_14274,N_14715);
or UO_987 (O_987,N_14617,N_14494);
xor UO_988 (O_988,N_14276,N_14409);
nor UO_989 (O_989,N_14255,N_14298);
and UO_990 (O_990,N_14940,N_14369);
nand UO_991 (O_991,N_14466,N_14987);
nand UO_992 (O_992,N_14109,N_14025);
or UO_993 (O_993,N_14278,N_14986);
xnor UO_994 (O_994,N_14307,N_14856);
nor UO_995 (O_995,N_14084,N_14377);
nand UO_996 (O_996,N_14333,N_14435);
or UO_997 (O_997,N_14681,N_14224);
and UO_998 (O_998,N_14368,N_14141);
nor UO_999 (O_999,N_14184,N_14534);
nor UO_1000 (O_1000,N_14266,N_14482);
nor UO_1001 (O_1001,N_14889,N_14732);
xnor UO_1002 (O_1002,N_14742,N_14398);
and UO_1003 (O_1003,N_14504,N_14403);
nand UO_1004 (O_1004,N_14698,N_14992);
or UO_1005 (O_1005,N_14138,N_14986);
xnor UO_1006 (O_1006,N_14696,N_14013);
nand UO_1007 (O_1007,N_14714,N_14673);
or UO_1008 (O_1008,N_14538,N_14364);
nand UO_1009 (O_1009,N_14623,N_14475);
nor UO_1010 (O_1010,N_14029,N_14124);
and UO_1011 (O_1011,N_14908,N_14803);
and UO_1012 (O_1012,N_14894,N_14112);
or UO_1013 (O_1013,N_14153,N_14706);
nor UO_1014 (O_1014,N_14263,N_14193);
and UO_1015 (O_1015,N_14066,N_14063);
nor UO_1016 (O_1016,N_14068,N_14150);
nor UO_1017 (O_1017,N_14441,N_14470);
or UO_1018 (O_1018,N_14226,N_14431);
or UO_1019 (O_1019,N_14539,N_14099);
or UO_1020 (O_1020,N_14663,N_14940);
or UO_1021 (O_1021,N_14831,N_14665);
and UO_1022 (O_1022,N_14969,N_14972);
nor UO_1023 (O_1023,N_14264,N_14770);
and UO_1024 (O_1024,N_14657,N_14694);
or UO_1025 (O_1025,N_14159,N_14551);
nor UO_1026 (O_1026,N_14508,N_14399);
and UO_1027 (O_1027,N_14899,N_14265);
and UO_1028 (O_1028,N_14540,N_14957);
or UO_1029 (O_1029,N_14105,N_14264);
nand UO_1030 (O_1030,N_14061,N_14170);
or UO_1031 (O_1031,N_14594,N_14389);
or UO_1032 (O_1032,N_14977,N_14377);
and UO_1033 (O_1033,N_14123,N_14168);
and UO_1034 (O_1034,N_14842,N_14109);
xnor UO_1035 (O_1035,N_14134,N_14681);
or UO_1036 (O_1036,N_14081,N_14924);
nand UO_1037 (O_1037,N_14552,N_14328);
or UO_1038 (O_1038,N_14499,N_14758);
or UO_1039 (O_1039,N_14135,N_14730);
or UO_1040 (O_1040,N_14760,N_14046);
xnor UO_1041 (O_1041,N_14631,N_14717);
and UO_1042 (O_1042,N_14313,N_14784);
nor UO_1043 (O_1043,N_14005,N_14505);
nor UO_1044 (O_1044,N_14530,N_14227);
nor UO_1045 (O_1045,N_14258,N_14622);
nand UO_1046 (O_1046,N_14656,N_14865);
nor UO_1047 (O_1047,N_14593,N_14259);
nor UO_1048 (O_1048,N_14404,N_14980);
nor UO_1049 (O_1049,N_14624,N_14099);
and UO_1050 (O_1050,N_14100,N_14011);
and UO_1051 (O_1051,N_14438,N_14504);
nor UO_1052 (O_1052,N_14805,N_14237);
or UO_1053 (O_1053,N_14193,N_14052);
or UO_1054 (O_1054,N_14448,N_14647);
nand UO_1055 (O_1055,N_14299,N_14901);
and UO_1056 (O_1056,N_14353,N_14083);
xnor UO_1057 (O_1057,N_14671,N_14668);
and UO_1058 (O_1058,N_14873,N_14985);
nor UO_1059 (O_1059,N_14473,N_14937);
or UO_1060 (O_1060,N_14818,N_14669);
and UO_1061 (O_1061,N_14229,N_14300);
or UO_1062 (O_1062,N_14429,N_14945);
and UO_1063 (O_1063,N_14531,N_14832);
nand UO_1064 (O_1064,N_14243,N_14712);
nand UO_1065 (O_1065,N_14731,N_14591);
nor UO_1066 (O_1066,N_14132,N_14274);
nor UO_1067 (O_1067,N_14733,N_14203);
and UO_1068 (O_1068,N_14028,N_14999);
nand UO_1069 (O_1069,N_14723,N_14072);
nand UO_1070 (O_1070,N_14198,N_14366);
and UO_1071 (O_1071,N_14307,N_14607);
nor UO_1072 (O_1072,N_14137,N_14904);
nor UO_1073 (O_1073,N_14331,N_14894);
or UO_1074 (O_1074,N_14090,N_14829);
nor UO_1075 (O_1075,N_14663,N_14694);
nor UO_1076 (O_1076,N_14772,N_14641);
or UO_1077 (O_1077,N_14097,N_14770);
nand UO_1078 (O_1078,N_14536,N_14153);
nand UO_1079 (O_1079,N_14283,N_14989);
nor UO_1080 (O_1080,N_14761,N_14923);
nor UO_1081 (O_1081,N_14591,N_14483);
and UO_1082 (O_1082,N_14357,N_14529);
or UO_1083 (O_1083,N_14515,N_14918);
and UO_1084 (O_1084,N_14896,N_14528);
nor UO_1085 (O_1085,N_14823,N_14418);
and UO_1086 (O_1086,N_14258,N_14525);
or UO_1087 (O_1087,N_14754,N_14349);
xor UO_1088 (O_1088,N_14153,N_14753);
nor UO_1089 (O_1089,N_14147,N_14549);
xor UO_1090 (O_1090,N_14080,N_14738);
nand UO_1091 (O_1091,N_14176,N_14115);
nand UO_1092 (O_1092,N_14704,N_14123);
nor UO_1093 (O_1093,N_14512,N_14811);
or UO_1094 (O_1094,N_14179,N_14444);
nand UO_1095 (O_1095,N_14793,N_14569);
and UO_1096 (O_1096,N_14824,N_14317);
and UO_1097 (O_1097,N_14621,N_14426);
or UO_1098 (O_1098,N_14058,N_14082);
and UO_1099 (O_1099,N_14101,N_14694);
and UO_1100 (O_1100,N_14971,N_14059);
or UO_1101 (O_1101,N_14783,N_14632);
nand UO_1102 (O_1102,N_14576,N_14545);
and UO_1103 (O_1103,N_14481,N_14107);
nand UO_1104 (O_1104,N_14645,N_14413);
and UO_1105 (O_1105,N_14543,N_14090);
nor UO_1106 (O_1106,N_14413,N_14058);
and UO_1107 (O_1107,N_14626,N_14237);
or UO_1108 (O_1108,N_14973,N_14720);
nand UO_1109 (O_1109,N_14633,N_14867);
and UO_1110 (O_1110,N_14668,N_14484);
or UO_1111 (O_1111,N_14232,N_14888);
nand UO_1112 (O_1112,N_14878,N_14575);
and UO_1113 (O_1113,N_14360,N_14309);
or UO_1114 (O_1114,N_14257,N_14337);
or UO_1115 (O_1115,N_14029,N_14430);
nand UO_1116 (O_1116,N_14903,N_14973);
xnor UO_1117 (O_1117,N_14058,N_14018);
and UO_1118 (O_1118,N_14509,N_14437);
nand UO_1119 (O_1119,N_14957,N_14775);
nor UO_1120 (O_1120,N_14761,N_14658);
xnor UO_1121 (O_1121,N_14260,N_14276);
xor UO_1122 (O_1122,N_14267,N_14094);
xnor UO_1123 (O_1123,N_14028,N_14817);
nor UO_1124 (O_1124,N_14126,N_14636);
xor UO_1125 (O_1125,N_14337,N_14239);
or UO_1126 (O_1126,N_14227,N_14573);
and UO_1127 (O_1127,N_14510,N_14157);
nor UO_1128 (O_1128,N_14069,N_14705);
and UO_1129 (O_1129,N_14541,N_14139);
or UO_1130 (O_1130,N_14063,N_14424);
nand UO_1131 (O_1131,N_14576,N_14568);
nand UO_1132 (O_1132,N_14878,N_14238);
and UO_1133 (O_1133,N_14330,N_14956);
nand UO_1134 (O_1134,N_14843,N_14410);
or UO_1135 (O_1135,N_14055,N_14210);
and UO_1136 (O_1136,N_14860,N_14652);
or UO_1137 (O_1137,N_14498,N_14014);
nor UO_1138 (O_1138,N_14546,N_14889);
and UO_1139 (O_1139,N_14831,N_14578);
nand UO_1140 (O_1140,N_14061,N_14914);
nand UO_1141 (O_1141,N_14352,N_14252);
nand UO_1142 (O_1142,N_14576,N_14899);
nor UO_1143 (O_1143,N_14150,N_14274);
and UO_1144 (O_1144,N_14917,N_14562);
nor UO_1145 (O_1145,N_14728,N_14815);
nor UO_1146 (O_1146,N_14668,N_14298);
or UO_1147 (O_1147,N_14477,N_14806);
nor UO_1148 (O_1148,N_14765,N_14662);
nand UO_1149 (O_1149,N_14753,N_14510);
nand UO_1150 (O_1150,N_14211,N_14176);
and UO_1151 (O_1151,N_14208,N_14290);
nor UO_1152 (O_1152,N_14239,N_14805);
nor UO_1153 (O_1153,N_14026,N_14453);
or UO_1154 (O_1154,N_14198,N_14841);
nor UO_1155 (O_1155,N_14518,N_14645);
and UO_1156 (O_1156,N_14149,N_14990);
nor UO_1157 (O_1157,N_14361,N_14114);
and UO_1158 (O_1158,N_14686,N_14840);
or UO_1159 (O_1159,N_14856,N_14475);
nand UO_1160 (O_1160,N_14451,N_14987);
and UO_1161 (O_1161,N_14569,N_14450);
nor UO_1162 (O_1162,N_14294,N_14022);
and UO_1163 (O_1163,N_14633,N_14921);
nand UO_1164 (O_1164,N_14996,N_14683);
or UO_1165 (O_1165,N_14564,N_14890);
nor UO_1166 (O_1166,N_14895,N_14748);
nor UO_1167 (O_1167,N_14583,N_14201);
nand UO_1168 (O_1168,N_14519,N_14554);
and UO_1169 (O_1169,N_14552,N_14803);
nand UO_1170 (O_1170,N_14394,N_14701);
xor UO_1171 (O_1171,N_14745,N_14586);
or UO_1172 (O_1172,N_14863,N_14784);
and UO_1173 (O_1173,N_14239,N_14573);
and UO_1174 (O_1174,N_14058,N_14729);
or UO_1175 (O_1175,N_14385,N_14828);
and UO_1176 (O_1176,N_14047,N_14186);
nor UO_1177 (O_1177,N_14727,N_14970);
and UO_1178 (O_1178,N_14862,N_14871);
or UO_1179 (O_1179,N_14671,N_14672);
or UO_1180 (O_1180,N_14337,N_14630);
nand UO_1181 (O_1181,N_14315,N_14882);
and UO_1182 (O_1182,N_14157,N_14233);
or UO_1183 (O_1183,N_14307,N_14767);
nand UO_1184 (O_1184,N_14946,N_14362);
nor UO_1185 (O_1185,N_14908,N_14920);
and UO_1186 (O_1186,N_14172,N_14148);
nand UO_1187 (O_1187,N_14268,N_14372);
nor UO_1188 (O_1188,N_14819,N_14044);
nor UO_1189 (O_1189,N_14312,N_14572);
xnor UO_1190 (O_1190,N_14727,N_14690);
nand UO_1191 (O_1191,N_14062,N_14354);
nand UO_1192 (O_1192,N_14681,N_14772);
and UO_1193 (O_1193,N_14657,N_14398);
and UO_1194 (O_1194,N_14773,N_14210);
nand UO_1195 (O_1195,N_14441,N_14342);
or UO_1196 (O_1196,N_14307,N_14461);
nand UO_1197 (O_1197,N_14023,N_14007);
or UO_1198 (O_1198,N_14595,N_14399);
nor UO_1199 (O_1199,N_14265,N_14663);
xor UO_1200 (O_1200,N_14175,N_14807);
nand UO_1201 (O_1201,N_14282,N_14729);
and UO_1202 (O_1202,N_14291,N_14203);
nor UO_1203 (O_1203,N_14098,N_14476);
xor UO_1204 (O_1204,N_14619,N_14742);
nor UO_1205 (O_1205,N_14822,N_14401);
or UO_1206 (O_1206,N_14996,N_14993);
nor UO_1207 (O_1207,N_14105,N_14769);
or UO_1208 (O_1208,N_14176,N_14195);
nor UO_1209 (O_1209,N_14943,N_14647);
nand UO_1210 (O_1210,N_14776,N_14554);
or UO_1211 (O_1211,N_14698,N_14960);
or UO_1212 (O_1212,N_14010,N_14766);
and UO_1213 (O_1213,N_14928,N_14971);
nor UO_1214 (O_1214,N_14004,N_14268);
or UO_1215 (O_1215,N_14423,N_14522);
nand UO_1216 (O_1216,N_14742,N_14056);
nand UO_1217 (O_1217,N_14762,N_14144);
nand UO_1218 (O_1218,N_14988,N_14472);
and UO_1219 (O_1219,N_14993,N_14152);
or UO_1220 (O_1220,N_14960,N_14962);
xnor UO_1221 (O_1221,N_14827,N_14113);
nand UO_1222 (O_1222,N_14475,N_14646);
and UO_1223 (O_1223,N_14897,N_14492);
xor UO_1224 (O_1224,N_14747,N_14308);
and UO_1225 (O_1225,N_14855,N_14144);
nand UO_1226 (O_1226,N_14542,N_14693);
xor UO_1227 (O_1227,N_14556,N_14367);
or UO_1228 (O_1228,N_14542,N_14198);
and UO_1229 (O_1229,N_14733,N_14592);
nor UO_1230 (O_1230,N_14748,N_14419);
nor UO_1231 (O_1231,N_14923,N_14240);
and UO_1232 (O_1232,N_14740,N_14042);
or UO_1233 (O_1233,N_14640,N_14199);
or UO_1234 (O_1234,N_14586,N_14482);
and UO_1235 (O_1235,N_14769,N_14682);
nand UO_1236 (O_1236,N_14441,N_14212);
or UO_1237 (O_1237,N_14327,N_14453);
nand UO_1238 (O_1238,N_14741,N_14843);
nand UO_1239 (O_1239,N_14825,N_14153);
xor UO_1240 (O_1240,N_14269,N_14186);
xor UO_1241 (O_1241,N_14128,N_14837);
nor UO_1242 (O_1242,N_14910,N_14891);
xnor UO_1243 (O_1243,N_14239,N_14107);
or UO_1244 (O_1244,N_14056,N_14598);
or UO_1245 (O_1245,N_14327,N_14853);
nor UO_1246 (O_1246,N_14851,N_14928);
xor UO_1247 (O_1247,N_14048,N_14416);
or UO_1248 (O_1248,N_14351,N_14291);
xor UO_1249 (O_1249,N_14752,N_14848);
and UO_1250 (O_1250,N_14813,N_14982);
nor UO_1251 (O_1251,N_14863,N_14688);
or UO_1252 (O_1252,N_14977,N_14351);
and UO_1253 (O_1253,N_14138,N_14353);
nand UO_1254 (O_1254,N_14257,N_14323);
and UO_1255 (O_1255,N_14896,N_14168);
and UO_1256 (O_1256,N_14634,N_14562);
and UO_1257 (O_1257,N_14302,N_14380);
nand UO_1258 (O_1258,N_14557,N_14664);
or UO_1259 (O_1259,N_14392,N_14951);
nor UO_1260 (O_1260,N_14507,N_14653);
or UO_1261 (O_1261,N_14829,N_14497);
nor UO_1262 (O_1262,N_14998,N_14550);
or UO_1263 (O_1263,N_14749,N_14456);
or UO_1264 (O_1264,N_14855,N_14088);
nand UO_1265 (O_1265,N_14598,N_14952);
nor UO_1266 (O_1266,N_14779,N_14252);
and UO_1267 (O_1267,N_14291,N_14269);
and UO_1268 (O_1268,N_14539,N_14029);
nor UO_1269 (O_1269,N_14896,N_14651);
nor UO_1270 (O_1270,N_14826,N_14354);
nor UO_1271 (O_1271,N_14611,N_14489);
and UO_1272 (O_1272,N_14783,N_14838);
and UO_1273 (O_1273,N_14649,N_14070);
and UO_1274 (O_1274,N_14646,N_14003);
nand UO_1275 (O_1275,N_14533,N_14105);
or UO_1276 (O_1276,N_14918,N_14860);
nand UO_1277 (O_1277,N_14160,N_14997);
nor UO_1278 (O_1278,N_14873,N_14310);
nor UO_1279 (O_1279,N_14032,N_14137);
nand UO_1280 (O_1280,N_14958,N_14432);
xor UO_1281 (O_1281,N_14065,N_14197);
or UO_1282 (O_1282,N_14282,N_14605);
xnor UO_1283 (O_1283,N_14847,N_14329);
nand UO_1284 (O_1284,N_14202,N_14237);
and UO_1285 (O_1285,N_14929,N_14541);
or UO_1286 (O_1286,N_14903,N_14207);
or UO_1287 (O_1287,N_14523,N_14529);
nand UO_1288 (O_1288,N_14286,N_14761);
and UO_1289 (O_1289,N_14127,N_14318);
and UO_1290 (O_1290,N_14986,N_14560);
nor UO_1291 (O_1291,N_14973,N_14772);
nand UO_1292 (O_1292,N_14602,N_14054);
and UO_1293 (O_1293,N_14326,N_14618);
nand UO_1294 (O_1294,N_14373,N_14983);
nor UO_1295 (O_1295,N_14302,N_14382);
and UO_1296 (O_1296,N_14723,N_14411);
nand UO_1297 (O_1297,N_14410,N_14086);
or UO_1298 (O_1298,N_14963,N_14765);
xnor UO_1299 (O_1299,N_14820,N_14998);
xor UO_1300 (O_1300,N_14711,N_14717);
nor UO_1301 (O_1301,N_14630,N_14416);
and UO_1302 (O_1302,N_14066,N_14041);
and UO_1303 (O_1303,N_14463,N_14555);
or UO_1304 (O_1304,N_14380,N_14417);
or UO_1305 (O_1305,N_14078,N_14103);
and UO_1306 (O_1306,N_14968,N_14039);
or UO_1307 (O_1307,N_14836,N_14754);
or UO_1308 (O_1308,N_14345,N_14366);
or UO_1309 (O_1309,N_14356,N_14938);
nand UO_1310 (O_1310,N_14738,N_14168);
nand UO_1311 (O_1311,N_14923,N_14250);
nand UO_1312 (O_1312,N_14787,N_14530);
xnor UO_1313 (O_1313,N_14672,N_14516);
and UO_1314 (O_1314,N_14521,N_14885);
or UO_1315 (O_1315,N_14238,N_14914);
or UO_1316 (O_1316,N_14103,N_14557);
and UO_1317 (O_1317,N_14196,N_14974);
nor UO_1318 (O_1318,N_14665,N_14807);
nand UO_1319 (O_1319,N_14487,N_14883);
nor UO_1320 (O_1320,N_14783,N_14080);
and UO_1321 (O_1321,N_14799,N_14033);
xnor UO_1322 (O_1322,N_14311,N_14249);
and UO_1323 (O_1323,N_14799,N_14573);
nor UO_1324 (O_1324,N_14343,N_14154);
and UO_1325 (O_1325,N_14807,N_14572);
and UO_1326 (O_1326,N_14422,N_14437);
nor UO_1327 (O_1327,N_14184,N_14466);
nor UO_1328 (O_1328,N_14557,N_14804);
nor UO_1329 (O_1329,N_14414,N_14841);
and UO_1330 (O_1330,N_14525,N_14714);
and UO_1331 (O_1331,N_14552,N_14643);
nand UO_1332 (O_1332,N_14245,N_14528);
nand UO_1333 (O_1333,N_14435,N_14446);
nor UO_1334 (O_1334,N_14134,N_14654);
nor UO_1335 (O_1335,N_14422,N_14241);
nor UO_1336 (O_1336,N_14596,N_14873);
nor UO_1337 (O_1337,N_14203,N_14792);
nor UO_1338 (O_1338,N_14477,N_14368);
or UO_1339 (O_1339,N_14698,N_14421);
or UO_1340 (O_1340,N_14455,N_14294);
or UO_1341 (O_1341,N_14783,N_14649);
nand UO_1342 (O_1342,N_14873,N_14763);
and UO_1343 (O_1343,N_14957,N_14803);
or UO_1344 (O_1344,N_14811,N_14036);
nor UO_1345 (O_1345,N_14921,N_14889);
and UO_1346 (O_1346,N_14580,N_14253);
and UO_1347 (O_1347,N_14795,N_14712);
xor UO_1348 (O_1348,N_14410,N_14655);
and UO_1349 (O_1349,N_14253,N_14264);
and UO_1350 (O_1350,N_14250,N_14333);
and UO_1351 (O_1351,N_14203,N_14450);
and UO_1352 (O_1352,N_14828,N_14444);
or UO_1353 (O_1353,N_14344,N_14032);
nor UO_1354 (O_1354,N_14870,N_14024);
or UO_1355 (O_1355,N_14646,N_14883);
nor UO_1356 (O_1356,N_14991,N_14587);
and UO_1357 (O_1357,N_14850,N_14140);
and UO_1358 (O_1358,N_14631,N_14703);
xnor UO_1359 (O_1359,N_14206,N_14605);
and UO_1360 (O_1360,N_14434,N_14516);
and UO_1361 (O_1361,N_14968,N_14483);
xnor UO_1362 (O_1362,N_14800,N_14124);
xor UO_1363 (O_1363,N_14000,N_14784);
or UO_1364 (O_1364,N_14439,N_14944);
nand UO_1365 (O_1365,N_14949,N_14231);
and UO_1366 (O_1366,N_14345,N_14325);
nor UO_1367 (O_1367,N_14751,N_14933);
xnor UO_1368 (O_1368,N_14180,N_14386);
nand UO_1369 (O_1369,N_14635,N_14747);
nor UO_1370 (O_1370,N_14119,N_14717);
xor UO_1371 (O_1371,N_14733,N_14582);
nand UO_1372 (O_1372,N_14203,N_14909);
or UO_1373 (O_1373,N_14695,N_14148);
and UO_1374 (O_1374,N_14456,N_14155);
nand UO_1375 (O_1375,N_14152,N_14052);
or UO_1376 (O_1376,N_14535,N_14100);
and UO_1377 (O_1377,N_14751,N_14198);
or UO_1378 (O_1378,N_14300,N_14757);
and UO_1379 (O_1379,N_14684,N_14519);
nor UO_1380 (O_1380,N_14810,N_14568);
or UO_1381 (O_1381,N_14197,N_14264);
and UO_1382 (O_1382,N_14092,N_14170);
nor UO_1383 (O_1383,N_14506,N_14614);
nor UO_1384 (O_1384,N_14881,N_14036);
nor UO_1385 (O_1385,N_14335,N_14846);
xor UO_1386 (O_1386,N_14090,N_14900);
and UO_1387 (O_1387,N_14592,N_14601);
nand UO_1388 (O_1388,N_14486,N_14154);
or UO_1389 (O_1389,N_14062,N_14226);
nand UO_1390 (O_1390,N_14607,N_14000);
xnor UO_1391 (O_1391,N_14885,N_14605);
xnor UO_1392 (O_1392,N_14910,N_14790);
nor UO_1393 (O_1393,N_14349,N_14117);
nor UO_1394 (O_1394,N_14992,N_14774);
and UO_1395 (O_1395,N_14304,N_14483);
nor UO_1396 (O_1396,N_14805,N_14511);
or UO_1397 (O_1397,N_14769,N_14859);
and UO_1398 (O_1398,N_14476,N_14123);
xnor UO_1399 (O_1399,N_14348,N_14717);
and UO_1400 (O_1400,N_14778,N_14860);
or UO_1401 (O_1401,N_14770,N_14046);
nand UO_1402 (O_1402,N_14174,N_14673);
nand UO_1403 (O_1403,N_14814,N_14505);
and UO_1404 (O_1404,N_14300,N_14485);
or UO_1405 (O_1405,N_14989,N_14056);
and UO_1406 (O_1406,N_14239,N_14350);
xnor UO_1407 (O_1407,N_14286,N_14387);
nor UO_1408 (O_1408,N_14554,N_14829);
nor UO_1409 (O_1409,N_14755,N_14231);
and UO_1410 (O_1410,N_14741,N_14433);
or UO_1411 (O_1411,N_14157,N_14222);
nand UO_1412 (O_1412,N_14664,N_14405);
and UO_1413 (O_1413,N_14947,N_14278);
nor UO_1414 (O_1414,N_14030,N_14791);
or UO_1415 (O_1415,N_14278,N_14362);
or UO_1416 (O_1416,N_14823,N_14135);
nand UO_1417 (O_1417,N_14149,N_14288);
nor UO_1418 (O_1418,N_14822,N_14871);
nor UO_1419 (O_1419,N_14026,N_14050);
nand UO_1420 (O_1420,N_14823,N_14067);
and UO_1421 (O_1421,N_14827,N_14640);
and UO_1422 (O_1422,N_14396,N_14089);
nand UO_1423 (O_1423,N_14607,N_14357);
nand UO_1424 (O_1424,N_14264,N_14844);
and UO_1425 (O_1425,N_14313,N_14753);
nand UO_1426 (O_1426,N_14294,N_14111);
and UO_1427 (O_1427,N_14222,N_14486);
and UO_1428 (O_1428,N_14376,N_14440);
nand UO_1429 (O_1429,N_14781,N_14269);
or UO_1430 (O_1430,N_14804,N_14041);
or UO_1431 (O_1431,N_14952,N_14398);
or UO_1432 (O_1432,N_14928,N_14158);
and UO_1433 (O_1433,N_14234,N_14053);
nor UO_1434 (O_1434,N_14198,N_14706);
nand UO_1435 (O_1435,N_14062,N_14507);
nand UO_1436 (O_1436,N_14571,N_14215);
and UO_1437 (O_1437,N_14165,N_14041);
and UO_1438 (O_1438,N_14800,N_14834);
nand UO_1439 (O_1439,N_14655,N_14918);
or UO_1440 (O_1440,N_14573,N_14724);
nor UO_1441 (O_1441,N_14903,N_14856);
nor UO_1442 (O_1442,N_14262,N_14349);
nand UO_1443 (O_1443,N_14578,N_14344);
nand UO_1444 (O_1444,N_14235,N_14212);
nor UO_1445 (O_1445,N_14041,N_14906);
nor UO_1446 (O_1446,N_14655,N_14647);
and UO_1447 (O_1447,N_14795,N_14144);
or UO_1448 (O_1448,N_14592,N_14122);
nand UO_1449 (O_1449,N_14446,N_14466);
and UO_1450 (O_1450,N_14082,N_14539);
xnor UO_1451 (O_1451,N_14826,N_14714);
and UO_1452 (O_1452,N_14383,N_14287);
or UO_1453 (O_1453,N_14808,N_14764);
nor UO_1454 (O_1454,N_14544,N_14326);
or UO_1455 (O_1455,N_14337,N_14487);
nand UO_1456 (O_1456,N_14573,N_14526);
nand UO_1457 (O_1457,N_14164,N_14215);
xnor UO_1458 (O_1458,N_14623,N_14810);
nor UO_1459 (O_1459,N_14646,N_14159);
or UO_1460 (O_1460,N_14073,N_14851);
or UO_1461 (O_1461,N_14719,N_14223);
and UO_1462 (O_1462,N_14759,N_14719);
xor UO_1463 (O_1463,N_14225,N_14885);
xnor UO_1464 (O_1464,N_14783,N_14567);
nand UO_1465 (O_1465,N_14622,N_14099);
nand UO_1466 (O_1466,N_14588,N_14916);
and UO_1467 (O_1467,N_14909,N_14356);
or UO_1468 (O_1468,N_14027,N_14005);
nor UO_1469 (O_1469,N_14025,N_14235);
xor UO_1470 (O_1470,N_14628,N_14900);
or UO_1471 (O_1471,N_14921,N_14493);
nand UO_1472 (O_1472,N_14428,N_14001);
nand UO_1473 (O_1473,N_14456,N_14757);
nor UO_1474 (O_1474,N_14147,N_14350);
or UO_1475 (O_1475,N_14054,N_14564);
xnor UO_1476 (O_1476,N_14101,N_14205);
or UO_1477 (O_1477,N_14540,N_14437);
nand UO_1478 (O_1478,N_14420,N_14722);
xnor UO_1479 (O_1479,N_14737,N_14784);
nor UO_1480 (O_1480,N_14178,N_14625);
or UO_1481 (O_1481,N_14111,N_14957);
or UO_1482 (O_1482,N_14418,N_14177);
and UO_1483 (O_1483,N_14205,N_14783);
and UO_1484 (O_1484,N_14631,N_14684);
nand UO_1485 (O_1485,N_14732,N_14052);
nand UO_1486 (O_1486,N_14789,N_14303);
or UO_1487 (O_1487,N_14329,N_14092);
nor UO_1488 (O_1488,N_14651,N_14788);
nand UO_1489 (O_1489,N_14244,N_14840);
or UO_1490 (O_1490,N_14430,N_14240);
xnor UO_1491 (O_1491,N_14785,N_14208);
or UO_1492 (O_1492,N_14879,N_14645);
nor UO_1493 (O_1493,N_14014,N_14224);
or UO_1494 (O_1494,N_14833,N_14945);
or UO_1495 (O_1495,N_14394,N_14164);
and UO_1496 (O_1496,N_14521,N_14738);
nor UO_1497 (O_1497,N_14308,N_14499);
nor UO_1498 (O_1498,N_14871,N_14396);
and UO_1499 (O_1499,N_14583,N_14015);
and UO_1500 (O_1500,N_14806,N_14762);
and UO_1501 (O_1501,N_14819,N_14181);
nor UO_1502 (O_1502,N_14098,N_14236);
and UO_1503 (O_1503,N_14322,N_14285);
xnor UO_1504 (O_1504,N_14269,N_14438);
and UO_1505 (O_1505,N_14897,N_14463);
nand UO_1506 (O_1506,N_14056,N_14249);
and UO_1507 (O_1507,N_14329,N_14385);
nor UO_1508 (O_1508,N_14457,N_14323);
nor UO_1509 (O_1509,N_14137,N_14855);
nand UO_1510 (O_1510,N_14160,N_14892);
nor UO_1511 (O_1511,N_14113,N_14337);
xor UO_1512 (O_1512,N_14220,N_14237);
and UO_1513 (O_1513,N_14279,N_14988);
xor UO_1514 (O_1514,N_14522,N_14510);
nor UO_1515 (O_1515,N_14368,N_14203);
or UO_1516 (O_1516,N_14517,N_14338);
or UO_1517 (O_1517,N_14262,N_14631);
and UO_1518 (O_1518,N_14742,N_14510);
nand UO_1519 (O_1519,N_14937,N_14971);
or UO_1520 (O_1520,N_14473,N_14003);
nand UO_1521 (O_1521,N_14218,N_14844);
nor UO_1522 (O_1522,N_14438,N_14049);
nor UO_1523 (O_1523,N_14517,N_14226);
and UO_1524 (O_1524,N_14348,N_14743);
nand UO_1525 (O_1525,N_14865,N_14914);
and UO_1526 (O_1526,N_14191,N_14501);
and UO_1527 (O_1527,N_14525,N_14897);
nand UO_1528 (O_1528,N_14830,N_14332);
nor UO_1529 (O_1529,N_14828,N_14364);
or UO_1530 (O_1530,N_14432,N_14426);
nand UO_1531 (O_1531,N_14123,N_14085);
or UO_1532 (O_1532,N_14901,N_14553);
nand UO_1533 (O_1533,N_14869,N_14427);
xor UO_1534 (O_1534,N_14846,N_14540);
nor UO_1535 (O_1535,N_14942,N_14543);
and UO_1536 (O_1536,N_14945,N_14348);
and UO_1537 (O_1537,N_14412,N_14426);
and UO_1538 (O_1538,N_14531,N_14738);
and UO_1539 (O_1539,N_14161,N_14317);
nor UO_1540 (O_1540,N_14715,N_14514);
xnor UO_1541 (O_1541,N_14879,N_14178);
xor UO_1542 (O_1542,N_14830,N_14389);
and UO_1543 (O_1543,N_14411,N_14305);
xor UO_1544 (O_1544,N_14148,N_14224);
nor UO_1545 (O_1545,N_14567,N_14587);
and UO_1546 (O_1546,N_14063,N_14816);
nand UO_1547 (O_1547,N_14790,N_14200);
nand UO_1548 (O_1548,N_14183,N_14738);
nor UO_1549 (O_1549,N_14093,N_14408);
xnor UO_1550 (O_1550,N_14699,N_14843);
nand UO_1551 (O_1551,N_14327,N_14123);
nand UO_1552 (O_1552,N_14227,N_14039);
or UO_1553 (O_1553,N_14902,N_14400);
and UO_1554 (O_1554,N_14369,N_14705);
and UO_1555 (O_1555,N_14312,N_14685);
and UO_1556 (O_1556,N_14973,N_14054);
or UO_1557 (O_1557,N_14426,N_14690);
and UO_1558 (O_1558,N_14588,N_14073);
or UO_1559 (O_1559,N_14101,N_14666);
and UO_1560 (O_1560,N_14963,N_14520);
nand UO_1561 (O_1561,N_14716,N_14994);
nand UO_1562 (O_1562,N_14566,N_14446);
nand UO_1563 (O_1563,N_14522,N_14169);
and UO_1564 (O_1564,N_14728,N_14780);
and UO_1565 (O_1565,N_14188,N_14641);
or UO_1566 (O_1566,N_14604,N_14597);
xnor UO_1567 (O_1567,N_14152,N_14691);
nor UO_1568 (O_1568,N_14631,N_14722);
nand UO_1569 (O_1569,N_14543,N_14005);
or UO_1570 (O_1570,N_14624,N_14179);
nand UO_1571 (O_1571,N_14363,N_14554);
nor UO_1572 (O_1572,N_14060,N_14330);
and UO_1573 (O_1573,N_14670,N_14319);
and UO_1574 (O_1574,N_14995,N_14102);
nor UO_1575 (O_1575,N_14375,N_14516);
nor UO_1576 (O_1576,N_14561,N_14352);
and UO_1577 (O_1577,N_14525,N_14349);
or UO_1578 (O_1578,N_14712,N_14579);
nor UO_1579 (O_1579,N_14585,N_14535);
or UO_1580 (O_1580,N_14398,N_14532);
and UO_1581 (O_1581,N_14761,N_14210);
nor UO_1582 (O_1582,N_14448,N_14150);
nor UO_1583 (O_1583,N_14770,N_14191);
nand UO_1584 (O_1584,N_14844,N_14520);
or UO_1585 (O_1585,N_14674,N_14702);
or UO_1586 (O_1586,N_14712,N_14037);
nand UO_1587 (O_1587,N_14276,N_14564);
xor UO_1588 (O_1588,N_14534,N_14970);
and UO_1589 (O_1589,N_14847,N_14289);
and UO_1590 (O_1590,N_14169,N_14317);
and UO_1591 (O_1591,N_14548,N_14584);
nor UO_1592 (O_1592,N_14003,N_14847);
nand UO_1593 (O_1593,N_14291,N_14145);
or UO_1594 (O_1594,N_14015,N_14652);
or UO_1595 (O_1595,N_14679,N_14848);
xor UO_1596 (O_1596,N_14486,N_14562);
and UO_1597 (O_1597,N_14588,N_14887);
and UO_1598 (O_1598,N_14646,N_14927);
nor UO_1599 (O_1599,N_14136,N_14078);
xor UO_1600 (O_1600,N_14015,N_14570);
nand UO_1601 (O_1601,N_14731,N_14126);
nor UO_1602 (O_1602,N_14331,N_14991);
or UO_1603 (O_1603,N_14674,N_14574);
nor UO_1604 (O_1604,N_14545,N_14965);
nand UO_1605 (O_1605,N_14830,N_14529);
or UO_1606 (O_1606,N_14189,N_14031);
or UO_1607 (O_1607,N_14393,N_14328);
nand UO_1608 (O_1608,N_14744,N_14932);
nor UO_1609 (O_1609,N_14139,N_14570);
and UO_1610 (O_1610,N_14487,N_14140);
nand UO_1611 (O_1611,N_14214,N_14734);
or UO_1612 (O_1612,N_14436,N_14478);
or UO_1613 (O_1613,N_14753,N_14467);
nand UO_1614 (O_1614,N_14480,N_14265);
and UO_1615 (O_1615,N_14204,N_14611);
or UO_1616 (O_1616,N_14936,N_14838);
nand UO_1617 (O_1617,N_14344,N_14809);
nor UO_1618 (O_1618,N_14844,N_14243);
nor UO_1619 (O_1619,N_14459,N_14372);
nor UO_1620 (O_1620,N_14293,N_14934);
and UO_1621 (O_1621,N_14117,N_14305);
and UO_1622 (O_1622,N_14916,N_14092);
nand UO_1623 (O_1623,N_14440,N_14380);
or UO_1624 (O_1624,N_14559,N_14084);
nor UO_1625 (O_1625,N_14886,N_14505);
nand UO_1626 (O_1626,N_14699,N_14383);
nor UO_1627 (O_1627,N_14668,N_14363);
and UO_1628 (O_1628,N_14110,N_14415);
nand UO_1629 (O_1629,N_14555,N_14387);
nor UO_1630 (O_1630,N_14921,N_14098);
or UO_1631 (O_1631,N_14431,N_14098);
or UO_1632 (O_1632,N_14835,N_14489);
nand UO_1633 (O_1633,N_14035,N_14223);
or UO_1634 (O_1634,N_14777,N_14555);
nor UO_1635 (O_1635,N_14827,N_14333);
nand UO_1636 (O_1636,N_14792,N_14472);
nor UO_1637 (O_1637,N_14944,N_14201);
or UO_1638 (O_1638,N_14328,N_14543);
or UO_1639 (O_1639,N_14537,N_14477);
and UO_1640 (O_1640,N_14270,N_14014);
nand UO_1641 (O_1641,N_14095,N_14036);
or UO_1642 (O_1642,N_14703,N_14629);
and UO_1643 (O_1643,N_14286,N_14506);
nor UO_1644 (O_1644,N_14411,N_14447);
nand UO_1645 (O_1645,N_14101,N_14048);
nor UO_1646 (O_1646,N_14108,N_14581);
and UO_1647 (O_1647,N_14201,N_14237);
or UO_1648 (O_1648,N_14946,N_14904);
nor UO_1649 (O_1649,N_14677,N_14380);
nand UO_1650 (O_1650,N_14185,N_14695);
or UO_1651 (O_1651,N_14199,N_14184);
and UO_1652 (O_1652,N_14893,N_14157);
nand UO_1653 (O_1653,N_14112,N_14128);
nand UO_1654 (O_1654,N_14330,N_14114);
nand UO_1655 (O_1655,N_14041,N_14244);
nor UO_1656 (O_1656,N_14788,N_14519);
nor UO_1657 (O_1657,N_14177,N_14483);
nand UO_1658 (O_1658,N_14681,N_14739);
and UO_1659 (O_1659,N_14411,N_14674);
and UO_1660 (O_1660,N_14938,N_14859);
nor UO_1661 (O_1661,N_14617,N_14966);
nor UO_1662 (O_1662,N_14388,N_14688);
nor UO_1663 (O_1663,N_14573,N_14360);
or UO_1664 (O_1664,N_14213,N_14034);
nand UO_1665 (O_1665,N_14458,N_14774);
or UO_1666 (O_1666,N_14767,N_14810);
xnor UO_1667 (O_1667,N_14466,N_14705);
or UO_1668 (O_1668,N_14604,N_14246);
or UO_1669 (O_1669,N_14646,N_14393);
or UO_1670 (O_1670,N_14501,N_14001);
xnor UO_1671 (O_1671,N_14574,N_14416);
nand UO_1672 (O_1672,N_14926,N_14911);
or UO_1673 (O_1673,N_14076,N_14201);
and UO_1674 (O_1674,N_14846,N_14255);
nand UO_1675 (O_1675,N_14748,N_14897);
and UO_1676 (O_1676,N_14380,N_14083);
nand UO_1677 (O_1677,N_14549,N_14881);
and UO_1678 (O_1678,N_14095,N_14341);
or UO_1679 (O_1679,N_14006,N_14459);
nand UO_1680 (O_1680,N_14074,N_14253);
xnor UO_1681 (O_1681,N_14419,N_14148);
nor UO_1682 (O_1682,N_14900,N_14571);
or UO_1683 (O_1683,N_14438,N_14040);
and UO_1684 (O_1684,N_14755,N_14698);
nand UO_1685 (O_1685,N_14513,N_14850);
and UO_1686 (O_1686,N_14449,N_14081);
nand UO_1687 (O_1687,N_14643,N_14167);
nor UO_1688 (O_1688,N_14096,N_14742);
nor UO_1689 (O_1689,N_14748,N_14571);
nor UO_1690 (O_1690,N_14684,N_14587);
and UO_1691 (O_1691,N_14639,N_14499);
nor UO_1692 (O_1692,N_14167,N_14793);
and UO_1693 (O_1693,N_14392,N_14604);
or UO_1694 (O_1694,N_14791,N_14780);
and UO_1695 (O_1695,N_14017,N_14191);
nor UO_1696 (O_1696,N_14506,N_14643);
nand UO_1697 (O_1697,N_14058,N_14015);
or UO_1698 (O_1698,N_14937,N_14298);
nor UO_1699 (O_1699,N_14444,N_14477);
and UO_1700 (O_1700,N_14453,N_14355);
xor UO_1701 (O_1701,N_14388,N_14470);
nor UO_1702 (O_1702,N_14470,N_14624);
nand UO_1703 (O_1703,N_14748,N_14523);
nand UO_1704 (O_1704,N_14518,N_14281);
nand UO_1705 (O_1705,N_14729,N_14062);
xor UO_1706 (O_1706,N_14512,N_14972);
nand UO_1707 (O_1707,N_14412,N_14482);
nor UO_1708 (O_1708,N_14959,N_14826);
nand UO_1709 (O_1709,N_14261,N_14577);
xor UO_1710 (O_1710,N_14013,N_14627);
nand UO_1711 (O_1711,N_14613,N_14003);
nand UO_1712 (O_1712,N_14807,N_14108);
nor UO_1713 (O_1713,N_14465,N_14037);
or UO_1714 (O_1714,N_14421,N_14563);
and UO_1715 (O_1715,N_14992,N_14872);
nand UO_1716 (O_1716,N_14193,N_14771);
nand UO_1717 (O_1717,N_14157,N_14568);
and UO_1718 (O_1718,N_14139,N_14694);
nor UO_1719 (O_1719,N_14337,N_14273);
or UO_1720 (O_1720,N_14283,N_14970);
nand UO_1721 (O_1721,N_14573,N_14933);
nand UO_1722 (O_1722,N_14468,N_14950);
and UO_1723 (O_1723,N_14815,N_14408);
nand UO_1724 (O_1724,N_14947,N_14964);
nor UO_1725 (O_1725,N_14231,N_14310);
and UO_1726 (O_1726,N_14594,N_14642);
nand UO_1727 (O_1727,N_14591,N_14666);
xor UO_1728 (O_1728,N_14623,N_14943);
or UO_1729 (O_1729,N_14426,N_14867);
nand UO_1730 (O_1730,N_14649,N_14136);
and UO_1731 (O_1731,N_14798,N_14806);
xor UO_1732 (O_1732,N_14738,N_14501);
nand UO_1733 (O_1733,N_14603,N_14262);
xnor UO_1734 (O_1734,N_14732,N_14351);
nand UO_1735 (O_1735,N_14098,N_14643);
nand UO_1736 (O_1736,N_14213,N_14076);
and UO_1737 (O_1737,N_14934,N_14688);
or UO_1738 (O_1738,N_14835,N_14915);
nand UO_1739 (O_1739,N_14753,N_14283);
and UO_1740 (O_1740,N_14275,N_14237);
xnor UO_1741 (O_1741,N_14720,N_14426);
nor UO_1742 (O_1742,N_14090,N_14628);
and UO_1743 (O_1743,N_14915,N_14819);
nand UO_1744 (O_1744,N_14921,N_14479);
nand UO_1745 (O_1745,N_14590,N_14629);
nand UO_1746 (O_1746,N_14776,N_14244);
nand UO_1747 (O_1747,N_14062,N_14520);
nor UO_1748 (O_1748,N_14007,N_14907);
nor UO_1749 (O_1749,N_14845,N_14935);
nand UO_1750 (O_1750,N_14439,N_14907);
or UO_1751 (O_1751,N_14748,N_14500);
and UO_1752 (O_1752,N_14606,N_14328);
nand UO_1753 (O_1753,N_14764,N_14613);
nor UO_1754 (O_1754,N_14591,N_14099);
nand UO_1755 (O_1755,N_14442,N_14781);
or UO_1756 (O_1756,N_14531,N_14526);
or UO_1757 (O_1757,N_14703,N_14470);
and UO_1758 (O_1758,N_14236,N_14229);
and UO_1759 (O_1759,N_14705,N_14751);
xor UO_1760 (O_1760,N_14377,N_14130);
nand UO_1761 (O_1761,N_14725,N_14151);
or UO_1762 (O_1762,N_14465,N_14106);
and UO_1763 (O_1763,N_14290,N_14220);
nor UO_1764 (O_1764,N_14827,N_14877);
and UO_1765 (O_1765,N_14791,N_14519);
xnor UO_1766 (O_1766,N_14741,N_14539);
nor UO_1767 (O_1767,N_14666,N_14810);
nand UO_1768 (O_1768,N_14687,N_14943);
or UO_1769 (O_1769,N_14986,N_14987);
nand UO_1770 (O_1770,N_14197,N_14726);
xnor UO_1771 (O_1771,N_14433,N_14076);
or UO_1772 (O_1772,N_14404,N_14761);
nor UO_1773 (O_1773,N_14598,N_14263);
nor UO_1774 (O_1774,N_14652,N_14636);
or UO_1775 (O_1775,N_14197,N_14317);
nor UO_1776 (O_1776,N_14587,N_14657);
nor UO_1777 (O_1777,N_14585,N_14528);
and UO_1778 (O_1778,N_14835,N_14329);
nand UO_1779 (O_1779,N_14037,N_14827);
nand UO_1780 (O_1780,N_14181,N_14663);
and UO_1781 (O_1781,N_14221,N_14140);
or UO_1782 (O_1782,N_14892,N_14292);
and UO_1783 (O_1783,N_14822,N_14513);
nor UO_1784 (O_1784,N_14169,N_14999);
nand UO_1785 (O_1785,N_14490,N_14631);
nand UO_1786 (O_1786,N_14519,N_14352);
and UO_1787 (O_1787,N_14441,N_14570);
nand UO_1788 (O_1788,N_14636,N_14639);
nand UO_1789 (O_1789,N_14454,N_14712);
xnor UO_1790 (O_1790,N_14209,N_14670);
and UO_1791 (O_1791,N_14575,N_14433);
and UO_1792 (O_1792,N_14170,N_14411);
xnor UO_1793 (O_1793,N_14167,N_14135);
and UO_1794 (O_1794,N_14183,N_14211);
and UO_1795 (O_1795,N_14716,N_14695);
nor UO_1796 (O_1796,N_14616,N_14589);
xnor UO_1797 (O_1797,N_14615,N_14192);
or UO_1798 (O_1798,N_14591,N_14798);
and UO_1799 (O_1799,N_14917,N_14170);
nand UO_1800 (O_1800,N_14816,N_14460);
nand UO_1801 (O_1801,N_14420,N_14779);
nor UO_1802 (O_1802,N_14814,N_14444);
nand UO_1803 (O_1803,N_14690,N_14222);
and UO_1804 (O_1804,N_14265,N_14481);
xnor UO_1805 (O_1805,N_14996,N_14190);
nor UO_1806 (O_1806,N_14085,N_14541);
and UO_1807 (O_1807,N_14250,N_14029);
or UO_1808 (O_1808,N_14360,N_14983);
and UO_1809 (O_1809,N_14665,N_14096);
or UO_1810 (O_1810,N_14552,N_14405);
or UO_1811 (O_1811,N_14519,N_14084);
nor UO_1812 (O_1812,N_14995,N_14293);
nand UO_1813 (O_1813,N_14760,N_14643);
nor UO_1814 (O_1814,N_14330,N_14367);
nor UO_1815 (O_1815,N_14127,N_14636);
xor UO_1816 (O_1816,N_14057,N_14460);
or UO_1817 (O_1817,N_14201,N_14616);
nand UO_1818 (O_1818,N_14612,N_14875);
nor UO_1819 (O_1819,N_14359,N_14876);
or UO_1820 (O_1820,N_14149,N_14061);
nand UO_1821 (O_1821,N_14392,N_14436);
nand UO_1822 (O_1822,N_14938,N_14389);
or UO_1823 (O_1823,N_14363,N_14743);
nand UO_1824 (O_1824,N_14830,N_14305);
and UO_1825 (O_1825,N_14578,N_14694);
nand UO_1826 (O_1826,N_14506,N_14143);
and UO_1827 (O_1827,N_14763,N_14471);
or UO_1828 (O_1828,N_14689,N_14275);
nor UO_1829 (O_1829,N_14867,N_14792);
nand UO_1830 (O_1830,N_14541,N_14429);
or UO_1831 (O_1831,N_14976,N_14073);
or UO_1832 (O_1832,N_14935,N_14077);
nand UO_1833 (O_1833,N_14262,N_14322);
and UO_1834 (O_1834,N_14951,N_14495);
xnor UO_1835 (O_1835,N_14083,N_14386);
and UO_1836 (O_1836,N_14681,N_14924);
and UO_1837 (O_1837,N_14318,N_14875);
or UO_1838 (O_1838,N_14933,N_14330);
or UO_1839 (O_1839,N_14645,N_14231);
nand UO_1840 (O_1840,N_14797,N_14765);
and UO_1841 (O_1841,N_14655,N_14401);
nand UO_1842 (O_1842,N_14755,N_14101);
or UO_1843 (O_1843,N_14040,N_14819);
or UO_1844 (O_1844,N_14476,N_14797);
nor UO_1845 (O_1845,N_14826,N_14177);
nor UO_1846 (O_1846,N_14145,N_14992);
or UO_1847 (O_1847,N_14671,N_14837);
or UO_1848 (O_1848,N_14450,N_14963);
and UO_1849 (O_1849,N_14586,N_14527);
and UO_1850 (O_1850,N_14751,N_14793);
or UO_1851 (O_1851,N_14425,N_14415);
nor UO_1852 (O_1852,N_14553,N_14037);
nand UO_1853 (O_1853,N_14643,N_14559);
xor UO_1854 (O_1854,N_14906,N_14211);
xnor UO_1855 (O_1855,N_14166,N_14088);
and UO_1856 (O_1856,N_14004,N_14199);
or UO_1857 (O_1857,N_14168,N_14172);
nand UO_1858 (O_1858,N_14038,N_14982);
and UO_1859 (O_1859,N_14905,N_14192);
or UO_1860 (O_1860,N_14748,N_14608);
and UO_1861 (O_1861,N_14805,N_14999);
nand UO_1862 (O_1862,N_14677,N_14579);
nor UO_1863 (O_1863,N_14381,N_14052);
nand UO_1864 (O_1864,N_14490,N_14481);
nor UO_1865 (O_1865,N_14015,N_14540);
xor UO_1866 (O_1866,N_14121,N_14550);
nand UO_1867 (O_1867,N_14095,N_14013);
nand UO_1868 (O_1868,N_14401,N_14875);
or UO_1869 (O_1869,N_14467,N_14638);
nor UO_1870 (O_1870,N_14201,N_14175);
nor UO_1871 (O_1871,N_14893,N_14817);
nand UO_1872 (O_1872,N_14291,N_14614);
nor UO_1873 (O_1873,N_14589,N_14451);
nand UO_1874 (O_1874,N_14168,N_14988);
nor UO_1875 (O_1875,N_14620,N_14892);
nor UO_1876 (O_1876,N_14663,N_14571);
nand UO_1877 (O_1877,N_14649,N_14759);
or UO_1878 (O_1878,N_14157,N_14178);
or UO_1879 (O_1879,N_14958,N_14968);
nor UO_1880 (O_1880,N_14213,N_14891);
nand UO_1881 (O_1881,N_14771,N_14578);
and UO_1882 (O_1882,N_14673,N_14566);
nand UO_1883 (O_1883,N_14591,N_14901);
or UO_1884 (O_1884,N_14509,N_14799);
and UO_1885 (O_1885,N_14737,N_14038);
and UO_1886 (O_1886,N_14051,N_14425);
nor UO_1887 (O_1887,N_14433,N_14303);
xnor UO_1888 (O_1888,N_14157,N_14040);
nor UO_1889 (O_1889,N_14462,N_14522);
nand UO_1890 (O_1890,N_14072,N_14496);
nor UO_1891 (O_1891,N_14594,N_14427);
and UO_1892 (O_1892,N_14341,N_14785);
and UO_1893 (O_1893,N_14582,N_14927);
and UO_1894 (O_1894,N_14040,N_14146);
xor UO_1895 (O_1895,N_14721,N_14480);
nand UO_1896 (O_1896,N_14203,N_14154);
nand UO_1897 (O_1897,N_14400,N_14690);
nand UO_1898 (O_1898,N_14027,N_14950);
nand UO_1899 (O_1899,N_14041,N_14825);
and UO_1900 (O_1900,N_14382,N_14531);
nand UO_1901 (O_1901,N_14209,N_14230);
nand UO_1902 (O_1902,N_14477,N_14135);
nor UO_1903 (O_1903,N_14727,N_14407);
and UO_1904 (O_1904,N_14506,N_14541);
xnor UO_1905 (O_1905,N_14055,N_14453);
xnor UO_1906 (O_1906,N_14639,N_14934);
nor UO_1907 (O_1907,N_14704,N_14081);
or UO_1908 (O_1908,N_14398,N_14242);
and UO_1909 (O_1909,N_14862,N_14471);
or UO_1910 (O_1910,N_14281,N_14680);
nor UO_1911 (O_1911,N_14988,N_14761);
nor UO_1912 (O_1912,N_14429,N_14964);
nor UO_1913 (O_1913,N_14273,N_14830);
nor UO_1914 (O_1914,N_14898,N_14273);
and UO_1915 (O_1915,N_14947,N_14283);
nand UO_1916 (O_1916,N_14281,N_14718);
nor UO_1917 (O_1917,N_14121,N_14205);
or UO_1918 (O_1918,N_14752,N_14633);
xnor UO_1919 (O_1919,N_14598,N_14585);
nand UO_1920 (O_1920,N_14127,N_14501);
nand UO_1921 (O_1921,N_14297,N_14548);
nor UO_1922 (O_1922,N_14550,N_14557);
or UO_1923 (O_1923,N_14440,N_14563);
nand UO_1924 (O_1924,N_14211,N_14683);
nand UO_1925 (O_1925,N_14557,N_14170);
and UO_1926 (O_1926,N_14477,N_14337);
or UO_1927 (O_1927,N_14544,N_14895);
and UO_1928 (O_1928,N_14311,N_14770);
and UO_1929 (O_1929,N_14572,N_14737);
and UO_1930 (O_1930,N_14090,N_14174);
or UO_1931 (O_1931,N_14998,N_14492);
or UO_1932 (O_1932,N_14399,N_14023);
nand UO_1933 (O_1933,N_14202,N_14187);
or UO_1934 (O_1934,N_14894,N_14725);
nor UO_1935 (O_1935,N_14892,N_14987);
nor UO_1936 (O_1936,N_14902,N_14584);
or UO_1937 (O_1937,N_14295,N_14132);
and UO_1938 (O_1938,N_14049,N_14239);
nand UO_1939 (O_1939,N_14362,N_14126);
and UO_1940 (O_1940,N_14134,N_14207);
nand UO_1941 (O_1941,N_14018,N_14436);
and UO_1942 (O_1942,N_14160,N_14431);
or UO_1943 (O_1943,N_14083,N_14749);
nand UO_1944 (O_1944,N_14198,N_14813);
and UO_1945 (O_1945,N_14618,N_14176);
xor UO_1946 (O_1946,N_14133,N_14394);
and UO_1947 (O_1947,N_14710,N_14518);
and UO_1948 (O_1948,N_14510,N_14963);
nor UO_1949 (O_1949,N_14275,N_14378);
and UO_1950 (O_1950,N_14578,N_14210);
and UO_1951 (O_1951,N_14642,N_14610);
and UO_1952 (O_1952,N_14739,N_14731);
nor UO_1953 (O_1953,N_14691,N_14079);
and UO_1954 (O_1954,N_14864,N_14594);
or UO_1955 (O_1955,N_14533,N_14045);
or UO_1956 (O_1956,N_14076,N_14886);
and UO_1957 (O_1957,N_14488,N_14075);
or UO_1958 (O_1958,N_14260,N_14436);
nand UO_1959 (O_1959,N_14363,N_14705);
and UO_1960 (O_1960,N_14878,N_14216);
and UO_1961 (O_1961,N_14234,N_14452);
nor UO_1962 (O_1962,N_14795,N_14812);
and UO_1963 (O_1963,N_14955,N_14488);
nor UO_1964 (O_1964,N_14172,N_14438);
nand UO_1965 (O_1965,N_14076,N_14288);
nor UO_1966 (O_1966,N_14895,N_14107);
nor UO_1967 (O_1967,N_14927,N_14433);
or UO_1968 (O_1968,N_14443,N_14741);
nor UO_1969 (O_1969,N_14392,N_14535);
and UO_1970 (O_1970,N_14596,N_14648);
or UO_1971 (O_1971,N_14432,N_14854);
nor UO_1972 (O_1972,N_14047,N_14046);
and UO_1973 (O_1973,N_14233,N_14523);
and UO_1974 (O_1974,N_14633,N_14442);
nor UO_1975 (O_1975,N_14544,N_14381);
nor UO_1976 (O_1976,N_14265,N_14146);
nor UO_1977 (O_1977,N_14250,N_14576);
or UO_1978 (O_1978,N_14526,N_14746);
nor UO_1979 (O_1979,N_14923,N_14663);
and UO_1980 (O_1980,N_14729,N_14589);
xor UO_1981 (O_1981,N_14935,N_14411);
and UO_1982 (O_1982,N_14687,N_14270);
nand UO_1983 (O_1983,N_14254,N_14890);
or UO_1984 (O_1984,N_14247,N_14901);
and UO_1985 (O_1985,N_14497,N_14164);
nor UO_1986 (O_1986,N_14026,N_14494);
nand UO_1987 (O_1987,N_14438,N_14698);
or UO_1988 (O_1988,N_14215,N_14680);
or UO_1989 (O_1989,N_14914,N_14871);
and UO_1990 (O_1990,N_14203,N_14108);
nand UO_1991 (O_1991,N_14148,N_14483);
xor UO_1992 (O_1992,N_14867,N_14811);
nor UO_1993 (O_1993,N_14896,N_14140);
or UO_1994 (O_1994,N_14894,N_14223);
and UO_1995 (O_1995,N_14927,N_14343);
nor UO_1996 (O_1996,N_14923,N_14344);
nor UO_1997 (O_1997,N_14550,N_14735);
xor UO_1998 (O_1998,N_14963,N_14211);
or UO_1999 (O_1999,N_14789,N_14338);
endmodule