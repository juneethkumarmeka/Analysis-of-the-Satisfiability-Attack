module basic_5000_50000_5000_20_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
and U0 (N_0,In_4903,In_2742);
or U1 (N_1,In_3140,In_4956);
or U2 (N_2,In_4871,In_3184);
xnor U3 (N_3,In_2112,In_1801);
nand U4 (N_4,In_1406,In_3064);
nand U5 (N_5,In_3676,In_3263);
nor U6 (N_6,In_4378,In_1374);
nand U7 (N_7,In_3728,In_1389);
xor U8 (N_8,In_4425,In_4165);
nand U9 (N_9,In_1394,In_4277);
nor U10 (N_10,In_4401,In_3298);
or U11 (N_11,In_1852,In_1850);
xnor U12 (N_12,In_4839,In_1268);
and U13 (N_13,In_4914,In_2220);
xor U14 (N_14,In_4962,In_4854);
xnor U15 (N_15,In_2647,In_2033);
or U16 (N_16,In_1387,In_4122);
nand U17 (N_17,In_2453,In_1944);
xnor U18 (N_18,In_3190,In_4537);
xor U19 (N_19,In_2456,In_1802);
or U20 (N_20,In_1405,In_4883);
and U21 (N_21,In_3264,In_879);
and U22 (N_22,In_2982,In_3032);
nand U23 (N_23,In_1205,In_2744);
xnor U24 (N_24,In_1708,In_4028);
nand U25 (N_25,In_2165,In_1202);
nor U26 (N_26,In_3246,In_3565);
nand U27 (N_27,In_4761,In_3227);
nand U28 (N_28,In_666,In_3035);
xor U29 (N_29,In_1099,In_4197);
xnor U30 (N_30,In_4658,In_1867);
and U31 (N_31,In_4265,In_1919);
nand U32 (N_32,In_3285,In_3522);
nor U33 (N_33,In_3417,In_2531);
and U34 (N_34,In_2078,In_3974);
or U35 (N_35,In_4693,In_2351);
nor U36 (N_36,In_3614,In_2440);
and U37 (N_37,In_4105,In_3960);
and U38 (N_38,In_1547,In_1145);
nand U39 (N_39,In_244,In_1688);
and U40 (N_40,In_3454,In_3476);
nand U41 (N_41,In_76,In_1050);
and U42 (N_42,In_2523,In_2676);
and U43 (N_43,In_947,In_2208);
or U44 (N_44,In_3238,In_4167);
nand U45 (N_45,In_4697,In_2297);
xor U46 (N_46,In_4734,In_1669);
nand U47 (N_47,In_1682,In_4846);
nor U48 (N_48,In_119,In_4725);
nand U49 (N_49,In_882,In_2395);
and U50 (N_50,In_3374,In_1732);
and U51 (N_51,In_691,In_1165);
nor U52 (N_52,In_2049,In_2569);
xor U53 (N_53,In_3570,In_1827);
nor U54 (N_54,In_821,In_728);
and U55 (N_55,In_3529,In_3203);
xnor U56 (N_56,In_3860,In_1316);
nand U57 (N_57,In_2031,In_3633);
nand U58 (N_58,In_1844,In_1700);
nor U59 (N_59,In_4504,In_470);
and U60 (N_60,In_3211,In_3596);
nand U61 (N_61,In_1879,In_346);
nand U62 (N_62,In_1560,In_38);
xnor U63 (N_63,In_3581,In_4580);
xor U64 (N_64,In_1528,In_206);
nand U65 (N_65,In_1989,In_4745);
xnor U66 (N_66,In_1735,In_779);
and U67 (N_67,In_543,In_4226);
nand U68 (N_68,In_1445,In_521);
xnor U69 (N_69,In_4662,In_2872);
nor U70 (N_70,In_405,In_2232);
and U71 (N_71,In_4957,In_515);
xor U72 (N_72,In_2250,In_437);
and U73 (N_73,In_3471,In_3413);
or U74 (N_74,In_435,In_2589);
xnor U75 (N_75,In_1450,In_429);
xnor U76 (N_76,In_4615,In_4894);
or U77 (N_77,In_4251,In_4519);
nand U78 (N_78,In_1585,In_4332);
nor U79 (N_79,In_2741,In_3718);
or U80 (N_80,In_355,In_1131);
or U81 (N_81,In_4155,In_1550);
or U82 (N_82,In_1933,In_4361);
nor U83 (N_83,In_1414,In_4272);
nor U84 (N_84,In_4009,In_2255);
and U85 (N_85,In_3116,In_3863);
nand U86 (N_86,In_3143,In_4482);
nand U87 (N_87,In_2431,In_1460);
and U88 (N_88,In_3661,In_298);
nand U89 (N_89,In_4000,In_4427);
and U90 (N_90,In_3253,In_4083);
nand U91 (N_91,In_563,In_2796);
xor U92 (N_92,In_1102,In_3490);
or U93 (N_93,In_1346,In_265);
nor U94 (N_94,In_2190,In_3590);
or U95 (N_95,In_2672,In_1804);
nor U96 (N_96,In_2080,In_1592);
nor U97 (N_97,In_4162,In_3110);
nand U98 (N_98,In_4412,In_3392);
xor U99 (N_99,In_2187,In_2211);
xnor U100 (N_100,In_2681,In_1244);
and U101 (N_101,In_4780,In_1035);
nor U102 (N_102,In_2148,In_1261);
nand U103 (N_103,In_2203,In_3368);
or U104 (N_104,In_3346,In_1957);
or U105 (N_105,In_987,In_1794);
nand U106 (N_106,In_3220,In_3616);
xor U107 (N_107,In_4326,In_3435);
nor U108 (N_108,In_3158,In_1539);
or U109 (N_109,In_1631,In_1027);
xnor U110 (N_110,In_1437,In_1982);
or U111 (N_111,In_1410,In_96);
or U112 (N_112,In_3147,In_2519);
xnor U113 (N_113,In_2246,In_1074);
or U114 (N_114,In_4203,In_3039);
xnor U115 (N_115,In_4334,In_782);
xor U116 (N_116,In_796,In_712);
and U117 (N_117,In_502,In_4360);
xnor U118 (N_118,In_2280,In_2830);
xnor U119 (N_119,In_3390,In_3835);
xnor U120 (N_120,In_140,In_1606);
nor U121 (N_121,In_4639,In_4475);
xor U122 (N_122,In_2850,In_1505);
xor U123 (N_123,In_4,In_4984);
nand U124 (N_124,In_2882,In_2684);
nor U125 (N_125,In_1129,In_2483);
nand U126 (N_126,In_2310,In_3963);
xnor U127 (N_127,In_4436,In_4570);
and U128 (N_128,In_3630,In_406);
nor U129 (N_129,In_272,In_2918);
nand U130 (N_130,In_3037,In_2240);
xor U131 (N_131,In_2314,In_1004);
xnor U132 (N_132,In_3175,In_2450);
and U133 (N_133,In_1239,In_3946);
nand U134 (N_134,In_4999,In_3660);
or U135 (N_135,In_212,In_2798);
nor U136 (N_136,In_3913,In_2394);
nor U137 (N_137,In_1355,In_3840);
or U138 (N_138,In_1251,In_45);
and U139 (N_139,In_3329,In_2114);
xor U140 (N_140,In_234,In_952);
xnor U141 (N_141,In_104,In_575);
xnor U142 (N_142,In_2392,In_117);
nand U143 (N_143,In_304,In_3900);
or U144 (N_144,In_2467,In_2898);
and U145 (N_145,In_3875,In_2139);
or U146 (N_146,In_1079,In_1218);
nor U147 (N_147,In_3341,In_2058);
or U148 (N_148,In_3470,In_3343);
nor U149 (N_149,In_67,In_4524);
xnor U150 (N_150,In_3272,In_756);
nand U151 (N_151,In_3081,In_4297);
nand U152 (N_152,In_3154,In_2306);
nand U153 (N_153,In_3256,In_4595);
xnor U154 (N_154,In_3700,In_1098);
or U155 (N_155,In_511,In_2169);
and U156 (N_156,In_404,In_3168);
xor U157 (N_157,In_1266,In_1213);
and U158 (N_158,In_1292,In_4836);
or U159 (N_159,In_2299,In_711);
and U160 (N_160,In_939,In_3122);
or U161 (N_161,In_1956,In_4769);
xor U162 (N_162,In_548,In_282);
or U163 (N_163,In_602,In_936);
nor U164 (N_164,In_2085,In_601);
and U165 (N_165,In_4875,In_3832);
and U166 (N_166,In_428,In_3772);
and U167 (N_167,In_1705,In_1275);
and U168 (N_168,In_2891,In_3194);
and U169 (N_169,In_914,In_3048);
or U170 (N_170,In_2161,In_4055);
or U171 (N_171,In_1019,In_2752);
xnor U172 (N_172,In_1051,In_63);
nor U173 (N_173,In_4454,In_695);
xor U174 (N_174,In_1876,In_478);
and U175 (N_175,In_3381,In_3536);
xor U176 (N_176,In_4908,In_1716);
or U177 (N_177,In_4910,In_2677);
or U178 (N_178,In_1635,In_559);
and U179 (N_179,In_2097,In_2803);
nor U180 (N_180,In_2474,In_1734);
or U181 (N_181,In_3248,In_3905);
xnor U182 (N_182,In_4195,In_341);
or U183 (N_183,In_447,In_2194);
nand U184 (N_184,In_1461,In_4258);
and U185 (N_185,In_1568,In_3895);
and U186 (N_186,In_4629,In_2309);
or U187 (N_187,In_2035,In_2151);
or U188 (N_188,In_121,In_1122);
or U189 (N_189,In_2438,In_3199);
nand U190 (N_190,In_3911,In_4208);
or U191 (N_191,In_3903,In_2267);
or U192 (N_192,In_794,In_4045);
nand U193 (N_193,In_1358,In_3856);
nand U194 (N_194,In_710,In_2973);
nand U195 (N_195,In_1687,In_2880);
nand U196 (N_196,In_4492,In_3228);
and U197 (N_197,In_2350,In_860);
xor U198 (N_198,In_685,In_2132);
nor U199 (N_199,In_824,In_3178);
nor U200 (N_200,In_1111,In_269);
nor U201 (N_201,In_1357,In_2380);
and U202 (N_202,In_3339,In_2059);
xor U203 (N_203,In_2908,In_3153);
nor U204 (N_204,In_1337,In_2956);
xor U205 (N_205,In_1083,In_913);
nor U206 (N_206,In_3928,In_3210);
and U207 (N_207,In_761,In_1141);
nand U208 (N_208,In_3924,In_644);
xor U209 (N_209,In_815,In_825);
xor U210 (N_210,In_4490,In_2773);
xnor U211 (N_211,In_1230,In_3984);
or U212 (N_212,In_560,In_702);
nand U213 (N_213,In_2659,In_3366);
nand U214 (N_214,In_1820,In_1639);
nand U215 (N_215,In_3890,In_1272);
xnor U216 (N_216,In_1578,In_1863);
xor U217 (N_217,In_4461,In_4359);
or U218 (N_218,In_3371,In_1249);
or U219 (N_219,In_1726,In_2378);
nor U220 (N_220,In_1649,In_4606);
or U221 (N_221,In_1717,In_4784);
and U222 (N_222,In_1604,In_1000);
nor U223 (N_223,In_2176,In_1656);
xnor U224 (N_224,In_596,In_1685);
nor U225 (N_225,In_3815,In_1484);
nor U226 (N_226,In_3337,In_1676);
or U227 (N_227,In_4551,In_313);
nor U228 (N_228,In_4338,In_3767);
or U229 (N_229,In_1022,In_1628);
xnor U230 (N_230,In_3102,In_394);
nor U231 (N_231,In_1113,In_4937);
xor U232 (N_232,In_2279,In_3555);
xor U233 (N_233,In_3687,In_1285);
and U234 (N_234,In_3694,In_4145);
and U235 (N_235,In_725,In_3019);
or U236 (N_236,In_1882,In_3968);
or U237 (N_237,In_1215,In_102);
and U238 (N_238,In_3094,In_2144);
nor U239 (N_239,In_4317,In_2482);
xor U240 (N_240,In_3222,In_4523);
nand U241 (N_241,In_2814,In_3891);
nand U242 (N_242,In_3411,In_1817);
xor U243 (N_243,In_643,In_3934);
xor U244 (N_244,In_3010,In_4563);
nor U245 (N_245,In_2832,In_1830);
and U246 (N_246,In_1293,In_2191);
and U247 (N_247,In_4856,In_2278);
xor U248 (N_248,In_2641,In_866);
and U249 (N_249,In_4939,In_4421);
or U250 (N_250,In_1730,In_2466);
nand U251 (N_251,In_4952,In_4276);
or U252 (N_252,In_4770,In_1784);
and U253 (N_253,In_332,In_4690);
nand U254 (N_254,In_5,In_901);
and U255 (N_255,In_2905,In_3977);
and U256 (N_256,In_906,In_673);
or U257 (N_257,In_4178,In_2865);
or U258 (N_258,In_4295,In_2695);
or U259 (N_259,In_1370,In_4822);
or U260 (N_260,In_2414,In_2625);
nand U261 (N_261,In_4684,In_115);
nor U262 (N_262,In_1853,In_1482);
xor U263 (N_263,In_979,In_86);
or U264 (N_264,In_4241,In_3384);
nand U265 (N_265,In_3512,In_2717);
nand U266 (N_266,In_3301,In_2597);
and U267 (N_267,In_3050,In_3439);
or U268 (N_268,In_1227,In_1323);
nand U269 (N_269,In_1872,In_2719);
nand U270 (N_270,In_3882,In_2781);
xnor U271 (N_271,In_1948,In_3046);
xor U272 (N_272,In_1938,In_4816);
nand U273 (N_273,In_335,In_3123);
xnor U274 (N_274,In_2789,In_4656);
nor U275 (N_275,In_4699,In_3990);
nor U276 (N_276,In_607,In_327);
nand U277 (N_277,In_479,In_186);
and U278 (N_278,In_4592,In_1194);
or U279 (N_279,In_4456,In_142);
or U280 (N_280,In_780,In_2367);
nor U281 (N_281,In_4309,In_3855);
nand U282 (N_282,In_4131,In_742);
or U283 (N_283,In_382,In_4247);
or U284 (N_284,In_2439,In_2551);
and U285 (N_285,In_3732,In_2501);
and U286 (N_286,In_258,In_2291);
xor U287 (N_287,In_3598,In_708);
nand U288 (N_288,In_4054,In_3736);
nor U289 (N_289,In_3436,In_2166);
nor U290 (N_290,In_4588,In_3808);
nor U291 (N_291,In_4351,In_3502);
and U292 (N_292,In_1760,In_425);
nand U293 (N_293,In_3080,In_4527);
and U294 (N_294,In_2349,In_2635);
and U295 (N_295,In_3982,In_2019);
nand U296 (N_296,In_929,In_3790);
and U297 (N_297,In_1930,In_2428);
nand U298 (N_298,In_4892,In_3745);
or U299 (N_299,In_854,In_2312);
or U300 (N_300,In_1348,In_30);
xnor U301 (N_301,In_758,In_295);
xnor U302 (N_302,In_4749,In_3557);
nand U303 (N_303,In_1479,In_3171);
or U304 (N_304,In_1121,In_4802);
nand U305 (N_305,In_1080,In_2664);
xor U306 (N_306,In_2996,In_2769);
and U307 (N_307,In_3567,In_4765);
nor U308 (N_308,In_1819,In_1335);
or U309 (N_309,In_453,In_1049);
nand U310 (N_310,In_2831,In_2617);
and U311 (N_311,In_2041,In_3219);
nor U312 (N_312,In_3308,In_2845);
or U313 (N_313,In_1363,In_1373);
xor U314 (N_314,In_1318,In_2917);
and U315 (N_315,In_1652,In_2821);
nand U316 (N_316,In_1743,In_769);
and U317 (N_317,In_3132,In_1671);
or U318 (N_318,In_4949,In_3358);
or U319 (N_319,In_1514,In_627);
and U320 (N_320,In_2671,In_4261);
and U321 (N_321,In_25,In_2648);
xor U322 (N_322,In_3018,In_4535);
and U323 (N_323,In_1220,In_152);
xnor U324 (N_324,In_1324,In_2331);
xnor U325 (N_325,In_2311,In_3568);
nor U326 (N_326,In_4188,In_1090);
and U327 (N_327,In_413,In_3317);
xnor U328 (N_328,In_4845,In_1477);
or U329 (N_329,In_65,In_3867);
nand U330 (N_330,In_4096,In_922);
and U331 (N_331,In_4763,In_3088);
or U332 (N_332,In_2273,In_716);
or U333 (N_333,In_4095,In_3440);
nand U334 (N_334,In_4236,In_4798);
nand U335 (N_335,In_2300,In_1845);
xnor U336 (N_336,In_2774,In_3837);
or U337 (N_337,In_3484,In_2621);
nor U338 (N_338,In_1965,In_1892);
or U339 (N_339,In_3364,In_3532);
or U340 (N_340,In_320,In_783);
nand U341 (N_341,In_4479,In_2733);
and U342 (N_342,In_3193,In_3103);
nand U343 (N_343,In_944,In_3268);
xnor U344 (N_344,In_3187,In_4429);
nand U345 (N_345,In_583,In_4548);
and U346 (N_346,In_615,In_2063);
xnor U347 (N_347,In_3877,In_3);
and U348 (N_348,In_160,In_3709);
nand U349 (N_349,In_4638,In_565);
or U350 (N_350,In_463,In_4449);
xnor U351 (N_351,In_3431,In_2270);
or U352 (N_352,In_998,In_4774);
nand U353 (N_353,In_4224,In_4652);
xor U354 (N_354,In_1707,In_2925);
nor U355 (N_355,In_4576,In_2330);
nor U356 (N_356,In_2053,In_226);
nand U357 (N_357,In_2700,In_4969);
and U358 (N_358,In_81,In_4586);
or U359 (N_359,In_4736,In_985);
and U360 (N_360,In_2103,In_1470);
nand U361 (N_361,In_2003,In_540);
or U362 (N_362,In_2953,In_2708);
nand U363 (N_363,In_3061,In_991);
nand U364 (N_364,In_267,In_2199);
nand U365 (N_365,In_4737,In_878);
nor U366 (N_366,In_485,In_3109);
xor U367 (N_367,In_4597,In_1811);
xor U368 (N_368,In_4832,In_4710);
and U369 (N_369,In_735,In_4841);
nor U370 (N_370,In_4564,In_1926);
xnor U371 (N_371,In_223,In_1979);
or U372 (N_372,In_4422,In_1713);
or U373 (N_373,In_1331,In_3141);
or U374 (N_374,In_3259,In_1627);
or U375 (N_375,In_1025,In_344);
or U376 (N_376,In_150,In_908);
xnor U377 (N_377,In_2859,In_4315);
and U378 (N_378,In_3185,In_4591);
nor U379 (N_379,In_385,In_3022);
xor U380 (N_380,In_3218,In_4431);
xnor U381 (N_381,In_505,In_3697);
and U382 (N_382,In_1447,In_460);
and U383 (N_383,In_2907,In_3850);
nor U384 (N_384,In_4038,In_4803);
nor U385 (N_385,In_4171,In_1192);
or U386 (N_386,In_1431,In_2665);
or U387 (N_387,In_4930,In_2177);
nor U388 (N_388,In_3636,In_3741);
xor U389 (N_389,In_192,In_2772);
nor U390 (N_390,In_1548,In_4938);
xnor U391 (N_391,In_912,In_2079);
xnor U392 (N_392,In_1940,In_1672);
nand U393 (N_393,In_3245,In_83);
or U394 (N_394,In_3133,In_4311);
nand U395 (N_395,In_3229,In_2294);
or U396 (N_396,In_4389,In_4772);
nor U397 (N_397,In_1759,In_1991);
nand U398 (N_398,In_3011,In_233);
and U399 (N_399,In_4049,In_3995);
xor U400 (N_400,In_224,In_3281);
xor U401 (N_401,In_1088,In_3333);
and U402 (N_402,In_536,In_4630);
nor U403 (N_403,In_1920,In_4555);
or U404 (N_404,In_2933,In_2981);
or U405 (N_405,In_4363,In_3066);
or U406 (N_406,In_414,In_242);
xnor U407 (N_407,In_499,In_4445);
xnor U408 (N_408,In_4773,In_449);
xnor U409 (N_409,In_112,In_2469);
nor U410 (N_410,In_1923,In_2104);
or U411 (N_411,In_3847,In_88);
xnor U412 (N_412,In_3330,In_557);
xnor U413 (N_413,In_3313,In_2071);
nor U414 (N_414,In_1945,In_303);
nor U415 (N_415,In_2261,In_4810);
nor U416 (N_416,In_4817,In_4951);
xnor U417 (N_417,In_3593,In_1338);
and U418 (N_418,In_4062,In_2042);
and U419 (N_419,In_1265,In_668);
nand U420 (N_420,In_2629,In_3563);
or U421 (N_421,In_3964,In_4354);
or U422 (N_422,In_4681,In_1916);
and U423 (N_423,In_889,In_376);
and U424 (N_424,In_1958,In_730);
and U425 (N_425,In_1038,In_4603);
nor U426 (N_426,In_2034,In_1228);
xor U427 (N_427,In_4546,In_670);
nor U428 (N_428,In_1663,In_177);
and U429 (N_429,In_2040,In_4103);
nor U430 (N_430,In_4179,In_2028);
nand U431 (N_431,In_613,In_57);
nand U432 (N_432,In_345,In_3269);
nor U433 (N_433,In_1325,In_2256);
and U434 (N_434,In_667,In_194);
nor U435 (N_435,In_4391,In_4970);
nand U436 (N_436,In_1039,In_3943);
or U437 (N_437,In_1905,In_616);
xor U438 (N_438,In_2897,In_3530);
nor U439 (N_439,In_2919,In_4730);
nand U440 (N_440,In_2746,In_3997);
xor U441 (N_441,In_3070,In_2527);
or U442 (N_442,In_4279,In_3774);
nand U443 (N_443,In_935,In_4018);
and U444 (N_444,In_4807,In_2258);
and U445 (N_445,In_2408,In_302);
or U446 (N_446,In_3179,In_3483);
nor U447 (N_447,In_2579,In_475);
or U448 (N_448,In_4044,In_2492);
or U449 (N_449,In_4721,In_3385);
nand U450 (N_450,In_3627,In_785);
or U451 (N_451,In_1211,In_2459);
xnor U452 (N_452,In_2316,In_3671);
nand U453 (N_453,In_3005,In_950);
nand U454 (N_454,In_4943,In_3503);
or U455 (N_455,In_4210,In_200);
or U456 (N_456,In_1756,In_4166);
nor U457 (N_457,In_3812,In_474);
or U458 (N_458,In_4614,In_2572);
nand U459 (N_459,In_3397,In_545);
or U460 (N_460,In_4990,In_558);
nand U461 (N_461,In_412,In_1873);
and U462 (N_462,In_1931,In_1681);
nor U463 (N_463,In_1654,In_1362);
xnor U464 (N_464,In_790,In_240);
nor U465 (N_465,In_1674,In_4353);
xnor U466 (N_466,In_1327,In_649);
nor U467 (N_467,In_1104,In_1166);
or U468 (N_468,In_4627,In_4072);
nand U469 (N_469,In_3416,In_1466);
xnor U470 (N_470,In_175,In_2087);
or U471 (N_471,In_1549,In_4805);
xor U472 (N_472,In_1123,In_2811);
or U473 (N_473,In_2875,In_2039);
nor U474 (N_474,In_1946,In_1237);
or U475 (N_475,In_1524,In_997);
and U476 (N_476,In_3556,In_578);
nand U477 (N_477,In_378,In_4811);
xnor U478 (N_478,In_1253,In_4646);
xor U479 (N_479,In_1729,In_3197);
and U480 (N_480,In_386,In_4651);
nand U481 (N_481,In_2417,In_630);
nand U482 (N_482,In_876,In_2747);
nand U483 (N_483,In_2842,In_1345);
nor U484 (N_484,In_2336,In_1155);
nand U485 (N_485,In_2141,In_4882);
nand U486 (N_486,In_3780,In_2069);
nand U487 (N_487,In_1602,In_3487);
nand U488 (N_488,In_1320,In_2283);
xor U489 (N_489,In_1188,In_1260);
nor U490 (N_490,In_3315,In_1854);
nor U491 (N_491,In_85,In_4147);
and U492 (N_492,In_3566,In_1225);
xnor U493 (N_493,In_4117,In_1494);
nor U494 (N_494,In_315,In_2926);
and U495 (N_495,In_157,In_3146);
or U496 (N_496,In_904,In_1838);
or U497 (N_497,In_4835,In_198);
and U498 (N_498,In_533,In_3370);
nand U499 (N_499,In_1139,In_2990);
and U500 (N_500,In_2084,In_2765);
and U501 (N_501,In_1737,In_4888);
and U502 (N_502,In_4402,In_4568);
or U503 (N_503,In_4579,In_1009);
xnor U504 (N_504,In_3846,In_4488);
xor U505 (N_505,In_763,In_831);
nor U506 (N_506,In_3309,In_1392);
and U507 (N_507,In_4259,In_2782);
nand U508 (N_508,In_227,In_4233);
xor U509 (N_509,In_3340,In_1151);
and U510 (N_510,In_2958,In_2573);
nand U511 (N_511,In_4872,In_713);
xor U512 (N_512,In_2969,In_4995);
nor U513 (N_513,In_1810,In_4024);
or U514 (N_514,In_1290,In_1469);
or U515 (N_515,In_1334,In_684);
xnor U516 (N_516,In_767,In_937);
nand U517 (N_517,In_577,In_2251);
nand U518 (N_518,In_1463,In_4727);
and U519 (N_519,In_3336,In_1200);
xor U520 (N_520,In_892,In_4476);
nand U521 (N_521,In_3959,In_3674);
xnor U522 (N_522,In_1014,In_3996);
or U523 (N_523,In_692,In_4278);
or U524 (N_524,In_1806,In_3386);
nand U525 (N_525,In_529,In_3970);
or U526 (N_526,In_2340,In_2282);
nor U527 (N_527,In_4560,In_1599);
nor U528 (N_528,In_170,In_1427);
nor U529 (N_529,In_640,In_2333);
xor U530 (N_530,In_2620,In_1891);
xor U531 (N_531,In_3734,In_4696);
xor U532 (N_532,In_2015,In_2948);
xnor U533 (N_533,In_3786,In_4284);
nor U534 (N_534,In_103,In_2217);
xnor U535 (N_535,In_508,In_993);
and U536 (N_536,In_144,In_2720);
nand U537 (N_537,In_3498,In_2150);
nand U538 (N_538,In_4369,In_4577);
nand U539 (N_539,In_3517,In_2216);
xor U540 (N_540,In_364,In_3399);
and U541 (N_541,In_3603,In_4408);
xnor U542 (N_542,In_2657,In_4997);
nand U543 (N_543,In_293,In_4336);
and U544 (N_544,In_398,In_1715);
nand U545 (N_545,In_3721,In_1018);
nand U546 (N_546,In_1143,In_3091);
xnor U547 (N_547,In_4785,In_1193);
nand U548 (N_548,In_3305,In_4847);
nor U549 (N_549,In_2520,In_3007);
nor U550 (N_550,In_4321,In_166);
xor U551 (N_551,In_11,In_3534);
and U552 (N_552,In_2383,In_3807);
and U553 (N_553,In_14,In_2667);
nand U554 (N_554,In_1657,In_3625);
or U555 (N_555,In_1816,In_3239);
or U556 (N_556,In_2026,In_4176);
nor U557 (N_557,In_350,In_2398);
nor U558 (N_558,In_3876,In_4347);
or U559 (N_559,In_2287,In_4578);
nand U560 (N_560,In_680,In_1774);
and U561 (N_561,In_424,In_1961);
or U562 (N_562,In_1178,In_2442);
xnor U563 (N_563,In_257,In_330);
xnor U564 (N_564,In_3087,In_1645);
xnor U565 (N_565,In_2706,In_1222);
and U566 (N_566,In_4755,In_3788);
and U567 (N_567,In_3999,In_4331);
and U568 (N_568,In_2164,In_2939);
or U569 (N_569,In_1135,In_999);
xnor U570 (N_570,In_2458,In_4569);
or U571 (N_571,In_4626,In_1581);
nand U572 (N_572,In_1206,In_2396);
xor U573 (N_573,In_1977,In_3658);
or U574 (N_574,In_4762,In_3521);
xnor U575 (N_575,In_3072,In_3737);
nor U576 (N_576,In_806,In_3726);
and U577 (N_577,In_4517,In_841);
and U578 (N_578,In_1117,In_116);
nand U579 (N_579,In_4485,In_4474);
or U580 (N_580,In_4705,In_4613);
nor U581 (N_581,In_3858,In_4858);
nand U582 (N_582,In_731,In_4531);
and U583 (N_583,In_2012,In_3466);
xnor U584 (N_584,In_3443,In_4473);
nand U585 (N_585,In_148,In_4089);
nor U586 (N_586,In_4534,In_3872);
or U587 (N_587,In_1727,In_3117);
and U588 (N_588,In_941,In_809);
or U589 (N_589,In_3188,In_2661);
or U590 (N_590,In_4953,In_4175);
and U591 (N_591,In_4843,In_1543);
nand U592 (N_592,In_4812,In_1377);
and U593 (N_593,In_3829,In_1284);
nor U594 (N_594,In_3240,In_2567);
or U595 (N_595,In_4448,In_4157);
and U596 (N_596,In_2202,In_1864);
nor U597 (N_597,In_4254,In_1138);
xnor U598 (N_598,In_3931,In_2402);
nor U599 (N_599,In_4253,In_1443);
xor U600 (N_600,In_4394,In_1775);
xnor U601 (N_601,In_4102,In_4936);
or U602 (N_602,In_916,In_4285);
nor U603 (N_603,In_3628,In_4230);
nand U604 (N_604,In_2591,In_4998);
xnor U605 (N_605,In_3208,In_4051);
nor U606 (N_606,In_433,In_93);
nand U607 (N_607,In_1792,In_4400);
nand U608 (N_608,In_856,In_837);
nand U609 (N_609,In_274,In_56);
nor U610 (N_610,In_3849,In_1888);
xnor U611 (N_611,In_3981,In_3394);
nor U612 (N_612,In_3597,In_4139);
nor U613 (N_613,In_3015,In_3884);
nor U614 (N_614,In_2539,In_1423);
nand U615 (N_615,In_1455,In_4205);
or U616 (N_616,In_2844,In_209);
xnor U617 (N_617,In_4104,In_984);
nand U618 (N_618,In_4874,In_2673);
or U619 (N_619,In_2890,In_3031);
xnor U620 (N_620,In_1530,In_1673);
xnor U621 (N_621,In_1566,In_1219);
nand U622 (N_622,In_1189,In_3704);
and U623 (N_623,In_2236,In_2731);
or U624 (N_624,In_1824,In_603);
nor U625 (N_625,In_4621,In_3756);
and U626 (N_626,In_1791,In_4468);
nor U627 (N_627,In_4971,In_2393);
and U628 (N_628,In_4093,In_2698);
xnor U629 (N_629,In_4099,In_1796);
and U630 (N_630,In_4409,In_1583);
nor U631 (N_631,In_2468,In_1144);
nor U632 (N_632,In_2696,In_243);
or U633 (N_633,In_423,In_3499);
xnor U634 (N_634,In_1187,In_1515);
nor U635 (N_635,In_1630,In_3822);
nand U636 (N_636,In_4477,In_4246);
nor U637 (N_637,In_771,In_2984);
or U638 (N_638,In_2808,In_2518);
nand U639 (N_639,In_1601,In_122);
and U640 (N_640,In_3234,In_551);
xnor U641 (N_641,In_1747,In_3888);
nand U642 (N_642,In_2265,In_1458);
xnor U643 (N_643,In_2936,In_2264);
or U644 (N_644,In_1924,In_3169);
nor U645 (N_645,In_2054,In_1959);
and U646 (N_646,In_3130,In_1690);
nand U647 (N_647,In_2846,In_1094);
or U648 (N_648,In_393,In_4683);
or U649 (N_649,In_1295,In_1164);
xor U650 (N_650,In_552,In_1286);
nand U651 (N_651,In_1709,In_3059);
and U652 (N_652,In_2538,In_636);
xnor U653 (N_653,In_3693,In_43);
or U654 (N_654,In_881,In_2477);
and U655 (N_655,In_1929,In_2358);
nand U656 (N_656,In_4161,In_4237);
nor U657 (N_657,In_1063,In_2472);
nand U658 (N_658,In_3595,In_1686);
nand U659 (N_659,In_2125,In_4232);
and U660 (N_660,In_1739,In_4650);
nand U661 (N_661,In_4223,In_4017);
nor U662 (N_662,In_2915,In_108);
xor U663 (N_663,In_3635,In_1843);
and U664 (N_664,In_3511,In_873);
or U665 (N_665,In_638,In_448);
and U666 (N_666,In_835,In_99);
and U667 (N_667,In_803,In_772);
nor U668 (N_668,In_4349,In_3899);
nand U669 (N_669,In_1308,In_78);
nor U670 (N_670,In_3157,In_1429);
nand U671 (N_671,In_2871,In_4191);
nand U672 (N_672,In_2147,In_146);
nand U673 (N_673,In_3830,In_3865);
and U674 (N_674,In_3119,In_3294);
xnor U675 (N_675,In_50,In_1662);
and U676 (N_676,In_1638,In_4550);
or U677 (N_677,In_759,In_4298);
nand U678 (N_678,In_1821,In_2170);
xor U679 (N_679,In_2851,In_3507);
or U680 (N_680,In_4659,In_2476);
and U681 (N_681,In_2369,In_4257);
nor U682 (N_682,In_1170,In_196);
or U683 (N_683,In_3922,In_1551);
and U684 (N_684,In_1848,In_2913);
nand U685 (N_685,In_486,In_3344);
xor U686 (N_686,In_1990,In_3751);
or U687 (N_687,In_1963,In_1728);
nor U688 (N_688,In_1574,In_1340);
or U689 (N_689,In_4433,In_361);
and U690 (N_690,In_572,In_1495);
nand U691 (N_691,In_2344,In_4245);
nor U692 (N_692,In_902,In_1480);
or U693 (N_693,In_3617,In_3461);
nor U694 (N_694,In_3699,In_2685);
nor U695 (N_695,In_4915,In_452);
and U696 (N_696,In_4107,In_3388);
or U697 (N_697,In_4671,In_811);
nor U698 (N_698,In_4016,In_1941);
and U699 (N_699,In_1199,In_2375);
nand U700 (N_700,In_2086,In_147);
and U701 (N_701,In_3244,In_1214);
nor U702 (N_702,In_4977,In_3422);
xor U703 (N_703,In_3480,In_2870);
nor U704 (N_704,In_1908,In_3969);
nand U705 (N_705,In_3752,In_4163);
or U706 (N_706,In_1127,In_652);
nor U707 (N_707,In_960,In_1092);
or U708 (N_708,In_202,In_3941);
nand U709 (N_709,In_3768,In_3949);
xnor U710 (N_710,In_1353,In_2292);
xor U711 (N_711,In_465,In_4043);
nand U712 (N_712,In_1393,In_3092);
xor U713 (N_713,In_4601,In_2497);
or U714 (N_714,In_2849,In_3250);
nand U715 (N_715,In_4058,In_1181);
xor U716 (N_716,In_1943,In_4806);
and U717 (N_717,In_2616,In_2838);
xnor U718 (N_718,In_573,In_1288);
or U719 (N_719,In_1315,In_2991);
nand U720 (N_720,In_4035,In_1486);
xnor U721 (N_721,In_4030,In_172);
nor U722 (N_722,In_1825,In_3465);
nor U723 (N_723,In_2883,In_2182);
nor U724 (N_724,In_611,In_3235);
and U725 (N_725,In_3112,In_4037);
xnor U726 (N_726,In_4379,In_4916);
xnor U727 (N_727,In_4376,In_126);
nor U728 (N_728,In_3611,In_73);
and U729 (N_729,In_1757,In_4013);
nor U730 (N_730,In_1884,In_3373);
xor U731 (N_731,In_4558,In_331);
nor U732 (N_732,In_4484,In_988);
nand U733 (N_733,In_2212,In_1880);
nand U734 (N_734,In_2288,In_54);
or U735 (N_735,In_1397,In_3319);
or U736 (N_736,In_2454,In_3893);
or U737 (N_737,In_4444,In_2221);
xnor U738 (N_738,In_2575,In_663);
xnor U739 (N_739,In_2770,In_3372);
nand U740 (N_740,In_4631,In_2585);
nor U741 (N_741,In_1893,In_741);
and U742 (N_742,In_955,In_975);
nand U743 (N_743,In_3114,In_208);
xor U744 (N_744,In_2544,In_3580);
xor U745 (N_745,In_1378,In_2475);
nor U746 (N_746,In_2565,In_3505);
and U747 (N_747,In_1651,In_2411);
xor U748 (N_748,In_2721,In_1575);
nand U749 (N_749,In_3698,In_1420);
xor U750 (N_750,In_909,In_2533);
nand U751 (N_751,In_4031,In_1054);
and U752 (N_752,In_1970,In_1303);
and U753 (N_753,In_4876,In_2686);
xnor U754 (N_754,In_775,In_39);
nand U755 (N_755,In_2412,In_1622);
and U756 (N_756,In_4396,In_1311);
nor U757 (N_757,In_1015,In_1563);
and U758 (N_758,In_2013,In_2432);
xnor U759 (N_759,In_3302,In_1236);
nand U760 (N_760,In_4085,In_4446);
nand U761 (N_761,In_2096,In_3150);
xnor U762 (N_762,In_1234,In_317);
xor U763 (N_763,In_635,In_2109);
nand U764 (N_764,In_4098,In_1832);
nor U765 (N_765,In_1565,In_2574);
and U766 (N_766,In_2788,In_384);
and U767 (N_767,In_2318,In_4933);
nor U768 (N_768,In_2252,In_4795);
xnor U769 (N_769,In_3776,In_1869);
and U770 (N_770,In_4213,In_4891);
and U771 (N_771,In_66,In_1544);
nor U772 (N_772,In_2855,In_4032);
and U773 (N_773,In_2168,In_930);
nor U774 (N_774,In_2628,In_1537);
and U775 (N_775,In_4182,In_247);
xor U776 (N_776,In_2293,In_4689);
and U777 (N_777,In_2262,In_994);
or U778 (N_778,In_2348,In_4377);
or U779 (N_779,In_4238,In_2327);
xor U780 (N_780,In_2183,In_3001);
nor U781 (N_781,In_3071,In_134);
nand U782 (N_782,In_4982,In_4411);
nor U783 (N_783,In_311,In_792);
or U784 (N_784,In_656,In_2810);
nand U785 (N_785,In_4511,In_4917);
xnor U786 (N_786,In_1696,In_495);
xnor U787 (N_787,In_1859,In_1386);
nand U788 (N_788,In_1538,In_3766);
or U789 (N_789,In_326,In_4920);
xnor U790 (N_790,In_2372,In_554);
nand U791 (N_791,In_288,In_3131);
nand U792 (N_792,In_1922,In_4976);
nor U793 (N_793,In_1158,In_3004);
or U794 (N_794,In_4981,In_3802);
nand U795 (N_795,In_2214,In_1736);
and U796 (N_796,In_750,In_4455);
or U797 (N_797,In_1987,In_2600);
xnor U798 (N_798,In_1034,In_1438);
xor U799 (N_799,In_1925,In_4980);
nand U800 (N_800,In_1610,In_4164);
nand U801 (N_801,In_105,In_4451);
or U802 (N_802,In_219,In_1702);
xnor U803 (N_803,In_3600,In_592);
and U804 (N_804,In_923,In_3021);
or U805 (N_805,In_1949,In_3729);
xnor U806 (N_806,In_1289,In_1274);
xor U807 (N_807,In_69,In_276);
xnor U808 (N_808,In_736,In_3474);
and U809 (N_809,In_3448,In_3415);
nor U810 (N_810,In_4112,In_513);
and U811 (N_811,In_1823,In_3369);
and U812 (N_812,In_249,In_2371);
nand U813 (N_813,In_4267,In_374);
nand U814 (N_814,In_2512,In_4884);
or U815 (N_815,In_4190,In_1317);
or U816 (N_816,In_943,In_4335);
and U817 (N_817,In_1381,In_1906);
xnor U818 (N_818,In_2550,In_199);
nand U819 (N_819,In_4923,In_4186);
or U820 (N_820,In_581,In_1247);
and U821 (N_821,In_4678,In_3939);
nor U822 (N_822,In_2643,In_4244);
or U823 (N_823,In_2868,In_4647);
nand U824 (N_824,In_4547,In_671);
xnor U825 (N_825,In_4260,In_4960);
nor U826 (N_826,In_4074,In_2775);
or U827 (N_827,In_2513,In_2359);
xor U828 (N_828,In_1632,In_4830);
xnor U829 (N_829,In_4420,In_3014);
nor U830 (N_830,In_1142,In_3703);
nand U831 (N_831,In_2205,In_948);
xnor U832 (N_832,In_970,In_632);
nand U833 (N_833,In_1745,In_3084);
or U834 (N_834,In_1001,In_4758);
xor U835 (N_835,In_2403,In_1780);
or U836 (N_836,In_765,In_2374);
xnor U837 (N_837,In_1457,In_1516);
nand U838 (N_838,In_443,In_3966);
nor U839 (N_839,In_372,In_653);
and U840 (N_840,In_995,In_2833);
nand U841 (N_841,In_965,In_3307);
xnor U842 (N_842,In_4834,In_2559);
nor U843 (N_843,In_2413,In_703);
nand U844 (N_844,In_1641,In_1382);
nor U845 (N_845,In_2223,In_4229);
xor U846 (N_846,In_3144,In_679);
and U847 (N_847,In_1232,In_3562);
xnor U848 (N_848,In_3099,In_3172);
or U849 (N_849,In_3993,In_3673);
nor U850 (N_850,In_4264,In_164);
and U851 (N_851,In_2938,In_618);
nand U852 (N_852,In_4324,In_109);
or U853 (N_853,In_2675,In_2111);
and U854 (N_854,In_2829,In_4852);
nor U855 (N_855,In_4174,In_4864);
nand U856 (N_856,In_2937,In_4881);
nor U857 (N_857,In_4941,In_2461);
nand U858 (N_858,In_4130,In_2975);
or U859 (N_859,In_98,In_2419);
nor U860 (N_860,In_183,In_1998);
or U861 (N_861,In_3518,In_1701);
and U862 (N_862,In_2658,In_1203);
xor U863 (N_863,In_4642,In_4809);
nor U864 (N_864,In_845,In_1350);
nand U865 (N_865,In_4596,In_3657);
nor U866 (N_866,In_1660,In_4702);
or U867 (N_867,In_519,In_1148);
nand U868 (N_868,In_880,In_301);
and U869 (N_869,In_3286,In_3972);
and U870 (N_870,In_1800,In_740);
nand U871 (N_871,In_4491,In_4152);
nor U872 (N_872,In_1513,In_2809);
xnor U873 (N_873,In_2100,In_3864);
xnor U874 (N_874,In_2624,In_3252);
and U875 (N_875,In_2790,In_2503);
nor U876 (N_876,In_2674,In_1975);
nand U877 (N_877,In_1416,In_159);
xor U878 (N_878,In_2598,In_1501);
nor U879 (N_879,In_4633,In_3221);
and U880 (N_880,In_3396,In_1936);
or U881 (N_881,In_2536,In_1840);
nand U882 (N_882,In_2989,In_891);
xor U883 (N_883,In_1626,In_2480);
nor U884 (N_884,In_3074,In_3292);
xor U885 (N_885,In_4961,In_286);
nor U886 (N_886,In_4565,In_4410);
nor U887 (N_887,In_1742,In_963);
nor U888 (N_888,In_4071,In_2734);
nand U889 (N_889,In_4094,In_4447);
or U890 (N_890,In_799,In_855);
xnor U891 (N_891,In_2785,In_1607);
and U892 (N_892,In_2806,In_1992);
nand U893 (N_893,In_617,In_297);
nor U894 (N_894,In_3078,In_2072);
or U895 (N_895,In_2699,In_2180);
and U896 (N_896,In_689,In_681);
xor U897 (N_897,In_3631,In_48);
nand U898 (N_898,In_3491,In_4660);
or U899 (N_899,In_4815,In_3983);
nor U900 (N_900,In_348,In_934);
and U901 (N_901,In_3076,In_1449);
xnor U902 (N_902,In_1868,In_3787);
or U903 (N_903,In_3036,In_1510);
and U904 (N_904,In_1464,In_3257);
xor U905 (N_905,In_2797,In_1976);
and U906 (N_906,In_4239,In_4201);
and U907 (N_907,In_3409,In_1133);
and U908 (N_908,In_3376,In_3243);
and U909 (N_909,In_4180,In_19);
and U910 (N_910,In_3322,In_2269);
and U911 (N_911,In_2603,In_4217);
nor U912 (N_912,In_2564,In_3712);
and U913 (N_913,In_1981,In_2486);
nor U914 (N_914,In_584,In_1697);
xnor U915 (N_915,In_338,In_4505);
and U916 (N_916,In_1557,In_2532);
nand U917 (N_917,In_4645,In_2771);
and U918 (N_918,In_2307,In_4002);
nand U919 (N_919,In_2812,In_3800);
and U920 (N_920,In_1011,In_674);
and U921 (N_921,In_3026,In_1100);
nor U922 (N_922,In_1186,In_2922);
or U923 (N_923,In_510,In_2093);
xor U924 (N_924,In_4092,In_2997);
nand U925 (N_925,In_4177,In_2113);
or U926 (N_926,In_3446,In_377);
or U927 (N_927,In_1161,In_359);
xor U928 (N_928,In_2959,In_2834);
xor U929 (N_929,In_2347,In_4623);
nand U930 (N_930,In_4383,In_4863);
nor U931 (N_931,In_2435,In_2376);
or U932 (N_932,In_2345,In_4390);
nand U933 (N_933,In_3546,In_2614);
nand U934 (N_934,In_905,In_3944);
and U935 (N_935,In_296,In_1703);
nor U936 (N_936,In_1561,In_661);
nand U937 (N_937,In_12,In_2547);
or U938 (N_938,In_3531,In_2479);
nand U939 (N_939,In_4575,In_3054);
and U940 (N_940,In_3508,In_3785);
nor U941 (N_941,In_594,In_281);
nor U942 (N_942,In_4136,In_3753);
and U943 (N_943,In_1665,In_3423);
nand U944 (N_944,In_145,In_4169);
and U945 (N_945,In_2779,In_3873);
and U946 (N_946,In_4993,In_1597);
and U947 (N_947,In_40,In_1078);
xor U948 (N_948,In_2740,In_4133);
nand U949 (N_949,In_2888,In_4672);
xor U950 (N_950,In_3145,In_2756);
nand U951 (N_951,In_4108,In_619);
xor U952 (N_952,In_2444,In_4828);
nor U953 (N_953,In_4948,In_4275);
and U954 (N_954,In_3216,In_3550);
or U955 (N_955,In_3909,In_3897);
nor U956 (N_956,In_2006,In_3192);
and U957 (N_957,In_4452,In_4889);
or U958 (N_958,In_3923,In_2189);
xor U959 (N_959,In_701,In_614);
or U960 (N_960,In_798,In_4308);
xnor U961 (N_961,In_402,In_2401);
nand U962 (N_962,In_1109,In_3916);
xnor U963 (N_963,In_1874,In_2062);
and U964 (N_964,In_4235,In_4989);
nand U965 (N_965,In_3510,In_518);
xor U966 (N_966,In_1271,In_4052);
nand U967 (N_967,In_205,In_461);
nor U968 (N_968,In_1478,In_2776);
nand U969 (N_969,In_1424,In_1684);
and U970 (N_970,In_1582,In_3526);
and U971 (N_971,In_2387,In_1877);
nor U972 (N_972,In_804,In_277);
xnor U973 (N_973,In_155,In_3056);
nand U974 (N_974,In_3696,In_2030);
nor U975 (N_975,In_2175,In_690);
nand U976 (N_976,In_2385,In_787);
nor U977 (N_977,In_4946,In_1795);
or U978 (N_978,In_4712,In_426);
or U979 (N_979,In_254,In_3564);
and U980 (N_980,In_51,In_3098);
and U981 (N_981,In_2633,In_895);
and U982 (N_982,In_532,In_1006);
nor U983 (N_983,In_3806,In_1168);
nor U984 (N_984,In_1870,In_2943);
and U985 (N_985,In_4611,In_2787);
nand U986 (N_986,In_608,In_2678);
and U987 (N_987,In_665,In_1579);
xor U988 (N_988,In_2957,In_4572);
nor U989 (N_989,In_2886,In_264);
and U990 (N_990,In_4865,In_875);
nor U991 (N_991,In_1209,In_877);
or U992 (N_992,In_4299,In_1150);
and U993 (N_993,In_1369,In_3542);
nand U994 (N_994,In_1344,In_3623);
or U995 (N_995,In_2732,In_3514);
nor U996 (N_996,In_3545,In_3428);
xor U997 (N_997,In_1277,In_1500);
and U998 (N_998,In_3214,In_1896);
xnor U999 (N_999,In_2163,In_2305);
xnor U1000 (N_1000,In_2761,In_1444);
nor U1001 (N_1001,In_4509,In_1572);
nor U1002 (N_1002,In_401,In_2745);
nand U1003 (N_1003,In_4240,In_784);
and U1004 (N_1004,In_4728,In_1089);
xnor U1005 (N_1005,In_4711,In_3979);
xnor U1006 (N_1006,In_1073,In_1097);
nor U1007 (N_1007,In_682,In_932);
nor U1008 (N_1008,In_1086,In_4768);
xnor U1009 (N_1009,In_3629,In_4673);
nand U1010 (N_1010,In_893,In_1570);
nand U1011 (N_1011,In_1621,In_1554);
or U1012 (N_1012,In_766,In_4934);
or U1013 (N_1013,In_4075,In_535);
xor U1014 (N_1014,In_3028,In_1475);
nand U1015 (N_1015,In_2716,In_4604);
nor U1016 (N_1016,In_898,In_2687);
xor U1017 (N_1017,In_29,In_3331);
nor U1018 (N_1018,In_2697,In_4931);
and U1019 (N_1019,In_2606,In_92);
nand U1020 (N_1020,In_2556,In_380);
nand U1021 (N_1021,In_4533,In_3578);
nand U1022 (N_1022,In_2737,In_3664);
xor U1023 (N_1023,In_1615,In_4706);
nor U1024 (N_1024,In_74,In_4393);
or U1025 (N_1025,In_1506,In_2738);
xor U1026 (N_1026,In_2854,In_1384);
nor U1027 (N_1027,In_167,In_2196);
xnor U1028 (N_1028,In_2793,In_3265);
xnor U1029 (N_1029,In_2382,In_2186);
and U1030 (N_1030,In_3469,In_3927);
xnor U1031 (N_1031,In_894,In_1456);
or U1032 (N_1032,In_2074,In_1772);
nand U1033 (N_1033,In_4655,In_1754);
and U1034 (N_1034,In_1966,In_2881);
and U1035 (N_1035,In_4271,In_1040);
nand U1036 (N_1036,In_324,In_4859);
nor U1037 (N_1037,In_347,In_4126);
or U1038 (N_1038,In_1302,In_828);
nand U1039 (N_1039,In_1467,In_1711);
nor U1040 (N_1040,In_810,In_1831);
xnor U1041 (N_1041,In_2932,In_3090);
nor U1042 (N_1042,In_4718,In_0);
xnor U1043 (N_1043,In_4082,In_46);
nand U1044 (N_1044,In_858,In_2328);
xor U1045 (N_1045,In_4620,In_2587);
and U1046 (N_1046,In_3574,In_2802);
xnor U1047 (N_1047,In_1822,In_1184);
nor U1048 (N_1048,In_660,In_3702);
nor U1049 (N_1049,In_774,In_2666);
xor U1050 (N_1050,In_1398,In_2233);
or U1051 (N_1051,In_4269,In_1243);
xor U1052 (N_1052,In_4771,In_1573);
and U1053 (N_1053,In_2090,In_4137);
and U1054 (N_1054,In_1556,In_466);
xor U1055 (N_1055,In_4788,In_329);
nand U1056 (N_1056,In_2137,In_4355);
nand U1057 (N_1057,In_436,In_1856);
or U1058 (N_1058,In_2784,In_4719);
nor U1059 (N_1059,In_4986,In_633);
nand U1060 (N_1060,In_4185,In_4301);
nor U1061 (N_1061,In_250,In_3453);
nand U1062 (N_1062,In_396,In_1770);
nand U1063 (N_1063,In_2149,In_3820);
and U1064 (N_1064,In_872,In_4849);
nand U1065 (N_1065,In_3760,In_851);
and U1066 (N_1066,In_2944,In_544);
nor U1067 (N_1067,In_3575,In_1330);
nor U1068 (N_1068,In_650,In_2506);
or U1069 (N_1069,In_1107,In_3043);
nor U1070 (N_1070,In_35,In_55);
nand U1071 (N_1071,In_1176,In_1815);
nor U1072 (N_1072,In_4346,In_1208);
xor U1073 (N_1073,In_1385,In_464);
or U1074 (N_1074,In_1301,In_1985);
xor U1075 (N_1075,In_4064,In_1132);
nand U1076 (N_1076,In_4640,In_628);
nor U1077 (N_1077,In_4442,In_3407);
xor U1078 (N_1078,In_2622,In_158);
xnor U1079 (N_1079,In_4536,In_654);
or U1080 (N_1080,In_3482,In_1147);
nand U1081 (N_1081,In_4138,In_2105);
xnor U1082 (N_1082,In_3306,In_4450);
nand U1083 (N_1083,In_1813,In_4243);
nor U1084 (N_1084,In_1299,In_1503);
and U1085 (N_1085,In_4679,In_2595);
xnor U1086 (N_1086,In_4539,In_1667);
xor U1087 (N_1087,In_2824,In_1928);
xnor U1088 (N_1088,In_4632,In_333);
or U1089 (N_1089,In_2546,In_3573);
xnor U1090 (N_1090,In_791,In_1664);
or U1091 (N_1091,In_2452,In_4624);
nand U1092 (N_1092,In_595,In_3473);
and U1093 (N_1093,In_2940,In_3588);
and U1094 (N_1094,In_1740,In_4367);
or U1095 (N_1095,In_2712,In_2557);
xor U1096 (N_1096,In_4029,In_2612);
xor U1097 (N_1097,In_4905,In_2045);
nand U1098 (N_1098,In_6,In_3247);
or U1099 (N_1099,In_981,In_958);
xnor U1100 (N_1100,In_4819,In_1191);
and U1101 (N_1101,In_1298,In_4729);
and U1102 (N_1102,In_3582,In_3348);
or U1103 (N_1103,In_3324,In_2604);
nor U1104 (N_1104,In_4263,In_3326);
or U1105 (N_1105,In_4567,In_3290);
or U1106 (N_1106,In_4026,In_1179);
or U1107 (N_1107,In_4392,In_926);
and U1108 (N_1108,In_4512,In_967);
nand U1109 (N_1109,In_2578,In_1351);
and U1110 (N_1110,In_4305,In_4060);
or U1111 (N_1111,In_4430,In_1699);
or U1112 (N_1112,In_1305,In_4924);
or U1113 (N_1113,In_1769,In_1751);
and U1114 (N_1114,In_2653,In_1062);
and U1115 (N_1115,In_2852,In_770);
nor U1116 (N_1116,In_4760,In_2609);
nand U1117 (N_1117,In_3260,In_367);
and U1118 (N_1118,In_3801,In_3304);
nor U1119 (N_1119,In_1162,In_4041);
nor U1120 (N_1120,In_2247,In_1087);
nor U1121 (N_1121,In_3255,In_4362);
xor U1122 (N_1122,In_4214,In_3690);
xor U1123 (N_1123,In_1718,In_2902);
nor U1124 (N_1124,In_2500,In_4365);
or U1125 (N_1125,In_2478,In_1046);
nor U1126 (N_1126,In_2860,In_306);
and U1127 (N_1127,In_4310,In_289);
nand U1128 (N_1128,In_2651,In_4206);
or U1129 (N_1129,In_4722,In_795);
xor U1130 (N_1130,In_2117,In_3679);
and U1131 (N_1131,In_3215,In_1910);
nor U1132 (N_1132,In_1593,In_897);
nor U1133 (N_1133,In_3452,In_4753);
nand U1134 (N_1134,In_4777,In_3223);
nand U1135 (N_1135,In_2704,In_1356);
nor U1136 (N_1136,In_4199,In_2548);
and U1137 (N_1137,In_2901,In_818);
or U1138 (N_1138,In_1068,In_371);
xor U1139 (N_1139,In_2517,In_1282);
xnor U1140 (N_1140,In_2433,In_2923);
or U1141 (N_1141,In_1070,In_2056);
nand U1142 (N_1142,In_2952,In_4494);
xnor U1143 (N_1143,In_3610,In_1153);
nand U1144 (N_1144,In_395,In_2610);
nor U1145 (N_1145,In_1347,In_3525);
xor U1146 (N_1146,In_4499,In_3113);
xnor U1147 (N_1147,In_3353,In_2646);
nor U1148 (N_1148,In_4348,In_2108);
nor U1149 (N_1149,In_2593,In_3063);
nor U1150 (N_1150,In_4966,In_3468);
nand U1151 (N_1151,In_3523,In_2640);
nand U1152 (N_1152,In_3278,In_4842);
or U1153 (N_1153,In_4288,In_962);
nor U1154 (N_1154,In_1890,In_4716);
xnor U1155 (N_1155,In_4743,In_641);
xor U1156 (N_1156,In_4529,In_111);
xor U1157 (N_1157,In_3777,In_2543);
nand U1158 (N_1158,In_4067,In_1055);
xnor U1159 (N_1159,In_3289,In_2346);
nand U1160 (N_1160,In_2792,In_4921);
and U1161 (N_1161,In_1453,In_4005);
and U1162 (N_1162,In_3612,In_4211);
nor U1163 (N_1163,In_4792,In_4829);
and U1164 (N_1164,In_1182,In_59);
or U1165 (N_1165,In_1108,In_211);
nand U1166 (N_1166,In_862,In_1947);
or U1167 (N_1167,In_1955,In_3813);
or U1168 (N_1168,In_4735,In_3359);
or U1169 (N_1169,In_1474,In_2296);
nor U1170 (N_1170,In_1028,In_2615);
and U1171 (N_1171,In_3426,In_1617);
xnor U1172 (N_1172,In_1110,In_1069);
or U1173 (N_1173,In_1185,In_4731);
or U1174 (N_1174,In_1257,In_3670);
and U1175 (N_1175,In_4192,In_3641);
xnor U1176 (N_1176,In_2896,In_1471);
or U1177 (N_1177,In_222,In_4270);
and U1178 (N_1178,In_2912,In_2167);
nand U1179 (N_1179,In_3271,In_1217);
xnor U1180 (N_1180,In_169,In_3477);
and U1181 (N_1181,In_579,In_4766);
or U1182 (N_1182,In_2427,In_2154);
and U1183 (N_1183,In_471,In_977);
and U1184 (N_1184,In_1611,In_4500);
or U1185 (N_1185,In_1075,In_1488);
nand U1186 (N_1186,In_3749,In_3444);
and U1187 (N_1187,In_3083,In_973);
xor U1188 (N_1188,In_4073,In_1889);
nand U1189 (N_1189,In_3387,In_278);
or U1190 (N_1190,In_2184,In_3955);
or U1191 (N_1191,In_1600,In_168);
nand U1192 (N_1192,In_2098,In_2576);
or U1193 (N_1193,In_1116,In_3183);
nand U1194 (N_1194,In_4143,In_1541);
nor U1195 (N_1195,In_4790,In_3878);
xnor U1196 (N_1196,In_4501,In_1857);
nor U1197 (N_1197,In_2023,In_4384);
and U1198 (N_1198,In_2360,In_1881);
or U1199 (N_1199,In_2138,In_4426);
nand U1200 (N_1200,In_1846,In_3901);
nor U1201 (N_1201,In_3430,In_4974);
nand U1202 (N_1202,In_2089,In_1835);
or U1203 (N_1203,In_4955,In_4827);
or U1204 (N_1204,In_3295,In_136);
nand U1205 (N_1205,In_4453,In_3316);
nor U1206 (N_1206,In_1399,In_3492);
and U1207 (N_1207,In_899,In_3057);
or U1208 (N_1208,In_1252,In_2021);
and U1209 (N_1209,In_3975,In_2116);
xor U1210 (N_1210,In_2226,In_1552);
xnor U1211 (N_1211,In_3817,In_2553);
nor U1212 (N_1212,In_1058,In_1160);
xor U1213 (N_1213,In_284,In_4541);
or U1214 (N_1214,In_1609,In_366);
xnor U1215 (N_1215,In_4330,In_3938);
xor U1216 (N_1216,In_4813,In_762);
or U1217 (N_1217,In_2965,In_2662);
or U1218 (N_1218,In_2400,In_734);
nand U1219 (N_1219,In_4530,In_2326);
xnor U1220 (N_1220,In_2381,In_241);
xor U1221 (N_1221,In_4398,In_1559);
and U1222 (N_1222,In_4352,In_1712);
or U1223 (N_1223,In_2682,In_473);
nand U1224 (N_1224,In_801,In_4794);
nor U1225 (N_1225,In_1216,In_827);
xor U1226 (N_1226,In_2983,In_3205);
nor U1227 (N_1227,In_493,In_2768);
and U1228 (N_1228,In_1226,In_2521);
or U1229 (N_1229,In_2580,In_1002);
nand U1230 (N_1230,In_131,In_733);
nand U1231 (N_1231,In_3821,In_3648);
nand U1232 (N_1232,In_672,In_1724);
xnor U1233 (N_1233,In_2876,In_498);
nand U1234 (N_1234,In_720,In_4625);
xor U1235 (N_1235,In_416,In_3962);
or U1236 (N_1236,In_2722,In_1095);
xor U1237 (N_1237,In_2856,In_3456);
nor U1238 (N_1238,In_139,In_2008);
nor U1239 (N_1239,In_3236,In_42);
or U1240 (N_1240,In_2974,In_490);
nor U1241 (N_1241,In_4850,In_4906);
or U1242 (N_1242,In_4128,In_3902);
nor U1243 (N_1243,In_3986,In_4967);
or U1244 (N_1244,In_2397,In_2195);
xor U1245 (N_1245,In_2820,In_4559);
or U1246 (N_1246,In_3232,In_2315);
and U1247 (N_1247,In_4857,In_3334);
and U1248 (N_1248,In_700,In_4740);
nor U1249 (N_1249,In_2627,In_2725);
nand U1250 (N_1250,In_411,In_1254);
and U1251 (N_1251,In_838,In_4879);
or U1252 (N_1252,In_1934,In_3769);
and U1253 (N_1253,In_4911,In_2171);
and U1254 (N_1254,In_4300,In_1072);
nand U1255 (N_1255,In_2373,In_2757);
xnor U1256 (N_1256,In_751,In_1839);
or U1257 (N_1257,In_1951,In_4644);
nand U1258 (N_1258,In_3637,In_3935);
nor U1259 (N_1259,In_658,In_4739);
nand U1260 (N_1260,In_1173,In_3450);
nand U1261 (N_1261,In_2688,In_588);
xor U1262 (N_1262,In_4844,In_3206);
xnor U1263 (N_1263,In_1407,In_2955);
nor U1264 (N_1264,In_542,In_1999);
xor U1265 (N_1265,In_180,In_3101);
and U1266 (N_1266,In_3520,In_4676);
or U1267 (N_1267,In_4159,In_2878);
nor U1268 (N_1268,In_3988,In_743);
or U1269 (N_1269,In_706,In_4958);
or U1270 (N_1270,In_3608,In_3859);
or U1271 (N_1271,In_4056,In_1689);
nor U1272 (N_1272,In_2014,In_2455);
xnor U1273 (N_1273,In_3707,In_996);
nand U1274 (N_1274,In_4540,In_2356);
nand U1275 (N_1275,In_1670,In_1440);
and U1276 (N_1276,In_2510,In_1562);
and U1277 (N_1277,In_2899,In_1283);
xor U1278 (N_1278,In_2924,In_3950);
and U1279 (N_1279,In_3791,In_3120);
nor U1280 (N_1280,In_1678,In_2446);
nor U1281 (N_1281,In_4618,In_3463);
and U1282 (N_1282,In_321,In_1595);
nand U1283 (N_1283,In_4314,In_4713);
and U1284 (N_1284,In_3991,In_620);
nor U1285 (N_1285,In_204,In_1390);
nand U1286 (N_1286,In_516,In_896);
nand U1287 (N_1287,In_2416,In_1808);
nor U1288 (N_1288,In_3191,In_138);
and U1289 (N_1289,In_3515,In_4940);
xor U1290 (N_1290,In_915,In_4414);
and U1291 (N_1291,In_323,In_2701);
nand U1292 (N_1292,In_1085,In_1619);
nand U1293 (N_1293,In_237,In_647);
nor U1294 (N_1294,In_2894,In_480);
nor U1295 (N_1295,In_4415,In_3933);
or U1296 (N_1296,In_2133,In_207);
or U1297 (N_1297,In_3589,In_2560);
nand U1298 (N_1298,In_1174,In_444);
nand U1299 (N_1299,In_4554,In_3156);
nor U1300 (N_1300,In_1352,In_3881);
nor U1301 (N_1301,In_4127,In_2027);
nand U1302 (N_1302,In_2502,In_239);
nand U1303 (N_1303,In_781,In_786);
or U1304 (N_1304,In_2207,In_2817);
nor U1305 (N_1305,In_4610,In_3180);
nor U1306 (N_1306,In_1008,In_850);
nand U1307 (N_1307,In_4898,In_1140);
or U1308 (N_1308,In_3135,In_2805);
nand U1309 (N_1309,In_2181,In_4757);
or U1310 (N_1310,In_4014,In_467);
or U1311 (N_1311,In_3971,In_3127);
nand U1312 (N_1312,In_4387,In_420);
xor U1313 (N_1313,In_292,In_4039);
and U1314 (N_1314,In_570,In_4296);
nand U1315 (N_1315,In_3604,In_4814);
xnor U1316 (N_1316,In_4667,In_124);
or U1317 (N_1317,In_238,In_1125);
xor U1318 (N_1318,In_3789,In_1564);
xor U1319 (N_1319,In_4273,In_3280);
nand U1320 (N_1320,In_1616,In_2760);
and U1321 (N_1321,In_4675,In_2735);
or U1322 (N_1322,In_1983,In_3458);
nor U1323 (N_1323,In_4886,In_4373);
nand U1324 (N_1324,In_571,In_4747);
nor U1325 (N_1325,In_4219,In_4250);
xnor U1326 (N_1326,In_1518,In_3656);
nand U1327 (N_1327,In_778,In_1790);
or U1328 (N_1328,In_26,In_1468);
and U1329 (N_1329,In_87,In_3279);
nand U1330 (N_1330,In_553,In_3967);
nor U1331 (N_1331,In_2009,In_4386);
or U1332 (N_1332,In_123,In_1935);
or U1333 (N_1333,In_3558,In_3609);
and U1334 (N_1334,In_576,In_3775);
nand U1335 (N_1335,In_4076,In_3583);
nor U1336 (N_1336,In_2115,In_1430);
xor U1337 (N_1337,In_2464,In_388);
and U1338 (N_1338,In_1367,In_4146);
xor U1339 (N_1339,In_1969,In_2044);
xnor U1340 (N_1340,In_678,In_4542);
and U1341 (N_1341,In_2748,In_1589);
and U1342 (N_1342,In_2801,In_3952);
nor U1343 (N_1343,In_3682,In_3795);
or U1344 (N_1344,In_1833,In_2839);
nor U1345 (N_1345,In_1404,In_3842);
and U1346 (N_1346,In_1988,In_439);
nand U1347 (N_1347,In_1695,In_3410);
nor U1348 (N_1348,In_1504,In_2271);
nand U1349 (N_1349,In_4312,In_53);
or U1350 (N_1350,In_125,In_2537);
or U1351 (N_1351,In_2487,In_3195);
nand U1352 (N_1352,In_3809,In_823);
nand U1353 (N_1353,In_4878,In_2866);
nand U1354 (N_1354,In_3134,In_4184);
xnor U1355 (N_1355,In_3495,In_3166);
xor U1356 (N_1356,In_2407,In_812);
and U1357 (N_1357,In_3314,In_2127);
nand U1358 (N_1358,In_857,In_956);
xnor U1359 (N_1359,In_921,In_3479);
xor U1360 (N_1360,In_2052,In_455);
or U1361 (N_1361,In_3716,In_3408);
nor U1362 (N_1362,In_2967,In_1402);
nor U1363 (N_1363,In_808,In_1932);
nor U1364 (N_1364,In_4218,In_1465);
and U1365 (N_1365,In_1115,In_2337);
nand U1366 (N_1366,In_1473,In_3645);
nand U1367 (N_1367,In_4767,In_1558);
nand U1368 (N_1368,In_221,In_3961);
nand U1369 (N_1369,In_2322,In_1847);
nor U1370 (N_1370,In_959,In_3357);
nor U1371 (N_1371,In_1359,In_3038);
and U1372 (N_1372,In_3335,In_1041);
xnor U1373 (N_1373,In_1980,In_2692);
nand U1374 (N_1374,In_2130,In_4649);
nor U1375 (N_1375,In_3142,In_4432);
xnor U1376 (N_1376,In_4520,In_3237);
nor U1377 (N_1377,In_4944,In_3437);
nand U1378 (N_1378,In_2485,In_4848);
xnor U1379 (N_1379,In_1918,In_677);
nand U1380 (N_1380,In_1555,In_2715);
nor U1381 (N_1381,In_4087,In_2156);
or U1382 (N_1382,In_1448,In_4979);
xnor U1383 (N_1383,In_1105,In_2786);
and U1384 (N_1384,In_2588,In_4114);
or U1385 (N_1385,In_2645,In_969);
or U1386 (N_1386,In_4274,In_2102);
nand U1387 (N_1387,In_954,In_3770);
and U1388 (N_1388,In_1917,In_3980);
and U1389 (N_1389,In_3513,In_322);
and U1390 (N_1390,In_3162,In_3488);
nor U1391 (N_1391,In_1771,In_4751);
xor U1392 (N_1392,In_531,In_727);
xor U1393 (N_1393,In_3159,In_1967);
or U1394 (N_1394,In_3360,In_3506);
nor U1395 (N_1395,In_3201,In_3748);
or U1396 (N_1396,In_4698,In_541);
nor U1397 (N_1397,In_3058,In_2608);
nand U1398 (N_1398,In_1112,In_637);
nor U1399 (N_1399,In_1029,In_1451);
nand U1400 (N_1400,In_1309,In_4573);
and U1401 (N_1401,In_422,In_3605);
or U1402 (N_1402,In_4088,In_1623);
or U1403 (N_1403,In_1647,In_3926);
or U1404 (N_1404,In_3375,In_2276);
or U1405 (N_1405,In_3012,In_3069);
or U1406 (N_1406,In_3883,In_4521);
or U1407 (N_1407,In_538,In_3887);
or U1408 (N_1408,In_3125,In_1904);
nor U1409 (N_1409,In_1911,In_2451);
and U1410 (N_1410,In_1519,In_1865);
or U1411 (N_1411,In_4694,In_698);
nand U1412 (N_1412,In_22,In_2763);
and U1413 (N_1413,In_4302,In_4231);
xnor U1414 (N_1414,In_417,In_2355);
nor U1415 (N_1415,In_1061,In_4463);
or U1416 (N_1416,In_235,In_1306);
nor U1417 (N_1417,In_31,In_4113);
or U1418 (N_1418,In_2867,In_503);
xnor U1419 (N_1419,In_3695,In_4011);
nand U1420 (N_1420,In_1546,In_1594);
nand U1421 (N_1421,In_2554,In_3692);
nor U1422 (N_1422,In_2081,In_3262);
nor U1423 (N_1423,In_3323,In_709);
nand U1424 (N_1424,In_4115,In_900);
or U1425 (N_1425,In_4840,In_3592);
and U1426 (N_1426,In_4319,In_2909);
and U1427 (N_1427,In_62,In_3621);
and U1428 (N_1428,In_4483,In_1532);
nand U1429 (N_1429,In_777,In_397);
nor U1430 (N_1430,In_1047,In_20);
xnor U1431 (N_1431,In_1278,In_1375);
or U1432 (N_1432,In_1719,In_820);
or U1433 (N_1433,In_1973,In_3104);
nor U1434 (N_1434,In_2928,In_2050);
nor U1435 (N_1435,In_4419,In_3053);
or U1436 (N_1436,In_3065,In_325);
or U1437 (N_1437,In_566,In_3095);
or U1438 (N_1438,In_4228,In_4502);
nor U1439 (N_1439,In_3516,In_3904);
and U1440 (N_1440,In_1417,In_3009);
nor U1441 (N_1441,In_392,In_4078);
or U1442 (N_1442,In_3389,In_4368);
or U1443 (N_1443,In_3644,In_4778);
xnor U1444 (N_1444,In_4818,In_946);
xnor U1445 (N_1445,In_1201,In_4808);
xnor U1446 (N_1446,In_3778,In_2729);
nor U1447 (N_1447,In_3051,In_1368);
or U1448 (N_1448,In_3910,In_4877);
xor U1449 (N_1449,In_2581,In_968);
nor U1450 (N_1450,In_3449,In_606);
and U1451 (N_1451,In_4012,In_2611);
nor U1452 (N_1452,In_130,In_2357);
nor U1453 (N_1453,In_379,In_4148);
xor U1454 (N_1454,In_4220,In_2430);
nand U1455 (N_1455,In_4221,In_4256);
or U1456 (N_1456,In_3167,In_598);
nand U1457 (N_1457,In_21,In_2654);
nor U1458 (N_1458,In_2174,In_2869);
and U1459 (N_1459,In_1523,In_1871);
or U1460 (N_1460,In_755,In_1297);
and U1461 (N_1461,In_3541,In_555);
nor U1462 (N_1462,In_4487,In_2275);
xor U1463 (N_1463,In_1640,In_3651);
nand U1464 (N_1464,In_4833,In_848);
nand U1465 (N_1465,In_2317,In_2301);
xnor U1466 (N_1466,In_262,In_2140);
nand U1467 (N_1467,In_1978,In_4323);
nand U1468 (N_1468,In_2225,In_1786);
nor U1469 (N_1469,In_173,In_2249);
xor U1470 (N_1470,In_1183,In_2599);
nor U1471 (N_1471,In_1900,In_3655);
nor U1472 (N_1472,In_747,In_3797);
or U1473 (N_1473,In_813,In_4748);
nor U1474 (N_1474,In_830,In_3393);
nand U1475 (N_1475,In_3879,In_3017);
or U1476 (N_1476,In_1855,In_2529);
or U1477 (N_1477,In_128,In_1953);
nor U1478 (N_1478,In_1644,In_4682);
and U1479 (N_1479,In_816,In_869);
or U1480 (N_1480,In_4744,In_328);
nor U1481 (N_1481,In_3973,In_2342);
and U1482 (N_1482,In_2289,In_2244);
nor U1483 (N_1483,In_3427,In_2379);
and U1484 (N_1484,In_4129,In_4069);
or U1485 (N_1485,In_3880,In_3937);
xor U1486 (N_1486,In_2777,In_2319);
nor U1487 (N_1487,In_4036,In_3987);
nor U1488 (N_1488,In_890,In_2332);
or U1489 (N_1489,In_3196,In_3277);
nand U1490 (N_1490,In_4837,In_3462);
and U1491 (N_1491,In_1400,In_539);
nor U1492 (N_1492,In_3165,In_1082);
nor U1493 (N_1493,In_2807,In_4692);
and U1494 (N_1494,In_1646,In_3680);
nor U1495 (N_1495,In_4466,In_4413);
and U1496 (N_1496,In_488,In_1643);
or U1497 (N_1497,In_1698,In_4374);
and U1498 (N_1498,In_3814,In_822);
xnor U1499 (N_1499,In_1130,In_4034);
nand U1500 (N_1500,In_4460,In_2172);
and U1501 (N_1501,In_1785,In_362);
nor U1502 (N_1502,In_4196,In_2496);
and U1503 (N_1503,In_3160,In_3740);
xor U1504 (N_1504,In_1401,In_299);
nor U1505 (N_1505,In_4022,In_4797);
nor U1506 (N_1506,In_4423,In_1169);
xor U1507 (N_1507,In_4249,In_2422);
or U1508 (N_1508,In_840,In_4964);
and U1509 (N_1509,In_3624,In_1207);
nand U1510 (N_1510,In_2914,In_753);
or U1511 (N_1511,In_2693,In_2022);
nor U1512 (N_1512,In_1861,In_4996);
nand U1513 (N_1513,In_527,In_2123);
and U1514 (N_1514,In_4590,In_1608);
nor U1515 (N_1515,In_3489,In_3137);
and U1516 (N_1516,In_918,In_4869);
and U1517 (N_1517,In_693,In_4714);
or U1518 (N_1518,In_4010,In_2999);
nand U1519 (N_1519,In_58,In_3638);
xnor U1520 (N_1520,In_2423,In_3632);
and U1521 (N_1521,In_863,In_4100);
xnor U1522 (N_1522,In_1768,In_1614);
nor U1523 (N_1523,In_3896,In_4141);
and U1524 (N_1524,In_3833,In_149);
or U1525 (N_1525,In_2018,In_2966);
or U1526 (N_1526,In_4047,In_1818);
nand U1527 (N_1527,In_2011,In_4366);
xor U1528 (N_1528,In_3401,In_3233);
nand U1529 (N_1529,In_2122,In_639);
and U1530 (N_1530,In_4458,In_337);
and U1531 (N_1531,In_3731,In_4053);
nor U1532 (N_1532,In_1294,In_3475);
nand U1533 (N_1533,In_2368,In_1114);
and U1534 (N_1534,In_3677,In_717);
and U1535 (N_1535,In_3659,In_3738);
nor U1536 (N_1536,In_3033,In_1587);
and U1537 (N_1537,In_1634,In_2753);
xor U1538 (N_1538,In_1789,In_2522);
xnor U1539 (N_1539,In_3016,In_2055);
nor U1540 (N_1540,In_3400,In_852);
xnor U1541 (N_1541,In_2304,In_1521);
xnor U1542 (N_1542,In_1571,In_4901);
and U1543 (N_1543,In_604,In_231);
nor U1544 (N_1544,In_2911,In_4880);
nand U1545 (N_1545,In_972,In_2873);
or U1546 (N_1546,In_4497,In_524);
and U1547 (N_1547,In_2509,In_651);
and U1548 (N_1548,In_4170,In_3500);
nor U1549 (N_1549,In_1883,In_1279);
or U1550 (N_1550,In_1180,In_4403);
or U1551 (N_1551,In_1287,In_4909);
and U1552 (N_1552,In_1137,In_203);
and U1553 (N_1553,In_4913,In_351);
xor U1554 (N_1554,In_1491,In_4922);
nand U1555 (N_1555,In_2388,In_3755);
nand U1556 (N_1556,In_4912,In_3432);
xnor U1557 (N_1557,In_84,In_556);
nor U1558 (N_1558,In_3472,In_2142);
nor U1559 (N_1559,In_1291,In_1016);
nand U1560 (N_1560,In_2650,In_210);
and U1561 (N_1561,In_4918,In_4587);
nor U1562 (N_1562,In_992,In_4008);
and U1563 (N_1563,In_1596,In_427);
nor U1564 (N_1564,In_1618,In_1744);
xnor U1565 (N_1565,In_2024,In_2524);
nand U1566 (N_1566,In_2663,In_4459);
nor U1567 (N_1567,In_3030,In_4641);
xnor U1568 (N_1568,In_4356,In_3136);
and U1569 (N_1569,In_1212,In_1157);
or U1570 (N_1570,In_3029,In_2152);
nand U1571 (N_1571,In_4204,In_3380);
or U1572 (N_1572,In_1462,In_4571);
and U1573 (N_1573,In_3652,In_4897);
nor U1574 (N_1574,In_3906,In_4120);
and U1575 (N_1575,In_3124,In_2702);
nor U1576 (N_1576,In_4726,In_2329);
and U1577 (N_1577,In_4443,In_3992);
xor U1578 (N_1578,In_4821,In_2542);
xor U1579 (N_1579,In_4156,In_171);
nand U1580 (N_1580,In_4077,In_2281);
and U1581 (N_1581,In_1659,In_2961);
nand U1582 (N_1582,In_2995,In_3451);
xor U1583 (N_1583,In_1365,In_4518);
nand U1584 (N_1584,In_3539,In_2751);
or U1585 (N_1585,In_3108,In_3068);
and U1586 (N_1586,In_1428,In_3089);
and U1587 (N_1587,In_3722,In_2032);
nor U1588 (N_1588,In_2884,In_2157);
xnor U1589 (N_1589,In_4959,In_1598);
nor U1590 (N_1590,In_1383,In_2892);
or U1591 (N_1591,In_3486,In_352);
nor U1592 (N_1592,In_3105,In_2);
nand U1593 (N_1593,In_2660,In_3204);
or U1594 (N_1594,In_4200,In_2253);
and U1595 (N_1595,In_920,In_4025);
nand U1596 (N_1596,In_3276,In_2499);
nand U1597 (N_1597,In_2470,In_2920);
or U1598 (N_1598,In_23,In_4873);
xor U1599 (N_1599,In_1255,In_3024);
nor U1600 (N_1600,In_4600,In_2185);
xor U1601 (N_1601,In_2254,In_522);
or U1602 (N_1602,In_283,In_4080);
nor U1603 (N_1603,In_2106,In_737);
or U1604 (N_1604,In_887,In_3825);
or U1605 (N_1605,In_2848,In_1723);
xnor U1606 (N_1606,In_1886,In_3273);
nor U1607 (N_1607,In_1415,In_1101);
nand U1608 (N_1608,In_744,In_4212);
nor U1609 (N_1609,In_2552,In_2979);
nand U1610 (N_1610,In_1388,In_3560);
nor U1611 (N_1611,In_2200,In_2929);
nor U1612 (N_1612,In_2060,In_3293);
nor U1613 (N_1613,In_1304,In_3040);
and U1614 (N_1614,In_2998,In_2158);
nand U1615 (N_1615,In_4732,In_2601);
and U1616 (N_1616,In_1280,In_942);
nor U1617 (N_1617,In_2655,In_883);
xor U1618 (N_1618,In_739,In_3118);
or U1619 (N_1619,In_201,In_4738);
and U1620 (N_1620,In_1326,In_3773);
xnor U1621 (N_1621,In_1590,In_3559);
nor U1622 (N_1622,In_2795,In_340);
nor U1623 (N_1623,In_1238,In_2266);
nor U1624 (N_1624,In_3717,In_2134);
nand U1625 (N_1625,In_4503,In_4371);
nand U1626 (N_1626,In_4489,In_1360);
or U1627 (N_1627,In_68,In_697);
xnor U1628 (N_1628,In_3705,In_2583);
and U1629 (N_1629,In_4424,In_4216);
xnor U1630 (N_1630,In_4281,In_3857);
xor U1631 (N_1631,In_3310,In_2689);
nand U1632 (N_1632,In_4416,In_3096);
or U1633 (N_1633,In_1433,In_2963);
nor U1634 (N_1634,In_3382,In_1826);
and U1635 (N_1635,In_408,In_1636);
or U1636 (N_1636,In_2767,In_2530);
xor U1637 (N_1637,In_300,In_4553);
nand U1638 (N_1638,In_4441,In_151);
xnor U1639 (N_1639,In_3585,In_4935);
xnor U1640 (N_1640,In_2864,In_1134);
and U1641 (N_1641,In_3008,In_655);
xnor U1642 (N_1642,In_4189,In_1312);
nor U1643 (N_1643,In_3441,In_407);
or U1644 (N_1644,In_2068,In_459);
and U1645 (N_1645,In_2800,In_2323);
nand U1646 (N_1646,In_4318,In_2586);
and U1647 (N_1647,In_3845,In_4593);
nor U1648 (N_1648,In_2986,In_1993);
and U1649 (N_1649,In_381,In_4364);
nor U1650 (N_1650,In_3723,In_3851);
or U1651 (N_1651,In_925,In_4289);
nand U1652 (N_1652,In_3998,In_4904);
nor U1653 (N_1653,In_2447,In_4481);
nand U1654 (N_1654,In_197,In_75);
xnor U1655 (N_1655,In_590,In_2308);
or U1656 (N_1656,In_97,In_16);
and U1657 (N_1657,In_1103,In_2669);
xnor U1658 (N_1658,In_3544,In_4215);
or U1659 (N_1659,In_2613,In_1413);
and U1660 (N_1660,In_683,In_3954);
or U1661 (N_1661,In_586,In_2607);
or U1662 (N_1662,In_4407,In_919);
nand U1663 (N_1663,In_2584,In_4090);
and U1664 (N_1664,In_526,In_2906);
nor U1665 (N_1665,In_4562,In_305);
or U1666 (N_1666,In_343,In_1321);
or U1667 (N_1667,In_2082,In_1778);
nor U1668 (N_1668,In_230,In_931);
nor U1669 (N_1669,In_3231,In_4358);
nor U1670 (N_1670,In_1013,In_3810);
xor U1671 (N_1671,In_2036,In_3459);
xor U1672 (N_1672,In_1485,In_1809);
xnor U1673 (N_1673,In_1391,In_3225);
nor U1674 (N_1674,In_2110,In_600);
nor U1675 (N_1675,In_3111,In_867);
or U1676 (N_1676,In_4703,In_3419);
nor U1677 (N_1677,In_3075,In_4209);
nor U1678 (N_1678,In_2566,In_1692);
xnor U1679 (N_1679,In_1710,In_4382);
xor U1680 (N_1680,In_4742,In_4290);
and U1681 (N_1681,In_4242,In_4528);
nor U1682 (N_1682,In_3420,In_4608);
nand U1683 (N_1683,In_4804,In_4172);
xnor U1684 (N_1684,In_2822,In_3945);
xor U1685 (N_1685,In_2818,In_3942);
nand U1686 (N_1686,In_2237,In_3554);
nor U1687 (N_1687,In_3395,In_2571);
and U1688 (N_1688,In_989,In_3045);
xnor U1689 (N_1689,In_1655,In_3042);
nor U1690 (N_1690,In_1233,In_2465);
or U1691 (N_1691,In_1942,In_4754);
nor U1692 (N_1692,In_82,In_4283);
nor U1693 (N_1693,In_4544,In_246);
xor U1694 (N_1694,In_3347,In_354);
nor U1695 (N_1695,In_3683,In_44);
nor U1696 (N_1696,In_3052,In_60);
xor U1697 (N_1697,In_445,In_2568);
nor U1698 (N_1698,In_4994,In_1954);
and U1699 (N_1699,In_861,In_3552);
or U1700 (N_1700,In_3626,In_1057);
and U1701 (N_1701,In_4357,In_2980);
nand U1702 (N_1702,In_1248,In_1758);
xnor U1703 (N_1703,In_1322,In_1408);
nand U1704 (N_1704,In_4207,In_2493);
xnor U1705 (N_1705,In_2046,In_3327);
or U1706 (N_1706,In_1043,In_1235);
and U1707 (N_1707,In_2960,In_1897);
or U1708 (N_1708,In_3591,In_4079);
xnor U1709 (N_1709,In_2124,In_318);
and U1710 (N_1710,In_4061,In_4498);
xnor U1711 (N_1711,In_4987,In_1446);
nand U1712 (N_1712,In_1005,In_2626);
or U1713 (N_1713,In_1241,In_1364);
nand U1714 (N_1714,In_3445,In_3930);
and U1715 (N_1715,In_220,In_4928);
nor U1716 (N_1716,In_2636,In_567);
or U1717 (N_1717,In_4975,In_4255);
and U1718 (N_1718,In_3418,In_2858);
nor U1719 (N_1719,In_2511,In_2303);
nor U1720 (N_1720,In_3077,In_802);
and U1721 (N_1721,In_3318,In_3561);
xor U1722 (N_1722,In_2508,In_3733);
xnor U1723 (N_1723,In_686,In_2827);
and U1724 (N_1724,In_1502,In_1731);
and U1725 (N_1725,In_707,In_675);
nor U1726 (N_1726,In_2921,In_228);
and U1727 (N_1727,In_4907,In_494);
and U1728 (N_1728,In_3406,In_4325);
and U1729 (N_1729,In_622,In_3533);
and U1730 (N_1730,In_2179,In_4144);
nand U1731 (N_1731,In_4168,In_1270);
nand U1732 (N_1732,In_4111,In_4405);
xor U1733 (N_1733,In_4194,In_2826);
nor U1734 (N_1734,In_3383,In_1937);
xnor U1735 (N_1735,In_1010,In_2242);
and U1736 (N_1736,In_1056,In_3613);
nand U1737 (N_1737,In_190,In_3258);
or U1738 (N_1738,In_1017,In_4124);
nand U1739 (N_1739,In_1263,In_3866);
xor U1740 (N_1740,In_3496,In_4508);
nor U1741 (N_1741,In_185,In_2405);
nor U1742 (N_1742,In_2209,In_3675);
or U1743 (N_1743,In_1354,In_2399);
nor U1744 (N_1744,In_1542,In_3715);
nand U1745 (N_1745,In_4397,In_2457);
nand U1746 (N_1746,In_3871,In_4619);
xnor U1747 (N_1747,In_3300,In_534);
xor U1748 (N_1748,In_2642,In_3174);
and U1749 (N_1749,In_3622,In_61);
nor U1750 (N_1750,In_2076,In_2703);
and U1751 (N_1751,In_4983,In_3746);
nand U1752 (N_1752,In_2160,In_1066);
nand U1753 (N_1753,In_788,In_520);
xnor U1754 (N_1754,In_4003,In_2404);
nor U1755 (N_1755,In_2153,In_4106);
nor U1756 (N_1756,In_2841,In_430);
or U1757 (N_1757,In_101,In_1779);
nor U1758 (N_1758,In_4337,In_1240);
or U1759 (N_1759,In_1426,In_141);
nor U1760 (N_1760,In_2836,In_4515);
or U1761 (N_1761,In_657,In_928);
nor U1762 (N_1762,In_3602,In_3601);
and U1763 (N_1763,In_4385,In_4313);
nand U1764 (N_1764,In_1264,In_2363);
or U1765 (N_1765,In_415,In_2193);
xor U1766 (N_1766,In_826,In_440);
and U1767 (N_1767,In_3994,In_705);
xnor U1768 (N_1768,In_1336,In_4823);
and U1769 (N_1769,In_2498,In_2488);
nor U1770 (N_1770,In_2877,In_2713);
nand U1771 (N_1771,In_2992,In_2885);
and U1772 (N_1772,In_4040,In_434);
xor U1773 (N_1773,In_976,In_2162);
or U1774 (N_1774,In_2263,In_1007);
nand U1775 (N_1775,In_454,In_216);
xor U1776 (N_1776,In_1319,In_4708);
nor U1777 (N_1777,In_1921,In_2639);
nand U1778 (N_1778,In_3932,In_1126);
nor U1779 (N_1779,In_4750,In_3757);
or U1780 (N_1780,In_699,In_3251);
nand U1781 (N_1781,In_2131,In_4963);
xnor U1782 (N_1782,In_3000,In_389);
xnor U1783 (N_1783,In_3275,In_3100);
and U1784 (N_1784,In_4752,In_4307);
xnor U1785 (N_1785,In_2235,In_2025);
xnor U1786 (N_1786,In_1683,In_3391);
or U1787 (N_1787,In_517,In_3055);
and U1788 (N_1788,In_589,In_2230);
nor U1789 (N_1789,In_2862,In_1442);
nor U1790 (N_1790,In_3587,In_360);
and U1791 (N_1791,In_1960,In_746);
and U1792 (N_1792,In_2515,In_2420);
nor U1793 (N_1793,In_4950,In_718);
nor U1794 (N_1794,In_2324,In_1962);
and U1795 (N_1795,In_980,In_3478);
nand U1796 (N_1796,In_3838,In_1403);
nor U1797 (N_1797,In_1653,In_71);
nand U1798 (N_1798,In_4268,In_1907);
and U1799 (N_1799,In_3217,In_2762);
or U1800 (N_1800,In_4467,In_4781);
nor U1801 (N_1801,In_3823,In_2245);
xnor U1802 (N_1802,In_2895,In_2484);
and U1803 (N_1803,In_2558,In_1529);
xnor U1804 (N_1804,In_13,In_724);
and U1805 (N_1805,In_4065,In_4893);
or U1806 (N_1806,In_1994,In_2495);
xor U1807 (N_1807,In_3067,In_2016);
nor U1808 (N_1808,In_1223,In_4004);
and U1809 (N_1809,In_1511,In_3978);
or U1810 (N_1810,In_2619,In_4954);
nor U1811 (N_1811,In_2602,In_2934);
xnor U1812 (N_1812,In_1878,In_1481);
nor U1813 (N_1813,In_2690,In_3792);
or U1814 (N_1814,In_4866,In_3412);
nor U1815 (N_1815,In_2229,In_4691);
nor U1816 (N_1816,In_2436,In_4135);
or U1817 (N_1817,In_294,In_3824);
and U1818 (N_1818,In_2004,In_1836);
nand U1819 (N_1819,In_591,In_3093);
xnor U1820 (N_1820,In_2426,In_1841);
nor U1821 (N_1821,In_4465,In_2759);
and U1822 (N_1822,In_2095,In_4927);
or U1823 (N_1823,In_1535,In_1862);
nand U1824 (N_1824,In_911,In_3762);
or U1825 (N_1825,In_252,In_3425);
or U1826 (N_1826,In_441,In_1648);
and U1827 (N_1827,In_4717,In_4222);
xnor U1828 (N_1828,In_4399,In_3710);
nand U1829 (N_1829,In_1679,In_1733);
and U1830 (N_1830,In_489,In_990);
or U1831 (N_1831,In_2321,In_487);
and U1832 (N_1832,In_547,In_2361);
xnor U1833 (N_1833,In_309,In_1741);
xor U1834 (N_1834,In_4825,In_3861);
and U1835 (N_1835,In_587,In_2198);
or U1836 (N_1836,In_4899,In_3267);
nor U1837 (N_1837,In_3646,In_3685);
nor U1838 (N_1838,In_688,In_3782);
nor U1839 (N_1839,In_266,In_3577);
and U1840 (N_1840,In_3750,In_4786);
or U1841 (N_1841,In_2118,In_3455);
nand U1842 (N_1842,In_3352,In_49);
nand U1843 (N_1843,In_391,In_403);
xor U1844 (N_1844,In_2644,In_1986);
or U1845 (N_1845,In_1395,In_4123);
and U1846 (N_1846,In_3365,In_3818);
xor U1847 (N_1847,In_760,In_107);
or U1848 (N_1848,In_888,In_2555);
xnor U1849 (N_1849,In_1782,In_2286);
and U1850 (N_1850,In_2313,In_4583);
xnor U1851 (N_1851,In_4091,In_3919);
xnor U1852 (N_1852,In_1296,In_2549);
and U1853 (N_1853,In_1339,In_805);
nor U1854 (N_1854,In_127,In_694);
nor U1855 (N_1855,In_3434,In_3464);
xnor U1856 (N_1856,In_3328,In_2010);
nor U1857 (N_1857,In_3868,In_3958);
xnor U1858 (N_1858,In_3771,In_4333);
nor U1859 (N_1859,In_933,In_4972);
nor U1860 (N_1860,In_4942,In_3288);
nand U1861 (N_1861,In_1512,In_605);
nor U1862 (N_1862,In_91,In_2632);
or U1863 (N_1863,In_369,In_4023);
nor U1864 (N_1864,In_3599,In_1156);
nand U1865 (N_1865,In_2900,In_2272);
nand U1866 (N_1866,In_4294,In_2136);
or U1867 (N_1867,In_2364,In_4063);
nand U1868 (N_1868,In_2540,In_1971);
nor U1869 (N_1869,In_36,In_2410);
xnor U1870 (N_1870,In_3311,In_1492);
nand U1871 (N_1871,In_2728,In_2128);
nand U1872 (N_1872,In_1091,In_368);
nor U1873 (N_1873,In_4066,In_2623);
nor U1874 (N_1874,In_4525,In_4097);
nor U1875 (N_1875,In_4070,In_3129);
nand U1876 (N_1876,In_3442,In_4042);
xnor U1877 (N_1877,In_1517,In_400);
nor U1878 (N_1878,In_4605,In_1950);
nand U1879 (N_1879,In_1044,In_3320);
and U1880 (N_1880,In_1766,In_491);
nand U1881 (N_1881,In_358,In_3296);
and U1882 (N_1882,In_3870,In_2816);
nand U1883 (N_1883,In_1310,In_1793);
nor U1884 (N_1884,In_3921,In_3826);
nand U1885 (N_1885,In_797,In_3925);
nand U1886 (N_1886,In_1436,In_3853);
nand U1887 (N_1887,In_2219,In_2823);
and U1888 (N_1888,In_1106,In_2709);
or U1889 (N_1889,In_676,In_2863);
nor U1890 (N_1890,In_100,In_399);
or U1891 (N_1891,In_2268,In_4919);
nor U1892 (N_1892,In_1175,In_2206);
and U1893 (N_1893,In_496,In_4470);
xnor U1894 (N_1894,In_3662,In_280);
and U1895 (N_1895,In_442,In_120);
or U1896 (N_1896,In_3501,In_764);
xnor U1897 (N_1897,In_3013,In_2343);
nand U1898 (N_1898,In_1895,In_2146);
nand U1899 (N_1899,In_629,In_609);
and U1900 (N_1900,In_704,In_2791);
nand U1901 (N_1901,In_3155,In_2726);
nand U1902 (N_1902,In_4668,In_2945);
and U1903 (N_1903,In_1536,In_24);
xor U1904 (N_1904,In_776,In_2239);
nor U1905 (N_1905,In_3584,In_3799);
nand U1906 (N_1906,In_483,In_2516);
nand U1907 (N_1907,In_1694,In_1071);
nand U1908 (N_1908,In_1952,In_2727);
nor U1909 (N_1909,In_4723,In_2758);
and U1910 (N_1910,In_3367,In_1171);
nand U1911 (N_1911,In_3889,In_506);
nand U1912 (N_1912,In_2637,In_1750);
xor U1913 (N_1913,In_3497,In_1224);
nor U1914 (N_1914,In_1281,In_4001);
nand U1915 (N_1915,In_2192,In_3398);
nor U1916 (N_1916,In_3149,In_2228);
nor U1917 (N_1917,In_1761,In_1159);
or U1918 (N_1918,In_2057,In_1026);
and U1919 (N_1919,In_4985,In_2935);
nor U1920 (N_1920,In_3241,In_2652);
nor U1921 (N_1921,In_213,In_18);
nor U1922 (N_1922,In_2119,In_1412);
nand U1923 (N_1923,In_3852,In_3862);
nand U1924 (N_1924,In_4707,In_4779);
nor U1925 (N_1925,In_4327,In_179);
or U1926 (N_1926,In_940,In_2638);
nand U1927 (N_1927,In_163,In_3586);
nand U1928 (N_1928,In_4406,In_3957);
and U1929 (N_1929,In_2874,In_2494);
xnor U1930 (N_1930,In_2994,In_1314);
nand U1931 (N_1931,In_2962,In_4594);
or U1932 (N_1932,In_4116,In_4602);
xnor U1933 (N_1933,In_2386,In_1797);
xor U1934 (N_1934,In_664,In_853);
or U1935 (N_1935,In_3351,In_4782);
nand U1936 (N_1936,In_3885,In_2668);
xnor U1937 (N_1937,In_2284,In_1313);
nor U1938 (N_1938,In_1196,In_245);
and U1939 (N_1939,In_1231,In_287);
nand U1940 (N_1940,In_3325,In_3654);
and U1941 (N_1941,In_696,In_2290);
or U1942 (N_1942,In_3639,In_3667);
nor U1943 (N_1943,In_2971,In_1167);
nor U1944 (N_1944,In_874,In_3684);
nor U1945 (N_1945,In_314,In_3619);
nor U1946 (N_1946,In_3527,In_1060);
or U1947 (N_1947,In_4068,In_15);
nand U1948 (N_1948,In_562,In_189);
nand U1949 (N_1949,In_1704,In_469);
and U1950 (N_1950,In_2231,In_1620);
nand U1951 (N_1951,In_1968,In_2949);
nand U1952 (N_1952,In_4616,In_4293);
nand U1953 (N_1953,In_3843,In_2107);
xor U1954 (N_1954,In_1668,In_3844);
nor U1955 (N_1955,In_3377,In_1379);
nand U1956 (N_1956,In_431,In_3041);
and U1957 (N_1957,In_3720,In_2320);
and U1958 (N_1958,In_1163,In_263);
or U1959 (N_1959,In_4764,In_3643);
nand U1960 (N_1960,In_3739,In_270);
or U1961 (N_1961,In_1021,In_418);
and U1962 (N_1962,In_2126,In_1204);
nor U1963 (N_1963,In_4543,In_4715);
or U1964 (N_1964,In_3173,In_3230);
nand U1965 (N_1965,In_4868,In_181);
nand U1966 (N_1966,In_4287,In_834);
or U1967 (N_1967,In_1586,In_1531);
nand U1968 (N_1968,In_1807,In_4622);
xor U1969 (N_1969,In_375,In_446);
or U1970 (N_1970,In_525,In_849);
or U1971 (N_1971,In_2710,In_3402);
nand U1972 (N_1972,In_687,In_118);
nor U1973 (N_1973,In_768,In_4472);
nor U1974 (N_1974,In_1421,In_3576);
nand U1975 (N_1975,In_3989,In_2067);
nor U1976 (N_1976,In_4234,In_1246);
xor U1977 (N_1977,In_4121,In_4086);
nand U1978 (N_1978,In_2094,In_4119);
nand U1979 (N_1979,In_1814,In_1637);
nand U1980 (N_1980,In_1,In_3579);
or U1981 (N_1981,In_4316,In_2970);
nor U1982 (N_1982,In_2277,In_2406);
and U1983 (N_1983,In_458,In_3509);
nor U1984 (N_1984,In_4050,In_4661);
or U1985 (N_1985,In_624,In_3678);
or U1986 (N_1986,In_1927,In_1613);
and U1987 (N_1987,In_1837,In_2723);
nand U1988 (N_1988,In_2441,In_3170);
nor U1989 (N_1989,In_3765,In_2197);
and U1990 (N_1990,In_1093,In_3803);
xnor U1991 (N_1991,In_3948,In_1781);
nand U1992 (N_1992,In_4800,In_2210);
and U1993 (N_1993,In_1454,In_4225);
and U1994 (N_1994,In_251,In_2241);
or U1995 (N_1995,In_2705,In_1366);
xnor U1996 (N_1996,In_2879,In_451);
nand U1997 (N_1997,In_2341,In_4988);
xor U1998 (N_1998,In_2145,In_1901);
or U1999 (N_1999,In_2437,In_4648);
or U2000 (N_2000,In_4552,In_833);
xor U2001 (N_2001,In_3607,In_2941);
nor U2002 (N_2002,In_4838,In_1788);
xor U2003 (N_2003,In_4900,In_1522);
xor U2004 (N_2004,In_2443,In_4669);
nor U2005 (N_2005,In_1300,In_3634);
or U2006 (N_2006,In_4181,In_2630);
or U2007 (N_2007,In_1190,In_4895);
or U2008 (N_2008,In_3666,In_2631);
xor U2009 (N_2009,In_885,In_37);
nand U2010 (N_2010,In_4862,In_456);
xnor U2011 (N_2011,In_4478,In_2505);
or U2012 (N_2012,In_4248,In_2001);
nor U2013 (N_2013,In_3182,In_2489);
nor U2014 (N_2014,In_3342,In_3485);
nand U2015 (N_2015,In_1752,In_3783);
nor U2016 (N_2016,In_3528,In_3148);
xnor U2017 (N_2017,In_2215,In_4549);
xnor U2018 (N_2018,In_3424,In_4607);
nor U2019 (N_2019,In_253,In_2143);
or U2020 (N_2020,In_1422,In_4609);
or U2021 (N_2021,In_2159,In_4926);
nand U2022 (N_2022,In_3672,In_9);
and U2023 (N_2023,In_1198,In_2088);
nor U2024 (N_2024,In_79,In_143);
nand U2025 (N_2025,In_1118,In_4457);
and U2026 (N_2026,In_365,In_1584);
or U2027 (N_2027,In_4526,In_1154);
or U2028 (N_2028,In_1376,In_1030);
xnor U2029 (N_2029,In_574,In_1725);
xnor U2030 (N_2030,In_4507,In_4831);
nand U2031 (N_2031,In_2285,In_218);
and U2032 (N_2032,In_1441,In_2964);
and U2033 (N_2033,In_2525,In_4799);
nand U2034 (N_2034,In_2390,In_3956);
nor U2035 (N_2035,In_4154,In_749);
or U2036 (N_2036,In_2243,In_3283);
or U2037 (N_2037,In_3062,In_884);
nand U2038 (N_2038,In_4329,In_1434);
nor U2039 (N_2039,In_3781,In_1680);
or U2040 (N_2040,In_1875,In_2066);
or U2041 (N_2041,In_232,In_64);
or U2042 (N_2042,In_3701,In_3086);
xnor U2043 (N_2043,In_2339,In_1065);
nand U2044 (N_2044,In_1425,In_438);
nand U2045 (N_2045,In_4109,In_3758);
xnor U2046 (N_2046,In_1269,In_2577);
nand U2047 (N_2047,In_859,In_612);
and U2048 (N_2048,In_1439,In_1773);
and U2049 (N_2049,In_2047,In_95);
nor U2050 (N_2050,In_3976,In_1328);
nor U2051 (N_2051,In_1885,In_1753);
nand U2052 (N_2052,In_27,In_3549);
and U2053 (N_2053,In_349,In_3985);
xor U2054 (N_2054,In_2946,In_1858);
xnor U2055 (N_2055,In_132,In_2064);
nor U2056 (N_2056,In_3429,In_986);
xnor U2057 (N_2057,In_4791,In_4887);
and U2058 (N_2058,In_3663,In_593);
or U2059 (N_2059,In_174,In_4687);
nand U2060 (N_2060,In_363,In_721);
or U2061 (N_2061,In_2618,In_383);
or U2062 (N_2062,In_497,In_1828);
xor U2063 (N_2063,In_634,In_28);
and U2064 (N_2064,In_4635,In_745);
or U2065 (N_2065,In_4021,In_1691);
xnor U2066 (N_2066,In_1787,In_1048);
xor U2067 (N_2067,In_3794,In_4582);
xor U2068 (N_2068,In_4657,In_2260);
nand U2069 (N_2069,In_2061,In_482);
nor U2070 (N_2070,In_4945,In_3708);
nand U2071 (N_2071,In_4506,In_4855);
nand U2072 (N_2072,In_390,In_52);
and U2073 (N_2073,In_1693,In_757);
and U2074 (N_2074,In_2526,In_4380);
xnor U2075 (N_2075,In_7,In_3002);
nand U2076 (N_2076,In_1995,In_748);
or U2077 (N_2077,In_4227,In_3918);
xor U2078 (N_2078,In_839,In_1023);
nand U2079 (N_2079,In_4469,In_1540);
nand U2080 (N_2080,In_1642,In_4947);
xnor U2081 (N_2081,In_2366,In_484);
and U2082 (N_2082,In_410,In_4701);
or U2083 (N_2083,In_1765,In_564);
xnor U2084 (N_2084,In_2987,In_3649);
nand U2085 (N_2085,In_1031,In_4340);
nand U2086 (N_2086,In_4628,In_1533);
and U2087 (N_2087,In_3213,In_1764);
or U2088 (N_2088,In_2893,In_2473);
or U2089 (N_2089,In_1720,In_4252);
nor U2090 (N_2090,In_1177,In_3345);
nand U2091 (N_2091,In_3713,In_3457);
xnor U2092 (N_2092,In_4851,In_3547);
and U2093 (N_2093,In_2766,In_225);
and U2094 (N_2094,In_964,In_829);
or U2095 (N_2095,In_549,In_3540);
or U2096 (N_2096,In_2535,In_285);
or U2097 (N_2097,In_4643,In_4286);
nand U2098 (N_2098,In_2020,In_2120);
and U2099 (N_2099,In_1493,In_4733);
or U2100 (N_2100,In_3571,In_4666);
or U2101 (N_2101,In_2000,In_3827);
nand U2102 (N_2102,In_903,In_836);
nand U2103 (N_2103,In_2545,In_1798);
and U2104 (N_2104,In_1149,In_1012);
and U2105 (N_2105,In_4292,In_2425);
xor U2106 (N_2106,In_974,In_2679);
or U2107 (N_2107,In_3689,In_1534);
nand U2108 (N_2108,In_2448,In_870);
nor U2109 (N_2109,In_3284,In_2070);
nor U2110 (N_2110,In_4291,In_4187);
xor U2111 (N_2111,In_3034,In_2434);
or U2112 (N_2112,In_1866,In_3152);
nor U2113 (N_2113,In_3421,In_4464);
nor U2114 (N_2114,In_1197,In_817);
nor U2115 (N_2115,In_1996,In_3735);
and U2116 (N_2116,In_1612,In_945);
and U2117 (N_2117,In_2954,In_2927);
nor U2118 (N_2118,In_1650,In_162);
or U2119 (N_2119,In_1913,In_719);
or U2120 (N_2120,In_509,In_4599);
xor U2121 (N_2121,In_4968,In_3892);
nand U2122 (N_2122,In_1509,In_3681);
and U2123 (N_2123,In_3027,In_2743);
and U2124 (N_2124,In_550,In_3606);
nor U2125 (N_2125,In_1633,In_2853);
xor U2126 (N_2126,In_4493,In_659);
and U2127 (N_2127,In_182,In_1894);
xor U2128 (N_2128,In_3176,In_2605);
xnor U2129 (N_2129,In_1329,In_4700);
or U2130 (N_2130,In_2091,In_3044);
xnor U2131 (N_2131,In_1805,In_4418);
and U2132 (N_2132,In_2736,In_1974);
xnor U2133 (N_2133,In_3332,In_3242);
xor U2134 (N_2134,In_4581,In_133);
nand U2135 (N_2135,In_3349,In_1567);
nor U2136 (N_2136,In_3126,In_514);
or U2137 (N_2137,In_1706,In_1045);
nand U2138 (N_2138,In_1096,In_2449);
or U2139 (N_2139,In_773,In_353);
nor U2140 (N_2140,In_4437,In_3744);
and U2141 (N_2141,In_580,In_2418);
nand U2142 (N_2142,In_3730,In_4496);
nor U2143 (N_2143,In_4787,In_3481);
and U2144 (N_2144,In_832,In_4801);
xnor U2145 (N_2145,In_2274,In_2861);
and U2146 (N_2146,In_2755,In_4160);
nor U2147 (N_2147,In_983,In_1349);
and U2148 (N_2148,In_4439,In_2238);
and U2149 (N_2149,In_4929,In_3894);
xnor U2150 (N_2150,In_3198,In_1487);
and U2151 (N_2151,In_2462,In_3519);
and U2152 (N_2152,In_1452,In_1489);
nand U2153 (N_2153,In_1972,In_3356);
or U2154 (N_2154,In_4375,In_3686);
or U2155 (N_2155,In_3553,In_1851);
xor U2156 (N_2156,In_961,In_492);
or U2157 (N_2157,In_1912,In_2362);
or U2158 (N_2158,In_1124,In_3524);
nor U2159 (N_2159,In_1076,In_3003);
nor U2160 (N_2160,In_569,In_1432);
xor U2161 (N_2161,In_3023,In_4793);
nand U2162 (N_2162,In_3763,In_3761);
or U2163 (N_2163,In_1898,In_3724);
nand U2164 (N_2164,In_3362,In_2213);
nand U2165 (N_2165,In_4020,In_2739);
and U2166 (N_2166,In_4435,In_752);
nor U2167 (N_2167,In_3743,In_2780);
and U2168 (N_2168,In_2711,In_2077);
and U2169 (N_2169,In_3085,In_1396);
xnor U2170 (N_2170,In_1411,In_4027);
xor U2171 (N_2171,In_2415,In_3535);
or U2172 (N_2172,In_528,In_373);
xnor U2173 (N_2173,In_4686,In_2065);
nand U2174 (N_2174,In_4262,In_2302);
nor U2175 (N_2175,In_3742,In_4019);
nand U2176 (N_2176,In_1576,In_106);
and U2177 (N_2177,In_2365,In_3569);
nor U2178 (N_2178,In_971,In_2561);
xor U2179 (N_2179,In_3361,In_4556);
nor U2180 (N_2180,In_1128,In_715);
nor U2181 (N_2181,In_4902,In_4404);
and U2182 (N_2182,In_2976,In_3854);
nand U2183 (N_2183,In_1903,In_4634);
and U2184 (N_2184,In_2227,In_4783);
nor U2185 (N_2185,In_2038,In_1812);
nor U2186 (N_2186,In_4861,In_2592);
xor U2187 (N_2187,In_1496,In_3354);
nor U2188 (N_2188,In_4695,In_2257);
and U2189 (N_2189,In_789,In_279);
nor U2190 (N_2190,In_561,In_2562);
xor U2191 (N_2191,In_4173,In_4991);
xor U2192 (N_2192,In_261,In_2977);
and U2193 (N_2193,In_2694,In_4637);
and U2194 (N_2194,In_669,In_307);
xor U2195 (N_2195,In_77,In_3274);
and U2196 (N_2196,In_4674,In_1887);
nor U2197 (N_2197,In_156,In_1526);
and U2198 (N_2198,In_3828,In_1081);
xnor U2199 (N_2199,In_2188,In_4636);
and U2200 (N_2200,In_476,In_256);
or U2201 (N_2201,In_17,In_2017);
and U2202 (N_2202,In_2930,In_3254);
and U2203 (N_2203,In_4775,In_2916);
or U2204 (N_2204,In_729,In_2804);
xnor U2205 (N_2205,In_477,In_3151);
nand U2206 (N_2206,In_3908,In_129);
nor U2207 (N_2207,In_2835,In_4428);
or U2208 (N_2208,In_2384,In_1459);
and U2209 (N_2209,In_4153,In_3164);
nor U2210 (N_2210,In_2931,In_846);
nor U2211 (N_2211,In_626,In_793);
nand U2212 (N_2212,In_1342,In_1763);
or U2213 (N_2213,In_1829,In_3951);
and U2214 (N_2214,In_3121,In_3321);
nor U2215 (N_2215,In_4925,In_4685);
and U2216 (N_2216,In_807,In_4193);
or U2217 (N_2217,In_1052,In_3433);
nand U2218 (N_2218,In_4720,In_2857);
xnor U2219 (N_2219,In_4992,In_1624);
xor U2220 (N_2220,In_3202,In_94);
or U2221 (N_2221,In_260,In_32);
nand U2222 (N_2222,In_1520,In_191);
nand U2223 (N_2223,In_4183,In_4417);
nor U2224 (N_2224,In_4266,In_3784);
nor U2225 (N_2225,In_917,In_2338);
xor U2226 (N_2226,In_4057,In_312);
or U2227 (N_2227,In_1860,In_886);
nor U2228 (N_2228,In_215,In_1842);
xnor U2229 (N_2229,In_3414,In_1419);
xor U2230 (N_2230,In_2370,In_1834);
or U2231 (N_2231,In_1629,In_2670);
nor U2232 (N_2232,In_1749,In_3836);
nand U2233 (N_2233,In_3025,In_4978);
or U2234 (N_2234,In_1803,In_3548);
and U2235 (N_2235,In_1714,In_161);
xnor U2236 (N_2236,In_432,In_1343);
nor U2237 (N_2237,In_472,In_3200);
nor U2238 (N_2238,In_2947,In_3816);
or U2239 (N_2239,In_3754,In_316);
and U2240 (N_2240,In_2389,In_113);
xor U2241 (N_2241,In_2204,In_3572);
nand U2242 (N_2242,In_3350,In_4545);
nand U2243 (N_2243,In_3107,In_1059);
or U2244 (N_2244,In_4853,In_3551);
nor U2245 (N_2245,In_530,In_871);
nand U2246 (N_2246,In_165,In_1755);
nor U2247 (N_2247,In_2002,In_3936);
and U2248 (N_2248,In_1527,In_3711);
nand U2249 (N_2249,In_89,In_1997);
nor U2250 (N_2250,In_4796,In_1341);
nand U2251 (N_2251,In_585,In_308);
or U2252 (N_2252,In_2222,In_1067);
xnor U2253 (N_2253,In_2043,In_4664);
xnor U2254 (N_2254,In_4150,In_4612);
xnor U2255 (N_2255,In_4973,In_2813);
nor U2256 (N_2256,In_2334,In_3405);
nor U2257 (N_2257,In_356,In_1003);
nand U2258 (N_2258,In_4132,In_645);
xor U2259 (N_2259,In_1119,In_3006);
or U2260 (N_2260,In_3460,In_4589);
and U2261 (N_2261,In_4342,In_3226);
or U2262 (N_2262,In_1409,In_2048);
nand U2263 (N_2263,In_4824,In_3297);
nand U2264 (N_2264,In_4341,In_2491);
nor U2265 (N_2265,In_1221,In_3266);
or U2266 (N_2266,In_2481,In_2950);
and U2267 (N_2267,In_1476,In_1380);
and U2268 (N_2268,In_4140,In_4557);
or U2269 (N_2269,In_3139,In_1033);
and U2270 (N_2270,In_868,In_2828);
xnor U2271 (N_2271,In_3647,In_4885);
nor U2272 (N_2272,In_3299,In_723);
and U2273 (N_2273,In_195,In_1569);
or U2274 (N_2274,In_1746,In_4759);
and U2275 (N_2275,In_3714,In_623);
and U2276 (N_2276,In_3725,In_3620);
or U2277 (N_2277,In_924,In_4704);
or U2278 (N_2278,In_114,In_135);
xnor U2279 (N_2279,In_419,In_41);
or U2280 (N_2280,In_2730,In_4372);
or U2281 (N_2281,In_2051,In_949);
and U2282 (N_2282,In_4306,In_336);
or U2283 (N_2283,In_1136,In_2825);
or U2284 (N_2284,In_273,In_1172);
nor U2285 (N_2285,In_2942,In_3282);
nand U2286 (N_2286,In_1553,In_2843);
nor U2287 (N_2287,In_4495,In_1077);
or U2288 (N_2288,In_4101,In_4282);
or U2289 (N_2289,In_800,In_2037);
nor U2290 (N_2290,In_4826,In_4510);
xor U2291 (N_2291,In_2445,In_3207);
or U2292 (N_2292,In_2029,In_4471);
or U2293 (N_2293,In_1210,In_3642);
or U2294 (N_2294,In_2968,In_4084);
nand U2295 (N_2295,In_4134,In_2421);
and U2296 (N_2296,In_4280,In_3537);
and U2297 (N_2297,In_2534,In_1799);
and U2298 (N_2298,In_3161,In_2135);
and U2299 (N_2299,In_3706,In_1661);
nor U2300 (N_2300,In_3494,In_3106);
nand U2301 (N_2301,In_3312,In_3047);
nand U2302 (N_2302,In_3804,In_1472);
and U2303 (N_2303,In_4110,In_3186);
nor U2304 (N_2304,In_1964,In_1914);
or U2305 (N_2305,In_4617,In_1256);
and U2306 (N_2306,In_1666,In_2783);
or U2307 (N_2307,In_1036,In_3886);
xor U2308 (N_2308,In_342,In_2092);
and U2309 (N_2309,In_2724,In_844);
nor U2310 (N_2310,In_1361,In_229);
nor U2311 (N_2311,In_370,In_1371);
xor U2312 (N_2312,In_2582,In_1605);
and U2313 (N_2313,In_4440,In_726);
and U2314 (N_2314,In_3209,In_33);
nand U2315 (N_2315,In_1591,In_2754);
nor U2316 (N_2316,In_3929,In_3953);
and U2317 (N_2317,In_2298,In_1849);
xnor U2318 (N_2318,In_1332,In_4584);
xnor U2319 (N_2319,In_1037,In_4046);
or U2320 (N_2320,In_582,In_3079);
xnor U2321 (N_2321,In_2887,In_4538);
nor U2322 (N_2322,In_2234,In_4516);
nor U2323 (N_2323,In_4033,In_938);
and U2324 (N_2324,In_4007,In_3798);
nand U2325 (N_2325,In_2749,In_2910);
and U2326 (N_2326,In_3874,In_1721);
nand U2327 (N_2327,In_2353,In_3261);
xor U2328 (N_2328,In_3355,In_648);
nand U2329 (N_2329,In_4566,In_3403);
nor U2330 (N_2330,In_72,In_953);
nand U2331 (N_2331,In_4345,In_3618);
xnor U2332 (N_2332,In_2683,In_1909);
xor U2333 (N_2333,In_4370,In_4677);
or U2334 (N_2334,In_754,In_2490);
nand U2335 (N_2335,In_1020,In_1273);
nor U2336 (N_2336,In_4339,In_319);
nor U2337 (N_2337,In_2847,In_2764);
nor U2338 (N_2338,In_3128,In_1603);
xor U2339 (N_2339,In_2507,In_1053);
and U2340 (N_2340,In_1262,In_4059);
nor U2341 (N_2341,In_2073,In_631);
xnor U2342 (N_2342,In_2099,In_3665);
nor U2343 (N_2343,In_290,In_1120);
or U2344 (N_2344,In_819,In_3650);
nand U2345 (N_2345,In_3615,In_236);
nor U2346 (N_2346,In_4006,In_2750);
xor U2347 (N_2347,In_4434,In_4151);
and U2348 (N_2348,In_3378,In_1577);
and U2349 (N_2349,In_1625,In_2409);
and U2350 (N_2350,In_2594,In_4322);
and U2351 (N_2351,In_3834,In_421);
xnor U2352 (N_2352,In_927,In_184);
or U2353 (N_2353,In_4149,In_3965);
nand U2354 (N_2354,In_110,In_4125);
nor U2355 (N_2355,In_1195,In_4304);
or U2356 (N_2356,In_259,In_450);
or U2357 (N_2357,In_1545,In_3404);
and U2358 (N_2358,In_248,In_3917);
nand U2359 (N_2359,In_3224,In_2514);
nor U2360 (N_2360,In_188,In_982);
nor U2361 (N_2361,In_978,In_1146);
and U2362 (N_2362,In_2224,In_3138);
or U2363 (N_2363,In_1677,In_1498);
and U2364 (N_2364,In_2904,In_662);
or U2365 (N_2365,In_2714,In_4142);
nor U2366 (N_2366,In_4514,In_3212);
nor U2367 (N_2367,In_732,In_714);
or U2368 (N_2368,In_268,In_4789);
or U2369 (N_2369,In_2083,In_1307);
xnor U2370 (N_2370,In_2707,In_4870);
or U2371 (N_2371,In_3727,In_3020);
nor U2372 (N_2372,In_646,In_4343);
nand U2373 (N_2373,In_2951,In_1675);
or U2374 (N_2374,In_4303,In_3764);
and U2375 (N_2375,In_3287,In_2173);
nor U2376 (N_2376,In_1777,In_625);
xor U2377 (N_2377,In_176,In_2985);
nor U2378 (N_2378,In_1490,In_568);
xnor U2379 (N_2379,In_457,In_3363);
nand U2380 (N_2380,In_2903,In_3163);
nand U2381 (N_2381,In_1722,In_3796);
nor U2382 (N_2382,In_3914,In_4724);
or U2383 (N_2383,In_4965,In_3940);
and U2384 (N_2384,In_2541,In_910);
xor U2385 (N_2385,In_3819,In_2978);
nand U2386 (N_2386,In_4585,In_3060);
or U2387 (N_2387,In_500,In_3668);
nor U2388 (N_2388,In_1242,In_1776);
xnor U2389 (N_2389,In_1738,In_1276);
xor U2390 (N_2390,In_2596,In_1499);
nand U2391 (N_2391,In_537,In_4158);
xor U2392 (N_2392,In_3653,In_34);
nand U2393 (N_2393,In_1032,In_214);
or U2394 (N_2394,In_3839,In_3073);
or U2395 (N_2395,In_2889,In_1024);
xnor U2396 (N_2396,In_217,In_4118);
or U2397 (N_2397,In_966,In_4480);
nand U2398 (N_2398,In_3915,In_2325);
and U2399 (N_2399,In_2993,In_409);
and U2400 (N_2400,In_2429,In_2649);
nand U2401 (N_2401,In_3831,In_2007);
xnor U2402 (N_2402,In_1250,In_4688);
xnor U2403 (N_2403,In_4598,In_4522);
nor U2404 (N_2404,In_2335,In_3082);
nor U2405 (N_2405,In_3805,In_2988);
nor U2406 (N_2406,In_4741,In_2680);
and U2407 (N_2407,In_2528,In_3097);
nand U2408 (N_2408,In_1497,In_2590);
and U2409 (N_2409,In_1762,In_4709);
nand U2410 (N_2410,In_4081,In_2218);
xor U2411 (N_2411,In_842,In_1507);
nor U2412 (N_2412,In_1229,In_481);
nand U2413 (N_2413,In_4561,In_597);
or U2414 (N_2414,In_357,In_3688);
and U2415 (N_2415,In_4320,In_1508);
nor U2416 (N_2416,In_334,In_722);
and U2417 (N_2417,In_3779,In_3759);
xnor U2418 (N_2418,In_275,In_2504);
or U2419 (N_2419,In_599,In_137);
xnor U2420 (N_2420,In_3438,In_512);
nor U2421 (N_2421,In_3691,In_1064);
nor U2422 (N_2422,In_3303,In_1915);
xor U2423 (N_2423,In_2129,In_3181);
or U2424 (N_2424,In_1588,In_4756);
xnor U2425 (N_2425,In_814,In_2471);
nand U2426 (N_2426,In_4350,In_865);
and U2427 (N_2427,In_4574,In_4867);
nand U2428 (N_2428,In_3291,In_3177);
xnor U2429 (N_2429,In_4890,In_4438);
xnor U2430 (N_2430,In_4015,In_1084);
and U2431 (N_2431,In_1783,In_951);
xnor U2432 (N_2432,In_4202,In_153);
nor U2433 (N_2433,In_847,In_3947);
and U2434 (N_2434,In_1580,In_80);
and U2435 (N_2435,In_4328,In_3594);
xor U2436 (N_2436,In_4395,In_2972);
and U2437 (N_2437,In_271,In_3848);
xnor U2438 (N_2438,In_2178,In_462);
nor U2439 (N_2439,In_1372,In_864);
nor U2440 (N_2440,In_523,In_504);
or U2441 (N_2441,In_4513,In_2155);
nand U2442 (N_2442,In_1748,In_1042);
or U2443 (N_2443,In_3747,In_2778);
xor U2444 (N_2444,In_2840,In_2718);
xnor U2445 (N_2445,In_2248,In_47);
xnor U2446 (N_2446,In_3189,In_4654);
or U2447 (N_2447,In_1902,In_1333);
nor U2448 (N_2448,In_4776,In_4746);
and U2449 (N_2449,In_3338,In_621);
nor U2450 (N_2450,In_843,In_3493);
and U2451 (N_2451,In_2799,In_3719);
xor U2452 (N_2452,In_2295,In_1525);
or U2453 (N_2453,In_4820,In_2121);
xnor U2454 (N_2454,In_1259,In_610);
and U2455 (N_2455,In_3841,In_3270);
or U2456 (N_2456,In_10,In_2819);
nand U2457 (N_2457,In_255,In_1435);
and U2458 (N_2458,In_3538,In_2354);
or U2459 (N_2459,In_3898,In_387);
xor U2460 (N_2460,In_4198,In_291);
and U2461 (N_2461,In_1152,In_4680);
nor U2462 (N_2462,In_187,In_2656);
or U2463 (N_2463,In_1418,In_3467);
and U2464 (N_2464,In_339,In_3049);
nand U2465 (N_2465,In_154,In_2424);
nand U2466 (N_2466,In_2794,In_957);
or U2467 (N_2467,In_310,In_1245);
nor U2468 (N_2468,In_4665,In_4462);
or U2469 (N_2469,In_178,In_1658);
nand U2470 (N_2470,In_2634,In_4532);
and U2471 (N_2471,In_2201,In_3811);
or U2472 (N_2472,In_1899,In_2259);
xnor U2473 (N_2473,In_3504,In_501);
xor U2474 (N_2474,In_1984,In_468);
nand U2475 (N_2475,In_1939,In_2463);
or U2476 (N_2476,In_2101,In_2005);
nor U2477 (N_2477,In_4653,In_2570);
or U2478 (N_2478,In_4048,In_2563);
nand U2479 (N_2479,In_507,In_3249);
or U2480 (N_2480,In_90,In_3907);
xnor U2481 (N_2481,In_642,In_4663);
or U2482 (N_2482,In_2352,In_4896);
and U2483 (N_2483,In_3869,In_1483);
or U2484 (N_2484,In_3447,In_4344);
xnor U2485 (N_2485,In_4932,In_546);
nand U2486 (N_2486,In_3793,In_907);
nand U2487 (N_2487,In_4388,In_1258);
and U2488 (N_2488,In_2691,In_3640);
nand U2489 (N_2489,In_193,In_2075);
nand U2490 (N_2490,In_2837,In_8);
xor U2491 (N_2491,In_1267,In_2391);
xnor U2492 (N_2492,In_3669,In_3920);
nor U2493 (N_2493,In_4381,In_3115);
or U2494 (N_2494,In_4670,In_1767);
xor U2495 (N_2495,In_3379,In_4486);
xnor U2496 (N_2496,In_3543,In_2377);
or U2497 (N_2497,In_4860,In_738);
nand U2498 (N_2498,In_70,In_3912);
and U2499 (N_2499,In_2815,In_2460);
or U2500 (N_2500,N_909,N_1178);
nand U2501 (N_2501,N_850,N_1255);
nor U2502 (N_2502,N_71,N_290);
xor U2503 (N_2503,N_159,N_99);
xor U2504 (N_2504,N_687,N_1960);
nor U2505 (N_2505,N_123,N_566);
nand U2506 (N_2506,N_673,N_2339);
and U2507 (N_2507,N_1706,N_914);
nor U2508 (N_2508,N_2449,N_1689);
nand U2509 (N_2509,N_2210,N_374);
xnor U2510 (N_2510,N_2180,N_2322);
and U2511 (N_2511,N_1498,N_584);
nor U2512 (N_2512,N_1595,N_2133);
and U2513 (N_2513,N_1412,N_1929);
or U2514 (N_2514,N_1572,N_240);
nor U2515 (N_2515,N_379,N_1897);
and U2516 (N_2516,N_518,N_1793);
xor U2517 (N_2517,N_1359,N_1239);
and U2518 (N_2518,N_1446,N_2331);
nor U2519 (N_2519,N_2438,N_1494);
nor U2520 (N_2520,N_1371,N_1829);
and U2521 (N_2521,N_597,N_1490);
or U2522 (N_2522,N_1280,N_2475);
nor U2523 (N_2523,N_1373,N_1584);
or U2524 (N_2524,N_1386,N_416);
nand U2525 (N_2525,N_1089,N_1704);
nand U2526 (N_2526,N_1822,N_2398);
nand U2527 (N_2527,N_152,N_1390);
xnor U2528 (N_2528,N_2254,N_1661);
xnor U2529 (N_2529,N_1070,N_1059);
xnor U2530 (N_2530,N_1582,N_1886);
nor U2531 (N_2531,N_2484,N_522);
nand U2532 (N_2532,N_915,N_1741);
nand U2533 (N_2533,N_721,N_2122);
nand U2534 (N_2534,N_2059,N_1838);
and U2535 (N_2535,N_622,N_972);
nor U2536 (N_2536,N_1105,N_2186);
xor U2537 (N_2537,N_312,N_1121);
or U2538 (N_2538,N_2196,N_1338);
nand U2539 (N_2539,N_1214,N_1755);
xor U2540 (N_2540,N_1229,N_1055);
nand U2541 (N_2541,N_155,N_1348);
and U2542 (N_2542,N_1614,N_1443);
xor U2543 (N_2543,N_579,N_1631);
xor U2544 (N_2544,N_2417,N_1870);
nor U2545 (N_2545,N_2213,N_1890);
nand U2546 (N_2546,N_2234,N_1213);
and U2547 (N_2547,N_541,N_2300);
nor U2548 (N_2548,N_2263,N_790);
nor U2549 (N_2549,N_1778,N_29);
xor U2550 (N_2550,N_2230,N_1786);
xnor U2551 (N_2551,N_1128,N_223);
and U2552 (N_2552,N_1200,N_2402);
nand U2553 (N_2553,N_1097,N_248);
nor U2554 (N_2554,N_777,N_1516);
xnor U2555 (N_2555,N_1108,N_1647);
xor U2556 (N_2556,N_425,N_169);
nand U2557 (N_2557,N_979,N_1468);
xor U2558 (N_2558,N_1609,N_2400);
nand U2559 (N_2559,N_457,N_1035);
nand U2560 (N_2560,N_1326,N_2242);
and U2561 (N_2561,N_179,N_2321);
nor U2562 (N_2562,N_1707,N_1459);
nand U2563 (N_2563,N_399,N_308);
or U2564 (N_2564,N_745,N_1884);
nor U2565 (N_2565,N_2212,N_734);
nor U2566 (N_2566,N_2482,N_1841);
nand U2567 (N_2567,N_11,N_1159);
or U2568 (N_2568,N_2481,N_1362);
nor U2569 (N_2569,N_918,N_641);
nand U2570 (N_2570,N_750,N_276);
nor U2571 (N_2571,N_2315,N_217);
nand U2572 (N_2572,N_774,N_2163);
and U2573 (N_2573,N_807,N_1651);
or U2574 (N_2574,N_1976,N_1279);
or U2575 (N_2575,N_815,N_1915);
nand U2576 (N_2576,N_229,N_516);
xnor U2577 (N_2577,N_209,N_1283);
nand U2578 (N_2578,N_974,N_203);
and U2579 (N_2579,N_1204,N_2266);
or U2580 (N_2580,N_1478,N_508);
and U2581 (N_2581,N_1856,N_1228);
and U2582 (N_2582,N_221,N_1221);
nand U2583 (N_2583,N_2256,N_968);
xnor U2584 (N_2584,N_1470,N_1534);
or U2585 (N_2585,N_268,N_401);
or U2586 (N_2586,N_449,N_2349);
and U2587 (N_2587,N_250,N_2167);
xnor U2588 (N_2588,N_297,N_266);
or U2589 (N_2589,N_1501,N_836);
or U2590 (N_2590,N_231,N_978);
xnor U2591 (N_2591,N_162,N_1570);
nand U2592 (N_2592,N_1457,N_594);
nor U2593 (N_2593,N_166,N_1126);
and U2594 (N_2594,N_2022,N_2053);
or U2595 (N_2595,N_608,N_1286);
or U2596 (N_2596,N_2499,N_1546);
xor U2597 (N_2597,N_793,N_2393);
and U2598 (N_2598,N_2024,N_1678);
or U2599 (N_2599,N_1317,N_323);
and U2600 (N_2600,N_2420,N_1766);
xnor U2601 (N_2601,N_1690,N_1530);
xor U2602 (N_2602,N_356,N_1505);
or U2603 (N_2603,N_2013,N_693);
nand U2604 (N_2604,N_683,N_106);
or U2605 (N_2605,N_1549,N_1482);
or U2606 (N_2606,N_1119,N_477);
and U2607 (N_2607,N_1816,N_148);
and U2608 (N_2608,N_262,N_1571);
or U2609 (N_2609,N_1917,N_1529);
or U2610 (N_2610,N_277,N_2286);
nand U2611 (N_2611,N_444,N_1807);
nand U2612 (N_2612,N_831,N_1575);
nor U2613 (N_2613,N_1106,N_624);
nand U2614 (N_2614,N_1852,N_453);
xor U2615 (N_2615,N_94,N_232);
and U2616 (N_2616,N_171,N_1653);
and U2617 (N_2617,N_716,N_1940);
nand U2618 (N_2618,N_275,N_220);
nor U2619 (N_2619,N_945,N_860);
xor U2620 (N_2620,N_1994,N_325);
nor U2621 (N_2621,N_2343,N_1389);
xor U2622 (N_2622,N_332,N_722);
or U2623 (N_2623,N_2463,N_222);
nor U2624 (N_2624,N_822,N_1698);
nand U2625 (N_2625,N_908,N_950);
or U2626 (N_2626,N_156,N_1695);
xor U2627 (N_2627,N_56,N_135);
xor U2628 (N_2628,N_2176,N_1439);
or U2629 (N_2629,N_2363,N_1919);
xor U2630 (N_2630,N_922,N_1720);
nand U2631 (N_2631,N_208,N_2293);
xnor U2632 (N_2632,N_855,N_1319);
nand U2633 (N_2633,N_2302,N_2245);
xnor U2634 (N_2634,N_103,N_1088);
nand U2635 (N_2635,N_785,N_780);
nor U2636 (N_2636,N_853,N_2269);
nor U2637 (N_2637,N_633,N_1589);
xnor U2638 (N_2638,N_1834,N_1471);
nand U2639 (N_2639,N_581,N_554);
and U2640 (N_2640,N_1329,N_126);
and U2641 (N_2641,N_35,N_1835);
nand U2642 (N_2642,N_2221,N_435);
xnor U2643 (N_2643,N_1010,N_2088);
xnor U2644 (N_2644,N_576,N_2003);
nor U2645 (N_2645,N_2413,N_1564);
nand U2646 (N_2646,N_2277,N_625);
nor U2647 (N_2647,N_969,N_1650);
or U2648 (N_2648,N_2289,N_539);
and U2649 (N_2649,N_452,N_1368);
and U2650 (N_2650,N_489,N_1957);
nor U2651 (N_2651,N_821,N_2427);
or U2652 (N_2652,N_1504,N_799);
and U2653 (N_2653,N_2103,N_1869);
or U2654 (N_2654,N_747,N_600);
or U2655 (N_2655,N_1692,N_3);
or U2656 (N_2656,N_2419,N_2032);
and U2657 (N_2657,N_2169,N_344);
nor U2658 (N_2658,N_309,N_1056);
nand U2659 (N_2659,N_770,N_863);
xnor U2660 (N_2660,N_1710,N_2442);
and U2661 (N_2661,N_2008,N_1183);
nor U2662 (N_2662,N_1811,N_703);
nor U2663 (N_2663,N_238,N_2480);
xnor U2664 (N_2664,N_787,N_963);
or U2665 (N_2665,N_376,N_768);
xor U2666 (N_2666,N_1462,N_2428);
nand U2667 (N_2667,N_1515,N_2365);
xor U2668 (N_2668,N_1166,N_23);
or U2669 (N_2669,N_2185,N_475);
nand U2670 (N_2670,N_1023,N_810);
xor U2671 (N_2671,N_505,N_1627);
nor U2672 (N_2672,N_384,N_2236);
nor U2673 (N_2673,N_726,N_966);
and U2674 (N_2674,N_744,N_1274);
xor U2675 (N_2675,N_1987,N_2358);
or U2676 (N_2676,N_1218,N_928);
and U2677 (N_2677,N_841,N_797);
xor U2678 (N_2678,N_940,N_2430);
nor U2679 (N_2679,N_769,N_1644);
or U2680 (N_2680,N_1448,N_2392);
nand U2681 (N_2681,N_1768,N_1536);
nand U2682 (N_2682,N_136,N_1618);
and U2683 (N_2683,N_1007,N_1230);
nor U2684 (N_2684,N_1879,N_1270);
nand U2685 (N_2685,N_2492,N_1261);
and U2686 (N_2686,N_251,N_1580);
and U2687 (N_2687,N_424,N_2173);
nor U2688 (N_2688,N_2435,N_57);
nand U2689 (N_2689,N_2182,N_65);
nand U2690 (N_2690,N_611,N_1949);
and U2691 (N_2691,N_194,N_1406);
and U2692 (N_2692,N_271,N_1115);
xor U2693 (N_2693,N_143,N_2247);
and U2694 (N_2694,N_2389,N_341);
and U2695 (N_2695,N_1712,N_1563);
or U2696 (N_2696,N_1970,N_1956);
or U2697 (N_2697,N_41,N_2165);
or U2698 (N_2698,N_1713,N_1107);
and U2699 (N_2699,N_1938,N_827);
nor U2700 (N_2700,N_1747,N_613);
and U2701 (N_2701,N_1892,N_2011);
and U2702 (N_2702,N_652,N_2062);
and U2703 (N_2703,N_858,N_236);
or U2704 (N_2704,N_2267,N_2487);
or U2705 (N_2705,N_32,N_2127);
xnor U2706 (N_2706,N_134,N_852);
nor U2707 (N_2707,N_733,N_102);
xor U2708 (N_2708,N_2136,N_1012);
nor U2709 (N_2709,N_2474,N_2399);
nand U2710 (N_2710,N_1775,N_939);
and U2711 (N_2711,N_1544,N_259);
and U2712 (N_2712,N_1091,N_1281);
or U2713 (N_2713,N_2423,N_1154);
and U2714 (N_2714,N_691,N_1437);
xor U2715 (N_2715,N_2191,N_2327);
or U2716 (N_2716,N_1477,N_2052);
or U2717 (N_2717,N_2206,N_524);
and U2718 (N_2718,N_1854,N_1637);
xor U2719 (N_2719,N_514,N_732);
and U2720 (N_2720,N_50,N_2498);
nor U2721 (N_2721,N_1765,N_619);
or U2722 (N_2722,N_1199,N_1265);
nor U2723 (N_2723,N_568,N_183);
xor U2724 (N_2724,N_1723,N_87);
nand U2725 (N_2725,N_2066,N_1846);
nand U2726 (N_2726,N_1287,N_2189);
and U2727 (N_2727,N_390,N_484);
and U2728 (N_2728,N_953,N_2275);
nor U2729 (N_2729,N_854,N_1761);
nand U2730 (N_2730,N_748,N_2068);
xnor U2731 (N_2731,N_1728,N_544);
or U2732 (N_2732,N_1782,N_218);
xnor U2733 (N_2733,N_1875,N_583);
or U2734 (N_2734,N_2425,N_235);
or U2735 (N_2735,N_1352,N_1951);
nor U2736 (N_2736,N_2406,N_656);
nand U2737 (N_2737,N_96,N_2380);
xor U2738 (N_2738,N_2395,N_450);
and U2739 (N_2739,N_359,N_752);
xnor U2740 (N_2740,N_1377,N_1292);
xor U2741 (N_2741,N_172,N_402);
nor U2742 (N_2742,N_127,N_1150);
nor U2743 (N_2743,N_1821,N_1000);
nor U2744 (N_2744,N_174,N_1005);
nor U2745 (N_2745,N_1903,N_1052);
nor U2746 (N_2746,N_1509,N_371);
nand U2747 (N_2747,N_2273,N_1020);
nor U2748 (N_2748,N_1111,N_809);
xnor U2749 (N_2749,N_669,N_1933);
xor U2750 (N_2750,N_1797,N_1655);
nand U2751 (N_2751,N_2055,N_519);
or U2752 (N_2752,N_1624,N_1163);
and U2753 (N_2753,N_2067,N_2007);
xor U2754 (N_2754,N_1688,N_1048);
or U2755 (N_2755,N_936,N_2243);
and U2756 (N_2756,N_988,N_320);
or U2757 (N_2757,N_663,N_101);
and U2758 (N_2758,N_2458,N_2489);
nand U2759 (N_2759,N_1525,N_1717);
and U2760 (N_2760,N_832,N_2453);
nor U2761 (N_2761,N_2057,N_636);
xnor U2762 (N_2762,N_789,N_382);
nor U2763 (N_2763,N_1619,N_1353);
xor U2764 (N_2764,N_1559,N_912);
nand U2765 (N_2765,N_1885,N_1735);
or U2766 (N_2766,N_365,N_666);
or U2767 (N_2767,N_383,N_2290);
and U2768 (N_2768,N_2382,N_531);
nor U2769 (N_2769,N_1606,N_779);
nor U2770 (N_2770,N_1585,N_1641);
or U2771 (N_2771,N_2328,N_1794);
or U2772 (N_2772,N_2356,N_2312);
nand U2773 (N_2773,N_1962,N_2366);
and U2774 (N_2774,N_2126,N_1422);
xor U2775 (N_2775,N_2050,N_1551);
xor U2776 (N_2776,N_2376,N_949);
nand U2777 (N_2777,N_1664,N_1672);
or U2778 (N_2778,N_1812,N_137);
nand U2779 (N_2779,N_696,N_2405);
nand U2780 (N_2780,N_1250,N_1764);
or U2781 (N_2781,N_1302,N_1535);
or U2782 (N_2782,N_2421,N_82);
nand U2783 (N_2783,N_555,N_158);
nand U2784 (N_2784,N_1050,N_2285);
or U2785 (N_2785,N_1165,N_980);
and U2786 (N_2786,N_2394,N_1438);
or U2787 (N_2787,N_49,N_2340);
and U2788 (N_2788,N_1864,N_1784);
or U2789 (N_2789,N_1074,N_496);
xor U2790 (N_2790,N_1420,N_1931);
nand U2791 (N_2791,N_1288,N_336);
or U2792 (N_2792,N_2369,N_196);
nand U2793 (N_2793,N_2037,N_527);
and U2794 (N_2794,N_1959,N_386);
or U2795 (N_2795,N_1577,N_642);
or U2796 (N_2796,N_2351,N_108);
nor U2797 (N_2797,N_413,N_1634);
and U2798 (N_2798,N_2145,N_1136);
nor U2799 (N_2799,N_1853,N_1001);
and U2800 (N_2800,N_1944,N_4);
xnor U2801 (N_2801,N_274,N_2161);
nand U2802 (N_2802,N_1227,N_1145);
and U2803 (N_2803,N_1922,N_1351);
or U2804 (N_2804,N_72,N_2344);
and U2805 (N_2805,N_2171,N_2249);
xnor U2806 (N_2806,N_2432,N_1667);
nand U2807 (N_2807,N_1744,N_1324);
xor U2808 (N_2808,N_2486,N_758);
nor U2809 (N_2809,N_944,N_864);
nand U2810 (N_2810,N_177,N_2283);
xnor U2811 (N_2811,N_2459,N_987);
nand U2812 (N_2812,N_1349,N_2086);
or U2813 (N_2813,N_1135,N_1034);
nor U2814 (N_2814,N_881,N_1493);
or U2815 (N_2815,N_1289,N_1697);
nor U2816 (N_2816,N_125,N_133);
or U2817 (N_2817,N_783,N_2326);
nand U2818 (N_2818,N_898,N_24);
nand U2819 (N_2819,N_1560,N_671);
or U2820 (N_2820,N_364,N_2232);
and U2821 (N_2821,N_2317,N_110);
nor U2822 (N_2822,N_757,N_702);
nor U2823 (N_2823,N_2105,N_2426);
and U2824 (N_2824,N_367,N_160);
or U2825 (N_2825,N_1857,N_1923);
xor U2826 (N_2826,N_1431,N_537);
nor U2827 (N_2827,N_1485,N_1781);
and U2828 (N_2828,N_1346,N_1401);
and U2829 (N_2829,N_1855,N_1557);
and U2830 (N_2830,N_2143,N_1750);
nand U2831 (N_2831,N_1068,N_1888);
nand U2832 (N_2832,N_2454,N_926);
and U2833 (N_2833,N_948,N_1943);
xor U2834 (N_2834,N_919,N_628);
and U2835 (N_2835,N_2334,N_707);
nand U2836 (N_2836,N_894,N_812);
nand U2837 (N_2837,N_753,N_2391);
or U2838 (N_2838,N_1427,N_1926);
xnor U2839 (N_2839,N_1593,N_1341);
nand U2840 (N_2840,N_2350,N_1285);
and U2841 (N_2841,N_612,N_2109);
nand U2842 (N_2842,N_1837,N_478);
or U2843 (N_2843,N_615,N_1550);
nor U2844 (N_2844,N_1849,N_1451);
xor U2845 (N_2845,N_756,N_331);
xnor U2846 (N_2846,N_202,N_1964);
nor U2847 (N_2847,N_2306,N_515);
or U2848 (N_2848,N_2033,N_1918);
nand U2849 (N_2849,N_1263,N_1850);
xor U2850 (N_2850,N_2036,N_715);
or U2851 (N_2851,N_1298,N_1700);
and U2852 (N_2852,N_749,N_2381);
nand U2853 (N_2853,N_1632,N_645);
xor U2854 (N_2854,N_982,N_1969);
xnor U2855 (N_2855,N_1225,N_291);
xor U2856 (N_2856,N_1517,N_754);
or U2857 (N_2857,N_2259,N_1124);
or U2858 (N_2858,N_1830,N_1084);
or U2859 (N_2859,N_1612,N_471);
or U2860 (N_2860,N_2168,N_2412);
nand U2861 (N_2861,N_132,N_762);
or U2862 (N_2862,N_317,N_1998);
nand U2863 (N_2863,N_113,N_2114);
xor U2864 (N_2864,N_2462,N_1568);
nor U2865 (N_2865,N_2238,N_1629);
and U2866 (N_2866,N_1787,N_1952);
nor U2867 (N_2867,N_1907,N_714);
xor U2868 (N_2868,N_2305,N_557);
or U2869 (N_2869,N_1144,N_142);
or U2870 (N_2870,N_368,N_1920);
nor U2871 (N_2871,N_1848,N_1312);
or U2872 (N_2872,N_977,N_438);
nand U2873 (N_2873,N_362,N_662);
nand U2874 (N_2874,N_1311,N_1833);
nand U2875 (N_2875,N_2219,N_1681);
and U2876 (N_2876,N_2264,N_2104);
nand U2877 (N_2877,N_335,N_587);
or U2878 (N_2878,N_429,N_1963);
or U2879 (N_2879,N_1172,N_1520);
xor U2880 (N_2880,N_150,N_1566);
nand U2881 (N_2881,N_322,N_442);
and U2882 (N_2882,N_873,N_543);
and U2883 (N_2883,N_2288,N_128);
and U2884 (N_2884,N_1561,N_635);
nand U2885 (N_2885,N_742,N_2370);
nor U2886 (N_2886,N_660,N_2142);
and U2887 (N_2887,N_327,N_479);
and U2888 (N_2888,N_1212,N_1016);
nor U2889 (N_2889,N_1014,N_1461);
xnor U2890 (N_2890,N_1621,N_1540);
and U2891 (N_2891,N_440,N_140);
xnor U2892 (N_2892,N_2360,N_975);
and U2893 (N_2893,N_588,N_54);
or U2894 (N_2894,N_1394,N_616);
xnor U2895 (N_2895,N_2401,N_1992);
or U2896 (N_2896,N_73,N_1103);
nor U2897 (N_2897,N_995,N_2025);
nand U2898 (N_2898,N_1565,N_866);
xor U2899 (N_2899,N_1046,N_675);
or U2900 (N_2900,N_1125,N_892);
and U2901 (N_2901,N_2000,N_1981);
nor U2902 (N_2902,N_292,N_353);
nor U2903 (N_2903,N_303,N_1383);
nor U2904 (N_2904,N_736,N_1798);
nand U2905 (N_2905,N_2320,N_569);
or U2906 (N_2906,N_2457,N_1425);
and U2907 (N_2907,N_1411,N_361);
xor U2908 (N_2908,N_1148,N_1539);
nand U2909 (N_2909,N_788,N_283);
or U2910 (N_2910,N_1282,N_1098);
nor U2911 (N_2911,N_2108,N_617);
or U2912 (N_2912,N_2139,N_1308);
xnor U2913 (N_2913,N_760,N_324);
nand U2914 (N_2914,N_792,N_1814);
xor U2915 (N_2915,N_2010,N_1002);
and U2916 (N_2916,N_738,N_817);
xor U2917 (N_2917,N_1331,N_1259);
nand U2918 (N_2918,N_849,N_761);
and U2919 (N_2919,N_1616,N_534);
nand U2920 (N_2920,N_1521,N_1090);
or U2921 (N_2921,N_637,N_655);
and U2922 (N_2922,N_2079,N_800);
and U2923 (N_2923,N_1077,N_2026);
nand U2924 (N_2924,N_1599,N_2437);
or U2925 (N_2925,N_1615,N_418);
or U2926 (N_2926,N_574,N_163);
and U2927 (N_2927,N_84,N_801);
nor U2928 (N_2928,N_2129,N_2157);
nand U2929 (N_2929,N_1330,N_388);
nand U2930 (N_2930,N_1581,N_2237);
or U2931 (N_2931,N_2301,N_773);
or U2932 (N_2932,N_1979,N_91);
and U2933 (N_2933,N_1435,N_965);
or U2934 (N_2934,N_2071,N_985);
and U2935 (N_2935,N_1044,N_803);
nor U2936 (N_2936,N_2478,N_1210);
xnor U2937 (N_2937,N_2252,N_2205);
xor U2938 (N_2938,N_154,N_1300);
or U2939 (N_2939,N_431,N_2233);
nand U2940 (N_2940,N_1398,N_1416);
nand U2941 (N_2941,N_2470,N_2359);
or U2942 (N_2942,N_775,N_2496);
nand U2943 (N_2943,N_2411,N_621);
or U2944 (N_2944,N_1791,N_2319);
nand U2945 (N_2945,N_1184,N_2497);
and U2946 (N_2946,N_265,N_1973);
and U2947 (N_2947,N_1021,N_1305);
nand U2948 (N_2948,N_1640,N_1999);
and U2949 (N_2949,N_375,N_1466);
or U2950 (N_2950,N_2479,N_1924);
nand U2951 (N_2951,N_1232,N_443);
xor U2952 (N_2952,N_6,N_2132);
xor U2953 (N_2953,N_369,N_1009);
or U2954 (N_2954,N_517,N_1278);
and U2955 (N_2955,N_970,N_389);
xor U2956 (N_2956,N_875,N_1209);
and U2957 (N_2957,N_1909,N_1906);
xnor U2958 (N_2958,N_139,N_1284);
nand U2959 (N_2959,N_1902,N_1442);
and U2960 (N_2960,N_192,N_153);
nor U2961 (N_2961,N_772,N_242);
nand U2962 (N_2962,N_2016,N_258);
and U2963 (N_2963,N_1488,N_2451);
nor U2964 (N_2964,N_2063,N_1967);
nand U2965 (N_2965,N_2075,N_1407);
or U2966 (N_2966,N_1272,N_1036);
and U2967 (N_2967,N_596,N_1067);
nand U2968 (N_2968,N_2117,N_490);
xor U2969 (N_2969,N_1845,N_310);
or U2970 (N_2970,N_1739,N_2012);
xor U2971 (N_2971,N_536,N_2258);
xor U2972 (N_2972,N_1388,N_1642);
and U2973 (N_2973,N_2092,N_1134);
xnor U2974 (N_2974,N_109,N_403);
or U2975 (N_2975,N_1513,N_2031);
nor U2976 (N_2976,N_2134,N_1017);
nand U2977 (N_2977,N_816,N_1235);
nand U2978 (N_2978,N_37,N_935);
and U2979 (N_2979,N_2078,N_244);
xor U2980 (N_2980,N_649,N_1731);
nor U2981 (N_2981,N_571,N_2342);
or U2982 (N_2982,N_937,N_2183);
xor U2983 (N_2983,N_823,N_1452);
xor U2984 (N_2984,N_167,N_89);
nand U2985 (N_2985,N_2323,N_2061);
and U2986 (N_2986,N_427,N_1267);
or U2987 (N_2987,N_2082,N_1414);
xor U2988 (N_2988,N_2341,N_1531);
nor U2989 (N_2989,N_1809,N_207);
nand U2990 (N_2990,N_1365,N_2228);
or U2991 (N_2991,N_1487,N_377);
nand U2992 (N_2992,N_1122,N_751);
and U2993 (N_2993,N_609,N_1156);
or U2994 (N_2994,N_1109,N_905);
nor U2995 (N_2995,N_178,N_2130);
nand U2996 (N_2996,N_193,N_598);
nor U2997 (N_2997,N_2148,N_42);
xnor U2998 (N_2998,N_1719,N_2455);
nor U2999 (N_2999,N_2065,N_2076);
or U3000 (N_3000,N_766,N_339);
and U3001 (N_3001,N_2468,N_2215);
and U3002 (N_3002,N_657,N_107);
xor U3003 (N_3003,N_387,N_407);
xor U3004 (N_3004,N_412,N_114);
xor U3005 (N_3005,N_931,N_2379);
nor U3006 (N_3006,N_1481,N_877);
or U3007 (N_3007,N_2407,N_2388);
or U3008 (N_3008,N_45,N_701);
or U3009 (N_3009,N_629,N_795);
or U3010 (N_3010,N_157,N_1276);
or U3011 (N_3011,N_7,N_355);
or U3012 (N_3012,N_472,N_1939);
or U3013 (N_3013,N_906,N_771);
xnor U3014 (N_3014,N_1972,N_626);
xnor U3015 (N_3015,N_415,N_1669);
and U3016 (N_3016,N_2329,N_1169);
and U3017 (N_3017,N_1233,N_1188);
nand U3018 (N_3018,N_1541,N_958);
nor U3019 (N_3019,N_278,N_151);
nor U3020 (N_3020,N_2345,N_20);
nand U3021 (N_3021,N_1767,N_111);
xnor U3022 (N_3022,N_2098,N_706);
nand U3023 (N_3023,N_1323,N_2177);
nor U3024 (N_3024,N_1151,N_592);
or U3025 (N_3025,N_1583,N_562);
or U3026 (N_3026,N_436,N_565);
nor U3027 (N_3027,N_2051,N_589);
nor U3028 (N_3028,N_206,N_2146);
nand U3029 (N_3029,N_225,N_1075);
nor U3030 (N_3030,N_981,N_1360);
nor U3031 (N_3031,N_1162,N_1528);
nand U3032 (N_3032,N_1792,N_2260);
nor U3033 (N_3033,N_1060,N_381);
and U3034 (N_3034,N_1455,N_474);
and U3035 (N_3035,N_2035,N_346);
and U3036 (N_3036,N_195,N_104);
or U3037 (N_3037,N_667,N_2081);
nor U3038 (N_3038,N_454,N_575);
and U3039 (N_3039,N_2361,N_2039);
xor U3040 (N_3040,N_1019,N_464);
nand U3041 (N_3041,N_1260,N_1301);
and U3042 (N_3042,N_2138,N_1754);
or U3043 (N_3043,N_1527,N_1366);
and U3044 (N_3044,N_2152,N_808);
xnor U3045 (N_3045,N_2352,N_647);
nand U3046 (N_3046,N_394,N_2397);
or U3047 (N_3047,N_1824,N_1393);
nand U3048 (N_3048,N_907,N_2002);
nor U3049 (N_3049,N_318,N_1403);
or U3050 (N_3050,N_1054,N_2222);
nand U3051 (N_3051,N_838,N_2477);
xor U3052 (N_3052,N_746,N_1733);
or U3053 (N_3053,N_2083,N_345);
xnor U3054 (N_3054,N_1607,N_1553);
and U3055 (N_3055,N_1428,N_2330);
nand U3056 (N_3056,N_1079,N_1078);
and U3057 (N_3057,N_796,N_885);
or U3058 (N_3058,N_1757,N_2429);
xor U3059 (N_3059,N_741,N_1685);
nor U3060 (N_3060,N_164,N_470);
nor U3061 (N_3061,N_1454,N_902);
xnor U3062 (N_3062,N_879,N_1004);
nor U3063 (N_3063,N_233,N_1600);
xnor U3064 (N_3064,N_2390,N_763);
and U3065 (N_3065,N_1133,N_546);
nand U3066 (N_3066,N_538,N_1149);
nor U3067 (N_3067,N_227,N_1173);
xnor U3068 (N_3068,N_1950,N_1860);
xor U3069 (N_3069,N_2307,N_19);
nand U3070 (N_3070,N_165,N_279);
nor U3071 (N_3071,N_366,N_1586);
nand U3072 (N_3072,N_1226,N_1293);
nor U3073 (N_3073,N_711,N_2223);
or U3074 (N_3074,N_1249,N_2089);
or U3075 (N_3075,N_1769,N_12);
or U3076 (N_3076,N_2030,N_582);
and U3077 (N_3077,N_406,N_2488);
and U3078 (N_3078,N_901,N_1480);
xor U3079 (N_3079,N_2160,N_1257);
nor U3080 (N_3080,N_1913,N_993);
and U3081 (N_3081,N_1831,N_2207);
nand U3082 (N_3082,N_2313,N_632);
nand U3083 (N_3083,N_1175,N_674);
or U3084 (N_3084,N_1396,N_446);
nand U3085 (N_3085,N_1948,N_63);
and U3086 (N_3086,N_458,N_2113);
nand U3087 (N_3087,N_44,N_1803);
and U3088 (N_3088,N_311,N_116);
or U3089 (N_3089,N_1160,N_2135);
nor U3090 (N_3090,N_396,N_243);
nand U3091 (N_3091,N_1955,N_1198);
nor U3092 (N_3092,N_1484,N_1898);
nor U3093 (N_3093,N_665,N_1726);
xor U3094 (N_3094,N_830,N_859);
nand U3095 (N_3095,N_699,N_468);
xnor U3096 (N_3096,N_1339,N_2476);
nor U3097 (N_3097,N_1147,N_1779);
nand U3098 (N_3098,N_1718,N_2080);
nor U3099 (N_3099,N_2287,N_845);
nand U3100 (N_3100,N_2456,N_1186);
nand U3101 (N_3101,N_1800,N_1361);
and U3102 (N_3102,N_973,N_170);
nand U3103 (N_3103,N_578,N_1142);
or U3104 (N_3104,N_486,N_500);
xor U3105 (N_3105,N_1840,N_1780);
xor U3106 (N_3106,N_1673,N_547);
nand U3107 (N_3107,N_1668,N_1161);
nand U3108 (N_3108,N_1400,N_1828);
nand U3109 (N_3109,N_86,N_1993);
or U3110 (N_3110,N_481,N_1025);
xnor U3111 (N_3111,N_1727,N_1062);
xnor U3112 (N_3112,N_2096,N_1345);
xnor U3113 (N_3113,N_2311,N_1483);
or U3114 (N_3114,N_717,N_100);
nor U3115 (N_3115,N_679,N_1945);
nor U3116 (N_3116,N_1242,N_1086);
xnor U3117 (N_3117,N_319,N_1203);
or U3118 (N_3118,N_420,N_542);
and U3119 (N_3119,N_585,N_2216);
xnor U3120 (N_3120,N_261,N_451);
or U3121 (N_3121,N_2018,N_1876);
or U3122 (N_3122,N_487,N_2077);
nor U3123 (N_3123,N_88,N_98);
nor U3124 (N_3124,N_564,N_426);
and U3125 (N_3125,N_989,N_971);
or U3126 (N_3126,N_282,N_1350);
and U3127 (N_3127,N_392,N_482);
nor U3128 (N_3128,N_358,N_1240);
or U3129 (N_3129,N_2198,N_1871);
xor U3130 (N_3130,N_2046,N_1453);
xnor U3131 (N_3131,N_1355,N_1709);
xnor U3132 (N_3132,N_2038,N_2029);
and U3133 (N_3133,N_1666,N_1721);
or U3134 (N_3134,N_2452,N_1456);
xnor U3135 (N_3135,N_428,N_1802);
and U3136 (N_3136,N_1370,N_1610);
and U3137 (N_3137,N_2297,N_1063);
xor U3138 (N_3138,N_1506,N_213);
and U3139 (N_3139,N_603,N_2115);
or U3140 (N_3140,N_1574,N_828);
and U3141 (N_3141,N_1347,N_523);
nor U3142 (N_3142,N_495,N_2054);
and U3143 (N_3143,N_2015,N_1474);
and U3144 (N_3144,N_872,N_954);
nor U3145 (N_3145,N_943,N_1748);
or U3146 (N_3146,N_529,N_959);
and U3147 (N_3147,N_731,N_1381);
xor U3148 (N_3148,N_219,N_2192);
nand U3149 (N_3149,N_1878,N_1391);
and U3150 (N_3150,N_499,N_1788);
or U3151 (N_3151,N_1908,N_1654);
nand U3152 (N_3152,N_161,N_1708);
and U3153 (N_3153,N_2048,N_1185);
or U3154 (N_3154,N_2102,N_296);
nand U3155 (N_3155,N_1639,N_187);
nor U3156 (N_3156,N_370,N_1405);
or U3157 (N_3157,N_1153,N_1423);
xnor U3158 (N_3158,N_74,N_2009);
or U3159 (N_3159,N_1817,N_1497);
nand U3160 (N_3160,N_395,N_269);
xnor U3161 (N_3161,N_447,N_1927);
nand U3162 (N_3162,N_868,N_0);
nor U3163 (N_3163,N_1662,N_295);
xnor U3164 (N_3164,N_784,N_117);
nor U3165 (N_3165,N_373,N_272);
nor U3166 (N_3166,N_284,N_2373);
or U3167 (N_3167,N_2235,N_2120);
nand U3168 (N_3168,N_1804,N_2461);
xor U3169 (N_3169,N_1436,N_1789);
xnor U3170 (N_3170,N_34,N_1508);
xor U3171 (N_3171,N_2495,N_503);
nor U3172 (N_3172,N_1222,N_623);
or U3173 (N_3173,N_2353,N_511);
nor U3174 (N_3174,N_260,N_1426);
or U3175 (N_3175,N_1189,N_1152);
xnor U3176 (N_3176,N_1295,N_1752);
xor U3177 (N_3177,N_2158,N_273);
nand U3178 (N_3178,N_337,N_886);
and U3179 (N_3179,N_2375,N_498);
nor U3180 (N_3180,N_1714,N_1635);
nand U3181 (N_3181,N_560,N_932);
xnor U3182 (N_3182,N_2118,N_506);
xnor U3183 (N_3183,N_601,N_204);
xnor U3184 (N_3184,N_1116,N_39);
and U3185 (N_3185,N_239,N_781);
xor U3186 (N_3186,N_1127,N_144);
and U3187 (N_3187,N_2299,N_2485);
xor U3188 (N_3188,N_1219,N_1337);
or U3189 (N_3189,N_467,N_2005);
or U3190 (N_3190,N_708,N_804);
or U3191 (N_3191,N_27,N_2017);
nand U3192 (N_3192,N_690,N_512);
and U3193 (N_3193,N_1296,N_1065);
and U3194 (N_3194,N_301,N_1031);
or U3195 (N_3195,N_492,N_2491);
xnor U3196 (N_3196,N_305,N_806);
nand U3197 (N_3197,N_1357,N_720);
nor U3198 (N_3198,N_2229,N_1538);
nor U3199 (N_3199,N_1313,N_205);
xnor U3200 (N_3200,N_513,N_857);
and U3201 (N_3201,N_1071,N_1805);
or U3202 (N_3202,N_2418,N_680);
nand U3203 (N_3203,N_737,N_1315);
or U3204 (N_3204,N_729,N_1303);
and U3205 (N_3205,N_2308,N_480);
and U3206 (N_3206,N_1882,N_1573);
nor U3207 (N_3207,N_1971,N_2472);
and U3208 (N_3208,N_2409,N_302);
and U3209 (N_3209,N_1602,N_1363);
nor U3210 (N_3210,N_58,N_1170);
or U3211 (N_3211,N_1510,N_814);
nor U3212 (N_3212,N_2014,N_1340);
and U3213 (N_3213,N_844,N_1532);
xor U3214 (N_3214,N_1995,N_1702);
or U3215 (N_3215,N_1138,N_118);
or U3216 (N_3216,N_294,N_1399);
nor U3217 (N_3217,N_2153,N_408);
or U3218 (N_3218,N_1826,N_247);
or U3219 (N_3219,N_1638,N_1343);
and U3220 (N_3220,N_78,N_851);
and U3221 (N_3221,N_556,N_2211);
and U3222 (N_3222,N_1143,N_553);
xor U3223 (N_3223,N_1705,N_1057);
nand U3224 (N_3224,N_1310,N_740);
or U3225 (N_3225,N_445,N_946);
nor U3226 (N_3226,N_2253,N_129);
nand U3227 (N_3227,N_1003,N_1533);
and U3228 (N_3228,N_2203,N_1756);
xnor U3229 (N_3229,N_618,N_314);
xor U3230 (N_3230,N_181,N_648);
xor U3231 (N_3231,N_900,N_1562);
nor U3232 (N_3232,N_2355,N_1495);
or U3233 (N_3233,N_961,N_1968);
or U3234 (N_3234,N_2199,N_2006);
xor U3235 (N_3235,N_2314,N_33);
and U3236 (N_3236,N_321,N_1058);
nor U3237 (N_3237,N_1449,N_465);
nor U3238 (N_3238,N_423,N_723);
nand U3239 (N_3239,N_530,N_1215);
and U3240 (N_3240,N_895,N_1114);
and U3241 (N_3241,N_228,N_923);
nor U3242 (N_3242,N_1262,N_846);
xor U3243 (N_3243,N_1628,N_2362);
and U3244 (N_3244,N_2439,N_21);
nor U3245 (N_3245,N_55,N_1989);
xor U3246 (N_3246,N_1941,N_957);
nand U3247 (N_3247,N_307,N_2060);
nor U3248 (N_3248,N_257,N_1901);
nor U3249 (N_3249,N_559,N_990);
nor U3250 (N_3250,N_2044,N_2023);
nor U3251 (N_3251,N_1524,N_1177);
or U3252 (N_3252,N_393,N_920);
nor U3253 (N_3253,N_147,N_1984);
xor U3254 (N_3254,N_1201,N_1523);
and U3255 (N_3255,N_1013,N_1392);
nor U3256 (N_3256,N_315,N_570);
nand U3257 (N_3257,N_2445,N_1395);
nor U3258 (N_3258,N_1937,N_2);
nor U3259 (N_3259,N_1514,N_1237);
xnor U3260 (N_3260,N_1325,N_2251);
and U3261 (N_3261,N_1447,N_201);
and U3262 (N_3262,N_190,N_1157);
nor U3263 (N_3263,N_1623,N_26);
or U3264 (N_3264,N_304,N_1131);
and U3265 (N_3265,N_1519,N_2384);
and U3266 (N_3266,N_2121,N_2473);
xnor U3267 (N_3267,N_2164,N_1328);
xnor U3268 (N_3268,N_1930,N_929);
or U3269 (N_3269,N_1254,N_1608);
nand U3270 (N_3270,N_630,N_2184);
nor U3271 (N_3271,N_1072,N_1676);
nor U3272 (N_3272,N_2147,N_728);
and U3273 (N_3273,N_1660,N_46);
and U3274 (N_3274,N_1061,N_709);
nand U3275 (N_3275,N_1663,N_2443);
or U3276 (N_3276,N_298,N_567);
nor U3277 (N_3277,N_847,N_1649);
xor U3278 (N_3278,N_1243,N_2028);
nor U3279 (N_3279,N_2414,N_1397);
nor U3280 (N_3280,N_1087,N_333);
and U3281 (N_3281,N_1432,N_326);
xor U3282 (N_3282,N_404,N_264);
nand U3283 (N_3283,N_189,N_1332);
or U3284 (N_3284,N_684,N_1047);
and U3285 (N_3285,N_16,N_2284);
and U3286 (N_3286,N_216,N_639);
nor U3287 (N_3287,N_1935,N_79);
xor U3288 (N_3288,N_1877,N_1093);
nand U3289 (N_3289,N_840,N_2073);
and U3290 (N_3290,N_1548,N_904);
nand U3291 (N_3291,N_1671,N_1027);
nor U3292 (N_3292,N_843,N_2069);
nor U3293 (N_3293,N_1537,N_1472);
and U3294 (N_3294,N_2346,N_349);
nor U3295 (N_3295,N_13,N_2446);
xor U3296 (N_3296,N_2268,N_1460);
xnor U3297 (N_3297,N_507,N_285);
or U3298 (N_3298,N_1716,N_491);
or U3299 (N_3299,N_2072,N_533);
nand U3300 (N_3300,N_997,N_1430);
and U3301 (N_3301,N_1217,N_2123);
and U3302 (N_3302,N_2282,N_15);
nand U3303 (N_3303,N_2174,N_1440);
nand U3304 (N_3304,N_938,N_210);
and U3305 (N_3305,N_991,N_1771);
nand U3306 (N_3306,N_986,N_25);
xnor U3307 (N_3307,N_1576,N_93);
or U3308 (N_3308,N_956,N_561);
nand U3309 (N_3309,N_2279,N_1730);
xor U3310 (N_3310,N_1974,N_2466);
and U3311 (N_3311,N_1168,N_1429);
nor U3312 (N_3312,N_421,N_168);
nand U3313 (N_3313,N_64,N_1465);
or U3314 (N_3314,N_286,N_2460);
nand U3315 (N_3315,N_36,N_2444);
or U3316 (N_3316,N_2220,N_105);
nand U3317 (N_3317,N_1904,N_441);
or U3318 (N_3318,N_1404,N_1354);
and U3319 (N_3319,N_1722,N_461);
nand U3320 (N_3320,N_70,N_510);
and U3321 (N_3321,N_1785,N_638);
or U3322 (N_3322,N_876,N_197);
nand U3323 (N_3323,N_834,N_75);
xor U3324 (N_3324,N_1421,N_1759);
xnor U3325 (N_3325,N_1512,N_1045);
and U3326 (N_3326,N_1092,N_1264);
nand U3327 (N_3327,N_1110,N_61);
or U3328 (N_3328,N_141,N_1307);
xor U3329 (N_3329,N_1659,N_710);
and U3330 (N_3330,N_1912,N_640);
and U3331 (N_3331,N_357,N_1921);
or U3332 (N_3332,N_1975,N_398);
nor U3333 (N_3333,N_347,N_1380);
and U3334 (N_3334,N_1896,N_1051);
nor U3335 (N_3335,N_1832,N_725);
nor U3336 (N_3336,N_352,N_372);
and U3337 (N_3337,N_348,N_1123);
or U3338 (N_3338,N_1732,N_1299);
nand U3339 (N_3339,N_550,N_967);
nand U3340 (N_3340,N_175,N_927);
nor U3341 (N_3341,N_289,N_1191);
xnor U3342 (N_3342,N_880,N_2244);
nor U3343 (N_3343,N_2021,N_22);
nor U3344 (N_3344,N_2224,N_1889);
and U3345 (N_3345,N_299,N_2416);
nor U3346 (N_3346,N_1858,N_1740);
nor U3347 (N_3347,N_1648,N_1095);
or U3348 (N_3348,N_681,N_1626);
and U3349 (N_3349,N_1745,N_2131);
or U3350 (N_3350,N_835,N_535);
and U3351 (N_3351,N_2280,N_1772);
nor U3352 (N_3352,N_1865,N_1543);
nor U3353 (N_3353,N_1120,N_199);
and U3354 (N_3354,N_397,N_1985);
nand U3355 (N_3355,N_2162,N_1823);
and U3356 (N_3356,N_917,N_688);
nand U3357 (N_3357,N_1139,N_1132);
and U3358 (N_3358,N_2181,N_1476);
nand U3359 (N_3359,N_343,N_634);
xor U3360 (N_3360,N_405,N_1018);
or U3361 (N_3361,N_983,N_833);
nor U3362 (N_3362,N_672,N_1859);
nor U3363 (N_3363,N_1385,N_1309);
or U3364 (N_3364,N_659,N_2357);
xnor U3365 (N_3365,N_924,N_115);
nand U3366 (N_3366,N_1502,N_1934);
nand U3367 (N_3367,N_1445,N_18);
or U3368 (N_3368,N_422,N_2156);
and U3369 (N_3369,N_1636,N_466);
xnor U3370 (N_3370,N_112,N_540);
xnor U3371 (N_3371,N_338,N_1463);
and U3372 (N_3372,N_1613,N_2387);
and U3373 (N_3373,N_2151,N_631);
and U3374 (N_3374,N_2187,N_1418);
or U3375 (N_3375,N_1321,N_842);
nor U3376 (N_3376,N_460,N_509);
or U3377 (N_3377,N_2217,N_1094);
nor U3378 (N_3378,N_59,N_182);
xnor U3379 (N_3379,N_2471,N_2441);
or U3380 (N_3380,N_1032,N_2149);
nor U3381 (N_3381,N_1,N_1522);
nor U3382 (N_3382,N_1467,N_1868);
or U3383 (N_3383,N_1587,N_2097);
and U3384 (N_3384,N_694,N_80);
and U3385 (N_3385,N_83,N_1806);
and U3386 (N_3386,N_921,N_1795);
xnor U3387 (N_3387,N_214,N_563);
nor U3388 (N_3388,N_1496,N_1900);
and U3389 (N_3389,N_485,N_1489);
or U3390 (N_3390,N_2041,N_1083);
and U3391 (N_3391,N_682,N_30);
nand U3392 (N_3392,N_1251,N_1749);
or U3393 (N_3393,N_1928,N_1356);
and U3394 (N_3394,N_947,N_17);
nor U3395 (N_3395,N_1367,N_493);
and U3396 (N_3396,N_215,N_1953);
nor U3397 (N_3397,N_1372,N_1819);
nor U3398 (N_3398,N_1202,N_865);
and U3399 (N_3399,N_1866,N_2019);
xnor U3400 (N_3400,N_664,N_2197);
nor U3401 (N_3401,N_776,N_419);
nor U3402 (N_3402,N_856,N_439);
xor U3403 (N_3403,N_1813,N_942);
or U3404 (N_3404,N_913,N_661);
or U3405 (N_3405,N_882,N_1883);
nor U3406 (N_3406,N_2226,N_504);
nor U3407 (N_3407,N_1965,N_1026);
or U3408 (N_3408,N_1657,N_964);
or U3409 (N_3409,N_2278,N_462);
or U3410 (N_3410,N_960,N_1194);
nor U3411 (N_3411,N_1895,N_765);
nand U3412 (N_3412,N_68,N_1171);
and U3413 (N_3413,N_1006,N_1441);
or U3414 (N_3414,N_874,N_614);
or U3415 (N_3415,N_130,N_695);
xor U3416 (N_3416,N_1208,N_903);
or U3417 (N_3417,N_653,N_2338);
and U3418 (N_3418,N_145,N_2386);
xnor U3419 (N_3419,N_211,N_916);
nor U3420 (N_3420,N_1734,N_1696);
and U3421 (N_3421,N_1433,N_1376);
xnor U3422 (N_3422,N_1675,N_411);
xnor U3423 (N_3423,N_313,N_1417);
or U3424 (N_3424,N_38,N_580);
nor U3425 (N_3425,N_1358,N_1318);
nor U3426 (N_3426,N_899,N_1693);
or U3427 (N_3427,N_1024,N_1751);
nand U3428 (N_3428,N_350,N_1977);
nor U3429 (N_3429,N_246,N_1763);
nor U3430 (N_3430,N_1049,N_724);
xnor U3431 (N_3431,N_1601,N_1997);
and U3432 (N_3432,N_1905,N_786);
and U3433 (N_3433,N_1746,N_606);
xnor U3434 (N_3434,N_558,N_782);
and U3435 (N_3435,N_552,N_778);
or U3436 (N_3436,N_360,N_2004);
and U3437 (N_3437,N_984,N_1861);
xnor U3438 (N_3438,N_1873,N_1241);
and U3439 (N_3439,N_2372,N_1674);
and U3440 (N_3440,N_2274,N_2194);
or U3441 (N_3441,N_2281,N_455);
or U3442 (N_3442,N_2040,N_1247);
or U3443 (N_3443,N_1117,N_825);
xor U3444 (N_3444,N_270,N_1894);
and U3445 (N_3445,N_1333,N_604);
or U3446 (N_3446,N_328,N_501);
or U3447 (N_3447,N_1387,N_1155);
nand U3448 (N_3448,N_2483,N_473);
nand U3449 (N_3449,N_1322,N_2494);
nand U3450 (N_3450,N_1682,N_1039);
and U3451 (N_3451,N_890,N_1113);
and U3452 (N_3452,N_678,N_1434);
nor U3453 (N_3453,N_1342,N_288);
or U3454 (N_3454,N_658,N_1670);
nor U3455 (N_3455,N_1102,N_1444);
nand U3456 (N_3456,N_1316,N_1643);
xnor U3457 (N_3457,N_549,N_955);
or U3458 (N_3458,N_287,N_2209);
xor U3459 (N_3459,N_1424,N_1028);
and U3460 (N_3460,N_433,N_1475);
xnor U3461 (N_3461,N_2195,N_1246);
nand U3462 (N_3462,N_1588,N_97);
nor U3463 (N_3463,N_2490,N_1179);
and U3464 (N_3464,N_2093,N_1146);
and U3465 (N_3465,N_551,N_813);
nand U3466 (N_3466,N_2225,N_1777);
nand U3467 (N_3467,N_802,N_1464);
and U3468 (N_3468,N_1645,N_521);
xnor U3469 (N_3469,N_2410,N_378);
nand U3470 (N_3470,N_1625,N_448);
nor U3471 (N_3471,N_1596,N_1665);
nand U3472 (N_3472,N_2137,N_2240);
nand U3473 (N_3473,N_1410,N_1043);
and U3474 (N_3474,N_930,N_1980);
nor U3475 (N_3475,N_910,N_2377);
xor U3476 (N_3476,N_888,N_1211);
nand U3477 (N_3477,N_66,N_1567);
xor U3478 (N_3478,N_1990,N_826);
xor U3479 (N_3479,N_1983,N_1851);
or U3480 (N_3480,N_1818,N_1419);
xor U3481 (N_3481,N_911,N_1862);
and U3482 (N_3482,N_2464,N_1836);
nand U3483 (N_3483,N_2208,N_2270);
or U3484 (N_3484,N_1622,N_2119);
or U3485 (N_3485,N_2292,N_698);
xor U3486 (N_3486,N_1244,N_340);
or U3487 (N_3487,N_1652,N_962);
or U3488 (N_3488,N_1526,N_85);
nand U3489 (N_3489,N_1776,N_1656);
nor U3490 (N_3490,N_2201,N_2020);
nor U3491 (N_3491,N_2295,N_1064);
nand U3492 (N_3492,N_2298,N_602);
nor U3493 (N_3493,N_976,N_705);
and U3494 (N_3494,N_1066,N_2128);
or U3495 (N_3495,N_1914,N_2255);
xor U3496 (N_3496,N_1492,N_410);
nor U3497 (N_3497,N_1252,N_925);
and U3498 (N_3498,N_1518,N_1167);
nand U3499 (N_3499,N_1910,N_2408);
nor U3500 (N_3500,N_77,N_2231);
and U3501 (N_3501,N_1334,N_2248);
nor U3502 (N_3502,N_1954,N_95);
xor U3503 (N_3503,N_2434,N_2190);
xor U3504 (N_3504,N_689,N_434);
nor U3505 (N_3505,N_1547,N_599);
and U3506 (N_3506,N_281,N_1008);
nor U3507 (N_3507,N_1022,N_933);
and U3508 (N_3508,N_300,N_692);
and U3509 (N_3509,N_2099,N_1774);
nand U3510 (N_3510,N_1839,N_607);
nor U3511 (N_3511,N_1137,N_40);
nand U3512 (N_3512,N_417,N_224);
xor U3513 (N_3513,N_1196,N_1597);
nand U3514 (N_3514,N_1699,N_1737);
nand U3515 (N_3515,N_1611,N_2465);
xnor U3516 (N_3516,N_848,N_1234);
xnor U3517 (N_3517,N_188,N_798);
or U3518 (N_3518,N_2367,N_2310);
nor U3519 (N_3519,N_380,N_342);
nor U3520 (N_3520,N_1594,N_2440);
nand U3521 (N_3521,N_2193,N_1542);
xor U3522 (N_3522,N_1266,N_532);
or U3523 (N_3523,N_1182,N_1140);
xor U3524 (N_3524,N_1499,N_878);
and U3525 (N_3525,N_2090,N_1683);
nor U3526 (N_3526,N_1503,N_1843);
or U3527 (N_3527,N_432,N_1181);
and U3528 (N_3528,N_1112,N_794);
xor U3529 (N_3529,N_494,N_245);
xor U3530 (N_3530,N_992,N_1847);
nor U3531 (N_3531,N_1469,N_591);
nor U3532 (N_3532,N_1630,N_124);
and U3533 (N_3533,N_2101,N_2469);
or U3534 (N_3534,N_1450,N_430);
nor U3535 (N_3535,N_759,N_253);
and U3536 (N_3536,N_1872,N_676);
and U3537 (N_3537,N_1096,N_1297);
xnor U3538 (N_3538,N_1724,N_255);
nand U3539 (N_3539,N_670,N_1658);
nand U3540 (N_3540,N_1402,N_2303);
xor U3541 (N_3541,N_2403,N_1554);
and U3542 (N_3542,N_119,N_81);
xnor U3543 (N_3543,N_2144,N_862);
nand U3544 (N_3544,N_1197,N_1335);
nand U3545 (N_3545,N_1207,N_483);
xor U3546 (N_3546,N_595,N_1694);
nor U3547 (N_3547,N_1076,N_718);
and U3548 (N_3548,N_1118,N_256);
or U3549 (N_3549,N_252,N_363);
or U3550 (N_3550,N_526,N_330);
xnor U3551 (N_3551,N_2246,N_2385);
nand U3552 (N_3552,N_829,N_2374);
xor U3553 (N_3553,N_2383,N_122);
or U3554 (N_3554,N_2124,N_1773);
and U3555 (N_3555,N_2070,N_1029);
xor U3556 (N_3556,N_1796,N_1224);
nand U3557 (N_3557,N_5,N_999);
nand U3558 (N_3558,N_2448,N_996);
and U3559 (N_3559,N_62,N_1790);
and U3560 (N_3560,N_2467,N_1269);
nor U3561 (N_3561,N_2265,N_1604);
and U3562 (N_3562,N_869,N_755);
xnor U3563 (N_3563,N_48,N_1306);
and U3564 (N_3564,N_2318,N_254);
and U3565 (N_3565,N_1738,N_1290);
nor U3566 (N_3566,N_528,N_2111);
nand U3567 (N_3567,N_897,N_1158);
and U3568 (N_3568,N_1880,N_1037);
or U3569 (N_3569,N_2085,N_941);
and U3570 (N_3570,N_677,N_2396);
and U3571 (N_3571,N_184,N_414);
or U3572 (N_3572,N_459,N_2094);
or U3573 (N_3573,N_1085,N_2100);
xnor U3574 (N_3574,N_2218,N_138);
nand U3575 (N_3575,N_889,N_191);
or U3576 (N_3576,N_861,N_2276);
nand U3577 (N_3577,N_1545,N_1378);
xnor U3578 (N_3578,N_200,N_893);
nor U3579 (N_3579,N_1190,N_2271);
and U3580 (N_3580,N_437,N_230);
nand U3581 (N_3581,N_1216,N_131);
nor U3582 (N_3582,N_1844,N_2202);
nor U3583 (N_3583,N_1986,N_1874);
and U3584 (N_3584,N_2112,N_1552);
nor U3585 (N_3585,N_1193,N_1936);
nand U3586 (N_3586,N_1760,N_627);
or U3587 (N_3587,N_1320,N_1038);
xnor U3588 (N_3588,N_1686,N_525);
nand U3589 (N_3589,N_2272,N_654);
nor U3590 (N_3590,N_1327,N_2493);
nand U3591 (N_3591,N_545,N_1379);
xnor U3592 (N_3592,N_43,N_1961);
and U3593 (N_3593,N_646,N_1996);
or U3594 (N_3594,N_1174,N_2316);
and U3595 (N_3595,N_2296,N_952);
nand U3596 (N_3596,N_1677,N_2332);
nand U3597 (N_3597,N_329,N_1081);
nand U3598 (N_3598,N_2261,N_2049);
nor U3599 (N_3599,N_2034,N_1409);
or U3600 (N_3600,N_121,N_1192);
nand U3601 (N_3601,N_1384,N_456);
and U3602 (N_3602,N_1591,N_743);
or U3603 (N_3603,N_887,N_824);
xor U3604 (N_3604,N_1291,N_1073);
nand U3605 (N_3605,N_1187,N_1273);
or U3606 (N_3606,N_2333,N_1579);
nand U3607 (N_3607,N_2368,N_1893);
and U3608 (N_3608,N_2064,N_1569);
nand U3609 (N_3609,N_2027,N_198);
nor U3610 (N_3610,N_51,N_2155);
or U3611 (N_3611,N_1479,N_668);
xnor U3612 (N_3612,N_52,N_610);
xor U3613 (N_3613,N_1304,N_2371);
nand U3614 (N_3614,N_2084,N_704);
xnor U3615 (N_3615,N_1491,N_735);
nand U3616 (N_3616,N_1129,N_712);
and U3617 (N_3617,N_149,N_1099);
nor U3618 (N_3618,N_643,N_385);
nand U3619 (N_3619,N_1680,N_1701);
nor U3620 (N_3620,N_488,N_870);
nor U3621 (N_3621,N_2074,N_2336);
nor U3622 (N_3622,N_463,N_334);
or U3623 (N_3623,N_2042,N_1881);
xor U3624 (N_3624,N_1810,N_2095);
or U3625 (N_3625,N_2045,N_2106);
or U3626 (N_3626,N_577,N_883);
nor U3627 (N_3627,N_1220,N_2047);
xor U3628 (N_3628,N_819,N_593);
nor U3629 (N_3629,N_180,N_1040);
and U3630 (N_3630,N_548,N_1294);
nor U3631 (N_3631,N_1041,N_1511);
nor U3632 (N_3632,N_951,N_1758);
and U3633 (N_3633,N_1742,N_1413);
nor U3634 (N_3634,N_605,N_1711);
nand U3635 (N_3635,N_1486,N_1982);
and U3636 (N_3636,N_14,N_1205);
xor U3637 (N_3637,N_1231,N_1256);
xor U3638 (N_3638,N_1245,N_994);
nand U3639 (N_3639,N_1887,N_316);
or U3640 (N_3640,N_293,N_820);
nand U3641 (N_3641,N_1176,N_146);
nor U3642 (N_3642,N_1268,N_2214);
and U3643 (N_3643,N_1080,N_2433);
and U3644 (N_3644,N_2424,N_1364);
or U3645 (N_3645,N_1947,N_2087);
xor U3646 (N_3646,N_1375,N_2172);
xnor U3647 (N_3647,N_497,N_1770);
or U3648 (N_3648,N_2001,N_1590);
nor U3649 (N_3649,N_1344,N_1736);
or U3650 (N_3650,N_2422,N_891);
or U3651 (N_3651,N_1238,N_2107);
xor U3652 (N_3652,N_92,N_837);
or U3653 (N_3653,N_1053,N_2324);
and U3654 (N_3654,N_1069,N_9);
or U3655 (N_3655,N_1687,N_2304);
and U3656 (N_3656,N_1473,N_2348);
or U3657 (N_3657,N_2170,N_934);
nand U3658 (N_3658,N_1277,N_1374);
xor U3659 (N_3659,N_1408,N_2091);
or U3660 (N_3660,N_1082,N_2140);
or U3661 (N_3661,N_1825,N_896);
and U3662 (N_3662,N_650,N_60);
nand U3663 (N_3663,N_1891,N_1801);
nand U3664 (N_3664,N_767,N_1679);
nor U3665 (N_3665,N_884,N_2309);
and U3666 (N_3666,N_520,N_1141);
or U3667 (N_3667,N_644,N_727);
and U3668 (N_3668,N_1275,N_1104);
nand U3669 (N_3669,N_2241,N_1592);
and U3670 (N_3670,N_1911,N_1867);
nand U3671 (N_3671,N_263,N_739);
nor U3672 (N_3672,N_1101,N_1715);
nor U3673 (N_3673,N_2347,N_2436);
nand U3674 (N_3674,N_1258,N_2141);
or U3675 (N_3675,N_1206,N_1743);
or U3676 (N_3676,N_1753,N_400);
nor U3677 (N_3677,N_1783,N_28);
nand U3678 (N_3678,N_2125,N_719);
nand U3679 (N_3679,N_1762,N_234);
nand U3680 (N_3680,N_1620,N_1271);
or U3681 (N_3681,N_1646,N_1942);
xnor U3682 (N_3682,N_2450,N_2335);
and U3683 (N_3683,N_267,N_2378);
or U3684 (N_3684,N_2262,N_1030);
xor U3685 (N_3685,N_685,N_2291);
and U3686 (N_3686,N_1369,N_818);
nand U3687 (N_3687,N_1684,N_1899);
nor U3688 (N_3688,N_1617,N_1815);
nand U3689 (N_3689,N_1916,N_2325);
nand U3690 (N_3690,N_1633,N_651);
and U3691 (N_3691,N_1223,N_10);
xor U3692 (N_3692,N_686,N_1703);
nor U3693 (N_3693,N_871,N_1033);
xnor U3694 (N_3694,N_2116,N_573);
and U3695 (N_3695,N_2364,N_226);
nor U3696 (N_3696,N_2250,N_1925);
nand U3697 (N_3697,N_1042,N_1556);
nor U3698 (N_3698,N_2404,N_791);
xor U3699 (N_3699,N_2239,N_1958);
nor U3700 (N_3700,N_1100,N_867);
nand U3701 (N_3701,N_1236,N_1253);
and U3702 (N_3702,N_1336,N_2337);
or U3703 (N_3703,N_1130,N_1991);
and U3704 (N_3704,N_185,N_120);
or U3705 (N_3705,N_2178,N_1314);
xor U3706 (N_3706,N_586,N_176);
and U3707 (N_3707,N_1978,N_998);
or U3708 (N_3708,N_53,N_1691);
nand U3709 (N_3709,N_249,N_590);
and U3710 (N_3710,N_1603,N_391);
xor U3711 (N_3711,N_2154,N_1820);
nand U3712 (N_3712,N_354,N_90);
xor U3713 (N_3713,N_620,N_1382);
nand U3714 (N_3714,N_1578,N_1248);
nor U3715 (N_3715,N_2447,N_409);
nand U3716 (N_3716,N_1799,N_730);
nand U3717 (N_3717,N_241,N_1195);
nor U3718 (N_3718,N_173,N_280);
nand U3719 (N_3719,N_1507,N_700);
and U3720 (N_3720,N_1015,N_31);
or U3721 (N_3721,N_2227,N_2431);
xnor U3722 (N_3722,N_2166,N_1500);
or U3723 (N_3723,N_1863,N_212);
nand U3724 (N_3724,N_2175,N_306);
nand U3725 (N_3725,N_2415,N_805);
nor U3726 (N_3726,N_502,N_1946);
nor U3727 (N_3727,N_237,N_469);
or U3728 (N_3728,N_811,N_2200);
nor U3729 (N_3729,N_476,N_1164);
or U3730 (N_3730,N_2354,N_351);
nor U3731 (N_3731,N_2159,N_1932);
nand U3732 (N_3732,N_1808,N_1415);
and U3733 (N_3733,N_1725,N_1011);
and U3734 (N_3734,N_1966,N_67);
xnor U3735 (N_3735,N_2056,N_1842);
xnor U3736 (N_3736,N_8,N_2257);
or U3737 (N_3737,N_1180,N_69);
or U3738 (N_3738,N_2179,N_839);
xnor U3739 (N_3739,N_697,N_1458);
or U3740 (N_3740,N_1605,N_1827);
and U3741 (N_3741,N_1729,N_47);
xor U3742 (N_3742,N_2110,N_1988);
nor U3743 (N_3743,N_2188,N_2294);
nor U3744 (N_3744,N_2058,N_2043);
xnor U3745 (N_3745,N_1558,N_2204);
nor U3746 (N_3746,N_2150,N_1598);
or U3747 (N_3747,N_572,N_186);
and U3748 (N_3748,N_764,N_76);
nand U3749 (N_3749,N_1555,N_713);
xnor U3750 (N_3750,N_2362,N_471);
xor U3751 (N_3751,N_643,N_1810);
or U3752 (N_3752,N_772,N_518);
xor U3753 (N_3753,N_1231,N_247);
and U3754 (N_3754,N_1528,N_2488);
nand U3755 (N_3755,N_1383,N_644);
nand U3756 (N_3756,N_878,N_2195);
xor U3757 (N_3757,N_1561,N_233);
xor U3758 (N_3758,N_1405,N_1186);
and U3759 (N_3759,N_645,N_2087);
nor U3760 (N_3760,N_643,N_2174);
nor U3761 (N_3761,N_497,N_1718);
and U3762 (N_3762,N_1490,N_1752);
and U3763 (N_3763,N_1380,N_1465);
nor U3764 (N_3764,N_394,N_410);
or U3765 (N_3765,N_2331,N_2437);
nor U3766 (N_3766,N_803,N_382);
or U3767 (N_3767,N_1064,N_724);
xor U3768 (N_3768,N_2214,N_2080);
and U3769 (N_3769,N_2026,N_2191);
xnor U3770 (N_3770,N_1895,N_2302);
nand U3771 (N_3771,N_614,N_1698);
and U3772 (N_3772,N_773,N_2249);
nand U3773 (N_3773,N_1278,N_1784);
and U3774 (N_3774,N_259,N_1658);
xnor U3775 (N_3775,N_1495,N_1378);
nand U3776 (N_3776,N_1133,N_665);
nor U3777 (N_3777,N_595,N_1229);
xor U3778 (N_3778,N_1767,N_1840);
or U3779 (N_3779,N_1669,N_832);
xor U3780 (N_3780,N_616,N_555);
and U3781 (N_3781,N_1391,N_1867);
and U3782 (N_3782,N_1047,N_1309);
xnor U3783 (N_3783,N_116,N_371);
xnor U3784 (N_3784,N_2203,N_116);
nand U3785 (N_3785,N_936,N_1058);
xor U3786 (N_3786,N_784,N_1499);
xnor U3787 (N_3787,N_653,N_423);
xnor U3788 (N_3788,N_941,N_810);
nand U3789 (N_3789,N_568,N_1630);
xnor U3790 (N_3790,N_1367,N_2288);
xor U3791 (N_3791,N_1229,N_646);
and U3792 (N_3792,N_171,N_675);
and U3793 (N_3793,N_884,N_216);
nand U3794 (N_3794,N_1288,N_324);
nor U3795 (N_3795,N_976,N_1949);
xor U3796 (N_3796,N_1392,N_1943);
nand U3797 (N_3797,N_1751,N_2430);
and U3798 (N_3798,N_1174,N_401);
xnor U3799 (N_3799,N_2487,N_1561);
and U3800 (N_3800,N_1952,N_1022);
xnor U3801 (N_3801,N_867,N_2044);
nor U3802 (N_3802,N_1818,N_1179);
xor U3803 (N_3803,N_820,N_2002);
or U3804 (N_3804,N_1372,N_491);
xor U3805 (N_3805,N_938,N_1310);
or U3806 (N_3806,N_2266,N_2014);
or U3807 (N_3807,N_1034,N_2003);
nor U3808 (N_3808,N_2280,N_2395);
nor U3809 (N_3809,N_768,N_1235);
or U3810 (N_3810,N_1543,N_1825);
nor U3811 (N_3811,N_839,N_1558);
nor U3812 (N_3812,N_177,N_40);
nor U3813 (N_3813,N_1619,N_383);
nand U3814 (N_3814,N_805,N_1293);
nor U3815 (N_3815,N_1313,N_776);
nor U3816 (N_3816,N_1877,N_1906);
and U3817 (N_3817,N_1341,N_15);
nor U3818 (N_3818,N_368,N_2120);
nand U3819 (N_3819,N_1805,N_795);
xor U3820 (N_3820,N_941,N_1002);
and U3821 (N_3821,N_1223,N_1520);
and U3822 (N_3822,N_2402,N_1449);
or U3823 (N_3823,N_1777,N_1779);
nor U3824 (N_3824,N_2469,N_788);
nand U3825 (N_3825,N_2259,N_1341);
nand U3826 (N_3826,N_911,N_1508);
nand U3827 (N_3827,N_2106,N_2377);
and U3828 (N_3828,N_493,N_744);
xnor U3829 (N_3829,N_293,N_2011);
nand U3830 (N_3830,N_1057,N_593);
and U3831 (N_3831,N_282,N_1978);
nor U3832 (N_3832,N_853,N_2459);
and U3833 (N_3833,N_792,N_1652);
nor U3834 (N_3834,N_2394,N_1256);
nand U3835 (N_3835,N_686,N_1627);
and U3836 (N_3836,N_663,N_2375);
or U3837 (N_3837,N_405,N_2113);
and U3838 (N_3838,N_2316,N_2133);
and U3839 (N_3839,N_2015,N_1503);
nor U3840 (N_3840,N_1035,N_226);
nor U3841 (N_3841,N_1362,N_200);
nand U3842 (N_3842,N_657,N_1126);
xnor U3843 (N_3843,N_712,N_1159);
xor U3844 (N_3844,N_775,N_363);
or U3845 (N_3845,N_687,N_904);
nor U3846 (N_3846,N_1058,N_1984);
nand U3847 (N_3847,N_1480,N_1290);
nor U3848 (N_3848,N_545,N_1457);
nand U3849 (N_3849,N_645,N_455);
or U3850 (N_3850,N_599,N_851);
nor U3851 (N_3851,N_1075,N_776);
nor U3852 (N_3852,N_637,N_1254);
nand U3853 (N_3853,N_84,N_1343);
nand U3854 (N_3854,N_688,N_1923);
or U3855 (N_3855,N_1590,N_1915);
nand U3856 (N_3856,N_306,N_1782);
xnor U3857 (N_3857,N_211,N_828);
nor U3858 (N_3858,N_1064,N_2302);
nand U3859 (N_3859,N_309,N_1462);
nor U3860 (N_3860,N_2096,N_1916);
xnor U3861 (N_3861,N_208,N_250);
or U3862 (N_3862,N_1701,N_2227);
nand U3863 (N_3863,N_1298,N_932);
nand U3864 (N_3864,N_1643,N_2225);
or U3865 (N_3865,N_1348,N_386);
and U3866 (N_3866,N_2121,N_799);
or U3867 (N_3867,N_1859,N_2288);
and U3868 (N_3868,N_165,N_1167);
nor U3869 (N_3869,N_418,N_2277);
nor U3870 (N_3870,N_1608,N_963);
or U3871 (N_3871,N_879,N_1403);
and U3872 (N_3872,N_952,N_37);
and U3873 (N_3873,N_979,N_1578);
and U3874 (N_3874,N_2259,N_2188);
or U3875 (N_3875,N_1669,N_1163);
nand U3876 (N_3876,N_1309,N_1920);
nor U3877 (N_3877,N_1839,N_155);
or U3878 (N_3878,N_348,N_2034);
nand U3879 (N_3879,N_922,N_2335);
nand U3880 (N_3880,N_1627,N_2482);
and U3881 (N_3881,N_1889,N_1037);
and U3882 (N_3882,N_2102,N_1625);
xor U3883 (N_3883,N_2050,N_51);
nor U3884 (N_3884,N_584,N_2295);
xnor U3885 (N_3885,N_1876,N_1977);
nand U3886 (N_3886,N_1212,N_1815);
nor U3887 (N_3887,N_96,N_2256);
and U3888 (N_3888,N_2428,N_2457);
nor U3889 (N_3889,N_1865,N_341);
nand U3890 (N_3890,N_683,N_2438);
or U3891 (N_3891,N_65,N_2405);
and U3892 (N_3892,N_621,N_1676);
xnor U3893 (N_3893,N_2239,N_591);
nand U3894 (N_3894,N_1097,N_1791);
or U3895 (N_3895,N_1838,N_1864);
or U3896 (N_3896,N_1455,N_2039);
nand U3897 (N_3897,N_241,N_9);
and U3898 (N_3898,N_1398,N_2401);
nor U3899 (N_3899,N_793,N_2443);
xor U3900 (N_3900,N_718,N_1152);
nand U3901 (N_3901,N_533,N_2196);
and U3902 (N_3902,N_317,N_1533);
and U3903 (N_3903,N_206,N_593);
and U3904 (N_3904,N_548,N_2042);
nand U3905 (N_3905,N_1040,N_542);
xnor U3906 (N_3906,N_417,N_1045);
nor U3907 (N_3907,N_454,N_2492);
xnor U3908 (N_3908,N_253,N_689);
nand U3909 (N_3909,N_1808,N_205);
nor U3910 (N_3910,N_918,N_1638);
nor U3911 (N_3911,N_1873,N_1960);
nand U3912 (N_3912,N_1162,N_63);
nor U3913 (N_3913,N_2140,N_2333);
nor U3914 (N_3914,N_585,N_1827);
nand U3915 (N_3915,N_796,N_281);
or U3916 (N_3916,N_103,N_2323);
or U3917 (N_3917,N_2388,N_781);
xnor U3918 (N_3918,N_1161,N_662);
and U3919 (N_3919,N_2242,N_1364);
nor U3920 (N_3920,N_1893,N_1022);
or U3921 (N_3921,N_601,N_1817);
and U3922 (N_3922,N_1875,N_1138);
and U3923 (N_3923,N_1945,N_1089);
nor U3924 (N_3924,N_1904,N_2332);
nor U3925 (N_3925,N_1749,N_1800);
or U3926 (N_3926,N_1649,N_163);
nand U3927 (N_3927,N_1367,N_1494);
xor U3928 (N_3928,N_1505,N_1602);
or U3929 (N_3929,N_2328,N_111);
nor U3930 (N_3930,N_1893,N_1261);
nor U3931 (N_3931,N_417,N_1342);
xor U3932 (N_3932,N_239,N_1499);
xor U3933 (N_3933,N_478,N_1929);
or U3934 (N_3934,N_1618,N_1741);
nor U3935 (N_3935,N_1247,N_401);
or U3936 (N_3936,N_104,N_2053);
or U3937 (N_3937,N_1995,N_205);
nand U3938 (N_3938,N_2195,N_490);
nand U3939 (N_3939,N_1299,N_933);
nor U3940 (N_3940,N_1299,N_278);
nor U3941 (N_3941,N_1285,N_1506);
and U3942 (N_3942,N_989,N_1342);
nand U3943 (N_3943,N_2493,N_1071);
nand U3944 (N_3944,N_2189,N_1430);
xnor U3945 (N_3945,N_1145,N_980);
nor U3946 (N_3946,N_238,N_1875);
nor U3947 (N_3947,N_1899,N_477);
xor U3948 (N_3948,N_799,N_1679);
xor U3949 (N_3949,N_723,N_1813);
or U3950 (N_3950,N_387,N_391);
nor U3951 (N_3951,N_1159,N_2217);
xnor U3952 (N_3952,N_1409,N_2049);
or U3953 (N_3953,N_2127,N_2157);
nor U3954 (N_3954,N_2069,N_808);
nor U3955 (N_3955,N_1564,N_2095);
or U3956 (N_3956,N_1256,N_1872);
nand U3957 (N_3957,N_0,N_544);
xnor U3958 (N_3958,N_718,N_814);
and U3959 (N_3959,N_545,N_765);
nor U3960 (N_3960,N_2286,N_238);
nor U3961 (N_3961,N_774,N_255);
or U3962 (N_3962,N_1111,N_2291);
nor U3963 (N_3963,N_832,N_1660);
and U3964 (N_3964,N_323,N_476);
xor U3965 (N_3965,N_1626,N_1033);
xor U3966 (N_3966,N_2025,N_2079);
nor U3967 (N_3967,N_161,N_849);
or U3968 (N_3968,N_914,N_1671);
or U3969 (N_3969,N_1221,N_1454);
and U3970 (N_3970,N_905,N_1237);
xor U3971 (N_3971,N_1792,N_398);
nor U3972 (N_3972,N_986,N_1841);
xnor U3973 (N_3973,N_1018,N_882);
nor U3974 (N_3974,N_842,N_1778);
nor U3975 (N_3975,N_1482,N_2313);
nor U3976 (N_3976,N_1484,N_2063);
and U3977 (N_3977,N_295,N_1961);
or U3978 (N_3978,N_993,N_2350);
nand U3979 (N_3979,N_2141,N_283);
and U3980 (N_3980,N_1569,N_1637);
xor U3981 (N_3981,N_1685,N_2040);
nor U3982 (N_3982,N_2496,N_1297);
or U3983 (N_3983,N_1024,N_1915);
or U3984 (N_3984,N_502,N_1520);
and U3985 (N_3985,N_1034,N_2030);
nand U3986 (N_3986,N_1497,N_203);
xnor U3987 (N_3987,N_1268,N_1707);
nand U3988 (N_3988,N_949,N_520);
and U3989 (N_3989,N_2006,N_1532);
xor U3990 (N_3990,N_2359,N_1073);
or U3991 (N_3991,N_1140,N_347);
xor U3992 (N_3992,N_1967,N_2226);
or U3993 (N_3993,N_1301,N_1688);
or U3994 (N_3994,N_1997,N_936);
or U3995 (N_3995,N_612,N_2035);
nor U3996 (N_3996,N_1757,N_228);
nor U3997 (N_3997,N_1465,N_1786);
nor U3998 (N_3998,N_1954,N_36);
nand U3999 (N_3999,N_1488,N_1757);
xor U4000 (N_4000,N_1996,N_277);
and U4001 (N_4001,N_585,N_884);
nor U4002 (N_4002,N_698,N_753);
and U4003 (N_4003,N_1775,N_1328);
nand U4004 (N_4004,N_279,N_1237);
xor U4005 (N_4005,N_1145,N_856);
or U4006 (N_4006,N_65,N_1175);
xor U4007 (N_4007,N_973,N_1504);
nand U4008 (N_4008,N_541,N_2205);
xnor U4009 (N_4009,N_785,N_2328);
xnor U4010 (N_4010,N_1180,N_437);
and U4011 (N_4011,N_2288,N_1097);
nand U4012 (N_4012,N_381,N_1870);
nor U4013 (N_4013,N_1084,N_1564);
xnor U4014 (N_4014,N_361,N_244);
nand U4015 (N_4015,N_1162,N_631);
nand U4016 (N_4016,N_1835,N_569);
xnor U4017 (N_4017,N_1979,N_2480);
nand U4018 (N_4018,N_294,N_732);
and U4019 (N_4019,N_266,N_473);
nand U4020 (N_4020,N_271,N_1990);
nor U4021 (N_4021,N_1812,N_1318);
or U4022 (N_4022,N_583,N_2362);
and U4023 (N_4023,N_1071,N_1916);
nor U4024 (N_4024,N_2456,N_2432);
nor U4025 (N_4025,N_774,N_2345);
or U4026 (N_4026,N_1568,N_909);
or U4027 (N_4027,N_350,N_1329);
and U4028 (N_4028,N_2285,N_1125);
nand U4029 (N_4029,N_2038,N_2124);
xnor U4030 (N_4030,N_2223,N_204);
nor U4031 (N_4031,N_1995,N_689);
nand U4032 (N_4032,N_2268,N_2405);
nor U4033 (N_4033,N_831,N_2122);
nor U4034 (N_4034,N_525,N_1765);
or U4035 (N_4035,N_1537,N_1694);
and U4036 (N_4036,N_2101,N_961);
and U4037 (N_4037,N_1794,N_1175);
nor U4038 (N_4038,N_2240,N_137);
xor U4039 (N_4039,N_1113,N_442);
nor U4040 (N_4040,N_2407,N_1453);
or U4041 (N_4041,N_855,N_663);
nor U4042 (N_4042,N_2451,N_2012);
nand U4043 (N_4043,N_1579,N_1193);
nand U4044 (N_4044,N_1032,N_443);
nand U4045 (N_4045,N_817,N_858);
nand U4046 (N_4046,N_2197,N_884);
nand U4047 (N_4047,N_2110,N_439);
xnor U4048 (N_4048,N_2175,N_488);
nand U4049 (N_4049,N_1810,N_1315);
nor U4050 (N_4050,N_68,N_599);
nand U4051 (N_4051,N_2133,N_1938);
and U4052 (N_4052,N_1096,N_828);
nor U4053 (N_4053,N_587,N_313);
xor U4054 (N_4054,N_1342,N_604);
and U4055 (N_4055,N_2360,N_1328);
and U4056 (N_4056,N_1643,N_184);
nand U4057 (N_4057,N_340,N_1637);
and U4058 (N_4058,N_2413,N_2447);
xor U4059 (N_4059,N_2324,N_366);
xor U4060 (N_4060,N_338,N_1071);
xor U4061 (N_4061,N_43,N_2069);
and U4062 (N_4062,N_231,N_2289);
and U4063 (N_4063,N_1813,N_250);
nor U4064 (N_4064,N_637,N_1687);
or U4065 (N_4065,N_1587,N_2261);
and U4066 (N_4066,N_315,N_372);
nor U4067 (N_4067,N_2089,N_760);
nand U4068 (N_4068,N_422,N_1190);
nor U4069 (N_4069,N_1809,N_86);
or U4070 (N_4070,N_2174,N_463);
or U4071 (N_4071,N_1775,N_1995);
xor U4072 (N_4072,N_2177,N_1929);
and U4073 (N_4073,N_1383,N_1977);
nor U4074 (N_4074,N_2426,N_1853);
xnor U4075 (N_4075,N_889,N_2117);
nor U4076 (N_4076,N_963,N_439);
and U4077 (N_4077,N_2216,N_1665);
xor U4078 (N_4078,N_714,N_168);
nor U4079 (N_4079,N_1598,N_1478);
xnor U4080 (N_4080,N_2415,N_2497);
or U4081 (N_4081,N_629,N_622);
or U4082 (N_4082,N_1135,N_1161);
nand U4083 (N_4083,N_1517,N_1845);
and U4084 (N_4084,N_2042,N_898);
nand U4085 (N_4085,N_1901,N_380);
xnor U4086 (N_4086,N_1494,N_130);
or U4087 (N_4087,N_1741,N_2370);
and U4088 (N_4088,N_336,N_2369);
or U4089 (N_4089,N_115,N_1965);
and U4090 (N_4090,N_2444,N_2342);
nand U4091 (N_4091,N_705,N_381);
nand U4092 (N_4092,N_141,N_797);
or U4093 (N_4093,N_2096,N_1076);
or U4094 (N_4094,N_2389,N_1476);
xnor U4095 (N_4095,N_1396,N_388);
and U4096 (N_4096,N_88,N_1886);
nor U4097 (N_4097,N_1721,N_1897);
nand U4098 (N_4098,N_442,N_1635);
nor U4099 (N_4099,N_339,N_1086);
or U4100 (N_4100,N_2373,N_1413);
nand U4101 (N_4101,N_164,N_1963);
or U4102 (N_4102,N_2244,N_1471);
and U4103 (N_4103,N_1873,N_411);
and U4104 (N_4104,N_2113,N_962);
and U4105 (N_4105,N_1381,N_184);
xnor U4106 (N_4106,N_1020,N_1478);
and U4107 (N_4107,N_1746,N_187);
or U4108 (N_4108,N_1637,N_903);
or U4109 (N_4109,N_2415,N_47);
or U4110 (N_4110,N_646,N_1571);
nor U4111 (N_4111,N_133,N_1637);
or U4112 (N_4112,N_2324,N_1615);
or U4113 (N_4113,N_2277,N_1993);
nand U4114 (N_4114,N_794,N_760);
xnor U4115 (N_4115,N_662,N_2368);
or U4116 (N_4116,N_951,N_2292);
nand U4117 (N_4117,N_1877,N_47);
nand U4118 (N_4118,N_1389,N_1022);
nand U4119 (N_4119,N_761,N_1948);
and U4120 (N_4120,N_1241,N_465);
and U4121 (N_4121,N_1613,N_289);
xor U4122 (N_4122,N_1076,N_115);
nand U4123 (N_4123,N_677,N_1875);
nor U4124 (N_4124,N_1487,N_778);
nor U4125 (N_4125,N_244,N_915);
xnor U4126 (N_4126,N_761,N_667);
nor U4127 (N_4127,N_1493,N_1045);
nor U4128 (N_4128,N_335,N_2474);
or U4129 (N_4129,N_284,N_2403);
or U4130 (N_4130,N_261,N_1347);
nand U4131 (N_4131,N_1845,N_588);
nor U4132 (N_4132,N_761,N_2138);
xnor U4133 (N_4133,N_2489,N_1945);
nand U4134 (N_4134,N_2274,N_792);
xor U4135 (N_4135,N_2105,N_1593);
or U4136 (N_4136,N_1212,N_746);
nor U4137 (N_4137,N_1257,N_2219);
xnor U4138 (N_4138,N_756,N_683);
and U4139 (N_4139,N_127,N_2299);
xnor U4140 (N_4140,N_306,N_727);
nor U4141 (N_4141,N_2449,N_852);
xor U4142 (N_4142,N_1937,N_327);
or U4143 (N_4143,N_2433,N_594);
or U4144 (N_4144,N_471,N_929);
and U4145 (N_4145,N_783,N_170);
xnor U4146 (N_4146,N_959,N_2024);
nand U4147 (N_4147,N_1026,N_2258);
nor U4148 (N_4148,N_1204,N_269);
and U4149 (N_4149,N_768,N_1830);
nor U4150 (N_4150,N_1868,N_1795);
nor U4151 (N_4151,N_2418,N_2314);
or U4152 (N_4152,N_262,N_1699);
nor U4153 (N_4153,N_228,N_1422);
xor U4154 (N_4154,N_200,N_753);
xnor U4155 (N_4155,N_2183,N_2313);
and U4156 (N_4156,N_775,N_339);
nand U4157 (N_4157,N_836,N_2196);
nand U4158 (N_4158,N_1774,N_333);
or U4159 (N_4159,N_1851,N_560);
nand U4160 (N_4160,N_1110,N_1238);
or U4161 (N_4161,N_665,N_2328);
or U4162 (N_4162,N_1617,N_1242);
and U4163 (N_4163,N_1849,N_242);
nand U4164 (N_4164,N_521,N_2128);
nor U4165 (N_4165,N_357,N_2411);
or U4166 (N_4166,N_132,N_40);
or U4167 (N_4167,N_194,N_2194);
nor U4168 (N_4168,N_507,N_70);
or U4169 (N_4169,N_1306,N_2163);
or U4170 (N_4170,N_448,N_290);
nor U4171 (N_4171,N_1982,N_1307);
nor U4172 (N_4172,N_1012,N_0);
nand U4173 (N_4173,N_51,N_778);
and U4174 (N_4174,N_780,N_1459);
and U4175 (N_4175,N_529,N_882);
xnor U4176 (N_4176,N_2384,N_599);
or U4177 (N_4177,N_1258,N_952);
xnor U4178 (N_4178,N_678,N_1317);
nor U4179 (N_4179,N_833,N_1704);
or U4180 (N_4180,N_721,N_2263);
xor U4181 (N_4181,N_1074,N_872);
and U4182 (N_4182,N_286,N_1719);
xnor U4183 (N_4183,N_1535,N_1525);
or U4184 (N_4184,N_40,N_390);
or U4185 (N_4185,N_778,N_2432);
or U4186 (N_4186,N_868,N_1821);
nand U4187 (N_4187,N_787,N_475);
nand U4188 (N_4188,N_1819,N_2135);
nand U4189 (N_4189,N_2157,N_113);
and U4190 (N_4190,N_1751,N_172);
and U4191 (N_4191,N_1728,N_9);
and U4192 (N_4192,N_459,N_1981);
or U4193 (N_4193,N_701,N_341);
nand U4194 (N_4194,N_2405,N_1577);
or U4195 (N_4195,N_991,N_1797);
or U4196 (N_4196,N_151,N_2361);
and U4197 (N_4197,N_2399,N_2310);
nor U4198 (N_4198,N_169,N_1818);
nand U4199 (N_4199,N_1554,N_714);
nand U4200 (N_4200,N_1725,N_1391);
nand U4201 (N_4201,N_2317,N_783);
and U4202 (N_4202,N_332,N_1134);
nor U4203 (N_4203,N_1862,N_614);
nor U4204 (N_4204,N_1525,N_1518);
nor U4205 (N_4205,N_1137,N_2192);
nand U4206 (N_4206,N_1741,N_172);
nand U4207 (N_4207,N_2051,N_1828);
nor U4208 (N_4208,N_1860,N_827);
xnor U4209 (N_4209,N_2444,N_1017);
nand U4210 (N_4210,N_1943,N_306);
or U4211 (N_4211,N_1369,N_2023);
nor U4212 (N_4212,N_2215,N_2285);
nand U4213 (N_4213,N_1069,N_2126);
and U4214 (N_4214,N_306,N_1234);
or U4215 (N_4215,N_1177,N_2143);
or U4216 (N_4216,N_1266,N_1344);
nor U4217 (N_4217,N_2347,N_241);
nand U4218 (N_4218,N_1949,N_775);
xor U4219 (N_4219,N_1710,N_1695);
nor U4220 (N_4220,N_66,N_1064);
xnor U4221 (N_4221,N_414,N_1232);
or U4222 (N_4222,N_1045,N_1688);
nand U4223 (N_4223,N_2086,N_1839);
and U4224 (N_4224,N_349,N_1801);
nor U4225 (N_4225,N_2395,N_713);
nand U4226 (N_4226,N_1899,N_2067);
nor U4227 (N_4227,N_1047,N_1069);
xnor U4228 (N_4228,N_364,N_2333);
nand U4229 (N_4229,N_866,N_1315);
or U4230 (N_4230,N_1253,N_236);
xor U4231 (N_4231,N_83,N_2191);
and U4232 (N_4232,N_2354,N_1855);
and U4233 (N_4233,N_429,N_1316);
and U4234 (N_4234,N_252,N_546);
nor U4235 (N_4235,N_996,N_28);
or U4236 (N_4236,N_2381,N_2051);
nor U4237 (N_4237,N_828,N_1743);
xnor U4238 (N_4238,N_1485,N_2001);
and U4239 (N_4239,N_499,N_360);
nand U4240 (N_4240,N_283,N_19);
or U4241 (N_4241,N_1117,N_562);
xor U4242 (N_4242,N_1223,N_1434);
nor U4243 (N_4243,N_2243,N_1994);
and U4244 (N_4244,N_497,N_1935);
xnor U4245 (N_4245,N_1873,N_1159);
and U4246 (N_4246,N_1417,N_1655);
and U4247 (N_4247,N_723,N_795);
xor U4248 (N_4248,N_708,N_1335);
xor U4249 (N_4249,N_1676,N_848);
nor U4250 (N_4250,N_1410,N_1752);
nor U4251 (N_4251,N_74,N_1165);
and U4252 (N_4252,N_2247,N_1071);
nor U4253 (N_4253,N_305,N_464);
xnor U4254 (N_4254,N_2456,N_2119);
xor U4255 (N_4255,N_564,N_339);
xor U4256 (N_4256,N_2391,N_586);
nor U4257 (N_4257,N_23,N_705);
nor U4258 (N_4258,N_1368,N_799);
or U4259 (N_4259,N_2394,N_9);
and U4260 (N_4260,N_2059,N_2371);
xor U4261 (N_4261,N_2311,N_166);
nand U4262 (N_4262,N_1773,N_601);
and U4263 (N_4263,N_1471,N_1945);
xor U4264 (N_4264,N_32,N_1130);
nor U4265 (N_4265,N_1972,N_1003);
nor U4266 (N_4266,N_2366,N_2153);
and U4267 (N_4267,N_190,N_2370);
nor U4268 (N_4268,N_1437,N_2102);
or U4269 (N_4269,N_428,N_1455);
nor U4270 (N_4270,N_1567,N_37);
and U4271 (N_4271,N_2202,N_767);
or U4272 (N_4272,N_2429,N_1146);
nand U4273 (N_4273,N_2232,N_305);
and U4274 (N_4274,N_1258,N_1830);
nand U4275 (N_4275,N_2349,N_1707);
xor U4276 (N_4276,N_455,N_787);
xor U4277 (N_4277,N_350,N_1702);
xnor U4278 (N_4278,N_2054,N_1837);
nor U4279 (N_4279,N_1219,N_1784);
and U4280 (N_4280,N_707,N_304);
nand U4281 (N_4281,N_2260,N_1861);
and U4282 (N_4282,N_676,N_1589);
nand U4283 (N_4283,N_1243,N_1538);
and U4284 (N_4284,N_1432,N_109);
nor U4285 (N_4285,N_1613,N_1713);
xnor U4286 (N_4286,N_611,N_1199);
or U4287 (N_4287,N_1570,N_1672);
xor U4288 (N_4288,N_2079,N_1256);
nor U4289 (N_4289,N_595,N_2074);
and U4290 (N_4290,N_1882,N_1345);
nand U4291 (N_4291,N_2081,N_173);
or U4292 (N_4292,N_402,N_1611);
or U4293 (N_4293,N_147,N_2073);
nor U4294 (N_4294,N_1223,N_2045);
nor U4295 (N_4295,N_1967,N_861);
nor U4296 (N_4296,N_1754,N_907);
nor U4297 (N_4297,N_2197,N_2170);
nand U4298 (N_4298,N_1505,N_2170);
xnor U4299 (N_4299,N_138,N_1581);
and U4300 (N_4300,N_1436,N_2471);
nor U4301 (N_4301,N_2024,N_2492);
and U4302 (N_4302,N_540,N_1384);
and U4303 (N_4303,N_725,N_917);
nand U4304 (N_4304,N_1053,N_424);
nand U4305 (N_4305,N_2236,N_1618);
nand U4306 (N_4306,N_1342,N_1608);
and U4307 (N_4307,N_1940,N_2460);
and U4308 (N_4308,N_1573,N_2493);
and U4309 (N_4309,N_696,N_377);
xor U4310 (N_4310,N_2039,N_1300);
nor U4311 (N_4311,N_27,N_2304);
xor U4312 (N_4312,N_1836,N_1136);
nand U4313 (N_4313,N_37,N_86);
nor U4314 (N_4314,N_757,N_1031);
nor U4315 (N_4315,N_2316,N_1530);
and U4316 (N_4316,N_2029,N_2147);
xor U4317 (N_4317,N_2260,N_2210);
nor U4318 (N_4318,N_2338,N_1059);
or U4319 (N_4319,N_525,N_1919);
or U4320 (N_4320,N_1743,N_2169);
nor U4321 (N_4321,N_1851,N_310);
or U4322 (N_4322,N_2480,N_2322);
and U4323 (N_4323,N_2252,N_2415);
or U4324 (N_4324,N_2447,N_988);
nand U4325 (N_4325,N_1494,N_747);
xnor U4326 (N_4326,N_1738,N_273);
and U4327 (N_4327,N_1490,N_777);
or U4328 (N_4328,N_2093,N_1437);
and U4329 (N_4329,N_135,N_1091);
nor U4330 (N_4330,N_1051,N_1617);
and U4331 (N_4331,N_2449,N_1215);
nand U4332 (N_4332,N_1597,N_331);
nand U4333 (N_4333,N_545,N_1123);
and U4334 (N_4334,N_1712,N_888);
nor U4335 (N_4335,N_579,N_395);
nand U4336 (N_4336,N_1499,N_2133);
xnor U4337 (N_4337,N_708,N_1126);
nor U4338 (N_4338,N_1244,N_2260);
and U4339 (N_4339,N_1779,N_1288);
and U4340 (N_4340,N_2410,N_2382);
nand U4341 (N_4341,N_79,N_323);
nor U4342 (N_4342,N_549,N_1622);
or U4343 (N_4343,N_541,N_520);
and U4344 (N_4344,N_1641,N_2107);
and U4345 (N_4345,N_1369,N_774);
xnor U4346 (N_4346,N_1143,N_1618);
nor U4347 (N_4347,N_837,N_2112);
and U4348 (N_4348,N_1425,N_2073);
nand U4349 (N_4349,N_110,N_89);
or U4350 (N_4350,N_385,N_316);
or U4351 (N_4351,N_416,N_31);
nor U4352 (N_4352,N_209,N_1487);
xor U4353 (N_4353,N_886,N_2498);
nor U4354 (N_4354,N_130,N_121);
nor U4355 (N_4355,N_917,N_1246);
nor U4356 (N_4356,N_1903,N_1148);
nor U4357 (N_4357,N_1917,N_2192);
nor U4358 (N_4358,N_1158,N_926);
nand U4359 (N_4359,N_892,N_972);
and U4360 (N_4360,N_1783,N_1566);
and U4361 (N_4361,N_1329,N_679);
and U4362 (N_4362,N_1771,N_1521);
nand U4363 (N_4363,N_1395,N_405);
and U4364 (N_4364,N_1523,N_2127);
xnor U4365 (N_4365,N_1487,N_320);
nand U4366 (N_4366,N_1102,N_1212);
or U4367 (N_4367,N_2224,N_1969);
nor U4368 (N_4368,N_1949,N_1055);
nand U4369 (N_4369,N_1569,N_2254);
and U4370 (N_4370,N_1525,N_618);
nand U4371 (N_4371,N_1391,N_684);
or U4372 (N_4372,N_839,N_1469);
nor U4373 (N_4373,N_747,N_2319);
or U4374 (N_4374,N_110,N_1830);
or U4375 (N_4375,N_2371,N_2246);
or U4376 (N_4376,N_2272,N_1098);
or U4377 (N_4377,N_2439,N_439);
xor U4378 (N_4378,N_1853,N_195);
xnor U4379 (N_4379,N_1336,N_1248);
nand U4380 (N_4380,N_440,N_661);
xor U4381 (N_4381,N_1434,N_1257);
or U4382 (N_4382,N_1461,N_471);
nor U4383 (N_4383,N_1602,N_259);
nand U4384 (N_4384,N_1143,N_16);
nand U4385 (N_4385,N_814,N_1776);
xnor U4386 (N_4386,N_182,N_1672);
and U4387 (N_4387,N_1453,N_552);
xor U4388 (N_4388,N_2387,N_1879);
or U4389 (N_4389,N_2189,N_298);
xnor U4390 (N_4390,N_1454,N_1672);
nor U4391 (N_4391,N_855,N_1922);
or U4392 (N_4392,N_1672,N_1769);
xor U4393 (N_4393,N_1393,N_1020);
or U4394 (N_4394,N_794,N_1179);
nor U4395 (N_4395,N_1505,N_2233);
nor U4396 (N_4396,N_2219,N_845);
nor U4397 (N_4397,N_87,N_183);
nor U4398 (N_4398,N_983,N_2454);
nor U4399 (N_4399,N_1534,N_382);
xor U4400 (N_4400,N_1146,N_1691);
nand U4401 (N_4401,N_8,N_944);
and U4402 (N_4402,N_53,N_476);
nor U4403 (N_4403,N_2,N_1320);
or U4404 (N_4404,N_2351,N_631);
nor U4405 (N_4405,N_1783,N_939);
or U4406 (N_4406,N_683,N_972);
xnor U4407 (N_4407,N_1959,N_980);
and U4408 (N_4408,N_178,N_1441);
nor U4409 (N_4409,N_2009,N_1497);
or U4410 (N_4410,N_936,N_2217);
nor U4411 (N_4411,N_172,N_1755);
and U4412 (N_4412,N_2149,N_702);
and U4413 (N_4413,N_1951,N_1099);
or U4414 (N_4414,N_1404,N_1432);
nor U4415 (N_4415,N_2421,N_385);
or U4416 (N_4416,N_1843,N_2492);
nand U4417 (N_4417,N_1700,N_2279);
and U4418 (N_4418,N_861,N_354);
nand U4419 (N_4419,N_173,N_931);
and U4420 (N_4420,N_798,N_1696);
nand U4421 (N_4421,N_2416,N_903);
nor U4422 (N_4422,N_1145,N_2084);
xnor U4423 (N_4423,N_435,N_325);
or U4424 (N_4424,N_1491,N_1828);
and U4425 (N_4425,N_1160,N_1390);
and U4426 (N_4426,N_928,N_629);
nand U4427 (N_4427,N_143,N_1425);
nand U4428 (N_4428,N_1763,N_1317);
nor U4429 (N_4429,N_428,N_1490);
nand U4430 (N_4430,N_2116,N_112);
nor U4431 (N_4431,N_1074,N_879);
nand U4432 (N_4432,N_71,N_1718);
xor U4433 (N_4433,N_1720,N_987);
nor U4434 (N_4434,N_1149,N_1614);
nor U4435 (N_4435,N_2335,N_1916);
xnor U4436 (N_4436,N_1772,N_1610);
nor U4437 (N_4437,N_630,N_876);
nor U4438 (N_4438,N_1614,N_2040);
nand U4439 (N_4439,N_937,N_487);
and U4440 (N_4440,N_847,N_2072);
and U4441 (N_4441,N_1109,N_1552);
nor U4442 (N_4442,N_2328,N_1305);
xnor U4443 (N_4443,N_569,N_1390);
or U4444 (N_4444,N_806,N_490);
and U4445 (N_4445,N_1601,N_17);
nor U4446 (N_4446,N_750,N_2217);
nor U4447 (N_4447,N_2376,N_1704);
and U4448 (N_4448,N_2209,N_1727);
nand U4449 (N_4449,N_916,N_2425);
nor U4450 (N_4450,N_473,N_290);
nor U4451 (N_4451,N_645,N_392);
nand U4452 (N_4452,N_1115,N_456);
nand U4453 (N_4453,N_2436,N_2306);
or U4454 (N_4454,N_1868,N_538);
and U4455 (N_4455,N_1240,N_1280);
or U4456 (N_4456,N_210,N_459);
or U4457 (N_4457,N_958,N_1509);
or U4458 (N_4458,N_553,N_683);
or U4459 (N_4459,N_1583,N_905);
and U4460 (N_4460,N_2358,N_2280);
nor U4461 (N_4461,N_2053,N_247);
nor U4462 (N_4462,N_602,N_1629);
nand U4463 (N_4463,N_1873,N_2268);
nand U4464 (N_4464,N_2180,N_126);
or U4465 (N_4465,N_1473,N_1168);
or U4466 (N_4466,N_2391,N_972);
or U4467 (N_4467,N_2168,N_1213);
nand U4468 (N_4468,N_468,N_2016);
nand U4469 (N_4469,N_1176,N_1006);
and U4470 (N_4470,N_368,N_2407);
or U4471 (N_4471,N_269,N_2209);
and U4472 (N_4472,N_1856,N_363);
xor U4473 (N_4473,N_2161,N_516);
and U4474 (N_4474,N_770,N_2453);
xnor U4475 (N_4475,N_338,N_959);
and U4476 (N_4476,N_2186,N_2097);
and U4477 (N_4477,N_2453,N_1649);
or U4478 (N_4478,N_700,N_1913);
and U4479 (N_4479,N_473,N_250);
nand U4480 (N_4480,N_1715,N_540);
or U4481 (N_4481,N_2274,N_356);
and U4482 (N_4482,N_2048,N_762);
nand U4483 (N_4483,N_1298,N_555);
xor U4484 (N_4484,N_1272,N_1812);
nand U4485 (N_4485,N_1436,N_528);
nor U4486 (N_4486,N_1071,N_1082);
and U4487 (N_4487,N_1764,N_162);
xor U4488 (N_4488,N_2269,N_2150);
or U4489 (N_4489,N_609,N_363);
nand U4490 (N_4490,N_2048,N_659);
or U4491 (N_4491,N_1038,N_300);
nand U4492 (N_4492,N_1353,N_2072);
or U4493 (N_4493,N_2496,N_825);
or U4494 (N_4494,N_871,N_459);
and U4495 (N_4495,N_1932,N_2381);
and U4496 (N_4496,N_701,N_1473);
nand U4497 (N_4497,N_1876,N_1593);
and U4498 (N_4498,N_660,N_1947);
or U4499 (N_4499,N_1462,N_300);
nor U4500 (N_4500,N_310,N_2175);
nor U4501 (N_4501,N_652,N_1008);
xnor U4502 (N_4502,N_2100,N_254);
nand U4503 (N_4503,N_642,N_1448);
nand U4504 (N_4504,N_2332,N_231);
nand U4505 (N_4505,N_700,N_1680);
nand U4506 (N_4506,N_2065,N_2083);
or U4507 (N_4507,N_1976,N_1429);
nor U4508 (N_4508,N_1111,N_1773);
nand U4509 (N_4509,N_1669,N_2134);
nand U4510 (N_4510,N_2029,N_782);
and U4511 (N_4511,N_625,N_1371);
xnor U4512 (N_4512,N_1166,N_2103);
nand U4513 (N_4513,N_1941,N_118);
xnor U4514 (N_4514,N_1197,N_279);
nor U4515 (N_4515,N_570,N_1531);
or U4516 (N_4516,N_57,N_1195);
nand U4517 (N_4517,N_1391,N_534);
xnor U4518 (N_4518,N_1516,N_1786);
xnor U4519 (N_4519,N_594,N_810);
or U4520 (N_4520,N_993,N_2071);
or U4521 (N_4521,N_743,N_1532);
nor U4522 (N_4522,N_1865,N_2219);
and U4523 (N_4523,N_838,N_110);
and U4524 (N_4524,N_1692,N_2326);
or U4525 (N_4525,N_764,N_294);
xnor U4526 (N_4526,N_731,N_1612);
and U4527 (N_4527,N_869,N_1856);
or U4528 (N_4528,N_180,N_2314);
or U4529 (N_4529,N_295,N_2460);
nor U4530 (N_4530,N_1487,N_1686);
or U4531 (N_4531,N_961,N_1775);
and U4532 (N_4532,N_293,N_601);
xor U4533 (N_4533,N_930,N_1603);
xnor U4534 (N_4534,N_1234,N_1808);
xnor U4535 (N_4535,N_1338,N_1816);
and U4536 (N_4536,N_1326,N_617);
or U4537 (N_4537,N_295,N_774);
and U4538 (N_4538,N_653,N_1335);
nand U4539 (N_4539,N_1509,N_2319);
or U4540 (N_4540,N_2009,N_867);
or U4541 (N_4541,N_1842,N_188);
xnor U4542 (N_4542,N_1637,N_1952);
nand U4543 (N_4543,N_935,N_2456);
and U4544 (N_4544,N_2217,N_16);
or U4545 (N_4545,N_486,N_2369);
nand U4546 (N_4546,N_959,N_2095);
and U4547 (N_4547,N_196,N_333);
or U4548 (N_4548,N_765,N_2435);
nor U4549 (N_4549,N_1607,N_1699);
nor U4550 (N_4550,N_230,N_416);
xor U4551 (N_4551,N_2160,N_754);
xnor U4552 (N_4552,N_1606,N_844);
xor U4553 (N_4553,N_884,N_1019);
xnor U4554 (N_4554,N_1169,N_2280);
xor U4555 (N_4555,N_243,N_744);
or U4556 (N_4556,N_1553,N_1345);
xor U4557 (N_4557,N_1855,N_1054);
nand U4558 (N_4558,N_1953,N_1082);
xor U4559 (N_4559,N_1784,N_1443);
xnor U4560 (N_4560,N_660,N_980);
xnor U4561 (N_4561,N_1514,N_1707);
nor U4562 (N_4562,N_278,N_1886);
nor U4563 (N_4563,N_1047,N_201);
and U4564 (N_4564,N_1632,N_2046);
or U4565 (N_4565,N_2302,N_821);
nand U4566 (N_4566,N_81,N_722);
nor U4567 (N_4567,N_2483,N_513);
and U4568 (N_4568,N_1306,N_138);
or U4569 (N_4569,N_2304,N_320);
and U4570 (N_4570,N_201,N_939);
nand U4571 (N_4571,N_1543,N_1153);
or U4572 (N_4572,N_1422,N_1421);
xor U4573 (N_4573,N_1500,N_1462);
and U4574 (N_4574,N_1044,N_1284);
and U4575 (N_4575,N_1984,N_384);
and U4576 (N_4576,N_313,N_1139);
nor U4577 (N_4577,N_1534,N_58);
xor U4578 (N_4578,N_38,N_1076);
nand U4579 (N_4579,N_766,N_507);
nand U4580 (N_4580,N_1739,N_1536);
nor U4581 (N_4581,N_2072,N_2348);
xnor U4582 (N_4582,N_1754,N_2313);
nand U4583 (N_4583,N_1252,N_1107);
nor U4584 (N_4584,N_1817,N_1292);
and U4585 (N_4585,N_2196,N_1277);
or U4586 (N_4586,N_1012,N_853);
nor U4587 (N_4587,N_2298,N_702);
xnor U4588 (N_4588,N_1669,N_2378);
xnor U4589 (N_4589,N_2254,N_673);
xor U4590 (N_4590,N_6,N_2199);
and U4591 (N_4591,N_1819,N_1021);
xnor U4592 (N_4592,N_1470,N_1621);
nand U4593 (N_4593,N_168,N_843);
nand U4594 (N_4594,N_1023,N_1041);
xnor U4595 (N_4595,N_864,N_259);
nor U4596 (N_4596,N_717,N_1840);
nand U4597 (N_4597,N_371,N_2066);
and U4598 (N_4598,N_1696,N_1337);
nor U4599 (N_4599,N_187,N_1916);
or U4600 (N_4600,N_251,N_148);
xor U4601 (N_4601,N_2192,N_1295);
nor U4602 (N_4602,N_1140,N_1898);
nor U4603 (N_4603,N_187,N_1611);
and U4604 (N_4604,N_2444,N_1570);
xnor U4605 (N_4605,N_2372,N_114);
and U4606 (N_4606,N_575,N_1836);
xnor U4607 (N_4607,N_1993,N_2460);
nor U4608 (N_4608,N_1066,N_1710);
and U4609 (N_4609,N_1740,N_111);
nand U4610 (N_4610,N_50,N_1174);
or U4611 (N_4611,N_1878,N_2237);
and U4612 (N_4612,N_1690,N_34);
or U4613 (N_4613,N_980,N_970);
xnor U4614 (N_4614,N_192,N_1773);
nor U4615 (N_4615,N_1582,N_1572);
nor U4616 (N_4616,N_452,N_2277);
xor U4617 (N_4617,N_1765,N_2314);
or U4618 (N_4618,N_2114,N_977);
or U4619 (N_4619,N_902,N_1227);
nor U4620 (N_4620,N_2231,N_2410);
xnor U4621 (N_4621,N_2253,N_1758);
nand U4622 (N_4622,N_159,N_1665);
nand U4623 (N_4623,N_423,N_1677);
or U4624 (N_4624,N_673,N_1161);
nor U4625 (N_4625,N_2179,N_2399);
xnor U4626 (N_4626,N_1320,N_300);
or U4627 (N_4627,N_763,N_897);
xnor U4628 (N_4628,N_1424,N_2290);
and U4629 (N_4629,N_985,N_2490);
nand U4630 (N_4630,N_698,N_1389);
and U4631 (N_4631,N_2317,N_1433);
nor U4632 (N_4632,N_676,N_22);
nand U4633 (N_4633,N_863,N_345);
and U4634 (N_4634,N_2341,N_404);
nor U4635 (N_4635,N_1834,N_512);
and U4636 (N_4636,N_233,N_691);
nand U4637 (N_4637,N_1678,N_1772);
nand U4638 (N_4638,N_1804,N_653);
nor U4639 (N_4639,N_936,N_1475);
nor U4640 (N_4640,N_2352,N_1396);
nor U4641 (N_4641,N_1800,N_241);
nand U4642 (N_4642,N_311,N_1588);
or U4643 (N_4643,N_1354,N_2315);
or U4644 (N_4644,N_1682,N_1146);
nand U4645 (N_4645,N_2084,N_1830);
nor U4646 (N_4646,N_652,N_1622);
and U4647 (N_4647,N_1222,N_2);
or U4648 (N_4648,N_2464,N_2477);
and U4649 (N_4649,N_1615,N_1553);
nor U4650 (N_4650,N_1134,N_41);
or U4651 (N_4651,N_1060,N_71);
nor U4652 (N_4652,N_34,N_178);
nand U4653 (N_4653,N_1495,N_1714);
or U4654 (N_4654,N_2205,N_201);
nand U4655 (N_4655,N_656,N_1155);
or U4656 (N_4656,N_1309,N_1198);
nand U4657 (N_4657,N_1607,N_2493);
and U4658 (N_4658,N_1091,N_1178);
or U4659 (N_4659,N_2428,N_1120);
nand U4660 (N_4660,N_442,N_115);
nand U4661 (N_4661,N_2324,N_775);
xnor U4662 (N_4662,N_1302,N_201);
and U4663 (N_4663,N_1695,N_904);
xnor U4664 (N_4664,N_180,N_594);
nand U4665 (N_4665,N_1383,N_1734);
or U4666 (N_4666,N_755,N_1081);
nand U4667 (N_4667,N_1823,N_2460);
or U4668 (N_4668,N_1290,N_1357);
xor U4669 (N_4669,N_1060,N_828);
or U4670 (N_4670,N_1918,N_911);
xnor U4671 (N_4671,N_1883,N_418);
xnor U4672 (N_4672,N_1794,N_837);
nor U4673 (N_4673,N_83,N_1545);
nand U4674 (N_4674,N_582,N_794);
nor U4675 (N_4675,N_1849,N_1540);
and U4676 (N_4676,N_589,N_957);
nor U4677 (N_4677,N_2178,N_805);
and U4678 (N_4678,N_1066,N_2150);
nor U4679 (N_4679,N_834,N_1283);
nand U4680 (N_4680,N_1341,N_1696);
and U4681 (N_4681,N_1877,N_403);
nor U4682 (N_4682,N_845,N_2216);
xnor U4683 (N_4683,N_734,N_1570);
xnor U4684 (N_4684,N_1213,N_963);
xor U4685 (N_4685,N_653,N_1409);
or U4686 (N_4686,N_2278,N_77);
and U4687 (N_4687,N_1674,N_195);
nor U4688 (N_4688,N_2250,N_86);
nor U4689 (N_4689,N_1114,N_1380);
or U4690 (N_4690,N_1993,N_1799);
or U4691 (N_4691,N_1230,N_2452);
nor U4692 (N_4692,N_2437,N_1902);
xor U4693 (N_4693,N_1452,N_1351);
xnor U4694 (N_4694,N_1999,N_1);
xor U4695 (N_4695,N_1883,N_963);
or U4696 (N_4696,N_1514,N_2100);
xor U4697 (N_4697,N_312,N_1081);
nor U4698 (N_4698,N_190,N_1259);
or U4699 (N_4699,N_702,N_1560);
xnor U4700 (N_4700,N_1598,N_595);
nor U4701 (N_4701,N_2222,N_2008);
xnor U4702 (N_4702,N_1808,N_1481);
or U4703 (N_4703,N_2071,N_1713);
nor U4704 (N_4704,N_2305,N_1565);
xor U4705 (N_4705,N_710,N_1988);
nand U4706 (N_4706,N_1094,N_2154);
or U4707 (N_4707,N_1364,N_234);
nor U4708 (N_4708,N_638,N_1433);
nand U4709 (N_4709,N_2082,N_1025);
or U4710 (N_4710,N_2101,N_712);
and U4711 (N_4711,N_1060,N_1459);
and U4712 (N_4712,N_12,N_1407);
or U4713 (N_4713,N_72,N_827);
xnor U4714 (N_4714,N_398,N_453);
xor U4715 (N_4715,N_1902,N_32);
and U4716 (N_4716,N_105,N_1827);
nor U4717 (N_4717,N_886,N_242);
or U4718 (N_4718,N_2021,N_2254);
and U4719 (N_4719,N_803,N_133);
nand U4720 (N_4720,N_1077,N_329);
or U4721 (N_4721,N_248,N_114);
xor U4722 (N_4722,N_787,N_2343);
nor U4723 (N_4723,N_1112,N_161);
nand U4724 (N_4724,N_2092,N_1565);
nor U4725 (N_4725,N_1765,N_2318);
nand U4726 (N_4726,N_1964,N_2134);
nand U4727 (N_4727,N_57,N_2495);
nor U4728 (N_4728,N_2248,N_1550);
xor U4729 (N_4729,N_1723,N_1476);
and U4730 (N_4730,N_2475,N_894);
xor U4731 (N_4731,N_686,N_935);
and U4732 (N_4732,N_1275,N_1674);
nand U4733 (N_4733,N_2108,N_1166);
nor U4734 (N_4734,N_167,N_2195);
xnor U4735 (N_4735,N_358,N_1301);
nand U4736 (N_4736,N_1702,N_759);
xnor U4737 (N_4737,N_1295,N_1635);
and U4738 (N_4738,N_1708,N_786);
or U4739 (N_4739,N_1180,N_95);
xnor U4740 (N_4740,N_583,N_756);
or U4741 (N_4741,N_1226,N_758);
xor U4742 (N_4742,N_464,N_1384);
nor U4743 (N_4743,N_621,N_1350);
or U4744 (N_4744,N_1546,N_1139);
nand U4745 (N_4745,N_193,N_1827);
xnor U4746 (N_4746,N_2229,N_2032);
nand U4747 (N_4747,N_1743,N_410);
and U4748 (N_4748,N_2100,N_737);
or U4749 (N_4749,N_201,N_1607);
and U4750 (N_4750,N_2492,N_2351);
xnor U4751 (N_4751,N_1870,N_2170);
or U4752 (N_4752,N_911,N_1345);
nand U4753 (N_4753,N_695,N_537);
and U4754 (N_4754,N_2245,N_542);
nor U4755 (N_4755,N_1981,N_2194);
nand U4756 (N_4756,N_515,N_133);
nand U4757 (N_4757,N_179,N_610);
nand U4758 (N_4758,N_633,N_463);
nand U4759 (N_4759,N_920,N_2104);
nand U4760 (N_4760,N_718,N_29);
and U4761 (N_4761,N_500,N_1912);
nand U4762 (N_4762,N_2287,N_407);
nand U4763 (N_4763,N_289,N_433);
or U4764 (N_4764,N_870,N_2346);
xnor U4765 (N_4765,N_2074,N_958);
nand U4766 (N_4766,N_2130,N_1617);
nor U4767 (N_4767,N_2173,N_1845);
xnor U4768 (N_4768,N_754,N_808);
and U4769 (N_4769,N_16,N_630);
nor U4770 (N_4770,N_2057,N_2175);
nand U4771 (N_4771,N_1240,N_2083);
or U4772 (N_4772,N_461,N_2351);
or U4773 (N_4773,N_1996,N_381);
nand U4774 (N_4774,N_452,N_646);
xor U4775 (N_4775,N_1587,N_867);
and U4776 (N_4776,N_897,N_2331);
xnor U4777 (N_4777,N_2276,N_1560);
xor U4778 (N_4778,N_824,N_199);
or U4779 (N_4779,N_1736,N_2117);
or U4780 (N_4780,N_1459,N_134);
and U4781 (N_4781,N_38,N_1696);
or U4782 (N_4782,N_1493,N_730);
xor U4783 (N_4783,N_774,N_397);
or U4784 (N_4784,N_668,N_393);
nor U4785 (N_4785,N_832,N_2023);
or U4786 (N_4786,N_36,N_723);
nand U4787 (N_4787,N_1255,N_1284);
and U4788 (N_4788,N_571,N_532);
or U4789 (N_4789,N_1970,N_799);
nor U4790 (N_4790,N_233,N_2407);
nor U4791 (N_4791,N_1797,N_1406);
or U4792 (N_4792,N_1902,N_1375);
nand U4793 (N_4793,N_55,N_2090);
nand U4794 (N_4794,N_440,N_99);
nor U4795 (N_4795,N_1824,N_2125);
xor U4796 (N_4796,N_325,N_545);
and U4797 (N_4797,N_1372,N_988);
nand U4798 (N_4798,N_1457,N_1619);
nand U4799 (N_4799,N_430,N_2295);
nor U4800 (N_4800,N_1316,N_952);
xor U4801 (N_4801,N_2062,N_2086);
and U4802 (N_4802,N_1185,N_2204);
nand U4803 (N_4803,N_1018,N_844);
nand U4804 (N_4804,N_1183,N_1026);
and U4805 (N_4805,N_1857,N_34);
xnor U4806 (N_4806,N_1785,N_254);
or U4807 (N_4807,N_517,N_875);
and U4808 (N_4808,N_2290,N_970);
nor U4809 (N_4809,N_1756,N_1307);
xnor U4810 (N_4810,N_1791,N_2086);
nand U4811 (N_4811,N_1484,N_2456);
or U4812 (N_4812,N_446,N_1494);
nor U4813 (N_4813,N_1966,N_1068);
nand U4814 (N_4814,N_1439,N_551);
xnor U4815 (N_4815,N_2486,N_727);
xnor U4816 (N_4816,N_1766,N_48);
nor U4817 (N_4817,N_1331,N_2210);
and U4818 (N_4818,N_1838,N_2109);
xnor U4819 (N_4819,N_1911,N_2267);
xor U4820 (N_4820,N_1778,N_2260);
xor U4821 (N_4821,N_370,N_1053);
xor U4822 (N_4822,N_1817,N_1041);
xnor U4823 (N_4823,N_208,N_1512);
or U4824 (N_4824,N_1880,N_2230);
or U4825 (N_4825,N_1640,N_212);
or U4826 (N_4826,N_979,N_30);
and U4827 (N_4827,N_1118,N_81);
nand U4828 (N_4828,N_1110,N_1562);
nor U4829 (N_4829,N_864,N_1830);
nor U4830 (N_4830,N_827,N_1656);
or U4831 (N_4831,N_1793,N_2391);
nor U4832 (N_4832,N_448,N_1147);
and U4833 (N_4833,N_1326,N_1247);
or U4834 (N_4834,N_1223,N_1644);
xor U4835 (N_4835,N_1988,N_735);
nand U4836 (N_4836,N_1043,N_1341);
nand U4837 (N_4837,N_775,N_2422);
xor U4838 (N_4838,N_497,N_514);
xnor U4839 (N_4839,N_1297,N_1529);
nor U4840 (N_4840,N_704,N_2113);
nor U4841 (N_4841,N_2473,N_1132);
nor U4842 (N_4842,N_2343,N_2103);
xor U4843 (N_4843,N_2015,N_1481);
nand U4844 (N_4844,N_1769,N_824);
or U4845 (N_4845,N_1676,N_1266);
or U4846 (N_4846,N_780,N_1406);
nand U4847 (N_4847,N_2086,N_1547);
or U4848 (N_4848,N_2292,N_972);
or U4849 (N_4849,N_399,N_151);
and U4850 (N_4850,N_772,N_528);
nand U4851 (N_4851,N_1694,N_374);
or U4852 (N_4852,N_472,N_367);
or U4853 (N_4853,N_961,N_552);
or U4854 (N_4854,N_150,N_1102);
nor U4855 (N_4855,N_1141,N_1854);
or U4856 (N_4856,N_138,N_807);
xor U4857 (N_4857,N_40,N_1225);
or U4858 (N_4858,N_344,N_222);
or U4859 (N_4859,N_2252,N_1914);
or U4860 (N_4860,N_564,N_2344);
or U4861 (N_4861,N_530,N_77);
or U4862 (N_4862,N_2146,N_2121);
xnor U4863 (N_4863,N_2319,N_1651);
and U4864 (N_4864,N_1145,N_863);
nor U4865 (N_4865,N_568,N_966);
nand U4866 (N_4866,N_758,N_1925);
nor U4867 (N_4867,N_274,N_347);
and U4868 (N_4868,N_1890,N_459);
xor U4869 (N_4869,N_1440,N_1247);
nand U4870 (N_4870,N_1255,N_1610);
xnor U4871 (N_4871,N_1571,N_751);
nand U4872 (N_4872,N_599,N_625);
xor U4873 (N_4873,N_457,N_1572);
nor U4874 (N_4874,N_1733,N_1019);
nor U4875 (N_4875,N_2461,N_2303);
nand U4876 (N_4876,N_1615,N_1331);
nor U4877 (N_4877,N_508,N_2303);
or U4878 (N_4878,N_2331,N_441);
nand U4879 (N_4879,N_456,N_1047);
or U4880 (N_4880,N_1922,N_1016);
or U4881 (N_4881,N_1381,N_2081);
or U4882 (N_4882,N_1173,N_1653);
or U4883 (N_4883,N_1460,N_304);
xor U4884 (N_4884,N_1350,N_2420);
and U4885 (N_4885,N_973,N_1029);
xor U4886 (N_4886,N_610,N_1800);
xor U4887 (N_4887,N_1518,N_1670);
or U4888 (N_4888,N_1548,N_117);
nand U4889 (N_4889,N_1467,N_2101);
and U4890 (N_4890,N_433,N_1628);
nor U4891 (N_4891,N_1240,N_0);
nor U4892 (N_4892,N_332,N_1894);
nor U4893 (N_4893,N_2013,N_2191);
or U4894 (N_4894,N_1090,N_2377);
xor U4895 (N_4895,N_628,N_962);
nand U4896 (N_4896,N_98,N_295);
and U4897 (N_4897,N_470,N_662);
xnor U4898 (N_4898,N_1100,N_62);
and U4899 (N_4899,N_1255,N_1948);
or U4900 (N_4900,N_2230,N_328);
nor U4901 (N_4901,N_45,N_2461);
or U4902 (N_4902,N_2099,N_125);
xor U4903 (N_4903,N_1531,N_193);
and U4904 (N_4904,N_1723,N_2045);
xnor U4905 (N_4905,N_912,N_200);
or U4906 (N_4906,N_2474,N_2309);
or U4907 (N_4907,N_1811,N_2155);
nor U4908 (N_4908,N_1666,N_1896);
and U4909 (N_4909,N_628,N_92);
nand U4910 (N_4910,N_183,N_1516);
nor U4911 (N_4911,N_2150,N_979);
and U4912 (N_4912,N_713,N_622);
nor U4913 (N_4913,N_2375,N_1621);
xor U4914 (N_4914,N_366,N_562);
and U4915 (N_4915,N_2305,N_1617);
or U4916 (N_4916,N_813,N_1569);
and U4917 (N_4917,N_1404,N_469);
and U4918 (N_4918,N_100,N_174);
nor U4919 (N_4919,N_1095,N_512);
xor U4920 (N_4920,N_166,N_2471);
and U4921 (N_4921,N_784,N_345);
nor U4922 (N_4922,N_1680,N_521);
xor U4923 (N_4923,N_122,N_2151);
xnor U4924 (N_4924,N_1617,N_723);
xnor U4925 (N_4925,N_1098,N_1900);
xnor U4926 (N_4926,N_1697,N_1608);
xor U4927 (N_4927,N_2451,N_2131);
nand U4928 (N_4928,N_1383,N_214);
and U4929 (N_4929,N_479,N_2232);
or U4930 (N_4930,N_544,N_1241);
and U4931 (N_4931,N_840,N_2060);
nand U4932 (N_4932,N_419,N_378);
nor U4933 (N_4933,N_1329,N_2434);
and U4934 (N_4934,N_982,N_1392);
or U4935 (N_4935,N_1578,N_1262);
nand U4936 (N_4936,N_1168,N_1804);
or U4937 (N_4937,N_2317,N_2220);
nor U4938 (N_4938,N_1909,N_1597);
nor U4939 (N_4939,N_478,N_1406);
or U4940 (N_4940,N_865,N_996);
and U4941 (N_4941,N_649,N_306);
xor U4942 (N_4942,N_1139,N_1347);
and U4943 (N_4943,N_1006,N_416);
nor U4944 (N_4944,N_1520,N_813);
nor U4945 (N_4945,N_516,N_348);
nor U4946 (N_4946,N_59,N_2401);
xor U4947 (N_4947,N_907,N_2089);
xor U4948 (N_4948,N_295,N_811);
or U4949 (N_4949,N_207,N_1300);
xor U4950 (N_4950,N_1717,N_434);
nand U4951 (N_4951,N_1901,N_312);
or U4952 (N_4952,N_1731,N_1445);
xor U4953 (N_4953,N_1612,N_936);
or U4954 (N_4954,N_2144,N_513);
and U4955 (N_4955,N_2026,N_1369);
nor U4956 (N_4956,N_1872,N_1659);
xnor U4957 (N_4957,N_1370,N_1265);
or U4958 (N_4958,N_1787,N_323);
or U4959 (N_4959,N_1780,N_2107);
nor U4960 (N_4960,N_985,N_1973);
or U4961 (N_4961,N_1566,N_909);
and U4962 (N_4962,N_1227,N_465);
nand U4963 (N_4963,N_694,N_1072);
nor U4964 (N_4964,N_1971,N_1267);
nor U4965 (N_4965,N_1639,N_1261);
nand U4966 (N_4966,N_2133,N_2006);
nand U4967 (N_4967,N_1452,N_2001);
nor U4968 (N_4968,N_1409,N_833);
xnor U4969 (N_4969,N_1722,N_1699);
nand U4970 (N_4970,N_2021,N_1743);
and U4971 (N_4971,N_1958,N_98);
or U4972 (N_4972,N_2404,N_2380);
nor U4973 (N_4973,N_1627,N_303);
xnor U4974 (N_4974,N_1714,N_849);
xnor U4975 (N_4975,N_1388,N_1679);
or U4976 (N_4976,N_1234,N_1838);
and U4977 (N_4977,N_1563,N_1517);
xnor U4978 (N_4978,N_621,N_2159);
nor U4979 (N_4979,N_276,N_786);
or U4980 (N_4980,N_1158,N_1902);
and U4981 (N_4981,N_992,N_900);
nand U4982 (N_4982,N_2385,N_1505);
nand U4983 (N_4983,N_562,N_2244);
or U4984 (N_4984,N_1611,N_1186);
nand U4985 (N_4985,N_900,N_762);
and U4986 (N_4986,N_1491,N_1975);
nor U4987 (N_4987,N_1371,N_1005);
nor U4988 (N_4988,N_1105,N_1044);
nand U4989 (N_4989,N_2120,N_1542);
nor U4990 (N_4990,N_389,N_13);
nor U4991 (N_4991,N_842,N_331);
nor U4992 (N_4992,N_353,N_946);
xor U4993 (N_4993,N_703,N_1937);
xor U4994 (N_4994,N_2153,N_2329);
xor U4995 (N_4995,N_2151,N_2382);
nor U4996 (N_4996,N_2497,N_2017);
xor U4997 (N_4997,N_86,N_495);
nand U4998 (N_4998,N_1705,N_1791);
or U4999 (N_4999,N_1468,N_1832);
and U5000 (N_5000,N_3923,N_4360);
and U5001 (N_5001,N_2628,N_4634);
nand U5002 (N_5002,N_3615,N_4259);
nor U5003 (N_5003,N_4680,N_3131);
nand U5004 (N_5004,N_3255,N_3281);
or U5005 (N_5005,N_3791,N_4286);
nand U5006 (N_5006,N_3513,N_3142);
or U5007 (N_5007,N_2866,N_2944);
or U5008 (N_5008,N_4105,N_3429);
and U5009 (N_5009,N_3945,N_4992);
nor U5010 (N_5010,N_2622,N_4130);
and U5011 (N_5011,N_4629,N_3064);
nor U5012 (N_5012,N_4198,N_4667);
xnor U5013 (N_5013,N_4582,N_4212);
nor U5014 (N_5014,N_3901,N_3022);
nor U5015 (N_5015,N_2845,N_3413);
or U5016 (N_5016,N_2935,N_3363);
nor U5017 (N_5017,N_3608,N_3486);
nor U5018 (N_5018,N_4632,N_4804);
and U5019 (N_5019,N_3378,N_4409);
nand U5020 (N_5020,N_3360,N_4700);
nand U5021 (N_5021,N_3437,N_2901);
nand U5022 (N_5022,N_3081,N_4319);
xnor U5023 (N_5023,N_4094,N_4496);
nor U5024 (N_5024,N_4605,N_4183);
xnor U5025 (N_5025,N_3013,N_4576);
nand U5026 (N_5026,N_3840,N_4065);
xor U5027 (N_5027,N_3578,N_4111);
nand U5028 (N_5028,N_2542,N_4792);
nand U5029 (N_5029,N_2800,N_4805);
nor U5030 (N_5030,N_4527,N_2985);
and U5031 (N_5031,N_2728,N_3158);
nor U5032 (N_5032,N_4144,N_4813);
nor U5033 (N_5033,N_4536,N_4169);
or U5034 (N_5034,N_3994,N_4981);
xor U5035 (N_5035,N_3720,N_4372);
nor U5036 (N_5036,N_2959,N_4455);
or U5037 (N_5037,N_2912,N_4693);
xnor U5038 (N_5038,N_3756,N_4980);
xnor U5039 (N_5039,N_2909,N_3166);
nor U5040 (N_5040,N_3477,N_4038);
nor U5041 (N_5041,N_2641,N_3082);
nand U5042 (N_5042,N_4067,N_3427);
or U5043 (N_5043,N_3277,N_4301);
or U5044 (N_5044,N_2822,N_3966);
and U5045 (N_5045,N_2829,N_4196);
xor U5046 (N_5046,N_3853,N_2864);
and U5047 (N_5047,N_3842,N_4084);
nor U5048 (N_5048,N_3792,N_4808);
nand U5049 (N_5049,N_4763,N_4614);
or U5050 (N_5050,N_4459,N_3249);
xnor U5051 (N_5051,N_4753,N_4015);
nor U5052 (N_5052,N_2741,N_3356);
or U5053 (N_5053,N_3491,N_4335);
or U5054 (N_5054,N_4546,N_2520);
or U5055 (N_5055,N_3447,N_3884);
and U5056 (N_5056,N_3212,N_4236);
xnor U5057 (N_5057,N_4171,N_4575);
and U5058 (N_5058,N_3334,N_4002);
or U5059 (N_5059,N_4976,N_3565);
nor U5060 (N_5060,N_3444,N_4456);
xor U5061 (N_5061,N_4504,N_2994);
nand U5062 (N_5062,N_4477,N_3926);
nor U5063 (N_5063,N_3112,N_4881);
nand U5064 (N_5064,N_3569,N_3471);
nor U5065 (N_5065,N_2662,N_4129);
and U5066 (N_5066,N_3071,N_4514);
or U5067 (N_5067,N_2993,N_3490);
xor U5068 (N_5068,N_4978,N_2750);
and U5069 (N_5069,N_3837,N_2565);
nor U5070 (N_5070,N_3958,N_2625);
nand U5071 (N_5071,N_4030,N_2519);
nor U5072 (N_5072,N_3711,N_4426);
and U5073 (N_5073,N_2821,N_4369);
xor U5074 (N_5074,N_4505,N_3001);
or U5075 (N_5075,N_4652,N_3521);
or U5076 (N_5076,N_3401,N_3902);
nand U5077 (N_5077,N_3929,N_3805);
nand U5078 (N_5078,N_4793,N_2646);
xnor U5079 (N_5079,N_3138,N_4288);
and U5080 (N_5080,N_4403,N_3391);
xor U5081 (N_5081,N_4469,N_2588);
nor U5082 (N_5082,N_2907,N_4012);
nand U5083 (N_5083,N_2804,N_3950);
and U5084 (N_5084,N_3306,N_3379);
or U5085 (N_5085,N_3388,N_2721);
and U5086 (N_5086,N_4098,N_2505);
xnor U5087 (N_5087,N_3612,N_3178);
or U5088 (N_5088,N_3193,N_3610);
nand U5089 (N_5089,N_2934,N_2884);
nand U5090 (N_5090,N_4449,N_3742);
nor U5091 (N_5091,N_3536,N_3523);
nand U5092 (N_5092,N_4585,N_4026);
or U5093 (N_5093,N_2963,N_4363);
nor U5094 (N_5094,N_4275,N_3492);
nand U5095 (N_5095,N_2808,N_3289);
or U5096 (N_5096,N_4701,N_3298);
nand U5097 (N_5097,N_3012,N_3554);
nand U5098 (N_5098,N_2958,N_3269);
nor U5099 (N_5099,N_2510,N_4247);
or U5100 (N_5100,N_4280,N_4079);
or U5101 (N_5101,N_4811,N_3392);
nand U5102 (N_5102,N_3267,N_4923);
or U5103 (N_5103,N_3888,N_3616);
and U5104 (N_5104,N_4194,N_3540);
xor U5105 (N_5105,N_3246,N_3182);
and U5106 (N_5106,N_4243,N_3149);
nand U5107 (N_5107,N_2862,N_3520);
and U5108 (N_5108,N_3896,N_4383);
xor U5109 (N_5109,N_3641,N_3383);
xnor U5110 (N_5110,N_3233,N_4187);
xor U5111 (N_5111,N_2514,N_3253);
and U5112 (N_5112,N_3900,N_3496);
nor U5113 (N_5113,N_3075,N_4491);
or U5114 (N_5114,N_3003,N_4151);
nor U5115 (N_5115,N_3783,N_3362);
nand U5116 (N_5116,N_2701,N_3596);
and U5117 (N_5117,N_3665,N_2924);
nor U5118 (N_5118,N_4666,N_4779);
or U5119 (N_5119,N_3949,N_4952);
or U5120 (N_5120,N_2870,N_4683);
nand U5121 (N_5121,N_3141,N_2850);
nand U5122 (N_5122,N_2962,N_3291);
nand U5123 (N_5123,N_3484,N_3262);
nor U5124 (N_5124,N_2785,N_4953);
and U5125 (N_5125,N_4088,N_3497);
xor U5126 (N_5126,N_4201,N_3635);
nor U5127 (N_5127,N_4966,N_3935);
xor U5128 (N_5128,N_4972,N_3323);
xor U5129 (N_5129,N_4176,N_2802);
xnor U5130 (N_5130,N_2516,N_4797);
and U5131 (N_5131,N_2773,N_4959);
nor U5132 (N_5132,N_4838,N_3442);
nor U5133 (N_5133,N_4934,N_2757);
nor U5134 (N_5134,N_2776,N_2562);
nand U5135 (N_5135,N_3609,N_3271);
or U5136 (N_5136,N_4764,N_4049);
xor U5137 (N_5137,N_4004,N_3780);
or U5138 (N_5138,N_3803,N_2723);
or U5139 (N_5139,N_4555,N_4896);
nor U5140 (N_5140,N_4298,N_3577);
xor U5141 (N_5141,N_3365,N_4836);
xor U5142 (N_5142,N_4907,N_4832);
nand U5143 (N_5143,N_4947,N_2610);
or U5144 (N_5144,N_2971,N_4495);
and U5145 (N_5145,N_3217,N_3708);
and U5146 (N_5146,N_3348,N_3710);
nand U5147 (N_5147,N_4780,N_4097);
xor U5148 (N_5148,N_4076,N_4149);
and U5149 (N_5149,N_4528,N_3647);
nand U5150 (N_5150,N_4862,N_4868);
or U5151 (N_5151,N_2584,N_3571);
and U5152 (N_5152,N_3525,N_4725);
nor U5153 (N_5153,N_4736,N_4810);
nor U5154 (N_5154,N_4005,N_3252);
nand U5155 (N_5155,N_4771,N_4530);
or U5156 (N_5156,N_2657,N_4150);
nand U5157 (N_5157,N_4599,N_4179);
nand U5158 (N_5158,N_3095,N_4317);
nor U5159 (N_5159,N_4277,N_3770);
nand U5160 (N_5160,N_3646,N_4690);
xnor U5161 (N_5161,N_3237,N_3913);
or U5162 (N_5162,N_4886,N_3113);
nand U5163 (N_5163,N_3371,N_4561);
and U5164 (N_5164,N_3152,N_2787);
xnor U5165 (N_5165,N_3036,N_4261);
and U5166 (N_5166,N_2508,N_3495);
xor U5167 (N_5167,N_4189,N_4675);
nand U5168 (N_5168,N_3656,N_3204);
nor U5169 (N_5169,N_3587,N_3802);
xnor U5170 (N_5170,N_4705,N_3136);
or U5171 (N_5171,N_2563,N_2927);
nand U5172 (N_5172,N_3181,N_3939);
nand U5173 (N_5173,N_4510,N_4917);
nand U5174 (N_5174,N_3468,N_3117);
nor U5175 (N_5175,N_4929,N_2941);
xnor U5176 (N_5176,N_3225,N_2856);
nor U5177 (N_5177,N_3586,N_2745);
or U5178 (N_5178,N_2846,N_4518);
nand U5179 (N_5179,N_4451,N_3592);
nand U5180 (N_5180,N_2975,N_4679);
nor U5181 (N_5181,N_3807,N_3983);
nand U5182 (N_5182,N_4995,N_4269);
or U5183 (N_5183,N_2583,N_3416);
nand U5184 (N_5184,N_2966,N_3076);
nand U5185 (N_5185,N_2697,N_2679);
nand U5186 (N_5186,N_3693,N_3874);
nor U5187 (N_5187,N_4345,N_3631);
or U5188 (N_5188,N_4148,N_2685);
nor U5189 (N_5189,N_3529,N_3368);
xnor U5190 (N_5190,N_3445,N_2801);
xor U5191 (N_5191,N_4356,N_4170);
and U5192 (N_5192,N_4658,N_3026);
and U5193 (N_5193,N_3432,N_4454);
xnor U5194 (N_5194,N_3029,N_4444);
nand U5195 (N_5195,N_2711,N_3299);
nand U5196 (N_5196,N_3015,N_4601);
or U5197 (N_5197,N_4028,N_3642);
or U5198 (N_5198,N_2521,N_3735);
or U5199 (N_5199,N_3698,N_3314);
nand U5200 (N_5200,N_3597,N_3895);
nor U5201 (N_5201,N_3589,N_2531);
xor U5202 (N_5202,N_2990,N_4070);
and U5203 (N_5203,N_3088,N_4054);
nand U5204 (N_5204,N_3806,N_2596);
nor U5205 (N_5205,N_3493,N_4651);
or U5206 (N_5206,N_4979,N_4205);
or U5207 (N_5207,N_4441,N_4722);
and U5208 (N_5208,N_4050,N_3366);
nand U5209 (N_5209,N_2806,N_4487);
nand U5210 (N_5210,N_2987,N_4726);
and U5211 (N_5211,N_3768,N_3175);
and U5212 (N_5212,N_4677,N_4931);
nor U5213 (N_5213,N_3917,N_2591);
nand U5214 (N_5214,N_4364,N_4948);
nand U5215 (N_5215,N_2938,N_3364);
and U5216 (N_5216,N_3727,N_4944);
or U5217 (N_5217,N_4964,N_4355);
and U5218 (N_5218,N_2817,N_4580);
nor U5219 (N_5219,N_3428,N_4627);
or U5220 (N_5220,N_2714,N_4579);
nor U5221 (N_5221,N_2707,N_3216);
and U5222 (N_5222,N_2736,N_2566);
or U5223 (N_5223,N_4075,N_2502);
or U5224 (N_5224,N_3165,N_3512);
nand U5225 (N_5225,N_3658,N_4106);
and U5226 (N_5226,N_4894,N_3730);
xor U5227 (N_5227,N_3111,N_3942);
nor U5228 (N_5228,N_2760,N_4022);
nor U5229 (N_5229,N_3914,N_3637);
or U5230 (N_5230,N_4562,N_4760);
or U5231 (N_5231,N_2857,N_3705);
nand U5232 (N_5232,N_3067,N_4209);
nor U5233 (N_5233,N_3679,N_4029);
nor U5234 (N_5234,N_2744,N_4545);
or U5235 (N_5235,N_4347,N_4937);
or U5236 (N_5236,N_4759,N_4628);
nand U5237 (N_5237,N_4738,N_4946);
or U5238 (N_5238,N_4548,N_3124);
nand U5239 (N_5239,N_4146,N_3527);
or U5240 (N_5240,N_3307,N_4963);
or U5241 (N_5241,N_4370,N_3580);
nand U5242 (N_5242,N_2501,N_3634);
or U5243 (N_5243,N_2546,N_4788);
xor U5244 (N_5244,N_3350,N_3263);
nand U5245 (N_5245,N_4322,N_2820);
or U5246 (N_5246,N_3753,N_4865);
and U5247 (N_5247,N_2556,N_2995);
or U5248 (N_5248,N_4252,N_2762);
or U5249 (N_5249,N_4720,N_4904);
xnor U5250 (N_5250,N_3184,N_3144);
and U5251 (N_5251,N_2636,N_2555);
nand U5252 (N_5252,N_4354,N_4107);
nor U5253 (N_5253,N_4271,N_2658);
xor U5254 (N_5254,N_4998,N_2983);
nand U5255 (N_5255,N_3930,N_4668);
nor U5256 (N_5256,N_3021,N_3723);
nor U5257 (N_5257,N_2605,N_3098);
or U5258 (N_5258,N_4604,N_3957);
nand U5259 (N_5259,N_3691,N_4711);
nor U5260 (N_5260,N_3568,N_3223);
or U5261 (N_5261,N_3984,N_4751);
and U5262 (N_5262,N_4968,N_4554);
xor U5263 (N_5263,N_3244,N_3800);
and U5264 (N_5264,N_4475,N_2602);
nor U5265 (N_5265,N_4816,N_2877);
or U5266 (N_5266,N_4202,N_3016);
and U5267 (N_5267,N_4912,N_4384);
xnor U5268 (N_5268,N_4860,N_3359);
or U5269 (N_5269,N_4197,N_4331);
xnor U5270 (N_5270,N_4279,N_3420);
nor U5271 (N_5271,N_3189,N_3582);
or U5272 (N_5272,N_2835,N_4297);
and U5273 (N_5273,N_3501,N_4213);
nand U5274 (N_5274,N_2836,N_4927);
xor U5275 (N_5275,N_3313,N_4276);
nor U5276 (N_5276,N_3759,N_2643);
nor U5277 (N_5277,N_3894,N_4134);
nand U5278 (N_5278,N_3606,N_4435);
nand U5279 (N_5279,N_3991,N_3352);
nand U5280 (N_5280,N_2621,N_2812);
or U5281 (N_5281,N_4965,N_4195);
nand U5282 (N_5282,N_4900,N_2706);
and U5283 (N_5283,N_4461,N_3228);
and U5284 (N_5284,N_3311,N_2917);
or U5285 (N_5285,N_4603,N_4359);
nand U5286 (N_5286,N_3941,N_4311);
and U5287 (N_5287,N_4436,N_3618);
or U5288 (N_5288,N_4040,N_3715);
nor U5289 (N_5289,N_4732,N_4296);
nand U5290 (N_5290,N_3393,N_4498);
nand U5291 (N_5291,N_2548,N_4997);
and U5292 (N_5292,N_3848,N_2704);
nand U5293 (N_5293,N_4513,N_4800);
or U5294 (N_5294,N_2549,N_4381);
or U5295 (N_5295,N_2718,N_3978);
xnor U5296 (N_5296,N_2891,N_2950);
nor U5297 (N_5297,N_3301,N_3947);
xnor U5298 (N_5298,N_4291,N_4342);
and U5299 (N_5299,N_3208,N_3555);
and U5300 (N_5300,N_4217,N_2922);
or U5301 (N_5301,N_4707,N_2998);
xor U5302 (N_5302,N_3153,N_4650);
or U5303 (N_5303,N_2897,N_4453);
and U5304 (N_5304,N_4165,N_4718);
or U5305 (N_5305,N_4433,N_2559);
or U5306 (N_5306,N_4737,N_4895);
and U5307 (N_5307,N_4227,N_2765);
xor U5308 (N_5308,N_3714,N_3040);
and U5309 (N_5309,N_3843,N_3514);
nor U5310 (N_5310,N_4293,N_4153);
nor U5311 (N_5311,N_3844,N_4787);
or U5312 (N_5312,N_2876,N_4299);
nand U5313 (N_5313,N_3077,N_4349);
nor U5314 (N_5314,N_4648,N_3732);
nand U5315 (N_5315,N_4919,N_4159);
and U5316 (N_5316,N_2522,N_4540);
nand U5317 (N_5317,N_4781,N_3174);
xor U5318 (N_5318,N_3406,N_4091);
nand U5319 (N_5319,N_2968,N_3517);
and U5320 (N_5320,N_2727,N_2888);
nor U5321 (N_5321,N_3018,N_3008);
nand U5322 (N_5322,N_3877,N_3054);
and U5323 (N_5323,N_3483,N_3801);
or U5324 (N_5324,N_3534,N_3159);
nor U5325 (N_5325,N_4871,N_3272);
xor U5326 (N_5326,N_4685,N_2567);
nor U5327 (N_5327,N_4366,N_2500);
or U5328 (N_5328,N_2933,N_3426);
nor U5329 (N_5329,N_2920,N_3719);
nor U5330 (N_5330,N_3147,N_2648);
or U5331 (N_5331,N_3810,N_4717);
or U5332 (N_5332,N_3275,N_3456);
nor U5333 (N_5333,N_2681,N_3200);
or U5334 (N_5334,N_2553,N_3954);
nand U5335 (N_5335,N_3910,N_3422);
nor U5336 (N_5336,N_4672,N_4192);
and U5337 (N_5337,N_2945,N_3948);
xor U5338 (N_5338,N_3296,N_4801);
nor U5339 (N_5339,N_4400,N_2809);
nand U5340 (N_5340,N_4138,N_4878);
nor U5341 (N_5341,N_2929,N_3157);
nor U5342 (N_5342,N_4289,N_4041);
or U5343 (N_5343,N_4141,N_3817);
nand U5344 (N_5344,N_2923,N_4786);
nor U5345 (N_5345,N_4689,N_4415);
xnor U5346 (N_5346,N_2504,N_4837);
nor U5347 (N_5347,N_3648,N_3762);
nand U5348 (N_5348,N_4733,N_4336);
nor U5349 (N_5349,N_4493,N_3229);
nand U5350 (N_5350,N_3583,N_3788);
xor U5351 (N_5351,N_4893,N_2590);
and U5352 (N_5352,N_2833,N_3214);
nand U5353 (N_5353,N_2587,N_4702);
nor U5354 (N_5354,N_2512,N_2843);
xor U5355 (N_5355,N_3660,N_4984);
and U5356 (N_5356,N_3607,N_4407);
and U5357 (N_5357,N_4284,N_3470);
xor U5358 (N_5358,N_3069,N_3031);
nand U5359 (N_5359,N_3668,N_3833);
or U5360 (N_5360,N_4913,N_4031);
xor U5361 (N_5361,N_3039,N_4873);
or U5362 (N_5362,N_3655,N_2530);
nor U5363 (N_5363,N_3411,N_3717);
nor U5364 (N_5364,N_3245,N_3572);
nor U5365 (N_5365,N_2709,N_3293);
or U5366 (N_5366,N_2665,N_3854);
nor U5367 (N_5367,N_2623,N_4147);
and U5368 (N_5368,N_4883,N_4140);
and U5369 (N_5369,N_2717,N_2732);
or U5370 (N_5370,N_4663,N_3969);
nor U5371 (N_5371,N_3130,N_3243);
or U5372 (N_5372,N_4468,N_3890);
nor U5373 (N_5373,N_4665,N_3057);
and U5374 (N_5374,N_3614,N_3503);
xnor U5375 (N_5375,N_3498,N_2577);
and U5376 (N_5376,N_3881,N_2581);
xor U5377 (N_5377,N_4292,N_3357);
nand U5378 (N_5378,N_4327,N_4330);
and U5379 (N_5379,N_4419,N_2989);
xnor U5380 (N_5380,N_2978,N_4656);
xnor U5381 (N_5381,N_3982,N_3099);
nor U5382 (N_5382,N_3774,N_4078);
or U5383 (N_5383,N_4000,N_4256);
and U5384 (N_5384,N_2979,N_4567);
or U5385 (N_5385,N_4290,N_2789);
or U5386 (N_5386,N_4118,N_2970);
nor U5387 (N_5387,N_4538,N_4282);
nor U5388 (N_5388,N_3358,N_3836);
or U5389 (N_5389,N_4758,N_2545);
and U5390 (N_5390,N_3654,N_4835);
nand U5391 (N_5391,N_3478,N_2654);
xnor U5392 (N_5392,N_3338,N_2614);
or U5393 (N_5393,N_3259,N_3686);
nand U5394 (N_5394,N_3302,N_4741);
nand U5395 (N_5395,N_3904,N_3516);
or U5396 (N_5396,N_3309,N_3889);
xnor U5397 (N_5397,N_4018,N_4664);
or U5398 (N_5398,N_3886,N_2572);
xnor U5399 (N_5399,N_4214,N_3198);
and U5400 (N_5400,N_4817,N_2595);
nand U5401 (N_5401,N_4180,N_3701);
nand U5402 (N_5402,N_2552,N_4861);
nand U5403 (N_5403,N_4373,N_3241);
and U5404 (N_5404,N_3731,N_4686);
xnor U5405 (N_5405,N_3505,N_4853);
nand U5406 (N_5406,N_3786,N_4714);
nand U5407 (N_5407,N_4464,N_3195);
and U5408 (N_5408,N_3125,N_2881);
and U5409 (N_5409,N_3532,N_3137);
nand U5410 (N_5410,N_3330,N_4523);
nor U5411 (N_5411,N_4077,N_4010);
nand U5412 (N_5412,N_2782,N_3955);
and U5413 (N_5413,N_3530,N_2982);
and U5414 (N_5414,N_3479,N_3871);
nand U5415 (N_5415,N_3893,N_3155);
nand U5416 (N_5416,N_4221,N_3559);
and U5417 (N_5417,N_4857,N_2842);
nor U5418 (N_5418,N_4938,N_2653);
nor U5419 (N_5419,N_4262,N_3453);
and U5420 (N_5420,N_4954,N_3489);
xor U5421 (N_5421,N_2631,N_3625);
nor U5422 (N_5422,N_3058,N_4386);
xor U5423 (N_5423,N_4594,N_4219);
or U5424 (N_5424,N_3541,N_4402);
and U5425 (N_5425,N_3102,N_4273);
and U5426 (N_5426,N_4230,N_4586);
or U5427 (N_5427,N_3795,N_3093);
xnor U5428 (N_5428,N_3928,N_4371);
nand U5429 (N_5429,N_2739,N_3740);
xnor U5430 (N_5430,N_3210,N_4610);
or U5431 (N_5431,N_2680,N_3985);
xnor U5432 (N_5432,N_2984,N_3177);
or U5433 (N_5433,N_2976,N_3100);
xor U5434 (N_5434,N_4774,N_3139);
xnor U5435 (N_5435,N_3769,N_2551);
and U5436 (N_5436,N_2981,N_4542);
xnor U5437 (N_5437,N_4945,N_4316);
or U5438 (N_5438,N_3068,N_3287);
nor U5439 (N_5439,N_2918,N_3767);
xnor U5440 (N_5440,N_3932,N_3304);
xor U5441 (N_5441,N_3603,N_3190);
nor U5442 (N_5442,N_3870,N_4785);
and U5443 (N_5443,N_4164,N_4987);
nand U5444 (N_5444,N_2585,N_3562);
and U5445 (N_5445,N_4820,N_3238);
nand U5446 (N_5446,N_2986,N_4389);
nand U5447 (N_5447,N_3997,N_3946);
or U5448 (N_5448,N_3461,N_3186);
or U5449 (N_5449,N_2637,N_4420);
nor U5450 (N_5450,N_3353,N_4458);
and U5451 (N_5451,N_4250,N_3355);
xnor U5452 (N_5452,N_4583,N_4588);
nand U5453 (N_5453,N_3838,N_2564);
nor U5454 (N_5454,N_3628,N_3337);
and U5455 (N_5455,N_3344,N_4391);
or U5456 (N_5456,N_4897,N_4511);
xnor U5457 (N_5457,N_3384,N_4818);
or U5458 (N_5458,N_3163,N_2582);
nand U5459 (N_5459,N_3687,N_3875);
and U5460 (N_5460,N_4157,N_2752);
or U5461 (N_5461,N_4595,N_4401);
and U5462 (N_5462,N_3509,N_4408);
nor U5463 (N_5463,N_3222,N_4184);
nor U5464 (N_5464,N_3123,N_3743);
nor U5465 (N_5465,N_3621,N_4237);
xnor U5466 (N_5466,N_4957,N_4925);
nor U5467 (N_5467,N_3974,N_3494);
and U5468 (N_5468,N_2908,N_4242);
nor U5469 (N_5469,N_3151,N_3316);
or U5470 (N_5470,N_2956,N_2532);
or U5471 (N_5471,N_3375,N_4199);
nor U5472 (N_5472,N_2754,N_4607);
and U5473 (N_5473,N_4709,N_4521);
nand U5474 (N_5474,N_2670,N_4678);
or U5475 (N_5475,N_3797,N_4566);
and U5476 (N_5476,N_4225,N_4003);
xnor U5477 (N_5477,N_3448,N_4254);
xor U5478 (N_5478,N_2777,N_2837);
or U5479 (N_5479,N_4844,N_4827);
nor U5480 (N_5480,N_2560,N_4855);
and U5481 (N_5481,N_3419,N_4739);
or U5482 (N_5482,N_4754,N_3972);
or U5483 (N_5483,N_4856,N_3257);
nor U5484 (N_5484,N_4684,N_4053);
nand U5485 (N_5485,N_3911,N_3037);
nor U5486 (N_5486,N_4670,N_3772);
or U5487 (N_5487,N_3303,N_3862);
nor U5488 (N_5488,N_4790,N_4543);
and U5489 (N_5489,N_4344,N_4274);
nand U5490 (N_5490,N_3466,N_3763);
xor U5491 (N_5491,N_3998,N_4220);
nand U5492 (N_5492,N_4885,N_3120);
xor U5493 (N_5493,N_4338,N_2533);
nand U5494 (N_5494,N_2650,N_4188);
or U5495 (N_5495,N_2571,N_4266);
nor U5496 (N_5496,N_3524,N_4626);
nand U5497 (N_5497,N_2951,N_3765);
xor U5498 (N_5498,N_2851,N_2738);
nand U5499 (N_5499,N_3755,N_3827);
nand U5500 (N_5500,N_4822,N_3162);
and U5501 (N_5501,N_2834,N_3282);
nand U5502 (N_5502,N_2682,N_2573);
xor U5503 (N_5503,N_3822,N_3140);
nor U5504 (N_5504,N_3482,N_2919);
nor U5505 (N_5505,N_3059,N_4395);
and U5506 (N_5506,N_2601,N_4257);
xor U5507 (N_5507,N_2865,N_4253);
or U5508 (N_5508,N_3038,N_3256);
or U5509 (N_5509,N_3652,N_4922);
nand U5510 (N_5510,N_3733,N_4425);
or U5511 (N_5511,N_4695,N_3602);
and U5512 (N_5512,N_3266,N_4564);
or U5513 (N_5513,N_4177,N_3661);
or U5514 (N_5514,N_2695,N_3782);
xnor U5515 (N_5515,N_4611,N_3127);
nor U5516 (N_5516,N_4674,N_3218);
nor U5517 (N_5517,N_3377,N_3996);
and U5518 (N_5518,N_4988,N_3114);
nor U5519 (N_5519,N_3027,N_3988);
nor U5520 (N_5520,N_3921,N_2816);
and U5521 (N_5521,N_2943,N_4593);
or U5522 (N_5522,N_4375,N_4826);
nand U5523 (N_5523,N_2847,N_4531);
nor U5524 (N_5524,N_4692,N_4112);
xnor U5525 (N_5525,N_2825,N_4204);
nor U5526 (N_5526,N_3812,N_4424);
or U5527 (N_5527,N_4509,N_4472);
xnor U5528 (N_5528,N_4208,N_3903);
nand U5529 (N_5529,N_2936,N_3258);
nand U5530 (N_5530,N_4719,N_3713);
nand U5531 (N_5531,N_4619,N_3273);
xnor U5532 (N_5532,N_3148,N_2557);
and U5533 (N_5533,N_2940,N_4647);
nand U5534 (N_5534,N_3231,N_3326);
and U5535 (N_5535,N_3906,N_4783);
and U5536 (N_5536,N_4642,N_4905);
nand U5537 (N_5537,N_3623,N_4044);
xor U5538 (N_5538,N_4819,N_3063);
and U5539 (N_5539,N_4233,N_2664);
xnor U5540 (N_5540,N_4346,N_3553);
and U5541 (N_5541,N_3161,N_3684);
and U5542 (N_5542,N_4597,N_4411);
xnor U5543 (N_5543,N_2753,N_2766);
or U5544 (N_5544,N_3779,N_4470);
or U5545 (N_5545,N_2818,N_4374);
and U5546 (N_5546,N_4600,N_2639);
nand U5547 (N_5547,N_3600,N_3374);
and U5548 (N_5548,N_4843,N_4854);
nor U5549 (N_5549,N_4501,N_2830);
nor U5550 (N_5550,N_3794,N_3891);
nand U5551 (N_5551,N_3626,N_4326);
nor U5552 (N_5552,N_4434,N_3773);
nand U5553 (N_5553,N_4902,N_3472);
or U5554 (N_5554,N_4085,N_3434);
or U5555 (N_5555,N_4522,N_2612);
nor U5556 (N_5556,N_2992,N_2538);
xor U5557 (N_5557,N_4210,N_3868);
nand U5558 (N_5558,N_2579,N_4887);
nor U5559 (N_5559,N_2769,N_4932);
xnor U5560 (N_5560,N_3290,N_4745);
and U5561 (N_5561,N_3024,N_3092);
or U5562 (N_5562,N_2638,N_4655);
or U5563 (N_5563,N_2613,N_3638);
nor U5564 (N_5564,N_3965,N_3170);
nor U5565 (N_5565,N_4592,N_4226);
nand U5566 (N_5566,N_4715,N_3866);
xnor U5567 (N_5567,N_4438,N_3270);
xnor U5568 (N_5568,N_4532,N_3405);
xor U5569 (N_5569,N_4606,N_3090);
and U5570 (N_5570,N_4768,N_4484);
and U5571 (N_5571,N_4133,N_3809);
xor U5572 (N_5572,N_3570,N_3590);
nand U5573 (N_5573,N_3469,N_3056);
xor U5574 (N_5574,N_4943,N_4361);
xor U5575 (N_5575,N_3938,N_4283);
nor U5576 (N_5576,N_3924,N_4870);
and U5577 (N_5577,N_4281,N_2931);
nor U5578 (N_5578,N_3361,N_2965);
nor U5579 (N_5579,N_3981,N_3134);
and U5580 (N_5580,N_4908,N_4450);
nor U5581 (N_5581,N_3396,N_3704);
and U5582 (N_5582,N_4248,N_3814);
xnor U5583 (N_5583,N_3808,N_4329);
and U5584 (N_5584,N_4161,N_2702);
nor U5585 (N_5585,N_4482,N_4609);
nor U5586 (N_5586,N_3399,N_4339);
and U5587 (N_5587,N_3083,N_3433);
nor U5588 (N_5588,N_3133,N_4069);
or U5589 (N_5589,N_2894,N_2747);
and U5590 (N_5590,N_3544,N_4698);
nor U5591 (N_5591,N_4486,N_2858);
or U5592 (N_5592,N_3934,N_4309);
xor U5593 (N_5593,N_4858,N_4307);
or U5594 (N_5594,N_4721,N_3084);
nand U5595 (N_5595,N_4617,N_4500);
xor U5596 (N_5596,N_3408,N_4499);
nand U5597 (N_5597,N_2576,N_4635);
nand U5598 (N_5598,N_2902,N_3667);
nor U5599 (N_5599,N_4382,N_2703);
nor U5600 (N_5600,N_2629,N_3815);
xnor U5601 (N_5601,N_4930,N_3639);
or U5602 (N_5602,N_4502,N_3051);
or U5603 (N_5603,N_2594,N_4190);
xor U5604 (N_5604,N_4011,N_3738);
and U5605 (N_5605,N_4613,N_3276);
nand U5606 (N_5606,N_2955,N_2660);
xor U5607 (N_5607,N_2860,N_4890);
xor U5608 (N_5608,N_3179,N_3633);
xnor U5609 (N_5609,N_3832,N_3004);
and U5610 (N_5610,N_2543,N_4108);
or U5611 (N_5611,N_3669,N_2913);
nor U5612 (N_5612,N_2722,N_2537);
nand U5613 (N_5613,N_2712,N_3053);
nor U5614 (N_5614,N_3087,N_3766);
and U5615 (N_5615,N_3049,N_4798);
nand U5616 (N_5616,N_4122,N_3725);
xor U5617 (N_5617,N_2759,N_3751);
or U5618 (N_5618,N_2674,N_4982);
and U5619 (N_5619,N_2698,N_2961);
and U5620 (N_5620,N_2859,N_2932);
or U5621 (N_5621,N_4682,N_4024);
xnor U5622 (N_5622,N_3678,N_3960);
or U5623 (N_5623,N_4767,N_4920);
nor U5624 (N_5624,N_4323,N_2668);
or U5625 (N_5625,N_4325,N_4406);
nor U5626 (N_5626,N_2778,N_4571);
xor U5627 (N_5627,N_3857,N_4043);
nor U5628 (N_5628,N_2529,N_4644);
nor U5629 (N_5629,N_2513,N_4646);
and U5630 (N_5630,N_4032,N_4761);
nor U5631 (N_5631,N_4396,N_2539);
or U5632 (N_5632,N_3709,N_4058);
nor U5633 (N_5633,N_3681,N_2726);
xnor U5634 (N_5634,N_3737,N_4525);
or U5635 (N_5635,N_4812,N_2640);
nand U5636 (N_5636,N_4019,N_3336);
or U5637 (N_5637,N_3515,N_4017);
nand U5638 (N_5638,N_3622,N_4313);
nand U5639 (N_5639,N_4710,N_4970);
nand U5640 (N_5640,N_3115,N_4777);
and U5641 (N_5641,N_4950,N_3487);
and U5642 (N_5642,N_3254,N_3020);
nand U5643 (N_5643,N_4872,N_2574);
or U5644 (N_5644,N_4497,N_3549);
nand U5645 (N_5645,N_4431,N_4727);
xor U5646 (N_5646,N_4160,N_4234);
and U5647 (N_5647,N_3695,N_2593);
xor U5648 (N_5648,N_4095,N_4973);
xor U5649 (N_5649,N_3085,N_3463);
nor U5650 (N_5650,N_3673,N_3909);
nand U5651 (N_5651,N_4660,N_4132);
and U5652 (N_5652,N_2731,N_4306);
and U5653 (N_5653,N_2734,N_2523);
nor U5654 (N_5654,N_4694,N_4831);
nand U5655 (N_5655,N_2879,N_4591);
and U5656 (N_5656,N_3729,N_4120);
or U5657 (N_5657,N_4127,N_4524);
xnor U5658 (N_5658,N_4688,N_2869);
or U5659 (N_5659,N_2954,N_3855);
nand U5660 (N_5660,N_3975,N_3407);
nand U5661 (N_5661,N_3680,N_3488);
nand U5662 (N_5662,N_4125,N_3697);
nor U5663 (N_5663,N_4119,N_3097);
or U5664 (N_5664,N_4222,N_3329);
xnor U5665 (N_5665,N_4882,N_3409);
nand U5666 (N_5666,N_2793,N_3331);
nand U5667 (N_5667,N_4463,N_3452);
or U5668 (N_5668,N_3164,N_3750);
nor U5669 (N_5669,N_3370,N_4551);
xnor U5670 (N_5670,N_3915,N_2667);
nor U5671 (N_5671,N_3160,N_2570);
nor U5672 (N_5672,N_4620,N_3689);
or U5673 (N_5673,N_4796,N_3688);
nand U5674 (N_5674,N_4806,N_2780);
nand U5675 (N_5675,N_4782,N_3858);
nand U5676 (N_5676,N_2630,N_4749);
nor U5677 (N_5677,N_4181,N_4967);
nor U5678 (N_5678,N_3963,N_3132);
or U5679 (N_5679,N_2541,N_2771);
xnor U5680 (N_5680,N_4928,N_2633);
and U5681 (N_5681,N_4128,N_3283);
and U5682 (N_5682,N_2854,N_3537);
or U5683 (N_5683,N_3699,N_2517);
and U5684 (N_5684,N_2634,N_3439);
and U5685 (N_5685,N_3703,N_3839);
nor U5686 (N_5686,N_2853,N_2875);
xnor U5687 (N_5687,N_4740,N_2823);
or U5688 (N_5688,N_4115,N_4047);
and U5689 (N_5689,N_2647,N_4071);
nor U5690 (N_5690,N_3504,N_3936);
nand U5691 (N_5691,N_4173,N_4113);
and U5692 (N_5692,N_4704,N_3265);
nand U5693 (N_5693,N_2507,N_2700);
nor U5694 (N_5694,N_3920,N_3573);
nor U5695 (N_5695,N_3122,N_4466);
and U5696 (N_5696,N_4544,N_4241);
and U5697 (N_5697,N_4587,N_3430);
nand U5698 (N_5698,N_4390,N_4899);
xor U5699 (N_5699,N_3232,N_3183);
nand U5700 (N_5700,N_2737,N_4062);
xnor U5701 (N_5701,N_3922,N_3404);
nor U5702 (N_5702,N_4263,N_2889);
nor U5703 (N_5703,N_3185,N_2768);
nand U5704 (N_5704,N_4848,N_4640);
or U5705 (N_5705,N_4145,N_4918);
or U5706 (N_5706,N_3599,N_4735);
and U5707 (N_5707,N_3074,N_4846);
nor U5708 (N_5708,N_3595,N_3781);
xnor U5709 (N_5709,N_4245,N_4770);
nor U5710 (N_5710,N_2957,N_4960);
and U5711 (N_5711,N_3197,N_4633);
and U5712 (N_5712,N_2885,N_3094);
nor U5713 (N_5713,N_4784,N_3457);
and U5714 (N_5714,N_3829,N_2964);
nand U5715 (N_5715,N_3078,N_2952);
or U5716 (N_5716,N_3518,N_2819);
xor U5717 (N_5717,N_4799,N_3883);
nand U5718 (N_5718,N_4624,N_2632);
nor U5719 (N_5719,N_3135,N_4748);
nor U5720 (N_5720,N_2807,N_3236);
or U5721 (N_5721,N_2914,N_3630);
nand U5722 (N_5722,N_4898,N_3443);
nand U5723 (N_5723,N_4016,N_3402);
nor U5724 (N_5724,N_3663,N_2725);
and U5725 (N_5725,N_3674,N_3107);
xor U5726 (N_5726,N_4752,N_3787);
and U5727 (N_5727,N_4892,N_4940);
xor U5728 (N_5728,N_2799,N_3180);
nand U5729 (N_5729,N_4572,N_4618);
nand U5730 (N_5730,N_2604,N_4852);
nor U5731 (N_5731,N_4909,N_3953);
or U5732 (N_5732,N_3898,N_4136);
nand U5733 (N_5733,N_3506,N_4168);
nor U5734 (N_5734,N_4013,N_3119);
xor U5735 (N_5735,N_3987,N_3899);
xor U5736 (N_5736,N_3335,N_4357);
and U5737 (N_5737,N_2861,N_3458);
or U5738 (N_5738,N_2794,N_2840);
and U5739 (N_5739,N_3171,N_4102);
or U5740 (N_5740,N_3349,N_2626);
nor U5741 (N_5741,N_4578,N_2844);
xnor U5742 (N_5742,N_3990,N_2550);
or U5743 (N_5743,N_4448,N_2848);
or U5744 (N_5744,N_3876,N_4445);
xor U5745 (N_5745,N_2568,N_4876);
nand U5746 (N_5746,N_3264,N_3436);
or U5747 (N_5747,N_3813,N_4052);
nor U5748 (N_5748,N_3191,N_4661);
nand U5749 (N_5749,N_3322,N_3066);
nand U5750 (N_5750,N_3539,N_3784);
nor U5751 (N_5751,N_4104,N_3467);
or U5752 (N_5752,N_3897,N_3702);
nand U5753 (N_5753,N_4224,N_2589);
xnor U5754 (N_5754,N_4063,N_2839);
and U5755 (N_5755,N_3627,N_3000);
xor U5756 (N_5756,N_4553,N_3227);
nor U5757 (N_5757,N_4803,N_3280);
or U5758 (N_5758,N_3372,N_2651);
and U5759 (N_5759,N_3819,N_3459);
xor U5760 (N_5760,N_4099,N_4825);
or U5761 (N_5761,N_3332,N_4691);
and U5762 (N_5762,N_3103,N_3864);
nor U5763 (N_5763,N_4488,N_4636);
xnor U5764 (N_5764,N_4413,N_4815);
nand U5765 (N_5765,N_3041,N_4962);
and U5766 (N_5766,N_3918,N_3431);
nand U5767 (N_5767,N_4517,N_4218);
nor U5768 (N_5768,N_4191,N_2873);
nand U5769 (N_5769,N_4295,N_3154);
or U5770 (N_5770,N_2867,N_2692);
or U5771 (N_5771,N_4958,N_4891);
nand U5772 (N_5772,N_3624,N_4795);
or U5773 (N_5773,N_4216,N_3499);
nor U5774 (N_5774,N_4343,N_4533);
or U5775 (N_5775,N_3234,N_4875);
xnor U5776 (N_5776,N_2705,N_4481);
nand U5777 (N_5777,N_3248,N_3869);
and U5778 (N_5778,N_4185,N_4440);
and U5779 (N_5779,N_4114,N_4009);
and U5780 (N_5780,N_2925,N_3653);
xor U5781 (N_5781,N_3047,N_2774);
or U5782 (N_5782,N_3598,N_4570);
nand U5783 (N_5783,N_4267,N_2673);
or U5784 (N_5784,N_3847,N_4240);
xnor U5785 (N_5785,N_3830,N_4791);
nand U5786 (N_5786,N_4851,N_3925);
nand U5787 (N_5787,N_3030,N_4207);
nor U5788 (N_5788,N_3108,N_4824);
xnor U5789 (N_5789,N_3425,N_4809);
nor U5790 (N_5790,N_3260,N_4547);
nor U5791 (N_5791,N_3050,N_2905);
or U5792 (N_5792,N_4310,N_3961);
xor U5793 (N_5793,N_2740,N_3211);
nor U5794 (N_5794,N_3574,N_3575);
nor U5795 (N_5795,N_4116,N_4087);
nand U5796 (N_5796,N_3239,N_3300);
and U5797 (N_5797,N_4367,N_4936);
nor U5798 (N_5798,N_3749,N_3278);
xor U5799 (N_5799,N_4203,N_4328);
xor U5800 (N_5800,N_4550,N_4746);
and U5801 (N_5801,N_2569,N_4847);
and U5802 (N_5802,N_4048,N_2751);
nand U5803 (N_5803,N_4139,N_2524);
nor U5804 (N_5804,N_3685,N_3345);
xor U5805 (N_5805,N_4124,N_4368);
nand U5806 (N_5806,N_2761,N_4474);
or U5807 (N_5807,N_4480,N_2729);
nor U5808 (N_5808,N_3105,N_2880);
or U5809 (N_5809,N_3118,N_3473);
and U5810 (N_5810,N_3173,N_4429);
or U5811 (N_5811,N_4834,N_3816);
and U5812 (N_5812,N_3346,N_3526);
or U5813 (N_5813,N_4669,N_3510);
xnor U5814 (N_5814,N_3292,N_4560);
nor U5815 (N_5815,N_4238,N_4534);
nor U5816 (N_5816,N_3907,N_3080);
or U5817 (N_5817,N_3799,N_4303);
or U5818 (N_5818,N_4457,N_3220);
xnor U5819 (N_5819,N_4649,N_4447);
nor U5820 (N_5820,N_4565,N_3519);
and U5821 (N_5821,N_3594,N_4452);
or U5822 (N_5822,N_2852,N_3672);
xor U5823 (N_5823,N_4991,N_4687);
xor U5824 (N_5824,N_3692,N_3880);
nor U5825 (N_5825,N_2910,N_4037);
xnor U5826 (N_5826,N_3286,N_4152);
nand U5827 (N_5827,N_2609,N_2947);
nand U5828 (N_5828,N_3754,N_3927);
and U5829 (N_5829,N_3645,N_4314);
xor U5830 (N_5830,N_3967,N_3683);
and U5831 (N_5831,N_3449,N_4612);
and U5832 (N_5832,N_2676,N_3522);
xnor U5833 (N_5833,N_3850,N_3230);
or U5834 (N_5834,N_4394,N_2689);
xnor U5835 (N_5835,N_2672,N_4742);
xor U5836 (N_5836,N_3604,N_3369);
and U5837 (N_5837,N_4716,N_2683);
or U5838 (N_5838,N_3101,N_4903);
and U5839 (N_5839,N_3042,N_4956);
nor U5840 (N_5840,N_3389,N_4332);
nor U5841 (N_5841,N_3511,N_4393);
nand U5842 (N_5842,N_4380,N_3308);
or U5843 (N_5843,N_4573,N_4703);
xor U5844 (N_5844,N_4387,N_4757);
or U5845 (N_5845,N_3700,N_2586);
or U5846 (N_5846,N_3546,N_2928);
xor U5847 (N_5847,N_2693,N_3670);
nor U5848 (N_5848,N_3215,N_3325);
xnor U5849 (N_5849,N_2988,N_3061);
or U5850 (N_5850,N_2694,N_3089);
xor U5851 (N_5851,N_3367,N_3146);
or U5852 (N_5852,N_2805,N_4414);
nand U5853 (N_5853,N_4163,N_4001);
and U5854 (N_5854,N_2838,N_4993);
nand U5855 (N_5855,N_2616,N_4059);
xor U5856 (N_5856,N_3011,N_2831);
and U5857 (N_5857,N_2784,N_4622);
nand U5858 (N_5858,N_4090,N_3288);
or U5859 (N_5859,N_4558,N_3295);
nand U5860 (N_5860,N_3340,N_4755);
xor U5861 (N_5861,N_4537,N_3055);
xnor U5862 (N_5862,N_2811,N_3438);
nand U5863 (N_5863,N_4731,N_2824);
or U5864 (N_5864,N_4708,N_4096);
nor U5865 (N_5865,N_3852,N_3662);
xor U5866 (N_5866,N_4623,N_3403);
xor U5867 (N_5867,N_4417,N_3297);
or U5868 (N_5868,N_4066,N_4494);
or U5869 (N_5869,N_2841,N_3475);
nor U5870 (N_5870,N_2997,N_2895);
or U5871 (N_5871,N_4333,N_3386);
nor U5872 (N_5872,N_4676,N_4270);
or U5873 (N_5873,N_2878,N_3129);
or U5874 (N_5874,N_4021,N_4589);
nand U5875 (N_5875,N_2688,N_4287);
or U5876 (N_5876,N_3418,N_4100);
or U5877 (N_5877,N_3760,N_3741);
and U5878 (N_5878,N_3315,N_4039);
or U5879 (N_5879,N_2764,N_4671);
or U5880 (N_5880,N_4641,N_3219);
xor U5881 (N_5881,N_4200,N_4175);
nor U5882 (N_5882,N_3417,N_3508);
nand U5883 (N_5883,N_4914,N_4418);
and U5884 (N_5884,N_3657,N_4789);
nor U5885 (N_5885,N_3644,N_2748);
nor U5886 (N_5886,N_3347,N_4556);
nand U5887 (N_5887,N_4353,N_4103);
nand U5888 (N_5888,N_3758,N_4584);
nand U5889 (N_5889,N_4643,N_4437);
nor U5890 (N_5890,N_2999,N_3485);
or U5891 (N_5891,N_3980,N_2611);
and U5892 (N_5892,N_3835,N_2509);
nor U5893 (N_5893,N_2903,N_4154);
or U5894 (N_5894,N_2649,N_3415);
xor U5895 (N_5895,N_3790,N_4228);
nand U5896 (N_5896,N_4086,N_4121);
and U5897 (N_5897,N_4051,N_3528);
xor U5898 (N_5898,N_2890,N_2506);
nand U5899 (N_5899,N_3611,N_4439);
and U5900 (N_5900,N_3006,N_4765);
or U5901 (N_5901,N_3194,N_4312);
nor U5902 (N_5902,N_4462,N_3979);
nand U5903 (N_5903,N_3390,N_2790);
or U5904 (N_5904,N_3834,N_4630);
xnor U5905 (N_5905,N_4446,N_3242);
xor U5906 (N_5906,N_4442,N_4045);
xor U5907 (N_5907,N_3579,N_4539);
nor U5908 (N_5908,N_3818,N_3992);
nor U5909 (N_5909,N_3872,N_4864);
nor U5910 (N_5910,N_2803,N_4421);
xnor U5911 (N_5911,N_3776,N_2663);
and U5912 (N_5912,N_2882,N_3919);
and U5913 (N_5913,N_2699,N_3224);
and U5914 (N_5914,N_2599,N_3109);
or U5915 (N_5915,N_3543,N_3319);
and U5916 (N_5916,N_4178,N_2939);
or U5917 (N_5917,N_2644,N_2916);
or U5918 (N_5918,N_2871,N_3395);
nor U5919 (N_5919,N_3952,N_3251);
nand U5920 (N_5920,N_4581,N_4552);
nor U5921 (N_5921,N_4880,N_2781);
nor U5922 (N_5922,N_3373,N_3188);
xor U5923 (N_5923,N_3312,N_3547);
or U5924 (N_5924,N_2716,N_4608);
and U5925 (N_5925,N_3716,N_2826);
and U5926 (N_5926,N_2696,N_4866);
nand U5927 (N_5927,N_4939,N_4025);
nand U5928 (N_5928,N_3560,N_3796);
xnor U5929 (N_5929,N_4485,N_3823);
nor U5930 (N_5930,N_3860,N_3168);
or U5931 (N_5931,N_4483,N_3424);
and U5932 (N_5932,N_2659,N_3856);
or U5933 (N_5933,N_2904,N_3905);
and U5934 (N_5934,N_4350,N_3712);
nand U5935 (N_5935,N_4519,N_2969);
nand U5936 (N_5936,N_3481,N_3636);
and U5937 (N_5937,N_3726,N_3172);
and U5938 (N_5938,N_4778,N_4135);
xor U5939 (N_5939,N_3339,N_2535);
and U5940 (N_5940,N_3268,N_4841);
xnor U5941 (N_5941,N_3828,N_2828);
or U5942 (N_5942,N_3465,N_3007);
xnor U5943 (N_5943,N_2575,N_2795);
nand U5944 (N_5944,N_2763,N_4068);
and U5945 (N_5945,N_2900,N_3746);
and U5946 (N_5946,N_3567,N_2960);
nand U5947 (N_5947,N_4467,N_3651);
xor U5948 (N_5948,N_4020,N_4251);
nor U5949 (N_5949,N_4596,N_4577);
and U5950 (N_5950,N_2973,N_4080);
nand U5951 (N_5951,N_4156,N_4162);
and U5952 (N_5952,N_2719,N_2730);
and U5953 (N_5953,N_3563,N_3968);
xor U5954 (N_5954,N_4926,N_3285);
nor U5955 (N_5955,N_3744,N_2892);
and U5956 (N_5956,N_4285,N_2906);
nor U5957 (N_5957,N_4014,N_3235);
or U5958 (N_5958,N_2708,N_3343);
nand U5959 (N_5959,N_2886,N_3535);
xnor U5960 (N_5960,N_3480,N_3203);
or U5961 (N_5961,N_4123,N_3321);
xnor U5962 (N_5962,N_4479,N_3588);
nor U5963 (N_5963,N_3126,N_2887);
xnor U5964 (N_5964,N_4639,N_3412);
nor U5965 (N_5965,N_2578,N_4916);
and U5966 (N_5966,N_3079,N_4879);
nor U5967 (N_5967,N_2796,N_4772);
or U5968 (N_5968,N_3677,N_4802);
xnor U5969 (N_5969,N_3908,N_3581);
or U5970 (N_5970,N_3351,N_2815);
nor U5971 (N_5971,N_2684,N_3354);
xnor U5972 (N_5972,N_4232,N_2720);
and U5973 (N_5973,N_4621,N_3169);
and U5974 (N_5974,N_2620,N_4645);
nand U5975 (N_5975,N_3014,N_4910);
nor U5976 (N_5976,N_3885,N_2788);
or U5977 (N_5977,N_3046,N_3724);
nor U5978 (N_5978,N_4971,N_2942);
and U5979 (N_5979,N_4625,N_3605);
xor U5980 (N_5980,N_4874,N_3043);
or U5981 (N_5981,N_2617,N_2948);
and U5982 (N_5982,N_2528,N_2678);
and U5983 (N_5983,N_4340,N_3956);
nor U5984 (N_5984,N_2618,N_4924);
nand U5985 (N_5985,N_3825,N_4476);
xnor U5986 (N_5986,N_4489,N_3005);
nand U5987 (N_5987,N_2603,N_3199);
and U5988 (N_5988,N_3538,N_4699);
and U5989 (N_5989,N_2598,N_3556);
nor U5990 (N_5990,N_4529,N_3464);
or U5991 (N_5991,N_4376,N_4142);
nor U5992 (N_5992,N_4884,N_4182);
nand U5993 (N_5993,N_2671,N_3202);
or U5994 (N_5994,N_3150,N_4712);
xnor U5995 (N_5995,N_2710,N_2911);
xnor U5996 (N_5996,N_3394,N_2915);
nor U5997 (N_5997,N_3973,N_4849);
or U5998 (N_5998,N_3044,N_3086);
or U5999 (N_5999,N_3032,N_4033);
nand U6000 (N_6000,N_4265,N_2735);
xnor U6001 (N_6001,N_3328,N_4072);
and U6002 (N_6002,N_3761,N_3849);
and U6003 (N_6003,N_4337,N_3034);
nand U6004 (N_6004,N_3878,N_3747);
or U6005 (N_6005,N_2642,N_3460);
and U6006 (N_6006,N_3629,N_4563);
or U6007 (N_6007,N_3091,N_2872);
and U6008 (N_6008,N_3706,N_4840);
xor U6009 (N_6009,N_2832,N_2775);
and U6010 (N_6010,N_3035,N_4061);
or U6011 (N_6011,N_4762,N_2770);
or U6012 (N_6012,N_3707,N_3664);
xnor U6013 (N_6013,N_4828,N_3682);
xnor U6014 (N_6014,N_2953,N_3284);
nor U6015 (N_6015,N_3410,N_4174);
nand U6016 (N_6016,N_4143,N_3887);
nand U6017 (N_6017,N_4057,N_4557);
and U6018 (N_6018,N_3867,N_4541);
nor U6019 (N_6019,N_3940,N_4126);
nor U6020 (N_6020,N_4008,N_2597);
and U6021 (N_6021,N_3247,N_2534);
xor U6022 (N_6022,N_3507,N_4990);
nor U6023 (N_6023,N_3718,N_4590);
nor U6024 (N_6024,N_4304,N_4830);
nand U6025 (N_6025,N_2792,N_4083);
xnor U6026 (N_6026,N_3002,N_4465);
or U6027 (N_6027,N_2921,N_3851);
or U6028 (N_6028,N_3116,N_3381);
and U6029 (N_6029,N_3048,N_3009);
xor U6030 (N_6030,N_4110,N_2898);
or U6031 (N_6031,N_4994,N_3128);
nand U6032 (N_6032,N_3736,N_4729);
or U6033 (N_6033,N_3561,N_4320);
and U6034 (N_6034,N_4308,N_4377);
nor U6035 (N_6035,N_4036,N_3446);
and U6036 (N_6036,N_4766,N_3826);
and U6037 (N_6037,N_3649,N_3201);
nor U6038 (N_6038,N_4559,N_3841);
nand U6039 (N_6039,N_4410,N_2949);
or U6040 (N_6040,N_2742,N_4574);
nand U6041 (N_6041,N_3104,N_4398);
or U6042 (N_6042,N_3440,N_2791);
or U6043 (N_6043,N_3145,N_4064);
nand U6044 (N_6044,N_4915,N_4568);
nor U6045 (N_6045,N_3072,N_3441);
xnor U6046 (N_6046,N_3221,N_3989);
nand U6047 (N_6047,N_2733,N_2608);
nor U6048 (N_6048,N_2874,N_3943);
nor U6049 (N_6049,N_4911,N_4404);
nand U6050 (N_6050,N_4951,N_4300);
xor U6051 (N_6051,N_3333,N_3798);
nand U6052 (N_6052,N_4794,N_3951);
or U6053 (N_6053,N_2863,N_4653);
or U6054 (N_6054,N_4034,N_2798);
and U6055 (N_6055,N_3863,N_4341);
nand U6056 (N_6056,N_3033,N_3324);
or U6057 (N_6057,N_3777,N_4723);
and U6058 (N_6058,N_3640,N_4775);
nor U6059 (N_6059,N_3976,N_4516);
nor U6060 (N_6060,N_2600,N_3620);
nand U6061 (N_6061,N_4166,N_4814);
nor U6062 (N_6062,N_3659,N_3831);
nand U6063 (N_6063,N_4056,N_2797);
nor U6064 (N_6064,N_3933,N_4508);
or U6065 (N_6065,N_3110,N_3734);
or U6066 (N_6066,N_2756,N_4901);
xnor U6067 (N_6067,N_3028,N_2518);
nor U6068 (N_6068,N_2627,N_4977);
xnor U6069 (N_6069,N_3250,N_3916);
or U6070 (N_6070,N_4503,N_3533);
nand U6071 (N_6071,N_4877,N_4869);
nor U6072 (N_6072,N_3062,N_2669);
nand U6073 (N_6073,N_4549,N_3728);
xor U6074 (N_6074,N_4921,N_3585);
and U6075 (N_6075,N_4697,N_2974);
and U6076 (N_6076,N_4602,N_4520);
or U6077 (N_6077,N_2749,N_3213);
nor U6078 (N_6078,N_4949,N_3745);
and U6079 (N_6079,N_2687,N_4315);
nor U6080 (N_6080,N_2893,N_2926);
and U6081 (N_6081,N_4131,N_3317);
xor U6082 (N_6082,N_3019,N_2515);
nand U6083 (N_6083,N_4696,N_2561);
xor U6084 (N_6084,N_3176,N_2619);
xor U6085 (N_6085,N_4507,N_4427);
nor U6086 (N_6086,N_4215,N_4235);
nor U6087 (N_6087,N_4863,N_4933);
or U6088 (N_6088,N_4231,N_3545);
or U6089 (N_6089,N_4526,N_4515);
and U6090 (N_6090,N_2715,N_4117);
or U6091 (N_6091,N_4823,N_2606);
or U6092 (N_6092,N_3591,N_4351);
nand U6093 (N_6093,N_3387,N_4615);
xor U6094 (N_6094,N_3593,N_3694);
nor U6095 (N_6095,N_2691,N_3977);
nand U6096 (N_6096,N_4807,N_4430);
xor U6097 (N_6097,N_3450,N_2813);
and U6098 (N_6098,N_4631,N_4773);
xor U6099 (N_6099,N_3882,N_2677);
nor U6100 (N_6100,N_4211,N_3995);
nor U6101 (N_6101,N_4258,N_3010);
or U6102 (N_6102,N_3564,N_4365);
and U6103 (N_6103,N_3778,N_3474);
nor U6104 (N_6104,N_3382,N_4941);
nor U6105 (N_6105,N_3398,N_2849);
nand U6106 (N_6106,N_4842,N_2743);
xor U6107 (N_6107,N_4186,N_4867);
or U6108 (N_6108,N_4046,N_4334);
nor U6109 (N_6109,N_3205,N_4985);
xor U6110 (N_6110,N_3143,N_3764);
or U6111 (N_6111,N_3073,N_3865);
and U6112 (N_6112,N_4734,N_2855);
nand U6113 (N_6113,N_2746,N_3192);
xnor U6114 (N_6114,N_3548,N_4744);
nand U6115 (N_6115,N_3206,N_3643);
or U6116 (N_6116,N_2755,N_3879);
nor U6117 (N_6117,N_3462,N_3748);
nor U6118 (N_6118,N_4268,N_4412);
nor U6119 (N_6119,N_4638,N_3421);
or U6120 (N_6120,N_3959,N_3619);
nand U6121 (N_6121,N_3310,N_4492);
xor U6122 (N_6122,N_4986,N_2713);
and U6123 (N_6123,N_2767,N_4302);
nand U6124 (N_6124,N_2511,N_3650);
nor U6125 (N_6125,N_4223,N_3675);
nor U6126 (N_6126,N_4352,N_3414);
nand U6127 (N_6127,N_3065,N_2624);
nand U6128 (N_6128,N_4428,N_3793);
nor U6129 (N_6129,N_4974,N_2868);
or U6130 (N_6130,N_4101,N_4397);
xnor U6131 (N_6131,N_2930,N_3671);
or U6132 (N_6132,N_3397,N_4074);
or U6133 (N_6133,N_3017,N_4379);
xnor U6134 (N_6134,N_4423,N_4839);
nand U6135 (N_6135,N_4569,N_4158);
and U6136 (N_6136,N_2652,N_2980);
nand U6137 (N_6137,N_3096,N_4405);
xor U6138 (N_6138,N_3121,N_3476);
nor U6139 (N_6139,N_4743,N_2772);
nor U6140 (N_6140,N_4681,N_4776);
and U6141 (N_6141,N_4167,N_4255);
nand U6142 (N_6142,N_3305,N_4244);
nand U6143 (N_6143,N_3859,N_4432);
nand U6144 (N_6144,N_3187,N_3789);
nand U6145 (N_6145,N_4239,N_3451);
or U6146 (N_6146,N_4833,N_4975);
nor U6147 (N_6147,N_2899,N_2827);
xor U6148 (N_6148,N_3550,N_4443);
xnor U6149 (N_6149,N_3261,N_4616);
or U6150 (N_6150,N_4229,N_4999);
or U6151 (N_6151,N_4055,N_3025);
nand U6152 (N_6152,N_4460,N_2724);
nand U6153 (N_6153,N_4249,N_2783);
nor U6154 (N_6154,N_3052,N_3294);
and U6155 (N_6155,N_3632,N_4473);
nand U6156 (N_6156,N_4137,N_2967);
nor U6157 (N_6157,N_3045,N_4348);
nor U6158 (N_6158,N_4035,N_2635);
or U6159 (N_6159,N_3873,N_3279);
nand U6160 (N_6160,N_2592,N_3584);
xnor U6161 (N_6161,N_4081,N_4654);
or U6162 (N_6162,N_4713,N_3617);
nor U6163 (N_6163,N_3993,N_2645);
and U6164 (N_6164,N_3341,N_4385);
nand U6165 (N_6165,N_3739,N_4392);
or U6166 (N_6166,N_3601,N_4193);
nor U6167 (N_6167,N_4756,N_3971);
and U6168 (N_6168,N_4662,N_4728);
and U6169 (N_6169,N_3804,N_4478);
nor U6170 (N_6170,N_3690,N_4318);
or U6171 (N_6171,N_3721,N_3023);
nand U6172 (N_6172,N_4172,N_3060);
nand U6173 (N_6173,N_3752,N_2615);
nand U6174 (N_6174,N_2547,N_3666);
xnor U6175 (N_6175,N_2558,N_4006);
nand U6176 (N_6176,N_4850,N_3156);
xor U6177 (N_6177,N_4324,N_3970);
nand U6178 (N_6178,N_4535,N_4747);
and U6179 (N_6179,N_4961,N_2544);
xor U6180 (N_6180,N_4471,N_3327);
and U6181 (N_6181,N_4422,N_3613);
nor U6182 (N_6182,N_2536,N_4769);
nand U6183 (N_6183,N_4416,N_3722);
nand U6184 (N_6184,N_2758,N_3811);
and U6185 (N_6185,N_3676,N_3912);
nor U6186 (N_6186,N_4750,N_2779);
and U6187 (N_6187,N_2526,N_4935);
or U6188 (N_6188,N_3435,N_2991);
nor U6189 (N_6189,N_3551,N_4264);
xnor U6190 (N_6190,N_3385,N_3240);
nor U6191 (N_6191,N_2503,N_2580);
nor U6192 (N_6192,N_3696,N_3196);
xor U6193 (N_6193,N_4362,N_4305);
nand U6194 (N_6194,N_4637,N_4027);
and U6195 (N_6195,N_2527,N_4089);
or U6196 (N_6196,N_3821,N_4023);
or U6197 (N_6197,N_3962,N_3845);
nor U6198 (N_6198,N_2786,N_2666);
and U6199 (N_6199,N_2937,N_2972);
and U6200 (N_6200,N_2661,N_3209);
xor U6201 (N_6201,N_2607,N_3775);
nor U6202 (N_6202,N_4092,N_4388);
or U6203 (N_6203,N_2814,N_3931);
nand U6204 (N_6204,N_2655,N_3106);
xor U6205 (N_6205,N_3318,N_4706);
and U6206 (N_6206,N_4399,N_3531);
xor U6207 (N_6207,N_3964,N_3566);
nor U6208 (N_6208,N_2675,N_4294);
xor U6209 (N_6209,N_3861,N_4859);
nand U6210 (N_6210,N_4073,N_3274);
xnor U6211 (N_6211,N_4598,N_4155);
nand U6212 (N_6212,N_4821,N_4060);
and U6213 (N_6213,N_3342,N_3576);
and U6214 (N_6214,N_2540,N_4321);
nor U6215 (N_6215,N_4007,N_3846);
nor U6216 (N_6216,N_4996,N_4093);
or U6217 (N_6217,N_4983,N_2690);
xnor U6218 (N_6218,N_2656,N_3502);
or U6219 (N_6219,N_3207,N_2883);
and U6220 (N_6220,N_3167,N_2977);
or U6221 (N_6221,N_3552,N_2810);
nor U6222 (N_6222,N_3226,N_3500);
or U6223 (N_6223,N_4889,N_4506);
and U6224 (N_6224,N_3455,N_4082);
and U6225 (N_6225,N_4989,N_4673);
nand U6226 (N_6226,N_4278,N_2686);
xor U6227 (N_6227,N_4378,N_4246);
and U6228 (N_6228,N_3558,N_4206);
nand U6229 (N_6229,N_3999,N_3785);
nand U6230 (N_6230,N_3892,N_2996);
or U6231 (N_6231,N_4845,N_4730);
xnor U6232 (N_6232,N_3944,N_4109);
nand U6233 (N_6233,N_4358,N_4272);
nand U6234 (N_6234,N_3557,N_4829);
xnor U6235 (N_6235,N_2554,N_4724);
xnor U6236 (N_6236,N_4906,N_3454);
xnor U6237 (N_6237,N_2525,N_4512);
nand U6238 (N_6238,N_3070,N_4942);
or U6239 (N_6239,N_4888,N_3423);
and U6240 (N_6240,N_3986,N_4969);
xnor U6241 (N_6241,N_3542,N_3824);
nor U6242 (N_6242,N_3376,N_3380);
or U6243 (N_6243,N_4042,N_2946);
or U6244 (N_6244,N_4657,N_2896);
and U6245 (N_6245,N_3937,N_4260);
nand U6246 (N_6246,N_4955,N_3400);
nand U6247 (N_6247,N_4490,N_4659);
xor U6248 (N_6248,N_3771,N_3320);
xnor U6249 (N_6249,N_3757,N_3820);
or U6250 (N_6250,N_4107,N_4139);
nor U6251 (N_6251,N_3353,N_4408);
nor U6252 (N_6252,N_4502,N_3490);
or U6253 (N_6253,N_4856,N_4722);
nor U6254 (N_6254,N_3592,N_2818);
nor U6255 (N_6255,N_4525,N_4708);
nor U6256 (N_6256,N_3758,N_2698);
xor U6257 (N_6257,N_2683,N_2836);
xnor U6258 (N_6258,N_3436,N_2893);
or U6259 (N_6259,N_3167,N_2956);
or U6260 (N_6260,N_3974,N_2711);
or U6261 (N_6261,N_2542,N_2527);
nand U6262 (N_6262,N_2744,N_3418);
xnor U6263 (N_6263,N_3206,N_4976);
nor U6264 (N_6264,N_4679,N_2661);
nor U6265 (N_6265,N_3696,N_4529);
or U6266 (N_6266,N_4758,N_4816);
and U6267 (N_6267,N_3339,N_2960);
and U6268 (N_6268,N_3088,N_3262);
xnor U6269 (N_6269,N_4997,N_4167);
nand U6270 (N_6270,N_2714,N_3572);
nor U6271 (N_6271,N_4066,N_3719);
nor U6272 (N_6272,N_4165,N_2900);
or U6273 (N_6273,N_2984,N_4134);
and U6274 (N_6274,N_2885,N_4977);
nand U6275 (N_6275,N_3732,N_3199);
nand U6276 (N_6276,N_4712,N_3461);
or U6277 (N_6277,N_4367,N_2865);
nand U6278 (N_6278,N_4308,N_4797);
nand U6279 (N_6279,N_4334,N_4908);
or U6280 (N_6280,N_4589,N_3991);
nor U6281 (N_6281,N_4410,N_4221);
nand U6282 (N_6282,N_2788,N_4001);
and U6283 (N_6283,N_4141,N_4096);
and U6284 (N_6284,N_3846,N_3942);
nor U6285 (N_6285,N_2539,N_4138);
and U6286 (N_6286,N_3006,N_2686);
xor U6287 (N_6287,N_2788,N_4319);
or U6288 (N_6288,N_3974,N_3610);
or U6289 (N_6289,N_3927,N_3007);
nor U6290 (N_6290,N_3416,N_4084);
nor U6291 (N_6291,N_3791,N_3640);
and U6292 (N_6292,N_3160,N_3205);
and U6293 (N_6293,N_3283,N_4456);
nand U6294 (N_6294,N_3708,N_2573);
or U6295 (N_6295,N_4385,N_2986);
xnor U6296 (N_6296,N_4390,N_2733);
xnor U6297 (N_6297,N_2939,N_3702);
and U6298 (N_6298,N_4273,N_2801);
xor U6299 (N_6299,N_4149,N_3028);
and U6300 (N_6300,N_3091,N_3147);
or U6301 (N_6301,N_3480,N_3252);
or U6302 (N_6302,N_4317,N_4809);
nand U6303 (N_6303,N_2963,N_4641);
and U6304 (N_6304,N_4121,N_4281);
and U6305 (N_6305,N_4049,N_3919);
and U6306 (N_6306,N_4062,N_3355);
or U6307 (N_6307,N_3813,N_2748);
nand U6308 (N_6308,N_3195,N_4007);
nor U6309 (N_6309,N_3114,N_4374);
nor U6310 (N_6310,N_2625,N_3168);
xor U6311 (N_6311,N_4952,N_4279);
xnor U6312 (N_6312,N_2507,N_4597);
nor U6313 (N_6313,N_4200,N_3417);
nand U6314 (N_6314,N_4963,N_4541);
or U6315 (N_6315,N_3624,N_3575);
xor U6316 (N_6316,N_4165,N_2997);
xnor U6317 (N_6317,N_3190,N_2969);
nor U6318 (N_6318,N_4195,N_2996);
xor U6319 (N_6319,N_3011,N_3590);
nor U6320 (N_6320,N_4178,N_4845);
xnor U6321 (N_6321,N_3252,N_3618);
nor U6322 (N_6322,N_3559,N_2865);
nand U6323 (N_6323,N_3578,N_4285);
or U6324 (N_6324,N_4184,N_4370);
nand U6325 (N_6325,N_2617,N_4243);
nand U6326 (N_6326,N_4634,N_4011);
nor U6327 (N_6327,N_4158,N_3913);
nor U6328 (N_6328,N_2650,N_3951);
and U6329 (N_6329,N_3491,N_3068);
and U6330 (N_6330,N_3183,N_3100);
and U6331 (N_6331,N_3223,N_4249);
and U6332 (N_6332,N_4822,N_4951);
xor U6333 (N_6333,N_4572,N_2636);
or U6334 (N_6334,N_3937,N_3134);
and U6335 (N_6335,N_3511,N_4545);
nor U6336 (N_6336,N_2993,N_3080);
nand U6337 (N_6337,N_3667,N_3908);
nand U6338 (N_6338,N_2572,N_2986);
or U6339 (N_6339,N_4689,N_3821);
or U6340 (N_6340,N_2507,N_2551);
nand U6341 (N_6341,N_3192,N_4052);
or U6342 (N_6342,N_3041,N_3990);
and U6343 (N_6343,N_2885,N_3626);
and U6344 (N_6344,N_3748,N_4280);
nor U6345 (N_6345,N_2773,N_3898);
nand U6346 (N_6346,N_3542,N_2971);
xor U6347 (N_6347,N_4037,N_4124);
or U6348 (N_6348,N_3717,N_3687);
nand U6349 (N_6349,N_4478,N_4830);
nand U6350 (N_6350,N_4751,N_4739);
xor U6351 (N_6351,N_4825,N_4264);
nor U6352 (N_6352,N_4092,N_2561);
nand U6353 (N_6353,N_4927,N_2826);
or U6354 (N_6354,N_3675,N_3530);
nand U6355 (N_6355,N_3464,N_3702);
nor U6356 (N_6356,N_4296,N_4505);
and U6357 (N_6357,N_3246,N_4823);
or U6358 (N_6358,N_2823,N_4472);
xnor U6359 (N_6359,N_3762,N_2996);
nor U6360 (N_6360,N_4544,N_2684);
and U6361 (N_6361,N_2561,N_2629);
xnor U6362 (N_6362,N_2627,N_3493);
xnor U6363 (N_6363,N_4060,N_4910);
nor U6364 (N_6364,N_3142,N_4929);
nor U6365 (N_6365,N_4032,N_2667);
and U6366 (N_6366,N_4823,N_3607);
and U6367 (N_6367,N_2638,N_3948);
and U6368 (N_6368,N_2799,N_4752);
xnor U6369 (N_6369,N_2794,N_3302);
or U6370 (N_6370,N_4254,N_4264);
nand U6371 (N_6371,N_3381,N_3132);
or U6372 (N_6372,N_3888,N_2968);
and U6373 (N_6373,N_3906,N_2614);
and U6374 (N_6374,N_3721,N_3015);
nor U6375 (N_6375,N_2897,N_3580);
nand U6376 (N_6376,N_4883,N_4252);
or U6377 (N_6377,N_3734,N_3997);
nand U6378 (N_6378,N_3829,N_3980);
and U6379 (N_6379,N_3849,N_3509);
nand U6380 (N_6380,N_4769,N_3342);
xnor U6381 (N_6381,N_4554,N_4547);
or U6382 (N_6382,N_4806,N_3005);
nand U6383 (N_6383,N_3780,N_3514);
xor U6384 (N_6384,N_3831,N_4562);
xor U6385 (N_6385,N_3057,N_3065);
nor U6386 (N_6386,N_4832,N_3485);
or U6387 (N_6387,N_3313,N_3970);
and U6388 (N_6388,N_4954,N_3889);
nand U6389 (N_6389,N_2652,N_3499);
nand U6390 (N_6390,N_2897,N_3247);
nand U6391 (N_6391,N_3521,N_4401);
or U6392 (N_6392,N_3333,N_3747);
nand U6393 (N_6393,N_3428,N_3158);
and U6394 (N_6394,N_3419,N_4075);
nand U6395 (N_6395,N_4745,N_4803);
nand U6396 (N_6396,N_3361,N_3463);
nor U6397 (N_6397,N_3658,N_4602);
or U6398 (N_6398,N_4533,N_3570);
or U6399 (N_6399,N_3675,N_4130);
nor U6400 (N_6400,N_3151,N_3333);
nor U6401 (N_6401,N_4222,N_3892);
or U6402 (N_6402,N_4387,N_3281);
or U6403 (N_6403,N_4668,N_2579);
nand U6404 (N_6404,N_2683,N_2897);
xnor U6405 (N_6405,N_4213,N_2637);
nor U6406 (N_6406,N_3258,N_4589);
or U6407 (N_6407,N_4158,N_4511);
and U6408 (N_6408,N_3375,N_4392);
and U6409 (N_6409,N_3049,N_4158);
nor U6410 (N_6410,N_2557,N_2912);
nor U6411 (N_6411,N_4973,N_4785);
nand U6412 (N_6412,N_2587,N_3099);
and U6413 (N_6413,N_4785,N_3050);
nand U6414 (N_6414,N_3450,N_4304);
xor U6415 (N_6415,N_4490,N_4994);
xnor U6416 (N_6416,N_3996,N_4922);
xor U6417 (N_6417,N_4341,N_3230);
and U6418 (N_6418,N_2936,N_4502);
xor U6419 (N_6419,N_3410,N_4138);
nor U6420 (N_6420,N_4344,N_2739);
or U6421 (N_6421,N_3491,N_4163);
nand U6422 (N_6422,N_2500,N_3589);
or U6423 (N_6423,N_4221,N_4739);
xnor U6424 (N_6424,N_4380,N_2767);
and U6425 (N_6425,N_4095,N_2971);
and U6426 (N_6426,N_3029,N_4641);
xnor U6427 (N_6427,N_3457,N_3610);
or U6428 (N_6428,N_3673,N_4395);
nor U6429 (N_6429,N_4028,N_3422);
nor U6430 (N_6430,N_4045,N_3748);
and U6431 (N_6431,N_3393,N_2903);
nor U6432 (N_6432,N_4299,N_3066);
xnor U6433 (N_6433,N_3667,N_3162);
or U6434 (N_6434,N_4344,N_3471);
nor U6435 (N_6435,N_2663,N_3936);
nor U6436 (N_6436,N_2712,N_2907);
xor U6437 (N_6437,N_3184,N_4918);
nand U6438 (N_6438,N_3208,N_4209);
nand U6439 (N_6439,N_3691,N_3396);
nor U6440 (N_6440,N_4017,N_3797);
and U6441 (N_6441,N_4019,N_3586);
and U6442 (N_6442,N_4916,N_3756);
xor U6443 (N_6443,N_3611,N_4953);
nor U6444 (N_6444,N_3647,N_4629);
nand U6445 (N_6445,N_4934,N_2820);
nand U6446 (N_6446,N_2979,N_4111);
nand U6447 (N_6447,N_2648,N_2846);
nand U6448 (N_6448,N_3339,N_2661);
and U6449 (N_6449,N_4687,N_3635);
nand U6450 (N_6450,N_4432,N_2969);
nor U6451 (N_6451,N_2821,N_3311);
nor U6452 (N_6452,N_3763,N_4364);
xnor U6453 (N_6453,N_4852,N_3788);
xnor U6454 (N_6454,N_4316,N_3113);
nor U6455 (N_6455,N_4631,N_2655);
nand U6456 (N_6456,N_4707,N_4817);
xnor U6457 (N_6457,N_2594,N_4419);
xnor U6458 (N_6458,N_2846,N_2574);
nor U6459 (N_6459,N_3996,N_3114);
or U6460 (N_6460,N_3176,N_2663);
nand U6461 (N_6461,N_4695,N_2907);
xor U6462 (N_6462,N_3835,N_3836);
or U6463 (N_6463,N_4909,N_3727);
and U6464 (N_6464,N_4322,N_2684);
nor U6465 (N_6465,N_4217,N_3089);
or U6466 (N_6466,N_4939,N_4537);
nand U6467 (N_6467,N_2825,N_4032);
xor U6468 (N_6468,N_4383,N_3038);
nand U6469 (N_6469,N_3036,N_3389);
nor U6470 (N_6470,N_3266,N_3087);
and U6471 (N_6471,N_3035,N_3640);
or U6472 (N_6472,N_2539,N_3336);
xor U6473 (N_6473,N_4275,N_2799);
xor U6474 (N_6474,N_3215,N_4075);
nor U6475 (N_6475,N_4542,N_4315);
nand U6476 (N_6476,N_4824,N_3373);
and U6477 (N_6477,N_4971,N_4196);
nand U6478 (N_6478,N_4927,N_4650);
nand U6479 (N_6479,N_4422,N_4119);
nand U6480 (N_6480,N_3261,N_4200);
xor U6481 (N_6481,N_4380,N_4030);
xor U6482 (N_6482,N_3081,N_4377);
or U6483 (N_6483,N_2609,N_3256);
xor U6484 (N_6484,N_4816,N_3127);
nor U6485 (N_6485,N_4512,N_4612);
or U6486 (N_6486,N_2831,N_4084);
nor U6487 (N_6487,N_3737,N_4259);
xnor U6488 (N_6488,N_4373,N_4831);
and U6489 (N_6489,N_4569,N_4701);
or U6490 (N_6490,N_3316,N_4841);
and U6491 (N_6491,N_4360,N_2594);
or U6492 (N_6492,N_3402,N_4074);
nor U6493 (N_6493,N_4574,N_2631);
and U6494 (N_6494,N_4740,N_2934);
or U6495 (N_6495,N_4478,N_2907);
nor U6496 (N_6496,N_4340,N_4911);
nor U6497 (N_6497,N_4321,N_4716);
xnor U6498 (N_6498,N_3373,N_3715);
or U6499 (N_6499,N_4138,N_2588);
nor U6500 (N_6500,N_4397,N_3004);
xor U6501 (N_6501,N_4443,N_3665);
nand U6502 (N_6502,N_3259,N_3591);
and U6503 (N_6503,N_2997,N_2976);
nor U6504 (N_6504,N_4045,N_3613);
xor U6505 (N_6505,N_4954,N_3229);
nand U6506 (N_6506,N_4459,N_4144);
nor U6507 (N_6507,N_4450,N_4362);
nand U6508 (N_6508,N_3421,N_2940);
nand U6509 (N_6509,N_4982,N_3487);
nor U6510 (N_6510,N_3713,N_4783);
xnor U6511 (N_6511,N_3884,N_3844);
nand U6512 (N_6512,N_4095,N_2776);
nor U6513 (N_6513,N_3253,N_4117);
nor U6514 (N_6514,N_4080,N_3298);
nor U6515 (N_6515,N_2802,N_3478);
or U6516 (N_6516,N_2746,N_3558);
nor U6517 (N_6517,N_3239,N_2711);
and U6518 (N_6518,N_4406,N_4698);
and U6519 (N_6519,N_3177,N_3478);
nand U6520 (N_6520,N_3177,N_3010);
and U6521 (N_6521,N_2812,N_3347);
or U6522 (N_6522,N_3406,N_3146);
nand U6523 (N_6523,N_3424,N_3948);
nor U6524 (N_6524,N_2898,N_3216);
nand U6525 (N_6525,N_3003,N_4972);
nand U6526 (N_6526,N_4265,N_2784);
or U6527 (N_6527,N_4624,N_2892);
nand U6528 (N_6528,N_3407,N_4640);
nor U6529 (N_6529,N_3954,N_3556);
xnor U6530 (N_6530,N_3940,N_4081);
nand U6531 (N_6531,N_4697,N_3531);
or U6532 (N_6532,N_3843,N_4437);
nor U6533 (N_6533,N_2624,N_3586);
or U6534 (N_6534,N_2733,N_4662);
nand U6535 (N_6535,N_3456,N_3254);
nor U6536 (N_6536,N_4956,N_2635);
and U6537 (N_6537,N_3646,N_3875);
xnor U6538 (N_6538,N_4468,N_4872);
nor U6539 (N_6539,N_2878,N_3753);
and U6540 (N_6540,N_4120,N_4190);
nand U6541 (N_6541,N_3040,N_4160);
or U6542 (N_6542,N_4188,N_3010);
and U6543 (N_6543,N_2521,N_3018);
xor U6544 (N_6544,N_3669,N_4911);
nor U6545 (N_6545,N_3477,N_4152);
xnor U6546 (N_6546,N_2504,N_4646);
xnor U6547 (N_6547,N_4660,N_3138);
and U6548 (N_6548,N_2905,N_3173);
nand U6549 (N_6549,N_3635,N_3150);
xor U6550 (N_6550,N_3556,N_3065);
or U6551 (N_6551,N_3338,N_3203);
or U6552 (N_6552,N_2853,N_4329);
or U6553 (N_6553,N_4526,N_4701);
nand U6554 (N_6554,N_3782,N_2775);
or U6555 (N_6555,N_3963,N_2591);
and U6556 (N_6556,N_3938,N_2805);
xnor U6557 (N_6557,N_4770,N_3237);
xnor U6558 (N_6558,N_4615,N_4045);
nor U6559 (N_6559,N_4402,N_2539);
xnor U6560 (N_6560,N_3465,N_2988);
or U6561 (N_6561,N_3761,N_3210);
xor U6562 (N_6562,N_3600,N_4977);
or U6563 (N_6563,N_4036,N_4591);
and U6564 (N_6564,N_4430,N_2862);
nor U6565 (N_6565,N_3342,N_3719);
xnor U6566 (N_6566,N_2985,N_3259);
nand U6567 (N_6567,N_3112,N_2533);
nand U6568 (N_6568,N_2598,N_2591);
or U6569 (N_6569,N_3071,N_3510);
xnor U6570 (N_6570,N_3728,N_2633);
or U6571 (N_6571,N_3056,N_3253);
nor U6572 (N_6572,N_4723,N_4900);
nand U6573 (N_6573,N_2964,N_3337);
nand U6574 (N_6574,N_3579,N_2715);
nand U6575 (N_6575,N_4211,N_2900);
or U6576 (N_6576,N_3859,N_4415);
nor U6577 (N_6577,N_4271,N_2736);
and U6578 (N_6578,N_3995,N_3773);
and U6579 (N_6579,N_2983,N_4129);
or U6580 (N_6580,N_3019,N_4577);
nand U6581 (N_6581,N_2585,N_4946);
nor U6582 (N_6582,N_2909,N_3724);
xnor U6583 (N_6583,N_4848,N_3743);
and U6584 (N_6584,N_3686,N_4767);
and U6585 (N_6585,N_3162,N_3636);
and U6586 (N_6586,N_3063,N_2769);
and U6587 (N_6587,N_3768,N_3326);
and U6588 (N_6588,N_2884,N_4507);
nor U6589 (N_6589,N_3392,N_2918);
or U6590 (N_6590,N_4170,N_4378);
or U6591 (N_6591,N_4510,N_3234);
nand U6592 (N_6592,N_3288,N_2729);
nor U6593 (N_6593,N_3930,N_2679);
nand U6594 (N_6594,N_4033,N_3416);
or U6595 (N_6595,N_3586,N_4208);
nand U6596 (N_6596,N_3728,N_4087);
and U6597 (N_6597,N_3649,N_3051);
xor U6598 (N_6598,N_4313,N_3093);
xor U6599 (N_6599,N_4667,N_4675);
nor U6600 (N_6600,N_2846,N_3679);
and U6601 (N_6601,N_3101,N_4527);
nor U6602 (N_6602,N_4077,N_2690);
and U6603 (N_6603,N_4893,N_2769);
nand U6604 (N_6604,N_3883,N_4239);
and U6605 (N_6605,N_3678,N_4392);
xor U6606 (N_6606,N_3415,N_4149);
and U6607 (N_6607,N_3735,N_4244);
nand U6608 (N_6608,N_3818,N_4950);
or U6609 (N_6609,N_2577,N_4112);
or U6610 (N_6610,N_3562,N_3057);
or U6611 (N_6611,N_4372,N_3701);
nor U6612 (N_6612,N_4869,N_3092);
nand U6613 (N_6613,N_3381,N_2919);
xnor U6614 (N_6614,N_4042,N_2658);
or U6615 (N_6615,N_4079,N_3881);
nand U6616 (N_6616,N_3375,N_4483);
nand U6617 (N_6617,N_4291,N_4403);
nor U6618 (N_6618,N_2614,N_2724);
nand U6619 (N_6619,N_4976,N_4239);
nor U6620 (N_6620,N_3821,N_4985);
nor U6621 (N_6621,N_4325,N_4359);
nor U6622 (N_6622,N_4295,N_4485);
nor U6623 (N_6623,N_3142,N_3986);
and U6624 (N_6624,N_3533,N_4059);
and U6625 (N_6625,N_3813,N_4500);
xor U6626 (N_6626,N_2853,N_2911);
xnor U6627 (N_6627,N_4429,N_4708);
and U6628 (N_6628,N_3782,N_4289);
or U6629 (N_6629,N_4745,N_4654);
nand U6630 (N_6630,N_4697,N_3802);
xnor U6631 (N_6631,N_4887,N_4817);
nand U6632 (N_6632,N_2826,N_3554);
or U6633 (N_6633,N_2981,N_4358);
nor U6634 (N_6634,N_3942,N_2783);
or U6635 (N_6635,N_4667,N_2750);
or U6636 (N_6636,N_4399,N_2887);
and U6637 (N_6637,N_3968,N_3144);
nor U6638 (N_6638,N_3136,N_3828);
and U6639 (N_6639,N_4867,N_4148);
nand U6640 (N_6640,N_4190,N_3425);
and U6641 (N_6641,N_4352,N_4619);
xnor U6642 (N_6642,N_3277,N_2961);
and U6643 (N_6643,N_2736,N_3206);
xor U6644 (N_6644,N_3153,N_4132);
or U6645 (N_6645,N_4740,N_2761);
nor U6646 (N_6646,N_3130,N_2948);
nand U6647 (N_6647,N_3656,N_4070);
or U6648 (N_6648,N_2693,N_4179);
and U6649 (N_6649,N_2637,N_3533);
nand U6650 (N_6650,N_4276,N_3271);
nand U6651 (N_6651,N_3526,N_4291);
or U6652 (N_6652,N_4385,N_2641);
nand U6653 (N_6653,N_4780,N_3616);
and U6654 (N_6654,N_3553,N_3526);
nand U6655 (N_6655,N_4182,N_4004);
and U6656 (N_6656,N_3736,N_3846);
and U6657 (N_6657,N_4116,N_4555);
nor U6658 (N_6658,N_4646,N_4605);
nor U6659 (N_6659,N_3290,N_3338);
and U6660 (N_6660,N_4324,N_2557);
and U6661 (N_6661,N_3373,N_2557);
and U6662 (N_6662,N_4842,N_3425);
nor U6663 (N_6663,N_3829,N_2846);
nand U6664 (N_6664,N_2698,N_3832);
nand U6665 (N_6665,N_3888,N_2663);
xnor U6666 (N_6666,N_2615,N_3171);
xnor U6667 (N_6667,N_4094,N_4424);
or U6668 (N_6668,N_2511,N_4185);
or U6669 (N_6669,N_3262,N_3662);
or U6670 (N_6670,N_4200,N_3428);
xor U6671 (N_6671,N_4266,N_3562);
nor U6672 (N_6672,N_3684,N_4347);
nand U6673 (N_6673,N_3517,N_3386);
and U6674 (N_6674,N_3074,N_4412);
nor U6675 (N_6675,N_3616,N_3278);
and U6676 (N_6676,N_4518,N_4678);
or U6677 (N_6677,N_3552,N_4484);
nor U6678 (N_6678,N_3038,N_4538);
nor U6679 (N_6679,N_4148,N_2530);
nor U6680 (N_6680,N_2622,N_4765);
or U6681 (N_6681,N_2876,N_4382);
xor U6682 (N_6682,N_2689,N_3956);
nand U6683 (N_6683,N_2653,N_3642);
nand U6684 (N_6684,N_4882,N_2565);
xor U6685 (N_6685,N_3851,N_3255);
and U6686 (N_6686,N_3353,N_2737);
nor U6687 (N_6687,N_3921,N_4722);
nand U6688 (N_6688,N_2726,N_4695);
nor U6689 (N_6689,N_3915,N_4467);
xor U6690 (N_6690,N_4703,N_4977);
nor U6691 (N_6691,N_4593,N_4579);
xor U6692 (N_6692,N_3646,N_4881);
and U6693 (N_6693,N_3822,N_2923);
xnor U6694 (N_6694,N_4638,N_4706);
or U6695 (N_6695,N_2840,N_4684);
or U6696 (N_6696,N_4936,N_3716);
xnor U6697 (N_6697,N_3891,N_3012);
nand U6698 (N_6698,N_4196,N_4495);
nand U6699 (N_6699,N_3837,N_4781);
nand U6700 (N_6700,N_3398,N_2679);
nand U6701 (N_6701,N_3513,N_3491);
xnor U6702 (N_6702,N_3017,N_4511);
xnor U6703 (N_6703,N_2578,N_3500);
xnor U6704 (N_6704,N_2822,N_3404);
or U6705 (N_6705,N_4034,N_2935);
or U6706 (N_6706,N_3087,N_4076);
or U6707 (N_6707,N_2657,N_3304);
nand U6708 (N_6708,N_3994,N_4585);
xor U6709 (N_6709,N_3087,N_2912);
xor U6710 (N_6710,N_3616,N_3934);
nand U6711 (N_6711,N_4419,N_3664);
xor U6712 (N_6712,N_3889,N_3135);
nand U6713 (N_6713,N_3230,N_3241);
or U6714 (N_6714,N_3089,N_4618);
nand U6715 (N_6715,N_2572,N_4425);
xor U6716 (N_6716,N_4508,N_4951);
nor U6717 (N_6717,N_4690,N_4324);
and U6718 (N_6718,N_2756,N_3948);
nand U6719 (N_6719,N_2804,N_3338);
xor U6720 (N_6720,N_2826,N_2573);
xor U6721 (N_6721,N_2623,N_4973);
nand U6722 (N_6722,N_3495,N_3191);
nor U6723 (N_6723,N_3798,N_3840);
and U6724 (N_6724,N_2712,N_4287);
nand U6725 (N_6725,N_3611,N_3798);
xnor U6726 (N_6726,N_3314,N_3688);
nand U6727 (N_6727,N_2942,N_3331);
nor U6728 (N_6728,N_3599,N_2632);
or U6729 (N_6729,N_3487,N_3863);
nand U6730 (N_6730,N_3610,N_4666);
xnor U6731 (N_6731,N_4787,N_3222);
nand U6732 (N_6732,N_3004,N_2975);
nand U6733 (N_6733,N_4385,N_4118);
nor U6734 (N_6734,N_3048,N_3869);
nor U6735 (N_6735,N_3929,N_4256);
nand U6736 (N_6736,N_3346,N_4681);
nand U6737 (N_6737,N_2980,N_2791);
xnor U6738 (N_6738,N_4168,N_2696);
xnor U6739 (N_6739,N_3564,N_4225);
and U6740 (N_6740,N_4493,N_2647);
and U6741 (N_6741,N_3289,N_4730);
nand U6742 (N_6742,N_4913,N_3335);
nor U6743 (N_6743,N_2629,N_3617);
nand U6744 (N_6744,N_4420,N_3071);
and U6745 (N_6745,N_3489,N_3173);
nand U6746 (N_6746,N_3537,N_3113);
xor U6747 (N_6747,N_3049,N_4883);
and U6748 (N_6748,N_3043,N_3902);
nor U6749 (N_6749,N_4105,N_3898);
or U6750 (N_6750,N_3328,N_4449);
and U6751 (N_6751,N_4228,N_2734);
nand U6752 (N_6752,N_4019,N_4161);
nand U6753 (N_6753,N_4300,N_4722);
nand U6754 (N_6754,N_3429,N_4429);
or U6755 (N_6755,N_3173,N_4336);
xor U6756 (N_6756,N_4983,N_4337);
nand U6757 (N_6757,N_3597,N_3097);
nand U6758 (N_6758,N_2969,N_4730);
and U6759 (N_6759,N_4855,N_2648);
and U6760 (N_6760,N_2787,N_4136);
and U6761 (N_6761,N_3735,N_2904);
or U6762 (N_6762,N_4064,N_2783);
nand U6763 (N_6763,N_3575,N_2529);
nand U6764 (N_6764,N_4418,N_3247);
xor U6765 (N_6765,N_2938,N_4356);
and U6766 (N_6766,N_3970,N_3713);
nand U6767 (N_6767,N_3409,N_4124);
nor U6768 (N_6768,N_4132,N_3556);
nor U6769 (N_6769,N_2690,N_2827);
nand U6770 (N_6770,N_4472,N_4909);
nand U6771 (N_6771,N_4470,N_3841);
or U6772 (N_6772,N_4623,N_2920);
and U6773 (N_6773,N_4324,N_4789);
or U6774 (N_6774,N_4586,N_4258);
nand U6775 (N_6775,N_2733,N_3537);
or U6776 (N_6776,N_4866,N_4151);
or U6777 (N_6777,N_2691,N_3978);
xor U6778 (N_6778,N_3853,N_4915);
and U6779 (N_6779,N_2934,N_4954);
xor U6780 (N_6780,N_4516,N_2565);
and U6781 (N_6781,N_3355,N_4042);
and U6782 (N_6782,N_3092,N_3255);
or U6783 (N_6783,N_4719,N_3186);
nand U6784 (N_6784,N_2707,N_3158);
nor U6785 (N_6785,N_3657,N_2917);
nand U6786 (N_6786,N_3006,N_2659);
or U6787 (N_6787,N_3393,N_3019);
or U6788 (N_6788,N_4948,N_3597);
xor U6789 (N_6789,N_4759,N_3021);
xor U6790 (N_6790,N_3101,N_3342);
and U6791 (N_6791,N_3549,N_4548);
or U6792 (N_6792,N_4250,N_4406);
or U6793 (N_6793,N_4450,N_3652);
or U6794 (N_6794,N_3775,N_2639);
xnor U6795 (N_6795,N_3476,N_3066);
xor U6796 (N_6796,N_4501,N_2679);
nor U6797 (N_6797,N_3746,N_3693);
nand U6798 (N_6798,N_4348,N_2598);
or U6799 (N_6799,N_3215,N_3951);
nand U6800 (N_6800,N_3254,N_3403);
and U6801 (N_6801,N_4769,N_3320);
or U6802 (N_6802,N_2588,N_2618);
nor U6803 (N_6803,N_3137,N_4140);
or U6804 (N_6804,N_4151,N_4976);
nor U6805 (N_6805,N_4337,N_4905);
and U6806 (N_6806,N_3194,N_3020);
xor U6807 (N_6807,N_4437,N_4607);
xor U6808 (N_6808,N_4374,N_3634);
nand U6809 (N_6809,N_4795,N_2810);
xor U6810 (N_6810,N_3262,N_3430);
or U6811 (N_6811,N_3838,N_4687);
and U6812 (N_6812,N_4525,N_4811);
and U6813 (N_6813,N_4323,N_4710);
and U6814 (N_6814,N_3949,N_4153);
xnor U6815 (N_6815,N_3405,N_4298);
xor U6816 (N_6816,N_4788,N_3448);
xnor U6817 (N_6817,N_2713,N_4707);
xnor U6818 (N_6818,N_2739,N_2874);
or U6819 (N_6819,N_4850,N_4385);
and U6820 (N_6820,N_4615,N_3964);
nand U6821 (N_6821,N_3082,N_2757);
nand U6822 (N_6822,N_3291,N_3033);
or U6823 (N_6823,N_4354,N_2519);
nand U6824 (N_6824,N_2886,N_4007);
nor U6825 (N_6825,N_2816,N_2646);
nand U6826 (N_6826,N_4441,N_2667);
and U6827 (N_6827,N_4740,N_3576);
and U6828 (N_6828,N_4113,N_3431);
nor U6829 (N_6829,N_4086,N_4588);
or U6830 (N_6830,N_2762,N_3262);
nor U6831 (N_6831,N_3930,N_2610);
nor U6832 (N_6832,N_3255,N_3311);
or U6833 (N_6833,N_4123,N_3896);
or U6834 (N_6834,N_4182,N_4858);
nand U6835 (N_6835,N_4409,N_4754);
xor U6836 (N_6836,N_2835,N_3837);
nand U6837 (N_6837,N_4255,N_3252);
nand U6838 (N_6838,N_3778,N_4061);
xnor U6839 (N_6839,N_4050,N_3961);
or U6840 (N_6840,N_3156,N_3427);
xor U6841 (N_6841,N_3567,N_4162);
or U6842 (N_6842,N_4800,N_3281);
or U6843 (N_6843,N_4522,N_3022);
and U6844 (N_6844,N_3186,N_4669);
and U6845 (N_6845,N_3924,N_4184);
and U6846 (N_6846,N_4999,N_2769);
xor U6847 (N_6847,N_4117,N_3319);
and U6848 (N_6848,N_3326,N_4944);
nand U6849 (N_6849,N_2747,N_3809);
and U6850 (N_6850,N_2639,N_3021);
and U6851 (N_6851,N_3694,N_4312);
xnor U6852 (N_6852,N_3135,N_4064);
and U6853 (N_6853,N_3676,N_4287);
nand U6854 (N_6854,N_2515,N_2904);
or U6855 (N_6855,N_3798,N_2970);
nand U6856 (N_6856,N_3990,N_4740);
xor U6857 (N_6857,N_3741,N_3415);
xnor U6858 (N_6858,N_4729,N_3451);
and U6859 (N_6859,N_3874,N_4318);
nor U6860 (N_6860,N_2972,N_3679);
xnor U6861 (N_6861,N_2810,N_4868);
or U6862 (N_6862,N_3856,N_3138);
xor U6863 (N_6863,N_4318,N_3650);
xor U6864 (N_6864,N_2767,N_4964);
xnor U6865 (N_6865,N_3767,N_3392);
nor U6866 (N_6866,N_4956,N_2623);
and U6867 (N_6867,N_4924,N_3518);
nand U6868 (N_6868,N_4507,N_4530);
and U6869 (N_6869,N_2554,N_3936);
nor U6870 (N_6870,N_3489,N_4003);
nor U6871 (N_6871,N_3902,N_3649);
and U6872 (N_6872,N_3947,N_4845);
and U6873 (N_6873,N_3186,N_2567);
or U6874 (N_6874,N_4885,N_3070);
nand U6875 (N_6875,N_4514,N_3253);
and U6876 (N_6876,N_3535,N_2571);
nand U6877 (N_6877,N_4422,N_4699);
nand U6878 (N_6878,N_4181,N_2903);
nor U6879 (N_6879,N_2634,N_4049);
and U6880 (N_6880,N_2530,N_2808);
or U6881 (N_6881,N_4539,N_4458);
nor U6882 (N_6882,N_2788,N_4903);
nand U6883 (N_6883,N_3918,N_4495);
and U6884 (N_6884,N_4314,N_4218);
xor U6885 (N_6885,N_3088,N_3515);
or U6886 (N_6886,N_3238,N_3787);
nor U6887 (N_6887,N_3927,N_2778);
xor U6888 (N_6888,N_3886,N_2949);
or U6889 (N_6889,N_3396,N_3120);
or U6890 (N_6890,N_3684,N_3547);
nor U6891 (N_6891,N_2652,N_3419);
nor U6892 (N_6892,N_3757,N_2682);
or U6893 (N_6893,N_3607,N_3393);
nand U6894 (N_6894,N_4340,N_4536);
nor U6895 (N_6895,N_4773,N_4058);
xnor U6896 (N_6896,N_3042,N_3047);
nand U6897 (N_6897,N_3429,N_4047);
or U6898 (N_6898,N_2708,N_4876);
or U6899 (N_6899,N_4373,N_3382);
nor U6900 (N_6900,N_4404,N_3494);
nand U6901 (N_6901,N_3016,N_2773);
and U6902 (N_6902,N_2947,N_2565);
nand U6903 (N_6903,N_2820,N_3778);
xnor U6904 (N_6904,N_3211,N_3509);
and U6905 (N_6905,N_3627,N_3982);
and U6906 (N_6906,N_4051,N_4582);
nor U6907 (N_6907,N_4949,N_2911);
nor U6908 (N_6908,N_2635,N_3923);
nor U6909 (N_6909,N_4107,N_4779);
nand U6910 (N_6910,N_2793,N_3881);
nand U6911 (N_6911,N_4876,N_4851);
or U6912 (N_6912,N_4668,N_3063);
or U6913 (N_6913,N_4016,N_2602);
nand U6914 (N_6914,N_4738,N_3580);
nor U6915 (N_6915,N_2618,N_4865);
or U6916 (N_6916,N_2529,N_2794);
or U6917 (N_6917,N_4650,N_4960);
nor U6918 (N_6918,N_3869,N_2686);
nand U6919 (N_6919,N_4601,N_3337);
and U6920 (N_6920,N_3281,N_4453);
nor U6921 (N_6921,N_4687,N_2520);
xor U6922 (N_6922,N_4444,N_4174);
or U6923 (N_6923,N_4674,N_3082);
nand U6924 (N_6924,N_3907,N_2775);
or U6925 (N_6925,N_3834,N_4137);
nand U6926 (N_6926,N_2630,N_4188);
nor U6927 (N_6927,N_4353,N_3642);
nor U6928 (N_6928,N_4598,N_3129);
xor U6929 (N_6929,N_4846,N_3245);
xnor U6930 (N_6930,N_4702,N_4346);
nand U6931 (N_6931,N_3342,N_4982);
and U6932 (N_6932,N_4545,N_4009);
or U6933 (N_6933,N_2727,N_3038);
xor U6934 (N_6934,N_2650,N_3158);
nand U6935 (N_6935,N_2521,N_2523);
xnor U6936 (N_6936,N_4345,N_2838);
nor U6937 (N_6937,N_4593,N_4638);
or U6938 (N_6938,N_3237,N_2610);
nand U6939 (N_6939,N_4889,N_4495);
or U6940 (N_6940,N_4042,N_4854);
xnor U6941 (N_6941,N_3575,N_3194);
and U6942 (N_6942,N_3482,N_4122);
or U6943 (N_6943,N_4724,N_2973);
nand U6944 (N_6944,N_3384,N_3573);
xnor U6945 (N_6945,N_4005,N_3155);
xor U6946 (N_6946,N_4381,N_4983);
nand U6947 (N_6947,N_2999,N_3499);
nand U6948 (N_6948,N_3423,N_2572);
nor U6949 (N_6949,N_3370,N_4918);
nand U6950 (N_6950,N_4800,N_2679);
xor U6951 (N_6951,N_3821,N_2634);
nand U6952 (N_6952,N_3231,N_4738);
or U6953 (N_6953,N_2715,N_3330);
nand U6954 (N_6954,N_3195,N_3591);
nor U6955 (N_6955,N_2744,N_4040);
nor U6956 (N_6956,N_3221,N_2908);
or U6957 (N_6957,N_3690,N_3404);
and U6958 (N_6958,N_4252,N_3748);
and U6959 (N_6959,N_4527,N_2736);
and U6960 (N_6960,N_2718,N_3809);
or U6961 (N_6961,N_3121,N_4606);
nor U6962 (N_6962,N_3427,N_2660);
and U6963 (N_6963,N_2561,N_4238);
or U6964 (N_6964,N_3869,N_4116);
or U6965 (N_6965,N_2558,N_2674);
nand U6966 (N_6966,N_4334,N_4877);
nor U6967 (N_6967,N_3374,N_2685);
or U6968 (N_6968,N_3120,N_2826);
nand U6969 (N_6969,N_3363,N_4571);
xnor U6970 (N_6970,N_3235,N_4343);
nor U6971 (N_6971,N_3897,N_3366);
xor U6972 (N_6972,N_3116,N_4808);
nor U6973 (N_6973,N_3263,N_3909);
nand U6974 (N_6974,N_4766,N_4068);
nand U6975 (N_6975,N_4030,N_3504);
and U6976 (N_6976,N_3460,N_3232);
nor U6977 (N_6977,N_3151,N_3414);
nor U6978 (N_6978,N_3269,N_2579);
or U6979 (N_6979,N_3435,N_3936);
and U6980 (N_6980,N_2732,N_3782);
and U6981 (N_6981,N_4997,N_3751);
nor U6982 (N_6982,N_4116,N_4839);
and U6983 (N_6983,N_3108,N_3736);
nand U6984 (N_6984,N_3797,N_4532);
nor U6985 (N_6985,N_2834,N_4991);
and U6986 (N_6986,N_4558,N_2763);
nor U6987 (N_6987,N_3924,N_2559);
nor U6988 (N_6988,N_4181,N_3868);
and U6989 (N_6989,N_3766,N_4330);
xnor U6990 (N_6990,N_4784,N_4019);
nor U6991 (N_6991,N_2887,N_4992);
xor U6992 (N_6992,N_2539,N_3416);
and U6993 (N_6993,N_3788,N_3218);
or U6994 (N_6994,N_3474,N_2529);
xor U6995 (N_6995,N_2871,N_4723);
and U6996 (N_6996,N_3081,N_3759);
nand U6997 (N_6997,N_4620,N_2810);
or U6998 (N_6998,N_3422,N_3396);
nor U6999 (N_6999,N_2897,N_4378);
and U7000 (N_7000,N_4130,N_4143);
xnor U7001 (N_7001,N_3408,N_4354);
and U7002 (N_7002,N_2512,N_4970);
nand U7003 (N_7003,N_3685,N_3985);
or U7004 (N_7004,N_4542,N_2556);
or U7005 (N_7005,N_3690,N_4098);
nor U7006 (N_7006,N_2544,N_4743);
nor U7007 (N_7007,N_4009,N_4572);
nor U7008 (N_7008,N_2829,N_4737);
or U7009 (N_7009,N_3493,N_4623);
or U7010 (N_7010,N_4877,N_3091);
nand U7011 (N_7011,N_4969,N_3624);
nor U7012 (N_7012,N_4070,N_3964);
xnor U7013 (N_7013,N_2958,N_3233);
xor U7014 (N_7014,N_4576,N_4326);
xor U7015 (N_7015,N_4396,N_4048);
nor U7016 (N_7016,N_4864,N_4475);
xor U7017 (N_7017,N_2865,N_2728);
nor U7018 (N_7018,N_3271,N_4008);
xnor U7019 (N_7019,N_4233,N_4146);
nand U7020 (N_7020,N_4703,N_3969);
xor U7021 (N_7021,N_3256,N_4234);
nand U7022 (N_7022,N_4482,N_2766);
or U7023 (N_7023,N_4034,N_3236);
or U7024 (N_7024,N_4605,N_2832);
and U7025 (N_7025,N_4491,N_3545);
and U7026 (N_7026,N_4428,N_3808);
nor U7027 (N_7027,N_3518,N_3230);
xor U7028 (N_7028,N_4166,N_3119);
and U7029 (N_7029,N_3143,N_4804);
and U7030 (N_7030,N_2820,N_4190);
and U7031 (N_7031,N_3890,N_3144);
nor U7032 (N_7032,N_2739,N_4221);
or U7033 (N_7033,N_4274,N_4527);
xnor U7034 (N_7034,N_2930,N_4848);
nand U7035 (N_7035,N_3178,N_2689);
xor U7036 (N_7036,N_4311,N_3683);
nor U7037 (N_7037,N_4301,N_3020);
nand U7038 (N_7038,N_4683,N_4299);
or U7039 (N_7039,N_2559,N_4721);
xor U7040 (N_7040,N_4923,N_4528);
xor U7041 (N_7041,N_3173,N_4333);
or U7042 (N_7042,N_3802,N_3273);
nand U7043 (N_7043,N_3349,N_3564);
nor U7044 (N_7044,N_4373,N_4744);
nor U7045 (N_7045,N_2549,N_4546);
nor U7046 (N_7046,N_2533,N_3799);
nand U7047 (N_7047,N_4169,N_3340);
xor U7048 (N_7048,N_3576,N_2909);
and U7049 (N_7049,N_2997,N_3095);
and U7050 (N_7050,N_2931,N_4349);
or U7051 (N_7051,N_3239,N_3581);
nor U7052 (N_7052,N_4714,N_4921);
nand U7053 (N_7053,N_4165,N_4458);
and U7054 (N_7054,N_4454,N_2581);
or U7055 (N_7055,N_4718,N_3212);
nor U7056 (N_7056,N_4444,N_4257);
or U7057 (N_7057,N_2795,N_3027);
and U7058 (N_7058,N_3362,N_3870);
and U7059 (N_7059,N_2973,N_4415);
nand U7060 (N_7060,N_3729,N_4634);
nor U7061 (N_7061,N_4218,N_2861);
or U7062 (N_7062,N_3268,N_3353);
and U7063 (N_7063,N_2518,N_3603);
xor U7064 (N_7064,N_2808,N_4426);
nor U7065 (N_7065,N_4154,N_4755);
nand U7066 (N_7066,N_4273,N_3899);
and U7067 (N_7067,N_4195,N_3828);
and U7068 (N_7068,N_2556,N_4433);
or U7069 (N_7069,N_4236,N_4844);
xnor U7070 (N_7070,N_3938,N_3026);
nand U7071 (N_7071,N_4656,N_3412);
nor U7072 (N_7072,N_4973,N_4581);
xor U7073 (N_7073,N_4864,N_4300);
and U7074 (N_7074,N_3032,N_3035);
nand U7075 (N_7075,N_2560,N_4017);
and U7076 (N_7076,N_4035,N_4083);
nand U7077 (N_7077,N_4710,N_4195);
or U7078 (N_7078,N_3095,N_3271);
xnor U7079 (N_7079,N_2540,N_2724);
or U7080 (N_7080,N_2558,N_4740);
and U7081 (N_7081,N_3717,N_3139);
nor U7082 (N_7082,N_3537,N_3552);
nor U7083 (N_7083,N_4633,N_4122);
xor U7084 (N_7084,N_3389,N_4230);
nand U7085 (N_7085,N_2730,N_2763);
xnor U7086 (N_7086,N_3085,N_4774);
and U7087 (N_7087,N_4437,N_2949);
and U7088 (N_7088,N_4145,N_2534);
nand U7089 (N_7089,N_2926,N_3092);
or U7090 (N_7090,N_4630,N_4178);
xnor U7091 (N_7091,N_4098,N_3600);
nor U7092 (N_7092,N_3051,N_4001);
or U7093 (N_7093,N_2749,N_3478);
nand U7094 (N_7094,N_3813,N_3768);
nand U7095 (N_7095,N_3553,N_3414);
nand U7096 (N_7096,N_3701,N_2999);
or U7097 (N_7097,N_3476,N_4526);
and U7098 (N_7098,N_4830,N_3858);
or U7099 (N_7099,N_3747,N_2538);
nor U7100 (N_7100,N_3742,N_4613);
nor U7101 (N_7101,N_2903,N_4139);
xor U7102 (N_7102,N_3258,N_4018);
nor U7103 (N_7103,N_4160,N_4999);
and U7104 (N_7104,N_4804,N_4115);
nor U7105 (N_7105,N_3502,N_4857);
nor U7106 (N_7106,N_3572,N_4443);
and U7107 (N_7107,N_3818,N_4418);
and U7108 (N_7108,N_2668,N_4301);
nor U7109 (N_7109,N_3339,N_4034);
xnor U7110 (N_7110,N_3536,N_3931);
xor U7111 (N_7111,N_4694,N_3345);
nor U7112 (N_7112,N_3912,N_2676);
or U7113 (N_7113,N_3906,N_4758);
nor U7114 (N_7114,N_4048,N_4910);
or U7115 (N_7115,N_4336,N_3941);
nor U7116 (N_7116,N_2918,N_3024);
nand U7117 (N_7117,N_2765,N_2661);
xor U7118 (N_7118,N_4597,N_3217);
or U7119 (N_7119,N_3888,N_4364);
nor U7120 (N_7120,N_4793,N_4101);
nor U7121 (N_7121,N_4655,N_3363);
and U7122 (N_7122,N_3275,N_4988);
xor U7123 (N_7123,N_3036,N_3330);
nor U7124 (N_7124,N_4854,N_4824);
nand U7125 (N_7125,N_2548,N_3235);
nor U7126 (N_7126,N_4426,N_4951);
or U7127 (N_7127,N_4255,N_4359);
nor U7128 (N_7128,N_4591,N_4854);
or U7129 (N_7129,N_4618,N_3504);
nor U7130 (N_7130,N_2636,N_3558);
or U7131 (N_7131,N_4720,N_2767);
nor U7132 (N_7132,N_2835,N_4092);
nor U7133 (N_7133,N_4182,N_2944);
or U7134 (N_7134,N_3984,N_3831);
nand U7135 (N_7135,N_2804,N_3336);
or U7136 (N_7136,N_3769,N_4671);
nor U7137 (N_7137,N_4955,N_3780);
nor U7138 (N_7138,N_3896,N_4138);
nor U7139 (N_7139,N_4143,N_4203);
and U7140 (N_7140,N_4671,N_3891);
and U7141 (N_7141,N_4778,N_2506);
xnor U7142 (N_7142,N_2935,N_4425);
xor U7143 (N_7143,N_3745,N_2877);
and U7144 (N_7144,N_2715,N_2745);
or U7145 (N_7145,N_2585,N_4627);
nand U7146 (N_7146,N_3055,N_3574);
or U7147 (N_7147,N_4938,N_3726);
or U7148 (N_7148,N_2694,N_4723);
or U7149 (N_7149,N_3636,N_4282);
and U7150 (N_7150,N_4265,N_3994);
nand U7151 (N_7151,N_3402,N_4920);
and U7152 (N_7152,N_4578,N_3068);
nor U7153 (N_7153,N_3322,N_3587);
nand U7154 (N_7154,N_4833,N_3472);
or U7155 (N_7155,N_4098,N_4951);
nand U7156 (N_7156,N_3037,N_3631);
nor U7157 (N_7157,N_4425,N_3200);
or U7158 (N_7158,N_3748,N_4856);
or U7159 (N_7159,N_4998,N_3413);
nand U7160 (N_7160,N_4277,N_3826);
or U7161 (N_7161,N_3782,N_4956);
nor U7162 (N_7162,N_4015,N_2694);
nand U7163 (N_7163,N_2872,N_2865);
nand U7164 (N_7164,N_4147,N_3512);
nor U7165 (N_7165,N_3936,N_4372);
or U7166 (N_7166,N_3281,N_4017);
and U7167 (N_7167,N_3482,N_2965);
xor U7168 (N_7168,N_3412,N_2893);
or U7169 (N_7169,N_4312,N_4881);
nand U7170 (N_7170,N_3193,N_4636);
or U7171 (N_7171,N_3545,N_3800);
and U7172 (N_7172,N_3436,N_2696);
nor U7173 (N_7173,N_2885,N_2568);
or U7174 (N_7174,N_3391,N_4233);
and U7175 (N_7175,N_2782,N_4994);
nor U7176 (N_7176,N_4983,N_4792);
nor U7177 (N_7177,N_3042,N_4936);
or U7178 (N_7178,N_4581,N_4330);
or U7179 (N_7179,N_4550,N_4130);
nor U7180 (N_7180,N_2954,N_4670);
nor U7181 (N_7181,N_3338,N_3734);
and U7182 (N_7182,N_3365,N_4022);
xnor U7183 (N_7183,N_4637,N_3648);
nand U7184 (N_7184,N_3765,N_2830);
nor U7185 (N_7185,N_3794,N_3556);
xor U7186 (N_7186,N_4310,N_4583);
nor U7187 (N_7187,N_4197,N_2701);
xnor U7188 (N_7188,N_3973,N_3225);
nand U7189 (N_7189,N_3942,N_2782);
nor U7190 (N_7190,N_2697,N_3395);
nand U7191 (N_7191,N_3821,N_3914);
nor U7192 (N_7192,N_2847,N_4180);
xnor U7193 (N_7193,N_2896,N_4739);
xor U7194 (N_7194,N_4205,N_4537);
nand U7195 (N_7195,N_3717,N_2657);
nand U7196 (N_7196,N_4745,N_3351);
xor U7197 (N_7197,N_2560,N_4417);
nand U7198 (N_7198,N_3063,N_2565);
xor U7199 (N_7199,N_4846,N_3768);
xnor U7200 (N_7200,N_3403,N_4634);
or U7201 (N_7201,N_2539,N_3040);
nand U7202 (N_7202,N_3900,N_2603);
and U7203 (N_7203,N_3997,N_2798);
nand U7204 (N_7204,N_2643,N_2612);
and U7205 (N_7205,N_2776,N_2749);
nand U7206 (N_7206,N_4555,N_4159);
and U7207 (N_7207,N_2653,N_4094);
and U7208 (N_7208,N_3861,N_4923);
or U7209 (N_7209,N_2964,N_3034);
nor U7210 (N_7210,N_3456,N_4899);
and U7211 (N_7211,N_4597,N_4941);
nand U7212 (N_7212,N_4878,N_4378);
xor U7213 (N_7213,N_4671,N_2914);
or U7214 (N_7214,N_3518,N_4516);
nor U7215 (N_7215,N_4672,N_3598);
or U7216 (N_7216,N_3992,N_3443);
or U7217 (N_7217,N_3997,N_3296);
nand U7218 (N_7218,N_4529,N_3834);
xor U7219 (N_7219,N_4226,N_3139);
xnor U7220 (N_7220,N_3227,N_3237);
nor U7221 (N_7221,N_2727,N_2822);
xor U7222 (N_7222,N_3746,N_3039);
and U7223 (N_7223,N_3334,N_3940);
nand U7224 (N_7224,N_4055,N_2778);
nand U7225 (N_7225,N_2697,N_4157);
and U7226 (N_7226,N_4093,N_4586);
nand U7227 (N_7227,N_3763,N_3929);
and U7228 (N_7228,N_3987,N_4710);
nand U7229 (N_7229,N_2924,N_4942);
or U7230 (N_7230,N_2598,N_3647);
xnor U7231 (N_7231,N_2966,N_4019);
or U7232 (N_7232,N_3333,N_4297);
or U7233 (N_7233,N_2601,N_3979);
or U7234 (N_7234,N_3648,N_4942);
xnor U7235 (N_7235,N_4816,N_3489);
nor U7236 (N_7236,N_4913,N_2905);
xnor U7237 (N_7237,N_2543,N_3780);
and U7238 (N_7238,N_4566,N_3067);
xor U7239 (N_7239,N_4029,N_2586);
nand U7240 (N_7240,N_3144,N_2953);
xor U7241 (N_7241,N_4768,N_3034);
nand U7242 (N_7242,N_4094,N_2955);
and U7243 (N_7243,N_4910,N_3796);
and U7244 (N_7244,N_3068,N_4713);
nand U7245 (N_7245,N_4696,N_4352);
nand U7246 (N_7246,N_4038,N_4608);
and U7247 (N_7247,N_3159,N_4118);
and U7248 (N_7248,N_4116,N_3721);
xor U7249 (N_7249,N_4537,N_4557);
xnor U7250 (N_7250,N_3235,N_4904);
and U7251 (N_7251,N_3799,N_2739);
xor U7252 (N_7252,N_3923,N_2685);
xor U7253 (N_7253,N_3357,N_3696);
nand U7254 (N_7254,N_3518,N_3397);
xor U7255 (N_7255,N_4336,N_4884);
xnor U7256 (N_7256,N_2915,N_4832);
nor U7257 (N_7257,N_3745,N_3100);
xnor U7258 (N_7258,N_2644,N_3809);
xnor U7259 (N_7259,N_3630,N_3891);
xor U7260 (N_7260,N_2984,N_3936);
nor U7261 (N_7261,N_3193,N_3708);
nand U7262 (N_7262,N_3813,N_2890);
nor U7263 (N_7263,N_2622,N_4257);
xor U7264 (N_7264,N_4481,N_2680);
nand U7265 (N_7265,N_4370,N_3259);
nor U7266 (N_7266,N_2817,N_3455);
nor U7267 (N_7267,N_4501,N_4748);
nand U7268 (N_7268,N_4295,N_4045);
nor U7269 (N_7269,N_3316,N_3918);
or U7270 (N_7270,N_3355,N_2682);
nand U7271 (N_7271,N_4824,N_3466);
nor U7272 (N_7272,N_2531,N_3756);
nor U7273 (N_7273,N_4613,N_4834);
nand U7274 (N_7274,N_4081,N_4623);
xnor U7275 (N_7275,N_3235,N_2995);
and U7276 (N_7276,N_4031,N_4568);
and U7277 (N_7277,N_3526,N_4935);
xnor U7278 (N_7278,N_4741,N_2546);
nor U7279 (N_7279,N_4245,N_3223);
or U7280 (N_7280,N_2606,N_2987);
nor U7281 (N_7281,N_2969,N_4414);
nand U7282 (N_7282,N_2669,N_3120);
nor U7283 (N_7283,N_4331,N_4206);
and U7284 (N_7284,N_4393,N_2790);
nand U7285 (N_7285,N_2943,N_4847);
nand U7286 (N_7286,N_3148,N_4470);
and U7287 (N_7287,N_4808,N_3477);
and U7288 (N_7288,N_2904,N_3420);
or U7289 (N_7289,N_4902,N_4321);
nor U7290 (N_7290,N_3672,N_2567);
nand U7291 (N_7291,N_2505,N_4604);
and U7292 (N_7292,N_3497,N_4982);
nor U7293 (N_7293,N_2819,N_4351);
xor U7294 (N_7294,N_3754,N_3260);
and U7295 (N_7295,N_3261,N_3419);
nor U7296 (N_7296,N_4262,N_4021);
or U7297 (N_7297,N_4051,N_3113);
xor U7298 (N_7298,N_2757,N_4199);
and U7299 (N_7299,N_4949,N_4033);
and U7300 (N_7300,N_3478,N_4334);
or U7301 (N_7301,N_3531,N_3950);
nor U7302 (N_7302,N_4372,N_3760);
and U7303 (N_7303,N_4953,N_2770);
or U7304 (N_7304,N_2586,N_4167);
or U7305 (N_7305,N_3069,N_4474);
and U7306 (N_7306,N_4824,N_3670);
or U7307 (N_7307,N_3996,N_3013);
or U7308 (N_7308,N_3684,N_3122);
or U7309 (N_7309,N_4948,N_3754);
nor U7310 (N_7310,N_4268,N_2690);
or U7311 (N_7311,N_4706,N_2517);
or U7312 (N_7312,N_4362,N_3952);
and U7313 (N_7313,N_3811,N_3404);
nand U7314 (N_7314,N_3310,N_4194);
and U7315 (N_7315,N_3018,N_4448);
nand U7316 (N_7316,N_3617,N_3676);
nor U7317 (N_7317,N_4468,N_3616);
and U7318 (N_7318,N_2750,N_4611);
nor U7319 (N_7319,N_4967,N_2626);
or U7320 (N_7320,N_3010,N_4636);
xor U7321 (N_7321,N_3092,N_3615);
and U7322 (N_7322,N_3485,N_3010);
or U7323 (N_7323,N_4752,N_4342);
or U7324 (N_7324,N_2916,N_4768);
xor U7325 (N_7325,N_2684,N_4341);
or U7326 (N_7326,N_2581,N_3629);
xnor U7327 (N_7327,N_4529,N_2512);
or U7328 (N_7328,N_3029,N_3870);
and U7329 (N_7329,N_3271,N_4932);
or U7330 (N_7330,N_4983,N_4911);
nand U7331 (N_7331,N_3121,N_4512);
xnor U7332 (N_7332,N_2696,N_4244);
xor U7333 (N_7333,N_3619,N_2954);
and U7334 (N_7334,N_4749,N_4537);
and U7335 (N_7335,N_3288,N_2992);
nand U7336 (N_7336,N_3035,N_4013);
or U7337 (N_7337,N_3885,N_2831);
or U7338 (N_7338,N_4471,N_2653);
xor U7339 (N_7339,N_3288,N_4218);
and U7340 (N_7340,N_3349,N_3656);
and U7341 (N_7341,N_4951,N_2617);
nor U7342 (N_7342,N_3357,N_4011);
nand U7343 (N_7343,N_2577,N_4628);
xnor U7344 (N_7344,N_4324,N_3465);
and U7345 (N_7345,N_3560,N_2932);
nand U7346 (N_7346,N_4015,N_3045);
or U7347 (N_7347,N_3210,N_2561);
xnor U7348 (N_7348,N_3455,N_3489);
and U7349 (N_7349,N_4211,N_3795);
or U7350 (N_7350,N_3432,N_3340);
nand U7351 (N_7351,N_4494,N_2730);
or U7352 (N_7352,N_2591,N_2895);
nand U7353 (N_7353,N_4041,N_3642);
nand U7354 (N_7354,N_3404,N_3699);
nor U7355 (N_7355,N_3154,N_3131);
nor U7356 (N_7356,N_2893,N_4469);
and U7357 (N_7357,N_4913,N_4932);
nor U7358 (N_7358,N_3913,N_3999);
nand U7359 (N_7359,N_3318,N_3052);
xor U7360 (N_7360,N_3711,N_3818);
or U7361 (N_7361,N_4599,N_4435);
and U7362 (N_7362,N_4436,N_4118);
nand U7363 (N_7363,N_3812,N_3523);
and U7364 (N_7364,N_4051,N_4226);
xnor U7365 (N_7365,N_4671,N_3131);
or U7366 (N_7366,N_2613,N_3115);
and U7367 (N_7367,N_3570,N_4060);
nor U7368 (N_7368,N_4837,N_4501);
or U7369 (N_7369,N_3885,N_3126);
and U7370 (N_7370,N_4579,N_3006);
xnor U7371 (N_7371,N_2736,N_3978);
and U7372 (N_7372,N_4475,N_3300);
nor U7373 (N_7373,N_3482,N_3456);
or U7374 (N_7374,N_3881,N_4559);
nor U7375 (N_7375,N_3396,N_2805);
xor U7376 (N_7376,N_2794,N_3410);
nor U7377 (N_7377,N_3181,N_3037);
or U7378 (N_7378,N_3667,N_3252);
xnor U7379 (N_7379,N_3061,N_4361);
nand U7380 (N_7380,N_4866,N_3601);
xnor U7381 (N_7381,N_2721,N_3664);
or U7382 (N_7382,N_4684,N_3613);
and U7383 (N_7383,N_3420,N_3400);
and U7384 (N_7384,N_3485,N_4763);
or U7385 (N_7385,N_2695,N_4546);
or U7386 (N_7386,N_4305,N_3251);
nand U7387 (N_7387,N_2915,N_4096);
and U7388 (N_7388,N_2777,N_2735);
and U7389 (N_7389,N_3998,N_3415);
and U7390 (N_7390,N_3786,N_3602);
nor U7391 (N_7391,N_3565,N_4817);
xor U7392 (N_7392,N_3165,N_2562);
nand U7393 (N_7393,N_4688,N_2885);
or U7394 (N_7394,N_3649,N_2859);
nand U7395 (N_7395,N_3447,N_2573);
nor U7396 (N_7396,N_3518,N_3140);
and U7397 (N_7397,N_3385,N_4207);
or U7398 (N_7398,N_2601,N_3307);
xnor U7399 (N_7399,N_4854,N_2844);
nand U7400 (N_7400,N_2619,N_3087);
xnor U7401 (N_7401,N_3173,N_2766);
and U7402 (N_7402,N_3251,N_4073);
or U7403 (N_7403,N_3604,N_4879);
and U7404 (N_7404,N_4765,N_3561);
nand U7405 (N_7405,N_3403,N_2954);
nand U7406 (N_7406,N_3596,N_3555);
and U7407 (N_7407,N_4126,N_2829);
nor U7408 (N_7408,N_2758,N_2642);
or U7409 (N_7409,N_3956,N_4296);
xor U7410 (N_7410,N_2725,N_4659);
nand U7411 (N_7411,N_4595,N_4393);
and U7412 (N_7412,N_4509,N_2684);
or U7413 (N_7413,N_3612,N_2950);
and U7414 (N_7414,N_4042,N_3793);
nand U7415 (N_7415,N_3479,N_3059);
nand U7416 (N_7416,N_2817,N_4655);
nor U7417 (N_7417,N_4532,N_4273);
nor U7418 (N_7418,N_3148,N_3133);
nor U7419 (N_7419,N_4337,N_2989);
nor U7420 (N_7420,N_2503,N_4468);
xnor U7421 (N_7421,N_2775,N_4764);
nand U7422 (N_7422,N_3683,N_2631);
nor U7423 (N_7423,N_3203,N_3761);
nand U7424 (N_7424,N_4751,N_3218);
and U7425 (N_7425,N_2860,N_4720);
nor U7426 (N_7426,N_2577,N_4528);
and U7427 (N_7427,N_3570,N_4178);
nand U7428 (N_7428,N_4849,N_3190);
nand U7429 (N_7429,N_4325,N_4278);
nor U7430 (N_7430,N_4506,N_2579);
and U7431 (N_7431,N_3011,N_4194);
or U7432 (N_7432,N_4278,N_3113);
nor U7433 (N_7433,N_4156,N_3755);
nor U7434 (N_7434,N_2800,N_3516);
nor U7435 (N_7435,N_4369,N_3580);
nand U7436 (N_7436,N_4832,N_4464);
nor U7437 (N_7437,N_2870,N_2897);
nor U7438 (N_7438,N_3352,N_2670);
xnor U7439 (N_7439,N_4230,N_4166);
or U7440 (N_7440,N_4236,N_3425);
nor U7441 (N_7441,N_3376,N_3818);
xor U7442 (N_7442,N_2983,N_3660);
or U7443 (N_7443,N_3730,N_4079);
and U7444 (N_7444,N_2822,N_3153);
xnor U7445 (N_7445,N_4725,N_4150);
or U7446 (N_7446,N_3742,N_3253);
nand U7447 (N_7447,N_3434,N_3079);
or U7448 (N_7448,N_4022,N_3812);
xnor U7449 (N_7449,N_3152,N_2870);
and U7450 (N_7450,N_4808,N_3964);
or U7451 (N_7451,N_4908,N_4152);
nor U7452 (N_7452,N_2824,N_3747);
and U7453 (N_7453,N_4208,N_4662);
nor U7454 (N_7454,N_3979,N_3063);
nor U7455 (N_7455,N_3774,N_4702);
and U7456 (N_7456,N_2601,N_3343);
xnor U7457 (N_7457,N_4461,N_3915);
nand U7458 (N_7458,N_3374,N_3653);
or U7459 (N_7459,N_3019,N_3949);
xor U7460 (N_7460,N_3643,N_2535);
nand U7461 (N_7461,N_4424,N_3534);
nor U7462 (N_7462,N_2501,N_4196);
xor U7463 (N_7463,N_2786,N_3311);
or U7464 (N_7464,N_3419,N_4840);
nand U7465 (N_7465,N_3004,N_4562);
or U7466 (N_7466,N_4231,N_4467);
xnor U7467 (N_7467,N_4672,N_4372);
or U7468 (N_7468,N_2654,N_4175);
nand U7469 (N_7469,N_2657,N_4964);
and U7470 (N_7470,N_4402,N_4549);
nor U7471 (N_7471,N_3155,N_3034);
nor U7472 (N_7472,N_2777,N_3599);
or U7473 (N_7473,N_3577,N_3149);
nor U7474 (N_7474,N_3815,N_3950);
nor U7475 (N_7475,N_4176,N_4719);
or U7476 (N_7476,N_3751,N_3133);
nand U7477 (N_7477,N_3829,N_2977);
and U7478 (N_7478,N_4168,N_3066);
xnor U7479 (N_7479,N_3890,N_3224);
xor U7480 (N_7480,N_3040,N_4907);
and U7481 (N_7481,N_4508,N_2520);
or U7482 (N_7482,N_3591,N_4166);
or U7483 (N_7483,N_3601,N_4963);
or U7484 (N_7484,N_3836,N_4789);
nand U7485 (N_7485,N_3716,N_4399);
xnor U7486 (N_7486,N_2928,N_2919);
nor U7487 (N_7487,N_3806,N_3694);
or U7488 (N_7488,N_4113,N_2764);
or U7489 (N_7489,N_3725,N_3855);
xor U7490 (N_7490,N_4932,N_3635);
nor U7491 (N_7491,N_4700,N_3176);
nand U7492 (N_7492,N_4531,N_3577);
or U7493 (N_7493,N_3422,N_3043);
or U7494 (N_7494,N_2517,N_3965);
xnor U7495 (N_7495,N_3393,N_2793);
nand U7496 (N_7496,N_3050,N_3410);
and U7497 (N_7497,N_2865,N_3787);
nor U7498 (N_7498,N_4925,N_4684);
xnor U7499 (N_7499,N_4690,N_4845);
nor U7500 (N_7500,N_6397,N_5060);
nand U7501 (N_7501,N_7192,N_5538);
nand U7502 (N_7502,N_5420,N_7045);
xnor U7503 (N_7503,N_7022,N_7158);
nand U7504 (N_7504,N_6983,N_6526);
and U7505 (N_7505,N_6509,N_7016);
nor U7506 (N_7506,N_6995,N_6233);
and U7507 (N_7507,N_5808,N_6144);
nand U7508 (N_7508,N_5260,N_5314);
nand U7509 (N_7509,N_6176,N_5346);
nand U7510 (N_7510,N_5331,N_5436);
or U7511 (N_7511,N_6858,N_6743);
and U7512 (N_7512,N_6820,N_5287);
nor U7513 (N_7513,N_6523,N_5716);
nand U7514 (N_7514,N_6985,N_7348);
and U7515 (N_7515,N_6211,N_6740);
nand U7516 (N_7516,N_5533,N_5893);
xnor U7517 (N_7517,N_6221,N_5304);
nand U7518 (N_7518,N_5862,N_6500);
nor U7519 (N_7519,N_5102,N_6992);
nand U7520 (N_7520,N_5568,N_5558);
nor U7521 (N_7521,N_6970,N_6531);
nor U7522 (N_7522,N_6905,N_5253);
and U7523 (N_7523,N_7445,N_6727);
and U7524 (N_7524,N_6598,N_5736);
nor U7525 (N_7525,N_7068,N_7433);
and U7526 (N_7526,N_7204,N_6096);
or U7527 (N_7527,N_7388,N_6404);
xor U7528 (N_7528,N_7049,N_6173);
and U7529 (N_7529,N_7131,N_6051);
and U7530 (N_7530,N_7205,N_5670);
nor U7531 (N_7531,N_5642,N_6689);
or U7532 (N_7532,N_6501,N_6507);
nand U7533 (N_7533,N_7404,N_5581);
nor U7534 (N_7534,N_7362,N_6936);
nor U7535 (N_7535,N_6043,N_6186);
or U7536 (N_7536,N_6941,N_5431);
nand U7537 (N_7537,N_5372,N_6587);
and U7538 (N_7538,N_5326,N_5173);
xor U7539 (N_7539,N_7415,N_6961);
or U7540 (N_7540,N_6105,N_6672);
or U7541 (N_7541,N_6636,N_5148);
xnor U7542 (N_7542,N_5891,N_7059);
and U7543 (N_7543,N_7402,N_6384);
xnor U7544 (N_7544,N_7499,N_5942);
nand U7545 (N_7545,N_7419,N_5035);
nand U7546 (N_7546,N_5203,N_6484);
and U7547 (N_7547,N_6889,N_5181);
nand U7548 (N_7548,N_5274,N_5805);
nor U7549 (N_7549,N_7467,N_7179);
and U7550 (N_7550,N_6447,N_5583);
nand U7551 (N_7551,N_5972,N_5960);
and U7552 (N_7552,N_7409,N_5498);
and U7553 (N_7553,N_6352,N_6213);
nand U7554 (N_7554,N_7309,N_5098);
or U7555 (N_7555,N_7458,N_5775);
or U7556 (N_7556,N_5537,N_6423);
nor U7557 (N_7557,N_5495,N_7232);
nand U7558 (N_7558,N_6470,N_5273);
nand U7559 (N_7559,N_6571,N_5439);
nor U7560 (N_7560,N_6456,N_5769);
nand U7561 (N_7561,N_5396,N_5467);
or U7562 (N_7562,N_5881,N_6100);
nor U7563 (N_7563,N_6007,N_6294);
nand U7564 (N_7564,N_7490,N_5167);
and U7565 (N_7565,N_5072,N_5363);
or U7566 (N_7566,N_7306,N_6282);
or U7567 (N_7567,N_5096,N_5466);
xor U7568 (N_7568,N_7399,N_6714);
and U7569 (N_7569,N_6957,N_5381);
or U7570 (N_7570,N_7082,N_5874);
xor U7571 (N_7571,N_5593,N_6111);
nand U7572 (N_7572,N_5021,N_5226);
nor U7573 (N_7573,N_7073,N_6094);
nand U7574 (N_7574,N_7237,N_5359);
nor U7575 (N_7575,N_5350,N_6769);
or U7576 (N_7576,N_6167,N_7225);
xnor U7577 (N_7577,N_5027,N_6859);
or U7578 (N_7578,N_5851,N_7254);
and U7579 (N_7579,N_7097,N_5632);
and U7580 (N_7580,N_6867,N_7035);
or U7581 (N_7581,N_6402,N_6067);
nand U7582 (N_7582,N_5379,N_5044);
nand U7583 (N_7583,N_6522,N_6826);
nor U7584 (N_7584,N_5634,N_6409);
nor U7585 (N_7585,N_6411,N_5463);
or U7586 (N_7586,N_5761,N_5286);
xnor U7587 (N_7587,N_6314,N_5054);
or U7588 (N_7588,N_7487,N_6909);
nand U7589 (N_7589,N_6506,N_5432);
and U7590 (N_7590,N_7211,N_7265);
and U7591 (N_7591,N_6641,N_6090);
xor U7592 (N_7592,N_6271,N_5600);
nand U7593 (N_7593,N_7349,N_5156);
nor U7594 (N_7594,N_5756,N_7485);
nand U7595 (N_7595,N_5180,N_5402);
nor U7596 (N_7596,N_5577,N_6442);
xnor U7597 (N_7597,N_6912,N_6882);
xnor U7598 (N_7598,N_6006,N_6567);
or U7599 (N_7599,N_6839,N_5742);
xnor U7600 (N_7600,N_7005,N_6750);
nor U7601 (N_7601,N_6316,N_6538);
xor U7602 (N_7602,N_6134,N_5366);
or U7603 (N_7603,N_6710,N_5841);
and U7604 (N_7604,N_5987,N_7367);
nor U7605 (N_7605,N_6130,N_5015);
and U7606 (N_7606,N_5609,N_6265);
nor U7607 (N_7607,N_6473,N_6788);
nand U7608 (N_7608,N_5418,N_7471);
nor U7609 (N_7609,N_6234,N_6573);
or U7610 (N_7610,N_6685,N_5394);
or U7611 (N_7611,N_6795,N_6181);
or U7612 (N_7612,N_6440,N_7406);
and U7613 (N_7613,N_7029,N_5790);
nand U7614 (N_7614,N_6003,N_6064);
or U7615 (N_7615,N_5678,N_5292);
nand U7616 (N_7616,N_6024,N_6058);
nor U7617 (N_7617,N_7238,N_6330);
or U7618 (N_7618,N_7377,N_5417);
and U7619 (N_7619,N_6155,N_5248);
xnor U7620 (N_7620,N_6548,N_6841);
nor U7621 (N_7621,N_5702,N_5852);
nor U7622 (N_7622,N_5190,N_6783);
and U7623 (N_7623,N_5585,N_7425);
xor U7624 (N_7624,N_5267,N_7241);
xnor U7625 (N_7625,N_6231,N_5689);
xor U7626 (N_7626,N_5848,N_7346);
or U7627 (N_7627,N_5205,N_7378);
and U7628 (N_7628,N_6774,N_6717);
nand U7629 (N_7629,N_5089,N_6785);
nor U7630 (N_7630,N_7261,N_6610);
nor U7631 (N_7631,N_5010,N_5921);
or U7632 (N_7632,N_5612,N_6516);
xnor U7633 (N_7633,N_5835,N_5022);
nand U7634 (N_7634,N_6150,N_5626);
nor U7635 (N_7635,N_7311,N_6421);
nand U7636 (N_7636,N_5816,N_6331);
and U7637 (N_7637,N_6419,N_5724);
or U7638 (N_7638,N_7114,N_5928);
nand U7639 (N_7639,N_5557,N_6428);
xnor U7640 (N_7640,N_7465,N_5582);
xor U7641 (N_7641,N_7001,N_6766);
or U7642 (N_7642,N_6949,N_7442);
xnor U7643 (N_7643,N_7017,N_6457);
nand U7644 (N_7644,N_7012,N_7075);
nand U7645 (N_7645,N_5038,N_5815);
and U7646 (N_7646,N_6990,N_5832);
nand U7647 (N_7647,N_6629,N_6278);
xnor U7648 (N_7648,N_6832,N_6799);
xor U7649 (N_7649,N_6373,N_5509);
nand U7650 (N_7650,N_5799,N_5513);
nand U7651 (N_7651,N_5449,N_5116);
nor U7652 (N_7652,N_7109,N_5643);
or U7653 (N_7653,N_6677,N_7120);
nand U7654 (N_7654,N_5317,N_5677);
or U7655 (N_7655,N_6805,N_7486);
nand U7656 (N_7656,N_5638,N_7496);
and U7657 (N_7657,N_5934,N_7356);
nor U7658 (N_7658,N_6078,N_7421);
nand U7659 (N_7659,N_5000,N_5947);
xor U7660 (N_7660,N_7278,N_6748);
nand U7661 (N_7661,N_5348,N_6301);
or U7662 (N_7662,N_6656,N_5965);
nor U7663 (N_7663,N_5143,N_5514);
or U7664 (N_7664,N_6227,N_6471);
nand U7665 (N_7665,N_7340,N_7498);
or U7666 (N_7666,N_5567,N_6008);
or U7667 (N_7667,N_5185,N_7376);
or U7668 (N_7668,N_7429,N_6873);
and U7669 (N_7669,N_6874,N_6813);
xor U7670 (N_7670,N_5145,N_5031);
nand U7671 (N_7671,N_6654,N_5327);
and U7672 (N_7672,N_5049,N_6308);
nor U7673 (N_7673,N_5081,N_6888);
xnor U7674 (N_7674,N_5788,N_5763);
and U7675 (N_7675,N_7247,N_6753);
nand U7676 (N_7676,N_5813,N_5201);
or U7677 (N_7677,N_5058,N_5887);
nor U7678 (N_7678,N_6232,N_7180);
nor U7679 (N_7679,N_6408,N_6482);
xnor U7680 (N_7680,N_5825,N_7361);
xor U7681 (N_7681,N_6448,N_5408);
xnor U7682 (N_7682,N_7121,N_5620);
or U7683 (N_7683,N_6153,N_7440);
and U7684 (N_7684,N_6978,N_6063);
nand U7685 (N_7685,N_5728,N_6102);
xor U7686 (N_7686,N_6074,N_6767);
nand U7687 (N_7687,N_5554,N_7470);
or U7688 (N_7688,N_7066,N_5545);
nor U7689 (N_7689,N_5768,N_5002);
and U7690 (N_7690,N_5536,N_6387);
xnor U7691 (N_7691,N_7056,N_6950);
and U7692 (N_7692,N_5275,N_6206);
nor U7693 (N_7693,N_6376,N_5871);
and U7694 (N_7694,N_6853,N_5047);
and U7695 (N_7695,N_5905,N_7010);
or U7696 (N_7696,N_7221,N_7391);
or U7697 (N_7697,N_5624,N_5265);
xnor U7698 (N_7698,N_5152,N_5877);
or U7699 (N_7699,N_7432,N_6147);
nand U7700 (N_7700,N_5555,N_5489);
xnor U7701 (N_7701,N_5320,N_5142);
nand U7702 (N_7702,N_5004,N_7149);
nand U7703 (N_7703,N_5720,N_5909);
and U7704 (N_7704,N_7087,N_7187);
or U7705 (N_7705,N_5045,N_6488);
nand U7706 (N_7706,N_6198,N_5935);
and U7707 (N_7707,N_6298,N_6116);
nand U7708 (N_7708,N_6542,N_7342);
xor U7709 (N_7709,N_7101,N_7305);
nand U7710 (N_7710,N_5783,N_6350);
nor U7711 (N_7711,N_6701,N_5884);
or U7712 (N_7712,N_5120,N_7090);
and U7713 (N_7713,N_5859,N_5809);
nor U7714 (N_7714,N_6117,N_5012);
and U7715 (N_7715,N_6259,N_5584);
or U7716 (N_7716,N_6603,N_6129);
nand U7717 (N_7717,N_5365,N_7230);
nand U7718 (N_7718,N_5801,N_6885);
and U7719 (N_7719,N_5594,N_5588);
xor U7720 (N_7720,N_7023,N_6989);
nor U7721 (N_7721,N_5491,N_7351);
nor U7722 (N_7722,N_6170,N_7042);
nor U7723 (N_7723,N_6215,N_6586);
and U7724 (N_7724,N_6268,N_5174);
and U7725 (N_7725,N_6709,N_5906);
and U7726 (N_7726,N_5944,N_5510);
or U7727 (N_7727,N_5607,N_5525);
xor U7728 (N_7728,N_5202,N_6216);
xnor U7729 (N_7729,N_6568,N_5666);
nand U7730 (N_7730,N_6830,N_5188);
and U7731 (N_7731,N_6029,N_6354);
or U7732 (N_7732,N_7046,N_5213);
nor U7733 (N_7733,N_6570,N_6017);
nor U7734 (N_7734,N_6158,N_5693);
or U7735 (N_7735,N_7366,N_6092);
and U7736 (N_7736,N_6791,N_5990);
xor U7737 (N_7737,N_5065,N_7151);
nor U7738 (N_7738,N_5302,N_7206);
and U7739 (N_7739,N_6236,N_5209);
xnor U7740 (N_7740,N_5014,N_5323);
xor U7741 (N_7741,N_7085,N_5685);
nand U7742 (N_7742,N_5461,N_6430);
nor U7743 (N_7743,N_7480,N_6264);
and U7744 (N_7744,N_6773,N_5738);
and U7745 (N_7745,N_5705,N_5611);
nor U7746 (N_7746,N_5914,N_7063);
or U7747 (N_7747,N_7285,N_6020);
nor U7748 (N_7748,N_5687,N_6368);
xnor U7749 (N_7749,N_7497,N_5223);
xnor U7750 (N_7750,N_5662,N_6427);
xnor U7751 (N_7751,N_5127,N_7092);
nor U7752 (N_7752,N_6337,N_5500);
or U7753 (N_7753,N_7474,N_6136);
and U7754 (N_7754,N_6599,N_6792);
and U7755 (N_7755,N_6393,N_5691);
and U7756 (N_7756,N_6422,N_7268);
nand U7757 (N_7757,N_5159,N_6938);
or U7758 (N_7758,N_5412,N_6347);
nor U7759 (N_7759,N_5970,N_7038);
or U7760 (N_7760,N_5817,N_6031);
nor U7761 (N_7761,N_6461,N_5648);
nor U7762 (N_7762,N_6048,N_6871);
xor U7763 (N_7763,N_7400,N_5373);
xnor U7764 (N_7764,N_5658,N_7369);
and U7765 (N_7765,N_5268,N_6417);
nand U7766 (N_7766,N_5541,N_6632);
nand U7767 (N_7767,N_5628,N_5748);
nor U7768 (N_7768,N_6786,N_7129);
xnor U7769 (N_7769,N_5590,N_7008);
and U7770 (N_7770,N_7084,N_6046);
xnor U7771 (N_7771,N_6551,N_6850);
or U7772 (N_7772,N_7272,N_5665);
and U7773 (N_7773,N_5196,N_6662);
nor U7774 (N_7774,N_5560,N_6412);
nand U7775 (N_7775,N_5401,N_6203);
nor U7776 (N_7776,N_5547,N_5855);
and U7777 (N_7777,N_5993,N_6565);
and U7778 (N_7778,N_6707,N_7181);
or U7779 (N_7779,N_5637,N_7252);
and U7780 (N_7780,N_6154,N_6295);
nand U7781 (N_7781,N_6975,N_6825);
nor U7782 (N_7782,N_6606,N_6686);
xor U7783 (N_7783,N_6544,N_5948);
xnor U7784 (N_7784,N_7488,N_6394);
nor U7785 (N_7785,N_7083,N_6763);
nand U7786 (N_7786,N_5645,N_5596);
xnor U7787 (N_7787,N_7080,N_5087);
and U7788 (N_7788,N_5849,N_6039);
nand U7789 (N_7789,N_6287,N_5169);
nand U7790 (N_7790,N_7191,N_6687);
xor U7791 (N_7791,N_7019,N_7395);
and U7792 (N_7792,N_5493,N_5225);
and U7793 (N_7793,N_7096,N_5200);
or U7794 (N_7794,N_5357,N_5591);
nor U7795 (N_7795,N_7267,N_7164);
and U7796 (N_7796,N_7276,N_5023);
or U7797 (N_7797,N_7177,N_6120);
and U7798 (N_7798,N_6680,N_5272);
nand U7799 (N_7799,N_6856,N_6252);
nand U7800 (N_7800,N_6380,N_6951);
xor U7801 (N_7801,N_5969,N_5669);
xnor U7802 (N_7802,N_6340,N_6730);
nor U7803 (N_7803,N_6256,N_6140);
xor U7804 (N_7804,N_5534,N_6351);
xor U7805 (N_7805,N_6266,N_5958);
nor U7806 (N_7806,N_6061,N_5562);
or U7807 (N_7807,N_5428,N_5258);
xor U7808 (N_7808,N_7363,N_6138);
xor U7809 (N_7809,N_7058,N_7152);
and U7810 (N_7810,N_5496,N_5499);
or U7811 (N_7811,N_6405,N_5369);
nand U7812 (N_7812,N_6212,N_6922);
xnor U7813 (N_7813,N_6794,N_5410);
nor U7814 (N_7814,N_5345,N_7455);
nor U7815 (N_7815,N_6353,N_7359);
xnor U7816 (N_7816,N_5903,N_5812);
nor U7817 (N_7817,N_7236,N_6016);
nor U7818 (N_7818,N_5179,N_5654);
and U7819 (N_7819,N_6625,N_5117);
nand U7820 (N_7820,N_7446,N_5351);
nor U7821 (N_7821,N_5422,N_5885);
nor U7822 (N_7822,N_6127,N_6612);
and U7823 (N_7823,N_6205,N_7479);
xnor U7824 (N_7824,N_5187,N_6512);
or U7825 (N_7825,N_6831,N_6238);
nand U7826 (N_7826,N_5967,N_6851);
nand U7827 (N_7827,N_6514,N_7318);
and U7828 (N_7828,N_5219,N_6431);
xor U7829 (N_7829,N_5975,N_6172);
nand U7830 (N_7830,N_5092,N_6892);
nand U7831 (N_7831,N_5186,N_7112);
xnor U7832 (N_7832,N_6944,N_6809);
or U7833 (N_7833,N_6403,N_5503);
or U7834 (N_7834,N_7463,N_6436);
xor U7835 (N_7835,N_7245,N_7472);
or U7836 (N_7836,N_6469,N_7341);
and U7837 (N_7837,N_5842,N_7466);
nand U7838 (N_7838,N_6503,N_6817);
nor U7839 (N_7839,N_6962,N_7482);
nand U7840 (N_7840,N_6081,N_7320);
nor U7841 (N_7841,N_6280,N_5563);
or U7842 (N_7842,N_6637,N_6998);
nand U7843 (N_7843,N_6269,N_5551);
or U7844 (N_7844,N_6835,N_6620);
and U7845 (N_7845,N_5542,N_5414);
nor U7846 (N_7846,N_5456,N_6114);
and U7847 (N_7847,N_6056,N_6908);
or U7848 (N_7848,N_6700,N_7155);
nand U7849 (N_7849,N_5690,N_6493);
nor U7850 (N_7850,N_6684,N_6323);
or U7851 (N_7851,N_7034,N_6933);
or U7852 (N_7852,N_5328,N_5476);
and U7853 (N_7853,N_5462,N_6787);
xnor U7854 (N_7854,N_5210,N_5195);
nor U7855 (N_7855,N_6375,N_5744);
or U7856 (N_7856,N_6665,N_7338);
and U7857 (N_7857,N_6622,N_5473);
and U7858 (N_7858,N_6285,N_7330);
nor U7859 (N_7859,N_5103,N_6183);
nor U7860 (N_7860,N_6192,N_5078);
or U7861 (N_7861,N_6217,N_7171);
nor U7862 (N_7862,N_5766,N_6987);
and U7863 (N_7863,N_5919,N_5356);
nand U7864 (N_7864,N_7064,N_6306);
nor U7865 (N_7865,N_5386,N_6000);
nor U7866 (N_7866,N_5233,N_5378);
and U7867 (N_7867,N_7235,N_7434);
nand U7868 (N_7868,N_5878,N_6521);
nand U7869 (N_7869,N_5288,N_6322);
and U7870 (N_7870,N_5251,N_6244);
nor U7871 (N_7871,N_6465,N_6847);
and U7872 (N_7872,N_5549,N_6073);
nor U7873 (N_7873,N_5130,N_6840);
and U7874 (N_7874,N_7405,N_6591);
or U7875 (N_7875,N_6091,N_5786);
or U7876 (N_7876,N_5646,N_6624);
xnor U7877 (N_7877,N_6108,N_5989);
xnor U7878 (N_7878,N_5943,N_5158);
xnor U7879 (N_7879,N_5968,N_7100);
and U7880 (N_7880,N_6865,N_6010);
nand U7881 (N_7881,N_5425,N_7300);
and U7882 (N_7882,N_5007,N_5112);
nand U7883 (N_7883,N_5349,N_5633);
or U7884 (N_7884,N_6284,N_6648);
or U7885 (N_7885,N_6060,N_6197);
xor U7886 (N_7886,N_5604,N_5811);
xor U7887 (N_7887,N_5316,N_6101);
and U7888 (N_7888,N_5168,N_6634);
nor U7889 (N_7889,N_7397,N_7195);
and U7890 (N_7890,N_5450,N_5552);
nor U7891 (N_7891,N_6142,N_7033);
nand U7892 (N_7892,N_7229,N_5505);
nand U7893 (N_7893,N_5937,N_5141);
nand U7894 (N_7894,N_7260,N_6343);
nand U7895 (N_7895,N_6566,N_6386);
xor U7896 (N_7896,N_7407,N_6906);
and U7897 (N_7897,N_7069,N_6149);
and U7898 (N_7898,N_5785,N_5310);
nand U7899 (N_7899,N_5754,N_5053);
and U7900 (N_7900,N_5732,N_5193);
xor U7901 (N_7901,N_7215,N_7098);
xor U7902 (N_7902,N_5189,N_5063);
and U7903 (N_7903,N_5207,N_6187);
nand U7904 (N_7904,N_5895,N_6804);
nor U7905 (N_7905,N_6711,N_5312);
or U7906 (N_7906,N_7089,N_5544);
xnor U7907 (N_7907,N_6939,N_6896);
xnor U7908 (N_7908,N_7134,N_5973);
nand U7909 (N_7909,N_7197,N_6728);
nor U7910 (N_7910,N_5247,N_6208);
and U7911 (N_7911,N_7250,N_5206);
and U7912 (N_7912,N_5270,N_5283);
and U7913 (N_7913,N_5644,N_6458);
or U7914 (N_7914,N_5427,N_5636);
and U7915 (N_7915,N_6462,N_6239);
or U7916 (N_7916,N_5299,N_5955);
nor U7917 (N_7917,N_5753,N_6658);
nor U7918 (N_7918,N_7344,N_6037);
or U7919 (N_7919,N_6608,N_7140);
nand U7920 (N_7920,N_5362,N_5030);
nor U7921 (N_7921,N_5639,N_6345);
and U7922 (N_7922,N_7459,N_7174);
or U7923 (N_7923,N_6455,N_5839);
or U7924 (N_7924,N_6319,N_5795);
nand U7925 (N_7925,N_5561,N_5668);
nand U7926 (N_7926,N_5172,N_6929);
nor U7927 (N_7927,N_6959,N_5191);
nor U7928 (N_7928,N_7118,N_6823);
nor U7929 (N_7929,N_5863,N_6644);
nand U7930 (N_7930,N_7313,N_6451);
or U7931 (N_7931,N_7283,N_5713);
and U7932 (N_7932,N_6971,N_6141);
or U7933 (N_7933,N_6574,N_5684);
or U7934 (N_7934,N_5986,N_5385);
nand U7935 (N_7935,N_5398,N_7025);
xor U7936 (N_7936,N_5249,N_7240);
xor U7937 (N_7937,N_6724,N_6655);
and U7938 (N_7938,N_5162,N_7288);
xnor U7939 (N_7939,N_6555,N_6148);
xor U7940 (N_7940,N_6434,N_5228);
or U7941 (N_7941,N_7036,N_6705);
nand U7942 (N_7942,N_6494,N_6619);
nand U7943 (N_7943,N_5576,N_5526);
and U7944 (N_7944,N_6775,N_5831);
and U7945 (N_7945,N_7186,N_5731);
nand U7946 (N_7946,N_5250,N_5999);
or U7947 (N_7947,N_5413,N_6812);
or U7948 (N_7948,N_6779,N_6675);
xnor U7949 (N_7949,N_6103,N_5478);
xor U7950 (N_7950,N_5411,N_7219);
or U7951 (N_7951,N_6535,N_6815);
or U7952 (N_7952,N_6475,N_6012);
or U7953 (N_7953,N_5111,N_7441);
or U7954 (N_7954,N_5959,N_5388);
xor U7955 (N_7955,N_7491,N_5559);
and U7956 (N_7956,N_6673,N_5681);
xnor U7957 (N_7957,N_5798,N_7161);
nor U7958 (N_7958,N_5184,N_5480);
nand U7959 (N_7959,N_5335,N_5695);
or U7960 (N_7960,N_7389,N_5377);
and U7961 (N_7961,N_7212,N_5471);
nor U7962 (N_7962,N_5957,N_6223);
xor U7963 (N_7963,N_6070,N_6161);
nor U7964 (N_7964,N_6879,N_7394);
or U7965 (N_7965,N_7325,N_7256);
xnor U7966 (N_7966,N_5289,N_5857);
and U7967 (N_7967,N_5627,N_6583);
xor U7968 (N_7968,N_6781,N_7427);
and U7969 (N_7969,N_6338,N_5619);
xor U7970 (N_7970,N_7207,N_6967);
nand U7971 (N_7971,N_5915,N_5936);
nand U7972 (N_7972,N_7358,N_6115);
and U7973 (N_7973,N_5086,N_5522);
or U7974 (N_7974,N_5869,N_6072);
nor U7975 (N_7975,N_6034,N_6713);
nand U7976 (N_7976,N_5897,N_5861);
or U7977 (N_7977,N_6023,N_5100);
nand U7978 (N_7978,N_5796,N_7263);
or U7979 (N_7979,N_6224,N_5828);
and U7980 (N_7980,N_5197,N_7431);
xor U7981 (N_7981,N_7021,N_6050);
nand U7982 (N_7982,N_7284,N_6777);
nand U7983 (N_7983,N_6923,N_6075);
and U7984 (N_7984,N_5548,N_6811);
nor U7985 (N_7985,N_5946,N_5523);
nor U7986 (N_7986,N_5565,N_5950);
nor U7987 (N_7987,N_5904,N_7384);
or U7988 (N_7988,N_5041,N_7122);
nand U7989 (N_7989,N_5652,N_7099);
nor U7990 (N_7990,N_5571,N_5170);
and U7991 (N_7991,N_6367,N_6911);
or U7992 (N_7992,N_7170,N_6175);
and U7993 (N_7993,N_6013,N_6429);
or U7994 (N_7994,N_6630,N_6616);
nor U7995 (N_7995,N_5256,N_5711);
or U7996 (N_7996,N_6868,N_6011);
or U7997 (N_7997,N_5484,N_6309);
nand U7998 (N_7998,N_6676,N_5515);
or U7999 (N_7999,N_7218,N_5793);
xnor U8000 (N_8000,N_5630,N_6560);
and U8001 (N_8001,N_6089,N_7253);
or U8002 (N_8002,N_6052,N_5052);
nor U8003 (N_8003,N_5866,N_5726);
or U8004 (N_8004,N_6229,N_6988);
xor U8005 (N_8005,N_5234,N_6479);
xnor U8006 (N_8006,N_7071,N_7373);
or U8007 (N_8007,N_6520,N_7018);
nor U8008 (N_8008,N_5888,N_7214);
and U8009 (N_8009,N_5527,N_5282);
xnor U8010 (N_8010,N_7128,N_5375);
nand U8011 (N_8011,N_5854,N_7242);
and U8012 (N_8012,N_6557,N_6047);
or U8013 (N_8013,N_5971,N_5067);
nand U8014 (N_8014,N_5380,N_6444);
or U8015 (N_8015,N_6366,N_5700);
xnor U8016 (N_8016,N_6055,N_5126);
nand U8017 (N_8017,N_6445,N_7452);
nand U8018 (N_8018,N_5784,N_5867);
or U8019 (N_8019,N_6916,N_5319);
nand U8020 (N_8020,N_6706,N_6897);
or U8021 (N_8021,N_7271,N_5198);
and U8022 (N_8022,N_6891,N_6018);
nand U8023 (N_8023,N_5823,N_5020);
and U8024 (N_8024,N_6098,N_6927);
nor U8025 (N_8025,N_6947,N_5929);
and U8026 (N_8026,N_5026,N_6401);
or U8027 (N_8027,N_7347,N_7013);
and U8028 (N_8028,N_5284,N_6802);
nand U8029 (N_8029,N_5334,N_6281);
nor U8030 (N_8030,N_6385,N_5718);
xor U8031 (N_8031,N_5907,N_7110);
and U8032 (N_8032,N_6901,N_6741);
nor U8033 (N_8033,N_6226,N_5782);
xnor U8034 (N_8034,N_5599,N_6716);
and U8035 (N_8035,N_5227,N_6803);
and U8036 (N_8036,N_6688,N_6245);
xnor U8037 (N_8037,N_5384,N_7148);
or U8038 (N_8038,N_5865,N_7493);
xor U8039 (N_8039,N_6601,N_6695);
or U8040 (N_8040,N_6605,N_5827);
xor U8041 (N_8041,N_5569,N_5192);
or U8042 (N_8042,N_6210,N_5107);
nor U8043 (N_8043,N_5019,N_6778);
nor U8044 (N_8044,N_6860,N_5743);
xnor U8045 (N_8045,N_7026,N_7386);
nor U8046 (N_8046,N_6814,N_5424);
or U8047 (N_8047,N_5028,N_5059);
nor U8048 (N_8048,N_6040,N_6782);
nand U8049 (N_8049,N_7116,N_5452);
nor U8050 (N_8050,N_6588,N_6201);
nand U8051 (N_8051,N_6476,N_6320);
xnor U8052 (N_8052,N_6135,N_7299);
nor U8053 (N_8053,N_5951,N_6534);
or U8054 (N_8054,N_6973,N_7166);
nor U8055 (N_8055,N_7165,N_6645);
nor U8056 (N_8056,N_6333,N_6876);
and U8057 (N_8057,N_6844,N_7130);
and U8058 (N_8058,N_7081,N_5709);
and U8059 (N_8059,N_6415,N_7416);
or U8060 (N_8060,N_6733,N_6099);
nand U8061 (N_8061,N_5898,N_5311);
xor U8062 (N_8062,N_7438,N_6647);
nand U8063 (N_8063,N_5740,N_6251);
nand U8064 (N_8064,N_5710,N_6722);
nor U8065 (N_8065,N_7292,N_6478);
xnor U8066 (N_8066,N_5077,N_6033);
nand U8067 (N_8067,N_6979,N_5546);
nand U8068 (N_8068,N_5163,N_7125);
nor U8069 (N_8069,N_6597,N_6755);
nor U8070 (N_8070,N_7428,N_6400);
and U8071 (N_8071,N_6307,N_7091);
xnor U8072 (N_8072,N_6862,N_6454);
xor U8073 (N_8073,N_5794,N_6821);
xor U8074 (N_8074,N_6877,N_5458);
or U8075 (N_8075,N_7061,N_5123);
xnor U8076 (N_8076,N_6009,N_5361);
xor U8077 (N_8077,N_5108,N_6125);
nor U8078 (N_8078,N_5339,N_5572);
nor U8079 (N_8079,N_7103,N_5403);
nor U8080 (N_8080,N_6977,N_5623);
nor U8081 (N_8081,N_5336,N_6768);
nand U8082 (N_8082,N_6038,N_6932);
nand U8083 (N_8083,N_6159,N_6248);
and U8084 (N_8084,N_7380,N_6549);
and U8085 (N_8085,N_5616,N_5305);
xor U8086 (N_8086,N_7043,N_7413);
or U8087 (N_8087,N_5920,N_5650);
or U8088 (N_8088,N_5792,N_6300);
and U8089 (N_8089,N_6982,N_7198);
or U8090 (N_8090,N_7435,N_5309);
or U8091 (N_8091,N_5985,N_5490);
or U8092 (N_8092,N_7477,N_7375);
or U8093 (N_8093,N_5635,N_6025);
nor U8094 (N_8094,N_7331,N_6807);
nand U8095 (N_8095,N_6362,N_5896);
and U8096 (N_8096,N_5997,N_6425);
and U8097 (N_8097,N_6533,N_5963);
xor U8098 (N_8098,N_7291,N_6855);
nand U8099 (N_8099,N_5486,N_5949);
nand U8100 (N_8100,N_6561,N_6432);
nor U8101 (N_8101,N_5229,N_5391);
nor U8102 (N_8102,N_6310,N_7321);
nor U8103 (N_8103,N_6952,N_7243);
nor U8104 (N_8104,N_6762,N_6972);
nor U8105 (N_8105,N_7312,N_6880);
nor U8106 (N_8106,N_5844,N_5008);
and U8107 (N_8107,N_6660,N_6243);
nand U8108 (N_8108,N_5128,N_6926);
nand U8109 (N_8109,N_6846,N_7248);
and U8110 (N_8110,N_6391,N_7410);
nand U8111 (N_8111,N_6121,N_6137);
and U8112 (N_8112,N_6541,N_5376);
or U8113 (N_8113,N_6255,N_6005);
xor U8114 (N_8114,N_5131,N_5257);
and U8115 (N_8115,N_5956,N_7138);
and U8116 (N_8116,N_5212,N_6691);
nor U8117 (N_8117,N_5176,N_6341);
or U8118 (N_8118,N_6650,N_7326);
xnor U8119 (N_8119,N_7412,N_5824);
xnor U8120 (N_8120,N_7454,N_5242);
xor U8121 (N_8121,N_5535,N_6563);
and U8122 (N_8122,N_6669,N_7355);
xnor U8123 (N_8123,N_5134,N_5430);
and U8124 (N_8124,N_5364,N_6004);
xor U8125 (N_8125,N_6921,N_5998);
xnor U8126 (N_8126,N_6168,N_7334);
nor U8127 (N_8127,N_6356,N_5610);
nand U8128 (N_8128,N_5755,N_5838);
nand U8129 (N_8129,N_5653,N_5082);
xnor U8130 (N_8130,N_6915,N_6132);
xnor U8131 (N_8131,N_7385,N_5502);
xnor U8132 (N_8132,N_6109,N_7217);
xor U8133 (N_8133,N_7436,N_5090);
xor U8134 (N_8134,N_6735,N_5083);
nor U8135 (N_8135,N_5132,N_6110);
xnor U8136 (N_8136,N_6837,N_6729);
or U8137 (N_8137,N_6784,N_6054);
nand U8138 (N_8138,N_5894,N_5344);
xnor U8139 (N_8139,N_5517,N_6663);
and U8140 (N_8140,N_7048,N_6866);
and U8141 (N_8141,N_7449,N_6474);
and U8142 (N_8142,N_7345,N_5733);
xnor U8143 (N_8143,N_5405,N_5760);
nor U8144 (N_8144,N_6027,N_5603);
nand U8145 (N_8145,N_5079,N_5995);
nor U8146 (N_8146,N_5419,N_6810);
or U8147 (N_8147,N_5009,N_5183);
nand U8148 (N_8148,N_7027,N_5468);
or U8149 (N_8149,N_6022,N_5237);
and U8150 (N_8150,N_7324,N_7447);
xnor U8151 (N_8151,N_5296,N_5750);
or U8152 (N_8152,N_5507,N_7319);
and U8153 (N_8153,N_5243,N_7213);
or U8154 (N_8154,N_6247,N_7115);
nor U8155 (N_8155,N_5013,N_6530);
nand U8156 (N_8156,N_7189,N_5781);
xor U8157 (N_8157,N_5797,N_5136);
or U8158 (N_8158,N_6241,N_6107);
xnor U8159 (N_8159,N_7117,N_5573);
xor U8160 (N_8160,N_7220,N_6002);
nor U8161 (N_8161,N_7343,N_6742);
or U8162 (N_8162,N_6664,N_5932);
xnor U8163 (N_8163,N_6481,N_7159);
nand U8164 (N_8164,N_6443,N_6359);
nand U8165 (N_8165,N_7202,N_7028);
or U8166 (N_8166,N_6537,N_5062);
and U8167 (N_8167,N_6696,N_5472);
xnor U8168 (N_8168,N_7047,N_7228);
or U8169 (N_8169,N_7178,N_6643);
xor U8170 (N_8170,N_6690,N_6539);
xnor U8171 (N_8171,N_5165,N_5124);
xor U8172 (N_8172,N_6738,N_5037);
or U8173 (N_8173,N_5830,N_6468);
and U8174 (N_8174,N_5445,N_6177);
and U8175 (N_8175,N_6702,N_6919);
xnor U8176 (N_8176,N_5688,N_7074);
nor U8177 (N_8177,N_5671,N_6536);
nor U8178 (N_8178,N_6228,N_5922);
xor U8179 (N_8179,N_5354,N_7460);
nand U8180 (N_8180,N_6450,N_7396);
or U8181 (N_8181,N_6553,N_5066);
xor U8182 (N_8182,N_6370,N_5370);
or U8183 (N_8183,N_5886,N_6899);
nand U8184 (N_8184,N_6613,N_5050);
nand U8185 (N_8185,N_7297,N_6934);
nand U8186 (N_8186,N_6954,N_6182);
or U8187 (N_8187,N_6834,N_5550);
nand U8188 (N_8188,N_5199,N_6683);
and U8189 (N_8189,N_6715,N_7357);
xor U8190 (N_8190,N_6062,N_7370);
xor U8191 (N_8191,N_7308,N_5029);
xor U8192 (N_8192,N_5901,N_5587);
nor U8193 (N_8193,N_7287,N_7188);
or U8194 (N_8194,N_5686,N_6044);
xnor U8195 (N_8195,N_6452,N_6633);
and U8196 (N_8196,N_5735,N_6057);
or U8197 (N_8197,N_7424,N_5084);
nor U8198 (N_8198,N_7364,N_6491);
nor U8199 (N_8199,N_5080,N_6704);
or U8200 (N_8200,N_5734,N_6928);
nor U8201 (N_8201,N_7332,N_6218);
nand U8202 (N_8202,N_6793,N_7423);
or U8203 (N_8203,N_5516,N_5789);
and U8204 (N_8204,N_5574,N_6326);
xor U8205 (N_8205,N_6953,N_7335);
nor U8206 (N_8206,N_5073,N_6900);
nand U8207 (N_8207,N_6996,N_5114);
xor U8208 (N_8208,N_7226,N_7328);
or U8209 (N_8209,N_7246,N_5488);
and U8210 (N_8210,N_6165,N_5390);
xnor U8211 (N_8211,N_6071,N_5622);
xnor U8212 (N_8212,N_5149,N_5374);
or U8213 (N_8213,N_5597,N_6734);
or U8214 (N_8214,N_5982,N_5217);
xor U8215 (N_8215,N_5075,N_6765);
and U8216 (N_8216,N_5451,N_5655);
or U8217 (N_8217,N_7365,N_5441);
xnor U8218 (N_8218,N_6966,N_5900);
nor U8219 (N_8219,N_5294,N_5976);
nand U8220 (N_8220,N_5368,N_6361);
nor U8221 (N_8221,N_6801,N_5404);
nand U8222 (N_8222,N_5821,N_7251);
and U8223 (N_8223,N_6325,N_6640);
or U8224 (N_8224,N_5532,N_5524);
nand U8225 (N_8225,N_5091,N_6968);
or U8226 (N_8226,N_5629,N_6477);
nor U8227 (N_8227,N_5121,N_5278);
xor U8228 (N_8228,N_5043,N_6088);
nor U8229 (N_8229,N_6194,N_5306);
nand U8230 (N_8230,N_5615,N_6260);
nand U8231 (N_8231,N_5218,N_6313);
or U8232 (N_8232,N_6719,N_5918);
nand U8233 (N_8233,N_7296,N_7208);
nor U8234 (N_8234,N_6554,N_5939);
or U8235 (N_8235,N_6139,N_6374);
nor U8236 (N_8236,N_5178,N_6582);
or U8237 (N_8237,N_5564,N_6355);
and U8238 (N_8238,N_7190,N_7430);
nand U8239 (N_8239,N_6937,N_6383);
nand U8240 (N_8240,N_7141,N_6410);
xor U8241 (N_8241,N_7014,N_6369);
and U8242 (N_8242,N_6974,N_6214);
nor U8243 (N_8243,N_6438,N_5826);
and U8244 (N_8244,N_5518,N_5618);
nand U8245 (N_8245,N_7294,N_7086);
and U8246 (N_8246,N_7303,N_5979);
xor U8247 (N_8247,N_5925,N_5290);
nor U8248 (N_8248,N_7329,N_6595);
or U8249 (N_8249,N_6459,N_6828);
nor U8250 (N_8250,N_7199,N_7289);
nor U8251 (N_8251,N_5850,N_6789);
xor U8252 (N_8252,N_5426,N_7076);
and U8253 (N_8253,N_5983,N_6790);
xnor U8254 (N_8254,N_7279,N_5981);
nand U8255 (N_8255,N_6956,N_5194);
nand U8256 (N_8256,N_6558,N_7132);
and U8257 (N_8257,N_6569,N_6379);
nor U8258 (N_8258,N_6065,N_6095);
xor U8259 (N_8259,N_6659,N_5340);
xnor U8260 (N_8260,N_7142,N_7107);
nor U8261 (N_8261,N_6240,N_6674);
nand U8262 (N_8262,N_5479,N_6564);
and U8263 (N_8263,N_5303,N_6496);
or U8264 (N_8264,N_6420,N_5679);
and U8265 (N_8265,N_6780,N_6209);
and U8266 (N_8266,N_6237,N_5438);
xor U8267 (N_8267,N_5964,N_5094);
nand U8268 (N_8268,N_5231,N_5703);
nor U8269 (N_8269,N_5927,N_6495);
or U8270 (N_8270,N_5460,N_6751);
and U8271 (N_8271,N_7280,N_5352);
or U8272 (N_8272,N_6594,N_7453);
nand U8273 (N_8273,N_5656,N_7403);
xor U8274 (N_8274,N_5696,N_6857);
or U8275 (N_8275,N_6649,N_5714);
nand U8276 (N_8276,N_5017,N_7000);
nand U8277 (N_8277,N_7108,N_6818);
xor U8278 (N_8278,N_5501,N_6806);
xor U8279 (N_8279,N_7464,N_6460);
and U8280 (N_8280,N_6652,N_5774);
and U8281 (N_8281,N_5721,N_5494);
or U8282 (N_8282,N_6424,N_7301);
nand U8283 (N_8283,N_7007,N_6678);
xnor U8284 (N_8284,N_5300,N_5940);
nand U8285 (N_8285,N_6960,N_5814);
xor U8286 (N_8286,N_5133,N_6745);
or U8287 (N_8287,N_6349,N_7448);
nor U8288 (N_8288,N_5382,N_6202);
nand U8289 (N_8289,N_6250,N_5220);
nand U8290 (N_8290,N_7360,N_5996);
xor U8291 (N_8291,N_5771,N_6191);
nand U8292 (N_8292,N_5994,N_5661);
nand U8293 (N_8293,N_7457,N_7126);
xor U8294 (N_8294,N_6626,N_6890);
xnor U8295 (N_8295,N_5106,N_5911);
nor U8296 (N_8296,N_6980,N_6193);
nand U8297 (N_8297,N_5659,N_7481);
or U8298 (N_8298,N_5407,N_5297);
nor U8299 (N_8299,N_6914,N_6607);
nand U8300 (N_8300,N_6312,N_5870);
nor U8301 (N_8301,N_5355,N_7032);
or U8302 (N_8302,N_5762,N_5153);
nand U8303 (N_8303,N_6253,N_6529);
nand U8304 (N_8304,N_6737,N_5429);
xor U8305 (N_8305,N_6196,N_5119);
nand U8306 (N_8306,N_5113,N_5046);
nor U8307 (N_8307,N_7476,N_6464);
or U8308 (N_8308,N_5845,N_5307);
xor U8309 (N_8309,N_6414,N_6948);
nand U8310 (N_8310,N_5836,N_5961);
nand U8311 (N_8311,N_7475,N_5125);
nand U8312 (N_8312,N_5791,N_5069);
nor U8313 (N_8313,N_6708,N_6833);
or U8314 (N_8314,N_7162,N_5211);
xor U8315 (N_8315,N_5770,N_5298);
nor U8316 (N_8316,N_6426,N_6291);
nor U8317 (N_8317,N_6562,N_6001);
nor U8318 (N_8318,N_6382,N_5055);
nand U8319 (N_8319,N_5492,N_6991);
nand U8320 (N_8320,N_5459,N_7295);
xnor U8321 (N_8321,N_5240,N_7275);
and U8322 (N_8322,N_5435,N_5676);
nand U8323 (N_8323,N_5566,N_7354);
nor U8324 (N_8324,N_6318,N_6943);
nand U8325 (N_8325,N_5807,N_6642);
nand U8326 (N_8326,N_5481,N_5974);
xnor U8327 (N_8327,N_6093,N_5325);
and U8328 (N_8328,N_5215,N_6463);
nand U8329 (N_8329,N_5261,N_5892);
or U8330 (N_8330,N_6019,N_6466);
and U8331 (N_8331,N_6519,N_7390);
nor U8332 (N_8332,N_6188,N_5011);
nand U8333 (N_8333,N_5262,N_6145);
or U8334 (N_8334,N_5085,N_6332);
nand U8335 (N_8335,N_7304,N_6045);
nand U8336 (N_8336,N_6653,N_5667);
xnor U8337 (N_8337,N_7469,N_6887);
or U8338 (N_8338,N_7054,N_6123);
or U8339 (N_8339,N_5723,N_5575);
xnor U8340 (N_8340,N_6066,N_5036);
xor U8341 (N_8341,N_6681,N_5991);
and U8342 (N_8342,N_5139,N_5680);
and U8343 (N_8343,N_6262,N_7070);
or U8344 (N_8344,N_7418,N_5802);
or U8345 (N_8345,N_6581,N_6504);
nor U8346 (N_8346,N_6082,N_6035);
nor U8347 (N_8347,N_6913,N_7143);
or U8348 (N_8348,N_6739,N_6163);
or U8349 (N_8349,N_5301,N_6032);
or U8350 (N_8350,N_5543,N_5704);
xor U8351 (N_8351,N_6467,N_6797);
xnor U8352 (N_8352,N_5729,N_6339);
nand U8353 (N_8353,N_5400,N_6335);
nand U8354 (N_8354,N_5751,N_6124);
nor U8355 (N_8355,N_6545,N_6747);
nand U8356 (N_8356,N_6028,N_6515);
or U8357 (N_8357,N_5216,N_5580);
or U8358 (N_8358,N_6246,N_6584);
xnor U8359 (N_8359,N_6059,N_6106);
nor U8360 (N_8360,N_6162,N_5847);
and U8361 (N_8361,N_7065,N_6731);
and U8362 (N_8362,N_6552,N_6272);
and U8363 (N_8363,N_7210,N_7182);
nor U8364 (N_8364,N_6392,N_6288);
nor U8365 (N_8365,N_6842,N_6772);
xnor U8366 (N_8366,N_7015,N_7264);
nor U8367 (N_8367,N_7106,N_6863);
nand U8368 (N_8368,N_6699,N_6030);
nand U8369 (N_8369,N_5749,N_6671);
or U8370 (N_8370,N_5135,N_6222);
xnor U8371 (N_8371,N_6993,N_6204);
nor U8372 (N_8372,N_6364,N_6235);
nand U8373 (N_8373,N_7478,N_6894);
and U8374 (N_8374,N_5367,N_7105);
nor U8375 (N_8375,N_7150,N_5347);
and U8376 (N_8376,N_5664,N_5730);
xor U8377 (N_8377,N_7426,N_6396);
xor U8378 (N_8378,N_6946,N_6069);
nor U8379 (N_8379,N_7079,N_6518);
xor U8380 (N_8380,N_5504,N_7145);
or U8381 (N_8381,N_6945,N_5663);
or U8382 (N_8382,N_7398,N_5980);
xnor U8383 (N_8383,N_6390,N_5440);
nand U8384 (N_8384,N_6771,N_5913);
xnor U8385 (N_8385,N_6112,N_5154);
or U8386 (N_8386,N_5707,N_5984);
nand U8387 (N_8387,N_6693,N_5931);
or U8388 (N_8388,N_6487,N_6254);
nand U8389 (N_8389,N_6602,N_5675);
and U8390 (N_8390,N_5293,N_5177);
and U8391 (N_8391,N_6439,N_6878);
xor U8392 (N_8392,N_6918,N_5511);
or U8393 (N_8393,N_6480,N_5917);
nand U8394 (N_8394,N_6286,N_6546);
or U8395 (N_8395,N_7310,N_7387);
and U8396 (N_8396,N_5070,N_6169);
or U8397 (N_8397,N_7323,N_6920);
xnor U8398 (N_8398,N_6041,N_5482);
and U8399 (N_8399,N_6550,N_5553);
xnor U8400 (N_8400,N_6133,N_6579);
nor U8401 (N_8401,N_5767,N_5337);
xnor U8402 (N_8402,N_6084,N_7060);
or U8403 (N_8403,N_5387,N_6618);
nand U8404 (N_8404,N_5570,N_6870);
nor U8405 (N_8405,N_6489,N_5161);
nand U8406 (N_8406,N_5613,N_7293);
nand U8407 (N_8407,N_5434,N_5423);
nand U8408 (N_8408,N_5592,N_5843);
or U8409 (N_8409,N_5595,N_7483);
xor U8410 (N_8410,N_7147,N_5833);
and U8411 (N_8411,N_5608,N_6907);
and U8412 (N_8412,N_6486,N_6021);
and U8413 (N_8413,N_5039,N_5752);
xnor U8414 (N_8414,N_6666,N_6883);
or U8415 (N_8415,N_6596,N_6754);
nand U8416 (N_8416,N_5764,N_6836);
or U8417 (N_8417,N_6378,N_7200);
or U8418 (N_8418,N_5586,N_5443);
nand U8419 (N_8419,N_6994,N_5692);
nand U8420 (N_8420,N_7111,N_5875);
nor U8421 (N_8421,N_5880,N_7078);
xor U8422 (N_8422,N_5001,N_5712);
or U8423 (N_8423,N_6752,N_6999);
or U8424 (N_8424,N_7053,N_6721);
nand U8425 (N_8425,N_5945,N_7462);
and U8426 (N_8426,N_5741,N_6053);
and U8427 (N_8427,N_5455,N_5674);
nor U8428 (N_8428,N_6258,N_5528);
nor U8429 (N_8429,N_5171,N_6651);
or U8430 (N_8430,N_6289,N_5399);
nor U8431 (N_8431,N_6263,N_6925);
nand U8432 (N_8432,N_5003,N_6732);
or U8433 (N_8433,N_6770,N_7372);
nand U8434 (N_8434,N_5719,N_5757);
and U8435 (N_8435,N_7154,N_6230);
and U8436 (N_8436,N_6958,N_5531);
nand U8437 (N_8437,N_5048,N_5280);
xor U8438 (N_8438,N_7282,N_5395);
nand U8439 (N_8439,N_5338,N_5397);
or U8440 (N_8440,N_6446,N_6184);
xor U8441 (N_8441,N_7062,N_5758);
or U8442 (N_8442,N_7031,N_6435);
or U8443 (N_8443,N_6483,N_5005);
nor U8444 (N_8444,N_5837,N_6524);
nor U8445 (N_8445,N_6490,N_6279);
and U8446 (N_8446,N_6854,N_5625);
or U8447 (N_8447,N_6930,N_5313);
and U8448 (N_8448,N_7044,N_6407);
nor U8449 (N_8449,N_7371,N_7368);
and U8450 (N_8450,N_5416,N_6152);
nand U8451 (N_8451,N_6087,N_5902);
nor U8452 (N_8452,N_5804,N_6590);
xor U8453 (N_8453,N_6305,N_5778);
nand U8454 (N_8454,N_7051,N_6604);
or U8455 (N_8455,N_5016,N_7055);
nand U8456 (N_8456,N_5076,N_7350);
nand U8457 (N_8457,N_5358,N_6189);
nand U8458 (N_8458,N_6249,N_6749);
and U8459 (N_8459,N_5151,N_5437);
or U8460 (N_8460,N_6559,N_7381);
xor U8461 (N_8461,N_7167,N_6157);
xor U8462 (N_8462,N_7274,N_5453);
nor U8463 (N_8463,N_6274,N_6348);
nor U8464 (N_8464,N_7411,N_5772);
or U8465 (N_8465,N_5222,N_7461);
nor U8466 (N_8466,N_6824,N_5115);
nand U8467 (N_8467,N_7153,N_5649);
xnor U8468 (N_8468,N_5876,N_6540);
xor U8469 (N_8469,N_6668,N_6360);
xor U8470 (N_8470,N_6976,N_5923);
and U8471 (N_8471,N_6614,N_6371);
and U8472 (N_8472,N_5341,N_6838);
and U8473 (N_8473,N_7157,N_6884);
or U8474 (N_8474,N_6621,N_6718);
nor U8475 (N_8475,N_6327,N_6667);
xnor U8476 (N_8476,N_7352,N_5579);
and U8477 (N_8477,N_5255,N_6869);
or U8478 (N_8478,N_7314,N_5787);
or U8479 (N_8479,N_7203,N_6819);
nand U8480 (N_8480,N_6843,N_7494);
and U8481 (N_8481,N_5617,N_6085);
xnor U8482 (N_8482,N_5739,N_6160);
and U8483 (N_8483,N_5602,N_6917);
xor U8484 (N_8484,N_5856,N_5271);
xnor U8485 (N_8485,N_5819,N_7495);
nor U8486 (N_8486,N_7422,N_6924);
and U8487 (N_8487,N_6042,N_6358);
or U8488 (N_8488,N_5487,N_7270);
and U8489 (N_8489,N_5853,N_6703);
xor U8490 (N_8490,N_5722,N_5144);
and U8491 (N_8491,N_5477,N_6963);
nor U8492 (N_8492,N_5024,N_5556);
nor U8493 (N_8493,N_7135,N_5465);
nand U8494 (N_8494,N_7374,N_7489);
nand U8495 (N_8495,N_6180,N_5329);
or U8496 (N_8496,N_6416,N_7004);
nand U8497 (N_8497,N_5601,N_6508);
and U8498 (N_8498,N_6498,N_6893);
or U8499 (N_8499,N_6299,N_6986);
nand U8500 (N_8500,N_5977,N_5099);
and U8501 (N_8501,N_6593,N_5640);
nand U8502 (N_8502,N_6580,N_7209);
xnor U8503 (N_8503,N_6334,N_5118);
nand U8504 (N_8504,N_5277,N_6872);
and U8505 (N_8505,N_7315,N_5025);
nor U8506 (N_8506,N_5530,N_6712);
nor U8507 (N_8507,N_7249,N_6086);
nor U8508 (N_8508,N_6113,N_6079);
nor U8509 (N_8509,N_5882,N_7224);
xor U8510 (N_8510,N_6623,N_6510);
and U8511 (N_8511,N_7172,N_5829);
nor U8512 (N_8512,N_7020,N_7113);
xor U8513 (N_8513,N_6171,N_5647);
nand U8514 (N_8514,N_5657,N_5088);
nand U8515 (N_8515,N_6126,N_6131);
nor U8516 (N_8516,N_5392,N_6543);
and U8517 (N_8517,N_5236,N_7322);
and U8518 (N_8518,N_6381,N_7223);
xnor U8519 (N_8519,N_7492,N_5056);
nand U8520 (N_8520,N_6627,N_6816);
or U8521 (N_8521,N_6499,N_6290);
xnor U8522 (N_8522,N_6800,N_6904);
xnor U8523 (N_8523,N_6128,N_6502);
nand U8524 (N_8524,N_7333,N_6881);
or U8525 (N_8525,N_7006,N_7104);
nor U8526 (N_8526,N_6736,N_5910);
and U8527 (N_8527,N_6517,N_6329);
nand U8528 (N_8528,N_5879,N_6174);
or U8529 (N_8529,N_5442,N_7039);
nor U8530 (N_8530,N_6200,N_6796);
nand U8531 (N_8531,N_5322,N_6219);
or U8532 (N_8532,N_7095,N_6984);
xor U8533 (N_8533,N_5916,N_7185);
xor U8534 (N_8534,N_7227,N_5064);
nor U8535 (N_8535,N_6372,N_7003);
nor U8536 (N_8536,N_6638,N_6592);
xnor U8537 (N_8537,N_6617,N_6311);
nor U8538 (N_8538,N_5899,N_7093);
nor U8539 (N_8539,N_6615,N_6746);
nor U8540 (N_8540,N_7302,N_5506);
nor U8541 (N_8541,N_7156,N_5061);
and U8542 (N_8542,N_6935,N_5806);
xnor U8543 (N_8543,N_7024,N_5926);
or U8544 (N_8544,N_5238,N_5520);
xor U8545 (N_8545,N_5765,N_6293);
nor U8546 (N_8546,N_5860,N_5138);
xnor U8547 (N_8547,N_6902,N_6199);
nor U8548 (N_8548,N_7175,N_5281);
xnor U8549 (N_8549,N_7163,N_7233);
xnor U8550 (N_8550,N_6336,N_5883);
nand U8551 (N_8551,N_5415,N_5810);
nor U8552 (N_8552,N_6026,N_5698);
or U8553 (N_8553,N_7201,N_5353);
xnor U8554 (N_8554,N_7136,N_5745);
nor U8555 (N_8555,N_6297,N_5912);
nor U8556 (N_8556,N_6575,N_6758);
and U8557 (N_8557,N_7298,N_5146);
or U8558 (N_8558,N_5308,N_5110);
nand U8559 (N_8559,N_6585,N_6726);
xnor U8560 (N_8560,N_7144,N_5706);
nand U8561 (N_8561,N_6437,N_6776);
and U8562 (N_8562,N_5259,N_7234);
nor U8563 (N_8563,N_5383,N_7231);
or U8564 (N_8564,N_6220,N_6679);
xor U8565 (N_8565,N_5454,N_5864);
nor U8566 (N_8566,N_5708,N_7277);
xor U8567 (N_8567,N_7258,N_5529);
and U8568 (N_8568,N_5241,N_7257);
nor U8569 (N_8569,N_6389,N_5006);
xor U8570 (N_8570,N_5137,N_5269);
nor U8571 (N_8571,N_6639,N_6692);
or U8572 (N_8572,N_7392,N_5444);
and U8573 (N_8573,N_5512,N_5175);
nor U8574 (N_8574,N_6118,N_6849);
nand U8575 (N_8575,N_5266,N_7317);
xor U8576 (N_8576,N_5157,N_7194);
xnor U8577 (N_8577,N_6848,N_7193);
or U8578 (N_8578,N_6273,N_7307);
nand U8579 (N_8579,N_5276,N_7255);
xor U8580 (N_8580,N_6346,N_7408);
xnor U8581 (N_8581,N_6146,N_5321);
or U8582 (N_8582,N_6694,N_5291);
xor U8583 (N_8583,N_5245,N_6698);
and U8584 (N_8584,N_6898,N_7286);
xnor U8585 (N_8585,N_5285,N_6395);
xor U8586 (N_8586,N_5475,N_5820);
nor U8587 (N_8587,N_6365,N_6940);
nor U8588 (N_8588,N_5846,N_5155);
nor U8589 (N_8589,N_5057,N_6864);
xnor U8590 (N_8590,N_5800,N_5954);
or U8591 (N_8591,N_6270,N_7336);
xor U8592 (N_8592,N_6532,N_6277);
and U8593 (N_8593,N_7030,N_7379);
or U8594 (N_8594,N_7067,N_5941);
nand U8595 (N_8595,N_7316,N_6388);
nor U8596 (N_8596,N_6910,N_5164);
and U8597 (N_8597,N_6485,N_5822);
and U8598 (N_8598,N_6611,N_6576);
nor U8599 (N_8599,N_5239,N_6761);
and U8600 (N_8600,N_7444,N_5727);
and U8601 (N_8601,N_5519,N_6303);
nand U8602 (N_8602,N_5447,N_5318);
nand U8603 (N_8603,N_5421,N_5101);
and U8604 (N_8604,N_7002,N_5780);
or U8605 (N_8605,N_6895,N_7473);
nand U8606 (N_8606,N_5508,N_5889);
or U8607 (N_8607,N_7244,N_6080);
and U8608 (N_8608,N_6760,N_6151);
nor U8609 (N_8609,N_7269,N_6723);
nand U8610 (N_8610,N_6344,N_6143);
or U8611 (N_8611,N_6635,N_5097);
or U8612 (N_8612,N_5224,N_7041);
nor U8613 (N_8613,N_5433,N_6399);
or U8614 (N_8614,N_7169,N_7353);
or U8615 (N_8615,N_7401,N_6511);
and U8616 (N_8616,N_6342,N_6969);
or U8617 (N_8617,N_6014,N_6321);
and U8618 (N_8618,N_7173,N_6472);
and U8619 (N_8619,N_7266,N_5071);
or U8620 (N_8620,N_7327,N_5343);
or U8621 (N_8621,N_5539,N_6097);
xor U8622 (N_8622,N_5464,N_6527);
nand U8623 (N_8623,N_7009,N_5933);
xnor U8624 (N_8624,N_5641,N_6453);
xor U8625 (N_8625,N_6441,N_6845);
nand U8626 (N_8626,N_7050,N_5182);
nand U8627 (N_8627,N_5737,N_6049);
nand U8628 (N_8628,N_5682,N_7456);
xor U8629 (N_8629,N_6822,N_5952);
nor U8630 (N_8630,N_5235,N_7137);
nand U8631 (N_8631,N_5930,N_7450);
xor U8632 (N_8632,N_5166,N_7420);
or U8633 (N_8633,N_5371,N_5992);
and U8634 (N_8634,N_5747,N_5924);
or U8635 (N_8635,N_7037,N_5858);
xor U8636 (N_8636,N_5122,N_5660);
and U8637 (N_8637,N_7439,N_5717);
nand U8638 (N_8638,N_5840,N_6119);
or U8639 (N_8639,N_5540,N_7383);
and U8640 (N_8640,N_5715,N_5051);
nand U8641 (N_8641,N_7183,N_6697);
xnor U8642 (N_8642,N_6292,N_5214);
xnor U8643 (N_8643,N_6178,N_6965);
nor U8644 (N_8644,N_6363,N_5773);
and U8645 (N_8645,N_6577,N_5332);
nor U8646 (N_8646,N_6257,N_7146);
xnor U8647 (N_8647,N_6646,N_5129);
and U8648 (N_8648,N_6756,N_5953);
or U8649 (N_8649,N_6572,N_6179);
xor U8650 (N_8650,N_5483,N_5589);
or U8651 (N_8651,N_6015,N_5694);
or U8652 (N_8652,N_6242,N_7168);
or U8653 (N_8653,N_5315,N_6122);
nor U8654 (N_8654,N_5389,N_5244);
and U8655 (N_8655,N_5651,N_7040);
xnor U8656 (N_8656,N_5160,N_6418);
nand U8657 (N_8657,N_7133,N_5699);
xor U8658 (N_8658,N_6328,N_5109);
and U8659 (N_8659,N_5469,N_7262);
or U8660 (N_8660,N_5042,N_6315);
or U8661 (N_8661,N_5606,N_5605);
xor U8662 (N_8662,N_6661,N_5746);
or U8663 (N_8663,N_7281,N_5485);
nand U8664 (N_8664,N_6757,N_5470);
nor U8665 (N_8665,N_6628,N_5095);
nand U8666 (N_8666,N_6267,N_6283);
or U8667 (N_8667,N_6547,N_6104);
nand U8668 (N_8668,N_6631,N_5033);
and U8669 (N_8669,N_5093,N_5777);
nand U8670 (N_8670,N_6600,N_6083);
and U8671 (N_8671,N_6497,N_7468);
or U8672 (N_8672,N_6525,N_5295);
or U8673 (N_8673,N_6166,N_5263);
xor U8674 (N_8674,N_7094,N_6942);
nor U8675 (N_8675,N_6324,N_5105);
nor U8676 (N_8676,N_5448,N_7484);
nor U8677 (N_8677,N_5938,N_6377);
or U8678 (N_8678,N_7176,N_6931);
nor U8679 (N_8679,N_7088,N_7339);
and U8680 (N_8680,N_7124,N_7011);
xor U8681 (N_8681,N_5776,N_7123);
nor U8682 (N_8682,N_7052,N_6759);
nand U8683 (N_8683,N_7184,N_6302);
and U8684 (N_8684,N_5342,N_5621);
nor U8685 (N_8685,N_6589,N_6852);
xnor U8686 (N_8686,N_6981,N_7337);
or U8687 (N_8687,N_5598,N_6903);
xnor U8688 (N_8688,N_6764,N_7414);
and U8689 (N_8689,N_6578,N_6725);
nand U8690 (N_8690,N_6261,N_7273);
or U8691 (N_8691,N_5140,N_5204);
or U8692 (N_8692,N_6492,N_5834);
nand U8693 (N_8693,N_7382,N_5966);
and U8694 (N_8694,N_6275,N_5497);
and U8695 (N_8695,N_5578,N_6276);
nor U8696 (N_8696,N_7160,N_7290);
nand U8697 (N_8697,N_6829,N_5074);
xor U8698 (N_8698,N_7119,N_5324);
and U8699 (N_8699,N_6861,N_6304);
and U8700 (N_8700,N_7057,N_6156);
xor U8701 (N_8701,N_5962,N_6808);
or U8702 (N_8702,N_7443,N_6357);
nand U8703 (N_8703,N_5279,N_6398);
or U8704 (N_8704,N_5803,N_6433);
and U8705 (N_8705,N_5614,N_5252);
nand U8706 (N_8706,N_5032,N_5759);
or U8707 (N_8707,N_5978,N_6997);
and U8708 (N_8708,N_5868,N_6556);
nor U8709 (N_8709,N_6720,N_6875);
xor U8710 (N_8710,N_7451,N_7072);
and U8711 (N_8711,N_7417,N_7393);
nor U8712 (N_8712,N_7102,N_5360);
xor U8713 (N_8713,N_5890,N_5446);
and U8714 (N_8714,N_6406,N_5150);
nor U8715 (N_8715,N_5232,N_6077);
or U8716 (N_8716,N_5254,N_5330);
or U8717 (N_8717,N_6744,N_5034);
nor U8718 (N_8718,N_6207,N_7139);
and U8719 (N_8719,N_6682,N_6036);
xor U8720 (N_8720,N_6528,N_5333);
nand U8721 (N_8721,N_6317,N_6296);
or U8722 (N_8722,N_7259,N_5873);
nor U8723 (N_8723,N_6225,N_5246);
or U8724 (N_8724,N_6413,N_5221);
xor U8725 (N_8725,N_5521,N_5872);
xor U8726 (N_8726,N_6657,N_6609);
and U8727 (N_8727,N_7196,N_6164);
and U8728 (N_8728,N_5631,N_5104);
nor U8729 (N_8729,N_5068,N_5393);
nor U8730 (N_8730,N_6827,N_5683);
nand U8731 (N_8731,N_7239,N_5701);
xor U8732 (N_8732,N_6505,N_5264);
nor U8733 (N_8733,N_6076,N_6964);
nand U8734 (N_8734,N_5230,N_5908);
xor U8735 (N_8735,N_7127,N_6670);
nor U8736 (N_8736,N_7216,N_7437);
nand U8737 (N_8737,N_5018,N_6513);
and U8738 (N_8738,N_5474,N_6449);
nor U8739 (N_8739,N_5725,N_5409);
or U8740 (N_8740,N_7077,N_5457);
nand U8741 (N_8741,N_6195,N_6886);
nand U8742 (N_8742,N_5672,N_5818);
nor U8743 (N_8743,N_5779,N_5147);
and U8744 (N_8744,N_6190,N_5208);
and U8745 (N_8745,N_5040,N_6185);
nand U8746 (N_8746,N_6955,N_5673);
nand U8747 (N_8747,N_6798,N_5988);
or U8748 (N_8748,N_6068,N_5697);
nand U8749 (N_8749,N_7222,N_5406);
nor U8750 (N_8750,N_6932,N_6228);
and U8751 (N_8751,N_5963,N_6351);
nand U8752 (N_8752,N_6568,N_6457);
nand U8753 (N_8753,N_5690,N_5867);
or U8754 (N_8754,N_5030,N_7099);
nand U8755 (N_8755,N_7436,N_6699);
or U8756 (N_8756,N_5742,N_6255);
nor U8757 (N_8757,N_6896,N_5392);
or U8758 (N_8758,N_6193,N_6273);
or U8759 (N_8759,N_7300,N_5498);
and U8760 (N_8760,N_5816,N_5591);
nand U8761 (N_8761,N_6017,N_5420);
and U8762 (N_8762,N_6533,N_6880);
and U8763 (N_8763,N_6982,N_6813);
nor U8764 (N_8764,N_5167,N_5696);
nor U8765 (N_8765,N_6021,N_7269);
and U8766 (N_8766,N_7135,N_7078);
nor U8767 (N_8767,N_6730,N_6930);
nand U8768 (N_8768,N_5425,N_7032);
nor U8769 (N_8769,N_5025,N_5023);
or U8770 (N_8770,N_6579,N_7488);
nor U8771 (N_8771,N_6029,N_6014);
nand U8772 (N_8772,N_5763,N_7012);
nand U8773 (N_8773,N_5401,N_5106);
or U8774 (N_8774,N_7215,N_7312);
nand U8775 (N_8775,N_7116,N_6894);
or U8776 (N_8776,N_6181,N_6368);
xor U8777 (N_8777,N_5366,N_5705);
nor U8778 (N_8778,N_5300,N_6047);
nand U8779 (N_8779,N_7261,N_5281);
nand U8780 (N_8780,N_7279,N_6913);
nor U8781 (N_8781,N_6057,N_5292);
nor U8782 (N_8782,N_5150,N_5807);
and U8783 (N_8783,N_5297,N_7162);
or U8784 (N_8784,N_7189,N_7143);
and U8785 (N_8785,N_7175,N_5098);
and U8786 (N_8786,N_7421,N_5846);
nand U8787 (N_8787,N_6273,N_5831);
nand U8788 (N_8788,N_5479,N_5796);
xnor U8789 (N_8789,N_5050,N_6546);
or U8790 (N_8790,N_5078,N_5765);
xor U8791 (N_8791,N_7486,N_6506);
and U8792 (N_8792,N_5660,N_7243);
nand U8793 (N_8793,N_7130,N_6967);
or U8794 (N_8794,N_6193,N_6556);
nand U8795 (N_8795,N_6259,N_5405);
or U8796 (N_8796,N_7216,N_6153);
nand U8797 (N_8797,N_6308,N_7198);
nor U8798 (N_8798,N_7230,N_6886);
and U8799 (N_8799,N_5064,N_6727);
or U8800 (N_8800,N_5269,N_7350);
xnor U8801 (N_8801,N_6953,N_6206);
nand U8802 (N_8802,N_5901,N_6178);
or U8803 (N_8803,N_5308,N_5860);
and U8804 (N_8804,N_6953,N_6748);
or U8805 (N_8805,N_6261,N_6145);
or U8806 (N_8806,N_7101,N_6025);
nor U8807 (N_8807,N_6990,N_6018);
or U8808 (N_8808,N_6232,N_5915);
nand U8809 (N_8809,N_6379,N_5172);
or U8810 (N_8810,N_5864,N_5146);
xnor U8811 (N_8811,N_5300,N_7130);
and U8812 (N_8812,N_6978,N_7204);
and U8813 (N_8813,N_5081,N_5829);
or U8814 (N_8814,N_5243,N_6465);
and U8815 (N_8815,N_7399,N_7465);
and U8816 (N_8816,N_5366,N_5721);
xnor U8817 (N_8817,N_6190,N_7364);
and U8818 (N_8818,N_6381,N_6282);
or U8819 (N_8819,N_5714,N_5495);
nor U8820 (N_8820,N_6713,N_6561);
or U8821 (N_8821,N_6836,N_7236);
nor U8822 (N_8822,N_6391,N_5272);
xnor U8823 (N_8823,N_7238,N_6490);
and U8824 (N_8824,N_5787,N_6048);
xor U8825 (N_8825,N_5185,N_5616);
and U8826 (N_8826,N_5414,N_5514);
nor U8827 (N_8827,N_6948,N_6510);
xnor U8828 (N_8828,N_6151,N_5878);
nor U8829 (N_8829,N_6638,N_7200);
or U8830 (N_8830,N_5343,N_7249);
xnor U8831 (N_8831,N_5382,N_5886);
nand U8832 (N_8832,N_6695,N_6067);
nor U8833 (N_8833,N_5541,N_5777);
or U8834 (N_8834,N_6012,N_5778);
or U8835 (N_8835,N_5290,N_7239);
nand U8836 (N_8836,N_6761,N_6591);
xor U8837 (N_8837,N_7415,N_5426);
nor U8838 (N_8838,N_7306,N_6560);
xor U8839 (N_8839,N_5206,N_7070);
or U8840 (N_8840,N_6960,N_5492);
xor U8841 (N_8841,N_6266,N_5094);
or U8842 (N_8842,N_5294,N_5720);
xor U8843 (N_8843,N_5607,N_5519);
xnor U8844 (N_8844,N_6746,N_7282);
and U8845 (N_8845,N_5146,N_7246);
and U8846 (N_8846,N_6678,N_6072);
nor U8847 (N_8847,N_6118,N_7488);
nand U8848 (N_8848,N_6175,N_7185);
nor U8849 (N_8849,N_6408,N_5307);
nand U8850 (N_8850,N_5536,N_7346);
and U8851 (N_8851,N_5778,N_6149);
xor U8852 (N_8852,N_5730,N_5826);
and U8853 (N_8853,N_7383,N_6094);
xnor U8854 (N_8854,N_7152,N_6649);
or U8855 (N_8855,N_5944,N_6211);
nand U8856 (N_8856,N_5842,N_5571);
and U8857 (N_8857,N_6476,N_5542);
and U8858 (N_8858,N_5958,N_7124);
nor U8859 (N_8859,N_6754,N_6057);
and U8860 (N_8860,N_7223,N_5508);
and U8861 (N_8861,N_5277,N_6304);
and U8862 (N_8862,N_6701,N_6431);
nor U8863 (N_8863,N_7473,N_5584);
nand U8864 (N_8864,N_6800,N_6673);
nand U8865 (N_8865,N_5533,N_6115);
nand U8866 (N_8866,N_7060,N_6412);
or U8867 (N_8867,N_5147,N_6411);
or U8868 (N_8868,N_5406,N_6531);
or U8869 (N_8869,N_6242,N_5904);
nand U8870 (N_8870,N_5891,N_6324);
xor U8871 (N_8871,N_6247,N_6203);
nor U8872 (N_8872,N_5839,N_5877);
and U8873 (N_8873,N_5324,N_7420);
nor U8874 (N_8874,N_6884,N_7308);
nor U8875 (N_8875,N_5342,N_5874);
xor U8876 (N_8876,N_6565,N_5114);
or U8877 (N_8877,N_7071,N_5415);
nor U8878 (N_8878,N_6990,N_6325);
xnor U8879 (N_8879,N_5236,N_6335);
and U8880 (N_8880,N_7394,N_5993);
nand U8881 (N_8881,N_5511,N_6575);
nor U8882 (N_8882,N_5778,N_7247);
nand U8883 (N_8883,N_5210,N_5073);
xnor U8884 (N_8884,N_6988,N_6924);
and U8885 (N_8885,N_6881,N_7052);
xor U8886 (N_8886,N_6042,N_6731);
nor U8887 (N_8887,N_5095,N_7256);
xnor U8888 (N_8888,N_5314,N_7219);
and U8889 (N_8889,N_5745,N_6883);
or U8890 (N_8890,N_6069,N_7440);
xor U8891 (N_8891,N_5848,N_7272);
xor U8892 (N_8892,N_7441,N_5491);
nor U8893 (N_8893,N_6687,N_5480);
nand U8894 (N_8894,N_6339,N_6694);
and U8895 (N_8895,N_6938,N_5457);
or U8896 (N_8896,N_5588,N_5956);
xor U8897 (N_8897,N_6727,N_6713);
nor U8898 (N_8898,N_5845,N_6916);
and U8899 (N_8899,N_7047,N_7478);
nor U8900 (N_8900,N_6102,N_5600);
or U8901 (N_8901,N_5655,N_5103);
nor U8902 (N_8902,N_7019,N_5655);
xor U8903 (N_8903,N_5766,N_5695);
or U8904 (N_8904,N_6433,N_6505);
nand U8905 (N_8905,N_6648,N_7079);
or U8906 (N_8906,N_6873,N_7080);
xnor U8907 (N_8907,N_5179,N_5669);
and U8908 (N_8908,N_5001,N_6502);
nand U8909 (N_8909,N_5717,N_5896);
or U8910 (N_8910,N_6113,N_5420);
and U8911 (N_8911,N_7051,N_5049);
xor U8912 (N_8912,N_6387,N_6361);
xnor U8913 (N_8913,N_6587,N_7288);
and U8914 (N_8914,N_6962,N_6550);
and U8915 (N_8915,N_6086,N_6465);
or U8916 (N_8916,N_7416,N_6543);
nor U8917 (N_8917,N_5402,N_5775);
nor U8918 (N_8918,N_5112,N_5479);
or U8919 (N_8919,N_5186,N_7036);
nor U8920 (N_8920,N_6772,N_6083);
or U8921 (N_8921,N_6561,N_7472);
nor U8922 (N_8922,N_5166,N_5062);
xnor U8923 (N_8923,N_5357,N_5369);
or U8924 (N_8924,N_6150,N_5552);
or U8925 (N_8925,N_6175,N_7157);
nor U8926 (N_8926,N_6242,N_5026);
nor U8927 (N_8927,N_6901,N_5125);
nand U8928 (N_8928,N_5570,N_5949);
nor U8929 (N_8929,N_5178,N_5376);
xnor U8930 (N_8930,N_6220,N_5523);
nor U8931 (N_8931,N_5938,N_6679);
nand U8932 (N_8932,N_6079,N_5059);
or U8933 (N_8933,N_5176,N_6370);
or U8934 (N_8934,N_5490,N_6005);
nand U8935 (N_8935,N_5363,N_5258);
xnor U8936 (N_8936,N_5549,N_5171);
xor U8937 (N_8937,N_6797,N_7284);
and U8938 (N_8938,N_7173,N_6106);
nand U8939 (N_8939,N_6185,N_5045);
or U8940 (N_8940,N_6683,N_6167);
or U8941 (N_8941,N_6035,N_6614);
nor U8942 (N_8942,N_5638,N_5396);
or U8943 (N_8943,N_6784,N_7001);
nand U8944 (N_8944,N_7087,N_7184);
nor U8945 (N_8945,N_6910,N_7142);
or U8946 (N_8946,N_6429,N_6437);
nand U8947 (N_8947,N_6711,N_7063);
or U8948 (N_8948,N_5687,N_7137);
nor U8949 (N_8949,N_5354,N_6367);
nand U8950 (N_8950,N_5472,N_6143);
xor U8951 (N_8951,N_6136,N_7264);
nor U8952 (N_8952,N_7066,N_5754);
xnor U8953 (N_8953,N_5873,N_7081);
or U8954 (N_8954,N_6661,N_6428);
nand U8955 (N_8955,N_6640,N_7132);
or U8956 (N_8956,N_7079,N_6011);
nor U8957 (N_8957,N_6447,N_6065);
nand U8958 (N_8958,N_6736,N_5208);
xor U8959 (N_8959,N_6810,N_6277);
nor U8960 (N_8960,N_5652,N_5320);
nor U8961 (N_8961,N_6383,N_7049);
nand U8962 (N_8962,N_7366,N_6882);
nor U8963 (N_8963,N_6210,N_6790);
or U8964 (N_8964,N_7024,N_5179);
nor U8965 (N_8965,N_5173,N_6003);
nand U8966 (N_8966,N_7477,N_5199);
nor U8967 (N_8967,N_6298,N_7258);
or U8968 (N_8968,N_6872,N_7459);
xor U8969 (N_8969,N_7490,N_5527);
and U8970 (N_8970,N_6141,N_5713);
or U8971 (N_8971,N_6373,N_6243);
or U8972 (N_8972,N_6936,N_7465);
and U8973 (N_8973,N_7342,N_6436);
nand U8974 (N_8974,N_6729,N_6827);
nand U8975 (N_8975,N_5603,N_5534);
or U8976 (N_8976,N_6966,N_7341);
and U8977 (N_8977,N_5525,N_6553);
nor U8978 (N_8978,N_6656,N_7351);
and U8979 (N_8979,N_6535,N_5269);
xnor U8980 (N_8980,N_6695,N_5764);
xnor U8981 (N_8981,N_7230,N_6164);
xor U8982 (N_8982,N_6217,N_6241);
and U8983 (N_8983,N_7390,N_5538);
xor U8984 (N_8984,N_6331,N_5168);
or U8985 (N_8985,N_5140,N_5366);
xor U8986 (N_8986,N_6218,N_6543);
nor U8987 (N_8987,N_6718,N_6823);
xor U8988 (N_8988,N_6688,N_6779);
nor U8989 (N_8989,N_5837,N_6832);
nand U8990 (N_8990,N_5813,N_6021);
and U8991 (N_8991,N_6943,N_7454);
nand U8992 (N_8992,N_6232,N_7155);
and U8993 (N_8993,N_6059,N_6911);
and U8994 (N_8994,N_5715,N_7220);
or U8995 (N_8995,N_6837,N_7432);
nor U8996 (N_8996,N_5276,N_6072);
xnor U8997 (N_8997,N_5150,N_6697);
nor U8998 (N_8998,N_6936,N_5515);
nor U8999 (N_8999,N_6511,N_5411);
nor U9000 (N_9000,N_6832,N_7065);
nand U9001 (N_9001,N_5329,N_6938);
nor U9002 (N_9002,N_6537,N_7248);
or U9003 (N_9003,N_7342,N_6030);
nor U9004 (N_9004,N_7304,N_6244);
xor U9005 (N_9005,N_6489,N_6959);
and U9006 (N_9006,N_6961,N_7319);
and U9007 (N_9007,N_6322,N_6422);
xor U9008 (N_9008,N_5449,N_7025);
nor U9009 (N_9009,N_6677,N_6585);
xnor U9010 (N_9010,N_7052,N_7499);
or U9011 (N_9011,N_6425,N_5376);
and U9012 (N_9012,N_6904,N_6857);
nand U9013 (N_9013,N_6641,N_7358);
nor U9014 (N_9014,N_5693,N_6370);
xor U9015 (N_9015,N_6527,N_5928);
nor U9016 (N_9016,N_7271,N_5325);
or U9017 (N_9017,N_5813,N_6796);
xor U9018 (N_9018,N_5984,N_7188);
xor U9019 (N_9019,N_7223,N_5707);
xnor U9020 (N_9020,N_5614,N_5756);
nor U9021 (N_9021,N_5960,N_6055);
nand U9022 (N_9022,N_5068,N_6379);
xor U9023 (N_9023,N_6859,N_5901);
and U9024 (N_9024,N_7215,N_7375);
or U9025 (N_9025,N_6725,N_6993);
and U9026 (N_9026,N_7203,N_6511);
and U9027 (N_9027,N_5284,N_6502);
and U9028 (N_9028,N_7455,N_7204);
or U9029 (N_9029,N_6422,N_5891);
xor U9030 (N_9030,N_5929,N_6753);
xor U9031 (N_9031,N_6347,N_6128);
and U9032 (N_9032,N_5323,N_6578);
or U9033 (N_9033,N_5666,N_5110);
or U9034 (N_9034,N_5106,N_6040);
or U9035 (N_9035,N_7042,N_5974);
or U9036 (N_9036,N_6372,N_7172);
nor U9037 (N_9037,N_7120,N_5150);
xor U9038 (N_9038,N_6847,N_7176);
xnor U9039 (N_9039,N_7453,N_5294);
nor U9040 (N_9040,N_5837,N_5824);
or U9041 (N_9041,N_6857,N_5540);
nor U9042 (N_9042,N_5244,N_5739);
nor U9043 (N_9043,N_5748,N_7496);
or U9044 (N_9044,N_5982,N_7213);
or U9045 (N_9045,N_6847,N_6455);
xnor U9046 (N_9046,N_7084,N_5238);
and U9047 (N_9047,N_5689,N_5302);
nor U9048 (N_9048,N_5752,N_6043);
or U9049 (N_9049,N_6778,N_6549);
nand U9050 (N_9050,N_6594,N_6340);
or U9051 (N_9051,N_5029,N_5565);
or U9052 (N_9052,N_5937,N_6734);
and U9053 (N_9053,N_6851,N_6714);
nand U9054 (N_9054,N_5982,N_6451);
and U9055 (N_9055,N_5735,N_5385);
or U9056 (N_9056,N_6337,N_7047);
or U9057 (N_9057,N_6959,N_5723);
nor U9058 (N_9058,N_5137,N_6956);
xnor U9059 (N_9059,N_6208,N_5936);
and U9060 (N_9060,N_6031,N_6068);
or U9061 (N_9061,N_5929,N_5622);
or U9062 (N_9062,N_6865,N_5021);
nor U9063 (N_9063,N_6373,N_7226);
xor U9064 (N_9064,N_6046,N_5502);
nor U9065 (N_9065,N_5033,N_5745);
nor U9066 (N_9066,N_7310,N_6539);
xor U9067 (N_9067,N_6477,N_6938);
nand U9068 (N_9068,N_5842,N_5537);
nor U9069 (N_9069,N_6735,N_7454);
and U9070 (N_9070,N_6814,N_5489);
or U9071 (N_9071,N_5547,N_6088);
nor U9072 (N_9072,N_7436,N_6598);
nor U9073 (N_9073,N_6812,N_5476);
nor U9074 (N_9074,N_5200,N_6901);
or U9075 (N_9075,N_6828,N_6942);
nor U9076 (N_9076,N_5229,N_5583);
and U9077 (N_9077,N_6831,N_7445);
nand U9078 (N_9078,N_7228,N_6524);
nor U9079 (N_9079,N_5039,N_5060);
nand U9080 (N_9080,N_6128,N_5417);
nor U9081 (N_9081,N_7104,N_6529);
nand U9082 (N_9082,N_7319,N_5539);
and U9083 (N_9083,N_6238,N_5884);
and U9084 (N_9084,N_6041,N_5975);
and U9085 (N_9085,N_6684,N_5267);
nand U9086 (N_9086,N_6967,N_6325);
nor U9087 (N_9087,N_5489,N_5928);
nor U9088 (N_9088,N_7318,N_6187);
or U9089 (N_9089,N_6406,N_6216);
xor U9090 (N_9090,N_5328,N_5195);
xor U9091 (N_9091,N_7091,N_6847);
xnor U9092 (N_9092,N_7182,N_7288);
xor U9093 (N_9093,N_5113,N_5602);
xnor U9094 (N_9094,N_6917,N_7138);
xnor U9095 (N_9095,N_5559,N_6125);
nor U9096 (N_9096,N_5156,N_5974);
nand U9097 (N_9097,N_7441,N_6195);
xnor U9098 (N_9098,N_5831,N_6014);
nor U9099 (N_9099,N_7205,N_5703);
xor U9100 (N_9100,N_6067,N_5787);
xor U9101 (N_9101,N_5507,N_5729);
or U9102 (N_9102,N_7438,N_5285);
nor U9103 (N_9103,N_7261,N_7473);
nand U9104 (N_9104,N_5015,N_6750);
or U9105 (N_9105,N_6598,N_6407);
xor U9106 (N_9106,N_6493,N_5023);
xnor U9107 (N_9107,N_6924,N_5456);
nand U9108 (N_9108,N_6897,N_5547);
nor U9109 (N_9109,N_5419,N_5873);
xnor U9110 (N_9110,N_6933,N_6785);
and U9111 (N_9111,N_6482,N_5614);
nand U9112 (N_9112,N_7093,N_5056);
or U9113 (N_9113,N_6398,N_5016);
or U9114 (N_9114,N_7239,N_5130);
nor U9115 (N_9115,N_6349,N_5614);
or U9116 (N_9116,N_6211,N_7047);
nand U9117 (N_9117,N_6280,N_7017);
nor U9118 (N_9118,N_5138,N_6634);
nor U9119 (N_9119,N_7472,N_7057);
or U9120 (N_9120,N_7380,N_5875);
nand U9121 (N_9121,N_7004,N_5659);
nor U9122 (N_9122,N_6519,N_7001);
or U9123 (N_9123,N_7360,N_5670);
or U9124 (N_9124,N_7239,N_6127);
xor U9125 (N_9125,N_6202,N_5973);
xnor U9126 (N_9126,N_7204,N_6959);
nor U9127 (N_9127,N_6559,N_5951);
or U9128 (N_9128,N_5261,N_6896);
nand U9129 (N_9129,N_6016,N_5731);
nand U9130 (N_9130,N_6832,N_7459);
and U9131 (N_9131,N_6912,N_5143);
xor U9132 (N_9132,N_5155,N_7117);
nand U9133 (N_9133,N_7089,N_5470);
or U9134 (N_9134,N_6129,N_6854);
or U9135 (N_9135,N_5415,N_5771);
or U9136 (N_9136,N_5245,N_6065);
nand U9137 (N_9137,N_5450,N_5162);
or U9138 (N_9138,N_6744,N_5292);
nand U9139 (N_9139,N_6937,N_6205);
and U9140 (N_9140,N_7171,N_6701);
xnor U9141 (N_9141,N_5485,N_7473);
nor U9142 (N_9142,N_5027,N_5114);
and U9143 (N_9143,N_6263,N_5897);
xor U9144 (N_9144,N_7067,N_5008);
and U9145 (N_9145,N_7498,N_5090);
and U9146 (N_9146,N_5628,N_6306);
or U9147 (N_9147,N_6590,N_7036);
or U9148 (N_9148,N_6741,N_5149);
and U9149 (N_9149,N_7090,N_6684);
nand U9150 (N_9150,N_5327,N_6418);
or U9151 (N_9151,N_5815,N_5446);
xnor U9152 (N_9152,N_6388,N_5933);
nor U9153 (N_9153,N_5032,N_7444);
xor U9154 (N_9154,N_5637,N_6250);
xor U9155 (N_9155,N_7175,N_5033);
and U9156 (N_9156,N_7158,N_6828);
xnor U9157 (N_9157,N_7272,N_6137);
nor U9158 (N_9158,N_6035,N_5585);
or U9159 (N_9159,N_7334,N_6390);
or U9160 (N_9160,N_5619,N_5446);
nor U9161 (N_9161,N_5767,N_5607);
or U9162 (N_9162,N_5427,N_5999);
and U9163 (N_9163,N_7383,N_6604);
xnor U9164 (N_9164,N_6207,N_7013);
nor U9165 (N_9165,N_6596,N_5317);
nor U9166 (N_9166,N_5330,N_7441);
nand U9167 (N_9167,N_5136,N_6635);
and U9168 (N_9168,N_6568,N_6524);
nand U9169 (N_9169,N_7067,N_5375);
nor U9170 (N_9170,N_7030,N_5444);
nor U9171 (N_9171,N_6931,N_5009);
and U9172 (N_9172,N_6087,N_7101);
and U9173 (N_9173,N_6265,N_5816);
and U9174 (N_9174,N_5184,N_5749);
and U9175 (N_9175,N_5413,N_6436);
and U9176 (N_9176,N_5154,N_6673);
xor U9177 (N_9177,N_7177,N_6116);
or U9178 (N_9178,N_5144,N_5023);
xor U9179 (N_9179,N_6400,N_5434);
and U9180 (N_9180,N_7422,N_7444);
xor U9181 (N_9181,N_6534,N_7319);
xor U9182 (N_9182,N_6291,N_6981);
nor U9183 (N_9183,N_6850,N_5885);
and U9184 (N_9184,N_6529,N_6149);
nand U9185 (N_9185,N_5233,N_5764);
xor U9186 (N_9186,N_5330,N_7052);
and U9187 (N_9187,N_6860,N_5502);
or U9188 (N_9188,N_6001,N_6543);
and U9189 (N_9189,N_5841,N_5991);
nand U9190 (N_9190,N_6816,N_5839);
nand U9191 (N_9191,N_5783,N_7034);
nor U9192 (N_9192,N_6965,N_5688);
and U9193 (N_9193,N_5039,N_6025);
xnor U9194 (N_9194,N_5011,N_6054);
xnor U9195 (N_9195,N_6213,N_5692);
and U9196 (N_9196,N_5511,N_7204);
and U9197 (N_9197,N_5716,N_6532);
and U9198 (N_9198,N_5251,N_5455);
nand U9199 (N_9199,N_5405,N_5808);
nand U9200 (N_9200,N_6782,N_5254);
nor U9201 (N_9201,N_7453,N_5252);
nand U9202 (N_9202,N_7246,N_6499);
or U9203 (N_9203,N_5570,N_6994);
xor U9204 (N_9204,N_6570,N_5256);
nor U9205 (N_9205,N_7061,N_6837);
xor U9206 (N_9206,N_5931,N_6770);
nand U9207 (N_9207,N_5331,N_5822);
nand U9208 (N_9208,N_5957,N_6862);
or U9209 (N_9209,N_5814,N_5433);
nand U9210 (N_9210,N_6123,N_5417);
or U9211 (N_9211,N_6822,N_5913);
and U9212 (N_9212,N_6722,N_5568);
nand U9213 (N_9213,N_6882,N_5726);
and U9214 (N_9214,N_6235,N_7435);
or U9215 (N_9215,N_7105,N_6522);
and U9216 (N_9216,N_5380,N_5196);
and U9217 (N_9217,N_6572,N_5771);
or U9218 (N_9218,N_5149,N_6532);
or U9219 (N_9219,N_5032,N_7348);
or U9220 (N_9220,N_5371,N_6428);
or U9221 (N_9221,N_7356,N_7282);
nand U9222 (N_9222,N_5533,N_6521);
or U9223 (N_9223,N_7072,N_5258);
or U9224 (N_9224,N_7184,N_6600);
xnor U9225 (N_9225,N_6094,N_6174);
and U9226 (N_9226,N_6769,N_7479);
xnor U9227 (N_9227,N_6478,N_6226);
nand U9228 (N_9228,N_6439,N_6706);
xnor U9229 (N_9229,N_6291,N_7434);
nand U9230 (N_9230,N_7308,N_6935);
xnor U9231 (N_9231,N_6723,N_5431);
and U9232 (N_9232,N_6656,N_6737);
nor U9233 (N_9233,N_6675,N_6034);
and U9234 (N_9234,N_7152,N_7197);
xnor U9235 (N_9235,N_7322,N_7429);
or U9236 (N_9236,N_5649,N_5333);
or U9237 (N_9237,N_6081,N_6127);
or U9238 (N_9238,N_5565,N_6611);
or U9239 (N_9239,N_5413,N_6768);
nand U9240 (N_9240,N_6744,N_6122);
xor U9241 (N_9241,N_6964,N_6132);
nand U9242 (N_9242,N_5778,N_5897);
xor U9243 (N_9243,N_7105,N_5545);
or U9244 (N_9244,N_6543,N_5888);
nor U9245 (N_9245,N_5401,N_7098);
nor U9246 (N_9246,N_7284,N_6453);
nand U9247 (N_9247,N_6518,N_7480);
and U9248 (N_9248,N_5765,N_5706);
nand U9249 (N_9249,N_7450,N_5234);
or U9250 (N_9250,N_5176,N_7315);
or U9251 (N_9251,N_5064,N_5014);
nor U9252 (N_9252,N_7101,N_5358);
or U9253 (N_9253,N_5168,N_5847);
nor U9254 (N_9254,N_6363,N_6490);
and U9255 (N_9255,N_5054,N_6608);
or U9256 (N_9256,N_5344,N_6922);
or U9257 (N_9257,N_5378,N_5833);
nor U9258 (N_9258,N_6375,N_5725);
or U9259 (N_9259,N_6503,N_6372);
xor U9260 (N_9260,N_6470,N_5397);
nor U9261 (N_9261,N_5187,N_6706);
and U9262 (N_9262,N_5714,N_5411);
nand U9263 (N_9263,N_6948,N_6425);
nand U9264 (N_9264,N_7468,N_7466);
xor U9265 (N_9265,N_6335,N_7432);
nor U9266 (N_9266,N_7379,N_6358);
and U9267 (N_9267,N_5145,N_6893);
or U9268 (N_9268,N_5284,N_5050);
xor U9269 (N_9269,N_7483,N_6083);
nand U9270 (N_9270,N_5032,N_7229);
and U9271 (N_9271,N_5947,N_6921);
and U9272 (N_9272,N_6317,N_5517);
or U9273 (N_9273,N_5523,N_7466);
nor U9274 (N_9274,N_6123,N_6682);
xor U9275 (N_9275,N_6199,N_5540);
nor U9276 (N_9276,N_6970,N_6057);
and U9277 (N_9277,N_6994,N_7067);
nor U9278 (N_9278,N_6917,N_5809);
nand U9279 (N_9279,N_6893,N_5128);
xnor U9280 (N_9280,N_6869,N_5424);
and U9281 (N_9281,N_6296,N_7238);
xnor U9282 (N_9282,N_5057,N_5545);
xor U9283 (N_9283,N_6137,N_7193);
nand U9284 (N_9284,N_6675,N_6776);
and U9285 (N_9285,N_5186,N_6023);
nor U9286 (N_9286,N_6135,N_5801);
xor U9287 (N_9287,N_5145,N_6038);
or U9288 (N_9288,N_5187,N_6902);
or U9289 (N_9289,N_6662,N_5001);
and U9290 (N_9290,N_5426,N_6348);
and U9291 (N_9291,N_6433,N_5103);
and U9292 (N_9292,N_5029,N_6798);
nor U9293 (N_9293,N_5820,N_7217);
xnor U9294 (N_9294,N_5250,N_7468);
and U9295 (N_9295,N_5581,N_7099);
nand U9296 (N_9296,N_7000,N_6402);
nand U9297 (N_9297,N_6252,N_6231);
or U9298 (N_9298,N_5032,N_5822);
nor U9299 (N_9299,N_6528,N_6377);
nor U9300 (N_9300,N_5515,N_5004);
xor U9301 (N_9301,N_5380,N_6966);
nor U9302 (N_9302,N_7455,N_6715);
or U9303 (N_9303,N_7215,N_5332);
xor U9304 (N_9304,N_6242,N_7414);
nand U9305 (N_9305,N_5552,N_5314);
nor U9306 (N_9306,N_7015,N_6696);
or U9307 (N_9307,N_6450,N_7295);
or U9308 (N_9308,N_6245,N_7111);
or U9309 (N_9309,N_6798,N_6449);
or U9310 (N_9310,N_5806,N_6189);
nand U9311 (N_9311,N_6110,N_5551);
or U9312 (N_9312,N_6442,N_5290);
or U9313 (N_9313,N_7473,N_6136);
xor U9314 (N_9314,N_5046,N_6896);
or U9315 (N_9315,N_7007,N_5380);
or U9316 (N_9316,N_7281,N_7421);
or U9317 (N_9317,N_5332,N_6067);
nor U9318 (N_9318,N_7364,N_6728);
nor U9319 (N_9319,N_6421,N_6481);
and U9320 (N_9320,N_5852,N_6389);
and U9321 (N_9321,N_5752,N_6199);
nor U9322 (N_9322,N_6694,N_5910);
nand U9323 (N_9323,N_5243,N_5571);
xor U9324 (N_9324,N_6395,N_6263);
or U9325 (N_9325,N_7065,N_5590);
xor U9326 (N_9326,N_6014,N_5979);
and U9327 (N_9327,N_6555,N_6189);
xor U9328 (N_9328,N_6414,N_6668);
nand U9329 (N_9329,N_7031,N_5557);
nor U9330 (N_9330,N_6731,N_6932);
or U9331 (N_9331,N_7085,N_6401);
nand U9332 (N_9332,N_6931,N_7442);
or U9333 (N_9333,N_6140,N_6932);
or U9334 (N_9334,N_6477,N_6464);
nor U9335 (N_9335,N_6769,N_6601);
nor U9336 (N_9336,N_6756,N_5372);
xor U9337 (N_9337,N_6465,N_5633);
or U9338 (N_9338,N_6481,N_6094);
nand U9339 (N_9339,N_6094,N_5976);
nand U9340 (N_9340,N_6917,N_5796);
or U9341 (N_9341,N_7257,N_7161);
or U9342 (N_9342,N_6560,N_5436);
nor U9343 (N_9343,N_6377,N_6889);
nor U9344 (N_9344,N_6845,N_6765);
or U9345 (N_9345,N_7310,N_6714);
nand U9346 (N_9346,N_6164,N_6703);
and U9347 (N_9347,N_6931,N_6250);
nand U9348 (N_9348,N_5038,N_7249);
nor U9349 (N_9349,N_7030,N_5120);
nor U9350 (N_9350,N_6560,N_6524);
nand U9351 (N_9351,N_5580,N_5349);
nor U9352 (N_9352,N_5966,N_5583);
nand U9353 (N_9353,N_6317,N_5121);
xnor U9354 (N_9354,N_7169,N_6318);
and U9355 (N_9355,N_5924,N_6014);
nand U9356 (N_9356,N_7016,N_6295);
or U9357 (N_9357,N_5102,N_6217);
nor U9358 (N_9358,N_6459,N_6279);
xnor U9359 (N_9359,N_7176,N_5592);
nor U9360 (N_9360,N_6729,N_6882);
nand U9361 (N_9361,N_6390,N_5804);
nand U9362 (N_9362,N_6433,N_6203);
nand U9363 (N_9363,N_7305,N_7471);
xnor U9364 (N_9364,N_5945,N_6400);
nand U9365 (N_9365,N_6338,N_5171);
nand U9366 (N_9366,N_5579,N_6964);
xor U9367 (N_9367,N_6217,N_6964);
or U9368 (N_9368,N_5251,N_7002);
or U9369 (N_9369,N_6222,N_6874);
nand U9370 (N_9370,N_5259,N_7373);
nor U9371 (N_9371,N_5257,N_5124);
xnor U9372 (N_9372,N_6046,N_7223);
nand U9373 (N_9373,N_5063,N_5754);
and U9374 (N_9374,N_5282,N_6369);
xnor U9375 (N_9375,N_7183,N_6090);
nand U9376 (N_9376,N_7394,N_5827);
xor U9377 (N_9377,N_5185,N_5691);
or U9378 (N_9378,N_6208,N_7487);
nor U9379 (N_9379,N_6354,N_5671);
nand U9380 (N_9380,N_6849,N_5098);
nor U9381 (N_9381,N_7221,N_5412);
xnor U9382 (N_9382,N_5119,N_6800);
nand U9383 (N_9383,N_5530,N_6001);
nand U9384 (N_9384,N_6664,N_5978);
nor U9385 (N_9385,N_5200,N_5680);
and U9386 (N_9386,N_5910,N_6316);
or U9387 (N_9387,N_5134,N_6803);
and U9388 (N_9388,N_5333,N_6270);
nor U9389 (N_9389,N_5403,N_6577);
xor U9390 (N_9390,N_7201,N_6745);
nor U9391 (N_9391,N_6885,N_5628);
or U9392 (N_9392,N_6765,N_7300);
xor U9393 (N_9393,N_7402,N_5140);
nor U9394 (N_9394,N_6271,N_5340);
xor U9395 (N_9395,N_7294,N_6232);
xor U9396 (N_9396,N_7174,N_6475);
nor U9397 (N_9397,N_6204,N_6700);
and U9398 (N_9398,N_5633,N_5782);
xnor U9399 (N_9399,N_7269,N_5100);
and U9400 (N_9400,N_6338,N_7126);
or U9401 (N_9401,N_7116,N_5680);
and U9402 (N_9402,N_5196,N_5847);
or U9403 (N_9403,N_5912,N_6399);
nor U9404 (N_9404,N_5457,N_6076);
xor U9405 (N_9405,N_6775,N_5642);
or U9406 (N_9406,N_6135,N_5423);
or U9407 (N_9407,N_5224,N_6560);
nor U9408 (N_9408,N_6006,N_7288);
xnor U9409 (N_9409,N_7275,N_6499);
nand U9410 (N_9410,N_5689,N_6012);
or U9411 (N_9411,N_6818,N_6926);
nand U9412 (N_9412,N_5998,N_6386);
and U9413 (N_9413,N_5178,N_5849);
xnor U9414 (N_9414,N_5122,N_5428);
xnor U9415 (N_9415,N_6372,N_7282);
nand U9416 (N_9416,N_5124,N_6621);
xnor U9417 (N_9417,N_6207,N_5736);
and U9418 (N_9418,N_5945,N_5917);
xor U9419 (N_9419,N_7337,N_5828);
nor U9420 (N_9420,N_6300,N_5259);
nand U9421 (N_9421,N_5046,N_6962);
nand U9422 (N_9422,N_5472,N_5405);
and U9423 (N_9423,N_5927,N_7038);
or U9424 (N_9424,N_5707,N_5842);
xnor U9425 (N_9425,N_6281,N_5401);
nor U9426 (N_9426,N_5089,N_7148);
xor U9427 (N_9427,N_7369,N_5722);
or U9428 (N_9428,N_6180,N_6005);
and U9429 (N_9429,N_5053,N_5713);
or U9430 (N_9430,N_5622,N_6656);
and U9431 (N_9431,N_6055,N_6378);
xnor U9432 (N_9432,N_6353,N_6848);
nor U9433 (N_9433,N_6064,N_6473);
and U9434 (N_9434,N_5691,N_7070);
nor U9435 (N_9435,N_5960,N_5051);
or U9436 (N_9436,N_6717,N_6012);
or U9437 (N_9437,N_6876,N_5111);
and U9438 (N_9438,N_5275,N_6419);
nor U9439 (N_9439,N_6671,N_5376);
nand U9440 (N_9440,N_5514,N_5901);
and U9441 (N_9441,N_5539,N_6072);
xnor U9442 (N_9442,N_5801,N_5539);
xor U9443 (N_9443,N_5806,N_6898);
nand U9444 (N_9444,N_6924,N_5573);
xnor U9445 (N_9445,N_5238,N_5652);
or U9446 (N_9446,N_6391,N_5958);
or U9447 (N_9447,N_5799,N_5759);
and U9448 (N_9448,N_6238,N_5876);
and U9449 (N_9449,N_6047,N_5260);
and U9450 (N_9450,N_6752,N_6261);
nor U9451 (N_9451,N_5201,N_5552);
or U9452 (N_9452,N_6147,N_5903);
nand U9453 (N_9453,N_6364,N_6225);
xor U9454 (N_9454,N_7317,N_7139);
or U9455 (N_9455,N_6084,N_6623);
and U9456 (N_9456,N_5155,N_5620);
or U9457 (N_9457,N_5918,N_6294);
and U9458 (N_9458,N_5417,N_6223);
xor U9459 (N_9459,N_6186,N_5299);
xor U9460 (N_9460,N_5617,N_6705);
and U9461 (N_9461,N_6387,N_5803);
or U9462 (N_9462,N_6466,N_5580);
or U9463 (N_9463,N_5933,N_5425);
or U9464 (N_9464,N_6753,N_6646);
nor U9465 (N_9465,N_6522,N_7491);
or U9466 (N_9466,N_7296,N_5096);
nand U9467 (N_9467,N_5988,N_5780);
nand U9468 (N_9468,N_5636,N_6561);
nand U9469 (N_9469,N_5899,N_5950);
or U9470 (N_9470,N_7417,N_7283);
nor U9471 (N_9471,N_6939,N_7337);
nor U9472 (N_9472,N_6863,N_5904);
nand U9473 (N_9473,N_6949,N_6856);
nor U9474 (N_9474,N_6575,N_7315);
xnor U9475 (N_9475,N_7302,N_6643);
nand U9476 (N_9476,N_6831,N_6307);
nor U9477 (N_9477,N_6643,N_5793);
or U9478 (N_9478,N_6011,N_5752);
or U9479 (N_9479,N_5498,N_7049);
nor U9480 (N_9480,N_6493,N_5002);
or U9481 (N_9481,N_5863,N_6863);
nand U9482 (N_9482,N_6027,N_6798);
nor U9483 (N_9483,N_7414,N_6103);
nor U9484 (N_9484,N_6642,N_7401);
or U9485 (N_9485,N_7094,N_6395);
nor U9486 (N_9486,N_5614,N_5961);
nand U9487 (N_9487,N_5532,N_6469);
nand U9488 (N_9488,N_5870,N_5582);
or U9489 (N_9489,N_6030,N_7269);
xnor U9490 (N_9490,N_7106,N_6859);
nand U9491 (N_9491,N_5923,N_7336);
xor U9492 (N_9492,N_5095,N_5558);
nand U9493 (N_9493,N_7138,N_6850);
nor U9494 (N_9494,N_6688,N_6431);
nor U9495 (N_9495,N_5778,N_6454);
xor U9496 (N_9496,N_6288,N_5028);
nand U9497 (N_9497,N_7427,N_7238);
nor U9498 (N_9498,N_7069,N_6154);
xnor U9499 (N_9499,N_5560,N_5227);
and U9500 (N_9500,N_6469,N_6240);
nand U9501 (N_9501,N_5048,N_6203);
nand U9502 (N_9502,N_7158,N_6772);
nand U9503 (N_9503,N_5980,N_5249);
xnor U9504 (N_9504,N_5819,N_7407);
or U9505 (N_9505,N_5634,N_6978);
xor U9506 (N_9506,N_6016,N_6861);
or U9507 (N_9507,N_5245,N_6746);
nor U9508 (N_9508,N_5861,N_7144);
nor U9509 (N_9509,N_5677,N_7287);
nand U9510 (N_9510,N_5587,N_5596);
or U9511 (N_9511,N_6866,N_5864);
xnor U9512 (N_9512,N_6473,N_5390);
nor U9513 (N_9513,N_5358,N_7078);
or U9514 (N_9514,N_5025,N_6118);
nand U9515 (N_9515,N_5403,N_5657);
nand U9516 (N_9516,N_5358,N_7055);
and U9517 (N_9517,N_6364,N_6846);
and U9518 (N_9518,N_5910,N_6118);
xor U9519 (N_9519,N_5737,N_6261);
nor U9520 (N_9520,N_5582,N_6499);
nand U9521 (N_9521,N_5578,N_7124);
nor U9522 (N_9522,N_5792,N_5923);
nor U9523 (N_9523,N_7264,N_5722);
and U9524 (N_9524,N_6910,N_5785);
or U9525 (N_9525,N_5071,N_6024);
nor U9526 (N_9526,N_7340,N_6519);
nand U9527 (N_9527,N_5952,N_6492);
nor U9528 (N_9528,N_5190,N_6426);
and U9529 (N_9529,N_5739,N_6946);
nor U9530 (N_9530,N_6158,N_5519);
nor U9531 (N_9531,N_5695,N_6891);
and U9532 (N_9532,N_6521,N_5734);
and U9533 (N_9533,N_5428,N_5846);
nand U9534 (N_9534,N_6524,N_5389);
nor U9535 (N_9535,N_6462,N_6576);
or U9536 (N_9536,N_6725,N_6611);
and U9537 (N_9537,N_5597,N_5544);
and U9538 (N_9538,N_7268,N_6096);
nand U9539 (N_9539,N_6992,N_5924);
nor U9540 (N_9540,N_7228,N_5207);
nand U9541 (N_9541,N_6855,N_6873);
nor U9542 (N_9542,N_6629,N_5000);
xnor U9543 (N_9543,N_6806,N_6631);
nor U9544 (N_9544,N_5699,N_6038);
nand U9545 (N_9545,N_5451,N_5441);
xor U9546 (N_9546,N_5587,N_5493);
and U9547 (N_9547,N_6743,N_7244);
xnor U9548 (N_9548,N_5092,N_5261);
xnor U9549 (N_9549,N_5081,N_7313);
nor U9550 (N_9550,N_6656,N_5613);
xnor U9551 (N_9551,N_6703,N_6717);
or U9552 (N_9552,N_5704,N_5247);
nand U9553 (N_9553,N_5407,N_7067);
xnor U9554 (N_9554,N_6929,N_6763);
nor U9555 (N_9555,N_5190,N_5502);
or U9556 (N_9556,N_6853,N_6483);
nor U9557 (N_9557,N_5231,N_5651);
and U9558 (N_9558,N_7179,N_5061);
xnor U9559 (N_9559,N_6407,N_7483);
nand U9560 (N_9560,N_6671,N_6821);
or U9561 (N_9561,N_5517,N_5228);
or U9562 (N_9562,N_5318,N_5898);
or U9563 (N_9563,N_7202,N_6052);
nand U9564 (N_9564,N_6756,N_5157);
or U9565 (N_9565,N_7317,N_5903);
xor U9566 (N_9566,N_5089,N_7421);
xor U9567 (N_9567,N_7461,N_6465);
xor U9568 (N_9568,N_6044,N_7261);
and U9569 (N_9569,N_5775,N_6626);
xor U9570 (N_9570,N_5297,N_5891);
or U9571 (N_9571,N_6113,N_6953);
xor U9572 (N_9572,N_5613,N_6429);
nand U9573 (N_9573,N_6095,N_5165);
nand U9574 (N_9574,N_5264,N_5980);
xor U9575 (N_9575,N_6876,N_6717);
and U9576 (N_9576,N_6382,N_7488);
nand U9577 (N_9577,N_6251,N_7297);
nand U9578 (N_9578,N_6061,N_5498);
nor U9579 (N_9579,N_5781,N_5668);
and U9580 (N_9580,N_5854,N_5317);
nand U9581 (N_9581,N_7047,N_6464);
xnor U9582 (N_9582,N_5418,N_6916);
nor U9583 (N_9583,N_7033,N_5245);
xnor U9584 (N_9584,N_5241,N_6808);
xnor U9585 (N_9585,N_7245,N_7371);
nor U9586 (N_9586,N_6261,N_6281);
or U9587 (N_9587,N_5090,N_5621);
nor U9588 (N_9588,N_7456,N_5651);
nand U9589 (N_9589,N_6960,N_5160);
xnor U9590 (N_9590,N_7464,N_5591);
nor U9591 (N_9591,N_5381,N_7171);
nor U9592 (N_9592,N_6156,N_5151);
and U9593 (N_9593,N_5897,N_5692);
nand U9594 (N_9594,N_5430,N_6578);
xor U9595 (N_9595,N_6391,N_5808);
nand U9596 (N_9596,N_5970,N_5709);
or U9597 (N_9597,N_5217,N_6632);
nand U9598 (N_9598,N_6266,N_6207);
nor U9599 (N_9599,N_7422,N_5345);
or U9600 (N_9600,N_6421,N_5409);
nor U9601 (N_9601,N_5963,N_5964);
or U9602 (N_9602,N_6941,N_5547);
nand U9603 (N_9603,N_6510,N_5681);
or U9604 (N_9604,N_6604,N_5528);
and U9605 (N_9605,N_5127,N_6026);
xnor U9606 (N_9606,N_7497,N_7120);
nor U9607 (N_9607,N_6760,N_5979);
and U9608 (N_9608,N_6938,N_5589);
and U9609 (N_9609,N_7271,N_6861);
xor U9610 (N_9610,N_6869,N_7221);
nor U9611 (N_9611,N_6167,N_6516);
and U9612 (N_9612,N_6456,N_7072);
nand U9613 (N_9613,N_5181,N_6815);
nand U9614 (N_9614,N_6002,N_5254);
nand U9615 (N_9615,N_6449,N_6116);
nand U9616 (N_9616,N_5444,N_5957);
nor U9617 (N_9617,N_7441,N_7306);
or U9618 (N_9618,N_5500,N_5407);
xnor U9619 (N_9619,N_7338,N_6333);
xnor U9620 (N_9620,N_6191,N_6767);
and U9621 (N_9621,N_6167,N_7289);
and U9622 (N_9622,N_7409,N_5941);
nor U9623 (N_9623,N_5236,N_6246);
nor U9624 (N_9624,N_5219,N_6537);
nor U9625 (N_9625,N_6503,N_5672);
nor U9626 (N_9626,N_5984,N_5702);
nand U9627 (N_9627,N_5653,N_5372);
nand U9628 (N_9628,N_6564,N_6086);
nor U9629 (N_9629,N_6901,N_7069);
or U9630 (N_9630,N_5912,N_5686);
xnor U9631 (N_9631,N_5761,N_6673);
and U9632 (N_9632,N_7117,N_7027);
nand U9633 (N_9633,N_5390,N_6205);
nor U9634 (N_9634,N_7111,N_6882);
nand U9635 (N_9635,N_7280,N_5912);
nand U9636 (N_9636,N_6222,N_7244);
xor U9637 (N_9637,N_7377,N_7265);
nor U9638 (N_9638,N_7471,N_5492);
nand U9639 (N_9639,N_5630,N_5270);
nand U9640 (N_9640,N_6968,N_5640);
or U9641 (N_9641,N_5829,N_6386);
xor U9642 (N_9642,N_5888,N_7166);
or U9643 (N_9643,N_5297,N_6381);
xnor U9644 (N_9644,N_7255,N_6198);
or U9645 (N_9645,N_7424,N_7315);
nor U9646 (N_9646,N_6968,N_5672);
nor U9647 (N_9647,N_5408,N_6452);
xnor U9648 (N_9648,N_6726,N_6312);
and U9649 (N_9649,N_6818,N_6385);
xnor U9650 (N_9650,N_6192,N_6639);
and U9651 (N_9651,N_5249,N_6763);
nor U9652 (N_9652,N_5877,N_6264);
xnor U9653 (N_9653,N_6144,N_6944);
and U9654 (N_9654,N_5563,N_7352);
nand U9655 (N_9655,N_6547,N_6654);
nand U9656 (N_9656,N_5567,N_5233);
and U9657 (N_9657,N_5009,N_6493);
nand U9658 (N_9658,N_6676,N_6034);
nor U9659 (N_9659,N_7355,N_7158);
nor U9660 (N_9660,N_5825,N_5739);
and U9661 (N_9661,N_5172,N_6856);
nor U9662 (N_9662,N_7091,N_5957);
xor U9663 (N_9663,N_5569,N_5700);
nand U9664 (N_9664,N_6887,N_7365);
nand U9665 (N_9665,N_5796,N_5524);
or U9666 (N_9666,N_5214,N_7194);
nand U9667 (N_9667,N_7272,N_5156);
nor U9668 (N_9668,N_5751,N_5572);
nand U9669 (N_9669,N_5303,N_5640);
nand U9670 (N_9670,N_5442,N_5206);
nor U9671 (N_9671,N_6048,N_6606);
and U9672 (N_9672,N_5224,N_5038);
nor U9673 (N_9673,N_5345,N_7094);
or U9674 (N_9674,N_5807,N_6626);
xor U9675 (N_9675,N_5685,N_6189);
xnor U9676 (N_9676,N_6794,N_6907);
nand U9677 (N_9677,N_6458,N_6400);
or U9678 (N_9678,N_5062,N_6044);
and U9679 (N_9679,N_5609,N_5125);
or U9680 (N_9680,N_7130,N_5167);
nor U9681 (N_9681,N_6141,N_5196);
and U9682 (N_9682,N_6813,N_7491);
nand U9683 (N_9683,N_6257,N_5833);
and U9684 (N_9684,N_5955,N_7175);
xor U9685 (N_9685,N_5710,N_5935);
and U9686 (N_9686,N_7309,N_6434);
xnor U9687 (N_9687,N_5479,N_7065);
nor U9688 (N_9688,N_5386,N_6012);
nand U9689 (N_9689,N_7495,N_5852);
nor U9690 (N_9690,N_7226,N_7409);
nor U9691 (N_9691,N_6761,N_6963);
xor U9692 (N_9692,N_6137,N_7148);
and U9693 (N_9693,N_6995,N_6365);
or U9694 (N_9694,N_5717,N_7142);
nand U9695 (N_9695,N_6946,N_5605);
and U9696 (N_9696,N_5499,N_7419);
nand U9697 (N_9697,N_6723,N_6323);
or U9698 (N_9698,N_6876,N_6868);
xnor U9699 (N_9699,N_7215,N_6656);
xnor U9700 (N_9700,N_6167,N_5164);
or U9701 (N_9701,N_6858,N_5890);
nor U9702 (N_9702,N_5717,N_6178);
and U9703 (N_9703,N_5024,N_5430);
nand U9704 (N_9704,N_6877,N_5839);
xnor U9705 (N_9705,N_6352,N_5693);
xor U9706 (N_9706,N_5321,N_6413);
xnor U9707 (N_9707,N_6127,N_6365);
xnor U9708 (N_9708,N_7137,N_5277);
nand U9709 (N_9709,N_7272,N_7401);
nand U9710 (N_9710,N_6018,N_6985);
and U9711 (N_9711,N_6936,N_7079);
or U9712 (N_9712,N_7439,N_6712);
xnor U9713 (N_9713,N_6121,N_5404);
nand U9714 (N_9714,N_7186,N_5468);
nor U9715 (N_9715,N_6250,N_7443);
xnor U9716 (N_9716,N_7257,N_5331);
and U9717 (N_9717,N_6757,N_6139);
or U9718 (N_9718,N_5143,N_5282);
xnor U9719 (N_9719,N_6055,N_6031);
nand U9720 (N_9720,N_7062,N_5988);
and U9721 (N_9721,N_6605,N_5276);
nand U9722 (N_9722,N_6512,N_5514);
nand U9723 (N_9723,N_6890,N_6107);
nand U9724 (N_9724,N_5979,N_5592);
nor U9725 (N_9725,N_6704,N_7367);
nor U9726 (N_9726,N_5498,N_5337);
nor U9727 (N_9727,N_5391,N_7103);
nor U9728 (N_9728,N_5784,N_6725);
xor U9729 (N_9729,N_5654,N_5690);
and U9730 (N_9730,N_6008,N_6162);
or U9731 (N_9731,N_7427,N_5204);
nor U9732 (N_9732,N_7369,N_5331);
nand U9733 (N_9733,N_5160,N_6217);
nor U9734 (N_9734,N_5320,N_6899);
xnor U9735 (N_9735,N_6095,N_5364);
xor U9736 (N_9736,N_6659,N_5054);
or U9737 (N_9737,N_5866,N_5053);
and U9738 (N_9738,N_7387,N_5281);
nor U9739 (N_9739,N_7499,N_7108);
xnor U9740 (N_9740,N_6312,N_7089);
nor U9741 (N_9741,N_5525,N_5399);
nor U9742 (N_9742,N_6440,N_6943);
xnor U9743 (N_9743,N_6276,N_6629);
nand U9744 (N_9744,N_5913,N_6767);
nand U9745 (N_9745,N_7128,N_5925);
or U9746 (N_9746,N_5753,N_5576);
and U9747 (N_9747,N_5843,N_5001);
or U9748 (N_9748,N_5096,N_5303);
or U9749 (N_9749,N_5685,N_7301);
nand U9750 (N_9750,N_5213,N_7179);
nand U9751 (N_9751,N_5256,N_6010);
xor U9752 (N_9752,N_6476,N_7121);
nor U9753 (N_9753,N_6731,N_7371);
and U9754 (N_9754,N_5185,N_6259);
xor U9755 (N_9755,N_5206,N_5508);
nand U9756 (N_9756,N_6790,N_5152);
or U9757 (N_9757,N_5056,N_6947);
nor U9758 (N_9758,N_7166,N_5191);
or U9759 (N_9759,N_7386,N_5791);
or U9760 (N_9760,N_5823,N_6002);
nor U9761 (N_9761,N_5980,N_5203);
xor U9762 (N_9762,N_7119,N_6372);
and U9763 (N_9763,N_5879,N_5463);
xnor U9764 (N_9764,N_7422,N_7248);
and U9765 (N_9765,N_6048,N_6389);
and U9766 (N_9766,N_5183,N_7489);
and U9767 (N_9767,N_5294,N_7448);
xnor U9768 (N_9768,N_6862,N_6864);
nand U9769 (N_9769,N_7201,N_6953);
or U9770 (N_9770,N_5524,N_7412);
nor U9771 (N_9771,N_6546,N_7277);
or U9772 (N_9772,N_7279,N_6165);
xnor U9773 (N_9773,N_5929,N_7290);
and U9774 (N_9774,N_7221,N_5532);
nand U9775 (N_9775,N_7451,N_6192);
or U9776 (N_9776,N_6945,N_6243);
or U9777 (N_9777,N_7467,N_5123);
nand U9778 (N_9778,N_6247,N_6290);
nand U9779 (N_9779,N_6959,N_6125);
xor U9780 (N_9780,N_5754,N_6279);
nor U9781 (N_9781,N_5267,N_5016);
nand U9782 (N_9782,N_5478,N_6607);
nor U9783 (N_9783,N_6841,N_5661);
xor U9784 (N_9784,N_5637,N_5332);
nand U9785 (N_9785,N_6861,N_5061);
nand U9786 (N_9786,N_6278,N_7064);
nor U9787 (N_9787,N_6332,N_6123);
xnor U9788 (N_9788,N_6079,N_7446);
nand U9789 (N_9789,N_6136,N_6309);
or U9790 (N_9790,N_6394,N_5624);
nand U9791 (N_9791,N_6023,N_6025);
nor U9792 (N_9792,N_5533,N_5021);
nor U9793 (N_9793,N_7366,N_6726);
xnor U9794 (N_9794,N_7037,N_5688);
xor U9795 (N_9795,N_7113,N_6550);
nor U9796 (N_9796,N_7329,N_5603);
nand U9797 (N_9797,N_6210,N_5570);
and U9798 (N_9798,N_6511,N_6892);
nor U9799 (N_9799,N_5158,N_6961);
and U9800 (N_9800,N_7451,N_5712);
and U9801 (N_9801,N_5674,N_6448);
nand U9802 (N_9802,N_6542,N_5692);
or U9803 (N_9803,N_5932,N_6782);
xnor U9804 (N_9804,N_6490,N_6141);
xnor U9805 (N_9805,N_5928,N_7095);
or U9806 (N_9806,N_7338,N_5928);
nand U9807 (N_9807,N_7288,N_6815);
nand U9808 (N_9808,N_5460,N_7147);
or U9809 (N_9809,N_5520,N_5117);
and U9810 (N_9810,N_5055,N_5446);
xor U9811 (N_9811,N_5545,N_6987);
xnor U9812 (N_9812,N_5562,N_5626);
nor U9813 (N_9813,N_6619,N_6340);
nand U9814 (N_9814,N_6720,N_7408);
and U9815 (N_9815,N_5312,N_6256);
and U9816 (N_9816,N_5613,N_5698);
and U9817 (N_9817,N_5161,N_6395);
or U9818 (N_9818,N_7056,N_5044);
xnor U9819 (N_9819,N_6391,N_7233);
and U9820 (N_9820,N_5092,N_6325);
nand U9821 (N_9821,N_6425,N_5494);
and U9822 (N_9822,N_6983,N_5599);
nor U9823 (N_9823,N_6708,N_5188);
xnor U9824 (N_9824,N_5515,N_5789);
nand U9825 (N_9825,N_5900,N_7238);
and U9826 (N_9826,N_6257,N_5247);
xor U9827 (N_9827,N_6032,N_5525);
nand U9828 (N_9828,N_5275,N_5199);
nand U9829 (N_9829,N_6056,N_5713);
and U9830 (N_9830,N_7111,N_7185);
or U9831 (N_9831,N_7211,N_6445);
xor U9832 (N_9832,N_5701,N_5238);
xnor U9833 (N_9833,N_5650,N_6267);
nor U9834 (N_9834,N_5636,N_6358);
xnor U9835 (N_9835,N_5794,N_5347);
nand U9836 (N_9836,N_5785,N_7259);
or U9837 (N_9837,N_5295,N_5071);
or U9838 (N_9838,N_5815,N_5372);
nand U9839 (N_9839,N_6233,N_7385);
nor U9840 (N_9840,N_7242,N_7355);
or U9841 (N_9841,N_6554,N_6516);
and U9842 (N_9842,N_6675,N_5178);
xnor U9843 (N_9843,N_7177,N_6770);
nor U9844 (N_9844,N_6684,N_5279);
and U9845 (N_9845,N_6857,N_6945);
xor U9846 (N_9846,N_5007,N_6676);
nand U9847 (N_9847,N_5464,N_7204);
and U9848 (N_9848,N_6057,N_6785);
xnor U9849 (N_9849,N_6800,N_6563);
and U9850 (N_9850,N_6249,N_6967);
nand U9851 (N_9851,N_7016,N_5167);
nor U9852 (N_9852,N_5099,N_7457);
and U9853 (N_9853,N_6665,N_7089);
xnor U9854 (N_9854,N_7036,N_6162);
xor U9855 (N_9855,N_5908,N_7381);
nand U9856 (N_9856,N_6644,N_7472);
or U9857 (N_9857,N_5166,N_7163);
nand U9858 (N_9858,N_5138,N_5187);
nand U9859 (N_9859,N_6897,N_5379);
or U9860 (N_9860,N_5645,N_7328);
nand U9861 (N_9861,N_6806,N_6775);
nand U9862 (N_9862,N_6764,N_7001);
and U9863 (N_9863,N_7407,N_5049);
or U9864 (N_9864,N_6204,N_5515);
nand U9865 (N_9865,N_7190,N_5468);
nand U9866 (N_9866,N_5316,N_6780);
xnor U9867 (N_9867,N_5655,N_5806);
and U9868 (N_9868,N_7267,N_6635);
nand U9869 (N_9869,N_5728,N_5678);
nor U9870 (N_9870,N_6723,N_6088);
xnor U9871 (N_9871,N_7203,N_5927);
and U9872 (N_9872,N_6920,N_5933);
nand U9873 (N_9873,N_7244,N_5274);
xnor U9874 (N_9874,N_5523,N_6802);
xor U9875 (N_9875,N_6917,N_5938);
xnor U9876 (N_9876,N_6357,N_5848);
xnor U9877 (N_9877,N_5233,N_5631);
and U9878 (N_9878,N_6342,N_7342);
nor U9879 (N_9879,N_5537,N_6376);
or U9880 (N_9880,N_6413,N_7264);
nand U9881 (N_9881,N_6637,N_5003);
and U9882 (N_9882,N_6280,N_7184);
and U9883 (N_9883,N_7030,N_6868);
nor U9884 (N_9884,N_5203,N_5716);
or U9885 (N_9885,N_5264,N_6681);
nand U9886 (N_9886,N_5245,N_6864);
or U9887 (N_9887,N_7228,N_6447);
xnor U9888 (N_9888,N_6282,N_6348);
nor U9889 (N_9889,N_6305,N_6254);
xnor U9890 (N_9890,N_5898,N_6614);
or U9891 (N_9891,N_7110,N_5289);
nor U9892 (N_9892,N_6920,N_6212);
or U9893 (N_9893,N_6722,N_5920);
and U9894 (N_9894,N_5914,N_5245);
nor U9895 (N_9895,N_5955,N_5446);
nor U9896 (N_9896,N_5410,N_5417);
nor U9897 (N_9897,N_5751,N_5970);
xnor U9898 (N_9898,N_6376,N_5487);
nor U9899 (N_9899,N_6845,N_5679);
nor U9900 (N_9900,N_7435,N_5093);
and U9901 (N_9901,N_7447,N_6035);
xnor U9902 (N_9902,N_5686,N_7192);
and U9903 (N_9903,N_6600,N_7112);
nor U9904 (N_9904,N_5456,N_7478);
nand U9905 (N_9905,N_7493,N_5127);
nand U9906 (N_9906,N_6486,N_5063);
or U9907 (N_9907,N_7273,N_5807);
and U9908 (N_9908,N_7359,N_5832);
nor U9909 (N_9909,N_6220,N_7160);
nand U9910 (N_9910,N_5549,N_6712);
nand U9911 (N_9911,N_6225,N_6500);
nand U9912 (N_9912,N_6044,N_5103);
xor U9913 (N_9913,N_5699,N_5782);
nor U9914 (N_9914,N_6795,N_6979);
xnor U9915 (N_9915,N_5967,N_5294);
nand U9916 (N_9916,N_6086,N_5824);
nand U9917 (N_9917,N_5785,N_5285);
nor U9918 (N_9918,N_6675,N_6683);
xnor U9919 (N_9919,N_6310,N_7241);
nand U9920 (N_9920,N_7435,N_5671);
or U9921 (N_9921,N_6974,N_7446);
and U9922 (N_9922,N_6626,N_5381);
and U9923 (N_9923,N_6932,N_6188);
nor U9924 (N_9924,N_6310,N_7222);
nand U9925 (N_9925,N_7377,N_6891);
xor U9926 (N_9926,N_5047,N_6512);
nor U9927 (N_9927,N_6120,N_5125);
xor U9928 (N_9928,N_5737,N_6046);
nor U9929 (N_9929,N_6162,N_5651);
xor U9930 (N_9930,N_6591,N_6739);
xnor U9931 (N_9931,N_5870,N_5303);
nor U9932 (N_9932,N_6167,N_6245);
and U9933 (N_9933,N_7353,N_6625);
xnor U9934 (N_9934,N_7181,N_6753);
and U9935 (N_9935,N_6648,N_6845);
or U9936 (N_9936,N_6312,N_6888);
nor U9937 (N_9937,N_5772,N_6097);
nor U9938 (N_9938,N_6025,N_6506);
xnor U9939 (N_9939,N_5656,N_6402);
or U9940 (N_9940,N_6297,N_7163);
nand U9941 (N_9941,N_5043,N_5827);
xnor U9942 (N_9942,N_5071,N_6420);
or U9943 (N_9943,N_7325,N_6743);
or U9944 (N_9944,N_5503,N_5645);
nand U9945 (N_9945,N_6048,N_5242);
and U9946 (N_9946,N_6032,N_6146);
nand U9947 (N_9947,N_6142,N_7433);
nor U9948 (N_9948,N_5905,N_6370);
or U9949 (N_9949,N_6685,N_6982);
nor U9950 (N_9950,N_5720,N_6543);
nand U9951 (N_9951,N_6808,N_5886);
nand U9952 (N_9952,N_6001,N_7473);
or U9953 (N_9953,N_7334,N_6109);
xor U9954 (N_9954,N_6596,N_7294);
nand U9955 (N_9955,N_5782,N_6575);
xnor U9956 (N_9956,N_5839,N_5265);
or U9957 (N_9957,N_5810,N_6714);
and U9958 (N_9958,N_5284,N_5504);
and U9959 (N_9959,N_7093,N_7119);
nand U9960 (N_9960,N_5743,N_5563);
xor U9961 (N_9961,N_5225,N_5753);
nand U9962 (N_9962,N_6697,N_6914);
and U9963 (N_9963,N_7180,N_5879);
nand U9964 (N_9964,N_6086,N_6357);
and U9965 (N_9965,N_6706,N_6962);
and U9966 (N_9966,N_5883,N_5080);
nand U9967 (N_9967,N_5673,N_5097);
nor U9968 (N_9968,N_5747,N_6393);
xor U9969 (N_9969,N_6857,N_5119);
or U9970 (N_9970,N_7173,N_5869);
and U9971 (N_9971,N_7086,N_5980);
and U9972 (N_9972,N_5757,N_5290);
xnor U9973 (N_9973,N_7446,N_6082);
and U9974 (N_9974,N_5675,N_6709);
and U9975 (N_9975,N_7369,N_6948);
nand U9976 (N_9976,N_6787,N_5051);
or U9977 (N_9977,N_5861,N_5400);
or U9978 (N_9978,N_6297,N_5692);
and U9979 (N_9979,N_5520,N_7350);
xnor U9980 (N_9980,N_5531,N_5872);
xor U9981 (N_9981,N_6644,N_6820);
nor U9982 (N_9982,N_5406,N_7046);
or U9983 (N_9983,N_7475,N_5253);
xnor U9984 (N_9984,N_5836,N_5216);
and U9985 (N_9985,N_6345,N_5771);
nand U9986 (N_9986,N_7062,N_5584);
nor U9987 (N_9987,N_6809,N_7285);
and U9988 (N_9988,N_6337,N_5260);
or U9989 (N_9989,N_7163,N_6849);
or U9990 (N_9990,N_6811,N_6063);
nand U9991 (N_9991,N_5318,N_5125);
xnor U9992 (N_9992,N_7396,N_7282);
xor U9993 (N_9993,N_5291,N_5110);
or U9994 (N_9994,N_6742,N_5306);
nand U9995 (N_9995,N_5308,N_6568);
xor U9996 (N_9996,N_5766,N_5414);
nand U9997 (N_9997,N_5639,N_6253);
or U9998 (N_9998,N_7499,N_7034);
and U9999 (N_9999,N_5699,N_6395);
or U10000 (N_10000,N_9699,N_9677);
and U10001 (N_10001,N_9347,N_8158);
xnor U10002 (N_10002,N_9458,N_7796);
nor U10003 (N_10003,N_9614,N_7713);
nor U10004 (N_10004,N_9781,N_8527);
xor U10005 (N_10005,N_8595,N_9240);
nor U10006 (N_10006,N_7693,N_8689);
nand U10007 (N_10007,N_8704,N_8440);
xnor U10008 (N_10008,N_7592,N_8938);
nor U10009 (N_10009,N_8063,N_8543);
or U10010 (N_10010,N_9535,N_9574);
and U10011 (N_10011,N_9715,N_8872);
xor U10012 (N_10012,N_8336,N_8651);
xnor U10013 (N_10013,N_7614,N_7945);
and U10014 (N_10014,N_9344,N_9595);
or U10015 (N_10015,N_7805,N_9890);
xnor U10016 (N_10016,N_8245,N_7867);
nand U10017 (N_10017,N_9943,N_8909);
xnor U10018 (N_10018,N_9519,N_7588);
xnor U10019 (N_10019,N_8427,N_9227);
and U10020 (N_10020,N_8801,N_8400);
nand U10021 (N_10021,N_9571,N_8284);
xor U10022 (N_10022,N_7966,N_9159);
nand U10023 (N_10023,N_9246,N_9467);
and U10024 (N_10024,N_7613,N_7608);
or U10025 (N_10025,N_7745,N_9705);
or U10026 (N_10026,N_7638,N_8764);
or U10027 (N_10027,N_9087,N_7985);
or U10028 (N_10028,N_9432,N_8627);
nor U10029 (N_10029,N_9049,N_9256);
nor U10030 (N_10030,N_8438,N_9929);
nand U10031 (N_10031,N_7685,N_8977);
xnor U10032 (N_10032,N_7850,N_9996);
nand U10033 (N_10033,N_7629,N_7542);
xor U10034 (N_10034,N_9094,N_9767);
xnor U10035 (N_10035,N_8496,N_8837);
and U10036 (N_10036,N_8673,N_8809);
and U10037 (N_10037,N_7816,N_8098);
nand U10038 (N_10038,N_8684,N_8469);
nand U10039 (N_10039,N_8424,N_8896);
or U10040 (N_10040,N_9731,N_8505);
nand U10041 (N_10041,N_9971,N_9418);
nor U10042 (N_10042,N_9865,N_9090);
nand U10043 (N_10043,N_8688,N_9913);
xnor U10044 (N_10044,N_9176,N_8827);
xnor U10045 (N_10045,N_8854,N_9386);
and U10046 (N_10046,N_8416,N_9839);
and U10047 (N_10047,N_8589,N_8575);
nor U10048 (N_10048,N_7936,N_9431);
nand U10049 (N_10049,N_8293,N_9590);
xor U10050 (N_10050,N_9204,N_9068);
and U10051 (N_10051,N_8934,N_9710);
and U10052 (N_10052,N_9026,N_9046);
or U10053 (N_10053,N_8492,N_7991);
nand U10054 (N_10054,N_8329,N_9529);
nor U10055 (N_10055,N_8932,N_8221);
or U10056 (N_10056,N_9345,N_9277);
xor U10057 (N_10057,N_8666,N_7730);
nand U10058 (N_10058,N_9324,N_8697);
and U10059 (N_10059,N_7659,N_8756);
or U10060 (N_10060,N_9258,N_9270);
and U10061 (N_10061,N_8136,N_8035);
nor U10062 (N_10062,N_9420,N_7690);
or U10063 (N_10063,N_9525,N_8487);
nand U10064 (N_10064,N_9106,N_8762);
or U10065 (N_10065,N_9138,N_9372);
xor U10066 (N_10066,N_8351,N_8774);
nand U10067 (N_10067,N_9442,N_9761);
and U10068 (N_10068,N_9000,N_7615);
or U10069 (N_10069,N_9294,N_8209);
xor U10070 (N_10070,N_9080,N_9904);
or U10071 (N_10071,N_7997,N_7533);
and U10072 (N_10072,N_8822,N_9764);
xor U10073 (N_10073,N_7898,N_9237);
and U10074 (N_10074,N_8460,N_9282);
and U10075 (N_10075,N_9945,N_8142);
xnor U10076 (N_10076,N_8632,N_9437);
nand U10077 (N_10077,N_9228,N_9663);
xnor U10078 (N_10078,N_8623,N_8449);
or U10079 (N_10079,N_8509,N_9422);
and U10080 (N_10080,N_8171,N_7522);
nand U10081 (N_10081,N_7746,N_7982);
and U10082 (N_10082,N_8728,N_9690);
xnor U10083 (N_10083,N_8444,N_8312);
xor U10084 (N_10084,N_8746,N_7950);
and U10085 (N_10085,N_9718,N_9393);
nor U10086 (N_10086,N_9735,N_8381);
nand U10087 (N_10087,N_9114,N_9544);
and U10088 (N_10088,N_9005,N_9889);
xnor U10089 (N_10089,N_9877,N_9275);
nor U10090 (N_10090,N_8213,N_8576);
xor U10091 (N_10091,N_8753,N_7649);
nand U10092 (N_10092,N_9615,N_8411);
xor U10093 (N_10093,N_8493,N_9626);
and U10094 (N_10094,N_7605,N_9668);
or U10095 (N_10095,N_7541,N_7590);
nor U10096 (N_10096,N_9619,N_9445);
nand U10097 (N_10097,N_7680,N_8302);
or U10098 (N_10098,N_7502,N_8160);
and U10099 (N_10099,N_7924,N_7820);
and U10100 (N_10100,N_8974,N_9694);
nand U10101 (N_10101,N_9105,N_9378);
nand U10102 (N_10102,N_7569,N_8920);
nand U10103 (N_10103,N_9370,N_8154);
and U10104 (N_10104,N_8795,N_9400);
or U10105 (N_10105,N_8625,N_9265);
or U10106 (N_10106,N_9888,N_9512);
nor U10107 (N_10107,N_7506,N_7549);
and U10108 (N_10108,N_9522,N_7666);
xor U10109 (N_10109,N_7989,N_8393);
nor U10110 (N_10110,N_9084,N_8436);
nor U10111 (N_10111,N_9513,N_8294);
nand U10112 (N_10112,N_8260,N_7813);
and U10113 (N_10113,N_9131,N_9536);
and U10114 (N_10114,N_8242,N_8707);
nand U10115 (N_10115,N_7594,N_8929);
or U10116 (N_10116,N_8007,N_8549);
xor U10117 (N_10117,N_8922,N_9464);
nand U10118 (N_10118,N_8499,N_9920);
or U10119 (N_10119,N_7915,N_8755);
nor U10120 (N_10120,N_7508,N_8188);
nor U10121 (N_10121,N_7926,N_8378);
or U10122 (N_10122,N_9340,N_8232);
nor U10123 (N_10123,N_7878,N_7849);
xor U10124 (N_10124,N_8249,N_9585);
and U10125 (N_10125,N_9686,N_8280);
or U10126 (N_10126,N_7951,N_9436);
xnor U10127 (N_10127,N_8374,N_7540);
xnor U10128 (N_10128,N_9381,N_8373);
nand U10129 (N_10129,N_8616,N_9992);
nand U10130 (N_10130,N_7869,N_7581);
xnor U10131 (N_10131,N_9855,N_9385);
xnor U10132 (N_10132,N_7505,N_8667);
xor U10133 (N_10133,N_7800,N_8330);
xnor U10134 (N_10134,N_9419,N_8129);
nor U10135 (N_10135,N_8803,N_8049);
nor U10136 (N_10136,N_9763,N_8453);
and U10137 (N_10137,N_9772,N_8092);
nand U10138 (N_10138,N_8268,N_8241);
xor U10139 (N_10139,N_8058,N_7977);
and U10140 (N_10140,N_8200,N_9142);
nor U10141 (N_10141,N_9773,N_8617);
or U10142 (N_10142,N_8364,N_9652);
nor U10143 (N_10143,N_7748,N_9933);
or U10144 (N_10144,N_8603,N_8586);
and U10145 (N_10145,N_8880,N_7510);
nor U10146 (N_10146,N_7828,N_8996);
nor U10147 (N_10147,N_9124,N_7759);
or U10148 (N_10148,N_8554,N_9955);
and U10149 (N_10149,N_8199,N_8950);
nor U10150 (N_10150,N_9112,N_7584);
xor U10151 (N_10151,N_9438,N_7794);
or U10152 (N_10152,N_9576,N_8788);
nor U10153 (N_10153,N_7689,N_9322);
xnor U10154 (N_10154,N_7777,N_9483);
nand U10155 (N_10155,N_8395,N_9244);
nand U10156 (N_10156,N_9852,N_8150);
xor U10157 (N_10157,N_9359,N_9175);
nor U10158 (N_10158,N_9739,N_9328);
and U10159 (N_10159,N_9061,N_7665);
or U10160 (N_10160,N_9791,N_9456);
nor U10161 (N_10161,N_9632,N_9224);
nand U10162 (N_10162,N_9880,N_7792);
or U10163 (N_10163,N_7607,N_7706);
xnor U10164 (N_10164,N_9448,N_9021);
nand U10165 (N_10165,N_9798,N_7988);
and U10166 (N_10166,N_8079,N_8958);
xnor U10167 (N_10167,N_8006,N_8478);
and U10168 (N_10168,N_8238,N_8301);
or U10169 (N_10169,N_8512,N_9274);
nand U10170 (N_10170,N_9681,N_7735);
nand U10171 (N_10171,N_9011,N_9104);
and U10172 (N_10172,N_9618,N_9493);
and U10173 (N_10173,N_9130,N_8966);
or U10174 (N_10174,N_7600,N_9495);
and U10175 (N_10175,N_7975,N_8005);
nand U10176 (N_10176,N_8733,N_8850);
and U10177 (N_10177,N_8708,N_9414);
or U10178 (N_10178,N_8531,N_9390);
nor U10179 (N_10179,N_8484,N_8779);
and U10180 (N_10180,N_8776,N_9022);
nand U10181 (N_10181,N_8626,N_9942);
and U10182 (N_10182,N_8610,N_7925);
nor U10183 (N_10183,N_9559,N_9169);
nor U10184 (N_10184,N_7998,N_8044);
and U10185 (N_10185,N_9696,N_7696);
or U10186 (N_10186,N_8672,N_8676);
or U10187 (N_10187,N_9064,N_8608);
and U10188 (N_10188,N_9266,N_8220);
nand U10189 (N_10189,N_7705,N_8437);
nand U10190 (N_10190,N_9081,N_8376);
nand U10191 (N_10191,N_9156,N_7655);
or U10192 (N_10192,N_9205,N_9801);
and U10193 (N_10193,N_8009,N_7577);
and U10194 (N_10194,N_7716,N_7625);
or U10195 (N_10195,N_9478,N_8816);
or U10196 (N_10196,N_9757,N_7532);
and U10197 (N_10197,N_7531,N_9332);
and U10198 (N_10198,N_9398,N_8725);
xor U10199 (N_10199,N_8352,N_9167);
nand U10200 (N_10200,N_9895,N_7793);
or U10201 (N_10201,N_8927,N_8555);
and U10202 (N_10202,N_8992,N_9617);
nor U10203 (N_10203,N_8088,N_7788);
or U10204 (N_10204,N_9966,N_8468);
and U10205 (N_10205,N_9160,N_7894);
nor U10206 (N_10206,N_7984,N_7664);
nor U10207 (N_10207,N_9222,N_9709);
xnor U10208 (N_10208,N_7809,N_8262);
nand U10209 (N_10209,N_7661,N_8569);
nand U10210 (N_10210,N_8291,N_8745);
nor U10211 (N_10211,N_9367,N_8017);
or U10212 (N_10212,N_7741,N_9999);
and U10213 (N_10213,N_9233,N_8955);
nand U10214 (N_10214,N_7518,N_7635);
nor U10215 (N_10215,N_9316,N_7775);
nor U10216 (N_10216,N_8326,N_9113);
nor U10217 (N_10217,N_8693,N_9285);
nand U10218 (N_10218,N_9582,N_8045);
or U10219 (N_10219,N_7683,N_9965);
or U10220 (N_10220,N_8450,N_7593);
or U10221 (N_10221,N_7598,N_7802);
and U10222 (N_10222,N_8240,N_7815);
nand U10223 (N_10223,N_9015,N_8075);
nor U10224 (N_10224,N_9994,N_9866);
and U10225 (N_10225,N_8462,N_7561);
nand U10226 (N_10226,N_8137,N_9778);
nor U10227 (N_10227,N_9125,N_9206);
nand U10228 (N_10228,N_9713,N_9726);
and U10229 (N_10229,N_7737,N_9701);
xor U10230 (N_10230,N_7524,N_7731);
nand U10231 (N_10231,N_9666,N_9982);
and U10232 (N_10232,N_9520,N_9981);
xor U10233 (N_10233,N_8897,N_9541);
xnor U10234 (N_10234,N_8784,N_7643);
or U10235 (N_10235,N_8338,N_8159);
xor U10236 (N_10236,N_8546,N_9162);
or U10237 (N_10237,N_9230,N_8204);
or U10238 (N_10238,N_8176,N_9546);
or U10239 (N_10239,N_7740,N_8838);
or U10240 (N_10240,N_8573,N_8208);
xor U10241 (N_10241,N_7896,N_8093);
or U10242 (N_10242,N_9411,N_8452);
nand U10243 (N_10243,N_8144,N_9872);
and U10244 (N_10244,N_9271,N_8180);
nand U10245 (N_10245,N_7993,N_9408);
xor U10246 (N_10246,N_8961,N_8128);
and U10247 (N_10247,N_9697,N_9181);
nand U10248 (N_10248,N_8706,N_8895);
or U10249 (N_10249,N_8490,N_8796);
xnor U10250 (N_10250,N_9995,N_9837);
xnor U10251 (N_10251,N_8466,N_9391);
and U10252 (N_10252,N_9262,N_7965);
and U10253 (N_10253,N_9504,N_7630);
nand U10254 (N_10254,N_8949,N_7776);
nand U10255 (N_10255,N_9521,N_9178);
or U10256 (N_10256,N_9816,N_8646);
nor U10257 (N_10257,N_8866,N_9315);
and U10258 (N_10258,N_9864,N_7931);
nand U10259 (N_10259,N_7606,N_8334);
or U10260 (N_10260,N_8973,N_8507);
nor U10261 (N_10261,N_8071,N_9292);
or U10262 (N_10262,N_7890,N_8047);
or U10263 (N_10263,N_8034,N_9330);
nand U10264 (N_10264,N_9514,N_9035);
or U10265 (N_10265,N_9631,N_8399);
nor U10266 (N_10266,N_7576,N_8864);
and U10267 (N_10267,N_8985,N_7960);
and U10268 (N_10268,N_7529,N_7546);
and U10269 (N_10269,N_9264,N_9691);
xnor U10270 (N_10270,N_9384,N_8924);
xor U10271 (N_10271,N_8313,N_8513);
nor U10272 (N_10272,N_9313,N_7801);
and U10273 (N_10273,N_9818,N_8102);
xnor U10274 (N_10274,N_9070,N_8739);
nor U10275 (N_10275,N_7919,N_8544);
or U10276 (N_10276,N_8723,N_7906);
nor U10277 (N_10277,N_7641,N_8463);
and U10278 (N_10278,N_8890,N_9883);
xor U10279 (N_10279,N_9100,N_8299);
nand U10280 (N_10280,N_7921,N_9314);
nand U10281 (N_10281,N_9812,N_7623);
xnor U10282 (N_10282,N_9202,N_9171);
nor U10283 (N_10283,N_8628,N_9191);
xnor U10284 (N_10284,N_7722,N_8681);
nand U10285 (N_10285,N_9479,N_9874);
or U10286 (N_10286,N_8067,N_8211);
or U10287 (N_10287,N_8911,N_9357);
xor U10288 (N_10288,N_8471,N_9117);
and U10289 (N_10289,N_9101,N_7647);
or U10290 (N_10290,N_8057,N_9916);
nor U10291 (N_10291,N_8138,N_8791);
or U10292 (N_10292,N_7891,N_9062);
and U10293 (N_10293,N_7912,N_8547);
xnor U10294 (N_10294,N_9789,N_9774);
nor U10295 (N_10295,N_9922,N_9607);
and U10296 (N_10296,N_8127,N_7574);
or U10297 (N_10297,N_8683,N_9008);
nor U10298 (N_10298,N_8679,N_8849);
or U10299 (N_10299,N_8821,N_8590);
nand U10300 (N_10300,N_9466,N_7612);
xor U10301 (N_10301,N_8968,N_8303);
nand U10302 (N_10302,N_9486,N_9579);
and U10303 (N_10303,N_9099,N_9402);
nor U10304 (N_10304,N_9291,N_7562);
nand U10305 (N_10305,N_9949,N_8808);
nand U10306 (N_10306,N_9148,N_9882);
nor U10307 (N_10307,N_8182,N_9803);
nor U10308 (N_10308,N_9564,N_9469);
xor U10309 (N_10309,N_9983,N_9517);
nand U10310 (N_10310,N_9901,N_8143);
nand U10311 (N_10311,N_9050,N_8514);
xor U10312 (N_10312,N_8644,N_8747);
xor U10313 (N_10313,N_8494,N_8223);
nor U10314 (N_10314,N_8168,N_7835);
nor U10315 (N_10315,N_7637,N_8883);
nor U10316 (N_10316,N_8935,N_9255);
or U10317 (N_10317,N_9986,N_9775);
nor U10318 (N_10318,N_9638,N_8570);
xor U10319 (N_10319,N_9675,N_8867);
nor U10320 (N_10320,N_7918,N_7628);
xnor U10321 (N_10321,N_7750,N_7855);
or U10322 (N_10322,N_9562,N_7553);
nand U10323 (N_10323,N_8542,N_7539);
or U10324 (N_10324,N_9443,N_8363);
nor U10325 (N_10325,N_9288,N_8852);
and U10326 (N_10326,N_9042,N_7787);
nor U10327 (N_10327,N_8674,N_9454);
nand U10328 (N_10328,N_9123,N_9948);
nor U10329 (N_10329,N_8271,N_8279);
nor U10330 (N_10330,N_7939,N_8042);
xor U10331 (N_10331,N_7969,N_7947);
or U10332 (N_10332,N_7871,N_9599);
nand U10333 (N_10333,N_8853,N_9079);
nor U10334 (N_10334,N_9001,N_9018);
and U10335 (N_10335,N_7956,N_7674);
xor U10336 (N_10336,N_9425,N_9656);
and U10337 (N_10337,N_8548,N_7856);
xnor U10338 (N_10338,N_7699,N_9056);
or U10339 (N_10339,N_8201,N_9847);
nand U10340 (N_10340,N_9980,N_9587);
nor U10341 (N_10341,N_8988,N_9034);
xor U10342 (N_10342,N_8141,N_8203);
xnor U10343 (N_10343,N_7917,N_8224);
xor U10344 (N_10344,N_9953,N_9251);
and U10345 (N_10345,N_8162,N_8076);
and U10346 (N_10346,N_9065,N_9349);
xor U10347 (N_10347,N_9896,N_8165);
nand U10348 (N_10348,N_8439,N_8314);
nand U10349 (N_10349,N_9024,N_9993);
or U10350 (N_10350,N_7587,N_8878);
xor U10351 (N_10351,N_8729,N_9932);
xor U10352 (N_10352,N_9811,N_8421);
xor U10353 (N_10353,N_9215,N_8435);
nor U10354 (N_10354,N_8842,N_9166);
xor U10355 (N_10355,N_7738,N_8031);
nand U10356 (N_10356,N_9412,N_8018);
nand U10357 (N_10357,N_7701,N_8670);
nor U10358 (N_10358,N_7648,N_9450);
and U10359 (N_10359,N_9762,N_7782);
nor U10360 (N_10360,N_8033,N_8173);
xor U10361 (N_10361,N_8701,N_9814);
or U10362 (N_10362,N_7718,N_9199);
and U10363 (N_10363,N_9527,N_8959);
nor U10364 (N_10364,N_7525,N_9293);
nand U10365 (N_10365,N_8823,N_8050);
and U10366 (N_10366,N_8323,N_7953);
nand U10367 (N_10367,N_7751,N_8792);
nor U10368 (N_10368,N_9241,N_7838);
xnor U10369 (N_10369,N_9613,N_7749);
xnor U10370 (N_10370,N_8412,N_7575);
xnor U10371 (N_10371,N_7824,N_8720);
or U10372 (N_10372,N_7538,N_8828);
and U10373 (N_10373,N_9635,N_9558);
or U10374 (N_10374,N_8010,N_8155);
nor U10375 (N_10375,N_9441,N_9195);
or U10376 (N_10376,N_7753,N_9433);
xnor U10377 (N_10377,N_9161,N_7762);
xor U10378 (N_10378,N_7513,N_8321);
nor U10379 (N_10379,N_8016,N_9609);
nand U10380 (N_10380,N_8954,N_9563);
xor U10381 (N_10381,N_9792,N_9914);
and U10382 (N_10382,N_8431,N_9484);
xnor U10383 (N_10383,N_9268,N_7865);
nand U10384 (N_10384,N_9845,N_7994);
or U10385 (N_10385,N_7876,N_8524);
nor U10386 (N_10386,N_9231,N_8658);
or U10387 (N_10387,N_7589,N_9339);
xnor U10388 (N_10388,N_7724,N_8552);
nor U10389 (N_10389,N_8675,N_9729);
xor U10390 (N_10390,N_8041,N_9144);
nor U10391 (N_10391,N_9962,N_9452);
or U10392 (N_10392,N_9586,N_9998);
nand U10393 (N_10393,N_8522,N_8454);
nand U10394 (N_10394,N_8122,N_7818);
nor U10395 (N_10395,N_8559,N_9250);
or U10396 (N_10396,N_7551,N_9006);
or U10397 (N_10397,N_8885,N_9236);
nand U10398 (N_10398,N_8698,N_8430);
nand U10399 (N_10399,N_7563,N_9537);
nand U10400 (N_10400,N_8078,N_7955);
or U10401 (N_10401,N_8773,N_9601);
nand U10402 (N_10402,N_8120,N_8389);
and U10403 (N_10403,N_7703,N_7842);
xnor U10404 (N_10404,N_9598,N_8802);
and U10405 (N_10405,N_7986,N_7946);
and U10406 (N_10406,N_8292,N_9620);
nor U10407 (N_10407,N_9926,N_9526);
and U10408 (N_10408,N_9040,N_8037);
nand U10409 (N_10409,N_9978,N_9790);
xor U10410 (N_10410,N_9930,N_9703);
xor U10411 (N_10411,N_9821,N_9232);
xor U10412 (N_10412,N_9780,N_7672);
nor U10413 (N_10413,N_8947,N_8163);
or U10414 (N_10414,N_7983,N_8624);
or U10415 (N_10415,N_9239,N_9854);
or U10416 (N_10416,N_9132,N_9766);
or U10417 (N_10417,N_9279,N_9216);
nor U10418 (N_10418,N_9891,N_8845);
and U10419 (N_10419,N_7515,N_8406);
or U10420 (N_10420,N_7814,N_9044);
nor U10421 (N_10421,N_9407,N_9333);
xor U10422 (N_10422,N_9047,N_8216);
nand U10423 (N_10423,N_8648,N_9426);
nor U10424 (N_10424,N_8342,N_8426);
and U10425 (N_10425,N_8053,N_7781);
nand U10426 (N_10426,N_9947,N_8653);
xor U10427 (N_10427,N_9145,N_9298);
or U10428 (N_10428,N_9665,N_8804);
nor U10429 (N_10429,N_9906,N_9146);
or U10430 (N_10430,N_7610,N_9894);
nand U10431 (N_10431,N_9730,N_9502);
nor U10432 (N_10432,N_8056,N_9405);
or U10433 (N_10433,N_9010,N_9187);
nand U10434 (N_10434,N_8497,N_9873);
and U10435 (N_10435,N_8072,N_8170);
and U10436 (N_10436,N_9606,N_7543);
nand U10437 (N_10437,N_8715,N_9941);
and U10438 (N_10438,N_9645,N_9281);
xnor U10439 (N_10439,N_9211,N_8059);
nand U10440 (N_10440,N_8761,N_8147);
and U10441 (N_10441,N_8353,N_8906);
nand U10442 (N_10442,N_9753,N_9720);
or U10443 (N_10443,N_9115,N_9136);
or U10444 (N_10444,N_8596,N_9155);
nand U10445 (N_10445,N_8811,N_9687);
xor U10446 (N_10446,N_8065,N_9312);
xor U10447 (N_10447,N_7893,N_7785);
or U10448 (N_10448,N_8664,N_8140);
or U10449 (N_10449,N_8630,N_8343);
nor U10450 (N_10450,N_8396,N_8545);
nand U10451 (N_10451,N_8486,N_8928);
nor U10452 (N_10452,N_8181,N_8479);
nor U10453 (N_10453,N_8686,N_8831);
nor U10454 (N_10454,N_8286,N_8978);
and U10455 (N_10455,N_8036,N_8488);
nor U10456 (N_10456,N_8750,N_8340);
xnor U10457 (N_10457,N_9154,N_8783);
or U10458 (N_10458,N_9179,N_8536);
xnor U10459 (N_10459,N_8498,N_7920);
xnor U10460 (N_10460,N_9083,N_8121);
and U10461 (N_10461,N_8807,N_9457);
nor U10462 (N_10462,N_7847,N_9908);
and U10463 (N_10463,N_8222,N_7821);
nor U10464 (N_10464,N_7653,N_9193);
nand U10465 (N_10465,N_8969,N_9556);
xnor U10466 (N_10466,N_8278,N_8726);
nand U10467 (N_10467,N_7725,N_8191);
and U10468 (N_10468,N_9515,N_7756);
nor U10469 (N_10469,N_9952,N_7678);
nor U10470 (N_10470,N_8682,N_8228);
xor U10471 (N_10471,N_7959,N_7761);
nand U10472 (N_10472,N_7857,N_9449);
or U10473 (N_10473,N_7790,N_9956);
nor U10474 (N_10474,N_9900,N_8981);
nor U10475 (N_10475,N_8477,N_8521);
nor U10476 (N_10476,N_9836,N_9698);
xor U10477 (N_10477,N_9267,N_9902);
nand U10478 (N_10478,N_9936,N_8465);
nand U10479 (N_10479,N_9884,N_8250);
and U10480 (N_10480,N_8769,N_9055);
and U10481 (N_10481,N_9487,N_9338);
nand U10482 (N_10482,N_9905,N_7688);
nand U10483 (N_10483,N_8282,N_7990);
or U10484 (N_10484,N_9724,N_7527);
nand U10485 (N_10485,N_7810,N_8881);
or U10486 (N_10486,N_8066,N_9575);
xnor U10487 (N_10487,N_9898,N_8384);
xnor U10488 (N_10488,N_9401,N_9572);
or U10489 (N_10489,N_8383,N_8556);
nand U10490 (N_10490,N_9122,N_9197);
nand U10491 (N_10491,N_9625,N_8350);
xor U10492 (N_10492,N_9168,N_9301);
or U10493 (N_10493,N_8873,N_8198);
xor U10494 (N_10494,N_8135,N_7866);
xnor U10495 (N_10495,N_9085,N_7772);
xnor U10496 (N_10496,N_9848,N_9406);
or U10497 (N_10497,N_7804,N_7864);
or U10498 (N_10498,N_7773,N_7719);
or U10499 (N_10499,N_8095,N_9334);
xor U10500 (N_10500,N_9499,N_9867);
nand U10501 (N_10501,N_7597,N_9033);
nand U10502 (N_10502,N_7884,N_8239);
or U10503 (N_10503,N_9743,N_7507);
or U10504 (N_10504,N_9610,N_8749);
and U10505 (N_10505,N_7654,N_9640);
nor U10506 (N_10506,N_7897,N_7870);
or U10507 (N_10507,N_8819,N_8660);
and U10508 (N_10508,N_7806,N_7798);
or U10509 (N_10509,N_9984,N_7684);
nand U10510 (N_10510,N_8022,N_8960);
nand U10511 (N_10511,N_9716,N_9069);
nor U10512 (N_10512,N_8923,N_8296);
or U10513 (N_10513,N_9799,N_9657);
and U10514 (N_10514,N_9152,N_9651);
xnor U10515 (N_10515,N_9004,N_7770);
and U10516 (N_10516,N_8711,N_7544);
xnor U10517 (N_10517,N_9972,N_8090);
xnor U10518 (N_10518,N_8540,N_9157);
nor U10519 (N_10519,N_9505,N_9082);
xor U10520 (N_10520,N_7651,N_9603);
xor U10521 (N_10521,N_8295,N_9283);
nand U10522 (N_10522,N_9832,N_9219);
and U10523 (N_10523,N_9793,N_8735);
and U10524 (N_10524,N_8613,N_9897);
nand U10525 (N_10525,N_8415,N_8495);
and U10526 (N_10526,N_7803,N_8834);
nor U10527 (N_10527,N_8003,N_8347);
xor U10528 (N_10528,N_9667,N_7545);
nand U10529 (N_10529,N_9350,N_9825);
nor U10530 (N_10530,N_8597,N_8967);
nand U10531 (N_10531,N_8306,N_8277);
nand U10532 (N_10532,N_8971,N_8101);
xor U10533 (N_10533,N_9560,N_9102);
xor U10534 (N_10534,N_8387,N_9455);
or U10535 (N_10535,N_8904,N_7779);
and U10536 (N_10536,N_9523,N_7836);
xor U10537 (N_10537,N_8775,N_7832);
nor U10538 (N_10538,N_9410,N_9850);
or U10539 (N_10539,N_7558,N_8585);
or U10540 (N_10540,N_8451,N_8768);
nor U10541 (N_10541,N_9485,N_9473);
nand U10542 (N_10542,N_9396,N_9353);
and U10543 (N_10543,N_7907,N_9352);
xor U10544 (N_10544,N_8337,N_7671);
nor U10545 (N_10545,N_9306,N_9118);
and U10546 (N_10546,N_9553,N_9462);
nand U10547 (N_10547,N_9247,N_9721);
nor U10548 (N_10548,N_9172,N_9403);
xor U10549 (N_10549,N_9822,N_7692);
and U10550 (N_10550,N_9428,N_9476);
or U10551 (N_10551,N_7889,N_9073);
nor U10552 (N_10552,N_9754,N_9838);
nor U10553 (N_10553,N_9950,N_8403);
nand U10554 (N_10554,N_9286,N_9565);
nor U10555 (N_10555,N_7769,N_8409);
nor U10556 (N_10556,N_8520,N_8328);
nor U10557 (N_10557,N_8917,N_9078);
nand U10558 (N_10558,N_9500,N_9800);
and U10559 (N_10559,N_9163,N_9459);
nand U10560 (N_10560,N_9689,N_8233);
and U10561 (N_10561,N_9654,N_8532);
and U10562 (N_10562,N_9795,N_8251);
and U10563 (N_10563,N_9758,N_9695);
or U10564 (N_10564,N_9899,N_8640);
nor U10565 (N_10565,N_9827,N_9133);
xnor U10566 (N_10566,N_7943,N_8738);
nand U10567 (N_10567,N_7941,N_9616);
and U10568 (N_10568,N_9810,N_8207);
or U10569 (N_10569,N_8040,N_9935);
nand U10570 (N_10570,N_7695,N_7922);
nand U10571 (N_10571,N_8609,N_9305);
xnor U10572 (N_10572,N_9508,N_8882);
or U10573 (N_10573,N_7667,N_7669);
and U10574 (N_10574,N_8357,N_7799);
nand U10575 (N_10575,N_9738,N_8744);
and U10576 (N_10576,N_9834,N_8841);
xnor U10577 (N_10577,N_9737,N_9057);
or U10578 (N_10578,N_9032,N_9321);
xnor U10579 (N_10579,N_9693,N_8618);
nor U10580 (N_10580,N_9659,N_9254);
or U10581 (N_10581,N_7662,N_8553);
or U10582 (N_10582,N_8107,N_9075);
xor U10583 (N_10583,N_9828,N_7712);
nand U10584 (N_10584,N_9573,N_7700);
nand U10585 (N_10585,N_7786,N_8826);
xor U10586 (N_10586,N_7521,N_9925);
nor U10587 (N_10587,N_9238,N_8273);
nand U10588 (N_10588,N_9538,N_9498);
and U10589 (N_10589,N_9351,N_8855);
nand U10590 (N_10590,N_8276,N_9550);
nand U10591 (N_10591,N_8702,N_9492);
nand U10592 (N_10592,N_8998,N_8694);
and U10593 (N_10593,N_9664,N_9875);
and U10594 (N_10594,N_8760,N_7642);
xor U10595 (N_10595,N_9819,N_7992);
nand U10596 (N_10596,N_8310,N_8951);
nand U10597 (N_10597,N_9600,N_8124);
and U10598 (N_10598,N_8870,N_7863);
nor U10599 (N_10599,N_8192,N_8943);
or U10600 (N_10600,N_8587,N_8269);
and U10601 (N_10601,N_7935,N_7783);
nor U10602 (N_10602,N_9088,N_8091);
and U10603 (N_10603,N_8259,N_9547);
nor U10604 (N_10604,N_9771,N_8069);
or U10605 (N_10605,N_7656,N_8080);
nand U10606 (N_10606,N_9964,N_9225);
and U10607 (N_10607,N_8705,N_8732);
nor U10608 (N_10608,N_8021,N_8964);
nor U10609 (N_10609,N_8111,N_9725);
xor U10610 (N_10610,N_9786,N_8606);
xnor U10611 (N_10611,N_9489,N_8741);
and U10612 (N_10612,N_7961,N_9346);
xnor U10613 (N_10613,N_8748,N_8846);
nor U10614 (N_10614,N_8386,N_7963);
or U10615 (N_10615,N_7973,N_8825);
xor U10616 (N_10616,N_7670,N_9869);
nand U10617 (N_10617,N_9229,N_8502);
and U10618 (N_10618,N_9658,N_9674);
or U10619 (N_10619,N_9253,N_9708);
xnor U10620 (N_10620,N_8461,N_7858);
or U10621 (N_10621,N_9649,N_8023);
nand U10622 (N_10622,N_8272,N_9967);
and U10623 (N_10623,N_8680,N_7578);
nand U10624 (N_10624,N_9141,N_8913);
nor U10625 (N_10625,N_9622,N_8533);
xnor U10626 (N_10626,N_9127,N_8936);
and U10627 (N_10627,N_7944,N_8480);
or U10628 (N_10628,N_7644,N_8563);
and U10629 (N_10629,N_7923,N_9361);
xnor U10630 (N_10630,N_8925,N_7624);
nand U10631 (N_10631,N_8794,N_7845);
nand U10632 (N_10632,N_9597,N_8025);
nor U10633 (N_10633,N_7837,N_9289);
xor U10634 (N_10634,N_8179,N_9427);
nor U10635 (N_10635,N_9509,N_8134);
or U10636 (N_10636,N_9209,N_8230);
or U10637 (N_10637,N_9714,N_8948);
xnor U10638 (N_10638,N_8264,N_9326);
and U10639 (N_10639,N_7682,N_8339);
nor U10640 (N_10640,N_9295,N_9309);
nor U10641 (N_10641,N_8026,N_8696);
or U10642 (N_10642,N_9077,N_8148);
nand U10643 (N_10643,N_9545,N_8261);
or U10644 (N_10644,N_9841,N_8118);
or U10645 (N_10645,N_8889,N_8902);
nand U10646 (N_10646,N_8254,N_9540);
xor U10647 (N_10647,N_7520,N_9806);
nor U10648 (N_10648,N_8641,N_8388);
nand U10649 (N_10649,N_8210,N_7631);
and U10650 (N_10650,N_7633,N_9488);
nor U10651 (N_10651,N_8857,N_7900);
or U10652 (N_10652,N_7668,N_8798);
or U10653 (N_10653,N_9912,N_8605);
nand U10654 (N_10654,N_7964,N_8839);
and U10655 (N_10655,N_8410,N_9276);
nor U10656 (N_10656,N_9465,N_9203);
nand U10657 (N_10657,N_8722,N_7789);
xnor U10658 (N_10658,N_9931,N_8511);
xnor U10659 (N_10659,N_9741,N_8263);
nand U10660 (N_10660,N_9824,N_9382);
and U10661 (N_10661,N_8805,N_8908);
xnor U10662 (N_10662,N_7566,N_9086);
nor U10663 (N_10663,N_9012,N_9712);
xor U10664 (N_10664,N_9570,N_8847);
nand U10665 (N_10665,N_9388,N_8117);
nand U10666 (N_10666,N_7851,N_8290);
nand U10667 (N_10667,N_9732,N_9747);
and U10668 (N_10668,N_9016,N_9060);
xnor U10669 (N_10669,N_8751,N_9581);
xnor U10670 (N_10670,N_7873,N_9496);
nand U10671 (N_10671,N_9542,N_7572);
nor U10672 (N_10672,N_8886,N_8903);
or U10673 (N_10673,N_9711,N_9568);
or U10674 (N_10674,N_8131,N_9969);
and U10675 (N_10675,N_9862,N_8106);
xor U10676 (N_10676,N_9303,N_9903);
xnor U10677 (N_10677,N_9680,N_7708);
nand U10678 (N_10678,N_9532,N_9461);
and U10679 (N_10679,N_8227,N_8650);
and U10680 (N_10680,N_8678,N_9921);
and U10681 (N_10681,N_8758,N_8275);
nor U10682 (N_10682,N_8377,N_9534);
xor U10683 (N_10683,N_9577,N_8614);
nand U10684 (N_10684,N_9280,N_9188);
and U10685 (N_10685,N_9444,N_9861);
xor U10686 (N_10686,N_8405,N_9503);
or U10687 (N_10687,N_9053,N_9752);
or U10688 (N_10688,N_7980,N_8517);
and U10689 (N_10689,N_8594,N_9924);
nand U10690 (N_10690,N_7780,N_8116);
nand U10691 (N_10691,N_9067,N_8446);
and U10692 (N_10692,N_8270,N_8584);
xor U10693 (N_10693,N_9988,N_9164);
nand U10694 (N_10694,N_8778,N_8862);
or U10695 (N_10695,N_9297,N_9863);
nor U10696 (N_10696,N_9642,N_8247);
and U10697 (N_10697,N_7620,N_9604);
and U10698 (N_10698,N_8473,N_8832);
nand U10699 (N_10699,N_9851,N_8962);
xor U10700 (N_10700,N_8900,N_8401);
or U10701 (N_10701,N_9137,N_9497);
and U10702 (N_10702,N_9387,N_9395);
or U10703 (N_10703,N_9915,N_8671);
and U10704 (N_10704,N_7948,N_8332);
nor U10705 (N_10705,N_7675,N_7854);
and U10706 (N_10706,N_8012,N_8887);
xnor U10707 (N_10707,N_9589,N_9003);
and U10708 (N_10708,N_7554,N_8763);
nand U10709 (N_10709,N_8086,N_9678);
or U10710 (N_10710,N_9052,N_9621);
nor U10711 (N_10711,N_8205,N_7503);
and U10712 (N_10712,N_7957,N_7978);
nor U10713 (N_10713,N_8829,N_7640);
xor U10714 (N_10714,N_7755,N_7679);
nand U10715 (N_10715,N_7710,N_8020);
and U10716 (N_10716,N_8196,N_8369);
nor U10717 (N_10717,N_7765,N_9071);
xor U10718 (N_10718,N_9036,N_7887);
nor U10719 (N_10719,N_9147,N_8244);
xnor U10720 (N_10720,N_7839,N_8077);
nor U10721 (N_10721,N_8183,N_7714);
and U10722 (N_10722,N_8109,N_8995);
xnor U10723 (N_10723,N_8248,N_8382);
and U10724 (N_10724,N_8235,N_7899);
nor U10725 (N_10725,N_9653,N_9910);
nand U10726 (N_10726,N_8177,N_9751);
xor U10727 (N_10727,N_7528,N_7739);
and U10728 (N_10728,N_7942,N_8429);
nand U10729 (N_10729,N_9629,N_8737);
nand U10730 (N_10730,N_8283,N_7727);
nand U10731 (N_10731,N_8476,N_9336);
xnor U10732 (N_10732,N_7846,N_7717);
nand U10733 (N_10733,N_7645,N_8024);
or U10734 (N_10734,N_8550,N_9923);
or U10735 (N_10735,N_8806,N_9296);
or U10736 (N_10736,N_7512,N_7868);
nor U10737 (N_10737,N_8202,N_9507);
and U10738 (N_10738,N_9027,N_8984);
and U10739 (N_10739,N_8407,N_9494);
and U10740 (N_10740,N_9787,N_8082);
xor U10741 (N_10741,N_8081,N_8089);
xnor U10742 (N_10742,N_8070,N_7530);
nand U10743 (N_10743,N_8631,N_9859);
nor U10744 (N_10744,N_8125,N_8032);
nand U10745 (N_10745,N_8356,N_8508);
nand U10746 (N_10746,N_8719,N_8145);
or U10747 (N_10747,N_7733,N_9769);
xnor U10748 (N_10748,N_8197,N_8515);
nor U10749 (N_10749,N_8068,N_9354);
or U10750 (N_10750,N_9415,N_8046);
nor U10751 (N_10751,N_7721,N_8433);
nand U10752 (N_10752,N_9954,N_7687);
nor U10753 (N_10753,N_9482,N_9856);
nand U10754 (N_10754,N_9961,N_7509);
and U10755 (N_10755,N_8912,N_9510);
and U10756 (N_10756,N_9784,N_9404);
xor U10757 (N_10757,N_9794,N_7559);
or U10758 (N_10758,N_9679,N_7547);
and U10759 (N_10759,N_8458,N_8234);
nor U10760 (N_10760,N_8836,N_9365);
nand U10761 (N_10761,N_7812,N_8190);
nand U10762 (N_10762,N_8108,N_7536);
and U10763 (N_10763,N_8856,N_8114);
nand U10764 (N_10764,N_9223,N_9551);
xnor U10765 (N_10765,N_9098,N_8483);
and U10766 (N_10766,N_8156,N_7715);
and U10767 (N_10767,N_8649,N_8419);
or U10768 (N_10768,N_8848,N_8564);
nand U10769 (N_10769,N_9569,N_9878);
nor U10770 (N_10770,N_9628,N_8304);
or U10771 (N_10771,N_9319,N_9634);
or U10772 (N_10772,N_7677,N_9180);
or U10773 (N_10773,N_8151,N_9472);
nand U10774 (N_10774,N_9655,N_8523);
and U10775 (N_10775,N_9746,N_8394);
nand U10776 (N_10776,N_9511,N_9259);
nand U10777 (N_10777,N_8786,N_8385);
xnor U10778 (N_10778,N_8742,N_9567);
xnor U10779 (N_10779,N_8976,N_9116);
nand U10780 (N_10780,N_8266,N_7952);
or U10781 (N_10781,N_9002,N_8274);
nand U10782 (N_10782,N_8957,N_8986);
or U10783 (N_10783,N_9424,N_8907);
or U10784 (N_10784,N_7859,N_9797);
nand U10785 (N_10785,N_8375,N_7599);
and U10786 (N_10786,N_8612,N_9421);
or U10787 (N_10787,N_9918,N_9300);
nor U10788 (N_10788,N_8219,N_9650);
or U10789 (N_10789,N_8939,N_8652);
nor U10790 (N_10790,N_9170,N_9038);
nand U10791 (N_10791,N_8074,N_8656);
nand U10792 (N_10792,N_8946,N_8331);
xnor U10793 (N_10793,N_8905,N_8534);
and U10794 (N_10794,N_7766,N_7888);
or U10795 (N_10795,N_8757,N_7875);
and U10796 (N_10796,N_9165,N_8311);
or U10797 (N_10797,N_7970,N_8952);
and U10798 (N_10798,N_9974,N_8333);
nand U10799 (N_10799,N_8583,N_7826);
and U10800 (N_10800,N_9733,N_9072);
or U10801 (N_10801,N_8607,N_7829);
nand U10802 (N_10802,N_8910,N_9661);
nand U10803 (N_10803,N_7743,N_9269);
and U10804 (N_10804,N_8379,N_8647);
xnor U10805 (N_10805,N_8100,N_9290);
nor U10806 (N_10806,N_9643,N_9226);
or U10807 (N_10807,N_9025,N_7711);
nand U10808 (N_10808,N_9091,N_7565);
and U10809 (N_10809,N_9881,N_9435);
and U10810 (N_10810,N_8562,N_9849);
and U10811 (N_10811,N_9566,N_9917);
and U10812 (N_10812,N_8434,N_9605);
nand U10813 (N_10813,N_8298,N_7582);
nand U10814 (N_10814,N_9979,N_9779);
and U10815 (N_10815,N_8456,N_8445);
nand U10816 (N_10816,N_8781,N_7744);
nor U10817 (N_10817,N_9977,N_8655);
and U10818 (N_10818,N_8178,N_8695);
and U10819 (N_10819,N_8253,N_7535);
or U10820 (N_10820,N_7673,N_9957);
and U10821 (N_10821,N_8225,N_9029);
and U10822 (N_10822,N_8366,N_9826);
nand U10823 (N_10823,N_9641,N_8677);
and U10824 (N_10824,N_9817,N_8073);
or U10825 (N_10825,N_8316,N_7516);
nand U10826 (N_10826,N_9468,N_8914);
xor U10827 (N_10827,N_8146,N_9463);
nor U10828 (N_10828,N_8372,N_9252);
and U10829 (N_10829,N_9842,N_8459);
and U10830 (N_10830,N_7736,N_9089);
nand U10831 (N_10831,N_9973,N_8348);
nand U10832 (N_10832,N_7879,N_9684);
nor U10833 (N_10833,N_7691,N_8236);
or U10834 (N_10834,N_7526,N_9063);
and U10835 (N_10835,N_9126,N_9648);
and U10836 (N_10836,N_9776,N_8716);
and U10837 (N_10837,N_8851,N_7702);
nor U10838 (N_10838,N_8997,N_8391);
nand U10839 (N_10839,N_8858,N_9121);
or U10840 (N_10840,N_7938,N_8759);
nand U10841 (N_10841,N_7910,N_7602);
nor U10842 (N_10842,N_9770,N_9765);
nor U10843 (N_10843,N_9139,N_9394);
and U10844 (N_10844,N_7619,N_8766);
xor U10845 (N_10845,N_9189,N_9660);
nor U10846 (N_10846,N_8861,N_9592);
or U10847 (N_10847,N_8731,N_8027);
or U10848 (N_10848,N_7720,N_8894);
nor U10849 (N_10849,N_8237,N_8055);
or U10850 (N_10850,N_9184,N_9759);
or U10851 (N_10851,N_8365,N_7591);
nand U10852 (N_10852,N_9054,N_7861);
xnor U10853 (N_10853,N_7841,N_7852);
or U10854 (N_10854,N_8317,N_8937);
xor U10855 (N_10855,N_8582,N_8620);
nor U10856 (N_10856,N_9612,N_9284);
nor U10857 (N_10857,N_7995,N_9278);
xor U10858 (N_10858,N_9870,N_9745);
xor U10859 (N_10859,N_9149,N_8551);
or U10860 (N_10860,N_7934,N_7817);
nand U10861 (N_10861,N_7937,N_9383);
or U10862 (N_10862,N_7811,N_9946);
and U10863 (N_10863,N_8185,N_8991);
nand U10864 (N_10864,N_7627,N_8579);
nand U10865 (N_10865,N_8112,N_9158);
nand U10866 (N_10866,N_7728,N_8038);
nor U10867 (N_10867,N_7504,N_7853);
nor U10868 (N_10868,N_9355,N_8714);
nor U10869 (N_10869,N_8898,N_8320);
nor U10870 (N_10870,N_9707,N_8231);
nand U10871 (N_10871,N_9477,N_8423);
and U10872 (N_10872,N_9939,N_8999);
and U10873 (N_10873,N_8919,N_8358);
xnor U10874 (N_10874,N_8565,N_9190);
nand U10875 (N_10875,N_8643,N_8130);
or U10876 (N_10876,N_8308,N_9907);
nor U10877 (N_10877,N_8859,N_9785);
and U10878 (N_10878,N_8944,N_8790);
or U10879 (N_10879,N_9263,N_8662);
or U10880 (N_10880,N_7905,N_8818);
or U10881 (N_10881,N_8061,N_8561);
and U10882 (N_10882,N_9524,N_7742);
nand U10883 (N_10883,N_8634,N_9201);
or U10884 (N_10884,N_7500,N_8398);
nor U10885 (N_10885,N_9325,N_8611);
or U10886 (N_10886,N_8428,N_9639);
and U10887 (N_10887,N_9093,N_8535);
or U10888 (N_10888,N_8051,N_8945);
xnor U10889 (N_10889,N_7784,N_9813);
nor U10890 (N_10890,N_8817,N_7650);
nand U10891 (N_10891,N_8891,N_9446);
xor U10892 (N_10892,N_8397,N_9366);
nand U10893 (N_10893,N_7676,N_9409);
or U10894 (N_10894,N_8420,N_8685);
nor U10895 (N_10895,N_9518,N_8577);
nand U10896 (N_10896,N_7697,N_9318);
xor U10897 (N_10897,N_8642,N_8104);
nor U10898 (N_10898,N_9471,N_9377);
nor U10899 (N_10899,N_8013,N_9976);
xor U10900 (N_10900,N_8820,N_7971);
and U10901 (N_10901,N_9804,N_8661);
xor U10902 (N_10902,N_8443,N_9058);
nand U10903 (N_10903,N_7560,N_7658);
and U10904 (N_10904,N_9702,N_9491);
or U10905 (N_10905,N_9375,N_9177);
xnor U10906 (N_10906,N_9583,N_9200);
nand U10907 (N_10907,N_9633,N_9682);
and U10908 (N_10908,N_9911,N_8622);
nor U10909 (N_10909,N_9611,N_8572);
and U10910 (N_10910,N_8710,N_9323);
or U10911 (N_10911,N_9379,N_8743);
and U10912 (N_10912,N_7732,N_8442);
nand U10913 (N_10913,N_9447,N_8448);
or U10914 (N_10914,N_8690,N_8489);
xor U10915 (N_10915,N_9207,N_8482);
nand U10916 (N_10916,N_8322,N_8506);
and U10917 (N_10917,N_8099,N_8193);
and U10918 (N_10918,N_7797,N_8700);
or U10919 (N_10919,N_9439,N_8004);
xnor U10920 (N_10920,N_8785,N_9212);
nor U10921 (N_10921,N_8994,N_8718);
nor U10922 (N_10922,N_9944,N_7962);
nand U10923 (N_10923,N_7807,N_9134);
and U10924 (N_10924,N_7621,N_8767);
or U10925 (N_10925,N_8619,N_7517);
xnor U10926 (N_10926,N_9019,N_7833);
xnor U10927 (N_10927,N_9533,N_8189);
xnor U10928 (N_10928,N_8169,N_9198);
nor U10929 (N_10929,N_7534,N_7987);
and U10930 (N_10930,N_8567,N_9453);
and U10931 (N_10931,N_7557,N_8588);
nor U10932 (N_10932,N_8892,N_9475);
nor U10933 (N_10933,N_7860,N_8481);
or U10934 (N_10934,N_7519,N_7514);
and U10935 (N_10935,N_8417,N_7862);
nor U10936 (N_10936,N_9220,N_9722);
nor U10937 (N_10937,N_9853,N_9221);
xor U10938 (N_10938,N_9013,N_9074);
nand U10939 (N_10939,N_9014,N_8218);
nor U10940 (N_10940,N_8327,N_8736);
or U10941 (N_10941,N_8987,N_9174);
and U10942 (N_10942,N_8503,N_7571);
and U10943 (N_10943,N_9342,N_8516);
nand U10944 (N_10944,N_8246,N_9051);
and U10945 (N_10945,N_8899,N_9304);
nand U10946 (N_10946,N_9153,N_7791);
and U10947 (N_10947,N_7734,N_9337);
xnor U10948 (N_10948,N_7639,N_7550);
xnor U10949 (N_10949,N_9272,N_9030);
nand U10950 (N_10950,N_9020,N_9963);
or U10951 (N_10951,N_9360,N_8447);
or U10952 (N_10952,N_9742,N_9397);
nand U10953 (N_10953,N_7747,N_9368);
nand U10954 (N_10954,N_8931,N_8011);
xor U10955 (N_10955,N_7564,N_7908);
nand U10956 (N_10956,N_8863,N_9673);
xor U10957 (N_10957,N_8730,N_9985);
xnor U10958 (N_10958,N_9860,N_8243);
nor U10959 (N_10959,N_9480,N_8267);
or U10960 (N_10960,N_7681,N_9417);
nand U10961 (N_10961,N_8518,N_8560);
and U10962 (N_10962,N_7949,N_8214);
nand U10963 (N_10963,N_8668,N_8770);
or U10964 (N_10964,N_9460,N_9987);
or U10965 (N_10965,N_7652,N_7583);
nand U10966 (N_10966,N_8598,N_9672);
and U10967 (N_10967,N_9555,N_8164);
or U10968 (N_10968,N_8793,N_8621);
nand U10969 (N_10969,N_8926,N_8345);
and U10970 (N_10970,N_8916,N_8028);
nor U10971 (N_10971,N_7913,N_9348);
and U10972 (N_10972,N_7892,N_7537);
xnor U10973 (N_10973,N_8325,N_7555);
nor U10974 (N_10974,N_7556,N_9310);
xor U10975 (N_10975,N_9755,N_9831);
or U10976 (N_10976,N_8982,N_9235);
and U10977 (N_10977,N_9887,N_8787);
nand U10978 (N_10978,N_9120,N_8709);
nand U10979 (N_10979,N_9343,N_8083);
or U10980 (N_10980,N_8015,N_8404);
nor U10981 (N_10981,N_8879,N_8390);
nor U10982 (N_10982,N_7843,N_8126);
and U10983 (N_10983,N_9490,N_7940);
and U10984 (N_10984,N_9968,N_9723);
nand U10985 (N_10985,N_8297,N_7707);
nor U10986 (N_10986,N_8087,N_7758);
nand U10987 (N_10987,N_8713,N_7840);
xor U10988 (N_10988,N_8472,N_8422);
nand U10989 (N_10989,N_8123,N_9846);
or U10990 (N_10990,N_8226,N_8812);
and U10991 (N_10991,N_8139,N_9588);
nor U10992 (N_10992,N_8604,N_7609);
nand U10993 (N_10993,N_7880,N_8989);
xnor U10994 (N_10994,N_8591,N_9561);
or U10995 (N_10995,N_7617,N_8833);
nand U10996 (N_10996,N_9717,N_9580);
xnor U10997 (N_10997,N_9103,N_9997);
or U10998 (N_10998,N_8287,N_9958);
xnor U10999 (N_10999,N_8915,N_8418);
nor U11000 (N_11000,N_8315,N_7901);
nor U11001 (N_11001,N_8965,N_8975);
xnor U11002 (N_11002,N_9670,N_8153);
or U11003 (N_11003,N_8300,N_8467);
nor U11004 (N_11004,N_8537,N_7604);
nand U11005 (N_11005,N_9990,N_7834);
or U11006 (N_11006,N_7585,N_9783);
nand U11007 (N_11007,N_7795,N_9893);
or U11008 (N_11008,N_7704,N_9892);
xor U11009 (N_11009,N_9970,N_7548);
nand U11010 (N_11010,N_8530,N_7872);
xnor U11011 (N_11011,N_8860,N_8048);
and U11012 (N_11012,N_9287,N_8600);
xor U11013 (N_11013,N_7844,N_7981);
nor U11014 (N_11014,N_8983,N_8413);
nor U11015 (N_11015,N_8187,N_9299);
xnor U11016 (N_11016,N_9596,N_8602);
or U11017 (N_11017,N_8184,N_9975);
or U11018 (N_11018,N_7825,N_8174);
nand U11019 (N_11019,N_7958,N_9501);
and U11020 (N_11020,N_8538,N_7771);
nand U11021 (N_11021,N_8875,N_8717);
nor U11022 (N_11022,N_8830,N_8663);
xor U11023 (N_11023,N_9807,N_8455);
xnor U11024 (N_11024,N_9317,N_7999);
xor U11025 (N_11025,N_8874,N_9037);
xor U11026 (N_11026,N_7928,N_8810);
or U11027 (N_11027,N_7573,N_7580);
and U11028 (N_11028,N_9756,N_8692);
xnor U11029 (N_11029,N_7874,N_7603);
or U11030 (N_11030,N_9919,N_8500);
nor U11031 (N_11031,N_8800,N_8571);
nor U11032 (N_11032,N_9991,N_8085);
or U11033 (N_11033,N_8578,N_9140);
nor U11034 (N_11034,N_9481,N_9676);
or U11035 (N_11035,N_9210,N_7570);
xnor U11036 (N_11036,N_7511,N_8659);
xnor U11037 (N_11037,N_8772,N_8771);
or U11038 (N_11038,N_9217,N_7634);
xnor U11039 (N_11039,N_8871,N_8869);
xor U11040 (N_11040,N_7646,N_9740);
nor U11041 (N_11041,N_9857,N_8638);
nor U11042 (N_11042,N_9692,N_8186);
nand U11043 (N_11043,N_9109,N_9185);
nand U11044 (N_11044,N_9830,N_9373);
and U11045 (N_11045,N_9835,N_8161);
or U11046 (N_11046,N_7657,N_8990);
or U11047 (N_11047,N_7916,N_7752);
and U11048 (N_11048,N_9637,N_7709);
nor U11049 (N_11049,N_9728,N_7886);
and U11050 (N_11050,N_7914,N_9734);
or U11051 (N_11051,N_8425,N_9369);
nand U11052 (N_11052,N_8485,N_7830);
or U11053 (N_11053,N_7909,N_9506);
and U11054 (N_11054,N_9744,N_9768);
nor U11055 (N_11055,N_8096,N_7663);
and U11056 (N_11056,N_8580,N_9429);
and U11057 (N_11057,N_8727,N_9876);
nor U11058 (N_11058,N_9243,N_8921);
nor U11059 (N_11059,N_7729,N_9362);
or U11060 (N_11060,N_9700,N_7967);
and U11061 (N_11061,N_8645,N_7764);
or U11062 (N_11062,N_8281,N_9320);
and U11063 (N_11063,N_8777,N_8008);
xnor U11064 (N_11064,N_7848,N_8941);
nor U11065 (N_11065,N_8639,N_8876);
xor U11066 (N_11066,N_7911,N_8593);
and U11067 (N_11067,N_8335,N_8637);
xor U11068 (N_11068,N_8528,N_9356);
xnor U11069 (N_11069,N_9805,N_9150);
or U11070 (N_11070,N_8474,N_8029);
and U11071 (N_11071,N_9135,N_7972);
and U11072 (N_11072,N_9430,N_8933);
or U11073 (N_11073,N_9959,N_8703);
xor U11074 (N_11074,N_8000,N_7622);
nand U11075 (N_11075,N_7996,N_8172);
or U11076 (N_11076,N_7881,N_9009);
nor U11077 (N_11077,N_8457,N_9928);
xor U11078 (N_11078,N_8359,N_8789);
or U11079 (N_11079,N_8843,N_8780);
and U11080 (N_11080,N_8113,N_9474);
nand U11081 (N_11081,N_8592,N_8344);
and U11082 (N_11082,N_8441,N_9039);
nor U11083 (N_11083,N_9311,N_9748);
and U11084 (N_11084,N_9248,N_9809);
nor U11085 (N_11085,N_7632,N_9548);
and U11086 (N_11086,N_8133,N_9097);
xor U11087 (N_11087,N_8432,N_7883);
or U11088 (N_11088,N_8529,N_9186);
nor U11089 (N_11089,N_8014,N_9671);
xor U11090 (N_11090,N_8318,N_9530);
and U11091 (N_11091,N_9066,N_9110);
and U11092 (N_11092,N_8993,N_8019);
xnor U11093 (N_11093,N_9934,N_8152);
nor U11094 (N_11094,N_7660,N_7595);
and U11095 (N_11095,N_8064,N_9095);
or U11096 (N_11096,N_9371,N_8258);
nand U11097 (N_11097,N_9192,N_9045);
or U11098 (N_11098,N_9208,N_8844);
nand U11099 (N_11099,N_8539,N_9543);
xnor U11100 (N_11100,N_8615,N_8166);
nor U11101 (N_11101,N_9683,N_7567);
and U11102 (N_11102,N_9196,N_7763);
nand U11103 (N_11103,N_9143,N_8566);
xor U11104 (N_11104,N_7694,N_7616);
nor U11105 (N_11105,N_9549,N_7827);
and U11106 (N_11106,N_8229,N_8252);
xor U11107 (N_11107,N_7754,N_8043);
xor U11108 (N_11108,N_9989,N_9886);
nor U11109 (N_11109,N_9434,N_9341);
xnor U11110 (N_11110,N_9844,N_9092);
xor U11111 (N_11111,N_9007,N_9584);
or U11112 (N_11112,N_8599,N_9706);
xnor U11113 (N_11113,N_9820,N_7954);
or U11114 (N_11114,N_9938,N_8062);
nor U11115 (N_11115,N_8402,N_8354);
or U11116 (N_11116,N_7774,N_9440);
nand U11117 (N_11117,N_8519,N_8361);
xnor U11118 (N_11118,N_9023,N_8765);
nand U11119 (N_11119,N_8355,N_8257);
and U11120 (N_11120,N_9591,N_8319);
xor U11121 (N_11121,N_7903,N_8884);
nand U11122 (N_11122,N_8002,N_7626);
or U11123 (N_11123,N_9646,N_8525);
nand U11124 (N_11124,N_9380,N_9937);
nor U11125 (N_11125,N_8132,N_8865);
xor U11126 (N_11126,N_9413,N_8001);
or U11127 (N_11127,N_9840,N_8568);
and U11128 (N_11128,N_8979,N_8712);
and U11129 (N_11129,N_7586,N_7976);
nand U11130 (N_11130,N_8501,N_8633);
nand U11131 (N_11131,N_9685,N_7757);
or U11132 (N_11132,N_9260,N_8368);
or U11133 (N_11133,N_8341,N_9307);
and U11134 (N_11134,N_9624,N_8510);
xnor U11135 (N_11135,N_9364,N_9119);
and U11136 (N_11136,N_9335,N_9593);
nand U11137 (N_11137,N_7501,N_8470);
nand U11138 (N_11138,N_8256,N_8799);
nand U11139 (N_11139,N_9399,N_9815);
nor U11140 (N_11140,N_9578,N_7698);
or U11141 (N_11141,N_9392,N_9096);
nor U11142 (N_11142,N_7552,N_9516);
nor U11143 (N_11143,N_8285,N_9214);
nand U11144 (N_11144,N_9802,N_8119);
xor U11145 (N_11145,N_7933,N_8740);
or U11146 (N_11146,N_8103,N_9028);
nand U11147 (N_11147,N_9719,N_8601);
nor U11148 (N_11148,N_9750,N_9940);
nor U11149 (N_11149,N_8963,N_8217);
or U11150 (N_11150,N_9782,N_9662);
nor U11151 (N_11151,N_8657,N_8380);
or U11152 (N_11152,N_9960,N_9183);
or U11153 (N_11153,N_8824,N_8175);
nand U11154 (N_11154,N_9249,N_9554);
nand U11155 (N_11155,N_8491,N_7895);
and U11156 (N_11156,N_8371,N_7979);
nand U11157 (N_11157,N_8930,N_9273);
xor U11158 (N_11158,N_7808,N_7636);
or U11159 (N_11159,N_9736,N_9173);
nor U11160 (N_11160,N_9389,N_8464);
and U11161 (N_11161,N_8901,N_9108);
or U11162 (N_11162,N_9048,N_9833);
nor U11163 (N_11163,N_7618,N_8105);
nor U11164 (N_11164,N_8060,N_8030);
xnor U11165 (N_11165,N_9076,N_9213);
nor U11166 (N_11166,N_8956,N_7885);
nand U11167 (N_11167,N_8734,N_8097);
or U11168 (N_11168,N_9151,N_9623);
nand U11169 (N_11169,N_9749,N_8754);
xor U11170 (N_11170,N_9329,N_9128);
xnor U11171 (N_11171,N_9552,N_8305);
xnor U11172 (N_11172,N_7768,N_8654);
and U11173 (N_11173,N_9302,N_9194);
and U11174 (N_11174,N_9627,N_7767);
nor U11175 (N_11175,N_8370,N_9868);
or U11176 (N_11176,N_9796,N_9871);
nor U11177 (N_11177,N_8408,N_8392);
and U11178 (N_11178,N_8167,N_9531);
nor U11179 (N_11179,N_8194,N_9327);
or U11180 (N_11180,N_9644,N_9594);
nand U11181 (N_11181,N_8206,N_8868);
xor U11182 (N_11182,N_9374,N_8265);
nor U11183 (N_11183,N_8721,N_8797);
or U11184 (N_11184,N_8669,N_8813);
or U11185 (N_11185,N_8157,N_9129);
xnor U11186 (N_11186,N_8691,N_9331);
or U11187 (N_11187,N_8215,N_9043);
and U11188 (N_11188,N_8307,N_8814);
xor U11189 (N_11189,N_7902,N_9669);
nand U11190 (N_11190,N_8877,N_9760);
nand U11191 (N_11191,N_9261,N_9858);
nor U11192 (N_11192,N_8629,N_8699);
nand U11193 (N_11193,N_8309,N_9218);
or U11194 (N_11194,N_8504,N_9376);
or U11195 (N_11195,N_8052,N_7601);
nor U11196 (N_11196,N_8362,N_8815);
xnor U11197 (N_11197,N_8110,N_9788);
and U11198 (N_11198,N_9416,N_9358);
xor U11199 (N_11199,N_8084,N_9704);
xnor U11200 (N_11200,N_8115,N_7760);
or U11201 (N_11201,N_9107,N_9927);
xor U11202 (N_11202,N_9470,N_9823);
or U11203 (N_11203,N_9451,N_8149);
or U11204 (N_11204,N_8918,N_9951);
nor U11205 (N_11205,N_8893,N_8840);
or U11206 (N_11206,N_7882,N_9539);
or U11207 (N_11207,N_9777,N_8970);
nor U11208 (N_11208,N_7819,N_8288);
xnor U11209 (N_11209,N_8752,N_9808);
xnor U11210 (N_11210,N_9017,N_8541);
xor U11211 (N_11211,N_8367,N_9630);
xor U11212 (N_11212,N_8665,N_8475);
nor U11213 (N_11213,N_9257,N_8835);
and U11214 (N_11214,N_8289,N_9111);
or U11215 (N_11215,N_8526,N_8557);
and U11216 (N_11216,N_8724,N_8953);
and U11217 (N_11217,N_7823,N_9423);
nand U11218 (N_11218,N_9909,N_9602);
nor U11219 (N_11219,N_7568,N_7686);
or U11220 (N_11220,N_9528,N_8195);
or U11221 (N_11221,N_7877,N_8360);
nor U11222 (N_11222,N_7596,N_8574);
and U11223 (N_11223,N_9245,N_8980);
and U11224 (N_11224,N_7523,N_7968);
nor U11225 (N_11225,N_7723,N_8782);
nor U11226 (N_11226,N_7611,N_8414);
nand U11227 (N_11227,N_9041,N_8940);
xnor U11228 (N_11228,N_9557,N_7932);
nand U11229 (N_11229,N_7831,N_9059);
xor U11230 (N_11230,N_8212,N_9843);
nor U11231 (N_11231,N_9829,N_9647);
xnor U11232 (N_11232,N_9885,N_8349);
nor U11233 (N_11233,N_8094,N_8888);
nor U11234 (N_11234,N_7778,N_8558);
or U11235 (N_11235,N_9234,N_8054);
xor U11236 (N_11236,N_8636,N_8039);
or U11237 (N_11237,N_9727,N_8255);
xnor U11238 (N_11238,N_8687,N_8942);
nand U11239 (N_11239,N_8972,N_7579);
xor U11240 (N_11240,N_9308,N_7822);
and U11241 (N_11241,N_7904,N_7927);
or U11242 (N_11242,N_8324,N_9608);
xnor U11243 (N_11243,N_9879,N_8346);
nand U11244 (N_11244,N_9242,N_9363);
nand U11245 (N_11245,N_7726,N_8635);
nor U11246 (N_11246,N_9182,N_7974);
nand U11247 (N_11247,N_8581,N_9688);
nor U11248 (N_11248,N_7929,N_9636);
or U11249 (N_11249,N_9031,N_7930);
nor U11250 (N_11250,N_7828,N_9910);
or U11251 (N_11251,N_8373,N_9910);
and U11252 (N_11252,N_9709,N_7808);
xor U11253 (N_11253,N_9295,N_8675);
nand U11254 (N_11254,N_9378,N_8973);
nor U11255 (N_11255,N_8064,N_8703);
nand U11256 (N_11256,N_8905,N_9561);
nor U11257 (N_11257,N_7650,N_8144);
xnor U11258 (N_11258,N_9086,N_9560);
xnor U11259 (N_11259,N_8294,N_7919);
nor U11260 (N_11260,N_7932,N_8606);
xnor U11261 (N_11261,N_9824,N_8894);
nand U11262 (N_11262,N_9984,N_8900);
nor U11263 (N_11263,N_9844,N_8588);
xor U11264 (N_11264,N_8150,N_9791);
or U11265 (N_11265,N_7767,N_9314);
or U11266 (N_11266,N_9448,N_9425);
xnor U11267 (N_11267,N_8465,N_8361);
or U11268 (N_11268,N_7935,N_8599);
or U11269 (N_11269,N_7818,N_7582);
or U11270 (N_11270,N_7980,N_9520);
nand U11271 (N_11271,N_8521,N_9181);
or U11272 (N_11272,N_9157,N_9293);
or U11273 (N_11273,N_8951,N_9450);
xnor U11274 (N_11274,N_9104,N_9034);
or U11275 (N_11275,N_8858,N_9533);
and U11276 (N_11276,N_8563,N_9570);
nand U11277 (N_11277,N_8166,N_8957);
nand U11278 (N_11278,N_9277,N_9117);
or U11279 (N_11279,N_8115,N_9282);
and U11280 (N_11280,N_8067,N_9077);
nor U11281 (N_11281,N_9971,N_8585);
nand U11282 (N_11282,N_8833,N_7779);
nand U11283 (N_11283,N_8860,N_8059);
or U11284 (N_11284,N_8947,N_9672);
or U11285 (N_11285,N_9473,N_9132);
nand U11286 (N_11286,N_8748,N_8871);
nand U11287 (N_11287,N_8823,N_8663);
or U11288 (N_11288,N_7843,N_9467);
xor U11289 (N_11289,N_7582,N_9492);
or U11290 (N_11290,N_7625,N_8466);
xor U11291 (N_11291,N_7936,N_7878);
nor U11292 (N_11292,N_7654,N_7607);
or U11293 (N_11293,N_8360,N_9864);
xnor U11294 (N_11294,N_9918,N_8814);
xnor U11295 (N_11295,N_8111,N_9945);
xnor U11296 (N_11296,N_9374,N_8184);
xnor U11297 (N_11297,N_9088,N_8905);
nor U11298 (N_11298,N_7738,N_8283);
xnor U11299 (N_11299,N_8278,N_9794);
or U11300 (N_11300,N_7820,N_9778);
nor U11301 (N_11301,N_9629,N_8581);
or U11302 (N_11302,N_8865,N_8364);
nor U11303 (N_11303,N_8087,N_8750);
and U11304 (N_11304,N_8476,N_8009);
or U11305 (N_11305,N_7842,N_9979);
or U11306 (N_11306,N_9568,N_8185);
and U11307 (N_11307,N_8668,N_7762);
nand U11308 (N_11308,N_9333,N_7981);
nand U11309 (N_11309,N_7822,N_8842);
nand U11310 (N_11310,N_7860,N_8876);
and U11311 (N_11311,N_9767,N_7918);
and U11312 (N_11312,N_8622,N_8492);
nand U11313 (N_11313,N_9179,N_8055);
nand U11314 (N_11314,N_8132,N_8289);
and U11315 (N_11315,N_7636,N_8406);
nand U11316 (N_11316,N_8746,N_8807);
nor U11317 (N_11317,N_9192,N_7582);
nor U11318 (N_11318,N_9311,N_8052);
or U11319 (N_11319,N_9460,N_8850);
xnor U11320 (N_11320,N_9970,N_7529);
nand U11321 (N_11321,N_7878,N_9933);
or U11322 (N_11322,N_7614,N_8589);
and U11323 (N_11323,N_8060,N_8502);
or U11324 (N_11324,N_9080,N_8933);
xnor U11325 (N_11325,N_8302,N_9897);
nor U11326 (N_11326,N_7821,N_9387);
nor U11327 (N_11327,N_8732,N_9842);
nor U11328 (N_11328,N_7826,N_9708);
nand U11329 (N_11329,N_9582,N_8751);
or U11330 (N_11330,N_8171,N_9459);
nor U11331 (N_11331,N_9723,N_8160);
or U11332 (N_11332,N_8616,N_7556);
or U11333 (N_11333,N_8201,N_9012);
or U11334 (N_11334,N_7765,N_8667);
or U11335 (N_11335,N_9555,N_8551);
nor U11336 (N_11336,N_7943,N_9645);
and U11337 (N_11337,N_8230,N_9203);
nand U11338 (N_11338,N_7944,N_9218);
nor U11339 (N_11339,N_9135,N_8291);
or U11340 (N_11340,N_8166,N_9397);
nor U11341 (N_11341,N_7523,N_8928);
and U11342 (N_11342,N_8657,N_8820);
nor U11343 (N_11343,N_8704,N_9288);
and U11344 (N_11344,N_8653,N_9981);
and U11345 (N_11345,N_8689,N_8440);
nand U11346 (N_11346,N_8208,N_8851);
nand U11347 (N_11347,N_8945,N_9399);
and U11348 (N_11348,N_9138,N_9531);
nand U11349 (N_11349,N_9090,N_9610);
nor U11350 (N_11350,N_7875,N_9073);
nor U11351 (N_11351,N_7687,N_8180);
xor U11352 (N_11352,N_9582,N_8934);
or U11353 (N_11353,N_9836,N_9822);
nor U11354 (N_11354,N_9269,N_8632);
and U11355 (N_11355,N_9190,N_7992);
nand U11356 (N_11356,N_9371,N_8514);
nor U11357 (N_11357,N_8694,N_8954);
nand U11358 (N_11358,N_9970,N_9259);
nand U11359 (N_11359,N_9144,N_8565);
xnor U11360 (N_11360,N_7723,N_9920);
nor U11361 (N_11361,N_7825,N_7580);
nand U11362 (N_11362,N_9689,N_9230);
nor U11363 (N_11363,N_7904,N_9017);
nor U11364 (N_11364,N_7696,N_8090);
xor U11365 (N_11365,N_8377,N_8971);
and U11366 (N_11366,N_7576,N_9891);
or U11367 (N_11367,N_9364,N_7548);
xnor U11368 (N_11368,N_9163,N_8499);
and U11369 (N_11369,N_9910,N_9028);
and U11370 (N_11370,N_8122,N_8322);
xor U11371 (N_11371,N_9529,N_8812);
and U11372 (N_11372,N_8094,N_9147);
nand U11373 (N_11373,N_8492,N_9178);
or U11374 (N_11374,N_7694,N_8452);
xor U11375 (N_11375,N_7616,N_9277);
nor U11376 (N_11376,N_9084,N_9512);
nor U11377 (N_11377,N_7539,N_9814);
nor U11378 (N_11378,N_9458,N_8105);
xor U11379 (N_11379,N_9449,N_9684);
and U11380 (N_11380,N_9144,N_8705);
nor U11381 (N_11381,N_8100,N_7887);
or U11382 (N_11382,N_9775,N_7871);
or U11383 (N_11383,N_8064,N_9287);
nor U11384 (N_11384,N_7941,N_8331);
xor U11385 (N_11385,N_9934,N_9302);
and U11386 (N_11386,N_9743,N_9929);
nand U11387 (N_11387,N_9897,N_8287);
xnor U11388 (N_11388,N_9101,N_9845);
and U11389 (N_11389,N_9846,N_9993);
or U11390 (N_11390,N_9722,N_9377);
or U11391 (N_11391,N_7833,N_9025);
and U11392 (N_11392,N_8385,N_8082);
and U11393 (N_11393,N_9004,N_8377);
and U11394 (N_11394,N_8430,N_8071);
nor U11395 (N_11395,N_8537,N_9482);
xor U11396 (N_11396,N_9654,N_9375);
nor U11397 (N_11397,N_8421,N_8971);
nor U11398 (N_11398,N_9346,N_8498);
xnor U11399 (N_11399,N_9650,N_9555);
nor U11400 (N_11400,N_8199,N_8944);
and U11401 (N_11401,N_7986,N_7988);
or U11402 (N_11402,N_7997,N_7780);
xor U11403 (N_11403,N_8347,N_7759);
and U11404 (N_11404,N_7602,N_9806);
and U11405 (N_11405,N_9276,N_7841);
xor U11406 (N_11406,N_7546,N_8597);
or U11407 (N_11407,N_9659,N_9463);
nand U11408 (N_11408,N_8363,N_8225);
nor U11409 (N_11409,N_9908,N_8891);
and U11410 (N_11410,N_8025,N_8902);
and U11411 (N_11411,N_7643,N_9100);
nor U11412 (N_11412,N_7984,N_9940);
or U11413 (N_11413,N_9821,N_7694);
and U11414 (N_11414,N_7957,N_8214);
xnor U11415 (N_11415,N_8323,N_7707);
nor U11416 (N_11416,N_7819,N_7827);
nor U11417 (N_11417,N_9607,N_7841);
nor U11418 (N_11418,N_7718,N_8165);
xnor U11419 (N_11419,N_9627,N_9226);
or U11420 (N_11420,N_7641,N_9943);
or U11421 (N_11421,N_7865,N_8403);
or U11422 (N_11422,N_9131,N_9663);
and U11423 (N_11423,N_9913,N_8097);
nor U11424 (N_11424,N_7517,N_9487);
xnor U11425 (N_11425,N_8315,N_9294);
or U11426 (N_11426,N_8909,N_9737);
and U11427 (N_11427,N_8958,N_8425);
nor U11428 (N_11428,N_9503,N_7823);
nor U11429 (N_11429,N_9510,N_9283);
xor U11430 (N_11430,N_7520,N_8493);
nand U11431 (N_11431,N_8813,N_7904);
nand U11432 (N_11432,N_9336,N_9295);
nor U11433 (N_11433,N_9214,N_7771);
or U11434 (N_11434,N_7996,N_8524);
xor U11435 (N_11435,N_9309,N_7895);
xor U11436 (N_11436,N_8838,N_9763);
and U11437 (N_11437,N_7821,N_9119);
nand U11438 (N_11438,N_8839,N_7873);
and U11439 (N_11439,N_8482,N_9623);
nand U11440 (N_11440,N_9130,N_8761);
nor U11441 (N_11441,N_7507,N_9074);
nand U11442 (N_11442,N_8449,N_8006);
nor U11443 (N_11443,N_8656,N_9105);
xnor U11444 (N_11444,N_8440,N_7929);
nor U11445 (N_11445,N_7783,N_9085);
nand U11446 (N_11446,N_9701,N_9650);
nor U11447 (N_11447,N_8616,N_7647);
or U11448 (N_11448,N_8506,N_8121);
nand U11449 (N_11449,N_8574,N_8890);
or U11450 (N_11450,N_9010,N_8902);
nand U11451 (N_11451,N_9189,N_9628);
or U11452 (N_11452,N_8232,N_8546);
or U11453 (N_11453,N_7533,N_7523);
nand U11454 (N_11454,N_7825,N_8532);
nor U11455 (N_11455,N_9817,N_9366);
xor U11456 (N_11456,N_8514,N_9903);
or U11457 (N_11457,N_8801,N_8558);
nor U11458 (N_11458,N_9769,N_9679);
xnor U11459 (N_11459,N_9746,N_9867);
and U11460 (N_11460,N_8076,N_9245);
and U11461 (N_11461,N_8867,N_8434);
and U11462 (N_11462,N_9562,N_9824);
or U11463 (N_11463,N_9298,N_9525);
or U11464 (N_11464,N_9174,N_7523);
nor U11465 (N_11465,N_7979,N_7922);
nor U11466 (N_11466,N_8321,N_7969);
and U11467 (N_11467,N_9744,N_8534);
nand U11468 (N_11468,N_8509,N_9559);
xor U11469 (N_11469,N_7957,N_9864);
nand U11470 (N_11470,N_8705,N_8606);
xor U11471 (N_11471,N_9272,N_7925);
xor U11472 (N_11472,N_8404,N_9616);
or U11473 (N_11473,N_8935,N_8077);
nor U11474 (N_11474,N_8253,N_7680);
xnor U11475 (N_11475,N_7961,N_9586);
nor U11476 (N_11476,N_9328,N_7579);
nor U11477 (N_11477,N_8838,N_9151);
or U11478 (N_11478,N_8881,N_8031);
or U11479 (N_11479,N_8620,N_7567);
nand U11480 (N_11480,N_8071,N_8291);
xnor U11481 (N_11481,N_7950,N_8968);
or U11482 (N_11482,N_9508,N_8368);
xor U11483 (N_11483,N_9094,N_7715);
or U11484 (N_11484,N_9640,N_8740);
nand U11485 (N_11485,N_8096,N_8328);
xnor U11486 (N_11486,N_8690,N_9763);
nand U11487 (N_11487,N_7941,N_8822);
nand U11488 (N_11488,N_7673,N_8663);
xnor U11489 (N_11489,N_9905,N_8591);
and U11490 (N_11490,N_9894,N_8088);
or U11491 (N_11491,N_8821,N_9158);
and U11492 (N_11492,N_9546,N_7682);
nor U11493 (N_11493,N_9778,N_8605);
xor U11494 (N_11494,N_8193,N_9234);
xor U11495 (N_11495,N_8178,N_9263);
and U11496 (N_11496,N_8480,N_8683);
nor U11497 (N_11497,N_9742,N_7917);
nand U11498 (N_11498,N_7675,N_8363);
and U11499 (N_11499,N_9016,N_9426);
and U11500 (N_11500,N_7647,N_9447);
and U11501 (N_11501,N_8668,N_8808);
nor U11502 (N_11502,N_8845,N_8329);
and U11503 (N_11503,N_9948,N_8405);
xnor U11504 (N_11504,N_8615,N_9049);
or U11505 (N_11505,N_8185,N_8942);
or U11506 (N_11506,N_9750,N_8658);
and U11507 (N_11507,N_8120,N_9382);
nor U11508 (N_11508,N_7743,N_8539);
nand U11509 (N_11509,N_9591,N_7620);
xnor U11510 (N_11510,N_8886,N_8944);
nor U11511 (N_11511,N_7925,N_9626);
xnor U11512 (N_11512,N_9763,N_9368);
or U11513 (N_11513,N_8948,N_7958);
and U11514 (N_11514,N_7548,N_9267);
and U11515 (N_11515,N_9268,N_8819);
or U11516 (N_11516,N_9026,N_9560);
and U11517 (N_11517,N_9247,N_9214);
nand U11518 (N_11518,N_7546,N_8683);
and U11519 (N_11519,N_8261,N_9836);
and U11520 (N_11520,N_8555,N_7802);
nand U11521 (N_11521,N_9341,N_8751);
and U11522 (N_11522,N_8559,N_9812);
and U11523 (N_11523,N_9338,N_8801);
or U11524 (N_11524,N_7804,N_8946);
nor U11525 (N_11525,N_7538,N_8031);
nor U11526 (N_11526,N_8510,N_8326);
nor U11527 (N_11527,N_9078,N_7996);
or U11528 (N_11528,N_8097,N_8401);
nor U11529 (N_11529,N_8867,N_8505);
xor U11530 (N_11530,N_8847,N_7849);
nor U11531 (N_11531,N_9553,N_8512);
nor U11532 (N_11532,N_8250,N_9789);
and U11533 (N_11533,N_9937,N_9013);
nand U11534 (N_11534,N_8025,N_9059);
nor U11535 (N_11535,N_9151,N_7733);
nand U11536 (N_11536,N_8698,N_9258);
and U11537 (N_11537,N_9048,N_7544);
nand U11538 (N_11538,N_7803,N_8642);
nand U11539 (N_11539,N_8683,N_8694);
nor U11540 (N_11540,N_7949,N_8659);
nand U11541 (N_11541,N_9161,N_7628);
nor U11542 (N_11542,N_9748,N_9894);
nor U11543 (N_11543,N_8817,N_8401);
and U11544 (N_11544,N_9309,N_7816);
or U11545 (N_11545,N_9814,N_9775);
nor U11546 (N_11546,N_8889,N_9474);
and U11547 (N_11547,N_9220,N_7793);
or U11548 (N_11548,N_9813,N_9562);
nand U11549 (N_11549,N_8101,N_9230);
nand U11550 (N_11550,N_8509,N_7552);
nor U11551 (N_11551,N_9369,N_8247);
nand U11552 (N_11552,N_7998,N_7860);
or U11553 (N_11553,N_7551,N_8710);
or U11554 (N_11554,N_8341,N_8109);
xnor U11555 (N_11555,N_9501,N_9227);
nor U11556 (N_11556,N_7539,N_7505);
or U11557 (N_11557,N_9177,N_8323);
or U11558 (N_11558,N_7657,N_8137);
nor U11559 (N_11559,N_9293,N_7905);
nor U11560 (N_11560,N_9433,N_9327);
or U11561 (N_11561,N_9069,N_9311);
and U11562 (N_11562,N_9035,N_9379);
nand U11563 (N_11563,N_8901,N_8285);
xnor U11564 (N_11564,N_8255,N_8536);
nor U11565 (N_11565,N_8712,N_8415);
or U11566 (N_11566,N_8119,N_7920);
xor U11567 (N_11567,N_9787,N_8758);
xor U11568 (N_11568,N_7915,N_8404);
nor U11569 (N_11569,N_8339,N_7554);
nor U11570 (N_11570,N_8145,N_8057);
nor U11571 (N_11571,N_8171,N_8457);
nor U11572 (N_11572,N_7757,N_9026);
nor U11573 (N_11573,N_8929,N_9720);
xor U11574 (N_11574,N_8378,N_9675);
nor U11575 (N_11575,N_8860,N_7988);
nor U11576 (N_11576,N_7785,N_9337);
nor U11577 (N_11577,N_7928,N_7754);
and U11578 (N_11578,N_9912,N_9650);
and U11579 (N_11579,N_8294,N_7946);
or U11580 (N_11580,N_9618,N_8383);
nand U11581 (N_11581,N_8405,N_8574);
nand U11582 (N_11582,N_7836,N_7626);
nor U11583 (N_11583,N_8027,N_7828);
or U11584 (N_11584,N_9470,N_9369);
or U11585 (N_11585,N_8466,N_8514);
or U11586 (N_11586,N_7635,N_9882);
or U11587 (N_11587,N_9459,N_8279);
nand U11588 (N_11588,N_7871,N_9652);
and U11589 (N_11589,N_8015,N_9861);
or U11590 (N_11590,N_8645,N_9439);
xnor U11591 (N_11591,N_8458,N_7703);
and U11592 (N_11592,N_8943,N_7581);
or U11593 (N_11593,N_8368,N_8173);
or U11594 (N_11594,N_8514,N_9899);
xor U11595 (N_11595,N_7857,N_9107);
or U11596 (N_11596,N_7909,N_8548);
or U11597 (N_11597,N_9851,N_7843);
and U11598 (N_11598,N_8911,N_7582);
and U11599 (N_11599,N_9740,N_7786);
and U11600 (N_11600,N_7748,N_9403);
and U11601 (N_11601,N_9145,N_8435);
xor U11602 (N_11602,N_9699,N_7893);
nor U11603 (N_11603,N_9146,N_8719);
xor U11604 (N_11604,N_9150,N_9966);
nand U11605 (N_11605,N_9526,N_9382);
nand U11606 (N_11606,N_9511,N_7534);
xnor U11607 (N_11607,N_8749,N_8177);
nand U11608 (N_11608,N_8008,N_8125);
and U11609 (N_11609,N_7966,N_9102);
xor U11610 (N_11610,N_9576,N_9305);
xor U11611 (N_11611,N_9144,N_8029);
xnor U11612 (N_11612,N_7507,N_7692);
or U11613 (N_11613,N_8428,N_9102);
nor U11614 (N_11614,N_7905,N_8562);
or U11615 (N_11615,N_7576,N_9041);
nand U11616 (N_11616,N_9417,N_8288);
or U11617 (N_11617,N_8143,N_7778);
and U11618 (N_11618,N_8911,N_8640);
xor U11619 (N_11619,N_8906,N_8939);
nor U11620 (N_11620,N_8615,N_9305);
xnor U11621 (N_11621,N_8471,N_9705);
xnor U11622 (N_11622,N_8472,N_7751);
or U11623 (N_11623,N_9882,N_9632);
or U11624 (N_11624,N_9826,N_7871);
nor U11625 (N_11625,N_8267,N_7906);
xor U11626 (N_11626,N_7868,N_9206);
and U11627 (N_11627,N_8925,N_7578);
or U11628 (N_11628,N_9385,N_8714);
or U11629 (N_11629,N_7897,N_9852);
nand U11630 (N_11630,N_8762,N_8989);
or U11631 (N_11631,N_7672,N_7829);
nand U11632 (N_11632,N_7983,N_8728);
nor U11633 (N_11633,N_9778,N_8980);
nor U11634 (N_11634,N_7558,N_8148);
nand U11635 (N_11635,N_9628,N_7551);
and U11636 (N_11636,N_8960,N_8585);
and U11637 (N_11637,N_7530,N_8408);
nor U11638 (N_11638,N_8790,N_7845);
xor U11639 (N_11639,N_7546,N_8344);
and U11640 (N_11640,N_8303,N_7799);
and U11641 (N_11641,N_7570,N_9163);
nor U11642 (N_11642,N_7636,N_9754);
xnor U11643 (N_11643,N_9100,N_9475);
or U11644 (N_11644,N_8924,N_9931);
or U11645 (N_11645,N_7844,N_8539);
xnor U11646 (N_11646,N_8998,N_8220);
and U11647 (N_11647,N_9444,N_9632);
or U11648 (N_11648,N_8384,N_9290);
nor U11649 (N_11649,N_9257,N_9341);
nor U11650 (N_11650,N_7724,N_8468);
or U11651 (N_11651,N_9496,N_7924);
nor U11652 (N_11652,N_9893,N_7986);
nand U11653 (N_11653,N_8713,N_7874);
and U11654 (N_11654,N_8644,N_7886);
nand U11655 (N_11655,N_8613,N_9277);
and U11656 (N_11656,N_9533,N_8112);
xnor U11657 (N_11657,N_8741,N_8745);
nand U11658 (N_11658,N_7564,N_8632);
or U11659 (N_11659,N_9440,N_9829);
xor U11660 (N_11660,N_9251,N_8190);
or U11661 (N_11661,N_9898,N_8847);
xnor U11662 (N_11662,N_9479,N_8749);
nor U11663 (N_11663,N_7966,N_9197);
xor U11664 (N_11664,N_9026,N_9996);
or U11665 (N_11665,N_8780,N_9411);
and U11666 (N_11666,N_8188,N_9497);
and U11667 (N_11667,N_9552,N_9960);
and U11668 (N_11668,N_9360,N_8207);
and U11669 (N_11669,N_8518,N_7948);
or U11670 (N_11670,N_9191,N_9105);
xnor U11671 (N_11671,N_9130,N_9187);
xnor U11672 (N_11672,N_9100,N_8612);
or U11673 (N_11673,N_8021,N_7519);
xnor U11674 (N_11674,N_8935,N_9725);
and U11675 (N_11675,N_8508,N_8398);
nor U11676 (N_11676,N_9232,N_9983);
nor U11677 (N_11677,N_9408,N_9040);
nand U11678 (N_11678,N_9833,N_9933);
or U11679 (N_11679,N_9712,N_9649);
xnor U11680 (N_11680,N_8281,N_8540);
nor U11681 (N_11681,N_9929,N_9181);
nand U11682 (N_11682,N_9390,N_8362);
or U11683 (N_11683,N_7503,N_9865);
xnor U11684 (N_11684,N_8753,N_9251);
nand U11685 (N_11685,N_7957,N_9145);
or U11686 (N_11686,N_8899,N_9932);
nor U11687 (N_11687,N_7552,N_9685);
xnor U11688 (N_11688,N_7737,N_8379);
nor U11689 (N_11689,N_9912,N_8839);
nor U11690 (N_11690,N_8245,N_8685);
nor U11691 (N_11691,N_8450,N_9415);
nand U11692 (N_11692,N_9677,N_9613);
and U11693 (N_11693,N_8733,N_8090);
nor U11694 (N_11694,N_8200,N_7778);
xnor U11695 (N_11695,N_8374,N_9400);
xnor U11696 (N_11696,N_9517,N_8842);
and U11697 (N_11697,N_8518,N_9685);
nor U11698 (N_11698,N_9412,N_7710);
xnor U11699 (N_11699,N_8478,N_9549);
xnor U11700 (N_11700,N_8722,N_7629);
nor U11701 (N_11701,N_9258,N_9727);
nor U11702 (N_11702,N_9297,N_8098);
xnor U11703 (N_11703,N_9564,N_8182);
or U11704 (N_11704,N_8539,N_9880);
nor U11705 (N_11705,N_7891,N_8486);
nand U11706 (N_11706,N_8477,N_9757);
nand U11707 (N_11707,N_8547,N_8110);
nand U11708 (N_11708,N_8984,N_8328);
nand U11709 (N_11709,N_8989,N_9317);
xnor U11710 (N_11710,N_9840,N_8599);
nand U11711 (N_11711,N_9541,N_7633);
or U11712 (N_11712,N_8200,N_9679);
or U11713 (N_11713,N_8235,N_9314);
nor U11714 (N_11714,N_9420,N_7962);
nand U11715 (N_11715,N_7928,N_9440);
xor U11716 (N_11716,N_7836,N_7592);
xor U11717 (N_11717,N_7570,N_7836);
xor U11718 (N_11718,N_9446,N_9934);
xnor U11719 (N_11719,N_9343,N_8466);
nand U11720 (N_11720,N_9657,N_9064);
xnor U11721 (N_11721,N_8402,N_9587);
xnor U11722 (N_11722,N_7575,N_9129);
nand U11723 (N_11723,N_8473,N_9032);
and U11724 (N_11724,N_9137,N_7617);
nor U11725 (N_11725,N_8187,N_9941);
nand U11726 (N_11726,N_8082,N_9823);
nand U11727 (N_11727,N_8662,N_9971);
or U11728 (N_11728,N_8563,N_9651);
xnor U11729 (N_11729,N_7728,N_9287);
or U11730 (N_11730,N_7824,N_8079);
or U11731 (N_11731,N_8941,N_9849);
nor U11732 (N_11732,N_7906,N_7893);
nand U11733 (N_11733,N_7839,N_9332);
nor U11734 (N_11734,N_9803,N_8511);
or U11735 (N_11735,N_9168,N_7668);
xor U11736 (N_11736,N_8470,N_9015);
nand U11737 (N_11737,N_7821,N_9030);
nor U11738 (N_11738,N_8157,N_9202);
xor U11739 (N_11739,N_9648,N_7928);
and U11740 (N_11740,N_9212,N_9528);
or U11741 (N_11741,N_9692,N_9477);
xor U11742 (N_11742,N_8478,N_8424);
and U11743 (N_11743,N_8291,N_7539);
xor U11744 (N_11744,N_8513,N_9464);
nor U11745 (N_11745,N_9589,N_8792);
xor U11746 (N_11746,N_8970,N_8324);
xor U11747 (N_11747,N_8150,N_8924);
nand U11748 (N_11748,N_9239,N_8292);
xnor U11749 (N_11749,N_7942,N_9553);
xnor U11750 (N_11750,N_7678,N_8666);
or U11751 (N_11751,N_8183,N_7699);
or U11752 (N_11752,N_7510,N_7900);
and U11753 (N_11753,N_8493,N_9720);
xnor U11754 (N_11754,N_9456,N_9244);
and U11755 (N_11755,N_7513,N_8154);
and U11756 (N_11756,N_8323,N_7732);
and U11757 (N_11757,N_7508,N_9166);
xor U11758 (N_11758,N_9954,N_8360);
nand U11759 (N_11759,N_8081,N_9875);
nand U11760 (N_11760,N_8006,N_7918);
and U11761 (N_11761,N_8785,N_9696);
nand U11762 (N_11762,N_9262,N_8791);
nand U11763 (N_11763,N_8233,N_8082);
and U11764 (N_11764,N_8010,N_8536);
and U11765 (N_11765,N_9777,N_7882);
nor U11766 (N_11766,N_8840,N_9084);
nor U11767 (N_11767,N_9711,N_8648);
and U11768 (N_11768,N_8965,N_9009);
or U11769 (N_11769,N_9211,N_8008);
nor U11770 (N_11770,N_9701,N_7931);
nand U11771 (N_11771,N_8194,N_9560);
and U11772 (N_11772,N_8084,N_8042);
or U11773 (N_11773,N_9754,N_9939);
or U11774 (N_11774,N_9321,N_8623);
and U11775 (N_11775,N_9059,N_7808);
nand U11776 (N_11776,N_7707,N_8939);
and U11777 (N_11777,N_7582,N_8586);
xnor U11778 (N_11778,N_7502,N_9044);
nor U11779 (N_11779,N_7856,N_9236);
nor U11780 (N_11780,N_9846,N_8557);
nor U11781 (N_11781,N_7627,N_9837);
and U11782 (N_11782,N_8317,N_8668);
nor U11783 (N_11783,N_8709,N_8936);
nand U11784 (N_11784,N_8841,N_9203);
and U11785 (N_11785,N_9872,N_8211);
xnor U11786 (N_11786,N_8283,N_9948);
xnor U11787 (N_11787,N_8973,N_9262);
nand U11788 (N_11788,N_9878,N_9639);
nor U11789 (N_11789,N_8362,N_8506);
nand U11790 (N_11790,N_9308,N_9533);
nor U11791 (N_11791,N_8447,N_7779);
xnor U11792 (N_11792,N_7780,N_8222);
nor U11793 (N_11793,N_9349,N_9548);
and U11794 (N_11794,N_9381,N_9872);
nor U11795 (N_11795,N_9397,N_8548);
and U11796 (N_11796,N_7843,N_9505);
nand U11797 (N_11797,N_8267,N_8482);
nor U11798 (N_11798,N_8155,N_8238);
or U11799 (N_11799,N_7937,N_8648);
xnor U11800 (N_11800,N_8371,N_7618);
nor U11801 (N_11801,N_8050,N_9458);
or U11802 (N_11802,N_7886,N_9996);
nor U11803 (N_11803,N_9728,N_8553);
nor U11804 (N_11804,N_9618,N_9081);
or U11805 (N_11805,N_8837,N_7716);
or U11806 (N_11806,N_8036,N_8402);
nor U11807 (N_11807,N_7520,N_9918);
or U11808 (N_11808,N_8963,N_7679);
nand U11809 (N_11809,N_8773,N_9464);
or U11810 (N_11810,N_8469,N_9104);
and U11811 (N_11811,N_7665,N_9386);
and U11812 (N_11812,N_9168,N_9985);
xnor U11813 (N_11813,N_8556,N_8479);
nand U11814 (N_11814,N_8275,N_8986);
or U11815 (N_11815,N_8859,N_9976);
or U11816 (N_11816,N_8393,N_9303);
and U11817 (N_11817,N_7912,N_9615);
xnor U11818 (N_11818,N_9834,N_8130);
nand U11819 (N_11819,N_8428,N_8398);
and U11820 (N_11820,N_9689,N_8724);
nand U11821 (N_11821,N_9522,N_9816);
or U11822 (N_11822,N_9405,N_9617);
xor U11823 (N_11823,N_7860,N_8379);
and U11824 (N_11824,N_8050,N_8951);
nor U11825 (N_11825,N_9514,N_8018);
xor U11826 (N_11826,N_9284,N_8299);
nand U11827 (N_11827,N_9844,N_9498);
nor U11828 (N_11828,N_9462,N_9571);
and U11829 (N_11829,N_7858,N_8925);
or U11830 (N_11830,N_8142,N_9877);
nor U11831 (N_11831,N_7706,N_9694);
or U11832 (N_11832,N_9335,N_8260);
and U11833 (N_11833,N_7920,N_8226);
nand U11834 (N_11834,N_8235,N_8885);
and U11835 (N_11835,N_8885,N_9990);
and U11836 (N_11836,N_8866,N_8382);
or U11837 (N_11837,N_8559,N_9425);
and U11838 (N_11838,N_9103,N_9975);
xor U11839 (N_11839,N_8383,N_8827);
or U11840 (N_11840,N_9536,N_8531);
and U11841 (N_11841,N_9590,N_8761);
xor U11842 (N_11842,N_9753,N_7551);
nor U11843 (N_11843,N_9756,N_9199);
xor U11844 (N_11844,N_9157,N_9370);
nand U11845 (N_11845,N_9652,N_8590);
nand U11846 (N_11846,N_8099,N_9813);
xnor U11847 (N_11847,N_8085,N_9833);
nand U11848 (N_11848,N_7775,N_9202);
and U11849 (N_11849,N_8187,N_8269);
xnor U11850 (N_11850,N_9498,N_7605);
nand U11851 (N_11851,N_9990,N_9757);
xnor U11852 (N_11852,N_7892,N_9064);
xor U11853 (N_11853,N_7582,N_9001);
xor U11854 (N_11854,N_9007,N_7607);
nor U11855 (N_11855,N_8554,N_7998);
or U11856 (N_11856,N_8125,N_9644);
nor U11857 (N_11857,N_7783,N_9534);
nor U11858 (N_11858,N_8903,N_8795);
nand U11859 (N_11859,N_9660,N_9061);
xnor U11860 (N_11860,N_8443,N_8986);
xor U11861 (N_11861,N_7689,N_9767);
nand U11862 (N_11862,N_8224,N_8092);
nand U11863 (N_11863,N_7925,N_9208);
or U11864 (N_11864,N_9264,N_9433);
xor U11865 (N_11865,N_8695,N_7968);
nor U11866 (N_11866,N_9649,N_7820);
xnor U11867 (N_11867,N_8531,N_8555);
or U11868 (N_11868,N_8256,N_9288);
nor U11869 (N_11869,N_8362,N_8889);
xnor U11870 (N_11870,N_9587,N_9938);
or U11871 (N_11871,N_8365,N_7620);
or U11872 (N_11872,N_9152,N_9097);
nor U11873 (N_11873,N_8405,N_9558);
or U11874 (N_11874,N_7725,N_8313);
nand U11875 (N_11875,N_8832,N_9441);
nor U11876 (N_11876,N_8976,N_8050);
or U11877 (N_11877,N_7715,N_9247);
and U11878 (N_11878,N_7611,N_7663);
nor U11879 (N_11879,N_9093,N_9132);
nor U11880 (N_11880,N_9408,N_7832);
nor U11881 (N_11881,N_9933,N_8611);
nor U11882 (N_11882,N_9098,N_7635);
or U11883 (N_11883,N_9091,N_8087);
and U11884 (N_11884,N_7770,N_9504);
xnor U11885 (N_11885,N_8511,N_8066);
and U11886 (N_11886,N_8003,N_9090);
or U11887 (N_11887,N_7986,N_8800);
nor U11888 (N_11888,N_8848,N_8596);
nand U11889 (N_11889,N_8673,N_8682);
xor U11890 (N_11890,N_9603,N_9454);
and U11891 (N_11891,N_7947,N_7943);
nand U11892 (N_11892,N_9092,N_8354);
nor U11893 (N_11893,N_8769,N_7883);
nor U11894 (N_11894,N_7653,N_7886);
xor U11895 (N_11895,N_8792,N_7578);
xnor U11896 (N_11896,N_9903,N_7642);
nor U11897 (N_11897,N_8811,N_8263);
and U11898 (N_11898,N_9751,N_7661);
and U11899 (N_11899,N_8538,N_8207);
nor U11900 (N_11900,N_7586,N_9912);
xor U11901 (N_11901,N_9049,N_8942);
nor U11902 (N_11902,N_8827,N_9686);
xnor U11903 (N_11903,N_8790,N_8115);
nand U11904 (N_11904,N_7505,N_9958);
xnor U11905 (N_11905,N_9294,N_8640);
and U11906 (N_11906,N_8355,N_7738);
or U11907 (N_11907,N_7841,N_8574);
xor U11908 (N_11908,N_8383,N_7725);
or U11909 (N_11909,N_8260,N_8519);
nor U11910 (N_11910,N_8350,N_8362);
xnor U11911 (N_11911,N_8353,N_9071);
nand U11912 (N_11912,N_7624,N_7706);
or U11913 (N_11913,N_8492,N_8193);
or U11914 (N_11914,N_8739,N_8010);
xor U11915 (N_11915,N_7648,N_9414);
xnor U11916 (N_11916,N_7604,N_7709);
or U11917 (N_11917,N_8245,N_8174);
nand U11918 (N_11918,N_8228,N_7568);
and U11919 (N_11919,N_7929,N_9558);
nand U11920 (N_11920,N_8038,N_8168);
nor U11921 (N_11921,N_8866,N_9523);
nor U11922 (N_11922,N_9697,N_9008);
xor U11923 (N_11923,N_9569,N_9785);
xnor U11924 (N_11924,N_8772,N_7730);
nand U11925 (N_11925,N_8257,N_8101);
nor U11926 (N_11926,N_9664,N_8518);
or U11927 (N_11927,N_8714,N_8603);
xor U11928 (N_11928,N_8156,N_9044);
nand U11929 (N_11929,N_9753,N_8610);
xor U11930 (N_11930,N_9175,N_9324);
nand U11931 (N_11931,N_8515,N_9332);
or U11932 (N_11932,N_7736,N_8503);
and U11933 (N_11933,N_8625,N_8630);
nand U11934 (N_11934,N_7719,N_9801);
or U11935 (N_11935,N_9568,N_8976);
and U11936 (N_11936,N_7791,N_7626);
nor U11937 (N_11937,N_8150,N_8101);
or U11938 (N_11938,N_7693,N_8061);
nand U11939 (N_11939,N_7914,N_8609);
or U11940 (N_11940,N_7766,N_9961);
xnor U11941 (N_11941,N_9824,N_8317);
nand U11942 (N_11942,N_8426,N_8379);
nor U11943 (N_11943,N_8656,N_7909);
nor U11944 (N_11944,N_7532,N_8419);
or U11945 (N_11945,N_9246,N_9918);
nor U11946 (N_11946,N_8298,N_8504);
and U11947 (N_11947,N_8730,N_8903);
nor U11948 (N_11948,N_8896,N_9531);
nand U11949 (N_11949,N_9210,N_9264);
and U11950 (N_11950,N_8021,N_8665);
nor U11951 (N_11951,N_8920,N_7724);
nand U11952 (N_11952,N_7860,N_9611);
or U11953 (N_11953,N_8998,N_8897);
and U11954 (N_11954,N_9015,N_8251);
nor U11955 (N_11955,N_9275,N_9043);
nand U11956 (N_11956,N_8740,N_7726);
nand U11957 (N_11957,N_7817,N_8448);
nand U11958 (N_11958,N_9193,N_9538);
nor U11959 (N_11959,N_9694,N_9453);
or U11960 (N_11960,N_8192,N_8556);
nand U11961 (N_11961,N_8541,N_9343);
and U11962 (N_11962,N_7804,N_8575);
xor U11963 (N_11963,N_8744,N_8238);
xor U11964 (N_11964,N_9982,N_9169);
xnor U11965 (N_11965,N_8184,N_9517);
xor U11966 (N_11966,N_8447,N_7707);
xnor U11967 (N_11967,N_9836,N_7722);
xnor U11968 (N_11968,N_9878,N_9699);
or U11969 (N_11969,N_8481,N_8073);
or U11970 (N_11970,N_9362,N_9868);
nor U11971 (N_11971,N_9981,N_8332);
nor U11972 (N_11972,N_7923,N_9166);
or U11973 (N_11973,N_7814,N_9160);
and U11974 (N_11974,N_9973,N_8048);
or U11975 (N_11975,N_8815,N_8159);
nand U11976 (N_11976,N_8323,N_9524);
xor U11977 (N_11977,N_8871,N_9724);
nand U11978 (N_11978,N_9576,N_9115);
nand U11979 (N_11979,N_8767,N_7757);
and U11980 (N_11980,N_8273,N_7572);
nor U11981 (N_11981,N_8331,N_7790);
nor U11982 (N_11982,N_8580,N_8961);
or U11983 (N_11983,N_8199,N_9872);
xor U11984 (N_11984,N_9701,N_8908);
and U11985 (N_11985,N_7670,N_7518);
nand U11986 (N_11986,N_9419,N_8271);
nor U11987 (N_11987,N_8957,N_9414);
xnor U11988 (N_11988,N_8380,N_8985);
and U11989 (N_11989,N_9291,N_9333);
or U11990 (N_11990,N_9052,N_7880);
nand U11991 (N_11991,N_8796,N_9275);
xor U11992 (N_11992,N_7864,N_8023);
or U11993 (N_11993,N_9240,N_8242);
nor U11994 (N_11994,N_9648,N_8556);
nand U11995 (N_11995,N_8414,N_9322);
nor U11996 (N_11996,N_8947,N_9862);
or U11997 (N_11997,N_8926,N_8655);
or U11998 (N_11998,N_7592,N_8178);
nand U11999 (N_11999,N_9116,N_9949);
or U12000 (N_12000,N_9369,N_9438);
or U12001 (N_12001,N_8783,N_9904);
xor U12002 (N_12002,N_8704,N_8414);
xor U12003 (N_12003,N_9261,N_7794);
and U12004 (N_12004,N_7938,N_9196);
or U12005 (N_12005,N_9705,N_9353);
nor U12006 (N_12006,N_9710,N_8788);
xor U12007 (N_12007,N_9959,N_8357);
and U12008 (N_12008,N_8618,N_9726);
and U12009 (N_12009,N_9728,N_7739);
or U12010 (N_12010,N_8648,N_9330);
xnor U12011 (N_12011,N_7560,N_9635);
xnor U12012 (N_12012,N_8205,N_8396);
nor U12013 (N_12013,N_9011,N_8492);
xor U12014 (N_12014,N_8935,N_9153);
and U12015 (N_12015,N_8945,N_8300);
or U12016 (N_12016,N_8082,N_9742);
nand U12017 (N_12017,N_9425,N_8767);
nor U12018 (N_12018,N_9164,N_8007);
and U12019 (N_12019,N_9579,N_7754);
nor U12020 (N_12020,N_7809,N_7758);
xor U12021 (N_12021,N_9501,N_9995);
or U12022 (N_12022,N_8119,N_8357);
or U12023 (N_12023,N_9443,N_9903);
nand U12024 (N_12024,N_8634,N_9777);
nor U12025 (N_12025,N_7935,N_8977);
or U12026 (N_12026,N_8043,N_8659);
xor U12027 (N_12027,N_9620,N_9262);
xnor U12028 (N_12028,N_7693,N_8474);
and U12029 (N_12029,N_9951,N_9061);
xor U12030 (N_12030,N_8144,N_9917);
nand U12031 (N_12031,N_9020,N_8155);
nor U12032 (N_12032,N_9465,N_8182);
and U12033 (N_12033,N_8604,N_7989);
nand U12034 (N_12034,N_8361,N_8111);
nor U12035 (N_12035,N_8895,N_9975);
or U12036 (N_12036,N_8942,N_9174);
nand U12037 (N_12037,N_9962,N_7849);
nor U12038 (N_12038,N_9349,N_9400);
nor U12039 (N_12039,N_9641,N_8460);
and U12040 (N_12040,N_7625,N_7770);
nor U12041 (N_12041,N_9457,N_9392);
xor U12042 (N_12042,N_8258,N_9764);
and U12043 (N_12043,N_9178,N_9578);
nor U12044 (N_12044,N_8635,N_8116);
and U12045 (N_12045,N_9662,N_8390);
or U12046 (N_12046,N_9265,N_9283);
and U12047 (N_12047,N_8185,N_8451);
nand U12048 (N_12048,N_8133,N_8910);
xor U12049 (N_12049,N_8358,N_9102);
xor U12050 (N_12050,N_8401,N_8873);
nor U12051 (N_12051,N_7569,N_8039);
nor U12052 (N_12052,N_8023,N_9801);
or U12053 (N_12053,N_9610,N_8653);
or U12054 (N_12054,N_8528,N_8646);
nand U12055 (N_12055,N_9341,N_7712);
nand U12056 (N_12056,N_8613,N_8137);
nand U12057 (N_12057,N_9515,N_8857);
nor U12058 (N_12058,N_8550,N_8445);
nor U12059 (N_12059,N_9131,N_9123);
xnor U12060 (N_12060,N_9708,N_8536);
and U12061 (N_12061,N_7788,N_9536);
or U12062 (N_12062,N_8079,N_7609);
or U12063 (N_12063,N_9810,N_7654);
xor U12064 (N_12064,N_7889,N_7637);
xnor U12065 (N_12065,N_9734,N_8815);
nor U12066 (N_12066,N_8727,N_9914);
nand U12067 (N_12067,N_8497,N_8576);
and U12068 (N_12068,N_8829,N_9707);
xor U12069 (N_12069,N_8766,N_8116);
and U12070 (N_12070,N_8980,N_7584);
or U12071 (N_12071,N_7824,N_7968);
nor U12072 (N_12072,N_9851,N_9170);
nor U12073 (N_12073,N_9755,N_8997);
xor U12074 (N_12074,N_8670,N_7788);
and U12075 (N_12075,N_7827,N_8029);
nand U12076 (N_12076,N_8509,N_7566);
and U12077 (N_12077,N_9940,N_9811);
or U12078 (N_12078,N_8251,N_8044);
or U12079 (N_12079,N_8214,N_8619);
and U12080 (N_12080,N_8019,N_8786);
or U12081 (N_12081,N_8373,N_9984);
and U12082 (N_12082,N_9415,N_9884);
and U12083 (N_12083,N_9194,N_9395);
nor U12084 (N_12084,N_9605,N_7697);
xor U12085 (N_12085,N_8991,N_8774);
xnor U12086 (N_12086,N_9218,N_7971);
nor U12087 (N_12087,N_9485,N_8404);
nor U12088 (N_12088,N_7511,N_7546);
nand U12089 (N_12089,N_9828,N_8152);
xnor U12090 (N_12090,N_8833,N_7679);
xnor U12091 (N_12091,N_7921,N_8360);
xnor U12092 (N_12092,N_8937,N_9460);
and U12093 (N_12093,N_8579,N_7921);
or U12094 (N_12094,N_8637,N_9345);
xor U12095 (N_12095,N_8681,N_7949);
or U12096 (N_12096,N_9920,N_8054);
nor U12097 (N_12097,N_7861,N_9925);
xnor U12098 (N_12098,N_8750,N_9557);
and U12099 (N_12099,N_9764,N_9106);
nand U12100 (N_12100,N_9903,N_8847);
or U12101 (N_12101,N_9677,N_8622);
or U12102 (N_12102,N_8717,N_8745);
nor U12103 (N_12103,N_9053,N_9551);
nor U12104 (N_12104,N_9761,N_8662);
nand U12105 (N_12105,N_8973,N_8989);
and U12106 (N_12106,N_9558,N_8027);
or U12107 (N_12107,N_7817,N_9843);
xor U12108 (N_12108,N_9350,N_8895);
nand U12109 (N_12109,N_9172,N_8841);
or U12110 (N_12110,N_9180,N_9978);
xor U12111 (N_12111,N_8486,N_9745);
or U12112 (N_12112,N_9260,N_7915);
xnor U12113 (N_12113,N_7501,N_7807);
xor U12114 (N_12114,N_8808,N_9696);
nor U12115 (N_12115,N_9392,N_7856);
or U12116 (N_12116,N_7872,N_8709);
or U12117 (N_12117,N_8056,N_9659);
and U12118 (N_12118,N_9846,N_9036);
nor U12119 (N_12119,N_8121,N_8034);
xor U12120 (N_12120,N_9461,N_7849);
and U12121 (N_12121,N_7725,N_9193);
nor U12122 (N_12122,N_8673,N_9473);
xnor U12123 (N_12123,N_9476,N_7669);
nor U12124 (N_12124,N_9688,N_9948);
xor U12125 (N_12125,N_8364,N_9989);
nand U12126 (N_12126,N_7754,N_9920);
nor U12127 (N_12127,N_7531,N_9013);
nand U12128 (N_12128,N_8086,N_8131);
nor U12129 (N_12129,N_8022,N_8214);
and U12130 (N_12130,N_7720,N_9227);
nor U12131 (N_12131,N_8018,N_8253);
xnor U12132 (N_12132,N_8329,N_8114);
nand U12133 (N_12133,N_8509,N_8684);
nor U12134 (N_12134,N_9000,N_9970);
or U12135 (N_12135,N_8988,N_9025);
or U12136 (N_12136,N_8539,N_9181);
nor U12137 (N_12137,N_7999,N_8660);
and U12138 (N_12138,N_8433,N_7517);
nand U12139 (N_12139,N_7719,N_8287);
or U12140 (N_12140,N_9421,N_9469);
nor U12141 (N_12141,N_9714,N_9428);
xor U12142 (N_12142,N_7888,N_9168);
nor U12143 (N_12143,N_9357,N_7643);
nor U12144 (N_12144,N_8050,N_8379);
and U12145 (N_12145,N_9999,N_9374);
or U12146 (N_12146,N_7876,N_7660);
or U12147 (N_12147,N_8192,N_8356);
nand U12148 (N_12148,N_8937,N_8489);
xor U12149 (N_12149,N_9541,N_9393);
or U12150 (N_12150,N_8292,N_7914);
xnor U12151 (N_12151,N_7778,N_8077);
nand U12152 (N_12152,N_7648,N_8901);
or U12153 (N_12153,N_7631,N_9894);
and U12154 (N_12154,N_7914,N_9003);
xnor U12155 (N_12155,N_9985,N_7595);
and U12156 (N_12156,N_7705,N_7868);
xnor U12157 (N_12157,N_8554,N_8786);
or U12158 (N_12158,N_9025,N_9078);
nand U12159 (N_12159,N_7720,N_9071);
or U12160 (N_12160,N_9615,N_9921);
or U12161 (N_12161,N_7896,N_9588);
nand U12162 (N_12162,N_9270,N_7519);
and U12163 (N_12163,N_9132,N_8939);
and U12164 (N_12164,N_8691,N_8630);
or U12165 (N_12165,N_8845,N_8674);
nand U12166 (N_12166,N_9377,N_9529);
and U12167 (N_12167,N_7921,N_8995);
or U12168 (N_12168,N_8947,N_7912);
nor U12169 (N_12169,N_7887,N_9119);
nor U12170 (N_12170,N_8704,N_7637);
nand U12171 (N_12171,N_8442,N_8292);
nand U12172 (N_12172,N_8999,N_9134);
and U12173 (N_12173,N_7835,N_8075);
xnor U12174 (N_12174,N_8282,N_9694);
nand U12175 (N_12175,N_8900,N_8881);
nand U12176 (N_12176,N_8955,N_9649);
and U12177 (N_12177,N_8767,N_8277);
and U12178 (N_12178,N_7720,N_9413);
or U12179 (N_12179,N_9122,N_8994);
and U12180 (N_12180,N_8932,N_9771);
or U12181 (N_12181,N_8475,N_9520);
or U12182 (N_12182,N_8641,N_8045);
and U12183 (N_12183,N_8432,N_9208);
nand U12184 (N_12184,N_9144,N_9340);
and U12185 (N_12185,N_9118,N_8791);
nor U12186 (N_12186,N_7545,N_8139);
nand U12187 (N_12187,N_9254,N_8891);
xnor U12188 (N_12188,N_9674,N_7603);
nand U12189 (N_12189,N_9219,N_8162);
nor U12190 (N_12190,N_9136,N_8891);
xnor U12191 (N_12191,N_7588,N_7849);
and U12192 (N_12192,N_8196,N_9183);
or U12193 (N_12193,N_9758,N_9052);
and U12194 (N_12194,N_9290,N_9222);
and U12195 (N_12195,N_8016,N_9319);
or U12196 (N_12196,N_9521,N_9073);
xnor U12197 (N_12197,N_9701,N_7855);
nor U12198 (N_12198,N_8901,N_8186);
nor U12199 (N_12199,N_8708,N_8836);
nor U12200 (N_12200,N_9735,N_8620);
nand U12201 (N_12201,N_7832,N_7901);
or U12202 (N_12202,N_7791,N_7672);
xor U12203 (N_12203,N_8261,N_9452);
and U12204 (N_12204,N_8163,N_9469);
xnor U12205 (N_12205,N_8032,N_9154);
or U12206 (N_12206,N_8241,N_8725);
nand U12207 (N_12207,N_9258,N_9112);
and U12208 (N_12208,N_9438,N_8133);
nor U12209 (N_12209,N_9874,N_8247);
and U12210 (N_12210,N_8232,N_8944);
or U12211 (N_12211,N_9243,N_8894);
nand U12212 (N_12212,N_9523,N_7956);
xor U12213 (N_12213,N_9239,N_8964);
and U12214 (N_12214,N_8320,N_9295);
xnor U12215 (N_12215,N_8913,N_7700);
or U12216 (N_12216,N_7830,N_8298);
nand U12217 (N_12217,N_9213,N_8248);
nor U12218 (N_12218,N_9120,N_9341);
and U12219 (N_12219,N_7560,N_8608);
and U12220 (N_12220,N_8290,N_9073);
and U12221 (N_12221,N_8285,N_8372);
xor U12222 (N_12222,N_7631,N_7777);
or U12223 (N_12223,N_9598,N_8394);
nand U12224 (N_12224,N_8948,N_9095);
nand U12225 (N_12225,N_8919,N_9673);
and U12226 (N_12226,N_9091,N_9530);
nand U12227 (N_12227,N_8158,N_8419);
xor U12228 (N_12228,N_9309,N_9503);
or U12229 (N_12229,N_8817,N_8829);
and U12230 (N_12230,N_9847,N_9003);
or U12231 (N_12231,N_9780,N_9633);
and U12232 (N_12232,N_9915,N_9154);
nor U12233 (N_12233,N_7861,N_9262);
xnor U12234 (N_12234,N_9284,N_9224);
nand U12235 (N_12235,N_8694,N_9769);
xnor U12236 (N_12236,N_7798,N_9008);
and U12237 (N_12237,N_8215,N_8288);
or U12238 (N_12238,N_8769,N_7942);
and U12239 (N_12239,N_7717,N_7897);
or U12240 (N_12240,N_8694,N_9249);
xnor U12241 (N_12241,N_7530,N_8878);
nor U12242 (N_12242,N_8418,N_9931);
nor U12243 (N_12243,N_7938,N_8980);
and U12244 (N_12244,N_9026,N_9167);
xnor U12245 (N_12245,N_7864,N_8318);
or U12246 (N_12246,N_8345,N_7506);
nor U12247 (N_12247,N_8348,N_7899);
nand U12248 (N_12248,N_9434,N_8994);
and U12249 (N_12249,N_8973,N_9876);
nand U12250 (N_12250,N_9363,N_8164);
or U12251 (N_12251,N_9115,N_8842);
and U12252 (N_12252,N_9519,N_8291);
xnor U12253 (N_12253,N_7670,N_8565);
or U12254 (N_12254,N_8708,N_7859);
or U12255 (N_12255,N_7668,N_9945);
nand U12256 (N_12256,N_9002,N_9098);
nor U12257 (N_12257,N_9705,N_9216);
and U12258 (N_12258,N_7558,N_8692);
or U12259 (N_12259,N_7547,N_9616);
nor U12260 (N_12260,N_7599,N_9338);
xnor U12261 (N_12261,N_9777,N_8261);
nand U12262 (N_12262,N_7930,N_7680);
nand U12263 (N_12263,N_9896,N_7591);
or U12264 (N_12264,N_8654,N_8296);
xor U12265 (N_12265,N_9174,N_8876);
nand U12266 (N_12266,N_7988,N_9245);
xnor U12267 (N_12267,N_8797,N_7952);
nand U12268 (N_12268,N_7937,N_7501);
nor U12269 (N_12269,N_8204,N_9844);
nand U12270 (N_12270,N_9901,N_8219);
or U12271 (N_12271,N_8563,N_8405);
xnor U12272 (N_12272,N_8273,N_9632);
or U12273 (N_12273,N_9849,N_9010);
nand U12274 (N_12274,N_8073,N_9679);
and U12275 (N_12275,N_9035,N_7627);
and U12276 (N_12276,N_7814,N_9232);
and U12277 (N_12277,N_8110,N_9376);
nor U12278 (N_12278,N_7757,N_7624);
nand U12279 (N_12279,N_8096,N_9447);
xor U12280 (N_12280,N_7849,N_7632);
xnor U12281 (N_12281,N_9943,N_8751);
or U12282 (N_12282,N_7781,N_9609);
xor U12283 (N_12283,N_9125,N_9977);
xor U12284 (N_12284,N_9847,N_7882);
or U12285 (N_12285,N_8305,N_8788);
nand U12286 (N_12286,N_9535,N_8680);
and U12287 (N_12287,N_8245,N_9297);
and U12288 (N_12288,N_9496,N_8627);
nor U12289 (N_12289,N_9653,N_8889);
xor U12290 (N_12290,N_9724,N_8191);
nor U12291 (N_12291,N_7891,N_8111);
xnor U12292 (N_12292,N_7521,N_7614);
xor U12293 (N_12293,N_7626,N_9229);
xnor U12294 (N_12294,N_7665,N_9752);
xnor U12295 (N_12295,N_7963,N_9946);
or U12296 (N_12296,N_9387,N_7731);
and U12297 (N_12297,N_9429,N_9953);
or U12298 (N_12298,N_8736,N_9343);
and U12299 (N_12299,N_7720,N_9954);
xnor U12300 (N_12300,N_7514,N_9153);
xor U12301 (N_12301,N_7710,N_7911);
nor U12302 (N_12302,N_8662,N_8561);
nor U12303 (N_12303,N_7827,N_7732);
and U12304 (N_12304,N_8090,N_9130);
or U12305 (N_12305,N_7690,N_7847);
nor U12306 (N_12306,N_9733,N_8504);
xnor U12307 (N_12307,N_9000,N_8153);
nand U12308 (N_12308,N_8866,N_9196);
and U12309 (N_12309,N_8037,N_8539);
nor U12310 (N_12310,N_9174,N_9878);
xnor U12311 (N_12311,N_9904,N_9215);
and U12312 (N_12312,N_8844,N_9556);
and U12313 (N_12313,N_9590,N_7936);
xnor U12314 (N_12314,N_8994,N_8231);
nor U12315 (N_12315,N_9022,N_9386);
xnor U12316 (N_12316,N_8141,N_7787);
nand U12317 (N_12317,N_7545,N_9474);
xor U12318 (N_12318,N_9643,N_9634);
nor U12319 (N_12319,N_7908,N_8375);
or U12320 (N_12320,N_7873,N_9816);
and U12321 (N_12321,N_8581,N_8863);
xnor U12322 (N_12322,N_9020,N_8269);
or U12323 (N_12323,N_9436,N_9205);
xor U12324 (N_12324,N_8727,N_9592);
xor U12325 (N_12325,N_9766,N_9374);
nand U12326 (N_12326,N_9357,N_7958);
or U12327 (N_12327,N_9179,N_9304);
or U12328 (N_12328,N_8153,N_8734);
nand U12329 (N_12329,N_9473,N_8521);
nand U12330 (N_12330,N_8863,N_8886);
xor U12331 (N_12331,N_9289,N_7534);
or U12332 (N_12332,N_8490,N_9851);
xor U12333 (N_12333,N_9325,N_9452);
or U12334 (N_12334,N_9212,N_8981);
nand U12335 (N_12335,N_8585,N_8650);
nor U12336 (N_12336,N_8686,N_9255);
nor U12337 (N_12337,N_7936,N_9310);
xnor U12338 (N_12338,N_7901,N_8440);
and U12339 (N_12339,N_9678,N_7823);
nor U12340 (N_12340,N_9367,N_9686);
nand U12341 (N_12341,N_9566,N_8387);
xor U12342 (N_12342,N_8471,N_7657);
xnor U12343 (N_12343,N_9724,N_9941);
or U12344 (N_12344,N_9492,N_7603);
nor U12345 (N_12345,N_9281,N_8612);
nand U12346 (N_12346,N_9961,N_8277);
nand U12347 (N_12347,N_8655,N_9937);
and U12348 (N_12348,N_9551,N_9386);
nor U12349 (N_12349,N_7528,N_9167);
xor U12350 (N_12350,N_9302,N_7919);
and U12351 (N_12351,N_8734,N_8199);
or U12352 (N_12352,N_7579,N_7976);
nor U12353 (N_12353,N_8602,N_9531);
or U12354 (N_12354,N_9524,N_9127);
or U12355 (N_12355,N_9571,N_8803);
nand U12356 (N_12356,N_8075,N_9245);
nand U12357 (N_12357,N_8886,N_8494);
nand U12358 (N_12358,N_9977,N_7946);
or U12359 (N_12359,N_8947,N_9204);
and U12360 (N_12360,N_9089,N_7633);
nand U12361 (N_12361,N_9537,N_9066);
nand U12362 (N_12362,N_8593,N_8930);
nor U12363 (N_12363,N_8417,N_8162);
and U12364 (N_12364,N_7619,N_8407);
or U12365 (N_12365,N_9231,N_8582);
or U12366 (N_12366,N_9350,N_7817);
nor U12367 (N_12367,N_9231,N_8153);
xor U12368 (N_12368,N_8969,N_9145);
or U12369 (N_12369,N_8269,N_9472);
or U12370 (N_12370,N_9208,N_7593);
xnor U12371 (N_12371,N_7602,N_7557);
nor U12372 (N_12372,N_8541,N_7881);
or U12373 (N_12373,N_9081,N_8723);
nor U12374 (N_12374,N_9042,N_7879);
nor U12375 (N_12375,N_8449,N_8015);
nor U12376 (N_12376,N_8305,N_8632);
xnor U12377 (N_12377,N_9407,N_8784);
and U12378 (N_12378,N_8799,N_9949);
nand U12379 (N_12379,N_8227,N_8028);
nor U12380 (N_12380,N_9683,N_7884);
xnor U12381 (N_12381,N_9707,N_8227);
nand U12382 (N_12382,N_9885,N_9893);
xor U12383 (N_12383,N_9608,N_8203);
nand U12384 (N_12384,N_8951,N_9464);
nor U12385 (N_12385,N_8655,N_9494);
or U12386 (N_12386,N_9814,N_9333);
or U12387 (N_12387,N_8389,N_9871);
xnor U12388 (N_12388,N_9943,N_9336);
or U12389 (N_12389,N_8401,N_7712);
nor U12390 (N_12390,N_8545,N_7500);
xnor U12391 (N_12391,N_7898,N_8917);
nor U12392 (N_12392,N_7732,N_8251);
nor U12393 (N_12393,N_9900,N_9712);
or U12394 (N_12394,N_9783,N_9817);
nor U12395 (N_12395,N_8995,N_9185);
or U12396 (N_12396,N_9930,N_9255);
nor U12397 (N_12397,N_9297,N_9818);
and U12398 (N_12398,N_7995,N_8054);
nand U12399 (N_12399,N_9658,N_8441);
nor U12400 (N_12400,N_9104,N_9507);
and U12401 (N_12401,N_8476,N_9909);
nand U12402 (N_12402,N_8562,N_8891);
nand U12403 (N_12403,N_8766,N_9351);
nand U12404 (N_12404,N_7758,N_7690);
and U12405 (N_12405,N_8871,N_9030);
nand U12406 (N_12406,N_7590,N_8707);
nor U12407 (N_12407,N_8914,N_7830);
xnor U12408 (N_12408,N_8824,N_8197);
xnor U12409 (N_12409,N_9574,N_9292);
or U12410 (N_12410,N_9648,N_8662);
and U12411 (N_12411,N_8434,N_9530);
nor U12412 (N_12412,N_9512,N_9240);
or U12413 (N_12413,N_7989,N_9570);
and U12414 (N_12414,N_8253,N_8915);
or U12415 (N_12415,N_9435,N_9692);
nor U12416 (N_12416,N_9941,N_9072);
and U12417 (N_12417,N_8523,N_9294);
and U12418 (N_12418,N_9300,N_8169);
or U12419 (N_12419,N_9386,N_7595);
and U12420 (N_12420,N_9147,N_7663);
xnor U12421 (N_12421,N_9419,N_8124);
nand U12422 (N_12422,N_7820,N_8102);
nand U12423 (N_12423,N_8230,N_8504);
nand U12424 (N_12424,N_9658,N_8622);
nand U12425 (N_12425,N_8522,N_9355);
and U12426 (N_12426,N_7788,N_8208);
xor U12427 (N_12427,N_8288,N_8925);
xnor U12428 (N_12428,N_7914,N_7860);
or U12429 (N_12429,N_7549,N_8080);
nor U12430 (N_12430,N_9154,N_8635);
and U12431 (N_12431,N_9033,N_8682);
nor U12432 (N_12432,N_8606,N_9393);
or U12433 (N_12433,N_8355,N_8150);
xor U12434 (N_12434,N_9097,N_7763);
nand U12435 (N_12435,N_9317,N_9312);
nand U12436 (N_12436,N_9186,N_8409);
and U12437 (N_12437,N_8026,N_9686);
nand U12438 (N_12438,N_9062,N_8660);
and U12439 (N_12439,N_8249,N_7542);
xnor U12440 (N_12440,N_9856,N_9587);
or U12441 (N_12441,N_9052,N_9794);
or U12442 (N_12442,N_7616,N_8238);
xnor U12443 (N_12443,N_7630,N_9359);
nand U12444 (N_12444,N_7587,N_9922);
and U12445 (N_12445,N_9267,N_9028);
and U12446 (N_12446,N_8655,N_8519);
nand U12447 (N_12447,N_7893,N_8291);
xnor U12448 (N_12448,N_7503,N_8287);
nor U12449 (N_12449,N_8664,N_8185);
nor U12450 (N_12450,N_9739,N_7728);
nor U12451 (N_12451,N_9444,N_9524);
xnor U12452 (N_12452,N_8888,N_8643);
xnor U12453 (N_12453,N_9027,N_9129);
xnor U12454 (N_12454,N_9518,N_9494);
or U12455 (N_12455,N_8725,N_8940);
nand U12456 (N_12456,N_8002,N_9143);
nand U12457 (N_12457,N_9412,N_7592);
nand U12458 (N_12458,N_9634,N_8617);
nand U12459 (N_12459,N_7634,N_8153);
xor U12460 (N_12460,N_7977,N_8883);
xor U12461 (N_12461,N_9825,N_7922);
or U12462 (N_12462,N_9008,N_9017);
nand U12463 (N_12463,N_9619,N_9563);
nor U12464 (N_12464,N_9759,N_8862);
xor U12465 (N_12465,N_7521,N_7533);
nand U12466 (N_12466,N_9295,N_7822);
nand U12467 (N_12467,N_8415,N_7525);
or U12468 (N_12468,N_9242,N_9618);
nor U12469 (N_12469,N_9460,N_9345);
and U12470 (N_12470,N_9936,N_8481);
nand U12471 (N_12471,N_9499,N_8703);
nand U12472 (N_12472,N_7817,N_9312);
nand U12473 (N_12473,N_9385,N_9354);
nand U12474 (N_12474,N_9537,N_8095);
xnor U12475 (N_12475,N_8778,N_8233);
nand U12476 (N_12476,N_9595,N_7852);
nor U12477 (N_12477,N_8188,N_7880);
and U12478 (N_12478,N_8516,N_7791);
nor U12479 (N_12479,N_9442,N_8337);
nor U12480 (N_12480,N_9131,N_7852);
or U12481 (N_12481,N_8032,N_8925);
nand U12482 (N_12482,N_8101,N_8175);
xor U12483 (N_12483,N_9140,N_8922);
nand U12484 (N_12484,N_8690,N_9567);
or U12485 (N_12485,N_8059,N_7918);
or U12486 (N_12486,N_9321,N_9833);
or U12487 (N_12487,N_8860,N_7694);
or U12488 (N_12488,N_7581,N_9289);
and U12489 (N_12489,N_8903,N_8072);
and U12490 (N_12490,N_7911,N_9254);
nor U12491 (N_12491,N_9876,N_9441);
nand U12492 (N_12492,N_9393,N_9490);
nor U12493 (N_12493,N_8837,N_9115);
or U12494 (N_12494,N_8351,N_8159);
and U12495 (N_12495,N_8180,N_9348);
and U12496 (N_12496,N_9037,N_9492);
xor U12497 (N_12497,N_8902,N_8487);
or U12498 (N_12498,N_8589,N_8159);
nand U12499 (N_12499,N_8488,N_8180);
nand U12500 (N_12500,N_12192,N_10962);
xor U12501 (N_12501,N_10544,N_10427);
or U12502 (N_12502,N_12161,N_10285);
nand U12503 (N_12503,N_10974,N_12345);
xor U12504 (N_12504,N_10837,N_11370);
nor U12505 (N_12505,N_10841,N_12404);
nand U12506 (N_12506,N_10626,N_10937);
and U12507 (N_12507,N_11995,N_10712);
and U12508 (N_12508,N_12180,N_10481);
or U12509 (N_12509,N_11878,N_10817);
and U12510 (N_12510,N_12163,N_10905);
or U12511 (N_12511,N_11169,N_11827);
nor U12512 (N_12512,N_12314,N_12168);
and U12513 (N_12513,N_10272,N_10090);
xnor U12514 (N_12514,N_12009,N_11004);
xnor U12515 (N_12515,N_12149,N_11932);
nand U12516 (N_12516,N_11633,N_11443);
nor U12517 (N_12517,N_10849,N_12238);
nand U12518 (N_12518,N_10382,N_10401);
nand U12519 (N_12519,N_11527,N_10972);
nand U12520 (N_12520,N_10995,N_10391);
or U12521 (N_12521,N_10643,N_10915);
nor U12522 (N_12522,N_11498,N_12291);
nand U12523 (N_12523,N_11456,N_10335);
nand U12524 (N_12524,N_11027,N_10771);
nand U12525 (N_12525,N_12209,N_10977);
nand U12526 (N_12526,N_11048,N_10204);
nand U12527 (N_12527,N_10205,N_11036);
or U12528 (N_12528,N_11903,N_11729);
nor U12529 (N_12529,N_10534,N_11865);
nand U12530 (N_12530,N_11256,N_11831);
and U12531 (N_12531,N_11340,N_10321);
or U12532 (N_12532,N_12006,N_11224);
nor U12533 (N_12533,N_10092,N_10264);
nand U12534 (N_12534,N_12427,N_11246);
xor U12535 (N_12535,N_10927,N_10958);
nor U12536 (N_12536,N_12351,N_11253);
or U12537 (N_12537,N_10323,N_10994);
or U12538 (N_12538,N_10519,N_10530);
nor U12539 (N_12539,N_12164,N_11901);
and U12540 (N_12540,N_10857,N_12109);
and U12541 (N_12541,N_12011,N_10338);
nor U12542 (N_12542,N_10606,N_10408);
nor U12543 (N_12543,N_12414,N_12426);
nor U12544 (N_12544,N_11471,N_11003);
xnor U12545 (N_12545,N_10402,N_10404);
and U12546 (N_12546,N_11136,N_12331);
and U12547 (N_12547,N_12022,N_10059);
and U12548 (N_12548,N_11118,N_10767);
nor U12549 (N_12549,N_11147,N_12096);
and U12550 (N_12550,N_10322,N_12460);
or U12551 (N_12551,N_10228,N_11701);
xor U12552 (N_12552,N_11117,N_10062);
nand U12553 (N_12553,N_10441,N_12432);
nor U12554 (N_12554,N_11488,N_12289);
and U12555 (N_12555,N_11356,N_10541);
or U12556 (N_12556,N_11294,N_11089);
or U12557 (N_12557,N_12230,N_12429);
nand U12558 (N_12558,N_10475,N_11475);
and U12559 (N_12559,N_11377,N_10799);
nor U12560 (N_12560,N_12493,N_10268);
or U12561 (N_12561,N_10906,N_11751);
xnor U12562 (N_12562,N_10439,N_10991);
nand U12563 (N_12563,N_11692,N_12008);
xor U12564 (N_12564,N_10941,N_11696);
and U12565 (N_12565,N_10627,N_12339);
or U12566 (N_12566,N_10640,N_11016);
xnor U12567 (N_12567,N_10975,N_12153);
or U12568 (N_12568,N_10951,N_11053);
and U12569 (N_12569,N_12295,N_12100);
or U12570 (N_12570,N_10527,N_11190);
and U12571 (N_12571,N_10503,N_10135);
or U12572 (N_12572,N_12128,N_10457);
or U12573 (N_12573,N_12073,N_10522);
xor U12574 (N_12574,N_10850,N_10586);
nand U12575 (N_12575,N_11544,N_11474);
nor U12576 (N_12576,N_11376,N_11541);
nor U12577 (N_12577,N_11449,N_12122);
nor U12578 (N_12578,N_10003,N_11677);
xnor U12579 (N_12579,N_11510,N_12489);
xor U12580 (N_12580,N_11746,N_10732);
and U12581 (N_12581,N_10159,N_10743);
xor U12582 (N_12582,N_10924,N_11805);
xor U12583 (N_12583,N_11402,N_11905);
xnor U12584 (N_12584,N_11359,N_10956);
xnor U12585 (N_12585,N_10892,N_10146);
or U12586 (N_12586,N_12341,N_10191);
xor U12587 (N_12587,N_10115,N_11912);
nand U12588 (N_12588,N_12055,N_10446);
xor U12589 (N_12589,N_11213,N_10845);
xnor U12590 (N_12590,N_10655,N_11508);
and U12591 (N_12591,N_10178,N_12320);
nand U12592 (N_12592,N_12391,N_10355);
xnor U12593 (N_12593,N_10594,N_11121);
nand U12594 (N_12594,N_11574,N_11973);
and U12595 (N_12595,N_11790,N_10934);
xor U12596 (N_12596,N_12157,N_10445);
nor U12597 (N_12597,N_10000,N_10584);
nor U12598 (N_12598,N_11872,N_10738);
nand U12599 (N_12599,N_11941,N_11324);
or U12600 (N_12600,N_11196,N_10020);
xor U12601 (N_12601,N_11276,N_10898);
and U12602 (N_12602,N_11731,N_11697);
or U12603 (N_12603,N_12202,N_12359);
xor U12604 (N_12604,N_10317,N_11342);
nand U12605 (N_12605,N_10834,N_10625);
xor U12606 (N_12606,N_11021,N_10926);
nand U12607 (N_12607,N_11210,N_12310);
and U12608 (N_12608,N_11465,N_11580);
xnor U12609 (N_12609,N_10303,N_12348);
and U12610 (N_12610,N_11312,N_10565);
nor U12611 (N_12611,N_10981,N_10557);
nand U12612 (N_12612,N_11575,N_10410);
xnor U12613 (N_12613,N_10966,N_11817);
nor U12614 (N_12614,N_10797,N_10703);
or U12615 (N_12615,N_10374,N_11200);
xnor U12616 (N_12616,N_11166,N_10669);
xnor U12617 (N_12617,N_10583,N_11238);
or U12618 (N_12618,N_11815,N_11594);
and U12619 (N_12619,N_11587,N_11774);
and U12620 (N_12620,N_10759,N_12448);
nor U12621 (N_12621,N_12329,N_11045);
nor U12622 (N_12622,N_12290,N_12330);
xnor U12623 (N_12623,N_12455,N_10870);
nor U12624 (N_12624,N_12268,N_10592);
nor U12625 (N_12625,N_11982,N_11066);
nor U12626 (N_12626,N_11298,N_10764);
xnor U12627 (N_12627,N_11682,N_11319);
nor U12628 (N_12628,N_11000,N_11345);
or U12629 (N_12629,N_10093,N_11137);
and U12630 (N_12630,N_11430,N_11519);
or U12631 (N_12631,N_10053,N_11185);
and U12632 (N_12632,N_12378,N_11693);
and U12633 (N_12633,N_10646,N_11821);
xor U12634 (N_12634,N_10883,N_11392);
nand U12635 (N_12635,N_10591,N_10256);
and U12636 (N_12636,N_10193,N_11440);
or U12637 (N_12637,N_12032,N_12306);
or U12638 (N_12638,N_10288,N_10513);
and U12639 (N_12639,N_11404,N_10710);
nand U12640 (N_12640,N_10242,N_11031);
nand U12641 (N_12641,N_10063,N_11482);
or U12642 (N_12642,N_10478,N_10024);
or U12643 (N_12643,N_10693,N_11424);
and U12644 (N_12644,N_11030,N_11269);
and U12645 (N_12645,N_11816,N_12449);
nor U12646 (N_12646,N_12467,N_11826);
xnor U12647 (N_12647,N_12041,N_10729);
nand U12648 (N_12648,N_10495,N_10673);
nor U12649 (N_12649,N_11748,N_11933);
nor U12650 (N_12650,N_12270,N_10246);
or U12651 (N_12651,N_12000,N_11739);
nor U12652 (N_12652,N_12471,N_10498);
nor U12653 (N_12653,N_12408,N_10846);
nand U12654 (N_12654,N_12037,N_10682);
nand U12655 (N_12655,N_10946,N_11212);
and U12656 (N_12656,N_10805,N_11001);
xnor U12657 (N_12657,N_12379,N_11057);
or U12658 (N_12658,N_10525,N_11942);
xnor U12659 (N_12659,N_12043,N_11078);
or U12660 (N_12660,N_10929,N_12420);
nor U12661 (N_12661,N_12077,N_12137);
or U12662 (N_12662,N_11785,N_12014);
and U12663 (N_12663,N_12374,N_11528);
nor U12664 (N_12664,N_11565,N_12316);
and U12665 (N_12665,N_10125,N_11271);
or U12666 (N_12666,N_10529,N_10843);
xnor U12667 (N_12667,N_11151,N_10684);
nor U12668 (N_12668,N_10051,N_10449);
nand U12669 (N_12669,N_12392,N_11434);
and U12670 (N_12670,N_10091,N_10572);
or U12671 (N_12671,N_11520,N_11895);
xor U12672 (N_12672,N_10201,N_10585);
nor U12673 (N_12673,N_12187,N_11242);
nand U12674 (N_12674,N_10031,N_10595);
xor U12675 (N_12675,N_11625,N_11499);
and U12676 (N_12676,N_11503,N_10025);
or U12677 (N_12677,N_11845,N_11496);
and U12678 (N_12678,N_10145,N_12367);
or U12679 (N_12679,N_10077,N_11222);
and U12680 (N_12680,N_11038,N_11661);
nor U12681 (N_12681,N_10749,N_10459);
nand U12682 (N_12682,N_11280,N_11622);
or U12683 (N_12683,N_10605,N_12039);
or U12684 (N_12684,N_12103,N_12297);
or U12685 (N_12685,N_10177,N_10683);
nand U12686 (N_12686,N_12213,N_11698);
nor U12687 (N_12687,N_10349,N_10027);
nand U12688 (N_12688,N_10774,N_12363);
nand U12689 (N_12689,N_12305,N_11409);
and U12690 (N_12690,N_10680,N_10875);
xor U12691 (N_12691,N_10083,N_11142);
and U12692 (N_12692,N_11733,N_11258);
nand U12693 (N_12693,N_10190,N_10181);
nor U12694 (N_12694,N_10444,N_11313);
xnor U12695 (N_12695,N_11561,N_10806);
xnor U12696 (N_12696,N_11960,N_10813);
or U12697 (N_12697,N_10533,N_11109);
xnor U12698 (N_12698,N_11640,N_11623);
and U12699 (N_12699,N_10989,N_11335);
xor U12700 (N_12700,N_10762,N_10987);
and U12701 (N_12701,N_11355,N_10599);
xor U12702 (N_12702,N_11135,N_11910);
nor U12703 (N_12703,N_11427,N_12051);
nor U12704 (N_12704,N_12382,N_12070);
and U12705 (N_12705,N_11768,N_11155);
nand U12706 (N_12706,N_12015,N_12152);
and U12707 (N_12707,N_12311,N_10287);
xnor U12708 (N_12708,N_11532,N_11154);
nor U12709 (N_12709,N_10865,N_10748);
and U12710 (N_12710,N_11876,N_11349);
or U12711 (N_12711,N_10950,N_11978);
xnor U12712 (N_12712,N_11899,N_10153);
xor U12713 (N_12713,N_11128,N_10550);
xnor U12714 (N_12714,N_10688,N_10563);
nand U12715 (N_12715,N_10096,N_10065);
nor U12716 (N_12716,N_10558,N_10095);
xor U12717 (N_12717,N_10198,N_10577);
nand U12718 (N_12718,N_11922,N_11466);
xor U12719 (N_12719,N_10353,N_11350);
or U12720 (N_12720,N_11996,N_11830);
nor U12721 (N_12721,N_10483,N_12170);
or U12722 (N_12722,N_12044,N_12013);
nor U12723 (N_12723,N_12113,N_10109);
and U12724 (N_12724,N_11299,N_10456);
nand U12725 (N_12725,N_10180,N_12045);
or U12726 (N_12726,N_12249,N_10465);
xnor U12727 (N_12727,N_10227,N_10071);
nand U12728 (N_12728,N_10289,N_11523);
nand U12729 (N_12729,N_10521,N_12244);
nor U12730 (N_12730,N_11384,N_10170);
or U12731 (N_12731,N_12365,N_10809);
and U12732 (N_12732,N_10796,N_11686);
xor U12733 (N_12733,N_10293,N_11863);
xnor U12734 (N_12734,N_12127,N_10363);
or U12735 (N_12735,N_11209,N_10366);
xnor U12736 (N_12736,N_12098,N_10903);
nand U12737 (N_12737,N_11833,N_10824);
and U12738 (N_12738,N_12254,N_11795);
or U12739 (N_12739,N_12487,N_12301);
nor U12740 (N_12740,N_11789,N_11553);
and U12741 (N_12741,N_11769,N_10328);
xor U12742 (N_12742,N_10454,N_10876);
nor U12743 (N_12743,N_12352,N_11669);
or U12744 (N_12744,N_11891,N_12498);
xnor U12745 (N_12745,N_11518,N_12129);
nor U12746 (N_12746,N_11913,N_10389);
and U12747 (N_12747,N_10021,N_12346);
nor U12748 (N_12748,N_10104,N_11691);
and U12749 (N_12749,N_10394,N_10219);
or U12750 (N_12750,N_10955,N_11619);
xnor U12751 (N_12751,N_12497,N_11537);
nor U12752 (N_12752,N_11002,N_11387);
nor U12753 (N_12753,N_11047,N_12199);
nor U12754 (N_12754,N_12402,N_12206);
or U12755 (N_12755,N_10756,N_12267);
nand U12756 (N_12756,N_10467,N_10306);
or U12757 (N_12757,N_11428,N_10925);
and U12758 (N_12758,N_10343,N_12237);
nand U12759 (N_12759,N_12018,N_11127);
xnor U12760 (N_12760,N_10775,N_10420);
nand U12761 (N_12761,N_12029,N_12495);
and U12762 (N_12762,N_12056,N_12376);
or U12763 (N_12763,N_12042,N_11517);
nand U12764 (N_12764,N_11763,N_11897);
xor U12765 (N_12765,N_10788,N_12433);
or U12766 (N_12766,N_12023,N_11857);
and U12767 (N_12767,N_11399,N_12095);
or U12768 (N_12768,N_11446,N_11801);
or U12769 (N_12769,N_10836,N_12280);
and U12770 (N_12770,N_11639,N_11998);
and U12771 (N_12771,N_10199,N_10019);
or U12772 (N_12772,N_11898,N_10510);
or U12773 (N_12773,N_12371,N_11171);
nand U12774 (N_12774,N_10280,N_10336);
and U12775 (N_12775,N_11195,N_11115);
and U12776 (N_12776,N_10725,N_11522);
and U12777 (N_12777,N_12231,N_12186);
nand U12778 (N_12778,N_10696,N_12084);
xor U12779 (N_12779,N_10140,N_11317);
nor U12780 (N_12780,N_12278,N_11656);
and U12781 (N_12781,N_11039,N_10458);
and U12782 (N_12782,N_10603,N_10081);
and U12783 (N_12783,N_11495,N_10935);
nor U12784 (N_12784,N_10361,N_12441);
and U12785 (N_12785,N_11668,N_11035);
and U12786 (N_12786,N_10760,N_10918);
nand U12787 (N_12787,N_11670,N_11835);
or U12788 (N_12788,N_11076,N_10888);
nor U12789 (N_12789,N_11162,N_11175);
nor U12790 (N_12790,N_11648,N_11197);
xor U12791 (N_12791,N_10225,N_11254);
nand U12792 (N_12792,N_11358,N_10502);
nor U12793 (N_12793,N_11323,N_12340);
nor U12794 (N_12794,N_11979,N_11695);
xnor U12795 (N_12795,N_12436,N_11540);
and U12796 (N_12796,N_10874,N_11679);
or U12797 (N_12797,N_10637,N_11414);
and U12798 (N_12798,N_11717,N_10678);
nand U12799 (N_12799,N_10014,N_12454);
or U12800 (N_12800,N_11156,N_10757);
nand U12801 (N_12801,N_10447,N_11564);
xnor U12802 (N_12802,N_12021,N_12285);
nand U12803 (N_12803,N_10909,N_10562);
nand U12804 (N_12804,N_10332,N_11153);
or U12805 (N_12805,N_11724,N_10316);
and U12806 (N_12806,N_10815,N_10517);
nor U12807 (N_12807,N_10149,N_12136);
and U12808 (N_12808,N_11255,N_10150);
or U12809 (N_12809,N_11552,N_12284);
and U12810 (N_12810,N_11451,N_11094);
and U12811 (N_12811,N_11013,N_10755);
xnor U12812 (N_12812,N_11132,N_12356);
nand U12813 (N_12813,N_11019,N_12182);
or U12814 (N_12814,N_10868,N_11316);
xor U12815 (N_12815,N_11107,N_12326);
nor U12816 (N_12816,N_11861,N_10136);
or U12817 (N_12817,N_10636,N_11685);
xnor U12818 (N_12818,N_12298,N_10147);
or U12819 (N_12819,N_10384,N_10663);
xnor U12820 (N_12820,N_11892,N_11265);
and U12821 (N_12821,N_10494,N_10474);
nand U12822 (N_12822,N_10214,N_10822);
nor U12823 (N_12823,N_11660,N_11725);
nand U12824 (N_12824,N_10524,N_11164);
nand U12825 (N_12825,N_12318,N_12174);
nand U12826 (N_12826,N_10183,N_11236);
xnor U12827 (N_12827,N_11969,N_12328);
nand U12828 (N_12828,N_11951,N_12124);
and U12829 (N_12829,N_12358,N_10976);
xnor U12830 (N_12830,N_11264,N_12089);
or U12831 (N_12831,N_12160,N_10436);
xor U12832 (N_12832,N_10393,N_12333);
or U12833 (N_12833,N_12119,N_10107);
xor U12834 (N_12834,N_10443,N_10587);
nand U12835 (N_12835,N_11919,N_12303);
or U12836 (N_12836,N_10079,N_11386);
nand U12837 (N_12837,N_11848,N_12144);
nand U12838 (N_12838,N_11653,N_10294);
nor U12839 (N_12839,N_10653,N_11343);
nor U12840 (N_12840,N_10614,N_11469);
nand U12841 (N_12841,N_11773,N_10238);
and U12842 (N_12842,N_11852,N_11814);
xor U12843 (N_12843,N_11902,N_11665);
and U12844 (N_12844,N_11046,N_12405);
and U12845 (N_12845,N_11344,N_11621);
or U12846 (N_12846,N_12184,N_11082);
xor U12847 (N_12847,N_11896,N_10831);
or U12848 (N_12848,N_10549,N_11944);
and U12849 (N_12849,N_11627,N_10699);
nand U12850 (N_12850,N_10895,N_11134);
xnor U12851 (N_12851,N_10327,N_11676);
xor U12852 (N_12852,N_11923,N_10161);
nor U12853 (N_12853,N_12417,N_11320);
xnor U12854 (N_12854,N_12189,N_12300);
nand U12855 (N_12855,N_10434,N_10485);
nor U12856 (N_12856,N_12395,N_11453);
nand U12857 (N_12857,N_12196,N_10241);
nor U12858 (N_12858,N_12431,N_10821);
nor U12859 (N_12859,N_10080,N_11573);
xnor U12860 (N_12860,N_12250,N_11487);
nor U12861 (N_12861,N_10641,N_11850);
nor U12862 (N_12862,N_11473,N_11441);
nand U12863 (N_12863,N_10432,N_12377);
or U12864 (N_12864,N_10901,N_12201);
and U12865 (N_12865,N_12437,N_10858);
or U12866 (N_12866,N_12194,N_11885);
and U12867 (N_12867,N_10952,N_11823);
nand U12868 (N_12868,N_12466,N_10388);
nand U12869 (N_12869,N_11678,N_11458);
or U12870 (N_12870,N_10820,N_11521);
nand U12871 (N_12871,N_11760,N_10270);
xor U12872 (N_12872,N_10087,N_11788);
xnor U12873 (N_12873,N_11567,N_11398);
nor U12874 (N_12874,N_10016,N_12275);
xor U12875 (N_12875,N_11592,N_10254);
nor U12876 (N_12876,N_11956,N_10372);
or U12877 (N_12877,N_10015,N_10041);
nand U12878 (N_12878,N_11477,N_12010);
xor U12879 (N_12879,N_11262,N_10209);
nand U12880 (N_12880,N_10647,N_11506);
xor U12881 (N_12881,N_10308,N_12204);
and U12882 (N_12882,N_10613,N_10315);
nor U12883 (N_12883,N_10378,N_10423);
nand U12884 (N_12884,N_12114,N_11244);
xor U12885 (N_12885,N_10597,N_11855);
nor U12886 (N_12886,N_10240,N_10986);
and U12887 (N_12887,N_10596,N_10542);
and U12888 (N_12888,N_11781,N_10826);
nor U12889 (N_12889,N_11173,N_12256);
nor U12890 (N_12890,N_10493,N_10780);
and U12891 (N_12891,N_11779,N_10724);
xnor U12892 (N_12892,N_12479,N_10997);
and U12893 (N_12893,N_10554,N_10677);
or U12894 (N_12894,N_11163,N_10968);
nor U12895 (N_12895,N_11369,N_11112);
xor U12896 (N_12896,N_11413,N_10904);
xnor U12897 (N_12897,N_11217,N_10546);
xnor U12898 (N_12898,N_10999,N_10723);
xnor U12899 (N_12899,N_11934,N_10894);
and U12900 (N_12900,N_10825,N_10279);
or U12901 (N_12901,N_10480,N_10878);
nor U12902 (N_12902,N_11208,N_10257);
or U12903 (N_12903,N_11292,N_12366);
or U12904 (N_12904,N_10333,N_11796);
nand U12905 (N_12905,N_11485,N_10884);
and U12906 (N_12906,N_10919,N_11229);
and U12907 (N_12907,N_10121,N_11886);
nor U12908 (N_12908,N_10963,N_10026);
nor U12909 (N_12909,N_10944,N_11362);
and U12910 (N_12910,N_11709,N_11732);
and U12911 (N_12911,N_11906,N_10169);
nand U12912 (N_12912,N_10127,N_12336);
nor U12913 (N_12913,N_11366,N_11921);
and U12914 (N_12914,N_12218,N_10064);
nand U12915 (N_12915,N_10621,N_10660);
and U12916 (N_12916,N_11509,N_10856);
nor U12917 (N_12917,N_10973,N_10112);
xnor U12918 (N_12918,N_10103,N_10429);
or U12919 (N_12919,N_10615,N_11308);
or U12920 (N_12920,N_10216,N_10790);
nand U12921 (N_12921,N_11787,N_11338);
and U12922 (N_12922,N_10574,N_10076);
xnor U12923 (N_12923,N_11674,N_11862);
xnor U12924 (N_12924,N_11705,N_11141);
or U12925 (N_12925,N_10278,N_10218);
xor U12926 (N_12926,N_10044,N_12389);
or U12927 (N_12927,N_10305,N_11176);
and U12928 (N_12928,N_12241,N_11099);
xor U12929 (N_12929,N_11975,N_11420);
xnor U12930 (N_12930,N_11794,N_12065);
nand U12931 (N_12931,N_10740,N_10564);
and U12932 (N_12932,N_12126,N_10292);
nand U12933 (N_12933,N_11990,N_12312);
nand U12934 (N_12934,N_10033,N_11505);
and U12935 (N_12935,N_11647,N_11551);
or U12936 (N_12936,N_11828,N_10034);
nor U12937 (N_12937,N_12229,N_10661);
nor U12938 (N_12938,N_11302,N_10383);
nand U12939 (N_12939,N_11026,N_11570);
or U12940 (N_12940,N_11328,N_11871);
xor U12941 (N_12941,N_11423,N_10812);
xor U12942 (N_12942,N_12442,N_11759);
nor U12943 (N_12943,N_11558,N_11703);
nor U12944 (N_12944,N_10276,N_10399);
nor U12945 (N_12945,N_11389,N_12067);
nor U12946 (N_12946,N_11707,N_10365);
or U12947 (N_12947,N_10017,N_10560);
nor U12948 (N_12948,N_11866,N_10094);
nand U12949 (N_12949,N_11372,N_11260);
and U12950 (N_12950,N_10867,N_11309);
nor U12951 (N_12951,N_10847,N_11306);
or U12952 (N_12952,N_11820,N_10325);
nand U12953 (N_12953,N_11450,N_11401);
nor U12954 (N_12954,N_10623,N_11008);
and U12955 (N_12955,N_12381,N_12191);
nor U12956 (N_12956,N_12026,N_10460);
or U12957 (N_12957,N_10887,N_12394);
and U12958 (N_12958,N_12058,N_12421);
nand U12959 (N_12959,N_12172,N_11526);
or U12960 (N_12960,N_12458,N_10154);
or U12961 (N_12961,N_11937,N_10861);
nor U12962 (N_12962,N_11680,N_11778);
and U12963 (N_12963,N_11334,N_11613);
xor U12964 (N_12964,N_10910,N_11864);
and U12965 (N_12965,N_10221,N_10890);
nor U12966 (N_12966,N_11877,N_11938);
and U12967 (N_12967,N_10672,N_12418);
xor U12968 (N_12968,N_11267,N_11318);
and U12969 (N_12969,N_10718,N_10864);
or U12970 (N_12970,N_11727,N_10551);
or U12971 (N_12971,N_11542,N_10784);
xnor U12972 (N_12972,N_10882,N_11178);
nand U12973 (N_12973,N_10505,N_10733);
xor U12974 (N_12974,N_11161,N_11361);
or U12975 (N_12975,N_11230,N_11216);
or U12976 (N_12976,N_11189,N_10250);
xor U12977 (N_12977,N_11616,N_11069);
and U12978 (N_12978,N_11330,N_10253);
xnor U12979 (N_12979,N_12370,N_11239);
nand U12980 (N_12980,N_11270,N_12279);
nor U12981 (N_12981,N_12227,N_11314);
or U12982 (N_12982,N_11716,N_10262);
and U12983 (N_12983,N_12296,N_11783);
nand U12984 (N_12984,N_12396,N_11548);
and U12985 (N_12985,N_11832,N_11168);
and U12986 (N_12986,N_11609,N_12216);
or U12987 (N_12987,N_11672,N_11662);
and U12988 (N_12988,N_10487,N_10873);
nand U12989 (N_12989,N_11749,N_11145);
or U12990 (N_12990,N_11829,N_11743);
or U12991 (N_12991,N_10472,N_10291);
xor U12992 (N_12992,N_11278,N_12108);
and U12993 (N_12993,N_12150,N_12111);
nor U12994 (N_12994,N_12302,N_11875);
and U12995 (N_12995,N_12483,N_10961);
and U12996 (N_12996,N_10631,N_11009);
or U12997 (N_12997,N_10168,N_12415);
nand U12998 (N_12998,N_11806,N_12193);
xnor U12999 (N_12999,N_12282,N_12470);
and U13000 (N_13000,N_11263,N_12078);
xnor U13001 (N_13001,N_11963,N_10223);
and U13002 (N_13002,N_12069,N_10842);
and U13003 (N_13003,N_11654,N_10568);
xnor U13004 (N_13004,N_10984,N_10967);
xnor U13005 (N_13005,N_10581,N_10182);
nor U13006 (N_13006,N_10965,N_11588);
nand U13007 (N_13007,N_10700,N_10039);
or U13008 (N_13008,N_12491,N_11747);
xor U13009 (N_13009,N_11873,N_10649);
or U13010 (N_13010,N_10761,N_10518);
nand U13011 (N_13011,N_11231,N_10188);
or U13012 (N_13012,N_11201,N_11900);
nor U13013 (N_13013,N_11494,N_11110);
and U13014 (N_13014,N_12179,N_10360);
nor U13015 (N_13015,N_10009,N_10543);
nor U13016 (N_13016,N_11452,N_10893);
or U13017 (N_13017,N_12390,N_10398);
nand U13018 (N_13018,N_11143,N_11415);
xnor U13019 (N_13019,N_10490,N_11106);
and U13020 (N_13020,N_11954,N_10629);
and U13021 (N_13021,N_11602,N_10284);
nor U13022 (N_13022,N_11481,N_10110);
nand U13023 (N_13023,N_12490,N_11437);
nor U13024 (N_13024,N_10113,N_11139);
nor U13025 (N_13025,N_12473,N_11764);
and U13026 (N_13026,N_11233,N_10097);
nor U13027 (N_13027,N_12259,N_11931);
or U13028 (N_13028,N_11569,N_12385);
or U13029 (N_13029,N_11044,N_11080);
xor U13030 (N_13030,N_12337,N_10616);
or U13031 (N_13031,N_10172,N_11600);
or U13032 (N_13032,N_10692,N_10851);
nand U13033 (N_13033,N_10368,N_10433);
nor U13034 (N_13034,N_12355,N_10235);
and U13035 (N_13035,N_11839,N_12154);
xor U13036 (N_13036,N_11840,N_10046);
or U13037 (N_13037,N_10252,N_11974);
and U13038 (N_13038,N_11432,N_10362);
or U13039 (N_13039,N_10832,N_11012);
nor U13040 (N_13040,N_11994,N_10450);
nor U13041 (N_13041,N_11591,N_12004);
nor U13042 (N_13042,N_11063,N_12177);
and U13043 (N_13043,N_10010,N_12401);
or U13044 (N_13044,N_11611,N_11412);
or U13045 (N_13045,N_10283,N_11416);
nor U13046 (N_13046,N_10100,N_10827);
and U13047 (N_13047,N_11348,N_11191);
or U13048 (N_13048,N_12446,N_12071);
nor U13049 (N_13049,N_11367,N_11237);
nor U13050 (N_13050,N_12185,N_10705);
nor U13051 (N_13051,N_11980,N_11364);
xnor U13052 (N_13052,N_11976,N_10913);
nor U13053 (N_13053,N_12323,N_10769);
xnor U13054 (N_13054,N_11985,N_12481);
xnor U13055 (N_13055,N_11586,N_12468);
nor U13056 (N_13056,N_12064,N_11712);
and U13057 (N_13057,N_11187,N_10711);
nor U13058 (N_13058,N_10220,N_12265);
nand U13059 (N_13059,N_11463,N_10695);
and U13060 (N_13060,N_12178,N_11643);
xor U13061 (N_13061,N_11915,N_11950);
nand U13062 (N_13062,N_12159,N_10763);
nor U13063 (N_13063,N_11360,N_11890);
nor U13064 (N_13064,N_10134,N_12048);
nand U13065 (N_13065,N_10773,N_12273);
nor U13066 (N_13066,N_11113,N_10607);
and U13067 (N_13067,N_10798,N_12287);
nor U13068 (N_13068,N_12452,N_10816);
nand U13069 (N_13069,N_10415,N_11754);
xnor U13070 (N_13070,N_12307,N_11149);
or U13071 (N_13071,N_11476,N_10381);
nor U13072 (N_13072,N_12324,N_12198);
or U13073 (N_13073,N_11215,N_10290);
nand U13074 (N_13074,N_12317,N_10930);
nand U13075 (N_13075,N_11177,N_11095);
nand U13076 (N_13076,N_10497,N_11381);
and U13077 (N_13077,N_10500,N_10698);
nor U13078 (N_13078,N_10304,N_10455);
nand U13079 (N_13079,N_10208,N_10897);
or U13080 (N_13080,N_11203,N_10215);
or U13081 (N_13081,N_10744,N_11808);
nand U13082 (N_13082,N_10949,N_12384);
and U13083 (N_13083,N_11273,N_10854);
and U13084 (N_13084,N_10392,N_12012);
or U13085 (N_13085,N_10721,N_10148);
or U13086 (N_13086,N_12322,N_12243);
nor U13087 (N_13087,N_12175,N_10129);
nor U13088 (N_13088,N_12001,N_11874);
xor U13089 (N_13089,N_11630,N_10889);
and U13090 (N_13090,N_12166,N_11557);
nor U13091 (N_13091,N_12074,N_12025);
xnor U13092 (N_13092,N_11859,N_10772);
nor U13093 (N_13093,N_12017,N_10492);
nor U13094 (N_13094,N_10891,N_10770);
and U13095 (N_13095,N_10514,N_10753);
or U13096 (N_13096,N_10345,N_10708);
and U13097 (N_13097,N_10055,N_12499);
or U13098 (N_13098,N_11363,N_10390);
and U13099 (N_13099,N_10697,N_10040);
nand U13100 (N_13100,N_11072,N_11198);
xnor U13101 (N_13101,N_12173,N_11967);
xor U13102 (N_13102,N_11457,N_11448);
and U13103 (N_13103,N_11949,N_11604);
xor U13104 (N_13104,N_11084,N_10570);
nand U13105 (N_13105,N_10128,N_12220);
nand U13106 (N_13106,N_10023,N_11911);
nor U13107 (N_13107,N_10982,N_10274);
or U13108 (N_13108,N_12138,N_10013);
nor U13109 (N_13109,N_11797,N_10671);
or U13110 (N_13110,N_10160,N_11418);
nand U13111 (N_13111,N_10043,N_11462);
nor U13112 (N_13112,N_10124,N_12360);
or U13113 (N_13113,N_10126,N_10879);
and U13114 (N_13114,N_12104,N_11098);
nor U13115 (N_13115,N_10665,N_11249);
and U13116 (N_13116,N_10230,N_12257);
xnor U13117 (N_13117,N_11916,N_12107);
or U13118 (N_13118,N_12030,N_12354);
xor U13119 (N_13119,N_10604,N_11411);
and U13120 (N_13120,N_12085,N_10656);
nor U13121 (N_13121,N_12246,N_11073);
or U13122 (N_13122,N_10061,N_11433);
and U13123 (N_13123,N_10413,N_11300);
xnor U13124 (N_13124,N_10309,N_11971);
and U13125 (N_13125,N_11767,N_10471);
xor U13126 (N_13126,N_10489,N_10800);
nor U13127 (N_13127,N_12422,N_10579);
xor U13128 (N_13128,N_10237,N_10520);
or U13129 (N_13129,N_11211,N_11221);
and U13130 (N_13130,N_10157,N_10689);
nand U13131 (N_13131,N_12334,N_12288);
and U13132 (N_13132,N_11493,N_11251);
nor U13133 (N_13133,N_12357,N_11819);
xnor U13134 (N_13134,N_12133,N_10358);
nand U13135 (N_13135,N_10789,N_12286);
nand U13136 (N_13136,N_12406,N_12299);
xor U13137 (N_13137,N_10667,N_11032);
nor U13138 (N_13138,N_11993,N_10866);
nand U13139 (N_13139,N_12082,N_11043);
and U13140 (N_13140,N_12428,N_10461);
nand U13141 (N_13141,N_11791,N_11713);
nand U13142 (N_13142,N_10477,N_10556);
xnor U13143 (N_13143,N_10569,N_10202);
xor U13144 (N_13144,N_10072,N_10814);
nor U13145 (N_13145,N_12261,N_10265);
nand U13146 (N_13146,N_11920,N_11745);
nor U13147 (N_13147,N_11535,N_12207);
xor U13148 (N_13148,N_11762,N_10648);
and U13149 (N_13149,N_11158,N_10038);
nand U13150 (N_13150,N_12118,N_10375);
nand U13151 (N_13151,N_11582,N_11059);
or U13152 (N_13152,N_10783,N_11385);
and U13153 (N_13153,N_11365,N_12140);
nor U13154 (N_13154,N_11657,N_11965);
nor U13155 (N_13155,N_11543,N_10844);
or U13156 (N_13156,N_10985,N_10200);
and U13157 (N_13157,N_12158,N_10679);
or U13158 (N_13158,N_11918,N_12245);
nor U13159 (N_13159,N_12130,N_11603);
or U13160 (N_13160,N_10249,N_12383);
nor U13161 (N_13161,N_10302,N_11388);
nor U13162 (N_13162,N_10589,N_10765);
or U13163 (N_13163,N_10869,N_11650);
nand U13164 (N_13164,N_11459,N_11097);
nand U13165 (N_13165,N_10726,N_10435);
xnor U13166 (N_13166,N_10715,N_10619);
nor U13167 (N_13167,N_11436,N_10818);
nand U13168 (N_13168,N_11822,N_11310);
xnor U13169 (N_13169,N_10954,N_12239);
nor U13170 (N_13170,N_10210,N_12375);
and U13171 (N_13171,N_11777,N_11718);
xor U13172 (N_13172,N_12347,N_10932);
or U13173 (N_13173,N_11227,N_11585);
or U13174 (N_13174,N_11977,N_11287);
and U13175 (N_13175,N_10707,N_11556);
and U13176 (N_13176,N_11186,N_11578);
xnor U13177 (N_13177,N_11460,N_10612);
and U13178 (N_13178,N_11125,N_11114);
nor U13179 (N_13179,N_10828,N_12373);
or U13180 (N_13180,N_12447,N_10400);
nand U13181 (N_13181,N_10473,N_10282);
and U13182 (N_13182,N_12066,N_10269);
nand U13183 (N_13183,N_10933,N_10185);
and U13184 (N_13184,N_12434,N_12190);
nor U13185 (N_13185,N_11533,N_11086);
nand U13186 (N_13186,N_11014,N_10036);
or U13187 (N_13187,N_11470,N_11800);
xor U13188 (N_13188,N_12283,N_10588);
or U13189 (N_13189,N_10638,N_11174);
nor U13190 (N_13190,N_10642,N_11394);
nand U13191 (N_13191,N_11930,N_10681);
nor U13192 (N_13192,N_10567,N_11742);
or U13193 (N_13193,N_10785,N_11028);
nand U13194 (N_13194,N_10491,N_12195);
xor U13195 (N_13195,N_10155,N_11706);
or U13196 (N_13196,N_10448,N_10633);
and U13197 (N_13197,N_11183,N_11041);
nor U13198 (N_13198,N_11525,N_10634);
or U13199 (N_13199,N_11811,N_11658);
nor U13200 (N_13200,N_10940,N_11846);
and U13201 (N_13201,N_10632,N_10084);
nand U13202 (N_13202,N_10561,N_10781);
nand U13203 (N_13203,N_12215,N_11804);
or U13204 (N_13204,N_11626,N_11307);
or U13205 (N_13205,N_11468,N_10735);
nor U13206 (N_13206,N_12183,N_11854);
nand U13207 (N_13207,N_11034,N_11375);
xor U13208 (N_13208,N_11397,N_10691);
nor U13209 (N_13209,N_10600,N_11925);
nor U13210 (N_13210,N_11571,N_10174);
nor U13211 (N_13211,N_10469,N_11935);
xor U13212 (N_13212,N_10983,N_10747);
nor U13213 (N_13213,N_12049,N_10658);
and U13214 (N_13214,N_11807,N_11371);
or U13215 (N_13215,N_10418,N_12309);
xnor U13216 (N_13216,N_10948,N_11478);
or U13217 (N_13217,N_11252,N_12171);
nand U13218 (N_13218,N_10706,N_11547);
and U13219 (N_13219,N_10523,N_12488);
or U13220 (N_13220,N_12224,N_10819);
xor U13221 (N_13221,N_10416,N_12258);
nand U13222 (N_13222,N_11501,N_10088);
and U13223 (N_13223,N_12321,N_12399);
and U13224 (N_13224,N_11704,N_10350);
nand U13225 (N_13225,N_10552,N_10324);
xor U13226 (N_13226,N_10468,N_12143);
xor U13227 (N_13227,N_10275,N_10426);
nand U13228 (N_13228,N_11225,N_10117);
nand U13229 (N_13229,N_10938,N_12380);
or U13230 (N_13230,N_12217,N_11576);
nor U13231 (N_13231,N_11917,N_10437);
nor U13232 (N_13232,N_12027,N_11516);
nand U13233 (N_13233,N_10339,N_11884);
xnor U13234 (N_13234,N_10348,N_11179);
nand U13235 (N_13235,N_10988,N_11512);
nand U13236 (N_13236,N_12210,N_11836);
xor U13237 (N_13237,N_11380,N_11953);
nor U13238 (N_13238,N_10992,N_10142);
xor U13239 (N_13239,N_11005,N_11737);
nand U13240 (N_13240,N_11987,N_10357);
and U13241 (N_13241,N_11711,N_10602);
and U13242 (N_13242,N_10840,N_12308);
and U13243 (N_13243,N_11929,N_11962);
xnor U13244 (N_13244,N_10440,N_12062);
nand U13245 (N_13245,N_11659,N_12102);
nor U13246 (N_13246,N_10635,N_10411);
nand U13247 (N_13247,N_11802,N_11029);
and U13248 (N_13248,N_10659,N_10920);
nand U13249 (N_13249,N_10582,N_11638);
nor U13250 (N_13250,N_10171,N_11948);
or U13251 (N_13251,N_11741,N_12223);
nor U13252 (N_13252,N_10971,N_11870);
xnor U13253 (N_13253,N_10299,N_11989);
nand U13254 (N_13254,N_12146,N_12016);
and U13255 (N_13255,N_10515,N_10751);
nand U13256 (N_13256,N_11406,N_10006);
or U13257 (N_13257,N_11579,N_11288);
nor U13258 (N_13258,N_11484,N_11006);
or U13259 (N_13259,N_11601,N_11295);
or U13260 (N_13260,N_10576,N_10421);
nor U13261 (N_13261,N_10508,N_11111);
nand U13262 (N_13262,N_11405,N_12407);
xor U13263 (N_13263,N_10376,N_10598);
or U13264 (N_13264,N_10247,N_12419);
and U13265 (N_13265,N_12142,N_10132);
nor U13266 (N_13266,N_11999,N_11927);
and U13267 (N_13267,N_11296,N_11914);
or U13268 (N_13268,N_12315,N_11595);
or U13269 (N_13269,N_10050,N_10830);
or U13270 (N_13270,N_10213,N_11634);
xor U13271 (N_13271,N_12086,N_11972);
xor U13272 (N_13272,N_12080,N_12457);
xor U13273 (N_13273,N_10234,N_10964);
xor U13274 (N_13274,N_12482,N_10045);
nor U13275 (N_13275,N_11536,N_10980);
or U13276 (N_13276,N_12132,N_10144);
xnor U13277 (N_13277,N_11284,N_11893);
nor U13278 (N_13278,N_12155,N_10320);
nand U13279 (N_13279,N_11664,N_12327);
xnor U13280 (N_13280,N_11798,N_10060);
xor U13281 (N_13281,N_10969,N_11144);
and U13282 (N_13282,N_11780,N_11710);
and U13283 (N_13283,N_11188,N_11124);
nor U13284 (N_13284,N_10803,N_10452);
xor U13285 (N_13285,N_11326,N_11074);
nor U13286 (N_13286,N_10959,N_11629);
xnor U13287 (N_13287,N_12416,N_11333);
nand U13288 (N_13288,N_11429,N_10464);
nor U13289 (N_13289,N_10008,N_11064);
nor U13290 (N_13290,N_10261,N_10571);
xnor U13291 (N_13291,N_10300,N_12156);
or U13292 (N_13292,N_10610,N_10067);
nand U13293 (N_13293,N_10835,N_10259);
nor U13294 (N_13294,N_11042,N_11842);
nand U13295 (N_13295,N_10507,N_10138);
nor U13296 (N_13296,N_11607,N_10922);
and U13297 (N_13297,N_10163,N_11250);
xor U13298 (N_13298,N_10371,N_11130);
and U13299 (N_13299,N_10086,N_10664);
nand U13300 (N_13300,N_10537,N_10939);
and U13301 (N_13301,N_10609,N_12181);
and U13302 (N_13302,N_12494,N_12092);
nand U13303 (N_13303,N_12075,N_10916);
nand U13304 (N_13304,N_12228,N_11395);
and U13305 (N_13305,N_11584,N_10931);
nor U13306 (N_13306,N_10255,N_10313);
xnor U13307 (N_13307,N_11926,N_12176);
nor U13308 (N_13308,N_11354,N_11379);
xnor U13309 (N_13309,N_10406,N_12020);
xnor U13310 (N_13310,N_12459,N_11882);
nor U13311 (N_13311,N_10617,N_11025);
nor U13312 (N_13312,N_11644,N_12242);
xor U13313 (N_13313,N_11894,N_11194);
nor U13314 (N_13314,N_11636,N_11617);
or U13315 (N_13315,N_11715,N_11202);
or U13316 (N_13316,N_11088,N_11615);
xnor U13317 (N_13317,N_11988,N_11765);
or U13318 (N_13318,N_10618,N_12477);
xnor U13319 (N_13319,N_11105,N_11529);
and U13320 (N_13320,N_11642,N_12167);
or U13321 (N_13321,N_11289,N_11782);
xor U13322 (N_13322,N_11614,N_12304);
or U13323 (N_13323,N_10318,N_11129);
nor U13324 (N_13324,N_10297,N_11497);
and U13325 (N_13325,N_12387,N_11560);
xnor U13326 (N_13326,N_11015,N_10566);
xor U13327 (N_13327,N_10802,N_11261);
nor U13328 (N_13328,N_11566,N_11728);
or U13329 (N_13329,N_11056,N_11723);
nand U13330 (N_13330,N_11240,N_11490);
nand U13331 (N_13331,N_12398,N_10396);
xor U13332 (N_13332,N_12464,N_11193);
or U13333 (N_13333,N_10624,N_11272);
nor U13334 (N_13334,N_12364,N_11513);
nor U13335 (N_13335,N_10122,N_11140);
nor U13336 (N_13336,N_12087,N_12450);
or U13337 (N_13337,N_12410,N_10176);
and U13338 (N_13338,N_11050,N_11880);
nand U13339 (N_13339,N_12386,N_11792);
and U13340 (N_13340,N_11438,N_10119);
nand U13341 (N_13341,N_12040,N_10486);
nand U13342 (N_13342,N_10479,N_10260);
nand U13343 (N_13343,N_12226,N_10212);
nand U13344 (N_13344,N_12372,N_11858);
or U13345 (N_13345,N_10342,N_10742);
xor U13346 (N_13346,N_11248,N_12465);
and U13347 (N_13347,N_11738,N_12456);
and U13348 (N_13348,N_11226,N_12342);
or U13349 (N_13349,N_12325,N_10717);
nor U13350 (N_13350,N_10341,N_11844);
xnor U13351 (N_13351,N_11285,N_12438);
nor U13352 (N_13352,N_11184,N_10233);
nand U13353 (N_13353,N_12281,N_11480);
nand U13354 (N_13354,N_11699,N_11422);
nor U13355 (N_13355,N_10752,N_12319);
xor U13356 (N_13356,N_12221,N_11981);
nand U13357 (N_13357,N_10151,N_10807);
xnor U13358 (N_13358,N_12236,N_12264);
and U13359 (N_13359,N_11756,N_10720);
xnor U13360 (N_13360,N_10804,N_10068);
xnor U13361 (N_13361,N_10476,N_10611);
or U13362 (N_13362,N_10578,N_12063);
nor U13363 (N_13363,N_10239,N_10979);
and U13364 (N_13364,N_11624,N_11022);
nor U13365 (N_13365,N_11148,N_11311);
nor U13366 (N_13366,N_10921,N_11081);
xnor U13367 (N_13367,N_10690,N_10593);
nor U13368 (N_13368,N_11282,N_11957);
nand U13369 (N_13369,N_11329,N_11853);
xnor U13370 (N_13370,N_11909,N_11058);
nor U13371 (N_13371,N_10786,N_11860);
nand U13372 (N_13372,N_10996,N_12060);
or U13373 (N_13373,N_11492,N_10741);
or U13374 (N_13374,N_10645,N_12294);
or U13375 (N_13375,N_11180,N_11581);
nand U13376 (N_13376,N_11390,N_11667);
or U13377 (N_13377,N_11841,N_11167);
and U13378 (N_13378,N_12047,N_10547);
nand U13379 (N_13379,N_10713,N_11959);
nand U13380 (N_13380,N_12338,N_12141);
or U13381 (N_13381,N_10650,N_12492);
nor U13382 (N_13382,N_10179,N_11770);
nand U13383 (N_13383,N_10886,N_10197);
nand U13384 (N_13384,N_10403,N_11631);
nor U13385 (N_13385,N_12225,N_11303);
and U13386 (N_13386,N_11952,N_10907);
xor U13387 (N_13387,N_11945,N_11374);
and U13388 (N_13388,N_12293,N_12430);
xor U13389 (N_13389,N_11301,N_11700);
xor U13390 (N_13390,N_10731,N_12052);
nor U13391 (N_13391,N_11924,N_11023);
or U13392 (N_13392,N_10970,N_11812);
nand U13393 (N_13393,N_10674,N_12094);
and U13394 (N_13394,N_12088,N_11138);
nor U13395 (N_13395,N_11593,N_10654);
and U13396 (N_13396,N_10352,N_11511);
and U13397 (N_13397,N_11992,N_10330);
or U13398 (N_13398,N_10011,N_12260);
and U13399 (N_13399,N_10164,N_11991);
xor U13400 (N_13400,N_11011,N_10195);
and U13401 (N_13401,N_11172,N_10496);
nor U13402 (N_13402,N_10545,N_10734);
nor U13403 (N_13403,N_12474,N_10057);
nor U13404 (N_13404,N_10296,N_12033);
and U13405 (N_13405,N_10853,N_12486);
nand U13406 (N_13406,N_11065,N_11096);
or U13407 (N_13407,N_12106,N_10258);
and U13408 (N_13408,N_10231,N_10377);
nor U13409 (N_13409,N_12034,N_11101);
nor U13410 (N_13410,N_10900,N_11247);
nor U13411 (N_13411,N_10810,N_11946);
xor U13412 (N_13412,N_11461,N_12024);
nand U13413 (N_13413,N_10947,N_10074);
nor U13414 (N_13414,N_12050,N_10211);
nor U13415 (N_13415,N_11708,N_10329);
and U13416 (N_13416,N_11887,N_11152);
and U13417 (N_13417,N_11431,N_12115);
xnor U13418 (N_13418,N_12131,N_11599);
or U13419 (N_13419,N_10754,N_11694);
nand U13420 (N_13420,N_12313,N_10451);
nor U13421 (N_13421,N_11702,N_10880);
or U13422 (N_13422,N_10116,N_12219);
nand U13423 (N_13423,N_11766,N_11157);
or U13424 (N_13424,N_11116,N_10651);
and U13425 (N_13425,N_11353,N_11550);
and U13426 (N_13426,N_12272,N_11775);
or U13427 (N_13427,N_10620,N_10359);
xnor U13428 (N_13428,N_12350,N_12147);
xnor U13429 (N_13429,N_11290,N_11572);
and U13430 (N_13430,N_12005,N_10194);
xnor U13431 (N_13431,N_10662,N_11939);
xnor U13432 (N_13432,N_10001,N_11383);
or U13433 (N_13433,N_11205,N_10331);
nand U13434 (N_13434,N_11663,N_11150);
nand U13435 (N_13435,N_11479,N_11281);
nor U13436 (N_13436,N_10002,N_10414);
xor U13437 (N_13437,N_11243,N_11486);
nor U13438 (N_13438,N_11799,N_11786);
nor U13439 (N_13439,N_11472,N_10945);
or U13440 (N_13440,N_11051,N_11218);
or U13441 (N_13441,N_12475,N_10657);
and U13442 (N_13442,N_10058,N_11123);
nor U13443 (N_13443,N_11843,N_10367);
or U13444 (N_13444,N_12072,N_10162);
xor U13445 (N_13445,N_10881,N_12057);
or U13446 (N_13446,N_10118,N_10860);
nor U13447 (N_13447,N_10801,N_10776);
or U13448 (N_13448,N_11228,N_11641);
nor U13449 (N_13449,N_12148,N_11847);
nand U13450 (N_13450,N_12123,N_11559);
nor U13451 (N_13451,N_10823,N_11206);
xnor U13452 (N_13452,N_11608,N_12120);
or U13453 (N_13453,N_11373,N_10337);
or U13454 (N_13454,N_11275,N_11964);
and U13455 (N_13455,N_12151,N_11291);
nor U13456 (N_13456,N_11598,N_10438);
nand U13457 (N_13457,N_12344,N_11286);
xor U13458 (N_13458,N_10224,N_10405);
xor U13459 (N_13459,N_11241,N_10271);
and U13460 (N_13460,N_11055,N_12453);
or U13461 (N_13461,N_10555,N_10998);
nand U13462 (N_13462,N_10217,N_11651);
nand U13463 (N_13463,N_12413,N_12369);
or U13464 (N_13464,N_10628,N_10340);
nand U13465 (N_13465,N_10351,N_11562);
and U13466 (N_13466,N_10943,N_12276);
nand U13467 (N_13467,N_11618,N_11018);
xnor U13468 (N_13468,N_11120,N_11093);
and U13469 (N_13469,N_11997,N_10425);
and U13470 (N_13470,N_10056,N_10838);
nand U13471 (N_13471,N_10018,N_10166);
and U13472 (N_13472,N_10356,N_11037);
nor U13473 (N_13473,N_10462,N_10029);
or U13474 (N_13474,N_10535,N_10936);
nand U13475 (N_13475,N_10042,N_11010);
nor U13476 (N_13476,N_10082,N_10099);
xor U13477 (N_13477,N_12445,N_10243);
or U13478 (N_13478,N_11947,N_12076);
nand U13479 (N_13479,N_11596,N_11351);
and U13480 (N_13480,N_11888,N_10911);
nand U13481 (N_13481,N_11332,N_10466);
nand U13482 (N_13482,N_11868,N_11403);
nand U13483 (N_13483,N_11958,N_11122);
xor U13484 (N_13484,N_10993,N_11293);
and U13485 (N_13485,N_10540,N_11771);
nand U13486 (N_13486,N_11784,N_10811);
and U13487 (N_13487,N_11635,N_12425);
nand U13488 (N_13488,N_11758,N_10499);
or U13489 (N_13489,N_10102,N_10839);
nand U13490 (N_13490,N_10791,N_11279);
nor U13491 (N_13491,N_11378,N_11435);
nand U13492 (N_13492,N_10244,N_10048);
nand U13493 (N_13493,N_11524,N_10192);
nor U13494 (N_13494,N_10120,N_12135);
or U13495 (N_13495,N_10196,N_12003);
nor U13496 (N_13496,N_10130,N_11426);
or U13497 (N_13497,N_10766,N_10139);
nor U13498 (N_13498,N_11590,N_12485);
and U13499 (N_13499,N_11730,N_11577);
nor U13500 (N_13500,N_10347,N_11160);
or U13501 (N_13501,N_11223,N_10266);
xnor U13502 (N_13502,N_12411,N_11199);
nand U13503 (N_13503,N_10778,N_11514);
and U13504 (N_13504,N_10953,N_10037);
xnor U13505 (N_13505,N_11357,N_11554);
or U13506 (N_13506,N_11352,N_11024);
xor U13507 (N_13507,N_11752,N_10165);
xnor U13508 (N_13508,N_10143,N_12101);
or U13509 (N_13509,N_10923,N_11075);
or U13510 (N_13510,N_11721,N_10622);
nand U13511 (N_13511,N_11108,N_12248);
or U13512 (N_13512,N_11407,N_11491);
and U13513 (N_13513,N_11555,N_10714);
or U13514 (N_13514,N_12214,N_11849);
xor U13515 (N_13515,N_12440,N_10409);
and U13516 (N_13516,N_11331,N_10686);
xor U13517 (N_13517,N_10787,N_11867);
and U13518 (N_13518,N_11268,N_11961);
or U13519 (N_13519,N_10899,N_10488);
and U13520 (N_13520,N_10277,N_10808);
nor U13521 (N_13521,N_11489,N_11881);
xor U13522 (N_13522,N_10482,N_10307);
nor U13523 (N_13523,N_10917,N_12203);
and U13524 (N_13524,N_11500,N_11612);
or U13525 (N_13525,N_12162,N_12240);
nand U13526 (N_13526,N_10206,N_12083);
nor U13527 (N_13527,N_10862,N_12002);
xor U13528 (N_13528,N_12400,N_11856);
and U13529 (N_13529,N_12139,N_11666);
and U13530 (N_13530,N_11104,N_10453);
xor U13531 (N_13531,N_11605,N_12125);
and U13532 (N_13532,N_12388,N_11943);
nor U13533 (N_13533,N_10222,N_10424);
nand U13534 (N_13534,N_11425,N_10859);
xnor U13535 (N_13535,N_11052,N_12169);
nor U13536 (N_13536,N_10052,N_10719);
nand U13537 (N_13537,N_11170,N_12134);
nor U13538 (N_13538,N_10745,N_10896);
xor U13539 (N_13539,N_10559,N_10704);
or U13540 (N_13540,N_11062,N_10412);
nor U13541 (N_13541,N_11968,N_10319);
nor U13542 (N_13542,N_10590,N_11714);
nand U13543 (N_13543,N_12361,N_11772);
or U13544 (N_13544,N_11539,N_10301);
xor U13545 (N_13545,N_10386,N_10463);
nor U13546 (N_13546,N_11719,N_10431);
nor U13547 (N_13547,N_11984,N_11327);
xor U13548 (N_13548,N_12393,N_10078);
nand U13549 (N_13549,N_11419,N_10675);
xnor U13550 (N_13550,N_11259,N_10908);
nand U13551 (N_13551,N_12222,N_10152);
or U13552 (N_13552,N_10158,N_10716);
xor U13553 (N_13553,N_11341,N_10310);
nor U13554 (N_13554,N_10573,N_11337);
or U13555 (N_13555,N_11454,N_11079);
nand U13556 (N_13556,N_10782,N_12079);
or U13557 (N_13557,N_11610,N_11092);
nand U13558 (N_13558,N_10273,N_11597);
xnor U13559 (N_13559,N_11531,N_12469);
nand U13560 (N_13560,N_12362,N_11722);
and U13561 (N_13561,N_10012,N_10668);
nand U13562 (N_13562,N_10877,N_11321);
or U13563 (N_13563,N_11283,N_10311);
nor U13564 (N_13564,N_12200,N_12349);
xor U13565 (N_13565,N_12476,N_11825);
nor U13566 (N_13566,N_11040,N_11091);
nand U13567 (N_13567,N_10701,N_10902);
nand U13568 (N_13568,N_11400,N_10314);
and U13569 (N_13569,N_11085,N_11546);
nor U13570 (N_13570,N_11908,N_10030);
nand U13571 (N_13571,N_10526,N_10141);
nand U13572 (N_13572,N_11220,N_11646);
xnor U13573 (N_13573,N_12368,N_10344);
or U13574 (N_13574,N_10175,N_12117);
nor U13575 (N_13575,N_11776,N_11671);
or U13576 (N_13576,N_10106,N_12091);
nor U13577 (N_13577,N_10912,N_11970);
or U13578 (N_13578,N_12439,N_12480);
nand U13579 (N_13579,N_10101,N_11688);
or U13580 (N_13580,N_11589,N_11408);
nand U13581 (N_13581,N_10511,N_10226);
nand U13582 (N_13582,N_10248,N_10630);
and U13583 (N_13583,N_10852,N_11736);
or U13584 (N_13584,N_11869,N_11146);
nand U13585 (N_13585,N_12081,N_12343);
nor U13586 (N_13586,N_10470,N_11315);
and U13587 (N_13587,N_10385,N_12353);
or U13588 (N_13588,N_11192,N_11297);
nand U13589 (N_13589,N_10005,N_12090);
nand U13590 (N_13590,N_12035,N_10442);
and U13591 (N_13591,N_10108,N_12496);
and U13592 (N_13592,N_10369,N_11100);
xnor U13593 (N_13593,N_10484,N_10346);
and U13594 (N_13594,N_10528,N_10957);
nand U13595 (N_13595,N_10295,N_12397);
or U13596 (N_13596,N_11266,N_11442);
or U13597 (N_13597,N_10085,N_10531);
or U13598 (N_13598,N_12038,N_12019);
nor U13599 (N_13599,N_10131,N_11675);
nand U13600 (N_13600,N_11563,N_11382);
or U13601 (N_13601,N_12277,N_10203);
nand U13602 (N_13602,N_11336,N_10267);
or U13603 (N_13603,N_11620,N_11060);
and U13604 (N_13604,N_11159,N_10848);
xnor U13605 (N_13605,N_10428,N_12335);
xnor U13606 (N_13606,N_11090,N_11445);
nand U13607 (N_13607,N_11119,N_11673);
or U13608 (N_13608,N_10173,N_11904);
xor U13609 (N_13609,N_11421,N_11214);
or U13610 (N_13610,N_11444,N_12208);
and U13611 (N_13611,N_11257,N_10379);
xnor U13612 (N_13612,N_11417,N_12463);
nor U13613 (N_13613,N_10187,N_10380);
or U13614 (N_13614,N_11017,N_11649);
or U13615 (N_13615,N_10666,N_11133);
xnor U13616 (N_13616,N_10069,N_10370);
or U13617 (N_13617,N_12093,N_11740);
or U13618 (N_13618,N_11347,N_10035);
and U13619 (N_13619,N_11907,N_11033);
or U13620 (N_13620,N_10768,N_10746);
and U13621 (N_13621,N_10795,N_12271);
xnor U13622 (N_13622,N_12028,N_10123);
nor U13623 (N_13623,N_11883,N_12112);
and U13624 (N_13624,N_10387,N_10580);
and U13625 (N_13625,N_12036,N_11690);
nand U13626 (N_13626,N_10516,N_11182);
nand U13627 (N_13627,N_10736,N_10990);
and U13628 (N_13628,N_11483,N_10022);
and U13629 (N_13629,N_11530,N_12061);
and U13630 (N_13630,N_12145,N_10373);
or U13631 (N_13631,N_12403,N_10105);
and U13632 (N_13632,N_10871,N_11504);
nor U13633 (N_13633,N_10501,N_10075);
and U13634 (N_13634,N_10028,N_11757);
nor U13635 (N_13635,N_11761,N_11103);
nor U13636 (N_13636,N_10793,N_10960);
nor U13637 (N_13637,N_11851,N_11181);
and U13638 (N_13638,N_11439,N_10730);
and U13639 (N_13639,N_11396,N_12234);
nand U13640 (N_13640,N_10536,N_10601);
xor U13641 (N_13641,N_10298,N_12233);
or U13642 (N_13642,N_11346,N_11837);
xnor U13643 (N_13643,N_12472,N_11207);
nand U13644 (N_13644,N_10702,N_10137);
xnor U13645 (N_13645,N_11545,N_10004);
or U13646 (N_13646,N_10709,N_11455);
and U13647 (N_13647,N_12251,N_11071);
xnor U13648 (N_13648,N_10073,N_10779);
or U13649 (N_13649,N_10928,N_11838);
and U13650 (N_13650,N_10111,N_12110);
and U13651 (N_13651,N_10054,N_11339);
or U13652 (N_13652,N_10286,N_12478);
and U13653 (N_13653,N_10407,N_11793);
nand U13654 (N_13654,N_10670,N_10397);
and U13655 (N_13655,N_11632,N_12031);
or U13656 (N_13656,N_12263,N_11067);
nor U13657 (N_13657,N_12232,N_10186);
nor U13658 (N_13658,N_11726,N_11232);
xor U13659 (N_13659,N_11824,N_12266);
or U13660 (N_13660,N_10548,N_11204);
xnor U13661 (N_13661,N_10430,N_12165);
nand U13662 (N_13662,N_11735,N_11753);
nand U13663 (N_13663,N_11070,N_11750);
nand U13664 (N_13664,N_10687,N_11077);
and U13665 (N_13665,N_11464,N_11131);
and U13666 (N_13666,N_10833,N_11606);
nand U13667 (N_13667,N_12211,N_11720);
nand U13668 (N_13668,N_10098,N_10728);
xor U13669 (N_13669,N_12099,N_10777);
and U13670 (N_13670,N_12205,N_11061);
nor U13671 (N_13671,N_11502,N_11744);
xnor U13672 (N_13672,N_11068,N_10608);
or U13673 (N_13673,N_10251,N_12462);
and U13674 (N_13674,N_12332,N_11049);
nand U13675 (N_13675,N_11391,N_11304);
nand U13676 (N_13676,N_11245,N_11368);
or U13677 (N_13677,N_10538,N_11689);
and U13678 (N_13678,N_10167,N_11447);
xor U13679 (N_13679,N_10114,N_10236);
and U13680 (N_13680,N_11583,N_12423);
and U13681 (N_13681,N_12274,N_10232);
or U13682 (N_13682,N_10049,N_11966);
nor U13683 (N_13683,N_10156,N_12255);
or U13684 (N_13684,N_11652,N_10509);
and U13685 (N_13685,N_11734,N_11102);
xor U13686 (N_13686,N_11810,N_11809);
and U13687 (N_13687,N_11277,N_10007);
or U13688 (N_13688,N_11834,N_10676);
or U13689 (N_13689,N_10639,N_10312);
nor U13690 (N_13690,N_11054,N_10089);
and U13691 (N_13691,N_10334,N_10354);
xor U13692 (N_13692,N_10722,N_11007);
nor U13693 (N_13693,N_12235,N_10737);
or U13694 (N_13694,N_12105,N_10207);
and U13695 (N_13695,N_10532,N_11393);
or U13696 (N_13696,N_12253,N_11515);
nor U13697 (N_13697,N_10229,N_10978);
nand U13698 (N_13698,N_10245,N_11568);
nand U13699 (N_13699,N_10727,N_11681);
nand U13700 (N_13700,N_10047,N_11087);
and U13701 (N_13701,N_12435,N_12007);
or U13702 (N_13702,N_10184,N_11645);
or U13703 (N_13703,N_12412,N_10885);
or U13704 (N_13704,N_12212,N_11637);
and U13705 (N_13705,N_11235,N_10685);
xor U13706 (N_13706,N_12046,N_12121);
nor U13707 (N_13707,N_10133,N_11410);
and U13708 (N_13708,N_10032,N_10364);
nor U13709 (N_13709,N_11020,N_11274);
xor U13710 (N_13710,N_12068,N_11126);
and U13711 (N_13711,N_10758,N_12116);
or U13712 (N_13712,N_11755,N_10539);
nor U13713 (N_13713,N_11986,N_11219);
and U13714 (N_13714,N_10942,N_12269);
xor U13715 (N_13715,N_12252,N_10750);
nand U13716 (N_13716,N_12262,N_10422);
nor U13717 (N_13717,N_11940,N_11928);
and U13718 (N_13718,N_11083,N_11955);
or U13719 (N_13719,N_10326,N_11818);
or U13720 (N_13720,N_11534,N_11889);
nand U13721 (N_13721,N_12424,N_12053);
nor U13722 (N_13722,N_12409,N_11628);
and U13723 (N_13723,N_12443,N_10644);
xnor U13724 (N_13724,N_10863,N_10914);
and U13725 (N_13725,N_12054,N_10189);
nor U13726 (N_13726,N_12451,N_11936);
and U13727 (N_13727,N_10553,N_11467);
nand U13728 (N_13728,N_10739,N_12444);
nand U13729 (N_13729,N_10652,N_11683);
nand U13730 (N_13730,N_10512,N_12461);
or U13731 (N_13731,N_12247,N_10506);
and U13732 (N_13732,N_11322,N_11549);
xnor U13733 (N_13733,N_11305,N_10575);
nand U13734 (N_13734,N_10794,N_10419);
nand U13735 (N_13735,N_11879,N_10829);
nor U13736 (N_13736,N_11687,N_11165);
and U13737 (N_13737,N_10855,N_11983);
and U13738 (N_13738,N_12197,N_10872);
nand U13739 (N_13739,N_10417,N_11655);
nand U13740 (N_13740,N_10070,N_11325);
nor U13741 (N_13741,N_11507,N_11234);
or U13742 (N_13742,N_11538,N_10281);
nor U13743 (N_13743,N_10263,N_10066);
or U13744 (N_13744,N_10792,N_10694);
and U13745 (N_13745,N_12484,N_12188);
nand U13746 (N_13746,N_12097,N_11684);
nor U13747 (N_13747,N_11813,N_10504);
nand U13748 (N_13748,N_12059,N_11803);
and U13749 (N_13749,N_10395,N_12292);
xnor U13750 (N_13750,N_10098,N_11427);
or U13751 (N_13751,N_10391,N_10212);
and U13752 (N_13752,N_11746,N_10776);
nor U13753 (N_13753,N_11480,N_11248);
nand U13754 (N_13754,N_11119,N_10836);
and U13755 (N_13755,N_11490,N_12411);
and U13756 (N_13756,N_11779,N_10299);
xor U13757 (N_13757,N_12313,N_11212);
nand U13758 (N_13758,N_10594,N_10904);
nor U13759 (N_13759,N_10305,N_11343);
nand U13760 (N_13760,N_12358,N_11765);
nor U13761 (N_13761,N_10326,N_10096);
xor U13762 (N_13762,N_11001,N_12341);
nor U13763 (N_13763,N_11657,N_11392);
nor U13764 (N_13764,N_10036,N_10304);
nor U13765 (N_13765,N_11068,N_10898);
xor U13766 (N_13766,N_10176,N_10262);
xor U13767 (N_13767,N_12353,N_11394);
nand U13768 (N_13768,N_11930,N_11628);
and U13769 (N_13769,N_10778,N_11894);
nor U13770 (N_13770,N_11516,N_11390);
xor U13771 (N_13771,N_11496,N_11614);
nor U13772 (N_13772,N_11837,N_12320);
or U13773 (N_13773,N_11154,N_12317);
or U13774 (N_13774,N_11363,N_11946);
nand U13775 (N_13775,N_11243,N_11415);
or U13776 (N_13776,N_11172,N_10656);
nand U13777 (N_13777,N_10172,N_10945);
nor U13778 (N_13778,N_10390,N_11334);
nor U13779 (N_13779,N_11180,N_12030);
xnor U13780 (N_13780,N_11500,N_11534);
nand U13781 (N_13781,N_11088,N_10236);
xnor U13782 (N_13782,N_10477,N_11119);
xor U13783 (N_13783,N_12267,N_12270);
xnor U13784 (N_13784,N_11683,N_11334);
or U13785 (N_13785,N_10696,N_11793);
nand U13786 (N_13786,N_10017,N_11247);
nand U13787 (N_13787,N_12111,N_10051);
or U13788 (N_13788,N_12257,N_10045);
nand U13789 (N_13789,N_11741,N_12016);
or U13790 (N_13790,N_11417,N_12066);
xor U13791 (N_13791,N_11128,N_11411);
nor U13792 (N_13792,N_11549,N_10347);
xnor U13793 (N_13793,N_11304,N_10636);
nand U13794 (N_13794,N_10910,N_11595);
nand U13795 (N_13795,N_10431,N_10173);
and U13796 (N_13796,N_10011,N_12425);
nand U13797 (N_13797,N_10389,N_10549);
xnor U13798 (N_13798,N_10719,N_11764);
nor U13799 (N_13799,N_11570,N_12110);
nand U13800 (N_13800,N_10915,N_12257);
and U13801 (N_13801,N_12361,N_10151);
and U13802 (N_13802,N_12367,N_11387);
or U13803 (N_13803,N_10678,N_10596);
nand U13804 (N_13804,N_11917,N_10763);
nor U13805 (N_13805,N_10175,N_11674);
nand U13806 (N_13806,N_11069,N_10396);
or U13807 (N_13807,N_10149,N_10410);
nand U13808 (N_13808,N_11430,N_11375);
or U13809 (N_13809,N_10656,N_11870);
nand U13810 (N_13810,N_11736,N_11053);
nor U13811 (N_13811,N_12337,N_10745);
nor U13812 (N_13812,N_11722,N_11376);
and U13813 (N_13813,N_10273,N_10286);
nor U13814 (N_13814,N_10560,N_11775);
nor U13815 (N_13815,N_12049,N_11093);
and U13816 (N_13816,N_12294,N_10502);
and U13817 (N_13817,N_12471,N_11369);
nand U13818 (N_13818,N_11709,N_11471);
or U13819 (N_13819,N_10257,N_10143);
xnor U13820 (N_13820,N_11108,N_10662);
and U13821 (N_13821,N_11957,N_12014);
and U13822 (N_13822,N_12371,N_11985);
or U13823 (N_13823,N_10346,N_12044);
nor U13824 (N_13824,N_12164,N_12077);
nor U13825 (N_13825,N_11399,N_10355);
and U13826 (N_13826,N_11729,N_10975);
xor U13827 (N_13827,N_11099,N_11293);
or U13828 (N_13828,N_11746,N_10358);
xor U13829 (N_13829,N_10809,N_10576);
nor U13830 (N_13830,N_12424,N_11207);
and U13831 (N_13831,N_10996,N_12294);
xor U13832 (N_13832,N_10851,N_11385);
nand U13833 (N_13833,N_11226,N_12343);
nor U13834 (N_13834,N_12258,N_12416);
nor U13835 (N_13835,N_12235,N_10399);
or U13836 (N_13836,N_11234,N_10554);
nand U13837 (N_13837,N_10420,N_11550);
and U13838 (N_13838,N_12441,N_10893);
nand U13839 (N_13839,N_11956,N_12298);
or U13840 (N_13840,N_11299,N_11693);
nor U13841 (N_13841,N_10483,N_12136);
nor U13842 (N_13842,N_10984,N_12229);
and U13843 (N_13843,N_11837,N_12208);
xnor U13844 (N_13844,N_10646,N_11952);
or U13845 (N_13845,N_11308,N_11903);
or U13846 (N_13846,N_12222,N_11720);
xor U13847 (N_13847,N_10386,N_11544);
nor U13848 (N_13848,N_11509,N_11278);
xnor U13849 (N_13849,N_11869,N_11153);
or U13850 (N_13850,N_10639,N_12255);
or U13851 (N_13851,N_12110,N_11382);
and U13852 (N_13852,N_11157,N_11459);
nor U13853 (N_13853,N_10907,N_11823);
nand U13854 (N_13854,N_11469,N_12326);
xor U13855 (N_13855,N_10681,N_10737);
xnor U13856 (N_13856,N_12302,N_10934);
and U13857 (N_13857,N_11179,N_10130);
or U13858 (N_13858,N_11587,N_10041);
or U13859 (N_13859,N_11330,N_12225);
nor U13860 (N_13860,N_10243,N_10529);
or U13861 (N_13861,N_11100,N_11553);
xor U13862 (N_13862,N_12339,N_10621);
or U13863 (N_13863,N_11741,N_10135);
and U13864 (N_13864,N_10647,N_12005);
or U13865 (N_13865,N_10763,N_12076);
xnor U13866 (N_13866,N_12470,N_11919);
and U13867 (N_13867,N_12045,N_12172);
nand U13868 (N_13868,N_11966,N_11386);
nor U13869 (N_13869,N_10899,N_11084);
nor U13870 (N_13870,N_10760,N_12138);
nand U13871 (N_13871,N_12442,N_10518);
nand U13872 (N_13872,N_12466,N_10906);
and U13873 (N_13873,N_11318,N_11052);
or U13874 (N_13874,N_10685,N_11401);
and U13875 (N_13875,N_12374,N_11140);
and U13876 (N_13876,N_10527,N_10807);
and U13877 (N_13877,N_11620,N_10325);
or U13878 (N_13878,N_11758,N_11349);
nand U13879 (N_13879,N_11651,N_11905);
nand U13880 (N_13880,N_10037,N_10024);
xnor U13881 (N_13881,N_10621,N_10915);
and U13882 (N_13882,N_10673,N_12217);
nand U13883 (N_13883,N_10606,N_10035);
and U13884 (N_13884,N_12280,N_10018);
and U13885 (N_13885,N_10019,N_10388);
or U13886 (N_13886,N_11514,N_11372);
xor U13887 (N_13887,N_10361,N_10247);
and U13888 (N_13888,N_10129,N_10250);
nand U13889 (N_13889,N_10167,N_10286);
or U13890 (N_13890,N_12337,N_10019);
or U13891 (N_13891,N_10175,N_10195);
nand U13892 (N_13892,N_12316,N_11085);
and U13893 (N_13893,N_11570,N_11951);
nor U13894 (N_13894,N_11000,N_11572);
or U13895 (N_13895,N_12033,N_12143);
nand U13896 (N_13896,N_11648,N_12293);
or U13897 (N_13897,N_10339,N_10010);
and U13898 (N_13898,N_11827,N_10162);
nand U13899 (N_13899,N_11492,N_12453);
nor U13900 (N_13900,N_10672,N_11476);
nor U13901 (N_13901,N_11038,N_10227);
or U13902 (N_13902,N_11021,N_11148);
nand U13903 (N_13903,N_10158,N_11632);
nand U13904 (N_13904,N_12338,N_10516);
and U13905 (N_13905,N_10205,N_10806);
nor U13906 (N_13906,N_11032,N_11738);
and U13907 (N_13907,N_10236,N_11002);
nor U13908 (N_13908,N_12142,N_11611);
nor U13909 (N_13909,N_11418,N_11535);
xor U13910 (N_13910,N_10887,N_10987);
nor U13911 (N_13911,N_11762,N_11022);
xor U13912 (N_13912,N_11325,N_10433);
or U13913 (N_13913,N_12327,N_11482);
nor U13914 (N_13914,N_11012,N_11570);
nand U13915 (N_13915,N_11690,N_10529);
xnor U13916 (N_13916,N_10159,N_10563);
nand U13917 (N_13917,N_10506,N_11349);
nor U13918 (N_13918,N_10829,N_12286);
or U13919 (N_13919,N_10139,N_12142);
nand U13920 (N_13920,N_10786,N_12159);
or U13921 (N_13921,N_10456,N_12229);
nor U13922 (N_13922,N_12450,N_10631);
nor U13923 (N_13923,N_12464,N_10006);
nand U13924 (N_13924,N_11060,N_11485);
nand U13925 (N_13925,N_10594,N_10031);
xnor U13926 (N_13926,N_11799,N_10124);
xnor U13927 (N_13927,N_10524,N_11282);
nand U13928 (N_13928,N_12116,N_11996);
or U13929 (N_13929,N_11228,N_10888);
nor U13930 (N_13930,N_10514,N_10571);
xor U13931 (N_13931,N_11601,N_11982);
xor U13932 (N_13932,N_10175,N_11237);
nor U13933 (N_13933,N_11184,N_11147);
nor U13934 (N_13934,N_12005,N_10320);
and U13935 (N_13935,N_10158,N_12020);
nand U13936 (N_13936,N_11454,N_10332);
xor U13937 (N_13937,N_11631,N_10145);
xnor U13938 (N_13938,N_10175,N_10328);
nand U13939 (N_13939,N_11235,N_10381);
xor U13940 (N_13940,N_12280,N_11950);
and U13941 (N_13941,N_10470,N_11301);
nor U13942 (N_13942,N_11414,N_11693);
and U13943 (N_13943,N_10070,N_11410);
or U13944 (N_13944,N_10189,N_11326);
or U13945 (N_13945,N_11156,N_10378);
xnor U13946 (N_13946,N_12419,N_11692);
or U13947 (N_13947,N_10243,N_10451);
nand U13948 (N_13948,N_10479,N_10462);
and U13949 (N_13949,N_11907,N_10172);
or U13950 (N_13950,N_11541,N_11701);
or U13951 (N_13951,N_11703,N_11472);
and U13952 (N_13952,N_11679,N_10431);
nand U13953 (N_13953,N_10242,N_11708);
and U13954 (N_13954,N_10637,N_10284);
nand U13955 (N_13955,N_10703,N_10745);
and U13956 (N_13956,N_10672,N_10155);
nor U13957 (N_13957,N_10721,N_12387);
or U13958 (N_13958,N_11158,N_12036);
nor U13959 (N_13959,N_12353,N_12443);
xor U13960 (N_13960,N_10957,N_10070);
xor U13961 (N_13961,N_10289,N_10615);
and U13962 (N_13962,N_11419,N_10232);
or U13963 (N_13963,N_11392,N_12140);
or U13964 (N_13964,N_11535,N_11649);
xor U13965 (N_13965,N_11022,N_10212);
xor U13966 (N_13966,N_10001,N_10963);
nand U13967 (N_13967,N_11890,N_11208);
nand U13968 (N_13968,N_11422,N_12294);
xor U13969 (N_13969,N_12452,N_10377);
xnor U13970 (N_13970,N_12302,N_10508);
and U13971 (N_13971,N_11473,N_12366);
and U13972 (N_13972,N_11370,N_10695);
or U13973 (N_13973,N_11394,N_11164);
and U13974 (N_13974,N_12010,N_12407);
nand U13975 (N_13975,N_11245,N_10781);
nor U13976 (N_13976,N_11094,N_11351);
xor U13977 (N_13977,N_11324,N_11555);
nor U13978 (N_13978,N_11807,N_10878);
nand U13979 (N_13979,N_12195,N_11876);
or U13980 (N_13980,N_10646,N_10353);
or U13981 (N_13981,N_11906,N_11057);
and U13982 (N_13982,N_11618,N_10270);
or U13983 (N_13983,N_11010,N_10386);
xor U13984 (N_13984,N_12202,N_10807);
nor U13985 (N_13985,N_10743,N_10734);
xnor U13986 (N_13986,N_10030,N_11541);
and U13987 (N_13987,N_10697,N_10524);
nand U13988 (N_13988,N_10109,N_11009);
or U13989 (N_13989,N_11554,N_12139);
or U13990 (N_13990,N_10969,N_11595);
and U13991 (N_13991,N_12294,N_10102);
nor U13992 (N_13992,N_11655,N_11950);
or U13993 (N_13993,N_10197,N_10290);
nand U13994 (N_13994,N_10206,N_11492);
or U13995 (N_13995,N_10760,N_11872);
nor U13996 (N_13996,N_10278,N_10660);
nand U13997 (N_13997,N_11249,N_11969);
and U13998 (N_13998,N_10398,N_11494);
and U13999 (N_13999,N_10750,N_12283);
nand U14000 (N_14000,N_10517,N_11042);
nand U14001 (N_14001,N_10523,N_11145);
and U14002 (N_14002,N_11105,N_11324);
and U14003 (N_14003,N_10095,N_11279);
nor U14004 (N_14004,N_10651,N_11393);
nor U14005 (N_14005,N_10877,N_12066);
xnor U14006 (N_14006,N_11029,N_10452);
and U14007 (N_14007,N_10242,N_12282);
nor U14008 (N_14008,N_10482,N_10122);
nand U14009 (N_14009,N_11006,N_12135);
or U14010 (N_14010,N_11549,N_10364);
xnor U14011 (N_14011,N_11962,N_11968);
xnor U14012 (N_14012,N_10032,N_11406);
nand U14013 (N_14013,N_10813,N_10253);
nand U14014 (N_14014,N_11623,N_10206);
xor U14015 (N_14015,N_12142,N_10697);
xor U14016 (N_14016,N_12044,N_10973);
and U14017 (N_14017,N_10600,N_11812);
nand U14018 (N_14018,N_10583,N_10389);
and U14019 (N_14019,N_11072,N_11745);
nand U14020 (N_14020,N_12178,N_11313);
nand U14021 (N_14021,N_10690,N_10940);
nand U14022 (N_14022,N_10056,N_12247);
xor U14023 (N_14023,N_12417,N_11790);
or U14024 (N_14024,N_10807,N_10981);
nor U14025 (N_14025,N_11158,N_10761);
xor U14026 (N_14026,N_11644,N_11059);
or U14027 (N_14027,N_10142,N_11239);
nand U14028 (N_14028,N_10696,N_12250);
nand U14029 (N_14029,N_11300,N_11823);
and U14030 (N_14030,N_11122,N_11421);
xor U14031 (N_14031,N_11876,N_11783);
nand U14032 (N_14032,N_11831,N_12046);
nand U14033 (N_14033,N_12077,N_11268);
or U14034 (N_14034,N_11764,N_10396);
or U14035 (N_14035,N_10149,N_12426);
nor U14036 (N_14036,N_11702,N_10594);
or U14037 (N_14037,N_11402,N_11305);
nand U14038 (N_14038,N_12497,N_10067);
or U14039 (N_14039,N_11523,N_12007);
and U14040 (N_14040,N_10565,N_12463);
nor U14041 (N_14041,N_12080,N_10758);
nand U14042 (N_14042,N_10132,N_10786);
or U14043 (N_14043,N_12227,N_12376);
nor U14044 (N_14044,N_11717,N_10545);
and U14045 (N_14045,N_10482,N_11410);
xnor U14046 (N_14046,N_12421,N_11853);
and U14047 (N_14047,N_11789,N_12292);
nand U14048 (N_14048,N_12083,N_11091);
nor U14049 (N_14049,N_12196,N_11957);
nand U14050 (N_14050,N_10521,N_10276);
nand U14051 (N_14051,N_10953,N_10416);
nand U14052 (N_14052,N_11430,N_11445);
and U14053 (N_14053,N_11399,N_10359);
or U14054 (N_14054,N_12266,N_10012);
or U14055 (N_14055,N_10415,N_10520);
xor U14056 (N_14056,N_11684,N_12292);
nor U14057 (N_14057,N_11671,N_11441);
xnor U14058 (N_14058,N_10356,N_11942);
nand U14059 (N_14059,N_11530,N_11072);
nor U14060 (N_14060,N_10195,N_10881);
or U14061 (N_14061,N_12271,N_12248);
or U14062 (N_14062,N_10912,N_12485);
nor U14063 (N_14063,N_11973,N_10120);
or U14064 (N_14064,N_11818,N_11555);
and U14065 (N_14065,N_11168,N_11242);
and U14066 (N_14066,N_11592,N_11467);
nor U14067 (N_14067,N_10668,N_11171);
nor U14068 (N_14068,N_10454,N_10410);
or U14069 (N_14069,N_10985,N_11455);
nand U14070 (N_14070,N_10500,N_11294);
xnor U14071 (N_14071,N_12446,N_11194);
xor U14072 (N_14072,N_11986,N_11233);
nor U14073 (N_14073,N_12302,N_11819);
and U14074 (N_14074,N_11245,N_11328);
or U14075 (N_14075,N_10544,N_11513);
nor U14076 (N_14076,N_10950,N_10271);
or U14077 (N_14077,N_10809,N_10525);
or U14078 (N_14078,N_10804,N_10229);
and U14079 (N_14079,N_11692,N_11195);
xor U14080 (N_14080,N_10729,N_11626);
and U14081 (N_14081,N_12416,N_12166);
nand U14082 (N_14082,N_12448,N_10721);
xor U14083 (N_14083,N_12038,N_10873);
or U14084 (N_14084,N_10279,N_10104);
nor U14085 (N_14085,N_12380,N_12270);
or U14086 (N_14086,N_11235,N_12219);
nand U14087 (N_14087,N_11007,N_12323);
xnor U14088 (N_14088,N_10472,N_10957);
and U14089 (N_14089,N_10442,N_11861);
nand U14090 (N_14090,N_12484,N_10593);
nand U14091 (N_14091,N_10877,N_12492);
nor U14092 (N_14092,N_10067,N_10640);
xor U14093 (N_14093,N_10123,N_11640);
nand U14094 (N_14094,N_11046,N_11221);
nand U14095 (N_14095,N_11386,N_11336);
nand U14096 (N_14096,N_11160,N_11887);
xnor U14097 (N_14097,N_10964,N_10142);
xnor U14098 (N_14098,N_10957,N_10965);
or U14099 (N_14099,N_11417,N_11846);
nor U14100 (N_14100,N_11187,N_10756);
nand U14101 (N_14101,N_12486,N_11250);
and U14102 (N_14102,N_11565,N_10285);
nand U14103 (N_14103,N_11744,N_10667);
xor U14104 (N_14104,N_10653,N_12207);
nand U14105 (N_14105,N_11431,N_11114);
nand U14106 (N_14106,N_10080,N_10613);
nand U14107 (N_14107,N_12031,N_11971);
nand U14108 (N_14108,N_11332,N_11833);
xnor U14109 (N_14109,N_10800,N_11165);
and U14110 (N_14110,N_10794,N_10548);
or U14111 (N_14111,N_11154,N_11462);
or U14112 (N_14112,N_12474,N_10680);
nor U14113 (N_14113,N_10797,N_10679);
xor U14114 (N_14114,N_11136,N_11254);
nand U14115 (N_14115,N_10741,N_12488);
nor U14116 (N_14116,N_11883,N_12030);
xor U14117 (N_14117,N_11469,N_10587);
nand U14118 (N_14118,N_10666,N_10911);
nor U14119 (N_14119,N_10244,N_11357);
nand U14120 (N_14120,N_11305,N_10467);
or U14121 (N_14121,N_10877,N_12093);
nand U14122 (N_14122,N_10794,N_11106);
nand U14123 (N_14123,N_11436,N_12122);
or U14124 (N_14124,N_10131,N_12448);
or U14125 (N_14125,N_11226,N_11515);
and U14126 (N_14126,N_11630,N_11302);
nor U14127 (N_14127,N_11724,N_12404);
or U14128 (N_14128,N_10488,N_11543);
nor U14129 (N_14129,N_10348,N_12087);
or U14130 (N_14130,N_12255,N_10562);
or U14131 (N_14131,N_12468,N_11553);
and U14132 (N_14132,N_11082,N_10960);
or U14133 (N_14133,N_10563,N_12433);
and U14134 (N_14134,N_10284,N_10368);
xnor U14135 (N_14135,N_10975,N_12066);
or U14136 (N_14136,N_11412,N_11588);
nor U14137 (N_14137,N_11401,N_11576);
xor U14138 (N_14138,N_10423,N_11118);
and U14139 (N_14139,N_11052,N_12079);
xor U14140 (N_14140,N_11006,N_10163);
and U14141 (N_14141,N_11001,N_11242);
or U14142 (N_14142,N_11543,N_11359);
or U14143 (N_14143,N_12038,N_12209);
xnor U14144 (N_14144,N_11362,N_12294);
xor U14145 (N_14145,N_11042,N_12071);
xnor U14146 (N_14146,N_12419,N_11843);
xnor U14147 (N_14147,N_10913,N_12079);
and U14148 (N_14148,N_10421,N_10879);
and U14149 (N_14149,N_10371,N_10765);
nor U14150 (N_14150,N_11380,N_12286);
or U14151 (N_14151,N_11707,N_12115);
and U14152 (N_14152,N_11299,N_10254);
or U14153 (N_14153,N_10483,N_12294);
xor U14154 (N_14154,N_10515,N_11123);
or U14155 (N_14155,N_11105,N_11276);
and U14156 (N_14156,N_11984,N_10389);
and U14157 (N_14157,N_12286,N_11548);
and U14158 (N_14158,N_11089,N_10383);
xnor U14159 (N_14159,N_11646,N_10684);
xnor U14160 (N_14160,N_11418,N_12389);
nor U14161 (N_14161,N_11066,N_11601);
or U14162 (N_14162,N_10805,N_12444);
and U14163 (N_14163,N_11594,N_10846);
nand U14164 (N_14164,N_12374,N_10735);
or U14165 (N_14165,N_10665,N_11299);
and U14166 (N_14166,N_10721,N_12183);
nor U14167 (N_14167,N_12247,N_11927);
and U14168 (N_14168,N_11982,N_10802);
and U14169 (N_14169,N_10695,N_11496);
and U14170 (N_14170,N_10611,N_10673);
or U14171 (N_14171,N_12356,N_11672);
and U14172 (N_14172,N_10557,N_12057);
and U14173 (N_14173,N_12334,N_10323);
xor U14174 (N_14174,N_11189,N_11025);
or U14175 (N_14175,N_10719,N_11808);
xnor U14176 (N_14176,N_11424,N_10941);
nand U14177 (N_14177,N_11000,N_11860);
nor U14178 (N_14178,N_12355,N_11668);
nand U14179 (N_14179,N_12246,N_12274);
or U14180 (N_14180,N_10952,N_12282);
nand U14181 (N_14181,N_10239,N_10625);
nor U14182 (N_14182,N_12455,N_10079);
xnor U14183 (N_14183,N_11669,N_11934);
nand U14184 (N_14184,N_12049,N_11136);
or U14185 (N_14185,N_10132,N_10609);
or U14186 (N_14186,N_10220,N_11433);
xnor U14187 (N_14187,N_10760,N_11862);
nor U14188 (N_14188,N_10316,N_11832);
nand U14189 (N_14189,N_12244,N_12468);
nand U14190 (N_14190,N_11960,N_11398);
xor U14191 (N_14191,N_11596,N_10889);
and U14192 (N_14192,N_11991,N_11969);
and U14193 (N_14193,N_10661,N_11712);
or U14194 (N_14194,N_10770,N_11972);
xor U14195 (N_14195,N_10216,N_10964);
xor U14196 (N_14196,N_10061,N_11714);
xnor U14197 (N_14197,N_12100,N_10819);
or U14198 (N_14198,N_10188,N_12156);
nor U14199 (N_14199,N_11213,N_12423);
and U14200 (N_14200,N_10763,N_10240);
nor U14201 (N_14201,N_10280,N_11225);
nand U14202 (N_14202,N_11729,N_11475);
xor U14203 (N_14203,N_11781,N_10139);
xor U14204 (N_14204,N_11640,N_10818);
xor U14205 (N_14205,N_12103,N_10426);
nand U14206 (N_14206,N_10554,N_10017);
nor U14207 (N_14207,N_10850,N_10790);
and U14208 (N_14208,N_10771,N_12420);
nand U14209 (N_14209,N_10333,N_10564);
xnor U14210 (N_14210,N_10074,N_12369);
nor U14211 (N_14211,N_10614,N_10713);
and U14212 (N_14212,N_12035,N_10663);
and U14213 (N_14213,N_11769,N_10454);
or U14214 (N_14214,N_11827,N_11218);
nand U14215 (N_14215,N_11465,N_10565);
nand U14216 (N_14216,N_10912,N_11916);
and U14217 (N_14217,N_12190,N_10364);
xor U14218 (N_14218,N_11740,N_12084);
xor U14219 (N_14219,N_11728,N_11803);
nand U14220 (N_14220,N_12239,N_12373);
or U14221 (N_14221,N_11099,N_10036);
or U14222 (N_14222,N_11002,N_11950);
nand U14223 (N_14223,N_11320,N_10658);
and U14224 (N_14224,N_10578,N_12031);
and U14225 (N_14225,N_10046,N_11974);
or U14226 (N_14226,N_10880,N_10953);
and U14227 (N_14227,N_11320,N_11238);
and U14228 (N_14228,N_12307,N_10367);
nand U14229 (N_14229,N_10446,N_10657);
and U14230 (N_14230,N_11754,N_11238);
or U14231 (N_14231,N_10501,N_12215);
nand U14232 (N_14232,N_12045,N_11777);
nor U14233 (N_14233,N_11041,N_10325);
or U14234 (N_14234,N_10663,N_11169);
and U14235 (N_14235,N_10101,N_10436);
or U14236 (N_14236,N_11426,N_12416);
or U14237 (N_14237,N_11819,N_10867);
nor U14238 (N_14238,N_11682,N_10435);
nand U14239 (N_14239,N_11306,N_11477);
or U14240 (N_14240,N_10127,N_11885);
and U14241 (N_14241,N_12357,N_11448);
and U14242 (N_14242,N_11506,N_10230);
and U14243 (N_14243,N_11875,N_11263);
and U14244 (N_14244,N_10088,N_12246);
or U14245 (N_14245,N_12228,N_10796);
nor U14246 (N_14246,N_11700,N_11343);
nor U14247 (N_14247,N_10780,N_11384);
xor U14248 (N_14248,N_10969,N_12253);
xnor U14249 (N_14249,N_12075,N_10700);
and U14250 (N_14250,N_11241,N_12251);
nand U14251 (N_14251,N_10144,N_11085);
or U14252 (N_14252,N_10845,N_11930);
and U14253 (N_14253,N_12469,N_12098);
or U14254 (N_14254,N_11687,N_10335);
nor U14255 (N_14255,N_10225,N_11298);
nand U14256 (N_14256,N_12197,N_10815);
nor U14257 (N_14257,N_11141,N_11830);
nand U14258 (N_14258,N_10876,N_11085);
xnor U14259 (N_14259,N_11618,N_11771);
nor U14260 (N_14260,N_10166,N_10603);
nor U14261 (N_14261,N_11576,N_11986);
xor U14262 (N_14262,N_10830,N_11961);
xnor U14263 (N_14263,N_12328,N_11368);
nand U14264 (N_14264,N_11044,N_10666);
or U14265 (N_14265,N_11554,N_11760);
nand U14266 (N_14266,N_11148,N_12384);
nor U14267 (N_14267,N_12073,N_10015);
and U14268 (N_14268,N_11738,N_10346);
and U14269 (N_14269,N_10259,N_10885);
xnor U14270 (N_14270,N_12248,N_11894);
nand U14271 (N_14271,N_11666,N_11670);
nand U14272 (N_14272,N_10552,N_11451);
and U14273 (N_14273,N_11074,N_10023);
nand U14274 (N_14274,N_10795,N_11641);
nor U14275 (N_14275,N_11019,N_11573);
xor U14276 (N_14276,N_10088,N_12126);
nand U14277 (N_14277,N_12260,N_11717);
nor U14278 (N_14278,N_12139,N_12341);
and U14279 (N_14279,N_11155,N_10890);
nor U14280 (N_14280,N_11477,N_11236);
nor U14281 (N_14281,N_10681,N_11090);
or U14282 (N_14282,N_11042,N_10202);
and U14283 (N_14283,N_10820,N_11884);
nand U14284 (N_14284,N_10795,N_11389);
xor U14285 (N_14285,N_11836,N_10670);
nor U14286 (N_14286,N_11075,N_12126);
or U14287 (N_14287,N_12250,N_12363);
or U14288 (N_14288,N_10726,N_10460);
or U14289 (N_14289,N_11100,N_11683);
xor U14290 (N_14290,N_11152,N_11481);
xor U14291 (N_14291,N_11425,N_10354);
or U14292 (N_14292,N_10283,N_11374);
nand U14293 (N_14293,N_11194,N_11224);
and U14294 (N_14294,N_11723,N_10914);
nor U14295 (N_14295,N_10805,N_12481);
xor U14296 (N_14296,N_10420,N_12476);
or U14297 (N_14297,N_10315,N_10482);
or U14298 (N_14298,N_10970,N_10165);
nand U14299 (N_14299,N_11192,N_10944);
or U14300 (N_14300,N_12485,N_11243);
and U14301 (N_14301,N_12343,N_10423);
or U14302 (N_14302,N_10248,N_12366);
nor U14303 (N_14303,N_10242,N_10144);
nand U14304 (N_14304,N_11940,N_10661);
and U14305 (N_14305,N_11118,N_10191);
and U14306 (N_14306,N_12238,N_11006);
or U14307 (N_14307,N_11335,N_12088);
or U14308 (N_14308,N_11376,N_11998);
or U14309 (N_14309,N_12212,N_11415);
nor U14310 (N_14310,N_11454,N_10196);
or U14311 (N_14311,N_12324,N_11845);
xor U14312 (N_14312,N_12401,N_12441);
or U14313 (N_14313,N_10786,N_11191);
nand U14314 (N_14314,N_11391,N_11990);
or U14315 (N_14315,N_10108,N_10773);
nand U14316 (N_14316,N_12021,N_12175);
or U14317 (N_14317,N_11406,N_10896);
or U14318 (N_14318,N_10304,N_11217);
nand U14319 (N_14319,N_10461,N_11660);
or U14320 (N_14320,N_11345,N_10885);
xor U14321 (N_14321,N_12344,N_11683);
nor U14322 (N_14322,N_11364,N_11544);
or U14323 (N_14323,N_10877,N_11264);
nand U14324 (N_14324,N_10981,N_12110);
nand U14325 (N_14325,N_10459,N_10339);
nor U14326 (N_14326,N_12484,N_10609);
nand U14327 (N_14327,N_11265,N_10710);
or U14328 (N_14328,N_11445,N_11225);
and U14329 (N_14329,N_10622,N_11457);
nand U14330 (N_14330,N_10193,N_11260);
nand U14331 (N_14331,N_11972,N_10916);
xnor U14332 (N_14332,N_12073,N_11033);
nand U14333 (N_14333,N_12055,N_11783);
and U14334 (N_14334,N_10003,N_11289);
nand U14335 (N_14335,N_12264,N_10317);
xnor U14336 (N_14336,N_11153,N_10563);
or U14337 (N_14337,N_10136,N_10161);
and U14338 (N_14338,N_11492,N_11699);
nand U14339 (N_14339,N_10814,N_11656);
nand U14340 (N_14340,N_11803,N_10661);
nor U14341 (N_14341,N_10528,N_10416);
nand U14342 (N_14342,N_12145,N_11745);
xor U14343 (N_14343,N_11125,N_12184);
nand U14344 (N_14344,N_10732,N_10625);
or U14345 (N_14345,N_12464,N_11344);
and U14346 (N_14346,N_10828,N_12392);
or U14347 (N_14347,N_10305,N_10174);
nor U14348 (N_14348,N_11264,N_11345);
nor U14349 (N_14349,N_11314,N_10757);
nor U14350 (N_14350,N_12036,N_11314);
nand U14351 (N_14351,N_10591,N_10336);
xnor U14352 (N_14352,N_10587,N_11232);
nand U14353 (N_14353,N_10071,N_10283);
nand U14354 (N_14354,N_10236,N_12275);
xnor U14355 (N_14355,N_12324,N_11783);
xnor U14356 (N_14356,N_10201,N_11591);
nor U14357 (N_14357,N_10208,N_11090);
nor U14358 (N_14358,N_10756,N_12075);
nand U14359 (N_14359,N_12297,N_10331);
or U14360 (N_14360,N_11201,N_10772);
xor U14361 (N_14361,N_10886,N_10349);
nor U14362 (N_14362,N_11155,N_10708);
or U14363 (N_14363,N_10776,N_10706);
nor U14364 (N_14364,N_10869,N_12093);
nand U14365 (N_14365,N_12119,N_11899);
and U14366 (N_14366,N_10480,N_12186);
nand U14367 (N_14367,N_12485,N_12087);
xnor U14368 (N_14368,N_12036,N_11900);
xnor U14369 (N_14369,N_12257,N_11117);
and U14370 (N_14370,N_11798,N_10132);
and U14371 (N_14371,N_11900,N_10984);
nor U14372 (N_14372,N_10253,N_11580);
nor U14373 (N_14373,N_10012,N_10227);
or U14374 (N_14374,N_10077,N_10045);
nor U14375 (N_14375,N_11815,N_12438);
xor U14376 (N_14376,N_11180,N_11115);
or U14377 (N_14377,N_11426,N_11397);
nand U14378 (N_14378,N_12494,N_10570);
or U14379 (N_14379,N_11385,N_10704);
or U14380 (N_14380,N_10956,N_12065);
nand U14381 (N_14381,N_11791,N_12064);
xor U14382 (N_14382,N_10054,N_11325);
or U14383 (N_14383,N_12284,N_11531);
nand U14384 (N_14384,N_10111,N_10036);
xnor U14385 (N_14385,N_10896,N_10250);
nand U14386 (N_14386,N_10207,N_10792);
nand U14387 (N_14387,N_11680,N_10387);
xnor U14388 (N_14388,N_11080,N_11624);
xor U14389 (N_14389,N_11983,N_10514);
nor U14390 (N_14390,N_11859,N_10489);
and U14391 (N_14391,N_11238,N_10212);
nor U14392 (N_14392,N_10947,N_10696);
or U14393 (N_14393,N_11563,N_12163);
nor U14394 (N_14394,N_11412,N_10795);
or U14395 (N_14395,N_10634,N_11519);
nand U14396 (N_14396,N_11780,N_10929);
and U14397 (N_14397,N_11136,N_10823);
or U14398 (N_14398,N_11377,N_11452);
or U14399 (N_14399,N_12064,N_12139);
nand U14400 (N_14400,N_10839,N_10373);
nand U14401 (N_14401,N_11253,N_12177);
and U14402 (N_14402,N_12150,N_11959);
nand U14403 (N_14403,N_10905,N_10390);
xor U14404 (N_14404,N_11155,N_10849);
or U14405 (N_14405,N_10960,N_12166);
nand U14406 (N_14406,N_12482,N_11376);
and U14407 (N_14407,N_11700,N_10136);
and U14408 (N_14408,N_10898,N_11152);
nand U14409 (N_14409,N_12454,N_10149);
and U14410 (N_14410,N_10813,N_11173);
nand U14411 (N_14411,N_11818,N_10143);
nor U14412 (N_14412,N_11860,N_12102);
nor U14413 (N_14413,N_10013,N_10734);
xor U14414 (N_14414,N_10805,N_11751);
or U14415 (N_14415,N_11707,N_11810);
xor U14416 (N_14416,N_11546,N_10242);
nand U14417 (N_14417,N_10625,N_10362);
nor U14418 (N_14418,N_10902,N_10183);
xnor U14419 (N_14419,N_12081,N_10228);
or U14420 (N_14420,N_11148,N_10654);
and U14421 (N_14421,N_10556,N_11562);
and U14422 (N_14422,N_10437,N_11876);
and U14423 (N_14423,N_11580,N_11979);
nor U14424 (N_14424,N_12084,N_12018);
and U14425 (N_14425,N_10641,N_11173);
nor U14426 (N_14426,N_10538,N_12208);
nor U14427 (N_14427,N_11288,N_10360);
nor U14428 (N_14428,N_11643,N_11273);
nor U14429 (N_14429,N_10150,N_11211);
xnor U14430 (N_14430,N_11602,N_11630);
xor U14431 (N_14431,N_11405,N_12288);
nor U14432 (N_14432,N_10914,N_12289);
or U14433 (N_14433,N_11023,N_11390);
xnor U14434 (N_14434,N_11916,N_11702);
or U14435 (N_14435,N_10209,N_11793);
xnor U14436 (N_14436,N_10564,N_11314);
nor U14437 (N_14437,N_10672,N_10070);
nand U14438 (N_14438,N_11859,N_12090);
nor U14439 (N_14439,N_12463,N_11341);
nand U14440 (N_14440,N_10529,N_10041);
nor U14441 (N_14441,N_12446,N_10937);
nand U14442 (N_14442,N_10761,N_10487);
nand U14443 (N_14443,N_11147,N_10557);
nor U14444 (N_14444,N_11450,N_11733);
and U14445 (N_14445,N_10271,N_10601);
nor U14446 (N_14446,N_10574,N_10758);
nor U14447 (N_14447,N_11451,N_11040);
xnor U14448 (N_14448,N_11647,N_10207);
or U14449 (N_14449,N_11402,N_12422);
nor U14450 (N_14450,N_11174,N_11798);
nand U14451 (N_14451,N_10636,N_12375);
nor U14452 (N_14452,N_10201,N_11787);
and U14453 (N_14453,N_11254,N_10610);
and U14454 (N_14454,N_11439,N_11835);
or U14455 (N_14455,N_11293,N_11211);
nor U14456 (N_14456,N_10556,N_11839);
xor U14457 (N_14457,N_10392,N_11528);
and U14458 (N_14458,N_11382,N_11014);
xor U14459 (N_14459,N_11560,N_11049);
or U14460 (N_14460,N_11247,N_10380);
nor U14461 (N_14461,N_12100,N_10687);
and U14462 (N_14462,N_11948,N_11038);
nor U14463 (N_14463,N_10967,N_10723);
or U14464 (N_14464,N_11555,N_11581);
nor U14465 (N_14465,N_10815,N_11780);
and U14466 (N_14466,N_10622,N_10258);
and U14467 (N_14467,N_12253,N_10250);
nor U14468 (N_14468,N_11243,N_12433);
nand U14469 (N_14469,N_12049,N_10241);
nand U14470 (N_14470,N_11595,N_11519);
or U14471 (N_14471,N_12249,N_10892);
and U14472 (N_14472,N_10002,N_10282);
nor U14473 (N_14473,N_10831,N_11734);
and U14474 (N_14474,N_10423,N_10262);
or U14475 (N_14475,N_10077,N_11026);
nor U14476 (N_14476,N_10748,N_12009);
nor U14477 (N_14477,N_11707,N_10393);
and U14478 (N_14478,N_11657,N_10487);
and U14479 (N_14479,N_12442,N_11090);
xor U14480 (N_14480,N_11671,N_10865);
or U14481 (N_14481,N_10245,N_10923);
or U14482 (N_14482,N_11999,N_10862);
nor U14483 (N_14483,N_10509,N_12163);
xnor U14484 (N_14484,N_11573,N_12179);
xor U14485 (N_14485,N_10234,N_11557);
and U14486 (N_14486,N_12444,N_12438);
and U14487 (N_14487,N_10695,N_11841);
and U14488 (N_14488,N_10452,N_10313);
nor U14489 (N_14489,N_10665,N_10222);
xnor U14490 (N_14490,N_11773,N_10257);
nand U14491 (N_14491,N_11856,N_10790);
nand U14492 (N_14492,N_10580,N_11338);
nor U14493 (N_14493,N_12217,N_12020);
nand U14494 (N_14494,N_11548,N_11126);
nand U14495 (N_14495,N_11314,N_11319);
nor U14496 (N_14496,N_10811,N_11614);
nor U14497 (N_14497,N_10421,N_10785);
xor U14498 (N_14498,N_11918,N_10791);
xor U14499 (N_14499,N_11547,N_11004);
or U14500 (N_14500,N_12228,N_11786);
nor U14501 (N_14501,N_10444,N_10012);
nor U14502 (N_14502,N_10530,N_11675);
xor U14503 (N_14503,N_11252,N_11542);
nor U14504 (N_14504,N_11328,N_10455);
and U14505 (N_14505,N_11775,N_12073);
or U14506 (N_14506,N_10707,N_10873);
or U14507 (N_14507,N_12222,N_10875);
or U14508 (N_14508,N_10260,N_10615);
xnor U14509 (N_14509,N_11045,N_10679);
or U14510 (N_14510,N_10623,N_10927);
nor U14511 (N_14511,N_10064,N_10151);
and U14512 (N_14512,N_10026,N_11654);
and U14513 (N_14513,N_11745,N_11442);
and U14514 (N_14514,N_11221,N_10499);
xnor U14515 (N_14515,N_12020,N_10348);
or U14516 (N_14516,N_11860,N_12108);
or U14517 (N_14517,N_11118,N_10698);
nor U14518 (N_14518,N_12161,N_11709);
and U14519 (N_14519,N_12396,N_11615);
and U14520 (N_14520,N_11581,N_12313);
nor U14521 (N_14521,N_12166,N_10180);
nand U14522 (N_14522,N_11574,N_12311);
nor U14523 (N_14523,N_10060,N_11925);
or U14524 (N_14524,N_10227,N_10341);
nand U14525 (N_14525,N_12458,N_11816);
xor U14526 (N_14526,N_10780,N_12369);
xnor U14527 (N_14527,N_11878,N_12330);
nand U14528 (N_14528,N_11342,N_12274);
and U14529 (N_14529,N_11838,N_11737);
and U14530 (N_14530,N_10766,N_11362);
xnor U14531 (N_14531,N_11623,N_12328);
xnor U14532 (N_14532,N_11829,N_11963);
nor U14533 (N_14533,N_11958,N_12025);
nand U14534 (N_14534,N_11984,N_10136);
nor U14535 (N_14535,N_10481,N_11220);
xnor U14536 (N_14536,N_10594,N_11812);
nand U14537 (N_14537,N_10815,N_10044);
xor U14538 (N_14538,N_12126,N_12353);
xnor U14539 (N_14539,N_12384,N_11019);
nand U14540 (N_14540,N_10422,N_10244);
nor U14541 (N_14541,N_11260,N_12083);
nand U14542 (N_14542,N_12397,N_10584);
xnor U14543 (N_14543,N_10941,N_10951);
and U14544 (N_14544,N_10340,N_11649);
nor U14545 (N_14545,N_10454,N_11234);
nor U14546 (N_14546,N_12207,N_11480);
and U14547 (N_14547,N_10842,N_10009);
nor U14548 (N_14548,N_10303,N_10467);
or U14549 (N_14549,N_12018,N_10145);
xor U14550 (N_14550,N_11882,N_11410);
nand U14551 (N_14551,N_12301,N_11938);
nand U14552 (N_14552,N_10563,N_11935);
nand U14553 (N_14553,N_10946,N_10322);
xor U14554 (N_14554,N_12226,N_12461);
nand U14555 (N_14555,N_11182,N_11934);
nor U14556 (N_14556,N_11246,N_12261);
nand U14557 (N_14557,N_11259,N_11245);
xnor U14558 (N_14558,N_11514,N_10664);
nand U14559 (N_14559,N_10454,N_11481);
or U14560 (N_14560,N_12039,N_12005);
or U14561 (N_14561,N_11784,N_11837);
or U14562 (N_14562,N_12093,N_11531);
or U14563 (N_14563,N_11209,N_10051);
and U14564 (N_14564,N_10911,N_10345);
xnor U14565 (N_14565,N_11204,N_10764);
nor U14566 (N_14566,N_10538,N_11005);
nor U14567 (N_14567,N_11411,N_11315);
and U14568 (N_14568,N_10492,N_11629);
or U14569 (N_14569,N_10867,N_12112);
or U14570 (N_14570,N_11503,N_12214);
or U14571 (N_14571,N_10148,N_10464);
xor U14572 (N_14572,N_11415,N_12069);
xor U14573 (N_14573,N_10719,N_10294);
nor U14574 (N_14574,N_11778,N_11000);
nor U14575 (N_14575,N_11411,N_11684);
or U14576 (N_14576,N_11836,N_12287);
or U14577 (N_14577,N_10392,N_10883);
nand U14578 (N_14578,N_10584,N_12056);
nor U14579 (N_14579,N_10775,N_11395);
and U14580 (N_14580,N_10008,N_11644);
xnor U14581 (N_14581,N_11528,N_10663);
xnor U14582 (N_14582,N_11486,N_11994);
nand U14583 (N_14583,N_11690,N_10618);
xor U14584 (N_14584,N_10875,N_11457);
nand U14585 (N_14585,N_12082,N_11883);
and U14586 (N_14586,N_10454,N_11439);
nand U14587 (N_14587,N_11961,N_11270);
nand U14588 (N_14588,N_10360,N_11474);
nor U14589 (N_14589,N_10793,N_11231);
and U14590 (N_14590,N_11371,N_10568);
nor U14591 (N_14591,N_11247,N_11335);
and U14592 (N_14592,N_11141,N_10775);
and U14593 (N_14593,N_10225,N_10702);
and U14594 (N_14594,N_11707,N_11176);
nand U14595 (N_14595,N_12297,N_11524);
or U14596 (N_14596,N_10441,N_11372);
or U14597 (N_14597,N_11280,N_12359);
or U14598 (N_14598,N_11839,N_10635);
nor U14599 (N_14599,N_10924,N_11799);
and U14600 (N_14600,N_11717,N_10653);
and U14601 (N_14601,N_11594,N_10818);
or U14602 (N_14602,N_10804,N_10049);
nand U14603 (N_14603,N_11304,N_11615);
or U14604 (N_14604,N_12233,N_10114);
and U14605 (N_14605,N_10417,N_10864);
nand U14606 (N_14606,N_12394,N_11808);
and U14607 (N_14607,N_11707,N_12499);
nand U14608 (N_14608,N_10514,N_10000);
and U14609 (N_14609,N_11757,N_11521);
nand U14610 (N_14610,N_10962,N_11606);
nor U14611 (N_14611,N_11953,N_11211);
or U14612 (N_14612,N_12277,N_10827);
nor U14613 (N_14613,N_10730,N_11723);
or U14614 (N_14614,N_10188,N_10594);
nor U14615 (N_14615,N_12135,N_11666);
and U14616 (N_14616,N_10513,N_11124);
nand U14617 (N_14617,N_11499,N_11240);
and U14618 (N_14618,N_10245,N_10159);
nor U14619 (N_14619,N_10312,N_11849);
xor U14620 (N_14620,N_10694,N_10477);
or U14621 (N_14621,N_11100,N_10451);
xnor U14622 (N_14622,N_12443,N_11032);
or U14623 (N_14623,N_11371,N_10880);
nor U14624 (N_14624,N_11479,N_10861);
xor U14625 (N_14625,N_10153,N_10667);
nor U14626 (N_14626,N_11572,N_10003);
xor U14627 (N_14627,N_10921,N_10235);
nand U14628 (N_14628,N_12296,N_11535);
nand U14629 (N_14629,N_11341,N_10101);
and U14630 (N_14630,N_10543,N_11395);
and U14631 (N_14631,N_10683,N_10005);
or U14632 (N_14632,N_11455,N_11780);
xnor U14633 (N_14633,N_11378,N_10293);
and U14634 (N_14634,N_12383,N_10126);
and U14635 (N_14635,N_12088,N_10371);
nand U14636 (N_14636,N_10003,N_11272);
nor U14637 (N_14637,N_10954,N_11679);
and U14638 (N_14638,N_11511,N_11369);
nor U14639 (N_14639,N_10220,N_12237);
nor U14640 (N_14640,N_10596,N_12370);
xor U14641 (N_14641,N_10234,N_10474);
nor U14642 (N_14642,N_12126,N_10306);
or U14643 (N_14643,N_12193,N_12099);
nor U14644 (N_14644,N_11936,N_12092);
nand U14645 (N_14645,N_10067,N_10413);
nor U14646 (N_14646,N_11624,N_10010);
nand U14647 (N_14647,N_12302,N_11881);
xor U14648 (N_14648,N_11008,N_11014);
nor U14649 (N_14649,N_11186,N_12248);
and U14650 (N_14650,N_10017,N_12455);
nor U14651 (N_14651,N_12467,N_10112);
xor U14652 (N_14652,N_12057,N_12300);
nor U14653 (N_14653,N_10999,N_11761);
nor U14654 (N_14654,N_12346,N_11348);
nor U14655 (N_14655,N_10415,N_11277);
nand U14656 (N_14656,N_11460,N_12224);
nor U14657 (N_14657,N_12452,N_11562);
nor U14658 (N_14658,N_10270,N_11024);
xnor U14659 (N_14659,N_11033,N_11931);
nor U14660 (N_14660,N_12036,N_11042);
nor U14661 (N_14661,N_10214,N_11367);
nand U14662 (N_14662,N_12301,N_12227);
xnor U14663 (N_14663,N_11418,N_10320);
and U14664 (N_14664,N_10536,N_10346);
and U14665 (N_14665,N_11928,N_12287);
and U14666 (N_14666,N_10711,N_11219);
and U14667 (N_14667,N_10163,N_11287);
nand U14668 (N_14668,N_10595,N_12089);
and U14669 (N_14669,N_11152,N_10736);
nor U14670 (N_14670,N_11013,N_10428);
xor U14671 (N_14671,N_10337,N_11040);
nor U14672 (N_14672,N_11163,N_11793);
or U14673 (N_14673,N_10420,N_11209);
nor U14674 (N_14674,N_12092,N_11533);
and U14675 (N_14675,N_12212,N_10355);
nand U14676 (N_14676,N_11921,N_12499);
xnor U14677 (N_14677,N_12176,N_11666);
nand U14678 (N_14678,N_12305,N_11565);
nand U14679 (N_14679,N_11585,N_10889);
or U14680 (N_14680,N_11302,N_11818);
and U14681 (N_14681,N_11706,N_11130);
xnor U14682 (N_14682,N_11821,N_10844);
or U14683 (N_14683,N_12288,N_10928);
xnor U14684 (N_14684,N_11017,N_10077);
nor U14685 (N_14685,N_10339,N_10446);
or U14686 (N_14686,N_10190,N_10173);
nand U14687 (N_14687,N_10402,N_10505);
nand U14688 (N_14688,N_10405,N_10595);
nor U14689 (N_14689,N_12086,N_11608);
and U14690 (N_14690,N_12170,N_10788);
and U14691 (N_14691,N_10033,N_10593);
xnor U14692 (N_14692,N_11535,N_10411);
or U14693 (N_14693,N_11755,N_12163);
and U14694 (N_14694,N_11854,N_12182);
xor U14695 (N_14695,N_10624,N_10598);
xnor U14696 (N_14696,N_10597,N_11652);
xor U14697 (N_14697,N_11566,N_10611);
xor U14698 (N_14698,N_11481,N_11889);
and U14699 (N_14699,N_11364,N_12311);
and U14700 (N_14700,N_12221,N_12115);
nand U14701 (N_14701,N_10001,N_11249);
nand U14702 (N_14702,N_11877,N_11152);
nor U14703 (N_14703,N_10279,N_11972);
or U14704 (N_14704,N_10918,N_10059);
or U14705 (N_14705,N_11054,N_12445);
or U14706 (N_14706,N_12079,N_12444);
and U14707 (N_14707,N_12087,N_12096);
nor U14708 (N_14708,N_11496,N_10654);
nand U14709 (N_14709,N_12397,N_10355);
xor U14710 (N_14710,N_10937,N_10596);
nand U14711 (N_14711,N_10667,N_10211);
and U14712 (N_14712,N_10053,N_10683);
nand U14713 (N_14713,N_10735,N_12325);
and U14714 (N_14714,N_11506,N_10403);
nand U14715 (N_14715,N_10445,N_11446);
nor U14716 (N_14716,N_10624,N_11802);
nand U14717 (N_14717,N_10994,N_11127);
nor U14718 (N_14718,N_10938,N_11060);
and U14719 (N_14719,N_12457,N_12477);
nand U14720 (N_14720,N_11670,N_10909);
nand U14721 (N_14721,N_12484,N_11972);
and U14722 (N_14722,N_10259,N_10509);
nor U14723 (N_14723,N_11139,N_11743);
or U14724 (N_14724,N_11960,N_11525);
nor U14725 (N_14725,N_11590,N_11263);
or U14726 (N_14726,N_10004,N_12321);
xnor U14727 (N_14727,N_11632,N_10195);
nand U14728 (N_14728,N_10377,N_10195);
nor U14729 (N_14729,N_11707,N_10312);
nor U14730 (N_14730,N_11819,N_12483);
nand U14731 (N_14731,N_10795,N_11170);
and U14732 (N_14732,N_11327,N_10847);
xor U14733 (N_14733,N_10573,N_10472);
nand U14734 (N_14734,N_11240,N_10073);
nand U14735 (N_14735,N_11805,N_11652);
nand U14736 (N_14736,N_10606,N_11641);
nand U14737 (N_14737,N_12468,N_11378);
nor U14738 (N_14738,N_10189,N_10215);
or U14739 (N_14739,N_10220,N_11297);
or U14740 (N_14740,N_10024,N_12298);
nor U14741 (N_14741,N_10223,N_10264);
nor U14742 (N_14742,N_11680,N_11221);
nor U14743 (N_14743,N_10562,N_10506);
xor U14744 (N_14744,N_10508,N_11953);
xor U14745 (N_14745,N_11750,N_11825);
nand U14746 (N_14746,N_10652,N_11137);
or U14747 (N_14747,N_11200,N_12189);
nor U14748 (N_14748,N_10925,N_10433);
nand U14749 (N_14749,N_10778,N_10296);
nand U14750 (N_14750,N_11084,N_10709);
and U14751 (N_14751,N_10483,N_10872);
nand U14752 (N_14752,N_11440,N_10798);
and U14753 (N_14753,N_11805,N_11780);
nand U14754 (N_14754,N_12453,N_10275);
and U14755 (N_14755,N_10359,N_12111);
nand U14756 (N_14756,N_11024,N_10168);
nand U14757 (N_14757,N_10109,N_12442);
nand U14758 (N_14758,N_10801,N_10891);
xnor U14759 (N_14759,N_10447,N_12280);
nor U14760 (N_14760,N_10609,N_11984);
and U14761 (N_14761,N_11859,N_10214);
or U14762 (N_14762,N_10635,N_11997);
nor U14763 (N_14763,N_10145,N_11406);
xnor U14764 (N_14764,N_11387,N_10262);
nand U14765 (N_14765,N_10987,N_10542);
and U14766 (N_14766,N_11216,N_11675);
and U14767 (N_14767,N_11815,N_10724);
nand U14768 (N_14768,N_11250,N_11685);
nand U14769 (N_14769,N_10985,N_12245);
xnor U14770 (N_14770,N_10810,N_12393);
or U14771 (N_14771,N_10257,N_10764);
nor U14772 (N_14772,N_12348,N_10155);
or U14773 (N_14773,N_11730,N_12304);
and U14774 (N_14774,N_12126,N_11737);
or U14775 (N_14775,N_10988,N_10329);
and U14776 (N_14776,N_10022,N_12036);
xnor U14777 (N_14777,N_11191,N_10214);
nor U14778 (N_14778,N_10343,N_10058);
and U14779 (N_14779,N_12432,N_10149);
or U14780 (N_14780,N_10640,N_11140);
xor U14781 (N_14781,N_10307,N_11384);
nor U14782 (N_14782,N_11174,N_10312);
nor U14783 (N_14783,N_10044,N_10981);
and U14784 (N_14784,N_11996,N_10933);
and U14785 (N_14785,N_11630,N_10759);
or U14786 (N_14786,N_10533,N_12423);
xnor U14787 (N_14787,N_11482,N_11576);
and U14788 (N_14788,N_11427,N_12243);
xnor U14789 (N_14789,N_10556,N_10320);
nand U14790 (N_14790,N_11712,N_11875);
nor U14791 (N_14791,N_11716,N_12060);
nor U14792 (N_14792,N_11796,N_10720);
xor U14793 (N_14793,N_10371,N_11057);
nand U14794 (N_14794,N_12440,N_11288);
and U14795 (N_14795,N_11490,N_11867);
nand U14796 (N_14796,N_11918,N_10056);
and U14797 (N_14797,N_11745,N_11032);
xnor U14798 (N_14798,N_10400,N_10173);
and U14799 (N_14799,N_11937,N_10195);
nand U14800 (N_14800,N_11406,N_10838);
and U14801 (N_14801,N_11592,N_10883);
xnor U14802 (N_14802,N_11992,N_10871);
nor U14803 (N_14803,N_10157,N_12350);
xor U14804 (N_14804,N_11206,N_10864);
or U14805 (N_14805,N_10537,N_12128);
nand U14806 (N_14806,N_10475,N_11877);
nand U14807 (N_14807,N_10319,N_11389);
or U14808 (N_14808,N_12490,N_12071);
and U14809 (N_14809,N_10586,N_10602);
nand U14810 (N_14810,N_11444,N_11705);
xnor U14811 (N_14811,N_11138,N_10995);
nand U14812 (N_14812,N_12311,N_11868);
nand U14813 (N_14813,N_11210,N_10732);
nor U14814 (N_14814,N_10063,N_12133);
nor U14815 (N_14815,N_10779,N_11335);
or U14816 (N_14816,N_10802,N_11197);
nand U14817 (N_14817,N_11735,N_10988);
and U14818 (N_14818,N_11104,N_10809);
or U14819 (N_14819,N_11071,N_11637);
nand U14820 (N_14820,N_12086,N_11330);
and U14821 (N_14821,N_11656,N_12181);
or U14822 (N_14822,N_10373,N_10722);
nand U14823 (N_14823,N_10404,N_11550);
and U14824 (N_14824,N_11834,N_12454);
or U14825 (N_14825,N_10098,N_12432);
nand U14826 (N_14826,N_11029,N_10943);
and U14827 (N_14827,N_11602,N_11073);
or U14828 (N_14828,N_11839,N_11684);
or U14829 (N_14829,N_12326,N_10984);
xnor U14830 (N_14830,N_11830,N_12249);
nor U14831 (N_14831,N_12327,N_11619);
xnor U14832 (N_14832,N_11318,N_11899);
and U14833 (N_14833,N_12440,N_11595);
nand U14834 (N_14834,N_11028,N_11553);
nor U14835 (N_14835,N_10128,N_10757);
and U14836 (N_14836,N_10784,N_10304);
nand U14837 (N_14837,N_12222,N_10407);
nand U14838 (N_14838,N_12483,N_11970);
nand U14839 (N_14839,N_10902,N_11389);
xor U14840 (N_14840,N_11947,N_11578);
nand U14841 (N_14841,N_11824,N_11314);
nand U14842 (N_14842,N_12414,N_10055);
nor U14843 (N_14843,N_12422,N_11567);
or U14844 (N_14844,N_10470,N_10909);
nand U14845 (N_14845,N_11191,N_12267);
and U14846 (N_14846,N_12115,N_12429);
nor U14847 (N_14847,N_10248,N_12336);
and U14848 (N_14848,N_12339,N_12468);
and U14849 (N_14849,N_11019,N_12284);
and U14850 (N_14850,N_11838,N_11659);
xor U14851 (N_14851,N_12103,N_10774);
xor U14852 (N_14852,N_12186,N_10068);
nand U14853 (N_14853,N_11180,N_10976);
and U14854 (N_14854,N_10659,N_12001);
nor U14855 (N_14855,N_10444,N_10140);
nand U14856 (N_14856,N_10540,N_11828);
xnor U14857 (N_14857,N_12416,N_11949);
nor U14858 (N_14858,N_11035,N_12197);
xor U14859 (N_14859,N_10849,N_11456);
or U14860 (N_14860,N_10962,N_11237);
or U14861 (N_14861,N_10721,N_12489);
and U14862 (N_14862,N_10768,N_11394);
nand U14863 (N_14863,N_11019,N_11807);
xnor U14864 (N_14864,N_10173,N_10363);
and U14865 (N_14865,N_10686,N_11707);
or U14866 (N_14866,N_12207,N_11257);
or U14867 (N_14867,N_12327,N_11800);
and U14868 (N_14868,N_11869,N_11059);
nor U14869 (N_14869,N_10683,N_11626);
xnor U14870 (N_14870,N_10315,N_12347);
nor U14871 (N_14871,N_10737,N_12345);
xor U14872 (N_14872,N_11956,N_11753);
nor U14873 (N_14873,N_10802,N_10686);
nand U14874 (N_14874,N_10282,N_10912);
and U14875 (N_14875,N_12426,N_11765);
or U14876 (N_14876,N_11860,N_10769);
xnor U14877 (N_14877,N_10451,N_10007);
or U14878 (N_14878,N_10262,N_11546);
xor U14879 (N_14879,N_12288,N_11977);
nor U14880 (N_14880,N_12281,N_10029);
xor U14881 (N_14881,N_11842,N_11758);
nand U14882 (N_14882,N_11574,N_12350);
and U14883 (N_14883,N_12227,N_10499);
or U14884 (N_14884,N_10161,N_11462);
xnor U14885 (N_14885,N_10454,N_11715);
xor U14886 (N_14886,N_12226,N_10898);
nor U14887 (N_14887,N_10922,N_10940);
nand U14888 (N_14888,N_10590,N_11409);
or U14889 (N_14889,N_11014,N_11386);
or U14890 (N_14890,N_11354,N_12122);
and U14891 (N_14891,N_11985,N_11425);
nand U14892 (N_14892,N_11010,N_11919);
and U14893 (N_14893,N_10991,N_10861);
nand U14894 (N_14894,N_11804,N_11058);
and U14895 (N_14895,N_10688,N_10039);
nor U14896 (N_14896,N_10556,N_11132);
xor U14897 (N_14897,N_11467,N_11715);
xor U14898 (N_14898,N_11679,N_11570);
and U14899 (N_14899,N_10418,N_11841);
nor U14900 (N_14900,N_10810,N_11569);
xnor U14901 (N_14901,N_12119,N_10567);
xnor U14902 (N_14902,N_10637,N_11811);
nand U14903 (N_14903,N_10663,N_11125);
nand U14904 (N_14904,N_10414,N_11736);
and U14905 (N_14905,N_11850,N_11241);
and U14906 (N_14906,N_11127,N_10172);
nor U14907 (N_14907,N_11836,N_12486);
and U14908 (N_14908,N_10066,N_10001);
and U14909 (N_14909,N_11847,N_10699);
xor U14910 (N_14910,N_10748,N_12269);
nor U14911 (N_14911,N_10842,N_12237);
nor U14912 (N_14912,N_12095,N_10031);
xor U14913 (N_14913,N_10651,N_10706);
or U14914 (N_14914,N_12484,N_10676);
nand U14915 (N_14915,N_11653,N_11060);
and U14916 (N_14916,N_10892,N_10387);
or U14917 (N_14917,N_11232,N_11142);
or U14918 (N_14918,N_12118,N_11141);
and U14919 (N_14919,N_12178,N_11862);
and U14920 (N_14920,N_11930,N_11530);
nor U14921 (N_14921,N_11083,N_11615);
or U14922 (N_14922,N_10853,N_11822);
nor U14923 (N_14923,N_10423,N_11211);
nand U14924 (N_14924,N_11387,N_10633);
or U14925 (N_14925,N_11163,N_10779);
xor U14926 (N_14926,N_12105,N_10295);
xor U14927 (N_14927,N_11773,N_12178);
or U14928 (N_14928,N_11133,N_11046);
xor U14929 (N_14929,N_11290,N_11591);
or U14930 (N_14930,N_12098,N_10129);
nand U14931 (N_14931,N_10303,N_10153);
and U14932 (N_14932,N_10872,N_10880);
or U14933 (N_14933,N_11918,N_10980);
and U14934 (N_14934,N_12392,N_10839);
nand U14935 (N_14935,N_10289,N_11379);
nand U14936 (N_14936,N_11398,N_11386);
xor U14937 (N_14937,N_10144,N_11475);
and U14938 (N_14938,N_10457,N_12235);
and U14939 (N_14939,N_11405,N_11797);
and U14940 (N_14940,N_11872,N_10795);
or U14941 (N_14941,N_10327,N_12159);
nand U14942 (N_14942,N_11014,N_10201);
nor U14943 (N_14943,N_12430,N_12244);
nand U14944 (N_14944,N_10204,N_10241);
nand U14945 (N_14945,N_12219,N_10392);
nor U14946 (N_14946,N_10543,N_10706);
and U14947 (N_14947,N_11404,N_10110);
nor U14948 (N_14948,N_10901,N_12167);
nor U14949 (N_14949,N_11079,N_12475);
nand U14950 (N_14950,N_10087,N_11645);
and U14951 (N_14951,N_10354,N_11586);
xor U14952 (N_14952,N_10648,N_11913);
nand U14953 (N_14953,N_12148,N_10574);
xor U14954 (N_14954,N_10593,N_11383);
and U14955 (N_14955,N_11551,N_12472);
or U14956 (N_14956,N_12226,N_10385);
nand U14957 (N_14957,N_10214,N_11414);
and U14958 (N_14958,N_12176,N_10534);
or U14959 (N_14959,N_10281,N_10139);
nand U14960 (N_14960,N_11677,N_10521);
and U14961 (N_14961,N_12000,N_12115);
nand U14962 (N_14962,N_10167,N_12202);
or U14963 (N_14963,N_12154,N_11757);
and U14964 (N_14964,N_10125,N_11787);
nor U14965 (N_14965,N_11618,N_10770);
and U14966 (N_14966,N_10103,N_12138);
or U14967 (N_14967,N_10319,N_10027);
nor U14968 (N_14968,N_10584,N_11346);
and U14969 (N_14969,N_11278,N_11870);
nor U14970 (N_14970,N_10243,N_10837);
nor U14971 (N_14971,N_12102,N_11535);
nand U14972 (N_14972,N_10401,N_10908);
nand U14973 (N_14973,N_11640,N_11708);
and U14974 (N_14974,N_11171,N_11907);
nor U14975 (N_14975,N_12094,N_11254);
nor U14976 (N_14976,N_10142,N_11077);
nor U14977 (N_14977,N_11615,N_10622);
nand U14978 (N_14978,N_10572,N_10852);
and U14979 (N_14979,N_11840,N_10416);
and U14980 (N_14980,N_11165,N_11789);
and U14981 (N_14981,N_12264,N_11792);
or U14982 (N_14982,N_10733,N_10826);
nand U14983 (N_14983,N_10757,N_10752);
or U14984 (N_14984,N_10304,N_11371);
nor U14985 (N_14985,N_10649,N_11926);
and U14986 (N_14986,N_11337,N_10208);
or U14987 (N_14987,N_11187,N_10459);
nand U14988 (N_14988,N_11125,N_11398);
and U14989 (N_14989,N_10760,N_11124);
and U14990 (N_14990,N_12460,N_10233);
xnor U14991 (N_14991,N_11899,N_10044);
or U14992 (N_14992,N_10564,N_11780);
xnor U14993 (N_14993,N_12183,N_10492);
nand U14994 (N_14994,N_10612,N_11853);
and U14995 (N_14995,N_12326,N_11256);
nand U14996 (N_14996,N_10717,N_12423);
xor U14997 (N_14997,N_10885,N_11881);
nand U14998 (N_14998,N_10457,N_11868);
nand U14999 (N_14999,N_10798,N_11304);
xnor U15000 (N_15000,N_13139,N_14990);
nor U15001 (N_15001,N_13357,N_13621);
or U15002 (N_15002,N_13093,N_14316);
nand U15003 (N_15003,N_14218,N_13441);
nand U15004 (N_15004,N_13838,N_13678);
xnor U15005 (N_15005,N_12647,N_13985);
xor U15006 (N_15006,N_13405,N_12667);
xor U15007 (N_15007,N_14894,N_13920);
and U15008 (N_15008,N_14390,N_14452);
nand U15009 (N_15009,N_14784,N_14070);
nor U15010 (N_15010,N_13254,N_13005);
or U15011 (N_15011,N_12632,N_13645);
nand U15012 (N_15012,N_13746,N_14392);
or U15013 (N_15013,N_13435,N_13605);
nor U15014 (N_15014,N_13651,N_13411);
and U15015 (N_15015,N_12851,N_13065);
nand U15016 (N_15016,N_14360,N_13836);
or U15017 (N_15017,N_12803,N_13190);
nor U15018 (N_15018,N_13818,N_14629);
and U15019 (N_15019,N_13545,N_12823);
nand U15020 (N_15020,N_14225,N_14433);
nor U15021 (N_15021,N_13560,N_12703);
nor U15022 (N_15022,N_13146,N_14168);
nand U15023 (N_15023,N_12527,N_14746);
or U15024 (N_15024,N_14011,N_14807);
nand U15025 (N_15025,N_13789,N_14210);
xor U15026 (N_15026,N_12742,N_13499);
nor U15027 (N_15027,N_14416,N_14120);
or U15028 (N_15028,N_14823,N_12809);
nand U15029 (N_15029,N_14204,N_13439);
and U15030 (N_15030,N_12955,N_14454);
and U15031 (N_15031,N_13432,N_13693);
nor U15032 (N_15032,N_13768,N_14728);
or U15033 (N_15033,N_14613,N_13370);
or U15034 (N_15034,N_14959,N_13506);
or U15035 (N_15035,N_14975,N_13373);
nor U15036 (N_15036,N_12746,N_14662);
or U15037 (N_15037,N_14865,N_13116);
and U15038 (N_15038,N_12951,N_13736);
nor U15039 (N_15039,N_14526,N_14772);
nor U15040 (N_15040,N_13615,N_13383);
nand U15041 (N_15041,N_13387,N_13580);
and U15042 (N_15042,N_14558,N_14549);
xor U15043 (N_15043,N_14188,N_13951);
nor U15044 (N_15044,N_13346,N_13997);
nand U15045 (N_15045,N_12774,N_14207);
nor U15046 (N_15046,N_12971,N_13739);
xor U15047 (N_15047,N_12923,N_14541);
and U15048 (N_15048,N_14622,N_14939);
nor U15049 (N_15049,N_14814,N_12592);
nor U15050 (N_15050,N_13793,N_14035);
or U15051 (N_15051,N_13835,N_13422);
xor U15052 (N_15052,N_12677,N_13688);
nand U15053 (N_15053,N_12570,N_12624);
and U15054 (N_15054,N_13899,N_13164);
and U15055 (N_15055,N_14376,N_13378);
or U15056 (N_15056,N_14811,N_13077);
nand U15057 (N_15057,N_14647,N_13599);
or U15058 (N_15058,N_12692,N_13953);
nand U15059 (N_15059,N_13394,N_14005);
nand U15060 (N_15060,N_14295,N_13434);
nand U15061 (N_15061,N_13250,N_12590);
nor U15062 (N_15062,N_13616,N_13869);
nand U15063 (N_15063,N_14201,N_13348);
nand U15064 (N_15064,N_13052,N_13967);
xor U15065 (N_15065,N_14173,N_12858);
xnor U15066 (N_15066,N_13812,N_12710);
or U15067 (N_15067,N_13202,N_13750);
nand U15068 (N_15068,N_13037,N_13548);
or U15069 (N_15069,N_13981,N_14477);
and U15070 (N_15070,N_14147,N_12654);
or U15071 (N_15071,N_14040,N_14502);
and U15072 (N_15072,N_13440,N_12818);
xor U15073 (N_15073,N_14182,N_14481);
and U15074 (N_15074,N_13166,N_14162);
xor U15075 (N_15075,N_13617,N_13211);
xnor U15076 (N_15076,N_14785,N_12531);
or U15077 (N_15077,N_14391,N_14499);
and U15078 (N_15078,N_13721,N_13229);
xnor U15079 (N_15079,N_13050,N_14642);
nor U15080 (N_15080,N_13004,N_13889);
nor U15081 (N_15081,N_13263,N_13572);
and U15082 (N_15082,N_14634,N_14194);
and U15083 (N_15083,N_14554,N_14082);
nor U15084 (N_15084,N_13762,N_14289);
xor U15085 (N_15085,N_14023,N_12612);
xor U15086 (N_15086,N_14618,N_13126);
xor U15087 (N_15087,N_13109,N_12901);
or U15088 (N_15088,N_14298,N_14859);
nand U15089 (N_15089,N_12772,N_14770);
or U15090 (N_15090,N_14694,N_13948);
nand U15091 (N_15091,N_13452,N_12698);
or U15092 (N_15092,N_14432,N_12944);
or U15093 (N_15093,N_14179,N_13585);
xnor U15094 (N_15094,N_12670,N_14435);
nand U15095 (N_15095,N_14062,N_14738);
and U15096 (N_15096,N_12773,N_14445);
or U15097 (N_15097,N_13702,N_13151);
or U15098 (N_15098,N_13063,N_13171);
nor U15099 (N_15099,N_14209,N_13749);
xnor U15100 (N_15100,N_14570,N_14565);
and U15101 (N_15101,N_12618,N_14259);
or U15102 (N_15102,N_13220,N_13887);
and U15103 (N_15103,N_12568,N_14925);
and U15104 (N_15104,N_12837,N_13026);
xnor U15105 (N_15105,N_14880,N_13729);
and U15106 (N_15106,N_13543,N_14739);
nor U15107 (N_15107,N_14796,N_13541);
nor U15108 (N_15108,N_13701,N_13694);
or U15109 (N_15109,N_12821,N_13815);
or U15110 (N_15110,N_14441,N_13034);
or U15111 (N_15111,N_13053,N_14603);
and U15112 (N_15112,N_14235,N_13087);
nand U15113 (N_15113,N_14605,N_13113);
and U15114 (N_15114,N_13578,N_12894);
xnor U15115 (N_15115,N_14666,N_14981);
nand U15116 (N_15116,N_14913,N_13354);
and U15117 (N_15117,N_14032,N_12993);
and U15118 (N_15118,N_13949,N_13282);
xor U15119 (N_15119,N_12844,N_14742);
xnor U15120 (N_15120,N_14214,N_14363);
nand U15121 (N_15121,N_12928,N_13960);
xnor U15122 (N_15122,N_12672,N_14243);
nor U15123 (N_15123,N_12927,N_13567);
nor U15124 (N_15124,N_14639,N_14139);
nand U15125 (N_15125,N_13814,N_13510);
and U15126 (N_15126,N_13245,N_13880);
nor U15127 (N_15127,N_14868,N_13956);
xor U15128 (N_15128,N_14081,N_13242);
nand U15129 (N_15129,N_13462,N_12855);
nor U15130 (N_15130,N_14787,N_14923);
and U15131 (N_15131,N_13902,N_14596);
and U15132 (N_15132,N_14983,N_12545);
nor U15133 (N_15133,N_12700,N_12828);
and U15134 (N_15134,N_12929,N_13860);
nand U15135 (N_15135,N_14248,N_14468);
nand U15136 (N_15136,N_13662,N_13994);
xor U15137 (N_15137,N_13196,N_14906);
nand U15138 (N_15138,N_13963,N_14703);
or U15139 (N_15139,N_14440,N_13327);
and U15140 (N_15140,N_13003,N_14150);
nand U15141 (N_15141,N_14765,N_13241);
and U15142 (N_15142,N_14372,N_14050);
nand U15143 (N_15143,N_12924,N_13794);
nor U15144 (N_15144,N_12622,N_13057);
or U15145 (N_15145,N_13334,N_14776);
and U15146 (N_15146,N_14767,N_13144);
and U15147 (N_15147,N_13283,N_14510);
or U15148 (N_15148,N_13904,N_12899);
nand U15149 (N_15149,N_14698,N_12542);
nand U15150 (N_15150,N_13366,N_13643);
nand U15151 (N_15151,N_13816,N_14043);
nand U15152 (N_15152,N_13658,N_13316);
and U15153 (N_15153,N_14963,N_13009);
and U15154 (N_15154,N_13206,N_13727);
nand U15155 (N_15155,N_13284,N_13266);
nor U15156 (N_15156,N_12599,N_12921);
or U15157 (N_15157,N_13879,N_14783);
xnor U15158 (N_15158,N_12969,N_13954);
nand U15159 (N_15159,N_12872,N_14230);
or U15160 (N_15160,N_12782,N_14068);
nor U15161 (N_15161,N_13748,N_13251);
xor U15162 (N_15162,N_14985,N_13160);
nor U15163 (N_15163,N_13074,N_14004);
xnor U15164 (N_15164,N_13897,N_14223);
nand U15165 (N_15165,N_13006,N_13374);
nor U15166 (N_15166,N_13168,N_13186);
or U15167 (N_15167,N_12603,N_13000);
nor U15168 (N_15168,N_14991,N_14381);
xnor U15169 (N_15169,N_13569,N_14205);
nor U15170 (N_15170,N_14436,N_13337);
or U15171 (N_15171,N_14505,N_14616);
and U15172 (N_15172,N_14350,N_14934);
or U15173 (N_15173,N_14041,N_14573);
nor U15174 (N_15174,N_14020,N_14231);
or U15175 (N_15175,N_14863,N_14103);
or U15176 (N_15176,N_14443,N_14491);
or U15177 (N_15177,N_12549,N_13025);
xnor U15178 (N_15178,N_14273,N_13756);
nand U15179 (N_15179,N_13349,N_14780);
nor U15180 (N_15180,N_13197,N_13757);
xnor U15181 (N_15181,N_14816,N_14157);
xor U15182 (N_15182,N_14971,N_13318);
nand U15183 (N_15183,N_14351,N_12817);
and U15184 (N_15184,N_14083,N_14266);
nor U15185 (N_15185,N_13375,N_13330);
or U15186 (N_15186,N_14160,N_14946);
or U15187 (N_15187,N_13042,N_13248);
and U15188 (N_15188,N_12835,N_13663);
and U15189 (N_15189,N_14504,N_13331);
nor U15190 (N_15190,N_14855,N_13364);
xor U15191 (N_15191,N_13384,N_14430);
or U15192 (N_15192,N_14591,N_13158);
xnor U15193 (N_15193,N_14978,N_13149);
xnor U15194 (N_15194,N_14487,N_13922);
xor U15195 (N_15195,N_14801,N_13226);
nor U15196 (N_15196,N_12995,N_12753);
and U15197 (N_15197,N_14951,N_12505);
xnor U15198 (N_15198,N_13563,N_14352);
or U15199 (N_15199,N_13068,N_14361);
xnor U15200 (N_15200,N_14878,N_12903);
nand U15201 (N_15201,N_13966,N_13041);
nor U15202 (N_15202,N_13368,N_12501);
nand U15203 (N_15203,N_13315,N_13217);
or U15204 (N_15204,N_14754,N_14810);
xnor U15205 (N_15205,N_13105,N_13905);
nand U15206 (N_15206,N_13517,N_14800);
and U15207 (N_15207,N_14084,N_12714);
and U15208 (N_15208,N_13177,N_12644);
nand U15209 (N_15209,N_14531,N_12546);
xor U15210 (N_15210,N_13076,N_14299);
xnor U15211 (N_15211,N_13033,N_14815);
and U15212 (N_15212,N_12631,N_13010);
and U15213 (N_15213,N_12691,N_13270);
xor U15214 (N_15214,N_13565,N_14701);
nor U15215 (N_15215,N_14842,N_12634);
and U15216 (N_15216,N_12966,N_13015);
and U15217 (N_15217,N_13125,N_13573);
nand U15218 (N_15218,N_13436,N_14314);
or U15219 (N_15219,N_14415,N_14654);
nor U15220 (N_15220,N_13021,N_13131);
xnor U15221 (N_15221,N_13401,N_13653);
or U15222 (N_15222,N_14095,N_14300);
and U15223 (N_15223,N_12619,N_14106);
and U15224 (N_15224,N_13511,N_14253);
nand U15225 (N_15225,N_14237,N_14758);
and U15226 (N_15226,N_14323,N_14533);
or U15227 (N_15227,N_13863,N_13508);
xor U15228 (N_15228,N_14485,N_13124);
or U15229 (N_15229,N_13408,N_12931);
and U15230 (N_15230,N_14385,N_14707);
and U15231 (N_15231,N_13837,N_13278);
and U15232 (N_15232,N_13145,N_13194);
and U15233 (N_15233,N_12932,N_12876);
xnor U15234 (N_15234,N_13853,N_14552);
or U15235 (N_15235,N_13800,N_13095);
or U15236 (N_15236,N_13728,N_13473);
xor U15237 (N_15237,N_13449,N_13970);
and U15238 (N_15238,N_13872,N_13276);
xor U15239 (N_15239,N_14817,N_14841);
xor U15240 (N_15240,N_14755,N_12831);
nor U15241 (N_15241,N_14358,N_13821);
and U15242 (N_15242,N_13478,N_14013);
or U15243 (N_15243,N_13342,N_12860);
or U15244 (N_15244,N_13649,N_12567);
or U15245 (N_15245,N_13100,N_14178);
and U15246 (N_15246,N_14760,N_12511);
nand U15247 (N_15247,N_14546,N_13118);
xnor U15248 (N_15248,N_14211,N_14753);
nand U15249 (N_15249,N_14805,N_12541);
and U15250 (N_15250,N_13751,N_14910);
xor U15251 (N_15251,N_12947,N_13082);
xnor U15252 (N_15252,N_13907,N_14635);
xnor U15253 (N_15253,N_13895,N_13367);
or U15254 (N_15254,N_12940,N_14292);
nand U15255 (N_15255,N_13603,N_14034);
nand U15256 (N_15256,N_12681,N_13822);
nand U15257 (N_15257,N_14625,N_12968);
nand U15258 (N_15258,N_13426,N_12979);
nand U15259 (N_15259,N_14079,N_12583);
nand U15260 (N_15260,N_14821,N_12723);
and U15261 (N_15261,N_13681,N_13371);
or U15262 (N_15262,N_13820,N_14886);
nor U15263 (N_15263,N_14076,N_14170);
or U15264 (N_15264,N_12608,N_13667);
or U15265 (N_15265,N_13023,N_14402);
or U15266 (N_15266,N_12830,N_14216);
nand U15267 (N_15267,N_14690,N_12640);
xor U15268 (N_15268,N_12715,N_14164);
and U15269 (N_15269,N_12999,N_13154);
and U15270 (N_15270,N_12617,N_12606);
xnor U15271 (N_15271,N_14759,N_13112);
and U15272 (N_15272,N_13598,N_13137);
or U15273 (N_15273,N_13081,N_14031);
nor U15274 (N_15274,N_13244,N_13141);
xor U15275 (N_15275,N_14832,N_14145);
and U15276 (N_15276,N_12996,N_12638);
nor U15277 (N_15277,N_13873,N_14893);
and U15278 (N_15278,N_12516,N_14954);
nor U15279 (N_15279,N_14217,N_14039);
and U15280 (N_15280,N_13036,N_13410);
and U15281 (N_15281,N_12810,N_14389);
and U15282 (N_15282,N_14782,N_13634);
nor U15283 (N_15283,N_12904,N_14597);
nor U15284 (N_15284,N_14332,N_13533);
nor U15285 (N_15285,N_14538,N_12633);
nor U15286 (N_15286,N_13490,N_13304);
and U15287 (N_15287,N_13183,N_13403);
and U15288 (N_15288,N_14046,N_13810);
or U15289 (N_15289,N_13461,N_13896);
nor U15290 (N_15290,N_13256,N_12839);
or U15291 (N_15291,N_13471,N_13636);
nor U15292 (N_15292,N_12561,N_12941);
or U15293 (N_15293,N_14420,N_13841);
xor U15294 (N_15294,N_14268,N_14374);
xor U15295 (N_15295,N_12641,N_14723);
nand U15296 (N_15296,N_13683,N_12643);
xnor U15297 (N_15297,N_14885,N_14426);
nor U15298 (N_15298,N_12659,N_14640);
xnor U15299 (N_15299,N_13279,N_14980);
nand U15300 (N_15300,N_14996,N_12768);
nor U15301 (N_15301,N_14064,N_12560);
xnor U15302 (N_15302,N_13732,N_14220);
xor U15303 (N_15303,N_13445,N_14924);
nand U15304 (N_15304,N_13507,N_14709);
and U15305 (N_15305,N_12987,N_13265);
and U15306 (N_15306,N_14444,N_14525);
xor U15307 (N_15307,N_12885,N_13798);
nand U15308 (N_15308,N_13935,N_14949);
nor U15309 (N_15309,N_12967,N_12558);
nor U15310 (N_15310,N_13467,N_14366);
nor U15311 (N_15311,N_14623,N_12792);
xor U15312 (N_15312,N_12827,N_13633);
and U15313 (N_15313,N_14492,N_12735);
nand U15314 (N_15314,N_13215,N_14371);
nand U15315 (N_15315,N_14917,N_12708);
and U15316 (N_15316,N_14853,N_14187);
xor U15317 (N_15317,N_12796,N_13776);
or U15318 (N_15318,N_13819,N_13677);
nor U15319 (N_15319,N_12676,N_13858);
or U15320 (N_15320,N_13952,N_14101);
nand U15321 (N_15321,N_12933,N_13919);
or U15322 (N_15322,N_14921,N_12994);
and U15323 (N_15323,N_14620,N_12520);
nor U15324 (N_15324,N_13574,N_14343);
nand U15325 (N_15325,N_14892,N_14711);
nor U15326 (N_15326,N_14691,N_13885);
and U15327 (N_15327,N_13546,N_14852);
and U15328 (N_15328,N_13385,N_13165);
xor U15329 (N_15329,N_13671,N_13641);
nand U15330 (N_15330,N_14524,N_13613);
nor U15331 (N_15331,N_14246,N_13965);
nand U15332 (N_15332,N_12820,N_13783);
nand U15333 (N_15333,N_14045,N_14519);
or U15334 (N_15334,N_13421,N_13995);
nor U15335 (N_15335,N_14534,N_13011);
nand U15336 (N_15336,N_12757,N_12939);
nand U15337 (N_15337,N_14869,N_14667);
and U15338 (N_15338,N_14850,N_13386);
xnor U15339 (N_15339,N_14422,N_13456);
xor U15340 (N_15340,N_13365,N_12635);
nand U15341 (N_15341,N_12816,N_12630);
and U15342 (N_15342,N_12705,N_13538);
nor U15343 (N_15343,N_14447,N_13975);
xor U15344 (N_15344,N_12719,N_13657);
xor U15345 (N_15345,N_13531,N_14812);
xor U15346 (N_15346,N_14875,N_14387);
and U15347 (N_15347,N_12988,N_13347);
or U15348 (N_15348,N_14606,N_12850);
and U15349 (N_15349,N_14719,N_14724);
xnor U15350 (N_15350,N_14896,N_12732);
nand U15351 (N_15351,N_13259,N_13974);
or U15352 (N_15352,N_13619,N_14152);
and U15353 (N_15353,N_14475,N_13909);
and U15354 (N_15354,N_13635,N_14583);
or U15355 (N_15355,N_13670,N_14818);
and U15356 (N_15356,N_13260,N_13504);
nand U15357 (N_15357,N_13515,N_14979);
xnor U15358 (N_15358,N_13884,N_12749);
nand U15359 (N_15359,N_13479,N_12865);
nand U15360 (N_15360,N_13703,N_14668);
or U15361 (N_15361,N_13391,N_13584);
xor U15362 (N_15362,N_14891,N_14966);
nand U15363 (N_15363,N_14055,N_12862);
xnor U15364 (N_15364,N_14423,N_14748);
or U15365 (N_15365,N_13308,N_14324);
or U15366 (N_15366,N_13274,N_13272);
and U15367 (N_15367,N_13632,N_13514);
nor U15368 (N_15368,N_12764,N_13993);
nor U15369 (N_15369,N_14633,N_14771);
and U15370 (N_15370,N_14998,N_12965);
nor U15371 (N_15371,N_12978,N_14108);
or U15372 (N_15372,N_12896,N_14294);
and U15373 (N_15373,N_13937,N_14912);
xnor U15374 (N_15374,N_13285,N_13071);
and U15375 (N_15375,N_12945,N_13682);
and U15376 (N_15376,N_12954,N_13777);
and U15377 (N_15377,N_13831,N_14143);
nor U15378 (N_15378,N_13811,N_14888);
or U15379 (N_15379,N_14006,N_13734);
nand U15380 (N_15380,N_13420,N_13390);
or U15381 (N_15381,N_13022,N_14594);
nor U15382 (N_15382,N_13977,N_14290);
nand U15383 (N_15383,N_14421,N_13428);
or U15384 (N_15384,N_13048,N_13163);
or U15385 (N_15385,N_14641,N_12841);
xor U15386 (N_15386,N_14676,N_13908);
or U15387 (N_15387,N_12806,N_12551);
nand U15388 (N_15388,N_13827,N_12625);
nor U15389 (N_15389,N_12696,N_12997);
xnor U15390 (N_15390,N_14601,N_14825);
xnor U15391 (N_15391,N_14022,N_13520);
xnor U15392 (N_15392,N_14099,N_13972);
or U15393 (N_15393,N_13759,N_14944);
and U15394 (N_15394,N_12819,N_13301);
xnor U15395 (N_15395,N_14488,N_14568);
and U15396 (N_15396,N_13059,N_14911);
xnor U15397 (N_15397,N_12871,N_12961);
or U15398 (N_15398,N_13817,N_12540);
and U15399 (N_15399,N_13224,N_14977);
or U15400 (N_15400,N_14689,N_12759);
nand U15401 (N_15401,N_14321,N_12727);
nor U15402 (N_15402,N_14592,N_14061);
and U15403 (N_15403,N_13659,N_12736);
and U15404 (N_15404,N_14014,N_13212);
or U15405 (N_15405,N_14704,N_14950);
or U15406 (N_15406,N_14529,N_13551);
nor U15407 (N_15407,N_12623,N_13468);
nor U15408 (N_15408,N_13766,N_12747);
nor U15409 (N_15409,N_14686,N_14769);
nor U15410 (N_15410,N_12521,N_12536);
nor U15411 (N_15411,N_13856,N_13110);
xnor U15412 (N_15412,N_14111,N_13291);
xor U15413 (N_15413,N_12718,N_13236);
nor U15414 (N_15414,N_12610,N_14283);
or U15415 (N_15415,N_13665,N_14523);
or U15416 (N_15416,N_13200,N_14631);
or U15417 (N_15417,N_12574,N_13961);
nor U15418 (N_15418,N_13775,N_12778);
and U15419 (N_15419,N_13135,N_13988);
nor U15420 (N_15420,N_12548,N_13791);
and U15421 (N_15421,N_14750,N_14658);
or U15422 (N_15422,N_13950,N_14446);
nor U15423 (N_15423,N_14947,N_14274);
and U15424 (N_15424,N_14213,N_12573);
xnor U15425 (N_15425,N_14241,N_14916);
or U15426 (N_15426,N_13877,N_14184);
xnor U15427 (N_15427,N_13028,N_13295);
or U15428 (N_15428,N_13795,N_14506);
and U15429 (N_15429,N_13313,N_14189);
xor U15430 (N_15430,N_12842,N_13894);
xor U15431 (N_15431,N_14478,N_14437);
or U15432 (N_15432,N_14405,N_14429);
or U15433 (N_15433,N_13724,N_14650);
or U15434 (N_15434,N_13142,N_13602);
or U15435 (N_15435,N_13881,N_14887);
nand U15436 (N_15436,N_14589,N_14411);
nand U15437 (N_15437,N_14696,N_12506);
xnor U15438 (N_15438,N_14325,N_14078);
nor U15439 (N_15439,N_14109,N_12614);
or U15440 (N_15440,N_13476,N_12777);
or U15441 (N_15441,N_14500,N_12717);
or U15442 (N_15442,N_14590,N_14119);
or U15443 (N_15443,N_14795,N_13097);
and U15444 (N_15444,N_13503,N_12722);
nand U15445 (N_15445,N_14773,N_13398);
xor U15446 (N_15446,N_14535,N_14219);
xor U15447 (N_15447,N_12713,N_12946);
xnor U15448 (N_15448,N_13044,N_13704);
nor U15449 (N_15449,N_14705,N_13485);
and U15450 (N_15450,N_14155,N_13870);
nand U15451 (N_15451,N_12678,N_12563);
and U15452 (N_15452,N_14907,N_14370);
nand U15453 (N_15453,N_13193,N_14542);
or U15454 (N_15454,N_14651,N_12991);
or U15455 (N_15455,N_13073,N_12970);
or U15456 (N_15456,N_14905,N_13646);
nand U15457 (N_15457,N_14025,N_13427);
xnor U15458 (N_15458,N_12507,N_12911);
and U15459 (N_15459,N_12581,N_12986);
xnor U15460 (N_15460,N_14560,N_14964);
or U15461 (N_15461,N_14958,N_13292);
or U15462 (N_15462,N_13806,N_14261);
xor U15463 (N_15463,N_14749,N_13223);
or U15464 (N_15464,N_13733,N_14834);
or U15465 (N_15465,N_12751,N_12985);
nor U15466 (N_15466,N_14090,N_13188);
and U15467 (N_15467,N_12528,N_14427);
or U15468 (N_15468,N_12565,N_13344);
xor U15469 (N_15469,N_13013,N_14918);
nor U15470 (N_15470,N_13941,N_12913);
or U15471 (N_15471,N_14379,N_13940);
nor U15472 (N_15472,N_13147,N_13589);
xor U15473 (N_15473,N_14265,N_13715);
nor U15474 (N_15474,N_13890,N_12600);
or U15475 (N_15475,N_12656,N_13361);
or U15476 (N_15476,N_14074,N_14607);
nand U15477 (N_15477,N_14576,N_14098);
or U15478 (N_15478,N_13779,N_13393);
or U15479 (N_15479,N_14028,N_14610);
nor U15480 (N_15480,N_12585,N_14382);
nor U15481 (N_15481,N_12509,N_12725);
nor U15482 (N_15482,N_14140,N_14751);
nor U15483 (N_15483,N_14763,N_12653);
xnor U15484 (N_15484,N_12651,N_12586);
xnor U15485 (N_15485,N_14581,N_13288);
nor U15486 (N_15486,N_13232,N_13329);
nand U15487 (N_15487,N_12992,N_14956);
nor U15488 (N_15488,N_14860,N_13720);
nand U15489 (N_15489,N_14858,N_14497);
and U15490 (N_15490,N_12642,N_13130);
and U15491 (N_15491,N_13257,N_14515);
and U15492 (N_15492,N_13607,N_13355);
or U15493 (N_15493,N_12752,N_14472);
nor U15494 (N_15494,N_14000,N_13017);
xnor U15495 (N_15495,N_13218,N_12662);
nor U15496 (N_15496,N_12980,N_14279);
or U15497 (N_15497,N_14967,N_13416);
xnor U15498 (N_15498,N_12834,N_13415);
nand U15499 (N_15499,N_13958,N_14926);
and U15500 (N_15500,N_13335,N_14344);
nand U15501 (N_15501,N_14333,N_12766);
nor U15502 (N_15502,N_12787,N_13929);
and U15503 (N_15503,N_14367,N_14752);
nand U15504 (N_15504,N_14786,N_12729);
or U15505 (N_15505,N_12878,N_12524);
and U15506 (N_15506,N_13305,N_12925);
and U15507 (N_15507,N_14054,N_14383);
or U15508 (N_15508,N_13433,N_14598);
and U15509 (N_15509,N_12731,N_12891);
nand U15510 (N_15510,N_14208,N_13417);
nor U15511 (N_15511,N_14609,N_14224);
nand U15512 (N_15512,N_14970,N_13859);
nand U15513 (N_15513,N_13099,N_14368);
and U15514 (N_15514,N_14007,N_13129);
or U15515 (N_15515,N_13611,N_12918);
xor U15516 (N_15516,N_14362,N_14577);
nand U15517 (N_15517,N_12769,N_12857);
and U15518 (N_15518,N_14038,N_14085);
xor U15519 (N_15519,N_14718,N_14089);
nand U15520 (N_15520,N_13523,N_13134);
nand U15521 (N_15521,N_14612,N_13045);
nor U15522 (N_15522,N_13512,N_13608);
or U15523 (N_15523,N_14854,N_14192);
nand U15524 (N_15524,N_13321,N_12569);
nand U15525 (N_15525,N_14992,N_13927);
nor U15526 (N_15526,N_14047,N_13092);
nor U15527 (N_15527,N_13978,N_14646);
and U15528 (N_15528,N_14669,N_13209);
and U15529 (N_15529,N_13119,N_13453);
or U15530 (N_15530,N_13309,N_13418);
and U15531 (N_15531,N_12897,N_14969);
nand U15532 (N_15532,N_12982,N_12781);
xor U15533 (N_15533,N_13700,N_12706);
and U15534 (N_15534,N_13592,N_12895);
xor U15535 (N_15535,N_14730,N_14808);
nor U15536 (N_15536,N_14473,N_14940);
nand U15537 (N_15537,N_13735,N_13983);
xnor U15538 (N_15538,N_14001,N_13055);
xnor U15539 (N_15539,N_13429,N_14569);
and U15540 (N_15540,N_14938,N_13326);
xnor U15541 (N_15541,N_14114,N_13012);
or U15542 (N_15542,N_13302,N_13926);
and U15543 (N_15543,N_12881,N_14086);
and U15544 (N_15544,N_13764,N_14928);
nor U15545 (N_15545,N_13489,N_14044);
and U15546 (N_15546,N_14574,N_13802);
or U15547 (N_15547,N_13943,N_14469);
xor U15548 (N_15548,N_12790,N_13123);
nor U15549 (N_15549,N_14424,N_12956);
nor U15550 (N_15550,N_13002,N_12663);
xor U15551 (N_15551,N_14355,N_13491);
and U15552 (N_15552,N_13201,N_13945);
nor U15553 (N_15553,N_13402,N_13656);
and U15554 (N_15554,N_14288,N_12906);
xor U15555 (N_15555,N_12646,N_13345);
xnor U15556 (N_15556,N_14263,N_14799);
nand U15557 (N_15557,N_14318,N_12660);
and U15558 (N_15558,N_12959,N_13207);
nand U15559 (N_15559,N_12902,N_14131);
and U15560 (N_15560,N_14584,N_13898);
and U15561 (N_15561,N_13618,N_13339);
xor U15562 (N_15562,N_12989,N_13901);
or U15563 (N_15563,N_13501,N_14675);
xnor U15564 (N_15564,N_13552,N_12519);
and U15565 (N_15565,N_14661,N_14024);
xor U15566 (N_15566,N_13356,N_12877);
nor U15567 (N_15567,N_13340,N_13064);
or U15568 (N_15568,N_13891,N_13472);
and U15569 (N_15569,N_13576,N_13180);
nand U15570 (N_15570,N_14448,N_12712);
or U15571 (N_15571,N_14556,N_14494);
and U15572 (N_15572,N_14655,N_12613);
or U15573 (N_15573,N_14281,N_14883);
or U15574 (N_15574,N_12566,N_12649);
xor U15575 (N_15575,N_13989,N_14678);
or U15576 (N_15576,N_14521,N_13593);
or U15577 (N_15577,N_14809,N_13024);
and U15578 (N_15578,N_12539,N_14196);
or U15579 (N_15579,N_12533,N_14334);
xnor U15580 (N_15580,N_14864,N_13079);
and U15581 (N_15581,N_13781,N_13866);
xor U15582 (N_15582,N_13824,N_13392);
or U15583 (N_15583,N_14792,N_14240);
and U15584 (N_15584,N_14460,N_13638);
and U15585 (N_15585,N_14575,N_14471);
nand U15586 (N_15586,N_12544,N_14404);
and U15587 (N_15587,N_14551,N_14797);
and U15588 (N_15588,N_14063,N_13406);
xnor U15589 (N_15589,N_12593,N_13400);
nand U15590 (N_15590,N_13103,N_12577);
nor U15591 (N_15591,N_14774,N_14904);
xor U15592 (N_15592,N_13723,N_13808);
and U15593 (N_15593,N_14158,N_14493);
xor U15594 (N_15594,N_14375,N_14806);
nor U15595 (N_15595,N_14929,N_12576);
nand U15596 (N_15596,N_14922,N_13362);
nand U15597 (N_15597,N_12780,N_14997);
or U15598 (N_15598,N_12887,N_14331);
or U15599 (N_15599,N_13829,N_13469);
and U15600 (N_15600,N_14483,N_13360);
nand U15601 (N_15601,N_13431,N_14315);
or U15602 (N_15602,N_13388,N_13091);
or U15603 (N_15603,N_14269,N_13219);
xnor U15604 (N_15604,N_13240,N_12733);
nand U15605 (N_15605,N_14463,N_14789);
nand U15606 (N_15606,N_14303,N_13062);
nand U15607 (N_15607,N_14663,N_12808);
or U15608 (N_15608,N_14710,N_13181);
nor U15609 (N_15609,N_13979,N_14136);
or U15610 (N_15610,N_12615,N_14457);
or U15611 (N_15611,N_14112,N_14093);
or U15612 (N_15612,N_14071,N_13871);
xnor U15613 (N_15613,N_13857,N_13610);
or U15614 (N_15614,N_13085,N_14304);
nor U15615 (N_15615,N_14313,N_14262);
nor U15616 (N_15616,N_14102,N_13121);
xnor U15617 (N_15617,N_14251,N_14995);
xor U15618 (N_15618,N_13397,N_14931);
and U15619 (N_15619,N_13570,N_13851);
xnor U15620 (N_15620,N_12503,N_14764);
nand U15621 (N_15621,N_14636,N_14087);
and U15622 (N_15622,N_13018,N_12760);
and U15623 (N_15623,N_13369,N_14348);
nand U15624 (N_15624,N_14509,N_14388);
xor U15625 (N_15625,N_14861,N_14465);
xor U15626 (N_15626,N_13848,N_14403);
and U15627 (N_15627,N_13622,N_14930);
and U15628 (N_15628,N_13492,N_14968);
nor U15629 (N_15629,N_13786,N_13101);
and U15630 (N_15630,N_14973,N_14238);
nor U15631 (N_15631,N_13550,N_12750);
or U15632 (N_15632,N_14067,N_14747);
and U15633 (N_15633,N_13143,N_13443);
and U15634 (N_15634,N_14960,N_12591);
nor U15635 (N_15635,N_12682,N_13535);
nand U15636 (N_15636,N_14122,N_13293);
xor U15637 (N_15637,N_14015,N_13625);
xnor U15638 (N_15638,N_14229,N_12795);
nor U15639 (N_15639,N_14125,N_13187);
or U15640 (N_15640,N_12500,N_12801);
and U15641 (N_15641,N_12550,N_12789);
or U15642 (N_15642,N_13271,N_12976);
nand U15643 (N_15643,N_13054,N_13275);
nand U15644 (N_15644,N_14008,N_13558);
or U15645 (N_15645,N_12597,N_13785);
xor U15646 (N_15646,N_14993,N_12765);
or U15647 (N_15647,N_13990,N_14359);
or U15648 (N_15648,N_12711,N_14110);
and U15649 (N_15649,N_12595,N_14715);
or U15650 (N_15650,N_13912,N_12856);
or U15651 (N_15651,N_14075,N_14721);
nor U15652 (N_15652,N_14245,N_14664);
or U15653 (N_15653,N_12579,N_13609);
nand U15654 (N_15654,N_14398,N_14222);
xnor U15655 (N_15655,N_14827,N_13767);
nor U15656 (N_15656,N_12611,N_14909);
nand U15657 (N_15657,N_14982,N_14884);
nor U15658 (N_15658,N_12972,N_13067);
nor U15659 (N_15659,N_13019,N_14898);
xor U15660 (N_15660,N_13205,N_14165);
xor U15661 (N_15661,N_12699,N_12843);
or U15662 (N_15662,N_14582,N_13483);
or U15663 (N_15663,N_13711,N_12832);
or U15664 (N_15664,N_13098,N_13932);
and U15665 (N_15665,N_12580,N_14682);
and U15666 (N_15666,N_13564,N_13454);
or U15667 (N_15667,N_13685,N_14354);
nor U15668 (N_15668,N_13088,N_12794);
nor U15669 (N_15669,N_13117,N_13001);
or U15670 (N_15670,N_12907,N_13962);
nor U15671 (N_15671,N_14802,N_14221);
and U15672 (N_15672,N_13038,N_14660);
or U15673 (N_15673,N_13807,N_14994);
xor U15674 (N_15674,N_14935,N_13716);
nand U15675 (N_15675,N_13253,N_14672);
nor U15676 (N_15676,N_12661,N_14227);
nand U15677 (N_15677,N_12754,N_13106);
nor U15678 (N_15678,N_13992,N_13277);
or U15679 (N_15679,N_13828,N_14459);
and U15680 (N_15680,N_12833,N_13849);
and U15681 (N_15681,N_14737,N_12804);
xor U15682 (N_15682,N_14937,N_14735);
nor U15683 (N_15683,N_12626,N_13933);
or U15684 (N_15684,N_12892,N_12917);
nand U15685 (N_15685,N_13225,N_13070);
and U15686 (N_15686,N_14804,N_13519);
nand U15687 (N_15687,N_12589,N_13726);
nor U15688 (N_15688,N_13122,N_13539);
xor U15689 (N_15689,N_14595,N_14673);
xor U15690 (N_15690,N_13676,N_14518);
nand U15691 (N_15691,N_13404,N_13695);
nor U15692 (N_15692,N_14113,N_13864);
and U15693 (N_15693,N_14626,N_13549);
and U15694 (N_15694,N_13928,N_14345);
or U15695 (N_15695,N_12952,N_14722);
xor U15696 (N_15696,N_13999,N_12936);
and U15697 (N_15697,N_13547,N_14226);
xnor U15698 (N_15698,N_12762,N_14461);
or U15699 (N_15699,N_13114,N_14181);
xor U15700 (N_15700,N_12534,N_13934);
or U15701 (N_15701,N_14734,N_14425);
nor U15702 (N_15702,N_13046,N_14408);
or U15703 (N_15703,N_14700,N_14185);
xnor U15704 (N_15704,N_12884,N_13846);
and U15705 (N_15705,N_12879,N_14681);
or U15706 (N_15706,N_13155,N_14151);
xnor U15707 (N_15707,N_14881,N_12826);
xor U15708 (N_15708,N_14779,N_14037);
nor U15709 (N_15709,N_13475,N_13148);
xor U15710 (N_15710,N_13032,N_13596);
nor U15711 (N_15711,N_14547,N_13203);
nor U15712 (N_15712,N_14824,N_12673);
nor U15713 (N_15713,N_14908,N_13796);
xor U15714 (N_15714,N_14234,N_13661);
nor U15715 (N_15715,N_13247,N_14708);
and U15716 (N_15716,N_12822,N_13246);
nand U15717 (N_15717,N_14154,N_13458);
and U15718 (N_15718,N_14149,N_14486);
and U15719 (N_15719,N_13424,N_13923);
nor U15720 (N_15720,N_13184,N_12522);
or U15721 (N_15721,N_12724,N_13921);
or U15722 (N_15722,N_14470,N_13069);
and U15723 (N_15723,N_14346,N_14790);
nand U15724 (N_15724,N_14857,N_12824);
xnor U15725 (N_15725,N_12767,N_12547);
nor U15726 (N_15726,N_13679,N_14585);
nand U15727 (N_15727,N_14056,N_14564);
nand U15728 (N_15728,N_13938,N_12686);
nor U15729 (N_15729,N_13799,N_14271);
nand U15730 (N_15730,N_14396,N_14123);
nand U15731 (N_15731,N_13918,N_14394);
nand U15732 (N_15732,N_14745,N_12665);
nor U15733 (N_15733,N_13761,N_14604);
xor U15734 (N_15734,N_14148,N_14495);
nand U15735 (N_15735,N_13874,N_13505);
or U15736 (N_15736,N_13030,N_13413);
nand U15737 (N_15737,N_14828,N_13460);
and U15738 (N_15738,N_13911,N_14693);
and U15739 (N_15739,N_12990,N_14830);
nor U15740 (N_15740,N_14260,N_14116);
nor U15741 (N_15741,N_14026,N_14528);
nand U15742 (N_15742,N_12845,N_14729);
xnor U15743 (N_15743,N_14835,N_13668);
nand U15744 (N_15744,N_14999,N_13568);
nand U15745 (N_15745,N_14066,N_13738);
and U15746 (N_15746,N_14456,N_12883);
or U15747 (N_15747,N_14309,N_14511);
nor U15748 (N_15748,N_13561,N_14627);
nor U15749 (N_15749,N_13089,N_14128);
nand U15750 (N_15750,N_12697,N_14322);
or U15751 (N_15751,N_14280,N_14349);
nand U15752 (N_15752,N_12755,N_13612);
or U15753 (N_15753,N_14899,N_14902);
xor U15754 (N_15754,N_13299,N_12588);
xor U15755 (N_15755,N_14927,N_14876);
or U15756 (N_15756,N_13773,N_13830);
or U15757 (N_15757,N_13035,N_13650);
nand U15758 (N_15758,N_12629,N_14513);
nand U15759 (N_15759,N_14480,N_12874);
xnor U15760 (N_15760,N_12882,N_14308);
and U15761 (N_15761,N_12815,N_13111);
nor U15762 (N_15762,N_14166,N_13423);
xnor U15763 (N_15763,N_14193,N_12934);
nand U15764 (N_15764,N_14826,N_14820);
and U15765 (N_15765,N_13844,N_13832);
xor U15766 (N_15766,N_14353,N_14692);
nand U15767 (N_15767,N_14153,N_14545);
and U15768 (N_15768,N_14016,N_14256);
xnor U15769 (N_15769,N_12805,N_12707);
xor U15770 (N_15770,N_14870,N_12849);
nor U15771 (N_15771,N_14048,N_12846);
nor U15772 (N_15772,N_12974,N_14890);
or U15773 (N_15773,N_13078,N_14232);
or U15774 (N_15774,N_12518,N_14236);
nand U15775 (N_15775,N_14733,N_14503);
or U15776 (N_15776,N_12607,N_14972);
xnor U15777 (N_15777,N_13058,N_14600);
or U15778 (N_15778,N_13480,N_12825);
xnor U15779 (N_15779,N_14134,N_12800);
nand U15780 (N_15780,N_13620,N_13982);
and U15781 (N_15781,N_13376,N_14611);
xor U15782 (N_15782,N_13379,N_12889);
or U15783 (N_15783,N_14418,N_13481);
and U15784 (N_15784,N_14163,N_13522);
nand U15785 (N_15785,N_12709,N_13778);
or U15786 (N_15786,N_14176,N_14839);
nor U15787 (N_15787,N_13900,N_13231);
nor U15788 (N_15788,N_13273,N_14788);
nor U15789 (N_15789,N_14837,N_12598);
xor U15790 (N_15790,N_14732,N_14100);
and U15791 (N_15791,N_14702,N_13698);
xor U15792 (N_15792,N_13628,N_12942);
and U15793 (N_15793,N_12508,N_12813);
xor U15794 (N_15794,N_12915,N_12687);
or U15795 (N_15795,N_13104,N_14027);
or U15796 (N_15796,N_12738,N_13639);
or U15797 (N_15797,N_13128,N_13591);
xor U15798 (N_15798,N_12922,N_13446);
nand U15799 (N_15799,N_13823,N_13850);
xor U15800 (N_15800,N_12745,N_12587);
or U15801 (N_15801,N_13644,N_14987);
nand U15802 (N_15802,N_13396,N_12620);
nand U15803 (N_15803,N_12880,N_12728);
nor U15804 (N_15804,N_14697,N_12758);
nor U15805 (N_15805,N_14104,N_13772);
and U15806 (N_15806,N_14657,N_13765);
and U15807 (N_15807,N_14052,N_13243);
or U15808 (N_15808,N_14397,N_12636);
or U15809 (N_15809,N_13840,N_13096);
or U15810 (N_15810,N_14286,N_14726);
and U15811 (N_15811,N_14539,N_12785);
and U15812 (N_15812,N_13233,N_14798);
or U15813 (N_15813,N_13199,N_12984);
and U15814 (N_15814,N_13680,N_12680);
xor U15815 (N_15815,N_12900,N_14490);
or U15816 (N_15816,N_14901,N_14129);
or U15817 (N_15817,N_14339,N_14267);
nor U15818 (N_15818,N_12893,N_12788);
nand U15819 (N_15819,N_13500,N_13675);
and U15820 (N_15820,N_14932,N_14637);
nor U15821 (N_15821,N_12775,N_13906);
nor U15822 (N_15822,N_13984,N_13939);
or U15823 (N_15823,N_13351,N_13300);
nor U15824 (N_15824,N_14974,N_13865);
nand U15825 (N_15825,N_14498,N_14451);
nor U15826 (N_15826,N_13752,N_12556);
nor U15827 (N_15827,N_13731,N_13524);
xnor U15828 (N_15828,N_14761,N_13448);
nor U15829 (N_15829,N_13261,N_13630);
and U15830 (N_15830,N_14347,N_12962);
nor U15831 (N_15831,N_14778,N_13297);
or U15832 (N_15832,N_13708,N_13132);
xnor U15833 (N_15833,N_12734,N_13915);
nand U15834 (N_15834,N_13986,N_12875);
nor U15835 (N_15835,N_14097,N_13172);
and U15836 (N_15836,N_13710,N_14848);
nand U15837 (N_15837,N_14141,N_13660);
nand U15838 (N_15838,N_13319,N_13627);
nand U15839 (N_15839,N_14307,N_14593);
nor U15840 (N_15840,N_13060,N_13213);
nand U15841 (N_15841,N_13447,N_13488);
nand U15842 (N_15842,N_13162,N_13287);
nor U15843 (N_15843,N_14228,N_14021);
nor U15844 (N_15844,N_12510,N_14175);
or U15845 (N_15845,N_14118,N_14638);
or U15846 (N_15846,N_12601,N_13640);
nor U15847 (N_15847,N_12683,N_13537);
xor U15848 (N_15848,N_14687,N_13372);
and U15849 (N_15849,N_13380,N_12829);
nor U15850 (N_15850,N_14665,N_13691);
nor U15851 (N_15851,N_12938,N_14671);
nand U15852 (N_15852,N_14599,N_13652);
xor U15853 (N_15853,N_14247,N_13425);
and U15854 (N_15854,N_13133,N_14553);
nor U15855 (N_15855,N_14467,N_12557);
nand U15856 (N_15856,N_14717,N_14458);
xor U15857 (N_15857,N_13350,N_14058);
nand U15858 (N_15858,N_14406,N_13336);
nor U15859 (N_15859,N_13655,N_13571);
nor U15860 (N_15860,N_13140,N_12721);
xnor U15861 (N_15861,N_12596,N_14578);
xnor U15862 (N_15862,N_13955,N_14195);
xnor U15863 (N_15863,N_14012,N_12958);
or U15864 (N_15864,N_13465,N_12525);
nor U15865 (N_15865,N_13959,N_13494);
nand U15866 (N_15866,N_14957,N_12863);
nand U15867 (N_15867,N_14378,N_12770);
nor U15868 (N_15868,N_13487,N_13258);
nor U15869 (N_15869,N_13825,N_13917);
xor U15870 (N_15870,N_13686,N_12741);
nor U15871 (N_15871,N_12852,N_13007);
and U15872 (N_15872,N_13707,N_13804);
nor U15873 (N_15873,N_13210,N_13696);
xnor U15874 (N_15874,N_14856,N_14137);
nand U15875 (N_15875,N_14419,N_13862);
nor U15876 (N_15876,N_12726,N_14285);
and U15877 (N_15877,N_13084,N_13861);
xnor U15878 (N_15878,N_12949,N_12537);
or U15879 (N_15879,N_12554,N_14844);
nand U15880 (N_15880,N_13637,N_14955);
nand U15881 (N_15881,N_13051,N_13239);
and U15882 (N_15882,N_14019,N_14688);
or U15883 (N_15883,N_13706,N_14051);
nand U15884 (N_15884,N_14952,N_13444);
xor U15885 (N_15885,N_13623,N_13230);
nor U15886 (N_15886,N_14757,N_14725);
or U15887 (N_15887,N_12693,N_14933);
nor U15888 (N_15888,N_13969,N_13179);
xor U15889 (N_15889,N_13782,N_14029);
or U15890 (N_15890,N_14146,N_13758);
and U15891 (N_15891,N_13582,N_13575);
and U15892 (N_15892,N_13061,N_14561);
nand U15893 (N_15893,N_14319,N_14277);
nand U15894 (N_15894,N_13883,N_13174);
xor U15895 (N_15895,N_13557,N_12744);
or U15896 (N_15896,N_14644,N_13826);
and U15897 (N_15897,N_14656,N_12776);
xor U15898 (N_15898,N_13234,N_14254);
xnor U15899 (N_15899,N_14121,N_14105);
nor U15900 (N_15900,N_14843,N_14548);
nand U15901 (N_15901,N_13601,N_12609);
and U15902 (N_15902,N_14069,N_13014);
or U15903 (N_15903,N_14057,N_14516);
nand U15904 (N_15904,N_13466,N_12669);
or U15905 (N_15905,N_14984,N_13407);
or U15906 (N_15906,N_13450,N_12578);
nand U15907 (N_15907,N_13040,N_14183);
xor U15908 (N_15908,N_13464,N_12793);
nor U15909 (N_15909,N_14849,N_14532);
xor U15910 (N_15910,N_12743,N_14002);
or U15911 (N_15911,N_13395,N_14756);
or U15912 (N_15912,N_14017,N_13031);
and U15913 (N_15913,N_13847,N_14264);
xor U15914 (N_15914,N_12504,N_13430);
xnor U15915 (N_15915,N_13509,N_14684);
and U15916 (N_15916,N_12671,N_13516);
and U15917 (N_15917,N_14030,N_13486);
nand U15918 (N_15918,N_13381,N_14291);
xnor U15919 (N_15919,N_14438,N_12701);
nor U15920 (N_15920,N_13744,N_14514);
xor U15921 (N_15921,N_13502,N_14305);
or U15922 (N_15922,N_13235,N_13753);
or U15923 (N_15923,N_12666,N_12853);
or U15924 (N_15924,N_13540,N_13867);
nand U15925 (N_15925,N_14948,N_14588);
or U15926 (N_15926,N_12926,N_12963);
nor U15927 (N_15927,N_12908,N_12756);
nor U15928 (N_15928,N_12530,N_13893);
xor U15929 (N_15929,N_12814,N_12869);
nand U15930 (N_15930,N_13323,N_13936);
nand U15931 (N_15931,N_12935,N_14608);
or U15932 (N_15932,N_14138,N_12532);
nand U15933 (N_15933,N_12628,N_14409);
nand U15934 (N_15934,N_13790,N_14685);
or U15935 (N_15935,N_12689,N_13980);
xnor U15936 (N_15936,N_14003,N_13886);
and U15937 (N_15937,N_12512,N_12847);
nand U15938 (N_15938,N_14794,N_13745);
xor U15939 (N_15939,N_13876,N_14680);
or U15940 (N_15940,N_14580,N_12983);
nor U15941 (N_15941,N_14233,N_14877);
or U15942 (N_15942,N_14275,N_14670);
and U15943 (N_15943,N_12664,N_14199);
nand U15944 (N_15944,N_14009,N_14819);
and U15945 (N_15945,N_13976,N_13968);
and U15946 (N_15946,N_13442,N_12535);
nor U15947 (N_15947,N_14479,N_14617);
nor U15948 (N_15948,N_14775,N_13414);
nor U15949 (N_15949,N_12645,N_13156);
xor U15950 (N_15950,N_14215,N_14365);
nand U15951 (N_15951,N_13153,N_12584);
and U15952 (N_15952,N_14276,N_13586);
xor U15953 (N_15953,N_14846,N_13496);
xnor U15954 (N_15954,N_13484,N_14699);
xor U15955 (N_15955,N_13016,N_13991);
xnor U15956 (N_15956,N_13971,N_13027);
nand U15957 (N_15957,N_14988,N_14257);
nand U15958 (N_15958,N_14450,N_14847);
and U15959 (N_15959,N_14871,N_12960);
and U15960 (N_15960,N_13208,N_13086);
nor U15961 (N_15961,N_14587,N_14417);
nand U15962 (N_15962,N_14628,N_14135);
and U15963 (N_15963,N_12898,N_12627);
or U15964 (N_15964,N_12838,N_13577);
nor U15965 (N_15965,N_13176,N_12916);
or U15966 (N_15966,N_12648,N_13389);
or U15967 (N_15967,N_13150,N_13513);
nor U15968 (N_15968,N_14555,N_14342);
or U15969 (N_15969,N_13115,N_14829);
or U15970 (N_15970,N_13451,N_14373);
nor U15971 (N_15971,N_12704,N_13699);
nand U15972 (N_15972,N_14096,N_13474);
nor U15973 (N_15973,N_13614,N_13269);
nand U15974 (N_15974,N_13353,N_14337);
nor U15975 (N_15975,N_14540,N_14889);
and U15976 (N_15976,N_13237,N_14840);
and U15977 (N_15977,N_13834,N_14439);
or U15978 (N_15978,N_13942,N_13238);
nand U15979 (N_15979,N_13214,N_14632);
or U15980 (N_15980,N_13047,N_13882);
and U15981 (N_15981,N_12981,N_12650);
and U15982 (N_15982,N_14172,N_14252);
xor U15983 (N_15983,N_12866,N_13996);
nor U15984 (N_15984,N_13264,N_12559);
nor U15985 (N_15985,N_13175,N_14873);
xor U15986 (N_15986,N_14652,N_14197);
nor U15987 (N_15987,N_13311,N_14272);
xnor U15988 (N_15988,N_14522,N_13771);
xor U15989 (N_15989,N_12802,N_13947);
nor U15990 (N_15990,N_14781,N_14965);
nand U15991 (N_15991,N_14586,N_13419);
nor U15992 (N_15992,N_14242,N_13957);
xor U15993 (N_15993,N_14614,N_14310);
xnor U15994 (N_15994,N_13249,N_14296);
nand U15995 (N_15995,N_14393,N_14572);
nor U15996 (N_15996,N_13438,N_14258);
nor U15997 (N_15997,N_13755,N_14159);
xor U15998 (N_15998,N_14049,N_13647);
nand U15999 (N_15999,N_12910,N_14706);
nor U16000 (N_16000,N_13566,N_13845);
and U16001 (N_16001,N_13189,N_13289);
or U16002 (N_16002,N_12716,N_13725);
nand U16003 (N_16003,N_14621,N_13312);
xor U16004 (N_16004,N_13709,N_13604);
and U16005 (N_16005,N_14903,N_13195);
nor U16006 (N_16006,N_14897,N_13973);
nand U16007 (N_16007,N_12694,N_13888);
or U16008 (N_16008,N_13072,N_13161);
nand U16009 (N_16009,N_14059,N_14833);
nor U16010 (N_16010,N_13294,N_14674);
and U16011 (N_16011,N_13470,N_13495);
nand U16012 (N_16012,N_13497,N_13747);
or U16013 (N_16013,N_13705,N_14036);
and U16014 (N_16014,N_12864,N_12912);
or U16015 (N_16015,N_13684,N_13944);
and U16016 (N_16016,N_12950,N_14803);
xnor U16017 (N_16017,N_13518,N_14092);
xor U16018 (N_16018,N_13600,N_14624);
nor U16019 (N_16019,N_13306,N_13157);
nor U16020 (N_16020,N_14619,N_14845);
xnor U16021 (N_16021,N_13286,N_13737);
nor U16022 (N_16022,N_13463,N_14683);
nor U16023 (N_16023,N_14400,N_13712);
nand U16024 (N_16024,N_14645,N_14169);
nand U16025 (N_16025,N_13553,N_12657);
and U16026 (N_16026,N_12937,N_12739);
xor U16027 (N_16027,N_14563,N_14330);
nand U16028 (N_16028,N_13298,N_13924);
nand U16029 (N_16029,N_12674,N_13075);
or U16030 (N_16030,N_14327,N_14566);
xnor U16031 (N_16031,N_13198,N_14512);
xnor U16032 (N_16032,N_13842,N_13774);
or U16033 (N_16033,N_12786,N_13352);
or U16034 (N_16034,N_14915,N_12582);
nor U16035 (N_16035,N_13136,N_12688);
nor U16036 (N_16036,N_13542,N_14401);
nor U16037 (N_16037,N_13910,N_14317);
xor U16038 (N_16038,N_13805,N_13673);
nor U16039 (N_16039,N_13792,N_12840);
or U16040 (N_16040,N_13648,N_14239);
nor U16041 (N_16041,N_13833,N_13107);
xor U16042 (N_16042,N_13343,N_13606);
xor U16043 (N_16043,N_13690,N_13854);
or U16044 (N_16044,N_14679,N_14177);
or U16045 (N_16045,N_14714,N_14484);
and U16046 (N_16046,N_12502,N_14287);
nor U16047 (N_16047,N_12975,N_14936);
nand U16048 (N_16048,N_14088,N_13173);
nor U16049 (N_16049,N_14862,N_14653);
xnor U16050 (N_16050,N_13916,N_14727);
nor U16051 (N_16051,N_12594,N_12812);
and U16052 (N_16052,N_14962,N_14414);
or U16053 (N_16053,N_12621,N_14326);
nand U16054 (N_16054,N_14144,N_14341);
nor U16055 (N_16055,N_14482,N_13056);
and U16056 (N_16056,N_14695,N_14250);
and U16057 (N_16057,N_12761,N_12517);
nor U16058 (N_16058,N_13382,N_13722);
or U16059 (N_16059,N_14527,N_14579);
and U16060 (N_16060,N_13094,N_12791);
xor U16061 (N_16061,N_14530,N_14867);
nor U16062 (N_16062,N_13562,N_13083);
xor U16063 (N_16063,N_13666,N_12799);
nor U16064 (N_16064,N_13455,N_14186);
or U16065 (N_16065,N_12695,N_14851);
xnor U16066 (N_16066,N_14356,N_14156);
nand U16067 (N_16067,N_14301,N_13998);
or U16068 (N_16068,N_12685,N_14132);
nor U16069 (N_16069,N_13281,N_13409);
xnor U16070 (N_16070,N_12668,N_12637);
nand U16071 (N_16071,N_13049,N_14130);
xnor U16072 (N_16072,N_14206,N_13152);
nor U16073 (N_16073,N_13412,N_13581);
nor U16074 (N_16074,N_13583,N_14413);
xor U16075 (N_16075,N_13167,N_14311);
nand U16076 (N_16076,N_14312,N_12763);
or U16077 (N_16077,N_12730,N_13120);
and U16078 (N_16078,N_12572,N_12783);
nand U16079 (N_16079,N_14117,N_12575);
and U16080 (N_16080,N_13227,N_14872);
nand U16081 (N_16081,N_14741,N_13556);
or U16082 (N_16082,N_14161,N_14449);
nor U16083 (N_16083,N_12515,N_14399);
xnor U16084 (N_16084,N_12890,N_13813);
nand U16085 (N_16085,N_12920,N_13521);
or U16086 (N_16086,N_14198,N_14943);
or U16087 (N_16087,N_14249,N_12529);
or U16088 (N_16088,N_12948,N_12888);
nand U16089 (N_16089,N_14203,N_14762);
and U16090 (N_16090,N_14407,N_14395);
nand U16091 (N_16091,N_13080,N_14986);
and U16092 (N_16092,N_13527,N_13555);
nor U16093 (N_16093,N_13221,N_14874);
or U16094 (N_16094,N_14127,N_13544);
xor U16095 (N_16095,N_13252,N_13743);
or U16096 (N_16096,N_14836,N_13332);
or U16097 (N_16097,N_14562,N_14060);
xor U16098 (N_16098,N_13534,N_13742);
nand U16099 (N_16099,N_13629,N_14643);
nor U16100 (N_16100,N_13377,N_12543);
nand U16101 (N_16101,N_14384,N_14212);
nor U16102 (N_16102,N_12779,N_12811);
and U16103 (N_16103,N_14284,N_14914);
xnor U16104 (N_16104,N_13868,N_14377);
nand U16105 (N_16105,N_13314,N_12639);
nor U16106 (N_16106,N_14649,N_14042);
nand U16107 (N_16107,N_13687,N_13296);
and U16108 (N_16108,N_14200,N_13913);
nor U16109 (N_16109,N_14571,N_14380);
nor U16110 (N_16110,N_13182,N_14094);
or U16111 (N_16111,N_12658,N_13482);
nor U16112 (N_16112,N_14793,N_13102);
and U16113 (N_16113,N_13741,N_14882);
or U16114 (N_16114,N_14895,N_13839);
or U16115 (N_16115,N_14434,N_13029);
xnor U16116 (N_16116,N_14961,N_13588);
nand U16117 (N_16117,N_12784,N_13108);
and U16118 (N_16118,N_13674,N_14442);
nand U16119 (N_16119,N_12909,N_13590);
or U16120 (N_16120,N_14364,N_14073);
or U16121 (N_16121,N_14520,N_12602);
or U16122 (N_16122,N_12604,N_13903);
or U16123 (N_16123,N_14297,N_14386);
xnor U16124 (N_16124,N_14126,N_12953);
nand U16125 (N_16125,N_13594,N_13579);
or U16126 (N_16126,N_14879,N_12702);
nor U16127 (N_16127,N_12919,N_14428);
xnor U16128 (N_16128,N_12848,N_13170);
and U16129 (N_16129,N_13185,N_12807);
and U16130 (N_16130,N_14953,N_14115);
or U16131 (N_16131,N_12737,N_14180);
nand U16132 (N_16132,N_14507,N_14712);
or U16133 (N_16133,N_13530,N_14369);
nor U16134 (N_16134,N_13780,N_14340);
xor U16135 (N_16135,N_13290,N_14293);
and U16136 (N_16136,N_13325,N_13852);
xor U16137 (N_16137,N_13358,N_14080);
or U16138 (N_16138,N_13204,N_14336);
and U16139 (N_16139,N_13714,N_13713);
xor U16140 (N_16140,N_12690,N_12605);
xnor U16141 (N_16141,N_13642,N_13307);
and U16142 (N_16142,N_12564,N_13654);
nand U16143 (N_16143,N_13320,N_14559);
nor U16144 (N_16144,N_14077,N_14550);
nor U16145 (N_16145,N_13697,N_13039);
or U16146 (N_16146,N_14107,N_14791);
xnor U16147 (N_16147,N_13090,N_12616);
xnor U16148 (N_16148,N_13457,N_14091);
xnor U16149 (N_16149,N_14716,N_14335);
and U16150 (N_16150,N_13892,N_12905);
or U16151 (N_16151,N_14329,N_13964);
nand U16152 (N_16152,N_13268,N_12957);
and U16153 (N_16153,N_12873,N_12797);
nand U16154 (N_16154,N_14476,N_14474);
and U16155 (N_16155,N_14190,N_13043);
or U16156 (N_16156,N_12861,N_13554);
nand U16157 (N_16157,N_14813,N_13493);
nand U16158 (N_16158,N_14065,N_13760);
and U16159 (N_16159,N_13946,N_13255);
and U16160 (N_16160,N_13784,N_13169);
nor U16161 (N_16161,N_14010,N_14320);
and U16162 (N_16162,N_12514,N_12538);
or U16163 (N_16163,N_13228,N_14306);
or U16164 (N_16164,N_13267,N_14743);
and U16165 (N_16165,N_12964,N_14466);
nor U16166 (N_16166,N_12562,N_14777);
nor U16167 (N_16167,N_14630,N_14900);
and U16168 (N_16168,N_13803,N_14736);
xnor U16169 (N_16169,N_12526,N_13719);
and U16170 (N_16170,N_14462,N_13754);
and U16171 (N_16171,N_14537,N_14544);
nand U16172 (N_16172,N_14501,N_12854);
or U16173 (N_16173,N_13399,N_13528);
nor U16174 (N_16174,N_14244,N_12555);
xor U16175 (N_16175,N_14018,N_13532);
and U16176 (N_16176,N_14831,N_13322);
and U16177 (N_16177,N_13875,N_13536);
nand U16178 (N_16178,N_13127,N_13262);
or U16179 (N_16179,N_13692,N_14412);
or U16180 (N_16180,N_13310,N_12867);
nand U16181 (N_16181,N_14543,N_13925);
nor U16182 (N_16182,N_12679,N_13718);
or U16183 (N_16183,N_13317,N_13178);
and U16184 (N_16184,N_13008,N_13459);
nor U16185 (N_16185,N_14976,N_13597);
nand U16186 (N_16186,N_13338,N_14124);
nand U16187 (N_16187,N_12836,N_12859);
nand U16188 (N_16188,N_12973,N_13664);
or U16189 (N_16189,N_14142,N_14677);
xor U16190 (N_16190,N_12930,N_13763);
xnor U16191 (N_16191,N_13303,N_14453);
or U16192 (N_16192,N_14302,N_14659);
or U16193 (N_16193,N_14455,N_13066);
and U16194 (N_16194,N_12870,N_14464);
and U16195 (N_16195,N_13324,N_14648);
nand U16196 (N_16196,N_14557,N_13280);
xor U16197 (N_16197,N_14768,N_14033);
xor U16198 (N_16198,N_14919,N_14338);
and U16199 (N_16199,N_13192,N_14945);
nand U16200 (N_16200,N_12552,N_14171);
xnor U16201 (N_16201,N_14167,N_13624);
nand U16202 (N_16202,N_14567,N_12798);
or U16203 (N_16203,N_13930,N_13855);
nand U16204 (N_16204,N_13559,N_13477);
nand U16205 (N_16205,N_13787,N_14838);
nor U16206 (N_16206,N_14489,N_14328);
nand U16207 (N_16207,N_13801,N_14920);
or U16208 (N_16208,N_13626,N_12914);
nor U16209 (N_16209,N_12513,N_13587);
xor U16210 (N_16210,N_13987,N_13359);
xor U16211 (N_16211,N_12571,N_14615);
nand U16212 (N_16212,N_13341,N_13769);
xnor U16213 (N_16213,N_14282,N_14270);
nand U16214 (N_16214,N_14766,N_13222);
nand U16215 (N_16215,N_13595,N_13809);
or U16216 (N_16216,N_12684,N_14278);
nand U16217 (N_16217,N_14740,N_13843);
nand U16218 (N_16218,N_12675,N_12652);
or U16219 (N_16219,N_14508,N_13437);
or U16220 (N_16220,N_12771,N_13878);
or U16221 (N_16221,N_13689,N_14410);
xor U16222 (N_16222,N_14517,N_14713);
nor U16223 (N_16223,N_13191,N_12868);
xnor U16224 (N_16224,N_13914,N_13363);
or U16225 (N_16225,N_14053,N_13525);
xor U16226 (N_16226,N_12886,N_14431);
nand U16227 (N_16227,N_13669,N_13788);
or U16228 (N_16228,N_13797,N_12720);
nand U16229 (N_16229,N_13333,N_14942);
and U16230 (N_16230,N_14357,N_14602);
or U16231 (N_16231,N_12977,N_12740);
xnor U16232 (N_16232,N_14496,N_13526);
xnor U16233 (N_16233,N_13740,N_13717);
or U16234 (N_16234,N_14202,N_14989);
or U16235 (N_16235,N_12553,N_14133);
and U16236 (N_16236,N_14866,N_13216);
xnor U16237 (N_16237,N_13631,N_14536);
xnor U16238 (N_16238,N_14191,N_13328);
and U16239 (N_16239,N_12523,N_13931);
nand U16240 (N_16240,N_14255,N_12748);
xor U16241 (N_16241,N_14720,N_12655);
nand U16242 (N_16242,N_13672,N_14744);
nand U16243 (N_16243,N_13770,N_12998);
or U16244 (N_16244,N_12943,N_14941);
xnor U16245 (N_16245,N_14731,N_14072);
nand U16246 (N_16246,N_13498,N_14174);
or U16247 (N_16247,N_13020,N_13529);
nor U16248 (N_16248,N_13138,N_13159);
nand U16249 (N_16249,N_13730,N_14822);
and U16250 (N_16250,N_14148,N_14881);
nand U16251 (N_16251,N_13839,N_13019);
nor U16252 (N_16252,N_14717,N_13502);
and U16253 (N_16253,N_12890,N_13479);
xor U16254 (N_16254,N_13714,N_14074);
nand U16255 (N_16255,N_13066,N_13107);
and U16256 (N_16256,N_14003,N_14648);
nand U16257 (N_16257,N_13467,N_12895);
nand U16258 (N_16258,N_12550,N_13977);
nand U16259 (N_16259,N_13310,N_14176);
nor U16260 (N_16260,N_13391,N_14254);
nor U16261 (N_16261,N_14886,N_14268);
nor U16262 (N_16262,N_13409,N_14184);
or U16263 (N_16263,N_14395,N_14910);
nand U16264 (N_16264,N_13152,N_13185);
or U16265 (N_16265,N_14726,N_12985);
nor U16266 (N_16266,N_13877,N_12754);
nand U16267 (N_16267,N_12705,N_14721);
nor U16268 (N_16268,N_14830,N_12596);
and U16269 (N_16269,N_14284,N_13947);
and U16270 (N_16270,N_13895,N_14994);
xnor U16271 (N_16271,N_13427,N_13299);
nand U16272 (N_16272,N_13179,N_13478);
nor U16273 (N_16273,N_13162,N_12859);
nand U16274 (N_16274,N_13509,N_14923);
nor U16275 (N_16275,N_13270,N_13628);
or U16276 (N_16276,N_13176,N_13556);
nand U16277 (N_16277,N_13216,N_14916);
nor U16278 (N_16278,N_13862,N_12988);
nor U16279 (N_16279,N_13658,N_13325);
xor U16280 (N_16280,N_12626,N_14015);
or U16281 (N_16281,N_13267,N_14662);
xor U16282 (N_16282,N_13542,N_13842);
and U16283 (N_16283,N_14133,N_14835);
nor U16284 (N_16284,N_14893,N_14250);
or U16285 (N_16285,N_14309,N_14291);
or U16286 (N_16286,N_13483,N_13024);
or U16287 (N_16287,N_12854,N_12673);
or U16288 (N_16288,N_13284,N_14043);
nor U16289 (N_16289,N_13209,N_13895);
and U16290 (N_16290,N_14967,N_12755);
nor U16291 (N_16291,N_13487,N_13315);
and U16292 (N_16292,N_14798,N_14468);
nor U16293 (N_16293,N_14330,N_13728);
and U16294 (N_16294,N_14734,N_13487);
xnor U16295 (N_16295,N_12796,N_14296);
nor U16296 (N_16296,N_12558,N_13049);
nand U16297 (N_16297,N_13603,N_13366);
xor U16298 (N_16298,N_14424,N_12571);
and U16299 (N_16299,N_14531,N_14222);
or U16300 (N_16300,N_13518,N_14050);
xnor U16301 (N_16301,N_13142,N_12602);
and U16302 (N_16302,N_12607,N_12675);
and U16303 (N_16303,N_12977,N_12868);
or U16304 (N_16304,N_14128,N_14001);
nand U16305 (N_16305,N_12861,N_13518);
and U16306 (N_16306,N_13719,N_14961);
xnor U16307 (N_16307,N_14824,N_13599);
or U16308 (N_16308,N_13282,N_14509);
or U16309 (N_16309,N_13924,N_13435);
or U16310 (N_16310,N_14531,N_12855);
nor U16311 (N_16311,N_13763,N_13622);
nand U16312 (N_16312,N_14608,N_14543);
and U16313 (N_16313,N_12545,N_14049);
nor U16314 (N_16314,N_14647,N_12966);
or U16315 (N_16315,N_13314,N_14601);
nand U16316 (N_16316,N_14297,N_14128);
xor U16317 (N_16317,N_12522,N_14616);
or U16318 (N_16318,N_13620,N_12795);
and U16319 (N_16319,N_13764,N_13753);
nor U16320 (N_16320,N_12714,N_13241);
and U16321 (N_16321,N_12648,N_14574);
or U16322 (N_16322,N_12990,N_13414);
and U16323 (N_16323,N_14280,N_13016);
and U16324 (N_16324,N_12773,N_12704);
xor U16325 (N_16325,N_14066,N_14204);
nand U16326 (N_16326,N_13445,N_14891);
and U16327 (N_16327,N_14723,N_13986);
nor U16328 (N_16328,N_13246,N_12799);
nor U16329 (N_16329,N_14039,N_14314);
xor U16330 (N_16330,N_14258,N_13454);
nor U16331 (N_16331,N_14774,N_12907);
xor U16332 (N_16332,N_14487,N_13782);
nand U16333 (N_16333,N_12729,N_14878);
or U16334 (N_16334,N_12894,N_12822);
nor U16335 (N_16335,N_13006,N_13621);
and U16336 (N_16336,N_13764,N_14510);
xor U16337 (N_16337,N_13265,N_14052);
nor U16338 (N_16338,N_13621,N_12679);
nor U16339 (N_16339,N_14441,N_14470);
and U16340 (N_16340,N_12581,N_14425);
nor U16341 (N_16341,N_14929,N_14461);
and U16342 (N_16342,N_13794,N_14230);
nand U16343 (N_16343,N_14499,N_13813);
nand U16344 (N_16344,N_14523,N_14917);
nand U16345 (N_16345,N_13047,N_13941);
nand U16346 (N_16346,N_13290,N_12879);
nor U16347 (N_16347,N_14251,N_13382);
xnor U16348 (N_16348,N_13466,N_13945);
and U16349 (N_16349,N_14417,N_13416);
nor U16350 (N_16350,N_12902,N_14205);
and U16351 (N_16351,N_13963,N_13384);
nor U16352 (N_16352,N_13800,N_13209);
nand U16353 (N_16353,N_13040,N_13192);
nand U16354 (N_16354,N_12878,N_12762);
and U16355 (N_16355,N_12994,N_13135);
and U16356 (N_16356,N_14295,N_13870);
or U16357 (N_16357,N_13627,N_14958);
and U16358 (N_16358,N_13892,N_13332);
nand U16359 (N_16359,N_12903,N_13023);
and U16360 (N_16360,N_13589,N_13692);
xor U16361 (N_16361,N_12938,N_12693);
nor U16362 (N_16362,N_13572,N_13442);
or U16363 (N_16363,N_13200,N_13737);
xor U16364 (N_16364,N_13093,N_12698);
and U16365 (N_16365,N_12915,N_14745);
or U16366 (N_16366,N_13738,N_13479);
xor U16367 (N_16367,N_14753,N_13897);
xnor U16368 (N_16368,N_14555,N_13023);
or U16369 (N_16369,N_14582,N_13272);
and U16370 (N_16370,N_13826,N_13410);
nand U16371 (N_16371,N_14421,N_14218);
nand U16372 (N_16372,N_12702,N_14666);
and U16373 (N_16373,N_14930,N_14301);
xor U16374 (N_16374,N_13381,N_12616);
and U16375 (N_16375,N_13729,N_12899);
nor U16376 (N_16376,N_14738,N_14405);
or U16377 (N_16377,N_13670,N_14531);
nor U16378 (N_16378,N_14900,N_14486);
or U16379 (N_16379,N_12780,N_12692);
nor U16380 (N_16380,N_13324,N_12550);
xnor U16381 (N_16381,N_12893,N_14951);
nor U16382 (N_16382,N_14082,N_14455);
and U16383 (N_16383,N_14385,N_14562);
xor U16384 (N_16384,N_13064,N_13001);
or U16385 (N_16385,N_14527,N_13339);
xnor U16386 (N_16386,N_13587,N_13212);
or U16387 (N_16387,N_14775,N_14670);
nor U16388 (N_16388,N_14528,N_13847);
and U16389 (N_16389,N_12582,N_13612);
nor U16390 (N_16390,N_12902,N_13833);
nor U16391 (N_16391,N_14751,N_14243);
and U16392 (N_16392,N_14475,N_13840);
nor U16393 (N_16393,N_14718,N_12996);
nor U16394 (N_16394,N_13080,N_12754);
xnor U16395 (N_16395,N_13734,N_14082);
and U16396 (N_16396,N_13608,N_12813);
nand U16397 (N_16397,N_12578,N_13361);
nand U16398 (N_16398,N_14075,N_13850);
or U16399 (N_16399,N_13658,N_14509);
nor U16400 (N_16400,N_13914,N_12862);
xor U16401 (N_16401,N_12674,N_13045);
xnor U16402 (N_16402,N_14101,N_12735);
nor U16403 (N_16403,N_14176,N_13353);
nand U16404 (N_16404,N_13188,N_13368);
nor U16405 (N_16405,N_14938,N_13831);
or U16406 (N_16406,N_13789,N_12806);
xnor U16407 (N_16407,N_13030,N_13187);
and U16408 (N_16408,N_12773,N_13058);
nor U16409 (N_16409,N_13239,N_13219);
and U16410 (N_16410,N_12909,N_13931);
nand U16411 (N_16411,N_14471,N_13682);
or U16412 (N_16412,N_13456,N_13204);
xor U16413 (N_16413,N_14542,N_13713);
and U16414 (N_16414,N_13859,N_13595);
nand U16415 (N_16415,N_14158,N_13328);
or U16416 (N_16416,N_14435,N_13715);
nand U16417 (N_16417,N_13138,N_12676);
and U16418 (N_16418,N_12644,N_13372);
nor U16419 (N_16419,N_12995,N_14038);
nand U16420 (N_16420,N_14953,N_13401);
xnor U16421 (N_16421,N_14119,N_12977);
nand U16422 (N_16422,N_13241,N_12775);
nor U16423 (N_16423,N_13199,N_13507);
nor U16424 (N_16424,N_13805,N_14948);
or U16425 (N_16425,N_13380,N_13255);
and U16426 (N_16426,N_14589,N_14739);
nand U16427 (N_16427,N_14350,N_12738);
xor U16428 (N_16428,N_14482,N_14006);
xor U16429 (N_16429,N_14616,N_12803);
xor U16430 (N_16430,N_14568,N_12892);
or U16431 (N_16431,N_12522,N_14195);
nand U16432 (N_16432,N_14882,N_14103);
xnor U16433 (N_16433,N_12568,N_12920);
and U16434 (N_16434,N_14510,N_12600);
or U16435 (N_16435,N_13393,N_13048);
xnor U16436 (N_16436,N_13548,N_12600);
nand U16437 (N_16437,N_14950,N_14093);
nand U16438 (N_16438,N_14929,N_14255);
xor U16439 (N_16439,N_13269,N_13426);
xnor U16440 (N_16440,N_12767,N_14630);
or U16441 (N_16441,N_14957,N_14409);
nand U16442 (N_16442,N_13937,N_13345);
xor U16443 (N_16443,N_12705,N_13617);
nand U16444 (N_16444,N_13990,N_13783);
and U16445 (N_16445,N_14990,N_12951);
nor U16446 (N_16446,N_13673,N_13058);
nor U16447 (N_16447,N_13486,N_12948);
and U16448 (N_16448,N_13270,N_14955);
or U16449 (N_16449,N_13774,N_14676);
nand U16450 (N_16450,N_14198,N_14157);
and U16451 (N_16451,N_12615,N_13872);
nand U16452 (N_16452,N_14456,N_14493);
nand U16453 (N_16453,N_14234,N_14779);
or U16454 (N_16454,N_12502,N_14773);
xor U16455 (N_16455,N_12685,N_13965);
xor U16456 (N_16456,N_12634,N_14567);
nand U16457 (N_16457,N_12982,N_13201);
or U16458 (N_16458,N_14453,N_13657);
nand U16459 (N_16459,N_13581,N_12503);
nand U16460 (N_16460,N_13073,N_14400);
nand U16461 (N_16461,N_14213,N_14236);
or U16462 (N_16462,N_12735,N_14510);
nand U16463 (N_16463,N_12665,N_13926);
nand U16464 (N_16464,N_13976,N_14956);
nand U16465 (N_16465,N_13371,N_14957);
or U16466 (N_16466,N_12791,N_14930);
nor U16467 (N_16467,N_14887,N_14093);
nor U16468 (N_16468,N_13824,N_12688);
nor U16469 (N_16469,N_13076,N_13837);
xor U16470 (N_16470,N_14696,N_13248);
or U16471 (N_16471,N_13752,N_13352);
and U16472 (N_16472,N_13282,N_13722);
nand U16473 (N_16473,N_14151,N_12806);
xor U16474 (N_16474,N_13009,N_13075);
or U16475 (N_16475,N_14887,N_13556);
nand U16476 (N_16476,N_14591,N_14140);
xnor U16477 (N_16477,N_12848,N_14902);
nor U16478 (N_16478,N_14354,N_13338);
or U16479 (N_16479,N_14815,N_14703);
nor U16480 (N_16480,N_13080,N_14409);
or U16481 (N_16481,N_14127,N_13806);
nand U16482 (N_16482,N_13795,N_14579);
nor U16483 (N_16483,N_13279,N_12573);
and U16484 (N_16484,N_14042,N_13961);
nor U16485 (N_16485,N_14929,N_14766);
xnor U16486 (N_16486,N_13978,N_14110);
and U16487 (N_16487,N_14360,N_12971);
and U16488 (N_16488,N_14537,N_12587);
xnor U16489 (N_16489,N_13844,N_13936);
and U16490 (N_16490,N_14869,N_12588);
or U16491 (N_16491,N_13298,N_12559);
nand U16492 (N_16492,N_13331,N_13089);
nor U16493 (N_16493,N_13969,N_14624);
nor U16494 (N_16494,N_13076,N_14889);
or U16495 (N_16495,N_13273,N_12835);
and U16496 (N_16496,N_14947,N_14328);
and U16497 (N_16497,N_14574,N_14490);
xor U16498 (N_16498,N_13590,N_14959);
nand U16499 (N_16499,N_13598,N_13641);
nor U16500 (N_16500,N_13433,N_13724);
nand U16501 (N_16501,N_14507,N_13965);
xnor U16502 (N_16502,N_13893,N_14397);
or U16503 (N_16503,N_14098,N_13880);
nor U16504 (N_16504,N_13964,N_14655);
or U16505 (N_16505,N_13976,N_13796);
xnor U16506 (N_16506,N_14183,N_13894);
xor U16507 (N_16507,N_13745,N_12866);
xnor U16508 (N_16508,N_14322,N_14483);
or U16509 (N_16509,N_14784,N_14486);
nand U16510 (N_16510,N_13355,N_14514);
and U16511 (N_16511,N_12537,N_12807);
nand U16512 (N_16512,N_14918,N_14368);
nand U16513 (N_16513,N_12779,N_14025);
and U16514 (N_16514,N_14070,N_13156);
nor U16515 (N_16515,N_14338,N_14376);
nand U16516 (N_16516,N_12822,N_13187);
xor U16517 (N_16517,N_14239,N_13755);
xnor U16518 (N_16518,N_13598,N_13682);
or U16519 (N_16519,N_12610,N_14507);
nand U16520 (N_16520,N_14459,N_14385);
nor U16521 (N_16521,N_13781,N_14979);
xor U16522 (N_16522,N_13040,N_12977);
xor U16523 (N_16523,N_13785,N_12870);
or U16524 (N_16524,N_13760,N_13822);
or U16525 (N_16525,N_13060,N_14122);
or U16526 (N_16526,N_14241,N_14370);
nor U16527 (N_16527,N_13023,N_13074);
or U16528 (N_16528,N_13246,N_14805);
and U16529 (N_16529,N_14187,N_14240);
nand U16530 (N_16530,N_13528,N_12979);
nand U16531 (N_16531,N_12774,N_13612);
or U16532 (N_16532,N_14363,N_12995);
or U16533 (N_16533,N_12802,N_13141);
nor U16534 (N_16534,N_14512,N_12501);
xnor U16535 (N_16535,N_13673,N_14239);
xor U16536 (N_16536,N_12876,N_13369);
and U16537 (N_16537,N_13241,N_13905);
nor U16538 (N_16538,N_13052,N_12641);
nor U16539 (N_16539,N_13668,N_12876);
nor U16540 (N_16540,N_14246,N_12788);
or U16541 (N_16541,N_12642,N_13166);
xnor U16542 (N_16542,N_13633,N_14967);
and U16543 (N_16543,N_13702,N_13871);
nor U16544 (N_16544,N_13703,N_14417);
or U16545 (N_16545,N_14234,N_14414);
or U16546 (N_16546,N_14050,N_13852);
nand U16547 (N_16547,N_13558,N_13583);
and U16548 (N_16548,N_12928,N_12678);
nand U16549 (N_16549,N_13401,N_13566);
xor U16550 (N_16550,N_12703,N_12601);
nand U16551 (N_16551,N_14473,N_14858);
nor U16552 (N_16552,N_14112,N_13553);
xnor U16553 (N_16553,N_13367,N_14721);
or U16554 (N_16554,N_13666,N_12588);
xnor U16555 (N_16555,N_13879,N_13494);
or U16556 (N_16556,N_13553,N_12987);
xnor U16557 (N_16557,N_14666,N_13171);
xor U16558 (N_16558,N_13662,N_14799);
or U16559 (N_16559,N_14336,N_14356);
nor U16560 (N_16560,N_14759,N_14869);
or U16561 (N_16561,N_13132,N_14802);
xor U16562 (N_16562,N_12988,N_13696);
nor U16563 (N_16563,N_13414,N_14052);
nand U16564 (N_16564,N_14595,N_14886);
nor U16565 (N_16565,N_14123,N_12583);
nand U16566 (N_16566,N_14901,N_14215);
xor U16567 (N_16567,N_13871,N_13721);
and U16568 (N_16568,N_14394,N_13606);
nand U16569 (N_16569,N_12816,N_13290);
and U16570 (N_16570,N_14266,N_14503);
nor U16571 (N_16571,N_13094,N_13939);
xor U16572 (N_16572,N_13066,N_14418);
nand U16573 (N_16573,N_13666,N_14393);
or U16574 (N_16574,N_12844,N_13386);
xnor U16575 (N_16575,N_12888,N_14896);
nor U16576 (N_16576,N_13557,N_14756);
and U16577 (N_16577,N_12924,N_14188);
and U16578 (N_16578,N_14670,N_14546);
or U16579 (N_16579,N_13291,N_13478);
or U16580 (N_16580,N_13136,N_12564);
nor U16581 (N_16581,N_13608,N_14174);
nor U16582 (N_16582,N_14713,N_12960);
or U16583 (N_16583,N_13857,N_14241);
or U16584 (N_16584,N_14262,N_14139);
or U16585 (N_16585,N_13194,N_13701);
nand U16586 (N_16586,N_14586,N_14366);
and U16587 (N_16587,N_14866,N_14054);
nand U16588 (N_16588,N_14444,N_14685);
nand U16589 (N_16589,N_14420,N_14216);
nand U16590 (N_16590,N_12672,N_13054);
nor U16591 (N_16591,N_13545,N_14944);
xnor U16592 (N_16592,N_14848,N_13440);
nor U16593 (N_16593,N_12715,N_14478);
nor U16594 (N_16594,N_14906,N_14206);
or U16595 (N_16595,N_14439,N_13485);
nand U16596 (N_16596,N_14274,N_14598);
nor U16597 (N_16597,N_14771,N_13645);
nor U16598 (N_16598,N_13361,N_12793);
and U16599 (N_16599,N_14143,N_13256);
nand U16600 (N_16600,N_14480,N_13172);
or U16601 (N_16601,N_12657,N_13573);
or U16602 (N_16602,N_14742,N_13651);
nand U16603 (N_16603,N_14783,N_13345);
xor U16604 (N_16604,N_14193,N_13798);
nand U16605 (N_16605,N_12521,N_12806);
xnor U16606 (N_16606,N_13711,N_14080);
nand U16607 (N_16607,N_14378,N_12999);
xnor U16608 (N_16608,N_14773,N_14303);
nand U16609 (N_16609,N_13678,N_12904);
nor U16610 (N_16610,N_12676,N_13839);
nor U16611 (N_16611,N_12730,N_13309);
and U16612 (N_16612,N_14248,N_14266);
or U16613 (N_16613,N_12713,N_14361);
or U16614 (N_16614,N_13832,N_14753);
or U16615 (N_16615,N_12997,N_12803);
nor U16616 (N_16616,N_14628,N_13717);
xor U16617 (N_16617,N_12939,N_14350);
xor U16618 (N_16618,N_12679,N_12509);
and U16619 (N_16619,N_13599,N_13159);
or U16620 (N_16620,N_14002,N_13069);
xor U16621 (N_16621,N_13854,N_12615);
and U16622 (N_16622,N_13029,N_13452);
and U16623 (N_16623,N_12647,N_14554);
nand U16624 (N_16624,N_13201,N_14553);
nor U16625 (N_16625,N_13164,N_14880);
nor U16626 (N_16626,N_14217,N_13654);
xnor U16627 (N_16627,N_12808,N_14360);
and U16628 (N_16628,N_12970,N_13845);
and U16629 (N_16629,N_13668,N_13486);
nor U16630 (N_16630,N_13535,N_14282);
or U16631 (N_16631,N_14479,N_14543);
or U16632 (N_16632,N_14683,N_14279);
nand U16633 (N_16633,N_14354,N_13884);
and U16634 (N_16634,N_14279,N_14074);
nor U16635 (N_16635,N_12869,N_13155);
nand U16636 (N_16636,N_13469,N_14835);
and U16637 (N_16637,N_14701,N_13240);
nand U16638 (N_16638,N_14190,N_14617);
or U16639 (N_16639,N_13900,N_12916);
nor U16640 (N_16640,N_13023,N_12632);
or U16641 (N_16641,N_14838,N_13754);
nor U16642 (N_16642,N_14717,N_12991);
nand U16643 (N_16643,N_13065,N_12636);
or U16644 (N_16644,N_12564,N_14282);
or U16645 (N_16645,N_14833,N_13228);
nand U16646 (N_16646,N_14070,N_13496);
nand U16647 (N_16647,N_12872,N_13565);
xnor U16648 (N_16648,N_14192,N_13932);
and U16649 (N_16649,N_13952,N_13712);
xor U16650 (N_16650,N_14608,N_13122);
xor U16651 (N_16651,N_14951,N_13909);
or U16652 (N_16652,N_14405,N_14236);
xnor U16653 (N_16653,N_13191,N_14527);
or U16654 (N_16654,N_13367,N_14118);
nand U16655 (N_16655,N_13185,N_13135);
nor U16656 (N_16656,N_14076,N_13079);
xnor U16657 (N_16657,N_13238,N_13499);
xor U16658 (N_16658,N_14528,N_13885);
nor U16659 (N_16659,N_14667,N_13248);
or U16660 (N_16660,N_12666,N_13980);
or U16661 (N_16661,N_13036,N_14961);
or U16662 (N_16662,N_13086,N_12953);
nand U16663 (N_16663,N_14623,N_13993);
nand U16664 (N_16664,N_13278,N_12924);
and U16665 (N_16665,N_12920,N_14264);
xor U16666 (N_16666,N_14086,N_12862);
nand U16667 (N_16667,N_12686,N_13639);
nor U16668 (N_16668,N_14668,N_12502);
nand U16669 (N_16669,N_13801,N_13057);
xnor U16670 (N_16670,N_12777,N_13928);
nand U16671 (N_16671,N_13986,N_13296);
xor U16672 (N_16672,N_14856,N_14226);
or U16673 (N_16673,N_13561,N_14251);
nand U16674 (N_16674,N_13226,N_13702);
nor U16675 (N_16675,N_13782,N_14445);
xnor U16676 (N_16676,N_13355,N_12690);
nor U16677 (N_16677,N_14021,N_12906);
nor U16678 (N_16678,N_13429,N_12764);
nor U16679 (N_16679,N_12954,N_14592);
and U16680 (N_16680,N_12676,N_13394);
nor U16681 (N_16681,N_13975,N_13842);
nor U16682 (N_16682,N_13776,N_13074);
nor U16683 (N_16683,N_14010,N_12878);
nand U16684 (N_16684,N_14903,N_12786);
xor U16685 (N_16685,N_14433,N_14553);
nand U16686 (N_16686,N_13573,N_12567);
and U16687 (N_16687,N_14593,N_14926);
nor U16688 (N_16688,N_12563,N_14378);
or U16689 (N_16689,N_13196,N_13017);
nor U16690 (N_16690,N_13040,N_13371);
nand U16691 (N_16691,N_14358,N_13994);
or U16692 (N_16692,N_13183,N_12536);
nand U16693 (N_16693,N_12858,N_13874);
or U16694 (N_16694,N_14215,N_13468);
or U16695 (N_16695,N_13968,N_14171);
xnor U16696 (N_16696,N_12512,N_14783);
xnor U16697 (N_16697,N_12644,N_13250);
xor U16698 (N_16698,N_14047,N_12803);
xnor U16699 (N_16699,N_14869,N_13483);
nand U16700 (N_16700,N_13875,N_14696);
or U16701 (N_16701,N_13923,N_13631);
xnor U16702 (N_16702,N_12657,N_13857);
nand U16703 (N_16703,N_13613,N_13097);
and U16704 (N_16704,N_12991,N_12671);
nand U16705 (N_16705,N_13890,N_12537);
xnor U16706 (N_16706,N_13843,N_12768);
xor U16707 (N_16707,N_12658,N_14862);
nor U16708 (N_16708,N_14523,N_13918);
nand U16709 (N_16709,N_12723,N_13506);
or U16710 (N_16710,N_12791,N_13089);
xor U16711 (N_16711,N_14746,N_14976);
or U16712 (N_16712,N_12543,N_14531);
nor U16713 (N_16713,N_13279,N_12539);
xor U16714 (N_16714,N_14859,N_14163);
xor U16715 (N_16715,N_13236,N_12547);
and U16716 (N_16716,N_14194,N_13483);
xnor U16717 (N_16717,N_14847,N_14620);
xnor U16718 (N_16718,N_14797,N_14331);
or U16719 (N_16719,N_14120,N_14473);
and U16720 (N_16720,N_12802,N_12761);
and U16721 (N_16721,N_14515,N_13894);
xnor U16722 (N_16722,N_13444,N_14940);
nor U16723 (N_16723,N_14805,N_12589);
xor U16724 (N_16724,N_13510,N_13095);
or U16725 (N_16725,N_13805,N_14544);
and U16726 (N_16726,N_13583,N_12587);
or U16727 (N_16727,N_13686,N_14744);
or U16728 (N_16728,N_13570,N_14657);
nand U16729 (N_16729,N_14771,N_14787);
nand U16730 (N_16730,N_14039,N_14658);
or U16731 (N_16731,N_13792,N_13454);
nand U16732 (N_16732,N_14139,N_12969);
or U16733 (N_16733,N_13456,N_13661);
nand U16734 (N_16734,N_12689,N_13983);
nand U16735 (N_16735,N_14496,N_13737);
nor U16736 (N_16736,N_13329,N_12568);
or U16737 (N_16737,N_14242,N_13679);
or U16738 (N_16738,N_13383,N_14118);
and U16739 (N_16739,N_14052,N_14391);
nand U16740 (N_16740,N_14565,N_13440);
nor U16741 (N_16741,N_14951,N_13082);
and U16742 (N_16742,N_13966,N_13367);
or U16743 (N_16743,N_14666,N_14194);
or U16744 (N_16744,N_12558,N_14157);
xnor U16745 (N_16745,N_12797,N_12940);
or U16746 (N_16746,N_13887,N_14452);
nand U16747 (N_16747,N_13372,N_14737);
or U16748 (N_16748,N_14422,N_13830);
nor U16749 (N_16749,N_13181,N_13551);
xor U16750 (N_16750,N_12775,N_13044);
xnor U16751 (N_16751,N_14096,N_13032);
or U16752 (N_16752,N_14657,N_12857);
nand U16753 (N_16753,N_14219,N_13681);
xor U16754 (N_16754,N_12720,N_14378);
nor U16755 (N_16755,N_13328,N_13037);
or U16756 (N_16756,N_13216,N_13681);
xnor U16757 (N_16757,N_14798,N_14485);
or U16758 (N_16758,N_12883,N_14869);
and U16759 (N_16759,N_14417,N_14007);
nand U16760 (N_16760,N_13942,N_13388);
xnor U16761 (N_16761,N_14908,N_13173);
xor U16762 (N_16762,N_13044,N_14344);
or U16763 (N_16763,N_13957,N_14817);
or U16764 (N_16764,N_13002,N_14250);
nand U16765 (N_16765,N_14721,N_12505);
xor U16766 (N_16766,N_12839,N_13038);
nand U16767 (N_16767,N_13385,N_12801);
and U16768 (N_16768,N_12566,N_12889);
nand U16769 (N_16769,N_14740,N_13810);
nor U16770 (N_16770,N_12779,N_13897);
nand U16771 (N_16771,N_13538,N_14877);
xnor U16772 (N_16772,N_12631,N_14104);
nand U16773 (N_16773,N_14159,N_13667);
nor U16774 (N_16774,N_13014,N_12949);
or U16775 (N_16775,N_14957,N_14160);
nand U16776 (N_16776,N_14650,N_13826);
nor U16777 (N_16777,N_13890,N_14601);
or U16778 (N_16778,N_13195,N_12514);
or U16779 (N_16779,N_13856,N_13432);
nor U16780 (N_16780,N_12811,N_14901);
nand U16781 (N_16781,N_13711,N_13010);
xor U16782 (N_16782,N_14928,N_14321);
xor U16783 (N_16783,N_13441,N_13805);
and U16784 (N_16784,N_13833,N_13713);
xnor U16785 (N_16785,N_13725,N_14472);
nand U16786 (N_16786,N_12530,N_13825);
nor U16787 (N_16787,N_14728,N_13040);
and U16788 (N_16788,N_13850,N_13205);
nand U16789 (N_16789,N_13148,N_14370);
xnor U16790 (N_16790,N_13274,N_12776);
or U16791 (N_16791,N_14948,N_13963);
nor U16792 (N_16792,N_14939,N_14400);
nand U16793 (N_16793,N_12995,N_12815);
nand U16794 (N_16794,N_12673,N_14771);
or U16795 (N_16795,N_14579,N_13057);
or U16796 (N_16796,N_14655,N_14895);
xnor U16797 (N_16797,N_13469,N_14073);
or U16798 (N_16798,N_14915,N_14821);
or U16799 (N_16799,N_13841,N_14969);
nand U16800 (N_16800,N_14919,N_14385);
xnor U16801 (N_16801,N_13459,N_12931);
xnor U16802 (N_16802,N_13616,N_14062);
xnor U16803 (N_16803,N_14229,N_12678);
or U16804 (N_16804,N_14202,N_13090);
nor U16805 (N_16805,N_14434,N_13307);
nand U16806 (N_16806,N_14501,N_13067);
or U16807 (N_16807,N_13178,N_13818);
nand U16808 (N_16808,N_14400,N_12529);
or U16809 (N_16809,N_14427,N_13317);
and U16810 (N_16810,N_14537,N_12740);
nand U16811 (N_16811,N_12773,N_14281);
nand U16812 (N_16812,N_14520,N_12926);
nand U16813 (N_16813,N_13082,N_13974);
nor U16814 (N_16814,N_14153,N_13884);
nand U16815 (N_16815,N_14801,N_13775);
xnor U16816 (N_16816,N_13992,N_13734);
nand U16817 (N_16817,N_14439,N_14360);
nor U16818 (N_16818,N_12890,N_13908);
xor U16819 (N_16819,N_13674,N_13901);
xnor U16820 (N_16820,N_13446,N_13822);
and U16821 (N_16821,N_14331,N_13813);
or U16822 (N_16822,N_12658,N_13900);
xnor U16823 (N_16823,N_13449,N_12748);
nor U16824 (N_16824,N_14168,N_14335);
nand U16825 (N_16825,N_13679,N_14297);
nor U16826 (N_16826,N_14683,N_13737);
nand U16827 (N_16827,N_12520,N_13601);
or U16828 (N_16828,N_13028,N_12880);
and U16829 (N_16829,N_13778,N_12942);
xor U16830 (N_16830,N_13436,N_14112);
and U16831 (N_16831,N_14372,N_12782);
nand U16832 (N_16832,N_14957,N_13506);
nand U16833 (N_16833,N_13601,N_13002);
or U16834 (N_16834,N_13931,N_13572);
and U16835 (N_16835,N_13166,N_14529);
or U16836 (N_16836,N_13279,N_12596);
nand U16837 (N_16837,N_13488,N_14926);
and U16838 (N_16838,N_14913,N_13456);
or U16839 (N_16839,N_14313,N_14952);
nand U16840 (N_16840,N_14253,N_14360);
and U16841 (N_16841,N_14493,N_12503);
or U16842 (N_16842,N_14675,N_13883);
nand U16843 (N_16843,N_13513,N_13531);
nor U16844 (N_16844,N_13929,N_13043);
nand U16845 (N_16845,N_14348,N_13710);
and U16846 (N_16846,N_14391,N_13363);
and U16847 (N_16847,N_13671,N_12562);
and U16848 (N_16848,N_12942,N_14530);
nand U16849 (N_16849,N_12717,N_13104);
xor U16850 (N_16850,N_14077,N_12737);
nor U16851 (N_16851,N_14084,N_13526);
or U16852 (N_16852,N_12611,N_14359);
nand U16853 (N_16853,N_13447,N_13390);
nand U16854 (N_16854,N_14745,N_12980);
and U16855 (N_16855,N_12678,N_13360);
and U16856 (N_16856,N_14825,N_14553);
or U16857 (N_16857,N_12810,N_13023);
and U16858 (N_16858,N_13549,N_14693);
nor U16859 (N_16859,N_12687,N_12832);
nor U16860 (N_16860,N_13859,N_13060);
or U16861 (N_16861,N_14596,N_12728);
or U16862 (N_16862,N_13816,N_12609);
nand U16863 (N_16863,N_13766,N_14258);
xnor U16864 (N_16864,N_12812,N_13552);
nand U16865 (N_16865,N_13131,N_13927);
and U16866 (N_16866,N_13649,N_14898);
nand U16867 (N_16867,N_14445,N_12517);
or U16868 (N_16868,N_12947,N_13254);
nor U16869 (N_16869,N_14887,N_13071);
nor U16870 (N_16870,N_14688,N_12899);
and U16871 (N_16871,N_13187,N_13461);
xor U16872 (N_16872,N_12972,N_14878);
xnor U16873 (N_16873,N_14678,N_14213);
xor U16874 (N_16874,N_14051,N_14551);
nor U16875 (N_16875,N_12862,N_13009);
nor U16876 (N_16876,N_13456,N_13741);
nor U16877 (N_16877,N_14081,N_13551);
and U16878 (N_16878,N_13674,N_13639);
and U16879 (N_16879,N_14822,N_12685);
xnor U16880 (N_16880,N_13984,N_13454);
nand U16881 (N_16881,N_13967,N_14916);
nand U16882 (N_16882,N_14289,N_13189);
or U16883 (N_16883,N_14269,N_13439);
nand U16884 (N_16884,N_13853,N_14487);
and U16885 (N_16885,N_13616,N_14522);
or U16886 (N_16886,N_14564,N_12809);
nor U16887 (N_16887,N_13737,N_13900);
nor U16888 (N_16888,N_13164,N_13169);
xnor U16889 (N_16889,N_13651,N_12846);
and U16890 (N_16890,N_14264,N_13355);
nand U16891 (N_16891,N_12976,N_14411);
or U16892 (N_16892,N_12611,N_13182);
and U16893 (N_16893,N_12969,N_13514);
or U16894 (N_16894,N_14438,N_12949);
nor U16895 (N_16895,N_13308,N_14859);
and U16896 (N_16896,N_13713,N_14427);
xor U16897 (N_16897,N_12938,N_14897);
and U16898 (N_16898,N_13659,N_13722);
nor U16899 (N_16899,N_13125,N_14516);
or U16900 (N_16900,N_14199,N_13711);
nor U16901 (N_16901,N_13629,N_14415);
xnor U16902 (N_16902,N_14390,N_14681);
and U16903 (N_16903,N_14715,N_13761);
and U16904 (N_16904,N_14060,N_14936);
nand U16905 (N_16905,N_14228,N_14734);
nor U16906 (N_16906,N_14973,N_12882);
or U16907 (N_16907,N_14424,N_14502);
or U16908 (N_16908,N_12935,N_14997);
nor U16909 (N_16909,N_14667,N_12616);
or U16910 (N_16910,N_12734,N_13070);
nand U16911 (N_16911,N_13029,N_13638);
nand U16912 (N_16912,N_13486,N_14532);
and U16913 (N_16913,N_12706,N_14663);
nand U16914 (N_16914,N_12782,N_14944);
nor U16915 (N_16915,N_14296,N_13252);
or U16916 (N_16916,N_12598,N_13325);
or U16917 (N_16917,N_14495,N_13186);
nor U16918 (N_16918,N_12930,N_13490);
nand U16919 (N_16919,N_14311,N_13376);
and U16920 (N_16920,N_13343,N_14270);
and U16921 (N_16921,N_12946,N_14009);
nand U16922 (N_16922,N_14122,N_12669);
and U16923 (N_16923,N_13549,N_13852);
and U16924 (N_16924,N_14590,N_14818);
xor U16925 (N_16925,N_12699,N_13178);
xor U16926 (N_16926,N_14242,N_13605);
nand U16927 (N_16927,N_13094,N_14802);
or U16928 (N_16928,N_14624,N_12670);
nand U16929 (N_16929,N_13038,N_14311);
and U16930 (N_16930,N_14750,N_13998);
and U16931 (N_16931,N_13903,N_12921);
xor U16932 (N_16932,N_14632,N_12551);
or U16933 (N_16933,N_13384,N_12914);
nand U16934 (N_16934,N_13486,N_12696);
nand U16935 (N_16935,N_14210,N_14692);
xnor U16936 (N_16936,N_13554,N_13893);
xor U16937 (N_16937,N_14480,N_12797);
nand U16938 (N_16938,N_14918,N_13228);
nor U16939 (N_16939,N_14603,N_13758);
nor U16940 (N_16940,N_13512,N_14076);
xnor U16941 (N_16941,N_14364,N_12828);
xor U16942 (N_16942,N_14499,N_13911);
or U16943 (N_16943,N_13619,N_12551);
or U16944 (N_16944,N_13090,N_14895);
xor U16945 (N_16945,N_14489,N_13326);
nand U16946 (N_16946,N_13822,N_13664);
and U16947 (N_16947,N_14613,N_13199);
or U16948 (N_16948,N_12921,N_13941);
or U16949 (N_16949,N_13470,N_14603);
nand U16950 (N_16950,N_14392,N_12771);
xnor U16951 (N_16951,N_14719,N_12835);
xor U16952 (N_16952,N_13214,N_14085);
or U16953 (N_16953,N_13158,N_14281);
xnor U16954 (N_16954,N_13033,N_12960);
xor U16955 (N_16955,N_13417,N_14293);
nor U16956 (N_16956,N_13702,N_12621);
or U16957 (N_16957,N_14240,N_12795);
nor U16958 (N_16958,N_13985,N_14728);
and U16959 (N_16959,N_13713,N_14580);
nor U16960 (N_16960,N_14876,N_13076);
or U16961 (N_16961,N_13190,N_14389);
nor U16962 (N_16962,N_14936,N_14393);
xor U16963 (N_16963,N_14665,N_13708);
xor U16964 (N_16964,N_14206,N_13566);
nand U16965 (N_16965,N_12662,N_13992);
nor U16966 (N_16966,N_14344,N_13726);
nor U16967 (N_16967,N_14581,N_14128);
nand U16968 (N_16968,N_14235,N_13879);
xor U16969 (N_16969,N_13925,N_13142);
xnor U16970 (N_16970,N_12626,N_12508);
or U16971 (N_16971,N_14244,N_14111);
nand U16972 (N_16972,N_13195,N_13038);
and U16973 (N_16973,N_12514,N_14390);
or U16974 (N_16974,N_13018,N_14113);
and U16975 (N_16975,N_14312,N_12976);
nor U16976 (N_16976,N_12645,N_14503);
or U16977 (N_16977,N_12885,N_13304);
or U16978 (N_16978,N_12727,N_12696);
nand U16979 (N_16979,N_13202,N_14545);
nor U16980 (N_16980,N_14113,N_13563);
nand U16981 (N_16981,N_12916,N_13273);
xor U16982 (N_16982,N_14414,N_14289);
nor U16983 (N_16983,N_13177,N_14813);
nand U16984 (N_16984,N_14724,N_14917);
or U16985 (N_16985,N_12983,N_13186);
nand U16986 (N_16986,N_13586,N_13697);
and U16987 (N_16987,N_12937,N_14936);
or U16988 (N_16988,N_13544,N_12527);
nor U16989 (N_16989,N_13732,N_13619);
and U16990 (N_16990,N_12626,N_12591);
xnor U16991 (N_16991,N_13100,N_13140);
or U16992 (N_16992,N_12759,N_13089);
and U16993 (N_16993,N_13311,N_14064);
or U16994 (N_16994,N_13814,N_14607);
xnor U16995 (N_16995,N_14664,N_14320);
nand U16996 (N_16996,N_12804,N_14963);
or U16997 (N_16997,N_14104,N_14362);
or U16998 (N_16998,N_13253,N_13660);
nand U16999 (N_16999,N_13205,N_14742);
or U17000 (N_17000,N_13606,N_14464);
nand U17001 (N_17001,N_13557,N_14133);
and U17002 (N_17002,N_13758,N_14929);
nor U17003 (N_17003,N_13417,N_12808);
nor U17004 (N_17004,N_12717,N_12716);
nand U17005 (N_17005,N_14516,N_14088);
nand U17006 (N_17006,N_12637,N_12916);
and U17007 (N_17007,N_13094,N_14490);
nor U17008 (N_17008,N_13357,N_13374);
or U17009 (N_17009,N_13066,N_12595);
and U17010 (N_17010,N_13188,N_13377);
nand U17011 (N_17011,N_14816,N_13696);
and U17012 (N_17012,N_14140,N_13715);
xnor U17013 (N_17013,N_14444,N_13071);
or U17014 (N_17014,N_12788,N_12797);
or U17015 (N_17015,N_13564,N_14157);
nand U17016 (N_17016,N_12594,N_14053);
xor U17017 (N_17017,N_14131,N_12514);
xnor U17018 (N_17018,N_12933,N_13019);
or U17019 (N_17019,N_14260,N_13613);
nand U17020 (N_17020,N_14870,N_13143);
nor U17021 (N_17021,N_14714,N_14200);
nand U17022 (N_17022,N_14901,N_12621);
xor U17023 (N_17023,N_14195,N_13076);
nor U17024 (N_17024,N_13268,N_13190);
xor U17025 (N_17025,N_13551,N_13977);
nand U17026 (N_17026,N_13429,N_13206);
nor U17027 (N_17027,N_12927,N_14991);
or U17028 (N_17028,N_14480,N_13063);
nor U17029 (N_17029,N_13528,N_13617);
xor U17030 (N_17030,N_12906,N_13059);
nor U17031 (N_17031,N_12753,N_13744);
or U17032 (N_17032,N_14225,N_14850);
and U17033 (N_17033,N_12814,N_13212);
or U17034 (N_17034,N_14300,N_13309);
nand U17035 (N_17035,N_12585,N_13896);
nand U17036 (N_17036,N_14913,N_14045);
or U17037 (N_17037,N_14658,N_14280);
nand U17038 (N_17038,N_13506,N_14881);
xor U17039 (N_17039,N_14927,N_13805);
xnor U17040 (N_17040,N_12537,N_14827);
nand U17041 (N_17041,N_14330,N_13608);
xor U17042 (N_17042,N_13582,N_13129);
nor U17043 (N_17043,N_14341,N_13777);
or U17044 (N_17044,N_14371,N_13713);
or U17045 (N_17045,N_13105,N_13854);
nor U17046 (N_17046,N_12562,N_13443);
and U17047 (N_17047,N_13087,N_14737);
and U17048 (N_17048,N_14662,N_12812);
nor U17049 (N_17049,N_14256,N_14462);
nand U17050 (N_17050,N_13293,N_13257);
nor U17051 (N_17051,N_13963,N_14256);
nand U17052 (N_17052,N_13604,N_13740);
and U17053 (N_17053,N_12634,N_13320);
nor U17054 (N_17054,N_13268,N_14873);
nor U17055 (N_17055,N_13947,N_14587);
and U17056 (N_17056,N_14755,N_14223);
nand U17057 (N_17057,N_14345,N_14837);
nand U17058 (N_17058,N_14008,N_13732);
or U17059 (N_17059,N_14437,N_14397);
and U17060 (N_17060,N_13425,N_14543);
and U17061 (N_17061,N_13694,N_13295);
xor U17062 (N_17062,N_12939,N_13733);
xor U17063 (N_17063,N_12866,N_13090);
xnor U17064 (N_17064,N_13913,N_12634);
xnor U17065 (N_17065,N_13327,N_14861);
and U17066 (N_17066,N_14000,N_14460);
nor U17067 (N_17067,N_14751,N_12653);
nor U17068 (N_17068,N_14875,N_13994);
and U17069 (N_17069,N_13427,N_14389);
xor U17070 (N_17070,N_13183,N_13609);
xor U17071 (N_17071,N_14697,N_14352);
or U17072 (N_17072,N_12575,N_14065);
or U17073 (N_17073,N_13111,N_13145);
nand U17074 (N_17074,N_13093,N_13937);
and U17075 (N_17075,N_14991,N_14947);
nand U17076 (N_17076,N_14867,N_14261);
or U17077 (N_17077,N_13217,N_14564);
or U17078 (N_17078,N_14376,N_14445);
or U17079 (N_17079,N_14501,N_14342);
nor U17080 (N_17080,N_14761,N_14079);
and U17081 (N_17081,N_12912,N_14611);
or U17082 (N_17082,N_13748,N_14779);
or U17083 (N_17083,N_13312,N_14224);
nor U17084 (N_17084,N_14353,N_13953);
nor U17085 (N_17085,N_12632,N_14681);
nor U17086 (N_17086,N_13322,N_14078);
xnor U17087 (N_17087,N_14564,N_13879);
nor U17088 (N_17088,N_13343,N_12966);
or U17089 (N_17089,N_13669,N_13628);
nand U17090 (N_17090,N_14078,N_13563);
nand U17091 (N_17091,N_13013,N_14333);
or U17092 (N_17092,N_14297,N_14929);
xnor U17093 (N_17093,N_12686,N_14878);
nor U17094 (N_17094,N_13934,N_14548);
xor U17095 (N_17095,N_14481,N_12640);
nand U17096 (N_17096,N_14268,N_14683);
nor U17097 (N_17097,N_14440,N_13740);
and U17098 (N_17098,N_14612,N_12856);
nand U17099 (N_17099,N_14644,N_13044);
nor U17100 (N_17100,N_12855,N_12509);
and U17101 (N_17101,N_14675,N_13928);
nor U17102 (N_17102,N_12757,N_14864);
nand U17103 (N_17103,N_12604,N_14333);
nor U17104 (N_17104,N_12637,N_13346);
nand U17105 (N_17105,N_13235,N_14614);
or U17106 (N_17106,N_13288,N_14634);
xnor U17107 (N_17107,N_14532,N_14178);
xor U17108 (N_17108,N_14845,N_13460);
xor U17109 (N_17109,N_14665,N_14735);
xnor U17110 (N_17110,N_13219,N_12836);
and U17111 (N_17111,N_13338,N_14109);
or U17112 (N_17112,N_14133,N_14144);
nor U17113 (N_17113,N_14228,N_12668);
or U17114 (N_17114,N_14378,N_14070);
xor U17115 (N_17115,N_14608,N_12755);
and U17116 (N_17116,N_14573,N_14459);
or U17117 (N_17117,N_14568,N_13020);
nor U17118 (N_17118,N_14142,N_13973);
and U17119 (N_17119,N_13102,N_13460);
and U17120 (N_17120,N_13533,N_12546);
and U17121 (N_17121,N_13174,N_14330);
nand U17122 (N_17122,N_13416,N_14161);
nor U17123 (N_17123,N_13855,N_12893);
or U17124 (N_17124,N_13876,N_13014);
nor U17125 (N_17125,N_13311,N_12826);
or U17126 (N_17126,N_13420,N_12635);
xnor U17127 (N_17127,N_14429,N_13273);
nor U17128 (N_17128,N_12995,N_14885);
xnor U17129 (N_17129,N_12795,N_12632);
xnor U17130 (N_17130,N_12869,N_14350);
nor U17131 (N_17131,N_14203,N_13256);
xnor U17132 (N_17132,N_12630,N_13552);
nand U17133 (N_17133,N_14035,N_13327);
xnor U17134 (N_17134,N_12787,N_14022);
xor U17135 (N_17135,N_12529,N_12615);
or U17136 (N_17136,N_14675,N_13609);
nor U17137 (N_17137,N_14115,N_14914);
nor U17138 (N_17138,N_14459,N_13912);
xor U17139 (N_17139,N_14814,N_14018);
nor U17140 (N_17140,N_14196,N_12790);
or U17141 (N_17141,N_14951,N_13182);
nor U17142 (N_17142,N_13214,N_13143);
and U17143 (N_17143,N_14369,N_14855);
xor U17144 (N_17144,N_14988,N_13592);
xnor U17145 (N_17145,N_14342,N_12586);
nor U17146 (N_17146,N_13128,N_14750);
xor U17147 (N_17147,N_14886,N_14195);
xor U17148 (N_17148,N_13547,N_14174);
or U17149 (N_17149,N_13450,N_14152);
and U17150 (N_17150,N_13043,N_13462);
nor U17151 (N_17151,N_14713,N_12957);
nor U17152 (N_17152,N_12996,N_12635);
and U17153 (N_17153,N_14003,N_14931);
nand U17154 (N_17154,N_14819,N_13492);
xor U17155 (N_17155,N_12636,N_14634);
nand U17156 (N_17156,N_13097,N_13493);
and U17157 (N_17157,N_14871,N_14191);
and U17158 (N_17158,N_14035,N_12782);
xor U17159 (N_17159,N_14385,N_14934);
xnor U17160 (N_17160,N_13156,N_14936);
xnor U17161 (N_17161,N_13684,N_13148);
nor U17162 (N_17162,N_14908,N_14880);
and U17163 (N_17163,N_13634,N_14572);
and U17164 (N_17164,N_14455,N_12666);
nor U17165 (N_17165,N_14258,N_13378);
and U17166 (N_17166,N_13678,N_12860);
nand U17167 (N_17167,N_13110,N_14474);
or U17168 (N_17168,N_12874,N_14730);
nand U17169 (N_17169,N_13419,N_14370);
or U17170 (N_17170,N_14717,N_14796);
nor U17171 (N_17171,N_12671,N_13680);
and U17172 (N_17172,N_14968,N_13939);
nand U17173 (N_17173,N_14731,N_14454);
or U17174 (N_17174,N_14675,N_13682);
xor U17175 (N_17175,N_13049,N_13789);
nand U17176 (N_17176,N_13798,N_14497);
nor U17177 (N_17177,N_12588,N_12866);
or U17178 (N_17178,N_13534,N_12794);
xor U17179 (N_17179,N_13972,N_14531);
xor U17180 (N_17180,N_14484,N_14653);
or U17181 (N_17181,N_12617,N_13504);
nand U17182 (N_17182,N_14773,N_14461);
xnor U17183 (N_17183,N_12744,N_13109);
xnor U17184 (N_17184,N_13738,N_13281);
nor U17185 (N_17185,N_12699,N_13948);
and U17186 (N_17186,N_13949,N_13984);
nor U17187 (N_17187,N_12597,N_13357);
or U17188 (N_17188,N_13803,N_14077);
nor U17189 (N_17189,N_13556,N_13958);
nor U17190 (N_17190,N_14165,N_14464);
nand U17191 (N_17191,N_13024,N_13617);
nor U17192 (N_17192,N_14699,N_14996);
and U17193 (N_17193,N_14122,N_14498);
xor U17194 (N_17194,N_14460,N_13131);
and U17195 (N_17195,N_13184,N_12628);
nor U17196 (N_17196,N_13165,N_12935);
nor U17197 (N_17197,N_14896,N_14020);
or U17198 (N_17198,N_13273,N_13065);
nor U17199 (N_17199,N_12816,N_14463);
or U17200 (N_17200,N_13635,N_14523);
or U17201 (N_17201,N_13570,N_12659);
and U17202 (N_17202,N_13763,N_14462);
nor U17203 (N_17203,N_12896,N_14202);
xnor U17204 (N_17204,N_14335,N_14651);
nand U17205 (N_17205,N_14130,N_14720);
or U17206 (N_17206,N_13641,N_14604);
nor U17207 (N_17207,N_13092,N_12517);
or U17208 (N_17208,N_14365,N_14807);
nand U17209 (N_17209,N_13249,N_13440);
nand U17210 (N_17210,N_13170,N_13568);
nand U17211 (N_17211,N_14896,N_12939);
and U17212 (N_17212,N_14966,N_13491);
and U17213 (N_17213,N_13698,N_14636);
or U17214 (N_17214,N_13261,N_13150);
or U17215 (N_17215,N_12533,N_13337);
nand U17216 (N_17216,N_12574,N_14791);
nand U17217 (N_17217,N_13172,N_14376);
or U17218 (N_17218,N_12550,N_13842);
nand U17219 (N_17219,N_13708,N_14317);
or U17220 (N_17220,N_13449,N_14457);
nor U17221 (N_17221,N_13962,N_14695);
xnor U17222 (N_17222,N_13373,N_14634);
xor U17223 (N_17223,N_14684,N_14236);
nor U17224 (N_17224,N_13766,N_14636);
or U17225 (N_17225,N_14523,N_14508);
and U17226 (N_17226,N_14645,N_12588);
nor U17227 (N_17227,N_14068,N_13683);
or U17228 (N_17228,N_12869,N_14366);
or U17229 (N_17229,N_14710,N_14896);
and U17230 (N_17230,N_13354,N_12509);
or U17231 (N_17231,N_14150,N_13955);
nor U17232 (N_17232,N_14768,N_13089);
and U17233 (N_17233,N_12899,N_14111);
xor U17234 (N_17234,N_12896,N_13298);
nand U17235 (N_17235,N_13608,N_12976);
nand U17236 (N_17236,N_12655,N_13308);
xor U17237 (N_17237,N_12670,N_13047);
or U17238 (N_17238,N_12543,N_14516);
and U17239 (N_17239,N_12898,N_13464);
nand U17240 (N_17240,N_12725,N_14141);
xor U17241 (N_17241,N_13480,N_14266);
xnor U17242 (N_17242,N_14535,N_12939);
nor U17243 (N_17243,N_12856,N_13011);
xor U17244 (N_17244,N_13311,N_13261);
and U17245 (N_17245,N_13722,N_14574);
nand U17246 (N_17246,N_13629,N_12937);
or U17247 (N_17247,N_14659,N_13333);
nand U17248 (N_17248,N_13654,N_13161);
nor U17249 (N_17249,N_14961,N_13200);
xor U17250 (N_17250,N_12682,N_14184);
and U17251 (N_17251,N_12721,N_14592);
xor U17252 (N_17252,N_13088,N_12692);
nand U17253 (N_17253,N_12695,N_13785);
or U17254 (N_17254,N_13421,N_13939);
nand U17255 (N_17255,N_13390,N_12753);
or U17256 (N_17256,N_12673,N_14214);
xor U17257 (N_17257,N_12985,N_13393);
nand U17258 (N_17258,N_13125,N_13787);
and U17259 (N_17259,N_13664,N_12981);
xnor U17260 (N_17260,N_14470,N_14387);
and U17261 (N_17261,N_13962,N_13229);
or U17262 (N_17262,N_13725,N_14627);
and U17263 (N_17263,N_13609,N_13861);
xnor U17264 (N_17264,N_14571,N_14749);
and U17265 (N_17265,N_14387,N_12880);
xor U17266 (N_17266,N_13889,N_14360);
xor U17267 (N_17267,N_14475,N_14298);
or U17268 (N_17268,N_13337,N_13805);
xor U17269 (N_17269,N_13323,N_14925);
nor U17270 (N_17270,N_13737,N_14094);
nor U17271 (N_17271,N_14746,N_13140);
nand U17272 (N_17272,N_14018,N_14077);
xnor U17273 (N_17273,N_13099,N_14561);
and U17274 (N_17274,N_14282,N_14149);
or U17275 (N_17275,N_13298,N_13401);
or U17276 (N_17276,N_13591,N_14813);
xnor U17277 (N_17277,N_13239,N_12934);
xnor U17278 (N_17278,N_13796,N_13878);
nand U17279 (N_17279,N_13956,N_14411);
xnor U17280 (N_17280,N_13759,N_14991);
nor U17281 (N_17281,N_13933,N_13353);
nand U17282 (N_17282,N_13543,N_13521);
nor U17283 (N_17283,N_13523,N_12816);
or U17284 (N_17284,N_12783,N_13493);
nand U17285 (N_17285,N_14905,N_14616);
nand U17286 (N_17286,N_13084,N_13879);
and U17287 (N_17287,N_14699,N_14295);
and U17288 (N_17288,N_13687,N_14446);
nor U17289 (N_17289,N_12730,N_14323);
or U17290 (N_17290,N_13039,N_13614);
nand U17291 (N_17291,N_13215,N_13698);
or U17292 (N_17292,N_13434,N_14098);
and U17293 (N_17293,N_14071,N_13831);
or U17294 (N_17294,N_14975,N_13371);
nand U17295 (N_17295,N_13373,N_14569);
nor U17296 (N_17296,N_14249,N_13368);
nor U17297 (N_17297,N_14671,N_13573);
nand U17298 (N_17298,N_13323,N_12619);
or U17299 (N_17299,N_13500,N_13073);
nand U17300 (N_17300,N_14838,N_14962);
and U17301 (N_17301,N_12515,N_13590);
xnor U17302 (N_17302,N_14767,N_13002);
and U17303 (N_17303,N_13379,N_12960);
nor U17304 (N_17304,N_14678,N_13013);
or U17305 (N_17305,N_14760,N_12883);
nor U17306 (N_17306,N_12679,N_13065);
nand U17307 (N_17307,N_14404,N_14118);
nand U17308 (N_17308,N_14863,N_13424);
nor U17309 (N_17309,N_12844,N_12621);
xor U17310 (N_17310,N_14186,N_14172);
nor U17311 (N_17311,N_12558,N_14930);
or U17312 (N_17312,N_14414,N_13954);
and U17313 (N_17313,N_13955,N_12694);
or U17314 (N_17314,N_12939,N_13721);
nand U17315 (N_17315,N_14095,N_12646);
nand U17316 (N_17316,N_13524,N_14295);
nand U17317 (N_17317,N_12724,N_13452);
xor U17318 (N_17318,N_12505,N_14416);
or U17319 (N_17319,N_14514,N_14533);
or U17320 (N_17320,N_13917,N_13932);
or U17321 (N_17321,N_13566,N_13352);
or U17322 (N_17322,N_14586,N_12613);
or U17323 (N_17323,N_13392,N_13680);
xnor U17324 (N_17324,N_12887,N_13339);
nor U17325 (N_17325,N_12772,N_13672);
or U17326 (N_17326,N_14712,N_14008);
nor U17327 (N_17327,N_12777,N_12905);
and U17328 (N_17328,N_13080,N_13567);
nand U17329 (N_17329,N_13679,N_14552);
nor U17330 (N_17330,N_13190,N_12556);
nor U17331 (N_17331,N_13886,N_13333);
or U17332 (N_17332,N_14560,N_13419);
or U17333 (N_17333,N_13127,N_12862);
and U17334 (N_17334,N_14106,N_14496);
and U17335 (N_17335,N_14988,N_14647);
xnor U17336 (N_17336,N_14697,N_13905);
or U17337 (N_17337,N_12758,N_14178);
or U17338 (N_17338,N_14345,N_14602);
xnor U17339 (N_17339,N_12692,N_13936);
xnor U17340 (N_17340,N_12698,N_12547);
nand U17341 (N_17341,N_13520,N_13376);
xnor U17342 (N_17342,N_13859,N_14361);
nand U17343 (N_17343,N_13387,N_13190);
nand U17344 (N_17344,N_12665,N_12908);
nor U17345 (N_17345,N_13484,N_12576);
nand U17346 (N_17346,N_12906,N_13333);
and U17347 (N_17347,N_13922,N_12786);
or U17348 (N_17348,N_12998,N_12713);
nor U17349 (N_17349,N_12516,N_13871);
nor U17350 (N_17350,N_14272,N_14189);
or U17351 (N_17351,N_13288,N_12918);
and U17352 (N_17352,N_13704,N_13151);
or U17353 (N_17353,N_13943,N_14003);
or U17354 (N_17354,N_13558,N_13187);
xor U17355 (N_17355,N_13358,N_14672);
and U17356 (N_17356,N_12623,N_13192);
nor U17357 (N_17357,N_13379,N_13369);
or U17358 (N_17358,N_14054,N_13969);
xnor U17359 (N_17359,N_14288,N_14497);
xor U17360 (N_17360,N_13357,N_13870);
xnor U17361 (N_17361,N_12642,N_13319);
or U17362 (N_17362,N_14477,N_13325);
nand U17363 (N_17363,N_14824,N_12573);
or U17364 (N_17364,N_12811,N_13841);
xnor U17365 (N_17365,N_12662,N_14501);
or U17366 (N_17366,N_12800,N_14288);
or U17367 (N_17367,N_14692,N_13195);
nand U17368 (N_17368,N_13795,N_13353);
or U17369 (N_17369,N_13588,N_14341);
and U17370 (N_17370,N_14839,N_14350);
xnor U17371 (N_17371,N_13800,N_13761);
nor U17372 (N_17372,N_14766,N_13793);
nor U17373 (N_17373,N_14471,N_12557);
and U17374 (N_17374,N_12885,N_13669);
nand U17375 (N_17375,N_12580,N_12957);
or U17376 (N_17376,N_13934,N_12589);
nor U17377 (N_17377,N_13560,N_12836);
or U17378 (N_17378,N_12979,N_14263);
nand U17379 (N_17379,N_14326,N_12850);
or U17380 (N_17380,N_13945,N_13605);
nand U17381 (N_17381,N_13732,N_13737);
or U17382 (N_17382,N_13482,N_14262);
and U17383 (N_17383,N_14541,N_14941);
or U17384 (N_17384,N_13035,N_14969);
or U17385 (N_17385,N_14690,N_13414);
nand U17386 (N_17386,N_12942,N_14706);
and U17387 (N_17387,N_14859,N_13361);
nor U17388 (N_17388,N_14047,N_14670);
xor U17389 (N_17389,N_14688,N_13107);
nor U17390 (N_17390,N_14820,N_14017);
and U17391 (N_17391,N_14677,N_13715);
nor U17392 (N_17392,N_13507,N_13482);
and U17393 (N_17393,N_13244,N_13193);
nor U17394 (N_17394,N_12975,N_12765);
and U17395 (N_17395,N_14669,N_14925);
nand U17396 (N_17396,N_12539,N_14065);
and U17397 (N_17397,N_14837,N_13991);
or U17398 (N_17398,N_12954,N_14831);
xnor U17399 (N_17399,N_12764,N_14743);
and U17400 (N_17400,N_14374,N_13451);
or U17401 (N_17401,N_14745,N_14017);
xor U17402 (N_17402,N_14066,N_13835);
nor U17403 (N_17403,N_12513,N_12806);
nor U17404 (N_17404,N_12767,N_13773);
nor U17405 (N_17405,N_13447,N_13761);
nand U17406 (N_17406,N_13876,N_14125);
xor U17407 (N_17407,N_14316,N_13375);
xor U17408 (N_17408,N_14150,N_14219);
xnor U17409 (N_17409,N_13061,N_12790);
or U17410 (N_17410,N_13626,N_13365);
and U17411 (N_17411,N_14603,N_14432);
nor U17412 (N_17412,N_14626,N_14808);
xnor U17413 (N_17413,N_12893,N_13919);
xor U17414 (N_17414,N_14027,N_14307);
and U17415 (N_17415,N_13928,N_14906);
nand U17416 (N_17416,N_13686,N_14964);
nand U17417 (N_17417,N_12672,N_13650);
nand U17418 (N_17418,N_14732,N_12833);
nand U17419 (N_17419,N_13039,N_14214);
nor U17420 (N_17420,N_14191,N_13797);
and U17421 (N_17421,N_13296,N_14485);
and U17422 (N_17422,N_13983,N_13458);
nand U17423 (N_17423,N_14279,N_14258);
and U17424 (N_17424,N_12933,N_14613);
and U17425 (N_17425,N_12911,N_14773);
nor U17426 (N_17426,N_13371,N_12667);
nand U17427 (N_17427,N_14285,N_13230);
nand U17428 (N_17428,N_13932,N_12677);
xor U17429 (N_17429,N_14013,N_14308);
xor U17430 (N_17430,N_13920,N_13699);
nand U17431 (N_17431,N_13302,N_14398);
and U17432 (N_17432,N_13976,N_13035);
and U17433 (N_17433,N_12801,N_14118);
or U17434 (N_17434,N_13219,N_14745);
and U17435 (N_17435,N_14706,N_13510);
or U17436 (N_17436,N_14850,N_14187);
nor U17437 (N_17437,N_12832,N_14369);
or U17438 (N_17438,N_14644,N_13985);
nor U17439 (N_17439,N_14689,N_13994);
xnor U17440 (N_17440,N_14330,N_14006);
and U17441 (N_17441,N_12596,N_13790);
nor U17442 (N_17442,N_12868,N_13825);
nand U17443 (N_17443,N_14470,N_12995);
nor U17444 (N_17444,N_12658,N_14335);
nand U17445 (N_17445,N_13755,N_13584);
nand U17446 (N_17446,N_12722,N_13218);
xor U17447 (N_17447,N_13272,N_12578);
and U17448 (N_17448,N_12923,N_14387);
nand U17449 (N_17449,N_14129,N_14103);
xnor U17450 (N_17450,N_14456,N_14300);
nor U17451 (N_17451,N_14483,N_14889);
nand U17452 (N_17452,N_12834,N_14788);
nand U17453 (N_17453,N_13046,N_13229);
nand U17454 (N_17454,N_12610,N_13238);
or U17455 (N_17455,N_13526,N_13782);
nand U17456 (N_17456,N_13047,N_13766);
and U17457 (N_17457,N_13884,N_12879);
or U17458 (N_17458,N_14599,N_13690);
and U17459 (N_17459,N_13000,N_12989);
and U17460 (N_17460,N_14414,N_13528);
and U17461 (N_17461,N_13415,N_13660);
nand U17462 (N_17462,N_14901,N_14574);
nand U17463 (N_17463,N_14553,N_12618);
and U17464 (N_17464,N_13477,N_14852);
and U17465 (N_17465,N_13564,N_13963);
and U17466 (N_17466,N_14276,N_13957);
nor U17467 (N_17467,N_14545,N_12973);
nor U17468 (N_17468,N_14509,N_14803);
and U17469 (N_17469,N_13356,N_13069);
nor U17470 (N_17470,N_13246,N_13768);
and U17471 (N_17471,N_13866,N_14499);
nand U17472 (N_17472,N_13083,N_13335);
nor U17473 (N_17473,N_12999,N_14260);
or U17474 (N_17474,N_13503,N_14081);
nor U17475 (N_17475,N_13667,N_13867);
nand U17476 (N_17476,N_13397,N_13374);
or U17477 (N_17477,N_13045,N_13572);
or U17478 (N_17478,N_12755,N_13480);
nand U17479 (N_17479,N_13451,N_13950);
nand U17480 (N_17480,N_14091,N_13520);
xnor U17481 (N_17481,N_13795,N_12543);
and U17482 (N_17482,N_12642,N_14698);
and U17483 (N_17483,N_13915,N_13708);
nand U17484 (N_17484,N_14318,N_14575);
or U17485 (N_17485,N_12909,N_13629);
or U17486 (N_17486,N_14183,N_13568);
nor U17487 (N_17487,N_13803,N_14453);
nor U17488 (N_17488,N_14399,N_14022);
and U17489 (N_17489,N_14849,N_13629);
nor U17490 (N_17490,N_13810,N_12593);
xnor U17491 (N_17491,N_14140,N_12785);
and U17492 (N_17492,N_13012,N_14187);
nand U17493 (N_17493,N_12964,N_13927);
and U17494 (N_17494,N_14556,N_14678);
or U17495 (N_17495,N_14532,N_12917);
or U17496 (N_17496,N_13574,N_14934);
nor U17497 (N_17497,N_14651,N_14313);
nand U17498 (N_17498,N_13359,N_13588);
nand U17499 (N_17499,N_14154,N_14858);
and U17500 (N_17500,N_16033,N_17193);
xnor U17501 (N_17501,N_16654,N_15768);
nor U17502 (N_17502,N_17463,N_16308);
and U17503 (N_17503,N_16766,N_16994);
and U17504 (N_17504,N_17179,N_16188);
or U17505 (N_17505,N_16622,N_17165);
or U17506 (N_17506,N_17414,N_16331);
nor U17507 (N_17507,N_15987,N_15847);
nand U17508 (N_17508,N_16614,N_15219);
nand U17509 (N_17509,N_15975,N_15422);
or U17510 (N_17510,N_15401,N_16703);
or U17511 (N_17511,N_16248,N_16442);
xnor U17512 (N_17512,N_15352,N_15076);
xor U17513 (N_17513,N_17181,N_17250);
and U17514 (N_17514,N_15146,N_15719);
xor U17515 (N_17515,N_17082,N_15537);
nor U17516 (N_17516,N_16446,N_15504);
xor U17517 (N_17517,N_15350,N_17262);
nor U17518 (N_17518,N_16548,N_16841);
and U17519 (N_17519,N_15115,N_15845);
nor U17520 (N_17520,N_15986,N_15641);
nor U17521 (N_17521,N_16128,N_16275);
or U17522 (N_17522,N_17091,N_16046);
nand U17523 (N_17523,N_16170,N_15091);
or U17524 (N_17524,N_15258,N_16891);
xnor U17525 (N_17525,N_16776,N_16850);
or U17526 (N_17526,N_16250,N_16296);
nor U17527 (N_17527,N_15682,N_15131);
nand U17528 (N_17528,N_16863,N_16177);
nand U17529 (N_17529,N_16943,N_15532);
and U17530 (N_17530,N_16484,N_15929);
xnor U17531 (N_17531,N_17290,N_16328);
nand U17532 (N_17532,N_15985,N_15229);
nand U17533 (N_17533,N_16745,N_17349);
xnor U17534 (N_17534,N_15110,N_16557);
nand U17535 (N_17535,N_15052,N_16110);
nor U17536 (N_17536,N_16507,N_17010);
and U17537 (N_17537,N_15180,N_16203);
and U17538 (N_17538,N_15775,N_15107);
nand U17539 (N_17539,N_17031,N_15758);
or U17540 (N_17540,N_15306,N_16349);
xor U17541 (N_17541,N_16431,N_15453);
or U17542 (N_17542,N_16474,N_15512);
and U17543 (N_17543,N_15857,N_17163);
xnor U17544 (N_17544,N_16939,N_16322);
and U17545 (N_17545,N_16695,N_16652);
nand U17546 (N_17546,N_15884,N_17231);
or U17547 (N_17547,N_15867,N_16213);
nand U17548 (N_17548,N_16993,N_17417);
or U17549 (N_17549,N_15982,N_16959);
or U17550 (N_17550,N_15676,N_16989);
xor U17551 (N_17551,N_17172,N_17470);
or U17552 (N_17552,N_15941,N_15441);
nand U17553 (N_17553,N_15232,N_16179);
and U17554 (N_17554,N_15741,N_16491);
xor U17555 (N_17555,N_17076,N_17190);
nor U17556 (N_17556,N_15816,N_15480);
nor U17557 (N_17557,N_16769,N_16343);
nor U17558 (N_17558,N_16635,N_16668);
nand U17559 (N_17559,N_15235,N_15157);
nor U17560 (N_17560,N_15151,N_16830);
or U17561 (N_17561,N_15317,N_15086);
xor U17562 (N_17562,N_16969,N_16547);
and U17563 (N_17563,N_16353,N_16027);
or U17564 (N_17564,N_16812,N_15438);
nand U17565 (N_17565,N_16590,N_16242);
nor U17566 (N_17566,N_15088,N_17473);
nand U17567 (N_17567,N_15749,N_17399);
nand U17568 (N_17568,N_16777,N_17438);
xor U17569 (N_17569,N_16999,N_15646);
nand U17570 (N_17570,N_16517,N_17089);
nor U17571 (N_17571,N_16187,N_17067);
or U17572 (N_17572,N_16166,N_16913);
and U17573 (N_17573,N_15804,N_16858);
nand U17574 (N_17574,N_16174,N_16335);
or U17575 (N_17575,N_16054,N_16161);
or U17576 (N_17576,N_16350,N_17126);
nor U17577 (N_17577,N_15835,N_17327);
xor U17578 (N_17578,N_15871,N_15283);
nand U17579 (N_17579,N_17061,N_15405);
and U17580 (N_17580,N_16092,N_15409);
or U17581 (N_17581,N_16230,N_17324);
xor U17582 (N_17582,N_15949,N_15234);
or U17583 (N_17583,N_16996,N_15527);
nor U17584 (N_17584,N_16060,N_16820);
nand U17585 (N_17585,N_17397,N_17107);
nor U17586 (N_17586,N_16219,N_15736);
xor U17587 (N_17587,N_17451,N_16411);
nand U17588 (N_17588,N_17162,N_16995);
nand U17589 (N_17589,N_16458,N_15842);
or U17590 (N_17590,N_17032,N_16937);
and U17591 (N_17591,N_15520,N_16782);
nor U17592 (N_17592,N_17015,N_16558);
or U17593 (N_17593,N_15491,N_16655);
and U17594 (N_17594,N_17467,N_15464);
and U17595 (N_17595,N_17127,N_15266);
and U17596 (N_17596,N_16261,N_16816);
nand U17597 (N_17597,N_16675,N_16220);
xor U17598 (N_17598,N_16665,N_15956);
xnor U17599 (N_17599,N_15497,N_15993);
or U17600 (N_17600,N_15068,N_16045);
or U17601 (N_17601,N_16511,N_17167);
and U17602 (N_17602,N_16382,N_15299);
and U17603 (N_17603,N_16566,N_17450);
nand U17604 (N_17604,N_15962,N_17045);
nor U17605 (N_17605,N_16029,N_16086);
nand U17606 (N_17606,N_16498,N_15057);
nand U17607 (N_17607,N_15353,N_16643);
and U17608 (N_17608,N_17355,N_16103);
nor U17609 (N_17609,N_16083,N_16537);
or U17610 (N_17610,N_15218,N_15097);
xnor U17611 (N_17611,N_15499,N_15034);
and U17612 (N_17612,N_15081,N_15495);
and U17613 (N_17613,N_16553,N_15386);
nand U17614 (N_17614,N_16581,N_15398);
or U17615 (N_17615,N_17444,N_15293);
and U17616 (N_17616,N_16157,N_15292);
nand U17617 (N_17617,N_15957,N_15319);
and U17618 (N_17618,N_17499,N_16818);
or U17619 (N_17619,N_16741,N_15139);
xnor U17620 (N_17620,N_16975,N_17175);
and U17621 (N_17621,N_16210,N_17445);
nor U17622 (N_17622,N_17209,N_16222);
or U17623 (N_17623,N_15140,N_16833);
nor U17624 (N_17624,N_16535,N_16181);
and U17625 (N_17625,N_15169,N_17459);
and U17626 (N_17626,N_17103,N_17096);
xor U17627 (N_17627,N_16062,N_16194);
and U17628 (N_17628,N_15150,N_16823);
nand U17629 (N_17629,N_16929,N_16737);
and U17630 (N_17630,N_15175,N_16567);
nor U17631 (N_17631,N_15814,N_16888);
nor U17632 (N_17632,N_16738,N_16360);
or U17633 (N_17633,N_17489,N_17353);
xor U17634 (N_17634,N_16512,N_16634);
and U17635 (N_17635,N_16319,N_16878);
xor U17636 (N_17636,N_16910,N_16066);
nand U17637 (N_17637,N_16619,N_15199);
nand U17638 (N_17638,N_17074,N_15083);
nor U17639 (N_17639,N_16272,N_15723);
nor U17640 (N_17640,N_15274,N_15851);
xnor U17641 (N_17641,N_15074,N_15357);
nor U17642 (N_17642,N_16361,N_15263);
or U17643 (N_17643,N_16167,N_17079);
nor U17644 (N_17644,N_15643,N_15481);
xor U17645 (N_17645,N_17288,N_16724);
nand U17646 (N_17646,N_15531,N_15567);
and U17647 (N_17647,N_15735,N_15800);
and U17648 (N_17648,N_16778,N_16490);
xor U17649 (N_17649,N_17068,N_15983);
nor U17650 (N_17650,N_17028,N_17111);
nand U17651 (N_17651,N_16716,N_17233);
xnor U17652 (N_17652,N_16928,N_15062);
and U17653 (N_17653,N_16692,N_15840);
nor U17654 (N_17654,N_15533,N_17035);
xor U17655 (N_17655,N_15012,N_15689);
nand U17656 (N_17656,N_15227,N_15554);
or U17657 (N_17657,N_15203,N_16726);
and U17658 (N_17658,N_15702,N_15466);
xnor U17659 (N_17659,N_16464,N_17384);
and U17660 (N_17660,N_16785,N_16415);
nor U17661 (N_17661,N_16405,N_16286);
or U17662 (N_17662,N_16666,N_15479);
or U17663 (N_17663,N_15112,N_15378);
nand U17664 (N_17664,N_16001,N_16529);
or U17665 (N_17665,N_16825,N_17310);
xnor U17666 (N_17666,N_17066,N_15449);
xnor U17667 (N_17667,N_15552,N_17346);
xnor U17668 (N_17668,N_15874,N_16217);
nor U17669 (N_17669,N_17457,N_15400);
xor U17670 (N_17670,N_16292,N_15577);
nor U17671 (N_17671,N_16224,N_16615);
xor U17672 (N_17672,N_15674,N_15490);
xnor U17673 (N_17673,N_16679,N_16199);
xor U17674 (N_17674,N_15542,N_16673);
or U17675 (N_17675,N_17157,N_15442);
xor U17676 (N_17676,N_16333,N_16043);
and U17677 (N_17677,N_16182,N_15233);
nor U17678 (N_17678,N_17282,N_15048);
nand U17679 (N_17679,N_16632,N_15320);
and U17680 (N_17680,N_15692,N_16425);
xnor U17681 (N_17681,N_15316,N_17350);
xor U17682 (N_17682,N_15767,N_15456);
or U17683 (N_17683,N_16662,N_16075);
nand U17684 (N_17684,N_16427,N_15436);
nand U17685 (N_17685,N_15226,N_16357);
nand U17686 (N_17686,N_16712,N_15372);
nand U17687 (N_17687,N_17478,N_15469);
xor U17688 (N_17688,N_15870,N_15955);
nand U17689 (N_17689,N_15657,N_16421);
and U17690 (N_17690,N_15889,N_16122);
nand U17691 (N_17691,N_15637,N_17276);
xnor U17692 (N_17692,N_16889,N_15318);
xnor U17693 (N_17693,N_17189,N_15358);
nand U17694 (N_17694,N_16258,N_16298);
nor U17695 (N_17695,N_16789,N_15925);
or U17696 (N_17696,N_15948,N_16400);
and U17697 (N_17697,N_15555,N_16836);
or U17698 (N_17698,N_16480,N_15731);
nor U17699 (N_17699,N_17090,N_17294);
nand U17700 (N_17700,N_16503,N_17483);
nand U17701 (N_17701,N_16905,N_15450);
xor U17702 (N_17702,N_16096,N_17016);
and U17703 (N_17703,N_17302,N_17249);
nor U17704 (N_17704,N_15311,N_15045);
and U17705 (N_17705,N_16014,N_15212);
xor U17706 (N_17706,N_16533,N_16306);
nand U17707 (N_17707,N_15943,N_16365);
and U17708 (N_17708,N_16051,N_17030);
nor U17709 (N_17709,N_17008,N_17306);
and U17710 (N_17710,N_17143,N_17370);
or U17711 (N_17711,N_16564,N_15394);
nor U17712 (N_17712,N_15668,N_15762);
nand U17713 (N_17713,N_16282,N_15451);
nand U17714 (N_17714,N_15678,N_16762);
xor U17715 (N_17715,N_16618,N_15772);
xnor U17716 (N_17716,N_17320,N_15244);
and U17717 (N_17717,N_17130,N_17460);
and U17718 (N_17718,N_16974,N_17264);
or U17719 (N_17719,N_15710,N_15715);
nor U17720 (N_17720,N_16031,N_15416);
xor U17721 (N_17721,N_15790,N_16388);
nand U17722 (N_17722,N_17206,N_15304);
and U17723 (N_17723,N_15006,N_17464);
nor U17724 (N_17724,N_16922,N_15653);
nand U17725 (N_17725,N_16853,N_16893);
xnor U17726 (N_17726,N_15765,N_15298);
nand U17727 (N_17727,N_15429,N_16926);
nand U17728 (N_17728,N_15435,N_15858);
or U17729 (N_17729,N_17319,N_15138);
nor U17730 (N_17730,N_17124,N_15652);
nand U17731 (N_17731,N_17495,N_16821);
and U17732 (N_17732,N_15265,N_15716);
xnor U17733 (N_17733,N_17223,N_16265);
nor U17734 (N_17734,N_15606,N_17252);
and U17735 (N_17735,N_17420,N_15954);
nand U17736 (N_17736,N_16805,N_16397);
xnor U17737 (N_17737,N_17094,N_17227);
nand U17738 (N_17738,N_17177,N_15005);
nor U17739 (N_17739,N_15132,N_16580);
and U17740 (N_17740,N_16918,N_17184);
and U17741 (N_17741,N_16753,N_17154);
nor U17742 (N_17742,N_16563,N_16208);
and U17743 (N_17743,N_16859,N_16664);
and U17744 (N_17744,N_17213,N_16460);
nand U17745 (N_17745,N_16793,N_17001);
nor U17746 (N_17746,N_16583,N_15739);
xnor U17747 (N_17747,N_15301,N_15486);
or U17748 (N_17748,N_17307,N_16587);
nand U17749 (N_17749,N_15341,N_17278);
nor U17750 (N_17750,N_15748,N_16794);
xor U17751 (N_17751,N_15043,N_15952);
xnor U17752 (N_17752,N_15037,N_16348);
nand U17753 (N_17753,N_17468,N_15694);
or U17754 (N_17754,N_17055,N_15278);
and U17755 (N_17755,N_17121,N_15620);
nor U17756 (N_17756,N_15902,N_15145);
nand U17757 (N_17757,N_17214,N_16534);
nand U17758 (N_17758,N_16815,N_17208);
xnor U17759 (N_17759,N_16351,N_15705);
or U17760 (N_17760,N_15404,N_15166);
and U17761 (N_17761,N_17312,N_17078);
nor U17762 (N_17762,N_16882,N_16118);
nand U17763 (N_17763,N_15868,N_16426);
nand U17764 (N_17764,N_17012,N_16002);
nand U17765 (N_17765,N_15246,N_17202);
nor U17766 (N_17766,N_15224,N_15573);
nor U17767 (N_17767,N_16585,N_15645);
xor U17768 (N_17768,N_17396,N_17337);
and U17769 (N_17769,N_15465,N_16921);
xnor U17770 (N_17770,N_16986,N_16711);
nor U17771 (N_17771,N_15025,N_16438);
xor U17772 (N_17772,N_16809,N_15369);
xor U17773 (N_17773,N_17421,N_17073);
nand U17774 (N_17774,N_15272,N_17474);
xnor U17775 (N_17775,N_15100,N_17205);
and U17776 (N_17776,N_16706,N_16621);
or U17777 (N_17777,N_16612,N_15934);
nor U17778 (N_17778,N_15104,N_17063);
nand U17779 (N_17779,N_16115,N_15393);
and U17780 (N_17780,N_15382,N_17149);
nand U17781 (N_17781,N_16617,N_15323);
nand U17782 (N_17782,N_16441,N_16339);
xnor U17783 (N_17783,N_17259,N_15011);
and U17784 (N_17784,N_16379,N_16672);
nand U17785 (N_17785,N_15594,N_16304);
nand U17786 (N_17786,N_16856,N_16920);
and U17787 (N_17787,N_15904,N_17338);
or U17788 (N_17788,N_16680,N_15519);
or U17789 (N_17789,N_15428,N_16952);
nand U17790 (N_17790,N_15467,N_15154);
nor U17791 (N_17791,N_16398,N_16964);
or U17792 (N_17792,N_16352,N_15658);
nor U17793 (N_17793,N_17007,N_15834);
or U17794 (N_17794,N_15707,N_16131);
nor U17795 (N_17795,N_16881,N_15538);
and U17796 (N_17796,N_16443,N_15782);
nand U17797 (N_17797,N_16895,N_17357);
xnor U17798 (N_17798,N_17148,N_17363);
and U17799 (N_17799,N_15918,N_15172);
and U17800 (N_17800,N_16984,N_16914);
xnor U17801 (N_17801,N_17038,N_16746);
xnor U17802 (N_17802,N_16731,N_17416);
nand U17803 (N_17803,N_15738,N_15628);
or U17804 (N_17804,N_15286,N_15970);
nand U17805 (N_17805,N_17486,N_16049);
xor U17806 (N_17806,N_16842,N_15873);
and U17807 (N_17807,N_17274,N_16908);
nand U17808 (N_17808,N_15002,N_16770);
nand U17809 (N_17809,N_15354,N_16288);
nand U17810 (N_17810,N_17328,N_15262);
and U17811 (N_17811,N_15066,N_15536);
and U17812 (N_17812,N_16671,N_16028);
nand U17813 (N_17813,N_15992,N_16477);
or U17814 (N_17814,N_15186,N_16467);
or U17815 (N_17815,N_15388,N_16890);
and U17816 (N_17816,N_16834,N_15410);
nand U17817 (N_17817,N_16356,N_15122);
or U17818 (N_17818,N_15756,N_16748);
or U17819 (N_17819,N_15093,N_16197);
nor U17820 (N_17820,N_15806,N_16932);
nor U17821 (N_17821,N_15377,N_16101);
xor U17822 (N_17822,N_15389,N_17442);
nand U17823 (N_17823,N_16325,N_15463);
xnor U17824 (N_17824,N_15528,N_16479);
or U17825 (N_17825,N_17062,N_16681);
or U17826 (N_17826,N_17323,N_16935);
xor U17827 (N_17827,N_17374,N_17358);
nand U17828 (N_17828,N_15271,N_15124);
xnor U17829 (N_17829,N_15908,N_15861);
or U17830 (N_17830,N_16779,N_16623);
nor U17831 (N_17831,N_15901,N_15371);
nand U17832 (N_17832,N_15725,N_17431);
nor U17833 (N_17833,N_16494,N_15510);
or U17834 (N_17834,N_16866,N_16252);
and U17835 (N_17835,N_15345,N_15050);
and U17836 (N_17836,N_15280,N_15018);
nor U17837 (N_17837,N_15558,N_16551);
and U17838 (N_17838,N_17301,N_15294);
nand U17839 (N_17839,N_16034,N_16301);
nor U17840 (N_17840,N_15875,N_15656);
nand U17841 (N_17841,N_16933,N_16981);
xnor U17842 (N_17842,N_16404,N_15004);
nand U17843 (N_17843,N_15055,N_16951);
xnor U17844 (N_17844,N_16368,N_15763);
nand U17845 (N_17845,N_16098,N_17222);
and U17846 (N_17846,N_16667,N_16297);
and U17847 (N_17847,N_15113,N_16663);
xor U17848 (N_17848,N_16829,N_16541);
xor U17849 (N_17849,N_16844,N_17427);
xnor U17850 (N_17850,N_17196,N_15644);
or U17851 (N_17851,N_16316,N_17492);
nor U17852 (N_17852,N_16649,N_15712);
or U17853 (N_17853,N_15213,N_15296);
or U17854 (N_17854,N_15133,N_15215);
nor U17855 (N_17855,N_16983,N_16992);
nand U17856 (N_17856,N_17439,N_17230);
xnor U17857 (N_17857,N_15604,N_16684);
or U17858 (N_17858,N_16150,N_15828);
nand U17859 (N_17859,N_15187,N_15195);
and U17860 (N_17860,N_15204,N_15717);
or U17861 (N_17861,N_15830,N_15667);
xnor U17862 (N_17862,N_17160,N_15448);
or U17863 (N_17863,N_17488,N_15333);
or U17864 (N_17864,N_17265,N_17248);
and U17865 (N_17865,N_15328,N_15361);
nand U17866 (N_17866,N_15826,N_17083);
and U17867 (N_17867,N_16659,N_16720);
and U17868 (N_17868,N_15118,N_15434);
nand U17869 (N_17869,N_17187,N_15489);
or U17870 (N_17870,N_16082,N_15757);
and U17871 (N_17871,N_16598,N_16119);
and U17872 (N_17872,N_15737,N_15297);
xor U17873 (N_17873,N_15780,N_15720);
and U17874 (N_17874,N_16912,N_16117);
and U17875 (N_17875,N_17097,N_16172);
nand U17876 (N_17876,N_16307,N_15427);
nand U17877 (N_17877,N_17108,N_15022);
xnor U17878 (N_17878,N_17064,N_17281);
xnor U17879 (N_17879,N_16709,N_15635);
nor U17880 (N_17880,N_15061,N_15496);
nand U17881 (N_17881,N_15421,N_16734);
nor U17882 (N_17882,N_15182,N_17191);
and U17883 (N_17883,N_16311,N_17119);
nor U17884 (N_17884,N_15245,N_16204);
or U17885 (N_17885,N_15363,N_15947);
nand U17886 (N_17886,N_15898,N_16790);
nand U17887 (N_17887,N_15075,N_16715);
nor U17888 (N_17888,N_15523,N_16056);
nor U17889 (N_17889,N_15634,N_17081);
nand U17890 (N_17890,N_16697,N_17471);
nand U17891 (N_17891,N_16246,N_15047);
nor U17892 (N_17892,N_15660,N_15220);
and U17893 (N_17893,N_16114,N_16302);
xnor U17894 (N_17894,N_16472,N_16211);
nor U17895 (N_17895,N_16931,N_16021);
xnor U17896 (N_17896,N_15815,N_16146);
or U17897 (N_17897,N_17405,N_17027);
and U17898 (N_17898,N_16257,N_17088);
and U17899 (N_17899,N_16120,N_16595);
nor U17900 (N_17900,N_16183,N_15193);
nand U17901 (N_17901,N_15788,N_17410);
or U17902 (N_17902,N_15196,N_16081);
xnor U17903 (N_17903,N_15778,N_17058);
nor U17904 (N_17904,N_15897,N_17135);
and U17905 (N_17905,N_15289,N_15582);
and U17906 (N_17906,N_16456,N_15773);
or U17907 (N_17907,N_16642,N_15032);
and U17908 (N_17908,N_16639,N_16729);
or U17909 (N_17909,N_16459,N_16018);
or U17910 (N_17910,N_17180,N_15953);
xor U17911 (N_17911,N_16900,N_17092);
xnor U17912 (N_17912,N_15273,N_16005);
nand U17913 (N_17913,N_17011,N_15882);
nor U17914 (N_17914,N_16269,N_15984);
nor U17915 (N_17915,N_15019,N_16420);
or U17916 (N_17916,N_17268,N_17455);
or U17917 (N_17917,N_15064,N_15202);
xnor U17918 (N_17918,N_16394,N_15664);
and U17919 (N_17919,N_16057,N_16239);
nor U17920 (N_17920,N_16254,N_17235);
xnor U17921 (N_17921,N_16806,N_15671);
xor U17922 (N_17922,N_17122,N_15521);
xnor U17923 (N_17923,N_15431,N_15769);
nand U17924 (N_17924,N_17398,N_15284);
or U17925 (N_17925,N_15614,N_17003);
xor U17926 (N_17926,N_16713,N_16875);
xnor U17927 (N_17927,N_17496,N_17228);
and U17928 (N_17928,N_16849,N_15515);
nor U17929 (N_17929,N_16055,N_17164);
nand U17930 (N_17930,N_16710,N_17217);
nand U17931 (N_17931,N_16963,N_15152);
or U17932 (N_17932,N_15507,N_16184);
nor U17933 (N_17933,N_17391,N_16604);
nand U17934 (N_17934,N_16136,N_15699);
nand U17935 (N_17935,N_16554,N_17137);
nand U17936 (N_17936,N_17448,N_17481);
and U17937 (N_17937,N_17037,N_15252);
or U17938 (N_17938,N_15197,N_15622);
or U17939 (N_17939,N_15566,N_15222);
xnor U17940 (N_17940,N_15572,N_15248);
nand U17941 (N_17941,N_17385,N_17215);
nor U17942 (N_17942,N_16127,N_15153);
or U17943 (N_17943,N_17330,N_16611);
and U17944 (N_17944,N_15534,N_15106);
nand U17945 (N_17945,N_16359,N_15960);
nand U17946 (N_17946,N_15726,N_17403);
nand U17947 (N_17947,N_16227,N_16589);
nor U17948 (N_17948,N_15506,N_15650);
or U17949 (N_17949,N_16445,N_16281);
nand U17950 (N_17950,N_15913,N_15267);
xor U17951 (N_17951,N_15129,N_16332);
nand U17952 (N_17952,N_16016,N_16530);
or U17953 (N_17953,N_15631,N_16670);
and U17954 (N_17954,N_15971,N_15755);
xnor U17955 (N_17955,N_17219,N_15470);
or U17956 (N_17956,N_16832,N_16638);
xor U17957 (N_17957,N_16685,N_16584);
nand U17958 (N_17958,N_16245,N_15355);
nor U17959 (N_17959,N_17388,N_16369);
nand U17960 (N_17960,N_15661,N_16429);
xnor U17961 (N_17961,N_17023,N_16837);
or U17962 (N_17962,N_16968,N_15885);
or U17963 (N_17963,N_17371,N_17277);
and U17964 (N_17964,N_16640,N_17321);
nand U17965 (N_17965,N_16510,N_16315);
nand U17966 (N_17966,N_17406,N_16473);
nor U17967 (N_17967,N_16138,N_16262);
and U17968 (N_17968,N_16897,N_15623);
xnor U17969 (N_17969,N_17053,N_16413);
and U17970 (N_17970,N_17435,N_16023);
nor U17971 (N_17971,N_16588,N_16887);
or U17972 (N_17972,N_17188,N_15633);
and U17973 (N_17973,N_15420,N_17367);
nand U17974 (N_17974,N_15397,N_15980);
nand U17975 (N_17975,N_17020,N_15223);
or U17976 (N_17976,N_16457,N_16972);
or U17977 (N_17977,N_16116,N_17113);
and U17978 (N_17978,N_15541,N_16380);
or U17979 (N_17979,N_15447,N_15415);
and U17980 (N_17980,N_17342,N_16153);
nor U17981 (N_17981,N_16527,N_16938);
and U17982 (N_17982,N_15303,N_16434);
and U17983 (N_17983,N_16078,N_16787);
or U17984 (N_17984,N_16085,N_16883);
and U17985 (N_17985,N_15040,N_16015);
nor U17986 (N_17986,N_17255,N_17234);
and U17987 (N_17987,N_16080,N_15348);
nor U17988 (N_17988,N_15513,N_15425);
xnor U17989 (N_17989,N_17174,N_15750);
nor U17990 (N_17990,N_15063,N_16259);
and U17991 (N_17991,N_16831,N_15094);
xor U17992 (N_17992,N_17253,N_17430);
nand U17993 (N_17993,N_16330,N_15001);
xor U17994 (N_17994,N_16641,N_16237);
or U17995 (N_17995,N_15879,N_16980);
or U17996 (N_17996,N_16965,N_16602);
nand U17997 (N_17997,N_16126,N_16044);
or U17998 (N_17998,N_15105,N_17243);
xor U17999 (N_17999,N_16280,N_15461);
and U18000 (N_18000,N_16496,N_16471);
xnor U18001 (N_18001,N_17144,N_15326);
xor U18002 (N_18002,N_15670,N_16020);
xnor U18003 (N_18003,N_15930,N_15862);
nand U18004 (N_18004,N_16971,N_17051);
xnor U18005 (N_18005,N_15454,N_16545);
and U18006 (N_18006,N_15825,N_16877);
or U18007 (N_18007,N_17014,N_16885);
nor U18008 (N_18008,N_15008,N_15684);
xor U18009 (N_18009,N_17364,N_17373);
xnor U18010 (N_18010,N_17043,N_17039);
and U18011 (N_18011,N_17436,N_15209);
or U18012 (N_18012,N_16156,N_17147);
nand U18013 (N_18013,N_15261,N_16030);
and U18014 (N_18014,N_17378,N_15939);
nand U18015 (N_18015,N_16579,N_16309);
or U18016 (N_18016,N_15609,N_17283);
and U18017 (N_18017,N_15230,N_15167);
and U18018 (N_18018,N_16218,N_16578);
nand U18019 (N_18019,N_16801,N_16097);
and U18020 (N_18020,N_16967,N_16189);
and U18021 (N_18021,N_16095,N_15214);
nand U18022 (N_18022,N_17019,N_16414);
and U18023 (N_18023,N_17198,N_15300);
xnor U18024 (N_18024,N_16267,N_16091);
or U18025 (N_18025,N_15777,N_16295);
and U18026 (N_18026,N_15524,N_16341);
nor U18027 (N_18027,N_15310,N_17070);
nand U18028 (N_18028,N_15811,N_15636);
xnor U18029 (N_18029,N_16958,N_15472);
or U18030 (N_18030,N_17212,N_15607);
or U18031 (N_18031,N_16163,N_16822);
and U18032 (N_18032,N_16752,N_15287);
nor U18033 (N_18033,N_16135,N_16861);
or U18034 (N_18034,N_15920,N_15909);
nor U18035 (N_18035,N_17024,N_16424);
nor U18036 (N_18036,N_16901,N_15424);
and U18037 (N_18037,N_15990,N_17360);
nor U18038 (N_18038,N_16810,N_17404);
nand U18039 (N_18039,N_17085,N_16293);
and U18040 (N_18040,N_15618,N_16728);
nand U18041 (N_18041,N_15482,N_15103);
nand U18042 (N_18042,N_15693,N_15231);
or U18043 (N_18043,N_15023,N_15648);
nor U18044 (N_18044,N_16176,N_15192);
xnor U18045 (N_18045,N_17054,N_16573);
or U18046 (N_18046,N_15994,N_17270);
nand U18047 (N_18047,N_16892,N_16990);
nor U18048 (N_18048,N_17299,N_15072);
nor U18049 (N_18049,N_16041,N_17341);
and U18050 (N_18050,N_16792,N_15584);
nor U18051 (N_18051,N_15312,N_15366);
or U18052 (N_18052,N_15959,N_15325);
nand U18053 (N_18053,N_15605,N_15189);
or U18054 (N_18054,N_16730,N_15170);
xnor U18055 (N_18055,N_15134,N_16575);
nand U18056 (N_18056,N_16979,N_15198);
and U18057 (N_18057,N_16466,N_16572);
nor U18058 (N_18058,N_17204,N_17491);
nor U18059 (N_18059,N_16513,N_15792);
nand U18060 (N_18060,N_16873,N_15168);
nand U18061 (N_18061,N_15242,N_16532);
nor U18062 (N_18062,N_15911,N_16804);
and U18063 (N_18063,N_16645,N_15540);
or U18064 (N_18064,N_15210,N_16334);
nor U18065 (N_18065,N_16102,N_17298);
xor U18066 (N_18066,N_17100,N_15797);
and U18067 (N_18067,N_15734,N_17484);
nand U18068 (N_18068,N_15374,N_15013);
or U18069 (N_18069,N_17221,N_15776);
or U18070 (N_18070,N_16318,N_17447);
or U18071 (N_18071,N_15251,N_16273);
or U18072 (N_18072,N_16207,N_16613);
nor U18073 (N_18073,N_16574,N_15697);
nor U18074 (N_18074,N_16616,N_17332);
nand U18075 (N_18075,N_15473,N_17247);
xor U18076 (N_18076,N_16470,N_15178);
and U18077 (N_18077,N_15877,N_15742);
nand U18078 (N_18078,N_15164,N_15277);
xnor U18079 (N_18079,N_15502,N_16698);
and U18080 (N_18080,N_16505,N_16898);
nand U18081 (N_18081,N_16053,N_16260);
or U18082 (N_18082,N_16371,N_17065);
nor U18083 (N_18083,N_17383,N_15663);
nor U18084 (N_18084,N_15850,N_17379);
xnor U18085 (N_18085,N_16828,N_16577);
or U18086 (N_18086,N_15881,N_16175);
xnor U18087 (N_18087,N_16363,N_15853);
and U18088 (N_18088,N_15935,N_15890);
nor U18089 (N_18089,N_15338,N_15360);
xnor U18090 (N_18090,N_16154,N_16462);
nand U18091 (N_18091,N_16063,N_17216);
and U18092 (N_18092,N_16549,N_15038);
and U18093 (N_18093,N_15854,N_15981);
and U18094 (N_18094,N_15493,N_15553);
nand U18095 (N_18095,N_15039,N_15989);
nand U18096 (N_18096,N_17146,N_16742);
and U18097 (N_18097,N_16482,N_17194);
xor U18098 (N_18098,N_16047,N_15621);
nand U18099 (N_18099,N_15795,N_17140);
nand U18100 (N_18100,N_15615,N_16651);
or U18101 (N_18101,N_16465,N_16597);
and U18102 (N_18102,N_15020,N_16463);
nor U18103 (N_18103,N_15883,N_16089);
nor U18104 (N_18104,N_15923,N_16855);
or U18105 (N_18105,N_16760,N_15514);
and U18106 (N_18106,N_16543,N_17344);
nor U18107 (N_18107,N_15938,N_16323);
nor U18108 (N_18108,N_17101,N_16236);
or U18109 (N_18109,N_15336,N_16771);
nor U18110 (N_18110,N_16907,N_16058);
and U18111 (N_18111,N_16406,N_15969);
nand U18112 (N_18112,N_16105,N_17411);
or U18113 (N_18113,N_16708,N_16106);
nor U18114 (N_18114,N_15880,N_17071);
nand U18115 (N_18115,N_17159,N_16283);
and U18116 (N_18116,N_15569,N_17443);
nand U18117 (N_18117,N_16940,N_17182);
and U18118 (N_18118,N_16303,N_15849);
nor U18119 (N_18119,N_16739,N_15373);
xnor U18120 (N_18120,N_15991,N_16608);
xnor U18121 (N_18121,N_16486,N_16763);
nor U18122 (N_18122,N_16266,N_16488);
and U18123 (N_18123,N_15056,N_17485);
nor U18124 (N_18124,N_15599,N_15340);
and U18125 (N_18125,N_16499,N_15078);
nor U18126 (N_18126,N_16233,N_16032);
nor U18127 (N_18127,N_15364,N_15407);
xnor U18128 (N_18128,N_17040,N_17348);
and U18129 (N_18129,N_16439,N_16234);
xor U18130 (N_18130,N_16290,N_17025);
or U18131 (N_18131,N_17236,N_16903);
and U18132 (N_18132,N_16757,N_15087);
and U18133 (N_18133,N_16291,N_15708);
nand U18134 (N_18134,N_15028,N_16727);
and U18135 (N_18135,N_16000,N_16559);
nand U18136 (N_18136,N_15839,N_15546);
xnor U18137 (N_18137,N_17308,N_17161);
xnor U18138 (N_18138,N_15574,N_16476);
and U18139 (N_18139,N_15787,N_15997);
xnor U18140 (N_18140,N_17075,N_16158);
nand U18141 (N_18141,N_16911,N_15116);
or U18142 (N_18142,N_15813,N_16469);
or U18143 (N_18143,N_17326,N_16509);
xor U18144 (N_18144,N_15827,N_15894);
or U18145 (N_18145,N_15525,N_15096);
nand U18146 (N_18146,N_17057,N_15185);
or U18147 (N_18147,N_16817,N_15276);
nand U18148 (N_18148,N_17400,N_16493);
or U18149 (N_18149,N_16489,N_16201);
and U18150 (N_18150,N_16300,N_15786);
nor U18151 (N_18151,N_17426,N_17077);
xor U18152 (N_18152,N_16141,N_16418);
nor U18153 (N_18153,N_15754,N_16690);
xnor U18154 (N_18154,N_17192,N_15383);
nor U18155 (N_18155,N_15906,N_16171);
xnor U18156 (N_18156,N_16338,N_16191);
xnor U18157 (N_18157,N_15201,N_15498);
nor U18158 (N_18158,N_15432,N_16276);
nand U18159 (N_18159,N_16342,N_15550);
xnor U18160 (N_18160,N_15126,N_17155);
or U18161 (N_18161,N_17395,N_15160);
or U18162 (N_18162,N_15024,N_17133);
nand U18163 (N_18163,N_15866,N_16132);
nand U18164 (N_18164,N_17380,N_15368);
or U18165 (N_18165,N_16137,N_16864);
nor U18166 (N_18166,N_16521,N_15119);
nor U18167 (N_18167,N_16838,N_15703);
nand U18168 (N_18168,N_17099,N_15900);
or U18169 (N_18169,N_15120,N_16998);
nor U18170 (N_18170,N_16991,N_17199);
and U18171 (N_18171,N_15396,N_16123);
xnor U18172 (N_18172,N_17238,N_16795);
xnor U18173 (N_18173,N_15331,N_15305);
or U18174 (N_18174,N_16228,N_15044);
and U18175 (N_18175,N_16090,N_16520);
nand U18176 (N_18176,N_17241,N_15114);
nor U18177 (N_18177,N_16764,N_15803);
and U18178 (N_18178,N_15624,N_16930);
xor U18179 (N_18179,N_15484,N_16310);
nand U18180 (N_18180,N_15015,N_15831);
and U18181 (N_18181,N_16383,N_17021);
xor U18182 (N_18182,N_16987,N_16109);
or U18183 (N_18183,N_15704,N_15090);
and U18184 (N_18184,N_16196,N_16270);
nand U18185 (N_18185,N_16165,N_15843);
or U18186 (N_18186,N_15337,N_16039);
nor U18187 (N_18187,N_16389,N_15586);
or U18188 (N_18188,N_17497,N_16658);
nor U18189 (N_18189,N_16797,N_16956);
nand U18190 (N_18190,N_16701,N_16880);
xnor U18191 (N_18191,N_17150,N_15417);
and U18192 (N_18192,N_17334,N_15070);
and U18193 (N_18193,N_16862,N_16774);
or U18194 (N_18194,N_15766,N_15964);
nand U18195 (N_18195,N_15142,N_17267);
or U18196 (N_18196,N_15642,N_15477);
or U18197 (N_18197,N_16289,N_17168);
and U18198 (N_18198,N_17359,N_15683);
and U18199 (N_18199,N_16786,N_15685);
xor U18200 (N_18200,N_16432,N_16159);
nand U18201 (N_18201,N_15207,N_15580);
or U18202 (N_18202,N_16483,N_16596);
xor U18203 (N_18203,N_16524,N_15746);
nor U18204 (N_18204,N_15996,N_16006);
nor U18205 (N_18205,N_17401,N_16072);
nand U18206 (N_18206,N_17331,N_15895);
nor U18207 (N_18207,N_17296,N_16042);
nor U18208 (N_18208,N_17289,N_16384);
or U18209 (N_18209,N_15988,N_15330);
nor U18210 (N_18210,N_15601,N_15492);
and U18211 (N_18211,N_15031,N_17313);
and U18212 (N_18212,N_16546,N_16628);
nand U18213 (N_18213,N_15433,N_17226);
nor U18214 (N_18214,N_16689,N_16190);
or U18215 (N_18215,N_15659,N_15608);
nor U18216 (N_18216,N_16839,N_17419);
or U18217 (N_18217,N_16802,N_16846);
and U18218 (N_18218,N_16871,N_17293);
or U18219 (N_18219,N_15452,N_17151);
and U18220 (N_18220,N_17106,N_16758);
xor U18221 (N_18221,N_17422,N_16947);
and U18222 (N_18222,N_16826,N_15332);
and U18223 (N_18223,N_17029,N_15603);
xor U18224 (N_18224,N_15543,N_16740);
nand U18225 (N_18225,N_16824,N_16783);
xor U18226 (N_18226,N_17449,N_17318);
nand U18227 (N_18227,N_15829,N_17240);
nand U18228 (N_18228,N_15165,N_16235);
nor U18229 (N_18229,N_17176,N_15560);
or U18230 (N_18230,N_16305,N_17458);
xnor U18231 (N_18231,N_17145,N_15927);
nor U18232 (N_18232,N_15695,N_15027);
xor U18233 (N_18233,N_15610,N_15680);
or U18234 (N_18234,N_15833,N_17138);
nand U18235 (N_18235,N_15077,N_17480);
nand U18236 (N_18236,N_15808,N_17263);
or U18237 (N_18237,N_15483,N_16605);
xor U18238 (N_18238,N_16693,N_16650);
nand U18239 (N_18239,N_16104,N_15109);
and U18240 (N_18240,N_17418,N_15375);
nor U18241 (N_18241,N_16791,N_16682);
nand U18242 (N_18242,N_16221,N_17272);
xor U18243 (N_18243,N_15753,N_17254);
xnor U18244 (N_18244,N_16447,N_17375);
nand U18245 (N_18245,N_16160,N_16683);
or U18246 (N_18246,N_15836,N_15740);
nor U18247 (N_18247,N_17434,N_16396);
and U18248 (N_18248,N_16966,N_15288);
and U18249 (N_18249,N_15700,N_17340);
nor U18250 (N_18250,N_15576,N_15439);
and U18251 (N_18251,N_15588,N_15250);
nand U18252 (N_18252,N_15067,N_17218);
and U18253 (N_18253,N_15099,N_17381);
nor U18254 (N_18254,N_15910,N_15359);
or U18255 (N_18255,N_15162,N_15551);
nor U18256 (N_18256,N_15191,N_16876);
xor U18257 (N_18257,N_17018,N_16955);
or U18258 (N_18258,N_17245,N_15914);
and U18259 (N_18259,N_15626,N_15108);
nand U18260 (N_18260,N_16851,N_15349);
and U18261 (N_18261,N_15101,N_16374);
nor U18262 (N_18262,N_17453,N_16847);
nor U18263 (N_18263,N_15822,N_17244);
nand U18264 (N_18264,N_15961,N_16401);
nor U18265 (N_18265,N_16759,N_16522);
nor U18266 (N_18266,N_15509,N_15007);
nand U18267 (N_18267,N_16501,N_15128);
nor U18268 (N_18268,N_16700,N_17178);
nand U18269 (N_18269,N_15619,N_16508);
xnor U18270 (N_18270,N_15974,N_15942);
nor U18271 (N_18271,N_16495,N_16751);
xnor U18272 (N_18272,N_15268,N_15446);
xnor U18273 (N_18273,N_16403,N_16518);
nand U18274 (N_18274,N_15721,N_15963);
nor U18275 (N_18275,N_15309,N_16884);
or U18276 (N_18276,N_15855,N_17120);
xor U18277 (N_18277,N_15125,N_17408);
nand U18278 (N_18278,N_17493,N_15256);
and U18279 (N_18279,N_16814,N_15821);
nor U18280 (N_18280,N_15084,N_16036);
nor U18281 (N_18281,N_16807,N_15595);
and U18282 (N_18282,N_15478,N_15687);
xnor U18283 (N_18283,N_15206,N_16223);
or U18284 (N_18284,N_15799,N_16630);
xor U18285 (N_18285,N_17297,N_15143);
nand U18286 (N_18286,N_16516,N_17225);
nor U18287 (N_18287,N_16362,N_16536);
and U18288 (N_18288,N_16694,N_16271);
xnor U18289 (N_18289,N_17139,N_16609);
nor U18290 (N_18290,N_17132,N_15809);
nand U18291 (N_18291,N_17232,N_16570);
nor U18292 (N_18292,N_15080,N_15290);
nor U18293 (N_18293,N_17413,N_16593);
or U18294 (N_18294,N_15972,N_15085);
or U18295 (N_18295,N_16377,N_15356);
and U18296 (N_18296,N_17372,N_16144);
and U18297 (N_18297,N_15518,N_16202);
and U18298 (N_18298,N_16780,N_15384);
and U18299 (N_18299,N_16544,N_17000);
or U18300 (N_18300,N_17017,N_15638);
xnor U18301 (N_18301,N_15590,N_15581);
nor U18302 (N_18302,N_15208,N_16827);
xnor U18303 (N_18303,N_15321,N_17386);
and U18304 (N_18304,N_15565,N_16594);
or U18305 (N_18305,N_16229,N_15269);
nand U18306 (N_18306,N_16448,N_15253);
xnor U18307 (N_18307,N_16927,N_17170);
nor U18308 (N_18308,N_16067,N_15852);
or U18309 (N_18309,N_16796,N_16390);
nand U18310 (N_18310,N_17220,N_16074);
or U18311 (N_18311,N_15082,N_15967);
xor U18312 (N_18312,N_15698,N_16069);
and U18313 (N_18313,N_15141,N_17498);
or U18314 (N_18314,N_16660,N_15471);
nor U18315 (N_18315,N_16656,N_15998);
nand U18316 (N_18316,N_17472,N_16416);
nand U18317 (N_18317,N_16133,N_17171);
nand U18318 (N_18318,N_15823,N_16327);
or U18319 (N_18319,N_15339,N_17432);
xor U18320 (N_18320,N_15733,N_15500);
nand U18321 (N_18321,N_15035,N_17246);
xnor U18322 (N_18322,N_15302,N_15238);
or U18323 (N_18323,N_16337,N_16084);
and U18324 (N_18324,N_16514,N_17466);
nor U18325 (N_18325,N_15474,N_15344);
or U18326 (N_18326,N_15859,N_15264);
xor U18327 (N_18327,N_15837,N_16013);
or U18328 (N_18328,N_15568,N_15784);
xor U18329 (N_18329,N_15958,N_16874);
and U18330 (N_18330,N_16699,N_16902);
xor U18331 (N_18331,N_15675,N_15136);
nor U18332 (N_18332,N_16215,N_15237);
nand U18333 (N_18333,N_15255,N_17153);
and U18334 (N_18334,N_17105,N_16487);
nor U18335 (N_18335,N_15403,N_16088);
nor U18336 (N_18336,N_16636,N_16093);
and U18337 (N_18337,N_15161,N_16285);
nor U18338 (N_18338,N_15183,N_17402);
nor U18339 (N_18339,N_15458,N_16870);
and U18340 (N_18340,N_17026,N_16648);
nor U18341 (N_18341,N_16244,N_16129);
or U18342 (N_18342,N_15010,N_16569);
nand U18343 (N_18343,N_15810,N_15445);
nand U18344 (N_18344,N_17446,N_15887);
xor U18345 (N_18345,N_17424,N_15722);
nand U18346 (N_18346,N_17125,N_16019);
nor U18347 (N_18347,N_15564,N_16399);
and U18348 (N_18348,N_16274,N_16231);
xnor U18349 (N_18349,N_15391,N_16702);
xnor U18350 (N_18350,N_16193,N_16139);
or U18351 (N_18351,N_15033,N_17368);
nand U18352 (N_18352,N_16743,N_16867);
xnor U18353 (N_18353,N_17087,N_17005);
nand U18354 (N_18354,N_15559,N_15916);
xor U18355 (N_18355,N_16313,N_15041);
or U18356 (N_18356,N_15759,N_16954);
nor U18357 (N_18357,N_15770,N_16022);
nor U18358 (N_18358,N_16284,N_16688);
and U18359 (N_18359,N_15291,N_15455);
nor U18360 (N_18360,N_16468,N_16433);
and U18361 (N_18361,N_16004,N_15095);
or U18362 (N_18362,N_16631,N_15443);
or U18363 (N_18363,N_16412,N_16904);
nand U18364 (N_18364,N_15488,N_15922);
or U18365 (N_18365,N_16925,N_17291);
nand U18366 (N_18366,N_15743,N_16003);
nor U18367 (N_18367,N_16677,N_16264);
and U18368 (N_18368,N_17044,N_15686);
nand U18369 (N_18369,N_16354,N_17475);
or U18370 (N_18370,N_16052,N_15426);
or U18371 (N_18371,N_15257,N_16099);
nand U18372 (N_18372,N_15216,N_15285);
and U18373 (N_18373,N_15647,N_16657);
and U18374 (N_18374,N_15460,N_15928);
nor U18375 (N_18375,N_17110,N_15713);
and U18376 (N_18376,N_15600,N_16358);
and U18377 (N_18377,N_15751,N_16808);
or U18378 (N_18378,N_16555,N_17048);
or U18379 (N_18379,N_17173,N_15593);
and U18380 (N_18380,N_17141,N_16601);
and U18381 (N_18381,N_15156,N_16761);
or U18382 (N_18382,N_16627,N_16732);
and U18383 (N_18383,N_17086,N_15915);
xnor U18384 (N_18384,N_15390,N_16894);
nand U18385 (N_18385,N_16531,N_16845);
nand U18386 (N_18386,N_15334,N_16916);
nor U18387 (N_18387,N_15530,N_15598);
nor U18388 (N_18388,N_16707,N_15783);
and U18389 (N_18389,N_17415,N_16025);
xor U18390 (N_18390,N_16592,N_17251);
or U18391 (N_18391,N_16568,N_16949);
xor U18392 (N_18392,N_15395,N_17412);
nand U18393 (N_18393,N_15807,N_16008);
nand U18394 (N_18394,N_16070,N_15791);
or U18395 (N_18395,N_15315,N_17098);
xnor U18396 (N_18396,N_16366,N_16287);
nand U18397 (N_18397,N_15159,N_15155);
or U18398 (N_18398,N_16750,N_16944);
and U18399 (N_18399,N_16781,N_16722);
xnor U18400 (N_18400,N_15228,N_16475);
nor U18401 (N_18401,N_15794,N_16705);
and U18402 (N_18402,N_17242,N_15098);
xor U18403 (N_18403,N_17041,N_17166);
or U18404 (N_18404,N_17009,N_16112);
nor U18405 (N_18405,N_15878,N_15149);
and U18406 (N_18406,N_16865,N_15709);
or U18407 (N_18407,N_15841,N_16556);
xnor U18408 (N_18408,N_16565,N_16872);
or U18409 (N_18409,N_15485,N_17452);
nand U18410 (N_18410,N_15526,N_15282);
xor U18411 (N_18411,N_15247,N_15548);
nor U18412 (N_18412,N_15819,N_16035);
or U18413 (N_18413,N_15539,N_16714);
xnor U18414 (N_18414,N_16582,N_15123);
nand U18415 (N_18415,N_17361,N_16436);
and U18416 (N_18416,N_16626,N_15365);
or U18417 (N_18417,N_15243,N_15950);
nand U18418 (N_18418,N_17152,N_16200);
or U18419 (N_18419,N_16919,N_15545);
or U18420 (N_18420,N_17022,N_15260);
or U18421 (N_18421,N_17046,N_15679);
xnor U18422 (N_18422,N_15651,N_16378);
nand U18423 (N_18423,N_15940,N_15069);
nor U18424 (N_18424,N_17060,N_16723);
or U18425 (N_18425,N_16633,N_15030);
nand U18426 (N_18426,N_15351,N_16329);
or U18427 (N_18427,N_15205,N_15596);
nand U18428 (N_18428,N_15440,N_17311);
or U18429 (N_18429,N_15423,N_17036);
and U18430 (N_18430,N_16408,N_16077);
and U18431 (N_18431,N_16735,N_17322);
nor U18432 (N_18432,N_16007,N_16982);
and U18433 (N_18433,N_17116,N_16143);
and U18434 (N_18434,N_16644,N_16367);
nor U18435 (N_18435,N_15681,N_16485);
and U18436 (N_18436,N_15575,N_15764);
or U18437 (N_18437,N_15917,N_15912);
and U18438 (N_18438,N_17042,N_16249);
xor U18439 (N_18439,N_16326,N_15163);
xor U18440 (N_18440,N_17056,N_15073);
nand U18441 (N_18441,N_16277,N_17002);
xor U18442 (N_18442,N_15585,N_17354);
nor U18443 (N_18443,N_16419,N_16946);
nand U18444 (N_18444,N_15399,N_16180);
nor U18445 (N_18445,N_16985,N_15174);
or U18446 (N_18446,N_15476,N_16637);
nand U18447 (N_18447,N_16906,N_15137);
nor U18448 (N_18448,N_16625,N_16647);
xor U18449 (N_18449,N_17197,N_16539);
nor U18450 (N_18450,N_16515,N_16765);
or U18451 (N_18451,N_16923,N_15430);
and U18452 (N_18452,N_16107,N_16226);
or U18453 (N_18453,N_16050,N_16373);
nand U18454 (N_18454,N_15217,N_17423);
and U18455 (N_18455,N_15677,N_15796);
nand U18456 (N_18456,N_16376,N_16347);
or U18457 (N_18457,N_17469,N_15817);
nor U18458 (N_18458,N_16212,N_17347);
and U18459 (N_18459,N_17052,N_15789);
nand U18460 (N_18460,N_15613,N_16526);
or U18461 (N_18461,N_15801,N_16599);
nor U18462 (N_18462,N_15844,N_16243);
xnor U18463 (N_18463,N_15501,N_17239);
nand U18464 (N_18464,N_16899,N_15194);
nand U18465 (N_18465,N_15893,N_16263);
or U18466 (N_18466,N_15812,N_16140);
nor U18467 (N_18467,N_16550,N_15583);
and U18468 (N_18468,N_15747,N_16773);
nor U18469 (N_18469,N_15779,N_15973);
xor U18470 (N_18470,N_17200,N_15270);
and U18471 (N_18471,N_17201,N_15188);
xor U18472 (N_18472,N_15176,N_17490);
or U18473 (N_18473,N_16444,N_15557);
and U18474 (N_18474,N_15249,N_16717);
nand U18475 (N_18475,N_17295,N_17104);
and U18476 (N_18476,N_15026,N_17115);
or U18477 (N_18477,N_16478,N_16370);
nor U18478 (N_18478,N_17479,N_16977);
and U18479 (N_18479,N_15016,N_16168);
xor U18480 (N_18480,N_15236,N_15872);
and U18481 (N_18481,N_16772,N_15933);
xnor U18482 (N_18482,N_16661,N_16299);
or U18483 (N_18483,N_15966,N_17275);
and U18484 (N_18484,N_16552,N_16504);
and U18485 (N_18485,N_16009,N_17237);
nand U18486 (N_18486,N_15864,N_16393);
nand U18487 (N_18487,N_16691,N_15000);
nor U18488 (N_18488,N_16962,N_17033);
nor U18489 (N_18489,N_15691,N_16733);
nor U18490 (N_18490,N_15065,N_16142);
and U18491 (N_18491,N_15999,N_16451);
and U18492 (N_18492,N_17069,N_15049);
nand U18493 (N_18493,N_16646,N_15630);
or U18494 (N_18494,N_16065,N_16113);
or U18495 (N_18495,N_17084,N_16209);
or U18496 (N_18496,N_16784,N_17134);
nand U18497 (N_18497,N_16718,N_15342);
or U18498 (N_18498,N_16011,N_15820);
nand U18499 (N_18499,N_15744,N_16997);
xor U18500 (N_18500,N_17425,N_15240);
and U18501 (N_18501,N_15281,N_16696);
xor U18502 (N_18502,N_15177,N_15547);
nor U18503 (N_18503,N_16148,N_16340);
xor U18504 (N_18504,N_16736,N_16519);
nand U18505 (N_18505,N_15259,N_15785);
xnor U18506 (N_18506,N_16960,N_17335);
nand U18507 (N_18507,N_17136,N_17428);
nand U18508 (N_18508,N_16173,N_16409);
and U18509 (N_18509,N_16094,N_15322);
and U18510 (N_18510,N_15617,N_15060);
nand U18511 (N_18511,N_16345,N_16542);
xnor U18512 (N_18512,N_15327,N_17393);
nor U18513 (N_18513,N_16988,N_15017);
nor U18514 (N_18514,N_15148,N_15561);
xor U18515 (N_18515,N_16195,N_15968);
nor U18516 (N_18516,N_16674,N_16452);
nor U18517 (N_18517,N_16978,N_17389);
nor U18518 (N_18518,N_16320,N_17114);
nand U18519 (N_18519,N_17261,N_17131);
and U18520 (N_18520,N_15079,N_16145);
nor U18521 (N_18521,N_15307,N_17093);
and U18522 (N_18522,N_16364,N_16038);
nand U18523 (N_18523,N_15937,N_15411);
xnor U18524 (N_18524,N_16386,N_15147);
nand U18525 (N_18525,N_15046,N_16450);
and U18526 (N_18526,N_17352,N_15578);
and U18527 (N_18527,N_16268,N_16840);
or U18528 (N_18528,N_17049,N_15059);
nand U18529 (N_18529,N_17462,N_17271);
xnor U18530 (N_18530,N_15184,N_16961);
and U18531 (N_18531,N_16048,N_16461);
or U18532 (N_18532,N_16917,N_15014);
or U18533 (N_18533,N_15752,N_15089);
and U18534 (N_18534,N_17482,N_17269);
nor U18535 (N_18535,N_16251,N_17461);
nand U18536 (N_18536,N_16819,N_15279);
and U18537 (N_18537,N_16941,N_16017);
and U18538 (N_18538,N_17343,N_15021);
nand U18539 (N_18539,N_15370,N_15931);
nand U18540 (N_18540,N_15522,N_17195);
and U18541 (N_18541,N_17387,N_15926);
and U18542 (N_18542,N_16279,N_15324);
and U18543 (N_18543,N_15724,N_16936);
xnor U18544 (N_18544,N_16147,N_15891);
nand U18545 (N_18545,N_15896,N_16026);
and U18546 (N_18546,N_16454,N_16240);
xor U18547 (N_18547,N_15696,N_15718);
nand U18548 (N_18548,N_15102,N_15612);
nor U18549 (N_18549,N_16100,N_17128);
nor U18550 (N_18550,N_15625,N_17377);
and U18551 (N_18551,N_15587,N_16391);
nor U18552 (N_18552,N_16800,N_16024);
xor U18553 (N_18553,N_15221,N_16079);
and U18554 (N_18554,N_17211,N_17257);
xor U18555 (N_18555,N_16435,N_16886);
nand U18556 (N_18556,N_17456,N_16059);
nand U18557 (N_18557,N_15730,N_16375);
or U18558 (N_18558,N_17183,N_15003);
nor U18559 (N_18559,N_15036,N_16803);
xor U18560 (N_18560,N_15144,N_16767);
nor U18561 (N_18561,N_15760,N_16788);
xnor U18562 (N_18562,N_17392,N_15173);
xor U18563 (N_18563,N_16811,N_16497);
xor U18564 (N_18564,N_15673,N_17407);
xnor U18565 (N_18565,N_15701,N_16813);
nor U18566 (N_18566,N_16040,N_16869);
and U18567 (N_18567,N_17314,N_17366);
and U18568 (N_18568,N_16957,N_17229);
xnor U18569 (N_18569,N_15556,N_16756);
nor U18570 (N_18570,N_16346,N_16481);
nand U18571 (N_18571,N_16879,N_17303);
nor U18572 (N_18572,N_15892,N_16754);
and U18573 (N_18573,N_17365,N_15562);
nand U18574 (N_18574,N_16186,N_16624);
and U18575 (N_18575,N_16942,N_15781);
and U18576 (N_18576,N_15419,N_16848);
nor U18577 (N_18577,N_17112,N_15860);
and U18578 (N_18578,N_16344,N_16125);
xor U18579 (N_18579,N_17454,N_17376);
nor U18580 (N_18580,N_15818,N_15042);
nor U18581 (N_18581,N_17210,N_17394);
nand U18582 (N_18582,N_17047,N_16169);
or U18583 (N_18583,N_15158,N_15459);
nand U18584 (N_18584,N_16909,N_17207);
nand U18585 (N_18585,N_17494,N_15414);
xnor U18586 (N_18586,N_17476,N_15632);
xor U18587 (N_18587,N_17292,N_16185);
xor U18588 (N_18588,N_17050,N_17382);
and U18589 (N_18589,N_16678,N_15629);
xor U18590 (N_18590,N_17129,N_16422);
nand U18591 (N_18591,N_15793,N_16747);
nor U18592 (N_18592,N_17156,N_16798);
nor U18593 (N_18593,N_17034,N_16238);
xnor U18594 (N_18594,N_15190,N_16164);
nand U18595 (N_18595,N_15592,N_15376);
or U18596 (N_18596,N_15899,N_15563);
and U18597 (N_18597,N_15627,N_16561);
nor U18598 (N_18598,N_15225,N_16915);
xnor U18599 (N_18599,N_15665,N_15976);
and U18600 (N_18600,N_15508,N_15579);
or U18601 (N_18601,N_16121,N_15381);
nand U18602 (N_18602,N_15856,N_15640);
xnor U18603 (N_18603,N_17345,N_17286);
xnor U18604 (N_18604,N_15903,N_15406);
nor U18605 (N_18605,N_17279,N_15798);
nand U18606 (N_18606,N_15688,N_16010);
xor U18607 (N_18607,N_15343,N_15051);
and U18608 (N_18608,N_16540,N_15308);
nor U18609 (N_18609,N_16721,N_17117);
xnor U18610 (N_18610,N_17006,N_15516);
nor U18611 (N_18611,N_16253,N_16835);
and U18612 (N_18612,N_17072,N_15706);
or U18613 (N_18613,N_16768,N_17203);
nand U18614 (N_18614,N_15529,N_15503);
xnor U18615 (N_18615,N_16449,N_16970);
xnor U18616 (N_18616,N_15475,N_15886);
and U18617 (N_18617,N_16704,N_16686);
nand U18618 (N_18618,N_16162,N_16744);
xor U18619 (N_18619,N_16973,N_17465);
and U18620 (N_18620,N_15254,N_16134);
or U18621 (N_18621,N_16108,N_15771);
and U18622 (N_18622,N_17013,N_16719);
xor U18623 (N_18623,N_15672,N_15335);
nand U18624 (N_18624,N_17256,N_15745);
nand U18625 (N_18625,N_15824,N_16068);
xnor U18626 (N_18626,N_15690,N_16455);
or U18627 (N_18627,N_16214,N_17158);
nand U18628 (N_18628,N_17309,N_15846);
nor U18629 (N_18629,N_15616,N_15662);
or U18630 (N_18630,N_15655,N_16620);
and U18631 (N_18631,N_15888,N_17316);
or U18632 (N_18632,N_17433,N_16506);
xnor U18633 (N_18633,N_17258,N_17284);
xnor U18634 (N_18634,N_16111,N_15802);
xnor U18635 (N_18635,N_17300,N_16178);
xor U18636 (N_18636,N_16216,N_16336);
xnor U18637 (N_18637,N_16061,N_15728);
or U18638 (N_18638,N_16948,N_15179);
nand U18639 (N_18639,N_15494,N_15367);
or U18640 (N_18640,N_16725,N_15649);
nor U18641 (N_18641,N_16130,N_16312);
nand U18642 (N_18642,N_15418,N_15379);
and U18643 (N_18643,N_16896,N_17351);
xnor U18644 (N_18644,N_15921,N_15669);
or U18645 (N_18645,N_15346,N_16392);
and U18646 (N_18646,N_16012,N_17169);
xor U18647 (N_18647,N_16206,N_16453);
or U18648 (N_18648,N_15387,N_15239);
nor U18649 (N_18649,N_16395,N_16247);
nor U18650 (N_18650,N_17362,N_17095);
nand U18651 (N_18651,N_16607,N_15727);
xnor U18652 (N_18652,N_15241,N_16586);
nor U18653 (N_18653,N_15774,N_15117);
xnor U18654 (N_18654,N_17004,N_15211);
and U18655 (N_18655,N_16064,N_16428);
and U18656 (N_18656,N_16192,N_17329);
nand U18657 (N_18657,N_17273,N_15729);
or U18658 (N_18658,N_15951,N_16073);
and U18659 (N_18659,N_17287,N_17118);
xor U18660 (N_18660,N_16676,N_15714);
nand U18661 (N_18661,N_15402,N_16653);
xnor U18662 (N_18662,N_16560,N_15392);
xnor U18663 (N_18663,N_16492,N_15029);
xnor U18664 (N_18664,N_16321,N_15945);
and U18665 (N_18665,N_15295,N_16417);
xnor U18666 (N_18666,N_15936,N_17260);
nand U18667 (N_18667,N_15570,N_16232);
xnor U18668 (N_18668,N_16151,N_16381);
and U18669 (N_18669,N_15924,N_16538);
nor U18670 (N_18670,N_16857,N_17123);
or U18671 (N_18671,N_15591,N_16205);
or U18672 (N_18672,N_16799,N_15869);
nand U18673 (N_18673,N_15462,N_15995);
nand U18674 (N_18674,N_15865,N_16198);
and U18675 (N_18675,N_15009,N_17285);
nand U18676 (N_18676,N_15666,N_15549);
and U18677 (N_18677,N_17333,N_15054);
and U18678 (N_18678,N_15805,N_17266);
and U18679 (N_18679,N_16860,N_16440);
nor U18680 (N_18680,N_15408,N_15977);
nand U18681 (N_18681,N_17477,N_17369);
nor U18682 (N_18682,N_15380,N_15329);
and U18683 (N_18683,N_17429,N_15444);
or U18684 (N_18684,N_16155,N_15135);
nand U18685 (N_18685,N_16576,N_17440);
xnor U18686 (N_18686,N_16600,N_15121);
and U18687 (N_18687,N_15058,N_17185);
nor U18688 (N_18688,N_17317,N_16843);
nor U18689 (N_18689,N_16437,N_15362);
nor U18690 (N_18690,N_15313,N_15761);
or U18691 (N_18691,N_16402,N_16387);
and U18692 (N_18692,N_16149,N_15314);
nand U18693 (N_18693,N_16629,N_15979);
or U18694 (N_18694,N_16924,N_15511);
or U18695 (N_18695,N_15838,N_17102);
nand U18696 (N_18696,N_17339,N_15571);
xnor U18697 (N_18697,N_17305,N_16324);
or U18698 (N_18698,N_15130,N_15468);
or U18699 (N_18699,N_16294,N_16124);
xnor U18700 (N_18700,N_15535,N_16953);
xor U18701 (N_18701,N_15946,N_15611);
or U18702 (N_18702,N_15092,N_16562);
and U18703 (N_18703,N_16423,N_15832);
nand U18704 (N_18704,N_16076,N_16945);
nand U18705 (N_18705,N_17325,N_17224);
xor U18706 (N_18706,N_15602,N_16755);
nand U18707 (N_18707,N_17437,N_16523);
or U18708 (N_18708,N_16500,N_15711);
and U18709 (N_18709,N_15907,N_16430);
and U18710 (N_18710,N_15171,N_15505);
nor U18711 (N_18711,N_16868,N_16255);
or U18712 (N_18712,N_16854,N_15275);
or U18713 (N_18713,N_16603,N_16749);
xnor U18714 (N_18714,N_15919,N_15385);
nand U18715 (N_18715,N_16669,N_15053);
nand U18716 (N_18716,N_15905,N_15457);
nand U18717 (N_18717,N_15487,N_17304);
xor U18718 (N_18718,N_16410,N_15517);
nor U18719 (N_18719,N_16775,N_17390);
and U18720 (N_18720,N_16687,N_16314);
nor U18721 (N_18721,N_15127,N_17059);
or U18722 (N_18722,N_16355,N_16372);
or U18723 (N_18723,N_16385,N_15181);
or U18724 (N_18724,N_15111,N_15071);
nor U18725 (N_18725,N_16071,N_17409);
nor U18726 (N_18726,N_15654,N_16950);
or U18727 (N_18727,N_17280,N_15597);
xor U18728 (N_18728,N_16225,N_17487);
nand U18729 (N_18729,N_17109,N_17186);
or U18730 (N_18730,N_15978,N_15965);
and U18731 (N_18731,N_16525,N_15732);
or U18732 (N_18732,N_15413,N_16037);
and U18733 (N_18733,N_15544,N_16528);
nor U18734 (N_18734,N_17441,N_15347);
or U18735 (N_18735,N_15848,N_16256);
nor U18736 (N_18736,N_16934,N_15437);
xor U18737 (N_18737,N_15589,N_15876);
and U18738 (N_18738,N_16317,N_16852);
or U18739 (N_18739,N_16976,N_16591);
and U18740 (N_18740,N_15932,N_16087);
or U18741 (N_18741,N_17315,N_16606);
or U18742 (N_18742,N_17080,N_16241);
and U18743 (N_18743,N_15863,N_16571);
or U18744 (N_18744,N_16502,N_16407);
xor U18745 (N_18745,N_17142,N_15412);
nor U18746 (N_18746,N_15944,N_17356);
nand U18747 (N_18747,N_16152,N_16278);
nand U18748 (N_18748,N_15639,N_16610);
xnor U18749 (N_18749,N_17336,N_15200);
or U18750 (N_18750,N_15795,N_16814);
nor U18751 (N_18751,N_15980,N_16619);
nand U18752 (N_18752,N_16437,N_15784);
and U18753 (N_18753,N_16937,N_16384);
and U18754 (N_18754,N_16563,N_15424);
nor U18755 (N_18755,N_16365,N_15780);
xor U18756 (N_18756,N_15439,N_16142);
nand U18757 (N_18757,N_16360,N_16895);
nor U18758 (N_18758,N_15509,N_15120);
xor U18759 (N_18759,N_15196,N_15847);
and U18760 (N_18760,N_16798,N_15711);
xor U18761 (N_18761,N_16017,N_15221);
nand U18762 (N_18762,N_16082,N_17063);
or U18763 (N_18763,N_15968,N_17439);
nor U18764 (N_18764,N_16050,N_16627);
nor U18765 (N_18765,N_15464,N_16879);
or U18766 (N_18766,N_17349,N_15142);
nand U18767 (N_18767,N_15306,N_17160);
and U18768 (N_18768,N_15649,N_15689);
nand U18769 (N_18769,N_15991,N_16569);
or U18770 (N_18770,N_16280,N_17327);
nand U18771 (N_18771,N_16940,N_15963);
and U18772 (N_18772,N_16566,N_15397);
or U18773 (N_18773,N_15828,N_16740);
nor U18774 (N_18774,N_17167,N_17027);
or U18775 (N_18775,N_17143,N_15346);
xnor U18776 (N_18776,N_16479,N_16239);
nand U18777 (N_18777,N_16439,N_15963);
nor U18778 (N_18778,N_16370,N_16447);
and U18779 (N_18779,N_15533,N_16183);
or U18780 (N_18780,N_16402,N_17288);
xnor U18781 (N_18781,N_15195,N_16952);
nor U18782 (N_18782,N_15729,N_16792);
xor U18783 (N_18783,N_16989,N_16681);
xnor U18784 (N_18784,N_17016,N_16327);
or U18785 (N_18785,N_17440,N_15049);
nor U18786 (N_18786,N_16434,N_15279);
and U18787 (N_18787,N_15015,N_15982);
and U18788 (N_18788,N_16935,N_17065);
and U18789 (N_18789,N_16055,N_15930);
xor U18790 (N_18790,N_15970,N_15081);
xor U18791 (N_18791,N_16322,N_17038);
and U18792 (N_18792,N_16050,N_16433);
nor U18793 (N_18793,N_15927,N_16834);
nand U18794 (N_18794,N_15991,N_16361);
nand U18795 (N_18795,N_16619,N_17149);
nor U18796 (N_18796,N_16108,N_15151);
or U18797 (N_18797,N_16666,N_16134);
nor U18798 (N_18798,N_15650,N_16181);
xor U18799 (N_18799,N_17323,N_16475);
and U18800 (N_18800,N_17328,N_15043);
or U18801 (N_18801,N_17494,N_17164);
xnor U18802 (N_18802,N_17126,N_16081);
or U18803 (N_18803,N_16260,N_15961);
xnor U18804 (N_18804,N_16531,N_15358);
nor U18805 (N_18805,N_17139,N_16969);
xor U18806 (N_18806,N_15589,N_16271);
xnor U18807 (N_18807,N_16556,N_16970);
and U18808 (N_18808,N_15368,N_15024);
and U18809 (N_18809,N_15437,N_16991);
and U18810 (N_18810,N_16236,N_15283);
xnor U18811 (N_18811,N_16511,N_17478);
nand U18812 (N_18812,N_16624,N_15775);
or U18813 (N_18813,N_15503,N_16675);
and U18814 (N_18814,N_17075,N_16840);
or U18815 (N_18815,N_15260,N_16065);
nand U18816 (N_18816,N_15458,N_17258);
xnor U18817 (N_18817,N_16538,N_17168);
nor U18818 (N_18818,N_17409,N_16916);
or U18819 (N_18819,N_15386,N_15463);
xnor U18820 (N_18820,N_17013,N_16530);
or U18821 (N_18821,N_15683,N_15691);
xor U18822 (N_18822,N_17390,N_16077);
nand U18823 (N_18823,N_15270,N_17249);
nor U18824 (N_18824,N_16551,N_16140);
xnor U18825 (N_18825,N_16390,N_15313);
nor U18826 (N_18826,N_16220,N_16537);
or U18827 (N_18827,N_15295,N_16024);
nor U18828 (N_18828,N_15062,N_16523);
nand U18829 (N_18829,N_15303,N_15588);
and U18830 (N_18830,N_15798,N_16377);
xor U18831 (N_18831,N_15251,N_16028);
nor U18832 (N_18832,N_16773,N_15904);
xnor U18833 (N_18833,N_16765,N_16821);
nand U18834 (N_18834,N_16996,N_15550);
xor U18835 (N_18835,N_16372,N_15931);
nor U18836 (N_18836,N_15896,N_17151);
and U18837 (N_18837,N_16833,N_15090);
nand U18838 (N_18838,N_16733,N_15217);
xnor U18839 (N_18839,N_15166,N_16562);
or U18840 (N_18840,N_15774,N_17219);
or U18841 (N_18841,N_16544,N_15979);
or U18842 (N_18842,N_15818,N_16499);
xor U18843 (N_18843,N_15716,N_15327);
xnor U18844 (N_18844,N_16962,N_17333);
nand U18845 (N_18845,N_15195,N_17499);
nor U18846 (N_18846,N_16655,N_16268);
or U18847 (N_18847,N_15094,N_15723);
nand U18848 (N_18848,N_15015,N_17136);
or U18849 (N_18849,N_17225,N_16163);
or U18850 (N_18850,N_17121,N_15333);
xnor U18851 (N_18851,N_16045,N_17497);
xor U18852 (N_18852,N_16703,N_15941);
nor U18853 (N_18853,N_16532,N_16260);
nand U18854 (N_18854,N_17136,N_16475);
nand U18855 (N_18855,N_15818,N_15088);
and U18856 (N_18856,N_17108,N_15697);
or U18857 (N_18857,N_17364,N_15118);
and U18858 (N_18858,N_17074,N_17435);
nand U18859 (N_18859,N_15074,N_16773);
or U18860 (N_18860,N_15234,N_16133);
xor U18861 (N_18861,N_17185,N_17224);
nor U18862 (N_18862,N_15811,N_15628);
and U18863 (N_18863,N_15506,N_16524);
or U18864 (N_18864,N_16837,N_17177);
and U18865 (N_18865,N_16167,N_15274);
or U18866 (N_18866,N_16217,N_16340);
xor U18867 (N_18867,N_15358,N_17438);
xor U18868 (N_18868,N_15411,N_16638);
or U18869 (N_18869,N_17079,N_16197);
nand U18870 (N_18870,N_16748,N_17129);
xor U18871 (N_18871,N_16304,N_16497);
and U18872 (N_18872,N_15094,N_16644);
xnor U18873 (N_18873,N_16529,N_15457);
and U18874 (N_18874,N_15551,N_17153);
xnor U18875 (N_18875,N_16684,N_15207);
xor U18876 (N_18876,N_16075,N_15559);
nand U18877 (N_18877,N_16205,N_17430);
nor U18878 (N_18878,N_15603,N_15820);
and U18879 (N_18879,N_16612,N_16917);
nand U18880 (N_18880,N_17264,N_15864);
xnor U18881 (N_18881,N_16020,N_16945);
xnor U18882 (N_18882,N_15011,N_17336);
nor U18883 (N_18883,N_15154,N_15404);
or U18884 (N_18884,N_16825,N_15024);
and U18885 (N_18885,N_16992,N_17382);
or U18886 (N_18886,N_15711,N_16025);
nor U18887 (N_18887,N_15785,N_16991);
nor U18888 (N_18888,N_16721,N_15596);
and U18889 (N_18889,N_15846,N_16893);
nand U18890 (N_18890,N_16457,N_15394);
and U18891 (N_18891,N_15289,N_16252);
and U18892 (N_18892,N_16092,N_15110);
nand U18893 (N_18893,N_16905,N_15820);
and U18894 (N_18894,N_15115,N_17389);
or U18895 (N_18895,N_15740,N_16747);
nor U18896 (N_18896,N_17367,N_15237);
xor U18897 (N_18897,N_17479,N_15224);
xnor U18898 (N_18898,N_16189,N_17296);
xor U18899 (N_18899,N_16895,N_17463);
nand U18900 (N_18900,N_16852,N_15258);
nand U18901 (N_18901,N_16897,N_15831);
xnor U18902 (N_18902,N_17225,N_15965);
nand U18903 (N_18903,N_16338,N_15221);
nor U18904 (N_18904,N_16582,N_15422);
or U18905 (N_18905,N_17379,N_17215);
or U18906 (N_18906,N_16739,N_15896);
and U18907 (N_18907,N_16212,N_17320);
nor U18908 (N_18908,N_16845,N_15779);
nand U18909 (N_18909,N_16963,N_16121);
xor U18910 (N_18910,N_15725,N_16233);
and U18911 (N_18911,N_17406,N_15418);
and U18912 (N_18912,N_15152,N_16343);
nand U18913 (N_18913,N_15467,N_16779);
xor U18914 (N_18914,N_16965,N_16281);
and U18915 (N_18915,N_15924,N_17295);
nand U18916 (N_18916,N_16252,N_16981);
nor U18917 (N_18917,N_16582,N_15710);
nor U18918 (N_18918,N_15173,N_15278);
xnor U18919 (N_18919,N_16306,N_17021);
xor U18920 (N_18920,N_17329,N_16323);
xnor U18921 (N_18921,N_16176,N_15660);
nor U18922 (N_18922,N_17351,N_16399);
nor U18923 (N_18923,N_16327,N_16191);
or U18924 (N_18924,N_16299,N_16448);
or U18925 (N_18925,N_17411,N_15858);
nor U18926 (N_18926,N_16341,N_17082);
and U18927 (N_18927,N_16529,N_17287);
nand U18928 (N_18928,N_16994,N_15425);
or U18929 (N_18929,N_17371,N_15025);
xor U18930 (N_18930,N_16542,N_16569);
or U18931 (N_18931,N_15209,N_15015);
or U18932 (N_18932,N_17015,N_16925);
nand U18933 (N_18933,N_15037,N_15030);
nor U18934 (N_18934,N_16815,N_17429);
xor U18935 (N_18935,N_15677,N_16340);
xor U18936 (N_18936,N_16763,N_15260);
or U18937 (N_18937,N_15929,N_16371);
nand U18938 (N_18938,N_15109,N_15281);
nand U18939 (N_18939,N_16835,N_16627);
nand U18940 (N_18940,N_15597,N_17385);
xor U18941 (N_18941,N_15474,N_17402);
nand U18942 (N_18942,N_15148,N_15769);
nand U18943 (N_18943,N_15088,N_16997);
xor U18944 (N_18944,N_16030,N_16703);
xor U18945 (N_18945,N_15741,N_16392);
or U18946 (N_18946,N_15663,N_15692);
xnor U18947 (N_18947,N_15098,N_16938);
and U18948 (N_18948,N_15961,N_15988);
nand U18949 (N_18949,N_15866,N_15999);
and U18950 (N_18950,N_15286,N_15216);
nor U18951 (N_18951,N_15053,N_16725);
nand U18952 (N_18952,N_17361,N_15665);
or U18953 (N_18953,N_16457,N_15469);
nand U18954 (N_18954,N_16073,N_16769);
and U18955 (N_18955,N_16538,N_15025);
nor U18956 (N_18956,N_16550,N_17227);
nor U18957 (N_18957,N_15791,N_16024);
and U18958 (N_18958,N_16762,N_16519);
xor U18959 (N_18959,N_16193,N_16270);
nor U18960 (N_18960,N_16883,N_17238);
and U18961 (N_18961,N_15954,N_16352);
nor U18962 (N_18962,N_15117,N_16413);
nor U18963 (N_18963,N_16373,N_15621);
or U18964 (N_18964,N_16601,N_15885);
xnor U18965 (N_18965,N_15005,N_16818);
or U18966 (N_18966,N_15397,N_15454);
nand U18967 (N_18967,N_16045,N_15036);
xor U18968 (N_18968,N_15883,N_16500);
and U18969 (N_18969,N_16210,N_15012);
nand U18970 (N_18970,N_17454,N_15208);
nand U18971 (N_18971,N_16091,N_17062);
xnor U18972 (N_18972,N_15224,N_16443);
and U18973 (N_18973,N_17378,N_17309);
nand U18974 (N_18974,N_15185,N_16742);
or U18975 (N_18975,N_15291,N_16845);
nand U18976 (N_18976,N_17460,N_16394);
nor U18977 (N_18977,N_16028,N_17447);
and U18978 (N_18978,N_15002,N_16188);
or U18979 (N_18979,N_16991,N_16893);
nand U18980 (N_18980,N_17314,N_15488);
nor U18981 (N_18981,N_16461,N_16695);
or U18982 (N_18982,N_16434,N_15509);
nand U18983 (N_18983,N_15713,N_17068);
nor U18984 (N_18984,N_16339,N_16939);
xor U18985 (N_18985,N_17189,N_15823);
nand U18986 (N_18986,N_15076,N_17325);
nor U18987 (N_18987,N_15924,N_15075);
or U18988 (N_18988,N_16139,N_15779);
or U18989 (N_18989,N_15685,N_16148);
and U18990 (N_18990,N_16502,N_17497);
nor U18991 (N_18991,N_16926,N_15638);
nor U18992 (N_18992,N_15291,N_15293);
xnor U18993 (N_18993,N_17262,N_16125);
and U18994 (N_18994,N_15562,N_16229);
nand U18995 (N_18995,N_15300,N_16765);
xnor U18996 (N_18996,N_17391,N_15824);
nand U18997 (N_18997,N_17459,N_16490);
and U18998 (N_18998,N_17460,N_15191);
xor U18999 (N_18999,N_16094,N_16533);
nor U19000 (N_19000,N_15474,N_15460);
nor U19001 (N_19001,N_16021,N_17065);
and U19002 (N_19002,N_16573,N_17087);
and U19003 (N_19003,N_15379,N_16882);
or U19004 (N_19004,N_15399,N_16490);
nand U19005 (N_19005,N_16211,N_15322);
or U19006 (N_19006,N_17386,N_16684);
nor U19007 (N_19007,N_16776,N_17404);
nor U19008 (N_19008,N_15353,N_17225);
and U19009 (N_19009,N_17225,N_17377);
or U19010 (N_19010,N_17218,N_15595);
and U19011 (N_19011,N_16858,N_16616);
and U19012 (N_19012,N_15020,N_15763);
and U19013 (N_19013,N_15418,N_16094);
and U19014 (N_19014,N_15858,N_15346);
or U19015 (N_19015,N_15873,N_15101);
and U19016 (N_19016,N_16531,N_16252);
xor U19017 (N_19017,N_15789,N_16520);
or U19018 (N_19018,N_15315,N_17328);
and U19019 (N_19019,N_15374,N_16829);
xor U19020 (N_19020,N_15275,N_17262);
nor U19021 (N_19021,N_15173,N_16753);
xnor U19022 (N_19022,N_17349,N_15374);
nand U19023 (N_19023,N_17448,N_15322);
and U19024 (N_19024,N_17289,N_15182);
and U19025 (N_19025,N_17223,N_16274);
xor U19026 (N_19026,N_17206,N_16006);
xnor U19027 (N_19027,N_16226,N_15990);
and U19028 (N_19028,N_17144,N_15401);
nor U19029 (N_19029,N_17273,N_17386);
or U19030 (N_19030,N_17092,N_15380);
or U19031 (N_19031,N_15210,N_16117);
nand U19032 (N_19032,N_16452,N_17188);
nor U19033 (N_19033,N_15642,N_15486);
and U19034 (N_19034,N_15584,N_17369);
nor U19035 (N_19035,N_17403,N_17124);
xor U19036 (N_19036,N_15328,N_17091);
nand U19037 (N_19037,N_17385,N_15016);
and U19038 (N_19038,N_16417,N_16227);
or U19039 (N_19039,N_16130,N_16637);
and U19040 (N_19040,N_16709,N_15704);
xnor U19041 (N_19041,N_16563,N_17044);
xnor U19042 (N_19042,N_16855,N_17018);
or U19043 (N_19043,N_15907,N_16277);
xor U19044 (N_19044,N_17486,N_16648);
xor U19045 (N_19045,N_15036,N_16325);
xor U19046 (N_19046,N_16691,N_16706);
xnor U19047 (N_19047,N_16377,N_16796);
nor U19048 (N_19048,N_15198,N_17069);
xnor U19049 (N_19049,N_17022,N_15435);
and U19050 (N_19050,N_16951,N_15087);
nor U19051 (N_19051,N_17236,N_16185);
nand U19052 (N_19052,N_15630,N_15170);
xor U19053 (N_19053,N_15038,N_16744);
and U19054 (N_19054,N_16089,N_15406);
xor U19055 (N_19055,N_15289,N_17164);
nand U19056 (N_19056,N_15740,N_16947);
or U19057 (N_19057,N_17479,N_17344);
or U19058 (N_19058,N_16994,N_16966);
or U19059 (N_19059,N_15972,N_16390);
or U19060 (N_19060,N_16924,N_16433);
or U19061 (N_19061,N_15515,N_15418);
nor U19062 (N_19062,N_17406,N_16279);
and U19063 (N_19063,N_16031,N_15190);
xnor U19064 (N_19064,N_16642,N_15172);
nor U19065 (N_19065,N_15920,N_15596);
and U19066 (N_19066,N_16938,N_15227);
nor U19067 (N_19067,N_16575,N_16908);
and U19068 (N_19068,N_15969,N_15583);
xor U19069 (N_19069,N_16205,N_16504);
or U19070 (N_19070,N_15805,N_17434);
nand U19071 (N_19071,N_16509,N_15358);
xor U19072 (N_19072,N_15766,N_16769);
nor U19073 (N_19073,N_17327,N_15237);
nand U19074 (N_19074,N_17352,N_15597);
xnor U19075 (N_19075,N_17220,N_17240);
and U19076 (N_19076,N_16228,N_15574);
and U19077 (N_19077,N_16692,N_15414);
and U19078 (N_19078,N_16243,N_15869);
or U19079 (N_19079,N_17385,N_17191);
xnor U19080 (N_19080,N_16169,N_15787);
nor U19081 (N_19081,N_15843,N_16477);
or U19082 (N_19082,N_16280,N_15724);
xnor U19083 (N_19083,N_16065,N_15288);
xor U19084 (N_19084,N_16488,N_16993);
and U19085 (N_19085,N_16034,N_16711);
and U19086 (N_19086,N_17060,N_16560);
and U19087 (N_19087,N_15445,N_15062);
nor U19088 (N_19088,N_15774,N_16513);
nor U19089 (N_19089,N_15946,N_16441);
or U19090 (N_19090,N_15168,N_15440);
nand U19091 (N_19091,N_16123,N_16828);
and U19092 (N_19092,N_16651,N_15543);
xnor U19093 (N_19093,N_15471,N_17179);
xor U19094 (N_19094,N_17497,N_15015);
nor U19095 (N_19095,N_15083,N_15844);
nand U19096 (N_19096,N_15674,N_16902);
or U19097 (N_19097,N_15307,N_15842);
nor U19098 (N_19098,N_15214,N_16113);
nor U19099 (N_19099,N_15951,N_16669);
or U19100 (N_19100,N_16965,N_15636);
or U19101 (N_19101,N_15583,N_16029);
nor U19102 (N_19102,N_16626,N_17377);
xor U19103 (N_19103,N_16410,N_16371);
nand U19104 (N_19104,N_16258,N_17459);
and U19105 (N_19105,N_15923,N_16270);
nand U19106 (N_19106,N_16553,N_16727);
xor U19107 (N_19107,N_15494,N_16432);
nand U19108 (N_19108,N_15585,N_16327);
nor U19109 (N_19109,N_15290,N_16124);
nand U19110 (N_19110,N_16486,N_15961);
nand U19111 (N_19111,N_15608,N_16193);
nand U19112 (N_19112,N_15880,N_15611);
nand U19113 (N_19113,N_15201,N_17100);
and U19114 (N_19114,N_15162,N_15076);
or U19115 (N_19115,N_17212,N_15150);
nand U19116 (N_19116,N_16736,N_15814);
xnor U19117 (N_19117,N_15599,N_15361);
xor U19118 (N_19118,N_16496,N_16939);
nor U19119 (N_19119,N_16311,N_16897);
xnor U19120 (N_19120,N_15591,N_15683);
xnor U19121 (N_19121,N_16025,N_15867);
nand U19122 (N_19122,N_15088,N_15471);
xnor U19123 (N_19123,N_17016,N_15516);
or U19124 (N_19124,N_17159,N_17060);
nand U19125 (N_19125,N_17147,N_15084);
xnor U19126 (N_19126,N_16067,N_15716);
or U19127 (N_19127,N_15390,N_16867);
xnor U19128 (N_19128,N_15787,N_16003);
or U19129 (N_19129,N_16137,N_17026);
xnor U19130 (N_19130,N_16979,N_15960);
nor U19131 (N_19131,N_15319,N_16429);
and U19132 (N_19132,N_17177,N_16141);
nor U19133 (N_19133,N_15432,N_16093);
xor U19134 (N_19134,N_16634,N_16538);
xnor U19135 (N_19135,N_16730,N_16283);
and U19136 (N_19136,N_16168,N_16293);
or U19137 (N_19137,N_16615,N_15731);
or U19138 (N_19138,N_15913,N_16341);
xnor U19139 (N_19139,N_15318,N_16784);
and U19140 (N_19140,N_16602,N_17488);
and U19141 (N_19141,N_17348,N_15440);
and U19142 (N_19142,N_16759,N_16995);
nor U19143 (N_19143,N_15826,N_16314);
nor U19144 (N_19144,N_16304,N_15389);
or U19145 (N_19145,N_16678,N_17195);
nor U19146 (N_19146,N_16665,N_16561);
nor U19147 (N_19147,N_15157,N_16111);
or U19148 (N_19148,N_15139,N_17418);
or U19149 (N_19149,N_16911,N_16090);
nand U19150 (N_19150,N_16289,N_16477);
or U19151 (N_19151,N_15370,N_16905);
nand U19152 (N_19152,N_16416,N_15375);
or U19153 (N_19153,N_16212,N_15873);
xnor U19154 (N_19154,N_16758,N_15028);
and U19155 (N_19155,N_17154,N_15351);
and U19156 (N_19156,N_15031,N_15341);
and U19157 (N_19157,N_15839,N_15232);
or U19158 (N_19158,N_15785,N_17302);
xnor U19159 (N_19159,N_15785,N_16096);
xor U19160 (N_19160,N_15199,N_17411);
nand U19161 (N_19161,N_15489,N_16267);
and U19162 (N_19162,N_16972,N_16724);
and U19163 (N_19163,N_15041,N_15812);
nor U19164 (N_19164,N_15230,N_15683);
nor U19165 (N_19165,N_15492,N_16331);
and U19166 (N_19166,N_17130,N_16058);
xnor U19167 (N_19167,N_17411,N_16641);
xnor U19168 (N_19168,N_16169,N_15252);
nand U19169 (N_19169,N_15945,N_16033);
xor U19170 (N_19170,N_15787,N_15854);
or U19171 (N_19171,N_15313,N_15447);
xnor U19172 (N_19172,N_15751,N_15362);
xnor U19173 (N_19173,N_17053,N_16754);
nand U19174 (N_19174,N_15273,N_15670);
or U19175 (N_19175,N_15721,N_16224);
xor U19176 (N_19176,N_16143,N_15797);
nand U19177 (N_19177,N_17199,N_17460);
nor U19178 (N_19178,N_17441,N_17207);
or U19179 (N_19179,N_16607,N_16569);
and U19180 (N_19180,N_17181,N_15982);
nand U19181 (N_19181,N_17034,N_16925);
and U19182 (N_19182,N_16941,N_15453);
nand U19183 (N_19183,N_15217,N_16969);
nor U19184 (N_19184,N_15199,N_16875);
and U19185 (N_19185,N_16333,N_16665);
nor U19186 (N_19186,N_16794,N_15941);
nor U19187 (N_19187,N_15756,N_15589);
xnor U19188 (N_19188,N_15640,N_17010);
nand U19189 (N_19189,N_16889,N_15127);
and U19190 (N_19190,N_15479,N_17001);
nor U19191 (N_19191,N_16487,N_16247);
nand U19192 (N_19192,N_17463,N_16015);
nor U19193 (N_19193,N_15643,N_15492);
and U19194 (N_19194,N_16907,N_16014);
and U19195 (N_19195,N_15206,N_16591);
nand U19196 (N_19196,N_15620,N_16594);
nand U19197 (N_19197,N_15969,N_15369);
xnor U19198 (N_19198,N_17288,N_15604);
and U19199 (N_19199,N_15335,N_15504);
nor U19200 (N_19200,N_15774,N_16274);
nor U19201 (N_19201,N_16946,N_16620);
or U19202 (N_19202,N_17450,N_16362);
xor U19203 (N_19203,N_16704,N_17055);
and U19204 (N_19204,N_16788,N_16157);
nand U19205 (N_19205,N_16247,N_15320);
nand U19206 (N_19206,N_16596,N_16864);
xnor U19207 (N_19207,N_17214,N_16330);
or U19208 (N_19208,N_17342,N_15985);
nor U19209 (N_19209,N_16124,N_16170);
or U19210 (N_19210,N_15221,N_16524);
xnor U19211 (N_19211,N_15800,N_15145);
nor U19212 (N_19212,N_16134,N_17214);
and U19213 (N_19213,N_15736,N_15152);
nor U19214 (N_19214,N_16936,N_15763);
xnor U19215 (N_19215,N_17092,N_17323);
xor U19216 (N_19216,N_15603,N_16509);
nand U19217 (N_19217,N_16850,N_17428);
nand U19218 (N_19218,N_16199,N_15898);
xnor U19219 (N_19219,N_17389,N_16940);
or U19220 (N_19220,N_17326,N_15616);
xnor U19221 (N_19221,N_16856,N_16595);
or U19222 (N_19222,N_17028,N_16117);
and U19223 (N_19223,N_16465,N_15233);
nor U19224 (N_19224,N_15500,N_17163);
and U19225 (N_19225,N_16543,N_16850);
or U19226 (N_19226,N_17432,N_16203);
or U19227 (N_19227,N_15608,N_16476);
and U19228 (N_19228,N_15360,N_17194);
or U19229 (N_19229,N_15416,N_16747);
and U19230 (N_19230,N_15511,N_17265);
xor U19231 (N_19231,N_17035,N_15730);
nor U19232 (N_19232,N_16465,N_15052);
nand U19233 (N_19233,N_15517,N_16478);
nand U19234 (N_19234,N_16519,N_15056);
xor U19235 (N_19235,N_15476,N_17457);
nand U19236 (N_19236,N_15769,N_17318);
or U19237 (N_19237,N_16275,N_15960);
xor U19238 (N_19238,N_15857,N_16456);
nand U19239 (N_19239,N_15514,N_16433);
and U19240 (N_19240,N_15666,N_17054);
nand U19241 (N_19241,N_16004,N_17158);
nand U19242 (N_19242,N_16362,N_17383);
and U19243 (N_19243,N_17258,N_15403);
nand U19244 (N_19244,N_16136,N_16928);
nor U19245 (N_19245,N_17361,N_16315);
nor U19246 (N_19246,N_15548,N_17435);
or U19247 (N_19247,N_16938,N_16480);
nand U19248 (N_19248,N_15721,N_15529);
or U19249 (N_19249,N_16946,N_16248);
or U19250 (N_19250,N_16919,N_15335);
and U19251 (N_19251,N_16667,N_15012);
nor U19252 (N_19252,N_16635,N_15415);
nor U19253 (N_19253,N_17098,N_16304);
nand U19254 (N_19254,N_16273,N_16129);
nor U19255 (N_19255,N_16713,N_17240);
nand U19256 (N_19256,N_15285,N_16925);
or U19257 (N_19257,N_17129,N_17328);
nor U19258 (N_19258,N_17127,N_15759);
and U19259 (N_19259,N_17369,N_16643);
xnor U19260 (N_19260,N_17264,N_16075);
or U19261 (N_19261,N_16492,N_16030);
and U19262 (N_19262,N_15008,N_15675);
nor U19263 (N_19263,N_16988,N_16004);
and U19264 (N_19264,N_15139,N_16688);
and U19265 (N_19265,N_17272,N_17311);
nand U19266 (N_19266,N_16746,N_15026);
or U19267 (N_19267,N_15725,N_17498);
nor U19268 (N_19268,N_15570,N_15343);
and U19269 (N_19269,N_17418,N_17241);
or U19270 (N_19270,N_15409,N_17409);
nand U19271 (N_19271,N_15227,N_16947);
nand U19272 (N_19272,N_16219,N_17000);
and U19273 (N_19273,N_16355,N_16941);
and U19274 (N_19274,N_15404,N_16861);
nand U19275 (N_19275,N_15933,N_15866);
or U19276 (N_19276,N_16068,N_17221);
or U19277 (N_19277,N_16576,N_16987);
nor U19278 (N_19278,N_15203,N_16707);
nor U19279 (N_19279,N_17245,N_15281);
nand U19280 (N_19280,N_15578,N_16086);
xor U19281 (N_19281,N_15772,N_16800);
or U19282 (N_19282,N_16003,N_16617);
nor U19283 (N_19283,N_17152,N_16074);
or U19284 (N_19284,N_15944,N_15444);
or U19285 (N_19285,N_15389,N_16299);
nand U19286 (N_19286,N_15718,N_15889);
nor U19287 (N_19287,N_16886,N_17407);
nor U19288 (N_19288,N_16429,N_15786);
or U19289 (N_19289,N_15367,N_17344);
nand U19290 (N_19290,N_16359,N_17243);
nor U19291 (N_19291,N_16565,N_16762);
nand U19292 (N_19292,N_16682,N_16219);
nor U19293 (N_19293,N_17096,N_17042);
or U19294 (N_19294,N_16771,N_15421);
or U19295 (N_19295,N_16775,N_17168);
or U19296 (N_19296,N_17363,N_17271);
nor U19297 (N_19297,N_17476,N_15844);
xnor U19298 (N_19298,N_15888,N_16989);
xor U19299 (N_19299,N_16424,N_16903);
and U19300 (N_19300,N_15695,N_16697);
xnor U19301 (N_19301,N_16625,N_16116);
nand U19302 (N_19302,N_17256,N_15075);
or U19303 (N_19303,N_16442,N_16009);
xor U19304 (N_19304,N_15755,N_17269);
and U19305 (N_19305,N_15751,N_16255);
or U19306 (N_19306,N_17048,N_17001);
or U19307 (N_19307,N_16830,N_17343);
xor U19308 (N_19308,N_16963,N_17127);
or U19309 (N_19309,N_15949,N_17322);
or U19310 (N_19310,N_15116,N_15772);
nand U19311 (N_19311,N_16329,N_15314);
or U19312 (N_19312,N_16867,N_15832);
xor U19313 (N_19313,N_15590,N_17205);
and U19314 (N_19314,N_15871,N_16935);
xnor U19315 (N_19315,N_16531,N_16798);
or U19316 (N_19316,N_16469,N_16434);
or U19317 (N_19317,N_15388,N_16432);
nand U19318 (N_19318,N_17441,N_17412);
nor U19319 (N_19319,N_15381,N_15373);
nor U19320 (N_19320,N_15689,N_17319);
or U19321 (N_19321,N_15547,N_15256);
or U19322 (N_19322,N_15994,N_15283);
xnor U19323 (N_19323,N_15631,N_16215);
and U19324 (N_19324,N_16188,N_16471);
xnor U19325 (N_19325,N_15130,N_17112);
xor U19326 (N_19326,N_15881,N_17021);
nand U19327 (N_19327,N_16853,N_15901);
nor U19328 (N_19328,N_17284,N_15552);
xor U19329 (N_19329,N_16529,N_15625);
xnor U19330 (N_19330,N_17244,N_17361);
nor U19331 (N_19331,N_15980,N_16121);
and U19332 (N_19332,N_15734,N_17111);
nand U19333 (N_19333,N_15408,N_15474);
nor U19334 (N_19334,N_17380,N_17326);
nand U19335 (N_19335,N_16233,N_15426);
nor U19336 (N_19336,N_17039,N_17266);
or U19337 (N_19337,N_15197,N_15272);
or U19338 (N_19338,N_17318,N_15548);
nand U19339 (N_19339,N_15580,N_15434);
nand U19340 (N_19340,N_16768,N_15924);
nand U19341 (N_19341,N_16852,N_15372);
nor U19342 (N_19342,N_15931,N_17238);
nand U19343 (N_19343,N_16153,N_16772);
xnor U19344 (N_19344,N_15514,N_16377);
or U19345 (N_19345,N_17368,N_15959);
xor U19346 (N_19346,N_15350,N_17236);
and U19347 (N_19347,N_16176,N_16829);
nand U19348 (N_19348,N_15011,N_16760);
or U19349 (N_19349,N_16257,N_16317);
nor U19350 (N_19350,N_15994,N_16616);
xor U19351 (N_19351,N_16570,N_17283);
nor U19352 (N_19352,N_15728,N_15051);
nor U19353 (N_19353,N_16533,N_15470);
nor U19354 (N_19354,N_16041,N_16918);
nand U19355 (N_19355,N_16122,N_16183);
nand U19356 (N_19356,N_15054,N_16055);
nor U19357 (N_19357,N_15970,N_17482);
or U19358 (N_19358,N_15963,N_15641);
nand U19359 (N_19359,N_17079,N_16219);
and U19360 (N_19360,N_15302,N_16707);
nor U19361 (N_19361,N_16618,N_17222);
nor U19362 (N_19362,N_16094,N_16876);
and U19363 (N_19363,N_15273,N_16632);
or U19364 (N_19364,N_17214,N_15263);
and U19365 (N_19365,N_15323,N_17416);
xor U19366 (N_19366,N_16423,N_15353);
and U19367 (N_19367,N_17162,N_16288);
nand U19368 (N_19368,N_15961,N_15583);
xor U19369 (N_19369,N_17325,N_17399);
and U19370 (N_19370,N_15399,N_17075);
and U19371 (N_19371,N_17324,N_16535);
and U19372 (N_19372,N_15559,N_16587);
nor U19373 (N_19373,N_16552,N_15197);
nand U19374 (N_19374,N_15588,N_15208);
xnor U19375 (N_19375,N_15293,N_16211);
nand U19376 (N_19376,N_15299,N_17207);
nand U19377 (N_19377,N_15535,N_17215);
xnor U19378 (N_19378,N_15848,N_17308);
or U19379 (N_19379,N_16386,N_17496);
or U19380 (N_19380,N_15378,N_16112);
or U19381 (N_19381,N_17049,N_17173);
and U19382 (N_19382,N_17395,N_17311);
xnor U19383 (N_19383,N_15435,N_16922);
nor U19384 (N_19384,N_16064,N_15868);
and U19385 (N_19385,N_16425,N_16236);
or U19386 (N_19386,N_15723,N_16574);
nor U19387 (N_19387,N_15442,N_15035);
xnor U19388 (N_19388,N_15563,N_15823);
or U19389 (N_19389,N_17042,N_17052);
nand U19390 (N_19390,N_17412,N_15785);
or U19391 (N_19391,N_15986,N_17138);
xnor U19392 (N_19392,N_16606,N_16880);
or U19393 (N_19393,N_16413,N_15844);
xor U19394 (N_19394,N_16374,N_15319);
xor U19395 (N_19395,N_16708,N_16088);
or U19396 (N_19396,N_16883,N_17168);
xnor U19397 (N_19397,N_17311,N_15506);
nand U19398 (N_19398,N_16064,N_15296);
and U19399 (N_19399,N_15407,N_17140);
nor U19400 (N_19400,N_15552,N_16703);
or U19401 (N_19401,N_16312,N_16211);
nor U19402 (N_19402,N_15099,N_17476);
and U19403 (N_19403,N_15168,N_15601);
xnor U19404 (N_19404,N_16021,N_16070);
and U19405 (N_19405,N_15637,N_16816);
nor U19406 (N_19406,N_16969,N_17096);
xnor U19407 (N_19407,N_16150,N_15010);
nor U19408 (N_19408,N_15608,N_15382);
nand U19409 (N_19409,N_16156,N_15623);
and U19410 (N_19410,N_15544,N_17246);
and U19411 (N_19411,N_15679,N_15513);
xor U19412 (N_19412,N_16242,N_15581);
and U19413 (N_19413,N_17323,N_15900);
or U19414 (N_19414,N_15214,N_15404);
and U19415 (N_19415,N_16515,N_17017);
xor U19416 (N_19416,N_17182,N_15154);
nand U19417 (N_19417,N_15769,N_16113);
or U19418 (N_19418,N_15950,N_16281);
nand U19419 (N_19419,N_15526,N_17424);
xor U19420 (N_19420,N_15376,N_15333);
nor U19421 (N_19421,N_15025,N_17059);
or U19422 (N_19422,N_17373,N_17350);
xor U19423 (N_19423,N_15597,N_16912);
xnor U19424 (N_19424,N_16604,N_17148);
or U19425 (N_19425,N_17121,N_15430);
xor U19426 (N_19426,N_16168,N_16328);
and U19427 (N_19427,N_15403,N_15890);
xnor U19428 (N_19428,N_17141,N_16509);
and U19429 (N_19429,N_15282,N_15132);
or U19430 (N_19430,N_16113,N_15599);
xor U19431 (N_19431,N_17405,N_15092);
nor U19432 (N_19432,N_15963,N_17324);
xnor U19433 (N_19433,N_17253,N_16201);
nor U19434 (N_19434,N_16378,N_16785);
or U19435 (N_19435,N_16152,N_15935);
xor U19436 (N_19436,N_16679,N_15782);
and U19437 (N_19437,N_15240,N_15767);
nand U19438 (N_19438,N_16010,N_15824);
xor U19439 (N_19439,N_16659,N_15471);
xor U19440 (N_19440,N_17309,N_16457);
and U19441 (N_19441,N_15951,N_15042);
or U19442 (N_19442,N_15997,N_15663);
nor U19443 (N_19443,N_15838,N_15912);
or U19444 (N_19444,N_15049,N_15118);
nand U19445 (N_19445,N_16071,N_17196);
nor U19446 (N_19446,N_15531,N_15362);
nor U19447 (N_19447,N_16685,N_16882);
or U19448 (N_19448,N_15775,N_15771);
xnor U19449 (N_19449,N_15386,N_16821);
xor U19450 (N_19450,N_16528,N_15287);
xor U19451 (N_19451,N_16458,N_16153);
nor U19452 (N_19452,N_16697,N_15983);
xnor U19453 (N_19453,N_16751,N_16181);
or U19454 (N_19454,N_16836,N_15406);
xnor U19455 (N_19455,N_16728,N_15009);
nand U19456 (N_19456,N_15425,N_16678);
xnor U19457 (N_19457,N_16632,N_15773);
or U19458 (N_19458,N_16962,N_16445);
or U19459 (N_19459,N_17361,N_15633);
and U19460 (N_19460,N_17407,N_15770);
nor U19461 (N_19461,N_17470,N_17175);
xnor U19462 (N_19462,N_15857,N_17450);
nor U19463 (N_19463,N_16519,N_15067);
and U19464 (N_19464,N_16820,N_15013);
or U19465 (N_19465,N_15699,N_16694);
nand U19466 (N_19466,N_17019,N_15433);
xnor U19467 (N_19467,N_16482,N_15080);
nor U19468 (N_19468,N_15545,N_16489);
or U19469 (N_19469,N_16508,N_15968);
or U19470 (N_19470,N_16525,N_17128);
or U19471 (N_19471,N_16779,N_15443);
or U19472 (N_19472,N_15132,N_15167);
xor U19473 (N_19473,N_16057,N_16727);
and U19474 (N_19474,N_15844,N_17394);
and U19475 (N_19475,N_16734,N_16943);
xor U19476 (N_19476,N_15462,N_15526);
nand U19477 (N_19477,N_15224,N_15081);
xnor U19478 (N_19478,N_17487,N_15509);
or U19479 (N_19479,N_17152,N_16242);
nor U19480 (N_19480,N_15008,N_16138);
xnor U19481 (N_19481,N_16956,N_15369);
nand U19482 (N_19482,N_16777,N_17144);
or U19483 (N_19483,N_16573,N_16284);
or U19484 (N_19484,N_16190,N_15018);
and U19485 (N_19485,N_16218,N_15875);
or U19486 (N_19486,N_16755,N_16828);
nand U19487 (N_19487,N_15577,N_16497);
or U19488 (N_19488,N_15677,N_16941);
and U19489 (N_19489,N_16231,N_17345);
and U19490 (N_19490,N_17007,N_15182);
nor U19491 (N_19491,N_16343,N_15631);
nand U19492 (N_19492,N_15863,N_17469);
or U19493 (N_19493,N_16810,N_17468);
or U19494 (N_19494,N_15915,N_16825);
xor U19495 (N_19495,N_15191,N_15737);
nor U19496 (N_19496,N_15329,N_15439);
nand U19497 (N_19497,N_15869,N_16490);
and U19498 (N_19498,N_16900,N_16541);
or U19499 (N_19499,N_17473,N_16220);
or U19500 (N_19500,N_15192,N_15746);
xnor U19501 (N_19501,N_15880,N_16968);
or U19502 (N_19502,N_15892,N_17197);
and U19503 (N_19503,N_16925,N_16781);
or U19504 (N_19504,N_15243,N_17150);
xor U19505 (N_19505,N_17362,N_15063);
nor U19506 (N_19506,N_16114,N_17408);
nand U19507 (N_19507,N_16333,N_16002);
nand U19508 (N_19508,N_16258,N_17096);
nand U19509 (N_19509,N_16244,N_16245);
or U19510 (N_19510,N_15110,N_17017);
xor U19511 (N_19511,N_16818,N_16191);
nor U19512 (N_19512,N_15631,N_17259);
or U19513 (N_19513,N_17105,N_16432);
and U19514 (N_19514,N_16109,N_15456);
nor U19515 (N_19515,N_15883,N_16087);
nand U19516 (N_19516,N_15086,N_16502);
nand U19517 (N_19517,N_15602,N_17296);
xor U19518 (N_19518,N_15946,N_16217);
xnor U19519 (N_19519,N_17087,N_15657);
xor U19520 (N_19520,N_16362,N_16748);
and U19521 (N_19521,N_15097,N_15653);
nand U19522 (N_19522,N_15960,N_15429);
nor U19523 (N_19523,N_16523,N_15136);
or U19524 (N_19524,N_16452,N_17059);
nor U19525 (N_19525,N_15488,N_16524);
and U19526 (N_19526,N_16965,N_16561);
nor U19527 (N_19527,N_17456,N_15992);
xor U19528 (N_19528,N_16474,N_17238);
nand U19529 (N_19529,N_17479,N_16345);
nand U19530 (N_19530,N_17436,N_15467);
or U19531 (N_19531,N_15843,N_16254);
nor U19532 (N_19532,N_15884,N_16994);
or U19533 (N_19533,N_17174,N_15977);
xnor U19534 (N_19534,N_16052,N_15284);
nor U19535 (N_19535,N_15035,N_16828);
xnor U19536 (N_19536,N_17203,N_15263);
xor U19537 (N_19537,N_16542,N_16625);
nand U19538 (N_19538,N_17328,N_16938);
xor U19539 (N_19539,N_15951,N_17216);
nand U19540 (N_19540,N_16857,N_15218);
nor U19541 (N_19541,N_15114,N_17050);
nand U19542 (N_19542,N_16997,N_16887);
nand U19543 (N_19543,N_15652,N_16797);
nand U19544 (N_19544,N_16420,N_15668);
xor U19545 (N_19545,N_16840,N_15567);
nand U19546 (N_19546,N_15542,N_15537);
xnor U19547 (N_19547,N_17218,N_17252);
and U19548 (N_19548,N_16716,N_16672);
xor U19549 (N_19549,N_16021,N_16821);
nor U19550 (N_19550,N_17018,N_16053);
xor U19551 (N_19551,N_16623,N_17264);
or U19552 (N_19552,N_15821,N_17118);
nor U19553 (N_19553,N_16827,N_16455);
xnor U19554 (N_19554,N_17314,N_17308);
xor U19555 (N_19555,N_15876,N_16129);
nor U19556 (N_19556,N_15299,N_15643);
nor U19557 (N_19557,N_16491,N_15932);
xnor U19558 (N_19558,N_15501,N_15709);
nor U19559 (N_19559,N_15021,N_17160);
or U19560 (N_19560,N_16142,N_16439);
and U19561 (N_19561,N_15105,N_16121);
and U19562 (N_19562,N_17010,N_16110);
nand U19563 (N_19563,N_15729,N_17042);
or U19564 (N_19564,N_16854,N_15909);
and U19565 (N_19565,N_15611,N_17146);
or U19566 (N_19566,N_15846,N_15695);
nor U19567 (N_19567,N_16603,N_17361);
or U19568 (N_19568,N_16884,N_15416);
nor U19569 (N_19569,N_17335,N_16164);
or U19570 (N_19570,N_15190,N_15742);
or U19571 (N_19571,N_15353,N_15160);
nand U19572 (N_19572,N_16657,N_15716);
nand U19573 (N_19573,N_15424,N_15335);
xnor U19574 (N_19574,N_15753,N_15287);
nand U19575 (N_19575,N_16827,N_15336);
and U19576 (N_19576,N_16256,N_17452);
nor U19577 (N_19577,N_15410,N_17343);
or U19578 (N_19578,N_15356,N_15262);
or U19579 (N_19579,N_16637,N_15915);
and U19580 (N_19580,N_16252,N_15455);
xnor U19581 (N_19581,N_15171,N_15442);
xor U19582 (N_19582,N_15467,N_15087);
or U19583 (N_19583,N_15273,N_15897);
and U19584 (N_19584,N_15909,N_17307);
and U19585 (N_19585,N_15941,N_16457);
or U19586 (N_19586,N_16802,N_16402);
or U19587 (N_19587,N_16772,N_16996);
xnor U19588 (N_19588,N_16602,N_16252);
or U19589 (N_19589,N_16682,N_15722);
or U19590 (N_19590,N_17265,N_16468);
nand U19591 (N_19591,N_16257,N_16847);
nor U19592 (N_19592,N_15477,N_17039);
nand U19593 (N_19593,N_16157,N_15480);
nor U19594 (N_19594,N_16590,N_15378);
nor U19595 (N_19595,N_15584,N_15903);
nor U19596 (N_19596,N_16803,N_15239);
and U19597 (N_19597,N_15963,N_16070);
xor U19598 (N_19598,N_15231,N_16997);
nor U19599 (N_19599,N_16863,N_15248);
and U19600 (N_19600,N_16792,N_16937);
xor U19601 (N_19601,N_16441,N_17312);
nand U19602 (N_19602,N_16074,N_16250);
nor U19603 (N_19603,N_15893,N_16122);
and U19604 (N_19604,N_15830,N_17495);
and U19605 (N_19605,N_15625,N_15129);
or U19606 (N_19606,N_17407,N_15846);
nor U19607 (N_19607,N_15199,N_17256);
nand U19608 (N_19608,N_17143,N_15606);
xnor U19609 (N_19609,N_16778,N_16780);
nand U19610 (N_19610,N_15154,N_16983);
and U19611 (N_19611,N_16793,N_15289);
nor U19612 (N_19612,N_17422,N_16967);
nand U19613 (N_19613,N_16610,N_16739);
nor U19614 (N_19614,N_15005,N_17208);
xnor U19615 (N_19615,N_16622,N_15450);
nor U19616 (N_19616,N_16950,N_15583);
nand U19617 (N_19617,N_16293,N_16146);
xnor U19618 (N_19618,N_17315,N_16251);
and U19619 (N_19619,N_16752,N_15244);
and U19620 (N_19620,N_16233,N_16396);
nor U19621 (N_19621,N_16000,N_15101);
or U19622 (N_19622,N_16867,N_17425);
xor U19623 (N_19623,N_16420,N_16599);
or U19624 (N_19624,N_16863,N_16777);
nand U19625 (N_19625,N_15928,N_16854);
and U19626 (N_19626,N_17303,N_16393);
nor U19627 (N_19627,N_15226,N_15016);
and U19628 (N_19628,N_15677,N_17231);
and U19629 (N_19629,N_16960,N_16522);
or U19630 (N_19630,N_15387,N_17291);
xnor U19631 (N_19631,N_15288,N_15910);
or U19632 (N_19632,N_15865,N_16801);
and U19633 (N_19633,N_17463,N_16088);
or U19634 (N_19634,N_17214,N_17000);
nand U19635 (N_19635,N_17023,N_16749);
or U19636 (N_19636,N_17020,N_15469);
nor U19637 (N_19637,N_16033,N_16541);
nor U19638 (N_19638,N_15259,N_17315);
nand U19639 (N_19639,N_15050,N_16688);
xor U19640 (N_19640,N_16221,N_16624);
nand U19641 (N_19641,N_16318,N_16080);
and U19642 (N_19642,N_15783,N_15889);
xor U19643 (N_19643,N_16187,N_16699);
nor U19644 (N_19644,N_17266,N_15831);
or U19645 (N_19645,N_16532,N_15542);
nand U19646 (N_19646,N_17106,N_17021);
nor U19647 (N_19647,N_15976,N_17221);
nand U19648 (N_19648,N_15437,N_16705);
and U19649 (N_19649,N_15687,N_16815);
nor U19650 (N_19650,N_15496,N_15278);
and U19651 (N_19651,N_16509,N_17160);
nor U19652 (N_19652,N_16392,N_15997);
nor U19653 (N_19653,N_15192,N_16037);
xor U19654 (N_19654,N_17424,N_15480);
nand U19655 (N_19655,N_15170,N_15505);
or U19656 (N_19656,N_16602,N_17174);
nand U19657 (N_19657,N_16910,N_16787);
xor U19658 (N_19658,N_15508,N_15075);
or U19659 (N_19659,N_17421,N_16166);
or U19660 (N_19660,N_15880,N_15368);
or U19661 (N_19661,N_16941,N_15707);
xor U19662 (N_19662,N_15189,N_15786);
or U19663 (N_19663,N_16900,N_16404);
nor U19664 (N_19664,N_15501,N_15820);
and U19665 (N_19665,N_16685,N_15818);
xnor U19666 (N_19666,N_15846,N_16513);
nor U19667 (N_19667,N_15536,N_16643);
and U19668 (N_19668,N_17089,N_17023);
and U19669 (N_19669,N_16884,N_15306);
nand U19670 (N_19670,N_15267,N_17330);
nor U19671 (N_19671,N_16177,N_17212);
nand U19672 (N_19672,N_15823,N_16158);
xnor U19673 (N_19673,N_17008,N_17009);
xor U19674 (N_19674,N_15312,N_17338);
and U19675 (N_19675,N_17203,N_15447);
xnor U19676 (N_19676,N_15930,N_15222);
nor U19677 (N_19677,N_16999,N_15008);
xor U19678 (N_19678,N_16604,N_17308);
and U19679 (N_19679,N_16658,N_16854);
and U19680 (N_19680,N_15637,N_15203);
xnor U19681 (N_19681,N_17098,N_16278);
and U19682 (N_19682,N_17276,N_16646);
xor U19683 (N_19683,N_16784,N_15221);
or U19684 (N_19684,N_16719,N_16805);
xor U19685 (N_19685,N_15949,N_16281);
and U19686 (N_19686,N_17016,N_15936);
and U19687 (N_19687,N_16936,N_15881);
nand U19688 (N_19688,N_17169,N_16893);
or U19689 (N_19689,N_16615,N_16173);
xnor U19690 (N_19690,N_16515,N_16977);
nor U19691 (N_19691,N_15360,N_15624);
nor U19692 (N_19692,N_17324,N_17201);
and U19693 (N_19693,N_16659,N_15321);
or U19694 (N_19694,N_15364,N_15581);
nor U19695 (N_19695,N_16917,N_15293);
nand U19696 (N_19696,N_16178,N_16924);
xor U19697 (N_19697,N_16531,N_16853);
and U19698 (N_19698,N_17292,N_16758);
xnor U19699 (N_19699,N_16918,N_16725);
xor U19700 (N_19700,N_17213,N_15998);
xnor U19701 (N_19701,N_15428,N_15900);
nand U19702 (N_19702,N_16095,N_16782);
and U19703 (N_19703,N_15004,N_16837);
nand U19704 (N_19704,N_15777,N_17251);
and U19705 (N_19705,N_16825,N_16752);
and U19706 (N_19706,N_15396,N_16721);
and U19707 (N_19707,N_15821,N_16229);
and U19708 (N_19708,N_16304,N_16659);
or U19709 (N_19709,N_15503,N_16837);
and U19710 (N_19710,N_15213,N_15750);
or U19711 (N_19711,N_15092,N_16290);
nor U19712 (N_19712,N_17487,N_15159);
nand U19713 (N_19713,N_15687,N_16160);
nand U19714 (N_19714,N_16683,N_15328);
xor U19715 (N_19715,N_16778,N_16960);
xnor U19716 (N_19716,N_16376,N_16430);
nand U19717 (N_19717,N_15612,N_16624);
xnor U19718 (N_19718,N_15008,N_15172);
xnor U19719 (N_19719,N_15103,N_15328);
nor U19720 (N_19720,N_15538,N_16884);
or U19721 (N_19721,N_16647,N_17187);
nand U19722 (N_19722,N_17439,N_15492);
nand U19723 (N_19723,N_17067,N_16001);
nor U19724 (N_19724,N_17466,N_16197);
or U19725 (N_19725,N_17046,N_17176);
and U19726 (N_19726,N_15991,N_16111);
and U19727 (N_19727,N_17283,N_15871);
nand U19728 (N_19728,N_15041,N_15780);
nand U19729 (N_19729,N_15512,N_16409);
or U19730 (N_19730,N_16468,N_16990);
or U19731 (N_19731,N_16572,N_15934);
and U19732 (N_19732,N_16349,N_15774);
nor U19733 (N_19733,N_16817,N_15916);
and U19734 (N_19734,N_15028,N_16931);
nor U19735 (N_19735,N_15018,N_15198);
xor U19736 (N_19736,N_15634,N_15053);
nor U19737 (N_19737,N_16052,N_17455);
or U19738 (N_19738,N_17167,N_15841);
and U19739 (N_19739,N_17043,N_16646);
nor U19740 (N_19740,N_15000,N_16493);
nor U19741 (N_19741,N_15845,N_16680);
or U19742 (N_19742,N_17067,N_16807);
or U19743 (N_19743,N_15077,N_15678);
xor U19744 (N_19744,N_15874,N_15442);
nor U19745 (N_19745,N_16365,N_15499);
nand U19746 (N_19746,N_16194,N_15744);
or U19747 (N_19747,N_15471,N_15603);
xnor U19748 (N_19748,N_16399,N_16939);
xnor U19749 (N_19749,N_16887,N_15183);
nor U19750 (N_19750,N_15896,N_17105);
nor U19751 (N_19751,N_15380,N_17052);
and U19752 (N_19752,N_15017,N_15122);
nor U19753 (N_19753,N_16229,N_15273);
and U19754 (N_19754,N_15585,N_16464);
and U19755 (N_19755,N_16620,N_15011);
xor U19756 (N_19756,N_16604,N_15744);
nor U19757 (N_19757,N_16790,N_15834);
or U19758 (N_19758,N_15753,N_15833);
and U19759 (N_19759,N_15122,N_16782);
or U19760 (N_19760,N_15243,N_16628);
nand U19761 (N_19761,N_16261,N_15955);
or U19762 (N_19762,N_17369,N_15692);
nand U19763 (N_19763,N_17068,N_17308);
nand U19764 (N_19764,N_17495,N_15613);
nand U19765 (N_19765,N_15304,N_15536);
xnor U19766 (N_19766,N_17313,N_16309);
nand U19767 (N_19767,N_15491,N_15713);
nor U19768 (N_19768,N_15945,N_16555);
or U19769 (N_19769,N_17047,N_15929);
or U19770 (N_19770,N_16881,N_15401);
xnor U19771 (N_19771,N_15697,N_16174);
nor U19772 (N_19772,N_16065,N_16257);
nand U19773 (N_19773,N_17108,N_15941);
nand U19774 (N_19774,N_16826,N_17367);
or U19775 (N_19775,N_17232,N_15356);
nand U19776 (N_19776,N_15562,N_15226);
nand U19777 (N_19777,N_15499,N_16750);
and U19778 (N_19778,N_16168,N_15365);
xor U19779 (N_19779,N_16733,N_15533);
nand U19780 (N_19780,N_15167,N_15656);
xnor U19781 (N_19781,N_15642,N_17249);
or U19782 (N_19782,N_16103,N_17048);
nand U19783 (N_19783,N_15798,N_16990);
xnor U19784 (N_19784,N_17042,N_15945);
and U19785 (N_19785,N_15902,N_16967);
nand U19786 (N_19786,N_15223,N_16680);
nand U19787 (N_19787,N_16192,N_15215);
and U19788 (N_19788,N_16291,N_16802);
nor U19789 (N_19789,N_15713,N_15804);
or U19790 (N_19790,N_16654,N_16055);
nor U19791 (N_19791,N_17106,N_15701);
nand U19792 (N_19792,N_17433,N_15427);
xnor U19793 (N_19793,N_15233,N_15567);
nand U19794 (N_19794,N_17480,N_17003);
xnor U19795 (N_19795,N_17437,N_16760);
nor U19796 (N_19796,N_17064,N_15476);
or U19797 (N_19797,N_16225,N_16540);
and U19798 (N_19798,N_16307,N_15506);
nand U19799 (N_19799,N_16933,N_15221);
or U19800 (N_19800,N_17409,N_17153);
nand U19801 (N_19801,N_15801,N_17336);
or U19802 (N_19802,N_17185,N_15816);
and U19803 (N_19803,N_17044,N_16748);
or U19804 (N_19804,N_16766,N_17065);
or U19805 (N_19805,N_16669,N_17109);
nand U19806 (N_19806,N_16942,N_15606);
nand U19807 (N_19807,N_15317,N_16122);
nor U19808 (N_19808,N_16038,N_15349);
or U19809 (N_19809,N_15674,N_16173);
and U19810 (N_19810,N_15017,N_16756);
nand U19811 (N_19811,N_15922,N_16852);
xnor U19812 (N_19812,N_16008,N_16797);
nand U19813 (N_19813,N_16882,N_15726);
xnor U19814 (N_19814,N_16445,N_15024);
nand U19815 (N_19815,N_17294,N_15446);
xnor U19816 (N_19816,N_17312,N_15021);
xnor U19817 (N_19817,N_16415,N_15161);
nor U19818 (N_19818,N_17278,N_15101);
or U19819 (N_19819,N_15184,N_15798);
and U19820 (N_19820,N_17221,N_17432);
nand U19821 (N_19821,N_16474,N_15653);
nand U19822 (N_19822,N_16694,N_17046);
and U19823 (N_19823,N_17209,N_16214);
xnor U19824 (N_19824,N_15183,N_17474);
xor U19825 (N_19825,N_16940,N_16445);
and U19826 (N_19826,N_17199,N_15608);
nor U19827 (N_19827,N_17153,N_15265);
xnor U19828 (N_19828,N_17407,N_16015);
and U19829 (N_19829,N_17115,N_16794);
xnor U19830 (N_19830,N_17360,N_16833);
xnor U19831 (N_19831,N_16922,N_16804);
xnor U19832 (N_19832,N_15214,N_16569);
and U19833 (N_19833,N_16847,N_17101);
nor U19834 (N_19834,N_16389,N_16707);
nand U19835 (N_19835,N_15978,N_15510);
xnor U19836 (N_19836,N_15637,N_16873);
nor U19837 (N_19837,N_16288,N_16174);
nor U19838 (N_19838,N_16905,N_16822);
and U19839 (N_19839,N_15498,N_16326);
nand U19840 (N_19840,N_15634,N_15474);
and U19841 (N_19841,N_15311,N_17158);
nand U19842 (N_19842,N_16985,N_15159);
nor U19843 (N_19843,N_17435,N_17395);
or U19844 (N_19844,N_15627,N_16227);
or U19845 (N_19845,N_17386,N_15027);
or U19846 (N_19846,N_16869,N_15840);
and U19847 (N_19847,N_17265,N_15086);
xor U19848 (N_19848,N_17324,N_15284);
nor U19849 (N_19849,N_15239,N_16575);
and U19850 (N_19850,N_17048,N_16898);
nand U19851 (N_19851,N_16261,N_17161);
nand U19852 (N_19852,N_16016,N_16926);
and U19853 (N_19853,N_15248,N_15587);
nand U19854 (N_19854,N_15409,N_15963);
nor U19855 (N_19855,N_17168,N_16778);
and U19856 (N_19856,N_16227,N_17330);
nor U19857 (N_19857,N_15055,N_16008);
or U19858 (N_19858,N_16975,N_15497);
nand U19859 (N_19859,N_16130,N_16785);
or U19860 (N_19860,N_17043,N_15809);
and U19861 (N_19861,N_16893,N_16250);
nor U19862 (N_19862,N_16121,N_16539);
nor U19863 (N_19863,N_16965,N_15009);
nand U19864 (N_19864,N_15036,N_15477);
nand U19865 (N_19865,N_16500,N_15743);
nor U19866 (N_19866,N_15115,N_15087);
and U19867 (N_19867,N_15243,N_16806);
nor U19868 (N_19868,N_17478,N_15911);
or U19869 (N_19869,N_15579,N_16319);
xnor U19870 (N_19870,N_15407,N_16488);
xnor U19871 (N_19871,N_16413,N_17334);
and U19872 (N_19872,N_15620,N_16865);
nand U19873 (N_19873,N_15231,N_17074);
nor U19874 (N_19874,N_15151,N_16729);
xnor U19875 (N_19875,N_17220,N_17246);
nand U19876 (N_19876,N_15412,N_17083);
or U19877 (N_19877,N_16730,N_16386);
nor U19878 (N_19878,N_16401,N_15959);
nor U19879 (N_19879,N_15106,N_15593);
nor U19880 (N_19880,N_15658,N_16017);
or U19881 (N_19881,N_15038,N_15323);
or U19882 (N_19882,N_15093,N_16193);
or U19883 (N_19883,N_16471,N_16539);
and U19884 (N_19884,N_16120,N_15939);
or U19885 (N_19885,N_15501,N_15532);
and U19886 (N_19886,N_16260,N_15131);
or U19887 (N_19887,N_17195,N_16371);
nor U19888 (N_19888,N_15763,N_15018);
nand U19889 (N_19889,N_17437,N_15816);
nand U19890 (N_19890,N_15251,N_17064);
and U19891 (N_19891,N_16706,N_15810);
and U19892 (N_19892,N_15504,N_15477);
nor U19893 (N_19893,N_17441,N_15483);
nor U19894 (N_19894,N_16039,N_16313);
and U19895 (N_19895,N_17219,N_16347);
or U19896 (N_19896,N_16084,N_16429);
xor U19897 (N_19897,N_16822,N_15541);
xnor U19898 (N_19898,N_16713,N_17272);
nand U19899 (N_19899,N_16294,N_17108);
nor U19900 (N_19900,N_16857,N_16734);
nor U19901 (N_19901,N_15726,N_17189);
xnor U19902 (N_19902,N_16040,N_15619);
and U19903 (N_19903,N_15675,N_15987);
and U19904 (N_19904,N_15724,N_16960);
xor U19905 (N_19905,N_16435,N_17209);
or U19906 (N_19906,N_15581,N_16095);
xor U19907 (N_19907,N_16021,N_16506);
and U19908 (N_19908,N_16032,N_16446);
nand U19909 (N_19909,N_15051,N_15033);
or U19910 (N_19910,N_16581,N_16695);
and U19911 (N_19911,N_16751,N_16741);
and U19912 (N_19912,N_16010,N_15502);
nor U19913 (N_19913,N_16214,N_16422);
xor U19914 (N_19914,N_16702,N_16413);
nor U19915 (N_19915,N_15206,N_16182);
and U19916 (N_19916,N_17111,N_15193);
xnor U19917 (N_19917,N_15247,N_15533);
xor U19918 (N_19918,N_16692,N_16928);
nor U19919 (N_19919,N_15274,N_15762);
xor U19920 (N_19920,N_15465,N_15560);
xor U19921 (N_19921,N_16101,N_16660);
xnor U19922 (N_19922,N_16377,N_15030);
nand U19923 (N_19923,N_15146,N_16953);
nor U19924 (N_19924,N_16611,N_16380);
nand U19925 (N_19925,N_16203,N_15733);
xnor U19926 (N_19926,N_17132,N_15571);
nor U19927 (N_19927,N_16158,N_16656);
and U19928 (N_19928,N_16884,N_16221);
and U19929 (N_19929,N_16503,N_15778);
and U19930 (N_19930,N_15686,N_16830);
and U19931 (N_19931,N_15639,N_15838);
nor U19932 (N_19932,N_17043,N_15404);
and U19933 (N_19933,N_15673,N_15130);
nor U19934 (N_19934,N_17229,N_17106);
xor U19935 (N_19935,N_16345,N_15178);
and U19936 (N_19936,N_17390,N_16025);
and U19937 (N_19937,N_15536,N_17252);
nand U19938 (N_19938,N_15839,N_15691);
nor U19939 (N_19939,N_16869,N_16520);
nor U19940 (N_19940,N_15514,N_15458);
xnor U19941 (N_19941,N_15763,N_16180);
xor U19942 (N_19942,N_15291,N_16616);
and U19943 (N_19943,N_16143,N_16190);
or U19944 (N_19944,N_15564,N_17363);
nand U19945 (N_19945,N_15351,N_15384);
nand U19946 (N_19946,N_17335,N_16483);
xnor U19947 (N_19947,N_15425,N_17133);
and U19948 (N_19948,N_15115,N_17168);
and U19949 (N_19949,N_15140,N_16611);
nand U19950 (N_19950,N_16400,N_16038);
xnor U19951 (N_19951,N_15065,N_17007);
or U19952 (N_19952,N_15981,N_17141);
nand U19953 (N_19953,N_15177,N_15093);
and U19954 (N_19954,N_15541,N_17344);
and U19955 (N_19955,N_15290,N_15774);
and U19956 (N_19956,N_17235,N_15517);
and U19957 (N_19957,N_15334,N_16165);
nand U19958 (N_19958,N_16555,N_16695);
and U19959 (N_19959,N_16622,N_15599);
or U19960 (N_19960,N_15015,N_16308);
or U19961 (N_19961,N_17298,N_15803);
or U19962 (N_19962,N_16099,N_17186);
nor U19963 (N_19963,N_16637,N_17159);
or U19964 (N_19964,N_16617,N_17000);
nand U19965 (N_19965,N_15187,N_16463);
nand U19966 (N_19966,N_16106,N_16322);
and U19967 (N_19967,N_15021,N_17218);
and U19968 (N_19968,N_15079,N_17105);
xnor U19969 (N_19969,N_15174,N_16341);
and U19970 (N_19970,N_15747,N_17076);
or U19971 (N_19971,N_15324,N_17051);
nand U19972 (N_19972,N_15669,N_16474);
and U19973 (N_19973,N_15800,N_16251);
or U19974 (N_19974,N_15823,N_16867);
nand U19975 (N_19975,N_15242,N_16399);
nor U19976 (N_19976,N_15978,N_15718);
xor U19977 (N_19977,N_15438,N_17153);
nand U19978 (N_19978,N_17315,N_17209);
and U19979 (N_19979,N_15942,N_15767);
and U19980 (N_19980,N_15124,N_17303);
or U19981 (N_19981,N_16004,N_15719);
nand U19982 (N_19982,N_15003,N_15267);
nand U19983 (N_19983,N_16829,N_16785);
nor U19984 (N_19984,N_15250,N_16153);
and U19985 (N_19985,N_16125,N_15626);
nand U19986 (N_19986,N_16893,N_17332);
and U19987 (N_19987,N_15342,N_16469);
nor U19988 (N_19988,N_17155,N_15155);
nand U19989 (N_19989,N_15015,N_16092);
xnor U19990 (N_19990,N_17159,N_16581);
xnor U19991 (N_19991,N_15977,N_16767);
and U19992 (N_19992,N_15182,N_15905);
nand U19993 (N_19993,N_15536,N_15155);
and U19994 (N_19994,N_15508,N_16285);
xor U19995 (N_19995,N_15496,N_16673);
xnor U19996 (N_19996,N_15540,N_15887);
nand U19997 (N_19997,N_16990,N_17198);
nor U19998 (N_19998,N_16756,N_15146);
xnor U19999 (N_19999,N_17270,N_15282);
and U20000 (N_20000,N_18380,N_18490);
or U20001 (N_20001,N_19583,N_17691);
nand U20002 (N_20002,N_19230,N_18275);
xor U20003 (N_20003,N_19571,N_19040);
nor U20004 (N_20004,N_19975,N_18202);
nor U20005 (N_20005,N_19067,N_18212);
nor U20006 (N_20006,N_18929,N_18952);
xor U20007 (N_20007,N_18297,N_19052);
and U20008 (N_20008,N_19661,N_18256);
xnor U20009 (N_20009,N_17969,N_18957);
nor U20010 (N_20010,N_18149,N_18999);
xor U20011 (N_20011,N_17783,N_19197);
xnor U20012 (N_20012,N_19989,N_17800);
nor U20013 (N_20013,N_18362,N_18540);
nor U20014 (N_20014,N_18290,N_18386);
xor U20015 (N_20015,N_19203,N_18532);
xnor U20016 (N_20016,N_18670,N_19075);
nand U20017 (N_20017,N_18280,N_18916);
nand U20018 (N_20018,N_17877,N_18026);
nor U20019 (N_20019,N_18176,N_18631);
nand U20020 (N_20020,N_18828,N_18864);
xor U20021 (N_20021,N_19106,N_18608);
nand U20022 (N_20022,N_19033,N_18397);
xnor U20023 (N_20023,N_17957,N_18955);
xnor U20024 (N_20024,N_19171,N_19003);
nand U20025 (N_20025,N_19678,N_19452);
xnor U20026 (N_20026,N_19167,N_18111);
or U20027 (N_20027,N_17580,N_18000);
nand U20028 (N_20028,N_18527,N_19775);
xnor U20029 (N_20029,N_18698,N_19814);
nor U20030 (N_20030,N_17671,N_18604);
and U20031 (N_20031,N_19994,N_18791);
nand U20032 (N_20032,N_19689,N_19290);
and U20033 (N_20033,N_19022,N_19313);
xnor U20034 (N_20034,N_18376,N_18882);
and U20035 (N_20035,N_17700,N_19972);
and U20036 (N_20036,N_18457,N_19114);
xnor U20037 (N_20037,N_19327,N_17899);
nand U20038 (N_20038,N_17790,N_18979);
nand U20039 (N_20039,N_19261,N_18143);
or U20040 (N_20040,N_19981,N_17587);
nor U20041 (N_20041,N_19800,N_17649);
and U20042 (N_20042,N_19468,N_19911);
and U20043 (N_20043,N_19978,N_19748);
and U20044 (N_20044,N_19785,N_19935);
and U20045 (N_20045,N_18968,N_17636);
xor U20046 (N_20046,N_18181,N_18492);
xnor U20047 (N_20047,N_17923,N_18807);
xnor U20048 (N_20048,N_19995,N_18482);
nand U20049 (N_20049,N_19716,N_18555);
xor U20050 (N_20050,N_17962,N_18217);
nor U20051 (N_20051,N_17904,N_19077);
nand U20052 (N_20052,N_19317,N_19427);
or U20053 (N_20053,N_18255,N_18034);
and U20054 (N_20054,N_18860,N_18767);
or U20055 (N_20055,N_18266,N_17801);
or U20056 (N_20056,N_17827,N_17832);
xnor U20057 (N_20057,N_19553,N_18182);
nand U20058 (N_20058,N_19915,N_19777);
and U20059 (N_20059,N_18675,N_19241);
or U20060 (N_20060,N_18095,N_17811);
and U20061 (N_20061,N_18312,N_18680);
nand U20062 (N_20062,N_18534,N_19130);
and U20063 (N_20063,N_18384,N_17606);
and U20064 (N_20064,N_18629,N_19474);
and U20065 (N_20065,N_19269,N_18300);
nand U20066 (N_20066,N_18552,N_18812);
nor U20067 (N_20067,N_18100,N_18461);
xor U20068 (N_20068,N_17753,N_17973);
or U20069 (N_20069,N_19168,N_18713);
and U20070 (N_20070,N_18684,N_18742);
nor U20071 (N_20071,N_19416,N_19840);
or U20072 (N_20072,N_18355,N_19532);
nor U20073 (N_20073,N_17975,N_18852);
and U20074 (N_20074,N_19201,N_19883);
or U20075 (N_20075,N_18031,N_18197);
and U20076 (N_20076,N_18502,N_17901);
or U20077 (N_20077,N_19219,N_19918);
nor U20078 (N_20078,N_18984,N_19023);
and U20079 (N_20079,N_18271,N_18654);
nand U20080 (N_20080,N_17559,N_18263);
nor U20081 (N_20081,N_18986,N_19070);
and U20082 (N_20082,N_18020,N_17946);
nor U20083 (N_20083,N_18792,N_19734);
xor U20084 (N_20084,N_17906,N_18706);
or U20085 (N_20085,N_19369,N_17803);
and U20086 (N_20086,N_19457,N_19148);
xnor U20087 (N_20087,N_18126,N_18806);
nor U20088 (N_20088,N_19929,N_19707);
nand U20089 (N_20089,N_19000,N_18514);
xnor U20090 (N_20090,N_18369,N_19374);
and U20091 (N_20091,N_19593,N_19854);
or U20092 (N_20092,N_18548,N_18880);
and U20093 (N_20093,N_19980,N_19617);
or U20094 (N_20094,N_19612,N_19899);
or U20095 (N_20095,N_18841,N_19969);
nand U20096 (N_20096,N_19503,N_17734);
nand U20097 (N_20097,N_18018,N_19709);
or U20098 (N_20098,N_18512,N_17555);
nor U20099 (N_20099,N_17537,N_17736);
nand U20100 (N_20100,N_17680,N_19309);
or U20101 (N_20101,N_19413,N_18752);
nand U20102 (N_20102,N_17908,N_19550);
xor U20103 (N_20103,N_19415,N_19527);
nand U20104 (N_20104,N_19046,N_18086);
nand U20105 (N_20105,N_19042,N_18106);
xnor U20106 (N_20106,N_19850,N_19486);
nor U20107 (N_20107,N_17586,N_19563);
nand U20108 (N_20108,N_17929,N_19875);
nor U20109 (N_20109,N_19712,N_17797);
and U20110 (N_20110,N_18282,N_19820);
nand U20111 (N_20111,N_17509,N_17521);
or U20112 (N_20112,N_17972,N_17704);
and U20113 (N_20113,N_17759,N_18774);
nor U20114 (N_20114,N_19178,N_17579);
and U20115 (N_20115,N_19485,N_18861);
nand U20116 (N_20116,N_19414,N_19897);
nor U20117 (N_20117,N_18189,N_18476);
and U20118 (N_20118,N_19343,N_18849);
and U20119 (N_20119,N_17958,N_19821);
and U20120 (N_20120,N_19892,N_19446);
or U20121 (N_20121,N_18959,N_17522);
nor U20122 (N_20122,N_19144,N_17510);
or U20123 (N_20123,N_17828,N_17590);
nand U20124 (N_20124,N_18711,N_19494);
nor U20125 (N_20125,N_18687,N_19439);
and U20126 (N_20126,N_18580,N_17993);
xnor U20127 (N_20127,N_19238,N_18493);
and U20128 (N_20128,N_19680,N_18001);
nor U20129 (N_20129,N_19641,N_19373);
nand U20130 (N_20130,N_18228,N_18617);
and U20131 (N_20131,N_19719,N_18153);
nor U20132 (N_20132,N_19429,N_19692);
xnor U20133 (N_20133,N_17733,N_19504);
nor U20134 (N_20134,N_19204,N_17868);
nor U20135 (N_20135,N_18993,N_19614);
xnor U20136 (N_20136,N_18344,N_17784);
xor U20137 (N_20137,N_18052,N_19728);
nand U20138 (N_20138,N_19254,N_18283);
nor U20139 (N_20139,N_18340,N_18649);
or U20140 (N_20140,N_18664,N_18685);
nor U20141 (N_20141,N_19530,N_17569);
nand U20142 (N_20142,N_19147,N_18786);
nor U20143 (N_20143,N_17727,N_18310);
nand U20144 (N_20144,N_19055,N_19973);
nand U20145 (N_20145,N_18480,N_18863);
nor U20146 (N_20146,N_19484,N_17755);
and U20147 (N_20147,N_17557,N_18700);
and U20148 (N_20148,N_18903,N_17843);
and U20149 (N_20149,N_19467,N_19252);
nor U20150 (N_20150,N_17792,N_19979);
nand U20151 (N_20151,N_19726,N_18139);
or U20152 (N_20152,N_17602,N_18976);
and U20153 (N_20153,N_18837,N_18392);
or U20154 (N_20154,N_19776,N_19516);
and U20155 (N_20155,N_18504,N_18789);
xor U20156 (N_20156,N_17694,N_19078);
xnor U20157 (N_20157,N_18808,N_19885);
nand U20158 (N_20158,N_19566,N_17740);
and U20159 (N_20159,N_19790,N_18773);
nand U20160 (N_20160,N_18611,N_18408);
nand U20161 (N_20161,N_18437,N_18822);
and U20162 (N_20162,N_18364,N_17977);
xnor U20163 (N_20163,N_19737,N_18980);
nand U20164 (N_20164,N_18305,N_17990);
nand U20165 (N_20165,N_17833,N_18130);
or U20166 (N_20166,N_19941,N_19587);
or U20167 (N_20167,N_19121,N_17853);
nand U20168 (N_20168,N_19035,N_17523);
nor U20169 (N_20169,N_19529,N_18356);
xor U20170 (N_20170,N_18569,N_19882);
nand U20171 (N_20171,N_18137,N_19592);
xnor U20172 (N_20172,N_18075,N_18761);
or U20173 (N_20173,N_19193,N_18198);
and U20174 (N_20174,N_18951,N_17830);
and U20175 (N_20175,N_17910,N_18393);
nand U20176 (N_20176,N_17572,N_19340);
xor U20177 (N_20177,N_18246,N_19381);
nand U20178 (N_20178,N_17931,N_18059);
nand U20179 (N_20179,N_17739,N_18798);
nor U20180 (N_20180,N_19630,N_19347);
nand U20181 (N_20181,N_19456,N_19827);
xnor U20182 (N_20182,N_17546,N_19830);
and U20183 (N_20183,N_18571,N_17944);
nand U20184 (N_20184,N_19064,N_17532);
or U20185 (N_20185,N_19893,N_19971);
nand U20186 (N_20186,N_19924,N_19358);
xnor U20187 (N_20187,N_18309,N_18438);
or U20188 (N_20188,N_19359,N_19319);
xnor U20189 (N_20189,N_19754,N_17789);
and U20190 (N_20190,N_19155,N_18602);
nand U20191 (N_20191,N_17779,N_19277);
xnor U20192 (N_20192,N_17631,N_17531);
xor U20193 (N_20193,N_17939,N_18695);
and U20194 (N_20194,N_18264,N_18030);
and U20195 (N_20195,N_18620,N_17541);
or U20196 (N_20196,N_19307,N_19874);
xor U20197 (N_20197,N_19202,N_19765);
nand U20198 (N_20198,N_19713,N_18598);
and U20199 (N_20199,N_18091,N_19225);
nor U20200 (N_20200,N_17777,N_17539);
nor U20201 (N_20201,N_19859,N_17534);
and U20202 (N_20202,N_19896,N_17641);
and U20203 (N_20203,N_18521,N_18636);
nand U20204 (N_20204,N_18445,N_18259);
nor U20205 (N_20205,N_17508,N_18832);
xnor U20206 (N_20206,N_18079,N_17743);
xnor U20207 (N_20207,N_18591,N_18082);
xor U20208 (N_20208,N_19888,N_18922);
nor U20209 (N_20209,N_18901,N_18730);
nand U20210 (N_20210,N_19634,N_18204);
nor U20211 (N_20211,N_17793,N_18164);
xor U20212 (N_20212,N_17568,N_17620);
nand U20213 (N_20213,N_19767,N_17750);
and U20214 (N_20214,N_17947,N_18988);
and U20215 (N_20215,N_19234,N_18316);
xor U20216 (N_20216,N_17699,N_18683);
and U20217 (N_20217,N_18574,N_19366);
or U20218 (N_20218,N_18399,N_19600);
nand U20219 (N_20219,N_18037,N_19557);
xor U20220 (N_20220,N_19598,N_17927);
or U20221 (N_20221,N_19295,N_17979);
or U20222 (N_20222,N_17924,N_19135);
nand U20223 (N_20223,N_19743,N_19293);
and U20224 (N_20224,N_18462,N_18920);
xnor U20225 (N_20225,N_18121,N_19001);
nand U20226 (N_20226,N_18589,N_19913);
or U20227 (N_20227,N_17761,N_18058);
and U20228 (N_20228,N_17670,N_18296);
or U20229 (N_20229,N_19750,N_19561);
xnor U20230 (N_20230,N_19338,N_17864);
nor U20231 (N_20231,N_19165,N_18339);
and U20232 (N_20232,N_18517,N_17989);
xnor U20233 (N_20233,N_18766,N_18811);
and U20234 (N_20234,N_18900,N_19968);
nand U20235 (N_20235,N_18085,N_18788);
nand U20236 (N_20236,N_18163,N_18178);
xnor U20237 (N_20237,N_18904,N_19390);
and U20238 (N_20238,N_18824,N_19879);
and U20239 (N_20239,N_19900,N_17693);
or U20240 (N_20240,N_19756,N_18314);
nor U20241 (N_20241,N_17511,N_18308);
or U20242 (N_20242,N_18835,N_18956);
nor U20243 (N_20243,N_18908,N_18307);
nor U20244 (N_20244,N_19610,N_18974);
xor U20245 (N_20245,N_18884,N_17858);
and U20246 (N_20246,N_19257,N_19872);
xnor U20247 (N_20247,N_19436,N_19585);
and U20248 (N_20248,N_18674,N_18734);
and U20249 (N_20249,N_18536,N_17506);
or U20250 (N_20250,N_19985,N_19442);
nand U20251 (N_20251,N_19517,N_18600);
nor U20252 (N_20252,N_18796,N_19944);
nand U20253 (N_20253,N_19423,N_19231);
nor U20254 (N_20254,N_17603,N_18120);
nor U20255 (N_20255,N_18732,N_19017);
xnor U20256 (N_20256,N_19596,N_19542);
and U20257 (N_20257,N_18220,N_19060);
nor U20258 (N_20258,N_18096,N_17664);
or U20259 (N_20259,N_18345,N_17849);
nand U20260 (N_20260,N_17562,N_17650);
and U20261 (N_20261,N_18293,N_17847);
nand U20262 (N_20262,N_19161,N_19722);
or U20263 (N_20263,N_18949,N_19597);
and U20264 (N_20264,N_18576,N_19117);
nand U20265 (N_20265,N_19488,N_17881);
or U20266 (N_20266,N_17945,N_18994);
or U20267 (N_20267,N_18686,N_18325);
or U20268 (N_20268,N_19301,N_19141);
and U20269 (N_20269,N_19648,N_19190);
nand U20270 (N_20270,N_17553,N_19316);
nor U20271 (N_20271,N_18699,N_18913);
nand U20272 (N_20272,N_17940,N_19966);
or U20273 (N_20273,N_19502,N_19438);
or U20274 (N_20274,N_18520,N_18579);
nand U20275 (N_20275,N_18644,N_19463);
xor U20276 (N_20276,N_19590,N_18754);
nor U20277 (N_20277,N_19235,N_19520);
nand U20278 (N_20278,N_18171,N_17854);
xnor U20279 (N_20279,N_18528,N_17985);
nor U20280 (N_20280,N_19051,N_18847);
nor U20281 (N_20281,N_19412,N_19922);
nor U20282 (N_20282,N_18216,N_19349);
nand U20283 (N_20283,N_19644,N_19156);
or U20284 (N_20284,N_17995,N_18374);
xor U20285 (N_20285,N_17961,N_17500);
nand U20286 (N_20286,N_19740,N_18329);
or U20287 (N_20287,N_19724,N_19250);
nor U20288 (N_20288,N_19365,N_19173);
nand U20289 (N_20289,N_18971,N_18247);
and U20290 (N_20290,N_17883,N_18691);
xnor U20291 (N_20291,N_17685,N_17794);
and U20292 (N_20292,N_19703,N_19096);
nand U20293 (N_20293,N_17869,N_19321);
and U20294 (N_20294,N_17712,N_18353);
nor U20295 (N_20295,N_19615,N_17630);
xnor U20296 (N_20296,N_19021,N_18161);
and U20297 (N_20297,N_18542,N_18759);
nor U20298 (N_20298,N_17809,N_19552);
xor U20299 (N_20299,N_19411,N_18193);
and U20300 (N_20300,N_18113,N_19746);
nor U20301 (N_20301,N_17676,N_18721);
nor U20302 (N_20302,N_19408,N_19873);
nor U20303 (N_20303,N_19531,N_18361);
nor U20304 (N_20304,N_18578,N_18475);
nand U20305 (N_20305,N_19196,N_18234);
nand U20306 (N_20306,N_18658,N_18545);
or U20307 (N_20307,N_18455,N_18078);
xnor U20308 (N_20308,N_18899,N_19669);
xnor U20309 (N_20309,N_19080,N_19731);
nor U20310 (N_20310,N_19914,N_18494);
or U20311 (N_20311,N_19246,N_19554);
nand U20312 (N_20312,N_18370,N_19472);
nor U20313 (N_20313,N_19940,N_19894);
nor U20314 (N_20314,N_18253,N_18823);
nand U20315 (N_20315,N_18122,N_19163);
nand U20316 (N_20316,N_17515,N_19714);
or U20317 (N_20317,N_19229,N_17760);
or U20318 (N_20318,N_18488,N_17719);
xor U20319 (N_20319,N_19222,N_19668);
nand U20320 (N_20320,N_19212,N_18505);
xnor U20321 (N_20321,N_19528,N_17971);
and U20322 (N_20322,N_17618,N_19586);
or U20323 (N_20323,N_17896,N_19673);
and U20324 (N_20324,N_17976,N_19526);
and U20325 (N_20325,N_18114,N_18021);
or U20326 (N_20326,N_19793,N_19342);
xnor U20327 (N_20327,N_18990,N_18817);
or U20328 (N_20328,N_19255,N_18626);
or U20329 (N_20329,N_19032,N_19864);
and U20330 (N_20330,N_18894,N_18472);
nand U20331 (N_20331,N_17730,N_19549);
xor U20332 (N_20332,N_18805,N_19510);
xnor U20333 (N_20333,N_18815,N_18775);
nor U20334 (N_20334,N_17963,N_19379);
or U20335 (N_20335,N_17932,N_18124);
and U20336 (N_20336,N_17624,N_19346);
nand U20337 (N_20337,N_17965,N_18983);
nand U20338 (N_20338,N_19727,N_19868);
nor U20339 (N_20339,N_19534,N_18735);
nand U20340 (N_20340,N_19514,N_17633);
xnor U20341 (N_20341,N_17874,N_18014);
xnor U20342 (N_20342,N_18939,N_17707);
or U20343 (N_20343,N_19997,N_17870);
or U20344 (N_20344,N_18035,N_19243);
and U20345 (N_20345,N_19133,N_18145);
nor U20346 (N_20346,N_17758,N_19666);
or U20347 (N_20347,N_17970,N_19902);
or U20348 (N_20348,N_17502,N_18601);
nand U20349 (N_20349,N_17623,N_19143);
xnor U20350 (N_20350,N_18042,N_18909);
or U20351 (N_20351,N_18332,N_19704);
nand U20352 (N_20352,N_18336,N_17974);
and U20353 (N_20353,N_17529,N_19258);
and U20354 (N_20354,N_19609,N_17518);
and U20355 (N_20355,N_18905,N_18200);
xor U20356 (N_20356,N_19251,N_18785);
or U20357 (N_20357,N_19524,N_19434);
xnor U20358 (N_20358,N_17720,N_19285);
xnor U20359 (N_20359,N_17613,N_18303);
or U20360 (N_20360,N_17710,N_18524);
nor U20361 (N_20361,N_18214,N_19419);
nor U20362 (N_20362,N_18388,N_17629);
nor U20363 (N_20363,N_18099,N_18655);
xor U20364 (N_20364,N_18288,N_18398);
xnor U20365 (N_20365,N_18666,N_19210);
or U20366 (N_20366,N_19927,N_18485);
and U20367 (N_20367,N_19620,N_18298);
nor U20368 (N_20368,N_18040,N_17735);
nand U20369 (N_20369,N_19091,N_18346);
or U20370 (N_20370,N_18450,N_17879);
and U20371 (N_20371,N_18004,N_19539);
or U20372 (N_20372,N_19013,N_17818);
nand U20373 (N_20373,N_17914,N_17878);
nand U20374 (N_20374,N_19843,N_18064);
xor U20375 (N_20375,N_18985,N_19742);
or U20376 (N_20376,N_17527,N_18365);
nand U20377 (N_20377,N_18405,N_18175);
or U20378 (N_20378,N_18010,N_17503);
and U20379 (N_20379,N_19833,N_18709);
nor U20380 (N_20380,N_18304,N_19705);
nand U20381 (N_20381,N_19856,N_17787);
or U20382 (N_20382,N_17536,N_19232);
and U20383 (N_20383,N_19651,N_17839);
nor U20384 (N_20384,N_17667,N_18186);
xnor U20385 (N_20385,N_17721,N_18413);
or U20386 (N_20386,N_17589,N_18201);
nand U20387 (N_20387,N_17612,N_18914);
xor U20388 (N_20388,N_17848,N_18714);
nor U20389 (N_20389,N_18779,N_17773);
or U20390 (N_20390,N_18128,N_19569);
nor U20391 (N_20391,N_18511,N_18481);
or U20392 (N_20392,N_18673,N_18727);
and U20393 (N_20393,N_18891,N_19282);
nor U20394 (N_20394,N_17997,N_18782);
or U20395 (N_20395,N_19890,N_18454);
or U20396 (N_20396,N_18898,N_18395);
xor U20397 (N_20397,N_19523,N_19236);
xor U20398 (N_20398,N_17892,N_19533);
nand U20399 (N_20399,N_19082,N_19266);
nand U20400 (N_20400,N_19410,N_19399);
nor U20401 (N_20401,N_18522,N_19912);
nand U20402 (N_20402,N_19142,N_19123);
and U20403 (N_20403,N_17614,N_17913);
xnor U20404 (N_20404,N_18751,N_18072);
nand U20405 (N_20405,N_18003,N_19109);
or U20406 (N_20406,N_18379,N_19352);
nand U20407 (N_20407,N_18606,N_18838);
xnor U20408 (N_20408,N_19331,N_19345);
nor U20409 (N_20409,N_19093,N_19946);
nor U20410 (N_20410,N_19140,N_19393);
nand U20411 (N_20411,N_18243,N_19448);
or U20412 (N_20412,N_18912,N_19807);
xor U20413 (N_20413,N_17814,N_19437);
and U20414 (N_20414,N_19395,N_18515);
and U20415 (N_20415,N_18769,N_18396);
xor U20416 (N_20416,N_17996,N_18150);
nor U20417 (N_20417,N_18292,N_19329);
or U20418 (N_20418,N_18378,N_19601);
nand U20419 (N_20419,N_18151,N_19676);
and U20420 (N_20420,N_18301,N_19525);
nand U20421 (N_20421,N_18705,N_18770);
and U20422 (N_20422,N_18302,N_18783);
nor U20423 (N_20423,N_19385,N_18337);
and U20424 (N_20424,N_18473,N_17824);
or U20425 (N_20425,N_18795,N_18158);
xor U20426 (N_20426,N_19487,N_19150);
xor U20427 (N_20427,N_18311,N_19454);
and U20428 (N_20428,N_17836,N_18746);
nor U20429 (N_20429,N_17655,N_17657);
and U20430 (N_20430,N_17808,N_17756);
xnor U20431 (N_20431,N_18237,N_18400);
and U20432 (N_20432,N_19752,N_19811);
nand U20433 (N_20433,N_17634,N_17695);
nand U20434 (N_20434,N_19594,N_19988);
nor U20435 (N_20435,N_19240,N_17862);
nor U20436 (N_20436,N_19054,N_19970);
nand U20437 (N_20437,N_17648,N_19747);
xnor U20438 (N_20438,N_19824,N_18516);
xnor U20439 (N_20439,N_19662,N_19447);
or U20440 (N_20440,N_18871,N_18827);
or U20441 (N_20441,N_17876,N_18453);
xnor U20442 (N_20442,N_18597,N_19443);
and U20443 (N_20443,N_18757,N_17742);
and U20444 (N_20444,N_18722,N_19482);
xnor U20445 (N_20445,N_18945,N_19172);
nand U20446 (N_20446,N_18236,N_18947);
xnor U20447 (N_20447,N_17900,N_18692);
nor U20448 (N_20448,N_17576,N_17949);
and U20449 (N_20449,N_19547,N_19270);
nor U20450 (N_20450,N_19402,N_18338);
nand U20451 (N_20451,N_19195,N_19819);
or U20452 (N_20452,N_19672,N_18431);
xnor U20453 (N_20453,N_19087,N_17852);
nor U20454 (N_20454,N_18508,N_18991);
and U20455 (N_20455,N_19268,N_18581);
nor U20456 (N_20456,N_17538,N_18351);
or U20457 (N_20457,N_19640,N_19421);
or U20458 (N_20458,N_18168,N_17807);
or U20459 (N_20459,N_18412,N_18132);
or U20460 (N_20460,N_18501,N_19160);
xor U20461 (N_20461,N_18170,N_18510);
nor U20462 (N_20462,N_18704,N_18474);
xor U20463 (N_20463,N_17860,N_18519);
and U20464 (N_20464,N_17841,N_18169);
nor U20465 (N_20465,N_18491,N_18466);
nor U20466 (N_20466,N_19066,N_17980);
xor U20467 (N_20467,N_19044,N_18530);
nand U20468 (N_20468,N_17955,N_19088);
nand U20469 (N_20469,N_19388,N_18270);
nand U20470 (N_20470,N_18109,N_18724);
xor U20471 (N_20471,N_19543,N_19702);
xnor U20472 (N_20472,N_17526,N_18816);
xor U20473 (N_20473,N_18140,N_19101);
or U20474 (N_20474,N_17686,N_18544);
nor U20475 (N_20475,N_18743,N_18420);
or U20476 (N_20476,N_19753,N_19787);
and U20477 (N_20477,N_18286,N_19397);
xor U20478 (N_20478,N_17942,N_18561);
or U20479 (N_20479,N_17565,N_19720);
and U20480 (N_20480,N_18818,N_18324);
or U20481 (N_20481,N_18103,N_19430);
nand U20482 (N_20482,N_19920,N_19336);
or U20483 (N_20483,N_19134,N_17838);
and U20484 (N_20484,N_19921,N_18219);
nand U20485 (N_20485,N_18289,N_19813);
nand U20486 (N_20486,N_17651,N_19848);
xor U20487 (N_20487,N_18469,N_17956);
nor U20488 (N_20488,N_17925,N_18953);
nor U20489 (N_20489,N_19223,N_18423);
nor U20490 (N_20490,N_18208,N_19732);
xnor U20491 (N_20491,N_18240,N_17654);
and U20492 (N_20492,N_19356,N_19845);
nor U20493 (N_20493,N_18486,N_18639);
and U20494 (N_20494,N_19009,N_19809);
nor U20495 (N_20495,N_18842,N_19466);
or U20496 (N_20496,N_18389,N_18933);
nand U20497 (N_20497,N_17857,N_19010);
and U20498 (N_20498,N_19224,N_18287);
and U20499 (N_20499,N_18192,N_19559);
and U20500 (N_20500,N_18593,N_18513);
and U20501 (N_20501,N_18294,N_19305);
nor U20502 (N_20502,N_17550,N_19908);
nand U20503 (N_20503,N_18467,N_17933);
or U20504 (N_20504,N_18005,N_19977);
and U20505 (N_20505,N_18007,N_19097);
xor U20506 (N_20506,N_19943,N_18230);
or U20507 (N_20507,N_19170,N_18931);
nand U20508 (N_20508,N_18184,N_18411);
nand U20509 (N_20509,N_19216,N_19084);
and U20510 (N_20510,N_19961,N_19567);
or U20511 (N_20511,N_19361,N_19215);
and U20512 (N_20512,N_19057,N_18634);
or U20513 (N_20513,N_19325,N_18652);
nor U20514 (N_20514,N_19136,N_18726);
and U20515 (N_20515,N_18222,N_18879);
nor U20516 (N_20516,N_17520,N_18738);
nor U20517 (N_20517,N_19842,N_17722);
xnor U20518 (N_20518,N_19296,N_19611);
xnor U20519 (N_20519,N_18657,N_17595);
xor U20520 (N_20520,N_18382,N_19878);
nand U20521 (N_20521,N_18129,N_17938);
or U20522 (N_20522,N_19694,N_18651);
nor U20523 (N_20523,N_19128,N_17563);
xor U20524 (N_20524,N_19544,N_17501);
or U20525 (N_20525,N_19061,N_19952);
xor U20526 (N_20526,N_18996,N_18720);
and U20527 (N_20527,N_18094,N_19930);
nor U20528 (N_20528,N_17764,N_18185);
xor U20529 (N_20529,N_19377,N_18367);
or U20530 (N_20530,N_19476,N_17585);
nor U20531 (N_20531,N_19118,N_18526);
nand U20532 (N_20532,N_18343,N_18147);
nor U20533 (N_20533,N_18758,N_18987);
nor U20534 (N_20534,N_19558,N_18633);
xor U20535 (N_20535,N_18554,N_19717);
and U20536 (N_20536,N_17672,N_17951);
and U20537 (N_20537,N_17598,N_18057);
nand U20538 (N_20538,N_17850,N_19099);
nand U20539 (N_20539,N_19233,N_19465);
and U20540 (N_20540,N_19992,N_18853);
nand U20541 (N_20541,N_18409,N_18209);
nor U20542 (N_20542,N_19916,N_17834);
nor U20543 (N_20543,N_17746,N_18549);
or U20544 (N_20544,N_17765,N_18183);
nand U20545 (N_20545,N_17726,N_18925);
and U20546 (N_20546,N_18349,N_18048);
xor U20547 (N_20547,N_19923,N_18717);
and U20548 (N_20548,N_18856,N_17702);
or U20549 (N_20549,N_17816,N_18242);
and U20550 (N_20550,N_17690,N_18123);
or U20551 (N_20551,N_19267,N_19621);
or U20552 (N_20552,N_19079,N_19891);
and U20553 (N_20553,N_18596,N_19877);
and U20554 (N_20554,N_19942,N_19288);
or U20555 (N_20555,N_18745,N_19623);
nand U20556 (N_20556,N_18981,N_17917);
and U20557 (N_20557,N_17635,N_18946);
nor U20558 (N_20558,N_19624,N_19176);
and U20559 (N_20559,N_18254,N_18723);
xnor U20560 (N_20560,N_19786,N_17802);
and U20561 (N_20561,N_19679,N_17600);
and U20562 (N_20562,N_19541,N_18321);
xnor U20563 (N_20563,N_18152,N_19622);
nor U20564 (N_20564,N_18276,N_19158);
or U20565 (N_20565,N_19367,N_18257);
nor U20566 (N_20566,N_18056,N_19322);
nand U20567 (N_20567,N_19433,N_18299);
or U20568 (N_20568,N_19249,N_19314);
xor U20569 (N_20569,N_18366,N_19209);
or U20570 (N_20570,N_17903,N_17825);
xnor U20571 (N_20571,N_19124,N_19667);
nand U20572 (N_20572,N_18223,N_17622);
nand U20573 (N_20573,N_17716,N_18013);
nor U20574 (N_20574,N_18826,N_18471);
nand U20575 (N_20575,N_17535,N_19284);
nor U20576 (N_20576,N_18235,N_19337);
xnor U20577 (N_20577,N_17645,N_18793);
and U20578 (N_20578,N_19248,N_18962);
xor U20579 (N_20579,N_19805,N_18317);
xnor U20580 (N_20580,N_18877,N_18105);
or U20581 (N_20581,N_18932,N_19218);
and U20582 (N_20582,N_19886,N_17751);
nor U20583 (N_20583,N_17582,N_17986);
nor U20584 (N_20584,N_19050,N_19764);
xor U20585 (N_20585,N_17813,N_19116);
or U20586 (N_20586,N_18964,N_18679);
or U20587 (N_20587,N_18537,N_18958);
nand U20588 (N_20588,N_19500,N_19828);
and U20589 (N_20589,N_17678,N_19449);
and U20590 (N_20590,N_18961,N_17855);
or U20591 (N_20591,N_18268,N_19028);
and U20592 (N_20592,N_19005,N_18930);
nor U20593 (N_20593,N_18110,N_18889);
or U20594 (N_20594,N_19418,N_17873);
nand U20595 (N_20595,N_18669,N_19876);
or U20596 (N_20596,N_17658,N_19303);
nor U20597 (N_20597,N_18046,N_19175);
nand U20598 (N_20598,N_17821,N_17588);
or U20599 (N_20599,N_19300,N_18028);
nand U20600 (N_20600,N_18433,N_19326);
nand U20601 (N_20601,N_18851,N_18375);
xor U20602 (N_20602,N_19431,N_18538);
xnor U20603 (N_20603,N_18277,N_19945);
xnor U20604 (N_20604,N_19862,N_19221);
nand U20605 (N_20605,N_18134,N_18509);
nor U20606 (N_20606,N_19462,N_18443);
or U20607 (N_20607,N_18448,N_19846);
xor U20608 (N_20608,N_18115,N_19901);
xnor U20609 (N_20609,N_19665,N_19403);
or U20610 (N_20610,N_19555,N_18002);
nand U20611 (N_20611,N_19495,N_17856);
xor U20612 (N_20612,N_19371,N_19847);
and U20613 (N_20613,N_19652,N_18756);
nor U20614 (N_20614,N_19518,N_19461);
xor U20615 (N_20615,N_18881,N_18897);
or U20616 (N_20616,N_19422,N_18074);
nand U20617 (N_20617,N_18998,N_18618);
and U20618 (N_20618,N_18155,N_18529);
xor U20619 (N_20619,N_18802,N_18982);
xor U20620 (N_20620,N_19451,N_17519);
or U20621 (N_20621,N_18207,N_19259);
and U20622 (N_20622,N_19265,N_17992);
nand U20623 (N_20623,N_18763,N_19291);
or U20624 (N_20624,N_18857,N_18281);
nand U20625 (N_20625,N_19745,N_19432);
xor U20626 (N_20626,N_19405,N_17513);
and U20627 (N_20627,N_18363,N_19884);
nor U20628 (N_20628,N_19211,N_18008);
and U20629 (N_20629,N_17796,N_19791);
or U20630 (N_20630,N_18954,N_19536);
xnor U20631 (N_20631,N_17916,N_17866);
nor U20632 (N_20632,N_19004,N_19089);
nand U20633 (N_20633,N_19762,N_18027);
xnor U20634 (N_20634,N_17610,N_18065);
or U20635 (N_20635,N_17647,N_19866);
or U20636 (N_20636,N_18421,N_17935);
nor U20637 (N_20637,N_18404,N_18499);
and U20638 (N_20638,N_18012,N_18320);
or U20639 (N_20639,N_19048,N_19453);
and U20640 (N_20640,N_18921,N_18646);
xnor U20641 (N_20641,N_18261,N_18659);
and U20642 (N_20642,N_19480,N_19110);
nand U20643 (N_20643,N_17752,N_19479);
nand U20644 (N_20644,N_17627,N_18190);
and U20645 (N_20645,N_18138,N_19625);
nor U20646 (N_20646,N_19368,N_19386);
and U20647 (N_20647,N_18019,N_18800);
or U20648 (N_20648,N_19605,N_19650);
nand U20649 (N_20649,N_19616,N_19145);
and U20650 (N_20650,N_18926,N_18348);
nor U20651 (N_20651,N_19049,N_18249);
nand U20652 (N_20652,N_19260,N_18410);
and U20653 (N_20653,N_18866,N_18747);
nand U20654 (N_20654,N_19782,N_17594);
and U20655 (N_20655,N_19025,N_19299);
nor U20656 (N_20656,N_18258,N_17540);
and U20657 (N_20657,N_17835,N_18553);
and U20658 (N_20658,N_17728,N_19655);
or U20659 (N_20659,N_18141,N_18352);
nand U20660 (N_20660,N_18650,N_17659);
nand U20661 (N_20661,N_19425,N_18432);
nor U20662 (N_20662,N_19656,N_19007);
or U20663 (N_20663,N_17905,N_18070);
and U20664 (N_20664,N_18506,N_17926);
or U20665 (N_20665,N_19058,N_19280);
and U20666 (N_20666,N_19792,N_18564);
xnor U20667 (N_20667,N_17748,N_19795);
xnor U20668 (N_20668,N_19398,N_19294);
nor U20669 (N_20669,N_19029,N_18381);
and U20670 (N_20670,N_18330,N_17573);
nand U20671 (N_20671,N_19955,N_19459);
and U20672 (N_20672,N_19507,N_19926);
xor U20673 (N_20673,N_18801,N_19682);
nor U20674 (N_20674,N_18133,N_18221);
and U20675 (N_20675,N_19244,N_17525);
nand U20676 (N_20676,N_18239,N_18621);
nand U20677 (N_20677,N_19853,N_18638);
or U20678 (N_20678,N_17786,N_18869);
or U20679 (N_20679,N_19681,N_17713);
nor U20680 (N_20680,N_19445,N_18794);
xnor U20681 (N_20681,N_18780,N_19174);
xor U20682 (N_20682,N_19928,N_19287);
nor U20683 (N_20683,N_19789,N_18458);
nand U20684 (N_20684,N_19967,N_18023);
xor U20685 (N_20685,N_19041,N_19318);
xor U20686 (N_20686,N_18119,N_17799);
nand U20687 (N_20687,N_19308,N_19636);
xor U20688 (N_20688,N_17911,N_17593);
nor U20689 (N_20689,N_18972,N_18797);
or U20690 (N_20690,N_17663,N_19330);
xor U20691 (N_20691,N_18360,N_19595);
nor U20692 (N_20692,N_18265,N_18690);
nor U20693 (N_20693,N_19126,N_19841);
nand U20694 (N_20694,N_17625,N_17882);
or U20695 (N_20695,N_17566,N_19217);
nand U20696 (N_20696,N_18551,N_17656);
and U20697 (N_20697,N_18326,N_17583);
and U20698 (N_20698,N_18765,N_19111);
or U20699 (N_20699,N_18595,N_19450);
nand U20700 (N_20700,N_18854,N_19629);
or U20701 (N_20701,N_17988,N_19286);
nand U20702 (N_20702,N_17596,N_17774);
or U20703 (N_20703,N_18825,N_19213);
xor U20704 (N_20704,N_18627,N_17718);
xnor U20705 (N_20705,N_17581,N_18728);
xnor U20706 (N_20706,N_19455,N_17564);
and U20707 (N_20707,N_18846,N_19687);
or U20708 (N_20708,N_19766,N_18665);
and U20709 (N_20709,N_18495,N_19376);
nor U20710 (N_20710,N_19324,N_18436);
and U20711 (N_20711,N_17895,N_19718);
nor U20712 (N_20712,N_19870,N_18858);
or U20713 (N_20713,N_18442,N_19157);
nor U20714 (N_20714,N_17768,N_17616);
and U20715 (N_20715,N_19607,N_18341);
nand U20716 (N_20716,N_18084,N_17548);
and U20717 (N_20717,N_19199,N_19253);
nor U20718 (N_20718,N_17884,N_19580);
and U20719 (N_20719,N_18768,N_19691);
xnor U20720 (N_20720,N_18915,N_18662);
and U20721 (N_20721,N_18011,N_18179);
nor U20722 (N_20722,N_18927,N_19417);
nand U20723 (N_20723,N_19104,N_17599);
or U20724 (N_20724,N_18619,N_18229);
or U20725 (N_20725,N_18590,N_19794);
and U20726 (N_20726,N_19643,N_17660);
and U20727 (N_20727,N_18449,N_19306);
nor U20728 (N_20728,N_18960,N_18444);
or U20729 (N_20729,N_17987,N_18870);
nand U20730 (N_20730,N_18592,N_18850);
nor U20731 (N_20731,N_19706,N_19986);
nand U20732 (N_20732,N_18496,N_19263);
xor U20733 (N_20733,N_17781,N_19822);
nor U20734 (N_20734,N_17507,N_19695);
or U20735 (N_20735,N_17675,N_18907);
nor U20736 (N_20736,N_18605,N_17845);
and U20737 (N_20737,N_19184,N_17805);
or U20738 (N_20738,N_19576,N_18044);
nand U20739 (N_20739,N_19741,N_17689);
and U20740 (N_20740,N_19604,N_17766);
nand U20741 (N_20741,N_17918,N_18563);
and U20742 (N_20742,N_18387,N_17617);
or U20743 (N_20743,N_18781,N_18372);
nor U20744 (N_20744,N_19700,N_17763);
or U20745 (N_20745,N_17894,N_17731);
or U20746 (N_20746,N_17782,N_19380);
xnor U20747 (N_20747,N_17517,N_18771);
xnor U20748 (N_20748,N_18359,N_17644);
nand U20749 (N_20749,N_17897,N_18539);
nor U20750 (N_20750,N_17646,N_19056);
xor U20751 (N_20751,N_18741,N_18306);
nand U20752 (N_20752,N_19844,N_17902);
and U20753 (N_20753,N_18997,N_17597);
nand U20754 (N_20754,N_18402,N_18682);
xor U20755 (N_20755,N_19570,N_17558);
and U20756 (N_20756,N_18678,N_19107);
or U20757 (N_20757,N_19063,N_19774);
nor U20758 (N_20758,N_19581,N_18087);
nand U20759 (N_20759,N_18295,N_18354);
and U20760 (N_20760,N_18117,N_18830);
nand U20761 (N_20761,N_18582,N_18090);
nand U20762 (N_20762,N_18635,N_19812);
or U20763 (N_20763,N_18016,N_19759);
xor U20764 (N_20764,N_19663,N_19857);
and U20765 (N_20765,N_19100,N_19383);
nand U20766 (N_20766,N_19932,N_17778);
xor U20767 (N_20767,N_19579,N_19491);
nand U20768 (N_20768,N_18224,N_19810);
or U20769 (N_20769,N_18572,N_18160);
xor U20770 (N_20770,N_17851,N_18350);
nand U20771 (N_20771,N_17937,N_19645);
xor U20772 (N_20772,N_18637,N_18910);
nand U20773 (N_20773,N_19186,N_19505);
and U20774 (N_20774,N_19113,N_19490);
nor U20775 (N_20775,N_19633,N_18531);
nand U20776 (N_20776,N_19816,N_18577);
or U20777 (N_20777,N_17822,N_19670);
and U20778 (N_20778,N_19906,N_19957);
and U20779 (N_20779,N_19990,N_17674);
xor U20780 (N_20780,N_18565,N_19936);
or U20781 (N_20781,N_17798,N_18562);
xor U20782 (N_20782,N_19721,N_19310);
nor U20783 (N_20783,N_18439,N_18896);
or U20784 (N_20784,N_17549,N_18567);
nand U20785 (N_20785,N_17861,N_18725);
or U20786 (N_20786,N_18570,N_19778);
xor U20787 (N_20787,N_17609,N_18948);
xor U20788 (N_20788,N_19698,N_19389);
nor U20789 (N_20789,N_19274,N_19799);
xnor U20790 (N_20790,N_19637,N_18556);
nand U20791 (N_20791,N_19798,N_17891);
xor U20792 (N_20792,N_19887,N_19683);
or U20793 (N_20793,N_19311,N_19355);
xnor U20794 (N_20794,N_19736,N_18989);
xor U20795 (N_20795,N_19372,N_18291);
and U20796 (N_20796,N_19991,N_17637);
and U20797 (N_20797,N_17984,N_17886);
nor U20798 (N_20798,N_18663,N_19839);
or U20799 (N_20799,N_18940,N_19638);
or U20800 (N_20800,N_18715,N_19513);
nand U20801 (N_20801,N_18104,N_19574);
xnor U20802 (N_20802,N_19577,N_18333);
nor U20803 (N_20803,N_19826,N_17888);
xnor U20804 (N_20804,N_19735,N_17543);
or U20805 (N_20805,N_17640,N_19723);
nand U20806 (N_20806,N_19441,N_17804);
and U20807 (N_20807,N_18422,N_17810);
xor U20808 (N_20808,N_18088,N_18965);
and U20809 (N_20809,N_18401,N_17776);
nor U20810 (N_20810,N_19496,N_19948);
nand U20811 (N_20811,N_18279,N_17889);
xnor U20812 (N_20812,N_19387,N_18107);
nor U20813 (N_20813,N_18165,N_18452);
nor U20814 (N_20814,N_19477,N_19768);
and U20815 (N_20815,N_18902,N_18862);
nand U20816 (N_20816,N_19642,N_18503);
nor U20817 (N_20817,N_17725,N_19823);
xor U20818 (N_20818,N_18417,N_18478);
nor U20819 (N_20819,N_18446,N_19584);
and U20820 (N_20820,N_19881,N_18039);
nor U20821 (N_20821,N_19085,N_18911);
or U20822 (N_20822,N_17653,N_19200);
or U20823 (N_20823,N_19889,N_17806);
xor U20824 (N_20824,N_17788,N_18045);
and U20825 (N_20825,N_17639,N_19351);
nand U20826 (N_20826,N_17780,N_19708);
or U20827 (N_20827,N_17863,N_18047);
xor U20828 (N_20828,N_17859,N_17605);
nand U20829 (N_20829,N_18188,N_17999);
nand U20830 (N_20830,N_18033,N_19262);
or U20831 (N_20831,N_19825,N_17998);
nor U20832 (N_20832,N_19956,N_19115);
or U20833 (N_20833,N_17865,N_19152);
nand U20834 (N_20834,N_19364,N_19191);
or U20835 (N_20835,N_18656,N_17967);
or U20836 (N_20836,N_18459,N_17757);
nand U20837 (N_20837,N_18583,N_19205);
nor U20838 (N_20838,N_18092,N_19758);
nand U20839 (N_20839,N_18648,N_19473);
and U20840 (N_20840,N_18667,N_17948);
and U20841 (N_20841,N_19304,N_18653);
xnor U20842 (N_20842,N_19919,N_18804);
and U20843 (N_20843,N_18829,N_18108);
nor U20844 (N_20844,N_18083,N_18995);
and U20845 (N_20845,N_19675,N_19038);
nand U20846 (N_20846,N_18893,N_18225);
and U20847 (N_20847,N_19685,N_19092);
or U20848 (N_20848,N_17683,N_18231);
or U20849 (N_20849,N_19458,N_18390);
nand U20850 (N_20850,N_18318,N_18777);
or U20851 (N_20851,N_17567,N_18718);
nor U20852 (N_20852,N_18383,N_18872);
and U20853 (N_20853,N_19016,N_19153);
and U20854 (N_20854,N_19671,N_19239);
nand U20855 (N_20855,N_18712,N_17723);
or U20856 (N_20856,N_17560,N_18876);
nand U20857 (N_20857,N_17652,N_18385);
or U20858 (N_20858,N_18622,N_18285);
nand U20859 (N_20859,N_19852,N_17978);
xor U20860 (N_20860,N_18146,N_18944);
and U20861 (N_20861,N_17673,N_17545);
nand U20862 (N_20862,N_18661,N_18547);
and U20863 (N_20863,N_18689,N_18377);
nand U20864 (N_20864,N_19725,N_19783);
xnor U20865 (N_20865,N_17547,N_19470);
and U20866 (N_20866,N_18919,N_18166);
nand U20867 (N_20867,N_19164,N_18707);
xnor U20868 (N_20868,N_17571,N_19582);
nor U20869 (N_20869,N_19618,N_18942);
and U20870 (N_20870,N_18575,N_18744);
nor U20871 (N_20871,N_19404,N_19788);
xor U20872 (N_20872,N_19965,N_19185);
xnor U20873 (N_20873,N_19072,N_19426);
and U20874 (N_20874,N_19710,N_18251);
nor U20875 (N_20875,N_17829,N_18963);
xor U20876 (N_20876,N_18029,N_19797);
nand U20877 (N_20877,N_19904,N_18820);
and U20878 (N_20878,N_19332,N_18628);
nor U20879 (N_20879,N_19635,N_19120);
and U20880 (N_20880,N_19861,N_18708);
and U20881 (N_20881,N_18697,N_19578);
or U20882 (N_20882,N_19664,N_17701);
and U20883 (N_20883,N_19228,N_18487);
xnor U20884 (N_20884,N_17754,N_18331);
xnor U20885 (N_20885,N_18238,N_19761);
xnor U20886 (N_20886,N_19492,N_17880);
or U20887 (N_20887,N_18233,N_18347);
nand U20888 (N_20888,N_19247,N_19315);
nand U20889 (N_20889,N_19982,N_19909);
nor U20890 (N_20890,N_19976,N_17994);
or U20891 (N_20891,N_19963,N_18440);
or U20892 (N_20892,N_19506,N_17872);
xor U20893 (N_20893,N_18017,N_19951);
nor U20894 (N_20894,N_19139,N_19159);
or U20895 (N_20895,N_19564,N_19498);
and U20896 (N_20896,N_18890,N_19562);
xnor U20897 (N_20897,N_18623,N_18935);
nor U20898 (N_20898,N_18844,N_17554);
or U20899 (N_20899,N_18603,N_18975);
nand U20900 (N_20900,N_18199,N_17920);
nor U20901 (N_20901,N_18191,N_18055);
nor U20902 (N_20902,N_19855,N_17607);
and U20903 (N_20903,N_18319,N_19226);
xnor U20904 (N_20904,N_18525,N_19018);
nand U20905 (N_20905,N_19588,N_18739);
nand U20906 (N_20906,N_18594,N_19696);
nor U20907 (N_20907,N_18368,N_18447);
nor U20908 (N_20908,N_18892,N_19939);
or U20909 (N_20909,N_18878,N_18992);
nand U20910 (N_20910,N_19659,N_19729);
nor U20911 (N_20911,N_18848,N_18834);
nor U20912 (N_20912,N_18607,N_17785);
nor U20913 (N_20913,N_19036,N_18273);
or U20914 (N_20914,N_19353,N_19273);
nor U20915 (N_20915,N_18032,N_19475);
xor U20916 (N_20916,N_18425,N_17692);
and U20917 (N_20917,N_19206,N_19556);
nor U20918 (N_20918,N_17514,N_18470);
and U20919 (N_20919,N_19804,N_17844);
nand U20920 (N_20920,N_17815,N_17964);
xnor U20921 (N_20921,N_19538,N_19481);
or U20922 (N_20922,N_18489,N_18357);
or U20923 (N_20923,N_19780,N_17762);
or U20924 (N_20924,N_18845,N_17542);
or U20925 (N_20925,N_18424,N_19189);
nand U20926 (N_20926,N_19074,N_17930);
and U20927 (N_20927,N_19573,N_17887);
nand U20928 (N_20928,N_19540,N_19836);
and U20929 (N_20929,N_18821,N_19938);
or U20930 (N_20930,N_18729,N_19953);
nand U20931 (N_20931,N_19715,N_19763);
nor U20932 (N_20932,N_18180,N_17608);
xor U20933 (N_20933,N_19545,N_18560);
and U20934 (N_20934,N_19925,N_19024);
or U20935 (N_20935,N_19108,N_18533);
nand U20936 (N_20936,N_19653,N_19281);
and U20937 (N_20937,N_19835,N_18764);
or U20938 (N_20938,N_19647,N_19801);
and U20939 (N_20939,N_18226,N_17551);
xor U20940 (N_20940,N_19069,N_18546);
xor U20941 (N_20941,N_18054,N_18787);
and U20942 (N_20942,N_19019,N_18642);
xor U20943 (N_20943,N_18162,N_17885);
xor U20944 (N_20944,N_17767,N_18803);
or U20945 (N_20945,N_19796,N_19535);
nor U20946 (N_20946,N_18762,N_18102);
and U20947 (N_20947,N_18062,N_19227);
and U20948 (N_20948,N_19483,N_19151);
and U20949 (N_20949,N_17533,N_19626);
nand U20950 (N_20950,N_18415,N_19537);
and U20951 (N_20951,N_17626,N_19194);
nand U20952 (N_20952,N_18641,N_17982);
and U20953 (N_20953,N_19858,N_18406);
nor U20954 (N_20954,N_19551,N_18895);
xnor U20955 (N_20955,N_17934,N_19428);
nand U20956 (N_20956,N_18419,N_18328);
and U20957 (N_20957,N_17867,N_18125);
and U20958 (N_20958,N_17643,N_19440);
nor U20959 (N_20959,N_18943,N_18036);
nand U20960 (N_20960,N_18843,N_17584);
and U20961 (N_20961,N_18051,N_18024);
nand U20962 (N_20962,N_19837,N_19508);
xor U20963 (N_20963,N_19784,N_18518);
nor U20964 (N_20964,N_19177,N_19565);
or U20965 (N_20965,N_18213,N_17749);
nand U20966 (N_20966,N_18609,N_17577);
nand U20967 (N_20967,N_18077,N_17666);
and U20968 (N_20968,N_19757,N_18274);
nor U20969 (N_20969,N_19619,N_19860);
or U20970 (N_20970,N_17959,N_17837);
nand U20971 (N_20971,N_19996,N_18371);
xor U20972 (N_20972,N_19382,N_18267);
or U20973 (N_20973,N_17684,N_19869);
nand U20974 (N_20974,N_17715,N_18394);
or U20975 (N_20975,N_18969,N_18599);
and U20976 (N_20976,N_18041,N_19053);
nor U20977 (N_20977,N_17890,N_17642);
nand U20978 (N_20978,N_19198,N_18855);
nand U20979 (N_20979,N_17952,N_19646);
xor U20980 (N_20980,N_19469,N_19772);
or U20981 (N_20981,N_18647,N_18918);
nand U20982 (N_20982,N_17960,N_17817);
nand U20983 (N_20983,N_19162,N_17770);
nor U20984 (N_20984,N_19086,N_19182);
xnor U20985 (N_20985,N_18131,N_18009);
nor U20986 (N_20986,N_19697,N_19220);
nand U20987 (N_20987,N_19180,N_18886);
or U20988 (N_20988,N_17615,N_18218);
xor U20989 (N_20989,N_17638,N_19435);
and U20990 (N_20990,N_19187,N_18073);
nor U20991 (N_20991,N_19179,N_18250);
and U20992 (N_20992,N_17504,N_19606);
xor U20993 (N_20993,N_18559,N_18749);
nor U20994 (N_20994,N_18566,N_17621);
xor U20995 (N_20995,N_17819,N_17611);
nor U20996 (N_20996,N_18696,N_19851);
nor U20997 (N_20997,N_18069,N_19898);
or U20998 (N_20998,N_17915,N_19802);
and U20999 (N_20999,N_18615,N_18731);
nor U21000 (N_21000,N_19002,N_18434);
nor U21001 (N_21001,N_18736,N_18498);
nor U21002 (N_21002,N_19335,N_18118);
nand U21003 (N_21003,N_19214,N_19103);
nand U21004 (N_21004,N_19131,N_19575);
and U21005 (N_21005,N_18067,N_19039);
or U21006 (N_21006,N_18252,N_18136);
or U21007 (N_21007,N_19515,N_19341);
xor U21008 (N_21008,N_18973,N_19125);
xor U21009 (N_21009,N_17922,N_18260);
xor U21010 (N_21010,N_17698,N_19073);
nand U21011 (N_21011,N_19964,N_18358);
or U21012 (N_21012,N_17682,N_19863);
and U21013 (N_21013,N_18694,N_18740);
xor U21014 (N_21014,N_18479,N_19960);
and U21015 (N_21015,N_19334,N_18142);
nand U21016 (N_21016,N_19690,N_18456);
nand U21017 (N_21017,N_19090,N_17950);
and U21018 (N_21018,N_19237,N_17516);
nor U21019 (N_21019,N_18887,N_19323);
and U21020 (N_21020,N_19632,N_17512);
or U21021 (N_21021,N_18748,N_19181);
or U21022 (N_21022,N_18865,N_19006);
nor U21023 (N_21023,N_19292,N_18672);
nand U21024 (N_21024,N_19907,N_18799);
nor U21025 (N_21025,N_17823,N_17907);
and U21026 (N_21026,N_18460,N_18660);
or U21027 (N_21027,N_17679,N_19760);
nand U21028 (N_21028,N_18839,N_17714);
nand U21029 (N_21029,N_18323,N_18327);
xnor U21030 (N_21030,N_18557,N_17703);
or U21031 (N_21031,N_18060,N_18558);
nand U21032 (N_21032,N_17936,N_18135);
nand U21033 (N_21033,N_18541,N_19998);
and U21034 (N_21034,N_17591,N_18157);
or U21035 (N_21035,N_17668,N_18241);
or U21036 (N_21036,N_17575,N_18195);
or U21037 (N_21037,N_18272,N_18210);
or U21038 (N_21038,N_19589,N_18643);
xor U21039 (N_21039,N_18484,N_19391);
nand U21040 (N_21040,N_19129,N_17708);
nand U21041 (N_21041,N_17893,N_19522);
nor U21042 (N_21042,N_19548,N_17530);
xnor U21043 (N_21043,N_18429,N_19362);
nor U21044 (N_21044,N_17744,N_18194);
and U21045 (N_21045,N_17846,N_18701);
or U21046 (N_21046,N_19409,N_18038);
xnor U21047 (N_21047,N_18543,N_17983);
nor U21048 (N_21048,N_19829,N_19344);
nor U21049 (N_21049,N_19298,N_18613);
nand U21050 (N_21050,N_18967,N_19815);
nand U21051 (N_21051,N_17665,N_19394);
or U21052 (N_21052,N_19603,N_19954);
or U21053 (N_21053,N_18507,N_18867);
nor U21054 (N_21054,N_19076,N_18203);
xor U21055 (N_21055,N_19871,N_18875);
and U21056 (N_21056,N_18427,N_19511);
or U21057 (N_21057,N_18414,N_18719);
xnor U21058 (N_21058,N_19420,N_19272);
nand U21059 (N_21059,N_19138,N_19931);
and U21060 (N_21060,N_18681,N_18174);
or U21061 (N_21061,N_19910,N_19962);
or U21062 (N_21062,N_18809,N_19684);
nand U21063 (N_21063,N_19102,N_19407);
and U21064 (N_21064,N_17826,N_17697);
xor U21065 (N_21065,N_17991,N_19572);
nand U21066 (N_21066,N_18430,N_19677);
xnor U21067 (N_21067,N_19654,N_19083);
xor U21068 (N_21068,N_19699,N_19781);
nor U21069 (N_21069,N_17732,N_18535);
xor U21070 (N_21070,N_18750,N_18245);
or U21071 (N_21071,N_18148,N_18970);
and U21072 (N_21072,N_17772,N_19027);
or U21073 (N_21073,N_18053,N_17524);
and U21074 (N_21074,N_18468,N_17968);
xor U21075 (N_21075,N_17820,N_19012);
or U21076 (N_21076,N_17604,N_19660);
nor U21077 (N_21077,N_18098,N_19613);
xor U21078 (N_21078,N_19363,N_19137);
and U21079 (N_21079,N_19030,N_19400);
nor U21080 (N_21080,N_19771,N_19357);
and U21081 (N_21081,N_19188,N_19937);
nand U21082 (N_21082,N_17561,N_18172);
xnor U21083 (N_21083,N_19127,N_19008);
or U21084 (N_21084,N_18342,N_17775);
or U21085 (N_21085,N_19987,N_19396);
or U21086 (N_21086,N_19501,N_17619);
or U21087 (N_21087,N_19701,N_19895);
or U21088 (N_21088,N_19999,N_18206);
nand U21089 (N_21089,N_17662,N_18612);
or U21090 (N_21090,N_17737,N_18588);
nand U21091 (N_21091,N_18403,N_19278);
xor U21092 (N_21092,N_19834,N_18043);
nor U21093 (N_21093,N_17919,N_19917);
nand U21094 (N_21094,N_19312,N_18645);
xor U21095 (N_21095,N_18585,N_17769);
xnor U21096 (N_21096,N_17578,N_18080);
and U21097 (N_21097,N_19657,N_18335);
xnor U21098 (N_21098,N_18772,N_17921);
and U21099 (N_21099,N_17505,N_18322);
or U21100 (N_21100,N_19686,N_18227);
or U21101 (N_21101,N_18874,N_18465);
and U21102 (N_21102,N_19094,N_19674);
nand U21103 (N_21103,N_18089,N_19958);
nand U21104 (N_21104,N_18063,N_18586);
xnor U21105 (N_21105,N_18610,N_18373);
and U21106 (N_21106,N_19627,N_18760);
or U21107 (N_21107,N_19880,N_18284);
nor U21108 (N_21108,N_19608,N_17556);
or U21109 (N_21109,N_17953,N_19112);
nor U21110 (N_21110,N_19169,N_17954);
or U21111 (N_21111,N_18859,N_19599);
and U21112 (N_21112,N_18187,N_19011);
nor U21113 (N_21113,N_18819,N_19242);
nor U21114 (N_21114,N_18737,N_18923);
nor U21115 (N_21115,N_18573,N_18677);
nand U21116 (N_21116,N_17709,N_19119);
and U21117 (N_21117,N_19711,N_19947);
nor U21118 (N_21118,N_18885,N_19546);
nand U21119 (N_21119,N_18624,N_18616);
nand U21120 (N_21120,N_18144,N_18888);
nor U21121 (N_21121,N_19905,N_17705);
nand U21122 (N_21122,N_19628,N_18416);
nor U21123 (N_21123,N_18568,N_19166);
xor U21124 (N_21124,N_19749,N_19031);
or U21125 (N_21125,N_19974,N_19499);
nand U21126 (N_21126,N_18966,N_17601);
nor U21127 (N_21127,N_18081,N_19770);
nand U21128 (N_21128,N_19302,N_19806);
nor U21129 (N_21129,N_18814,N_17661);
or U21130 (N_21130,N_19658,N_17875);
and U21131 (N_21131,N_18950,N_18938);
nand U21132 (N_21132,N_18211,N_19034);
nand U21133 (N_21133,N_18156,N_17741);
nand U21134 (N_21134,N_19631,N_19154);
nor U21135 (N_21135,N_19348,N_18391);
and U21136 (N_21136,N_19059,N_18248);
nor U21137 (N_21137,N_18671,N_19693);
nand U21138 (N_21138,N_18676,N_17688);
and U21139 (N_21139,N_19808,N_18101);
nand U21140 (N_21140,N_19509,N_18093);
xor U21141 (N_21141,N_18703,N_18315);
or U21142 (N_21142,N_18868,N_18269);
xor U21143 (N_21143,N_19098,N_19739);
nand U21144 (N_21144,N_18244,N_18068);
and U21145 (N_21145,N_19271,N_17747);
or U21146 (N_21146,N_19208,N_18840);
xnor U21147 (N_21147,N_19460,N_17724);
or U21148 (N_21148,N_18435,N_19803);
nand U21149 (N_21149,N_18934,N_17745);
xor U21150 (N_21150,N_18978,N_19065);
and U21151 (N_21151,N_19959,N_17570);
nor U21152 (N_21152,N_18167,N_19401);
or U21153 (N_21153,N_19497,N_19183);
nor U21154 (N_21154,N_19865,N_19993);
or U21155 (N_21155,N_18076,N_18936);
xnor U21156 (N_21156,N_17711,N_18334);
or U21157 (N_21157,N_17941,N_19649);
and U21158 (N_21158,N_18924,N_19384);
and U21159 (N_21159,N_18584,N_19512);
nor U21160 (N_21160,N_18710,N_19602);
or U21161 (N_21161,N_18196,N_18937);
nor U21162 (N_21162,N_18022,N_18640);
nand U21163 (N_21163,N_18464,N_17912);
and U21164 (N_21164,N_18790,N_18733);
and U21165 (N_21165,N_18977,N_18688);
and U21166 (N_21166,N_19289,N_18716);
nand U21167 (N_21167,N_17677,N_18061);
nor U21168 (N_21168,N_19779,N_18831);
and U21169 (N_21169,N_17552,N_19360);
xor U21170 (N_21170,N_19591,N_19279);
and U21171 (N_21171,N_19339,N_18483);
xnor U21172 (N_21172,N_19068,N_18778);
or U21173 (N_21173,N_17898,N_18451);
xor U21174 (N_21174,N_18668,N_19444);
nand U21175 (N_21175,N_19560,N_19014);
nor U21176 (N_21176,N_19493,N_18418);
nand U21177 (N_21177,N_19333,N_18127);
nand U21178 (N_21178,N_18784,N_18177);
xnor U21179 (N_21179,N_18917,N_19020);
xnor U21180 (N_21180,N_19026,N_19933);
and U21181 (N_21181,N_19867,N_19755);
or U21182 (N_21182,N_18232,N_19105);
nand U21183 (N_21183,N_19320,N_19519);
or U21184 (N_21184,N_19071,N_18463);
or U21185 (N_21185,N_18497,N_19751);
nand U21186 (N_21186,N_17628,N_18215);
nor U21187 (N_21187,N_17729,N_18154);
nand U21188 (N_21188,N_17928,N_17669);
or U21189 (N_21189,N_17966,N_18776);
nor U21190 (N_21190,N_19146,N_17831);
and U21191 (N_21191,N_18428,N_19849);
nand U21192 (N_21192,N_17812,N_19950);
xor U21193 (N_21193,N_18407,N_19489);
nand U21194 (N_21194,N_17842,N_18523);
xnor U21195 (N_21195,N_19934,N_19370);
xor U21196 (N_21196,N_19275,N_19378);
or U21197 (N_21197,N_19192,N_18159);
nand U21198 (N_21198,N_19062,N_18066);
nor U21199 (N_21199,N_19478,N_17717);
xnor U21200 (N_21200,N_18050,N_18049);
or U21201 (N_21201,N_19037,N_19568);
nor U21202 (N_21202,N_19122,N_19132);
and U21203 (N_21203,N_17791,N_17592);
or U21204 (N_21204,N_17706,N_18071);
xor U21205 (N_21205,N_18833,N_18015);
nor U21206 (N_21206,N_18173,N_18630);
nor U21207 (N_21207,N_18426,N_19015);
or U21208 (N_21208,N_19730,N_18006);
nor U21209 (N_21209,N_19375,N_17795);
nor U21210 (N_21210,N_19297,N_18025);
and U21211 (N_21211,N_18693,N_18813);
or U21212 (N_21212,N_17738,N_18625);
or U21213 (N_21213,N_19424,N_19903);
nor U21214 (N_21214,N_19350,N_18906);
and U21215 (N_21215,N_18262,N_19081);
nand U21216 (N_21216,N_19149,N_18441);
xnor U21217 (N_21217,N_19639,N_19264);
or U21218 (N_21218,N_18941,N_19818);
and U21219 (N_21219,N_18205,N_19744);
nand U21220 (N_21220,N_18116,N_19817);
or U21221 (N_21221,N_19283,N_17681);
or U21222 (N_21222,N_18097,N_19688);
xnor U21223 (N_21223,N_17632,N_19738);
xnor U21224 (N_21224,N_17943,N_18873);
and U21225 (N_21225,N_19984,N_19983);
and U21226 (N_21226,N_19047,N_18112);
and U21227 (N_21227,N_18632,N_17771);
nand U21228 (N_21228,N_18928,N_17687);
nand U21229 (N_21229,N_19471,N_19733);
nor U21230 (N_21230,N_19831,N_18883);
and U21231 (N_21231,N_18313,N_19354);
nand U21232 (N_21232,N_17696,N_19773);
nor U21233 (N_21233,N_17981,N_18587);
xor U21234 (N_21234,N_19832,N_18702);
nor U21235 (N_21235,N_18810,N_18755);
nand U21236 (N_21236,N_17871,N_18550);
and U21237 (N_21237,N_19838,N_19949);
and U21238 (N_21238,N_19256,N_19095);
and U21239 (N_21239,N_18500,N_19521);
nand U21240 (N_21240,N_18278,N_19045);
or U21241 (N_21241,N_19328,N_17840);
or U21242 (N_21242,N_19276,N_19043);
nand U21243 (N_21243,N_18836,N_17574);
nor U21244 (N_21244,N_19207,N_19392);
xnor U21245 (N_21245,N_19464,N_19245);
nor U21246 (N_21246,N_18614,N_17528);
nand U21247 (N_21247,N_17544,N_18753);
xor U21248 (N_21248,N_17909,N_19406);
or U21249 (N_21249,N_19769,N_18477);
nand U21250 (N_21250,N_19046,N_17997);
and U21251 (N_21251,N_19924,N_18933);
nor U21252 (N_21252,N_17873,N_18039);
xnor U21253 (N_21253,N_18728,N_19946);
and U21254 (N_21254,N_17833,N_19753);
nor U21255 (N_21255,N_19870,N_18964);
xor U21256 (N_21256,N_17941,N_18304);
xnor U21257 (N_21257,N_17590,N_19764);
and U21258 (N_21258,N_19302,N_18304);
nand U21259 (N_21259,N_19149,N_19805);
xor U21260 (N_21260,N_19505,N_19523);
nand U21261 (N_21261,N_17508,N_18082);
nor U21262 (N_21262,N_19380,N_18195);
nand U21263 (N_21263,N_18920,N_19633);
and U21264 (N_21264,N_19592,N_17623);
nor U21265 (N_21265,N_19144,N_19059);
xnor U21266 (N_21266,N_17751,N_19672);
and U21267 (N_21267,N_19040,N_19334);
xor U21268 (N_21268,N_18113,N_18090);
nand U21269 (N_21269,N_19023,N_18471);
and U21270 (N_21270,N_18124,N_18997);
or U21271 (N_21271,N_18053,N_19960);
or U21272 (N_21272,N_19757,N_18237);
or U21273 (N_21273,N_19812,N_19216);
and U21274 (N_21274,N_17745,N_19382);
xor U21275 (N_21275,N_18987,N_18206);
xnor U21276 (N_21276,N_17580,N_18837);
nand U21277 (N_21277,N_17582,N_18858);
nor U21278 (N_21278,N_18296,N_19505);
xnor U21279 (N_21279,N_18965,N_19376);
or U21280 (N_21280,N_17701,N_18596);
and U21281 (N_21281,N_17985,N_19186);
nand U21282 (N_21282,N_18975,N_19138);
or U21283 (N_21283,N_18434,N_18979);
or U21284 (N_21284,N_18075,N_17577);
nand U21285 (N_21285,N_18001,N_17584);
nand U21286 (N_21286,N_18472,N_19938);
xor U21287 (N_21287,N_18129,N_19125);
and U21288 (N_21288,N_18136,N_19919);
and U21289 (N_21289,N_19293,N_18445);
nand U21290 (N_21290,N_18534,N_19844);
or U21291 (N_21291,N_18712,N_19105);
nor U21292 (N_21292,N_18007,N_19938);
or U21293 (N_21293,N_17617,N_18537);
or U21294 (N_21294,N_17639,N_19326);
nor U21295 (N_21295,N_17574,N_17944);
xnor U21296 (N_21296,N_19994,N_19683);
xnor U21297 (N_21297,N_17534,N_18446);
and U21298 (N_21298,N_17946,N_18423);
xor U21299 (N_21299,N_19252,N_19518);
xnor U21300 (N_21300,N_18032,N_17741);
and U21301 (N_21301,N_19643,N_18893);
nor U21302 (N_21302,N_18398,N_18928);
nand U21303 (N_21303,N_19698,N_18267);
xnor U21304 (N_21304,N_19986,N_18636);
nand U21305 (N_21305,N_19848,N_19048);
or U21306 (N_21306,N_19469,N_18726);
nand U21307 (N_21307,N_19740,N_17801);
xnor U21308 (N_21308,N_19663,N_18981);
or U21309 (N_21309,N_19043,N_19873);
or U21310 (N_21310,N_18270,N_17504);
nand U21311 (N_21311,N_19573,N_18398);
or U21312 (N_21312,N_19944,N_19878);
or U21313 (N_21313,N_18457,N_18483);
xor U21314 (N_21314,N_19534,N_17786);
xor U21315 (N_21315,N_19769,N_18347);
or U21316 (N_21316,N_19489,N_18417);
or U21317 (N_21317,N_19460,N_18009);
or U21318 (N_21318,N_18358,N_18894);
xor U21319 (N_21319,N_17674,N_19720);
nand U21320 (N_21320,N_17781,N_19982);
nand U21321 (N_21321,N_19563,N_18044);
and U21322 (N_21322,N_19080,N_19255);
xnor U21323 (N_21323,N_18710,N_17896);
nor U21324 (N_21324,N_18693,N_19037);
nor U21325 (N_21325,N_17695,N_17517);
nand U21326 (N_21326,N_19204,N_19403);
and U21327 (N_21327,N_19497,N_19652);
nand U21328 (N_21328,N_17692,N_19576);
nand U21329 (N_21329,N_19202,N_18820);
xor U21330 (N_21330,N_17839,N_19796);
or U21331 (N_21331,N_18193,N_17512);
and U21332 (N_21332,N_17880,N_17863);
nor U21333 (N_21333,N_19296,N_18168);
xnor U21334 (N_21334,N_19336,N_19865);
xor U21335 (N_21335,N_19377,N_18165);
nor U21336 (N_21336,N_17693,N_19177);
nor U21337 (N_21337,N_19334,N_19632);
or U21338 (N_21338,N_18701,N_19102);
nor U21339 (N_21339,N_19049,N_18278);
and U21340 (N_21340,N_18895,N_18848);
nor U21341 (N_21341,N_18911,N_19359);
xnor U21342 (N_21342,N_19419,N_17760);
or U21343 (N_21343,N_18775,N_19038);
nor U21344 (N_21344,N_18437,N_19447);
and U21345 (N_21345,N_18252,N_19131);
nor U21346 (N_21346,N_18830,N_18350);
and U21347 (N_21347,N_18373,N_19348);
nand U21348 (N_21348,N_19988,N_19780);
and U21349 (N_21349,N_17574,N_17739);
nand U21350 (N_21350,N_18621,N_18795);
and U21351 (N_21351,N_18682,N_18546);
nand U21352 (N_21352,N_19905,N_19825);
xor U21353 (N_21353,N_19087,N_19023);
nor U21354 (N_21354,N_18388,N_18661);
xnor U21355 (N_21355,N_19436,N_19380);
nand U21356 (N_21356,N_18389,N_17680);
and U21357 (N_21357,N_18058,N_18799);
nor U21358 (N_21358,N_19655,N_19820);
nand U21359 (N_21359,N_17753,N_19831);
nand U21360 (N_21360,N_17670,N_17682);
xnor U21361 (N_21361,N_19303,N_19659);
and U21362 (N_21362,N_18103,N_18479);
xor U21363 (N_21363,N_19591,N_17782);
nand U21364 (N_21364,N_19716,N_19824);
or U21365 (N_21365,N_17993,N_18015);
or U21366 (N_21366,N_18777,N_19354);
and U21367 (N_21367,N_17765,N_18402);
or U21368 (N_21368,N_17841,N_18140);
nor U21369 (N_21369,N_18367,N_17685);
or U21370 (N_21370,N_18216,N_18012);
nand U21371 (N_21371,N_17986,N_19565);
xnor U21372 (N_21372,N_18984,N_17742);
or U21373 (N_21373,N_18824,N_18257);
nor U21374 (N_21374,N_18539,N_17628);
or U21375 (N_21375,N_19770,N_17693);
xor U21376 (N_21376,N_19747,N_18516);
and U21377 (N_21377,N_18197,N_18363);
nor U21378 (N_21378,N_18832,N_18302);
xor U21379 (N_21379,N_19822,N_18226);
and U21380 (N_21380,N_17694,N_19893);
or U21381 (N_21381,N_18153,N_17898);
nand U21382 (N_21382,N_18099,N_19203);
nor U21383 (N_21383,N_18577,N_18800);
and U21384 (N_21384,N_18931,N_19406);
nand U21385 (N_21385,N_18071,N_19538);
xnor U21386 (N_21386,N_18470,N_19707);
nor U21387 (N_21387,N_18872,N_19947);
xnor U21388 (N_21388,N_19970,N_19441);
nor U21389 (N_21389,N_17527,N_17649);
nand U21390 (N_21390,N_19665,N_18654);
nand U21391 (N_21391,N_18227,N_19518);
nor U21392 (N_21392,N_19757,N_17817);
nand U21393 (N_21393,N_18364,N_19474);
xor U21394 (N_21394,N_19097,N_19348);
nand U21395 (N_21395,N_19294,N_18956);
nor U21396 (N_21396,N_18003,N_17812);
or U21397 (N_21397,N_17851,N_19056);
nand U21398 (N_21398,N_19280,N_19728);
nor U21399 (N_21399,N_19096,N_18358);
or U21400 (N_21400,N_17852,N_19795);
nand U21401 (N_21401,N_18582,N_18133);
nand U21402 (N_21402,N_18869,N_18438);
and U21403 (N_21403,N_18670,N_18945);
or U21404 (N_21404,N_19094,N_18392);
xnor U21405 (N_21405,N_18932,N_18894);
xnor U21406 (N_21406,N_19787,N_17660);
and U21407 (N_21407,N_17530,N_19742);
nor U21408 (N_21408,N_18768,N_18570);
xor U21409 (N_21409,N_18688,N_18411);
or U21410 (N_21410,N_19356,N_18708);
and U21411 (N_21411,N_18199,N_17873);
and U21412 (N_21412,N_19517,N_17690);
nand U21413 (N_21413,N_19589,N_18390);
and U21414 (N_21414,N_18236,N_17698);
nand U21415 (N_21415,N_19148,N_19874);
nor U21416 (N_21416,N_18369,N_18483);
xnor U21417 (N_21417,N_18211,N_19141);
nand U21418 (N_21418,N_17937,N_19295);
or U21419 (N_21419,N_18973,N_19386);
or U21420 (N_21420,N_18512,N_17987);
nand U21421 (N_21421,N_18548,N_19476);
nor U21422 (N_21422,N_18155,N_17764);
and U21423 (N_21423,N_17936,N_19946);
and U21424 (N_21424,N_18434,N_17615);
nand U21425 (N_21425,N_17704,N_19058);
nor U21426 (N_21426,N_18845,N_18327);
or U21427 (N_21427,N_17778,N_19139);
nand U21428 (N_21428,N_19916,N_19943);
nor U21429 (N_21429,N_17959,N_17531);
or U21430 (N_21430,N_19277,N_19454);
and U21431 (N_21431,N_17755,N_19790);
xor U21432 (N_21432,N_18931,N_17887);
nor U21433 (N_21433,N_18664,N_18251);
xnor U21434 (N_21434,N_18708,N_19583);
nor U21435 (N_21435,N_19894,N_18264);
and U21436 (N_21436,N_19063,N_18214);
and U21437 (N_21437,N_18865,N_18314);
xnor U21438 (N_21438,N_18534,N_17786);
nand U21439 (N_21439,N_19762,N_19327);
and U21440 (N_21440,N_18963,N_19949);
and U21441 (N_21441,N_19416,N_19690);
xor U21442 (N_21442,N_18326,N_19107);
and U21443 (N_21443,N_18725,N_18283);
xor U21444 (N_21444,N_19391,N_19169);
xor U21445 (N_21445,N_19450,N_18118);
xor U21446 (N_21446,N_17611,N_18926);
and U21447 (N_21447,N_17507,N_18279);
and U21448 (N_21448,N_18619,N_18478);
and U21449 (N_21449,N_17517,N_17817);
xnor U21450 (N_21450,N_18422,N_18300);
nand U21451 (N_21451,N_19948,N_19936);
or U21452 (N_21452,N_18673,N_17577);
and U21453 (N_21453,N_19386,N_17847);
nor U21454 (N_21454,N_19848,N_18603);
or U21455 (N_21455,N_18003,N_18811);
or U21456 (N_21456,N_17515,N_18576);
or U21457 (N_21457,N_19247,N_19953);
or U21458 (N_21458,N_17629,N_18554);
nor U21459 (N_21459,N_18807,N_18247);
nand U21460 (N_21460,N_18047,N_19841);
nor U21461 (N_21461,N_18531,N_19940);
xnor U21462 (N_21462,N_18791,N_19644);
and U21463 (N_21463,N_19692,N_18201);
nor U21464 (N_21464,N_18902,N_18232);
xor U21465 (N_21465,N_18004,N_19566);
nand U21466 (N_21466,N_18408,N_17924);
xnor U21467 (N_21467,N_18171,N_17814);
xnor U21468 (N_21468,N_19480,N_18120);
and U21469 (N_21469,N_18254,N_18149);
nor U21470 (N_21470,N_19688,N_17630);
nor U21471 (N_21471,N_18894,N_19693);
nor U21472 (N_21472,N_19493,N_19393);
nand U21473 (N_21473,N_18415,N_17789);
nor U21474 (N_21474,N_18542,N_18061);
and U21475 (N_21475,N_18638,N_18910);
or U21476 (N_21476,N_17888,N_18876);
xor U21477 (N_21477,N_17626,N_19533);
nand U21478 (N_21478,N_18182,N_17591);
and U21479 (N_21479,N_18310,N_17636);
xnor U21480 (N_21480,N_18008,N_18870);
or U21481 (N_21481,N_19341,N_17752);
nand U21482 (N_21482,N_18975,N_18164);
and U21483 (N_21483,N_19850,N_18026);
nand U21484 (N_21484,N_19389,N_18113);
nand U21485 (N_21485,N_18949,N_19085);
and U21486 (N_21486,N_19684,N_19600);
nand U21487 (N_21487,N_18666,N_18909);
nor U21488 (N_21488,N_18756,N_19672);
xor U21489 (N_21489,N_19290,N_17579);
xor U21490 (N_21490,N_19953,N_18877);
nand U21491 (N_21491,N_17992,N_18202);
or U21492 (N_21492,N_19311,N_18997);
xnor U21493 (N_21493,N_18864,N_17551);
or U21494 (N_21494,N_19242,N_17998);
and U21495 (N_21495,N_18758,N_18831);
nor U21496 (N_21496,N_18487,N_19605);
and U21497 (N_21497,N_19277,N_18327);
nand U21498 (N_21498,N_17743,N_19508);
nand U21499 (N_21499,N_17704,N_17811);
xnor U21500 (N_21500,N_18053,N_19097);
and U21501 (N_21501,N_19415,N_17715);
nand U21502 (N_21502,N_19385,N_19077);
nand U21503 (N_21503,N_17828,N_17952);
xor U21504 (N_21504,N_17630,N_18039);
or U21505 (N_21505,N_18585,N_19043);
nand U21506 (N_21506,N_19354,N_19154);
nor U21507 (N_21507,N_18689,N_18697);
or U21508 (N_21508,N_18557,N_19821);
xnor U21509 (N_21509,N_19397,N_17962);
nand U21510 (N_21510,N_19474,N_18585);
and U21511 (N_21511,N_19849,N_19631);
or U21512 (N_21512,N_17920,N_19282);
nor U21513 (N_21513,N_18799,N_18028);
nor U21514 (N_21514,N_19905,N_19989);
nand U21515 (N_21515,N_18743,N_18863);
nor U21516 (N_21516,N_18015,N_17977);
or U21517 (N_21517,N_19995,N_17576);
xor U21518 (N_21518,N_19940,N_17604);
nor U21519 (N_21519,N_18423,N_18782);
and U21520 (N_21520,N_18729,N_17518);
or U21521 (N_21521,N_18665,N_19778);
xnor U21522 (N_21522,N_19038,N_18313);
xor U21523 (N_21523,N_19693,N_19299);
or U21524 (N_21524,N_17524,N_19917);
and U21525 (N_21525,N_17812,N_18494);
xnor U21526 (N_21526,N_18794,N_17716);
and U21527 (N_21527,N_19163,N_19254);
xnor U21528 (N_21528,N_18996,N_19567);
nand U21529 (N_21529,N_17692,N_18678);
or U21530 (N_21530,N_18511,N_17693);
nand U21531 (N_21531,N_17733,N_19990);
xnor U21532 (N_21532,N_19546,N_17819);
nand U21533 (N_21533,N_19894,N_19833);
nand U21534 (N_21534,N_18979,N_19284);
or U21535 (N_21535,N_18798,N_17667);
or U21536 (N_21536,N_18381,N_18098);
and U21537 (N_21537,N_19156,N_17609);
nor U21538 (N_21538,N_19015,N_17842);
and U21539 (N_21539,N_17764,N_17941);
xnor U21540 (N_21540,N_18643,N_17564);
xor U21541 (N_21541,N_19897,N_17646);
nor U21542 (N_21542,N_18250,N_18945);
nand U21543 (N_21543,N_19830,N_17693);
nand U21544 (N_21544,N_19096,N_17922);
nand U21545 (N_21545,N_19857,N_18934);
xor U21546 (N_21546,N_19653,N_19566);
xor U21547 (N_21547,N_19848,N_19156);
and U21548 (N_21548,N_19532,N_17567);
or U21549 (N_21549,N_18863,N_19738);
nand U21550 (N_21550,N_19617,N_18872);
and U21551 (N_21551,N_19772,N_18479);
or U21552 (N_21552,N_19779,N_18170);
xor U21553 (N_21553,N_17786,N_18178);
and U21554 (N_21554,N_19126,N_19565);
and U21555 (N_21555,N_18985,N_18360);
nand U21556 (N_21556,N_18736,N_18348);
or U21557 (N_21557,N_17984,N_18569);
nand U21558 (N_21558,N_18512,N_18535);
and U21559 (N_21559,N_18962,N_19601);
xnor U21560 (N_21560,N_18664,N_19879);
nand U21561 (N_21561,N_19741,N_18495);
nand U21562 (N_21562,N_18642,N_18385);
xnor U21563 (N_21563,N_19152,N_18310);
xor U21564 (N_21564,N_17898,N_19977);
and U21565 (N_21565,N_19431,N_19086);
and U21566 (N_21566,N_19965,N_18385);
xor U21567 (N_21567,N_19861,N_17988);
nand U21568 (N_21568,N_19151,N_19006);
and U21569 (N_21569,N_19983,N_17773);
nand U21570 (N_21570,N_18043,N_19868);
or U21571 (N_21571,N_19224,N_17861);
and U21572 (N_21572,N_19137,N_19229);
nor U21573 (N_21573,N_19197,N_19730);
xnor U21574 (N_21574,N_18548,N_19759);
xor U21575 (N_21575,N_18588,N_18565);
or U21576 (N_21576,N_18744,N_17933);
and U21577 (N_21577,N_18038,N_17693);
xor U21578 (N_21578,N_19338,N_19072);
xnor U21579 (N_21579,N_17729,N_18638);
nand U21580 (N_21580,N_19895,N_19256);
nor U21581 (N_21581,N_17532,N_18493);
nor U21582 (N_21582,N_18441,N_17577);
or U21583 (N_21583,N_18061,N_17854);
and U21584 (N_21584,N_17986,N_19082);
and U21585 (N_21585,N_18214,N_17656);
and U21586 (N_21586,N_18934,N_19682);
xor U21587 (N_21587,N_18829,N_19708);
xnor U21588 (N_21588,N_19907,N_18163);
xor U21589 (N_21589,N_19734,N_18431);
and U21590 (N_21590,N_19849,N_18429);
and U21591 (N_21591,N_18307,N_19404);
or U21592 (N_21592,N_17653,N_19636);
and U21593 (N_21593,N_18778,N_18091);
nand U21594 (N_21594,N_19402,N_17526);
nand U21595 (N_21595,N_18875,N_19349);
or U21596 (N_21596,N_19284,N_19001);
or U21597 (N_21597,N_19555,N_19719);
nand U21598 (N_21598,N_19730,N_19577);
xor U21599 (N_21599,N_18692,N_19398);
nor U21600 (N_21600,N_18771,N_18213);
or U21601 (N_21601,N_18959,N_19096);
and U21602 (N_21602,N_18710,N_19853);
xor U21603 (N_21603,N_18191,N_18399);
or U21604 (N_21604,N_19136,N_18782);
nand U21605 (N_21605,N_18595,N_19332);
xor U21606 (N_21606,N_18808,N_18769);
and U21607 (N_21607,N_18711,N_18081);
xnor U21608 (N_21608,N_18563,N_17932);
or U21609 (N_21609,N_17811,N_17816);
nor U21610 (N_21610,N_19971,N_18109);
or U21611 (N_21611,N_19792,N_19552);
xor U21612 (N_21612,N_18717,N_19389);
nor U21613 (N_21613,N_18022,N_19998);
nand U21614 (N_21614,N_17948,N_19798);
nor U21615 (N_21615,N_19285,N_18371);
and U21616 (N_21616,N_17642,N_19978);
and U21617 (N_21617,N_19139,N_18788);
xor U21618 (N_21618,N_18783,N_17560);
nand U21619 (N_21619,N_18445,N_18627);
nor U21620 (N_21620,N_18262,N_19110);
xnor U21621 (N_21621,N_19575,N_19696);
and U21622 (N_21622,N_18900,N_18993);
nor U21623 (N_21623,N_18992,N_19286);
xor U21624 (N_21624,N_19751,N_19790);
nand U21625 (N_21625,N_19721,N_18193);
xor U21626 (N_21626,N_19623,N_18612);
and U21627 (N_21627,N_18400,N_17598);
xnor U21628 (N_21628,N_19859,N_18574);
nand U21629 (N_21629,N_19092,N_17988);
and U21630 (N_21630,N_19614,N_17558);
or U21631 (N_21631,N_18423,N_17596);
xor U21632 (N_21632,N_18599,N_17801);
or U21633 (N_21633,N_18723,N_17784);
xor U21634 (N_21634,N_18995,N_17967);
nand U21635 (N_21635,N_19123,N_19151);
and U21636 (N_21636,N_18849,N_19324);
or U21637 (N_21637,N_18233,N_18479);
xor U21638 (N_21638,N_19492,N_19699);
and U21639 (N_21639,N_18871,N_17936);
nand U21640 (N_21640,N_19840,N_17935);
or U21641 (N_21641,N_18366,N_19464);
nor U21642 (N_21642,N_18644,N_18316);
nor U21643 (N_21643,N_19598,N_19906);
nand U21644 (N_21644,N_17606,N_18165);
nor U21645 (N_21645,N_19216,N_17513);
nand U21646 (N_21646,N_18682,N_19108);
nor U21647 (N_21647,N_19553,N_18796);
or U21648 (N_21648,N_18475,N_19820);
nand U21649 (N_21649,N_17688,N_18952);
nand U21650 (N_21650,N_19251,N_17924);
and U21651 (N_21651,N_18178,N_17531);
xnor U21652 (N_21652,N_17865,N_18567);
or U21653 (N_21653,N_18272,N_19825);
and U21654 (N_21654,N_19599,N_18532);
xor U21655 (N_21655,N_17666,N_19280);
and U21656 (N_21656,N_17982,N_18268);
nand U21657 (N_21657,N_18507,N_17516);
or U21658 (N_21658,N_19010,N_18537);
and U21659 (N_21659,N_18620,N_19459);
or U21660 (N_21660,N_18389,N_19695);
or U21661 (N_21661,N_19419,N_19341);
nand U21662 (N_21662,N_18263,N_17941);
nand U21663 (N_21663,N_18294,N_19905);
nand U21664 (N_21664,N_18067,N_17686);
nand U21665 (N_21665,N_17929,N_18557);
xor U21666 (N_21666,N_18803,N_18415);
nand U21667 (N_21667,N_19105,N_19555);
or U21668 (N_21668,N_18153,N_18234);
xnor U21669 (N_21669,N_19402,N_19774);
xor U21670 (N_21670,N_17954,N_18034);
or U21671 (N_21671,N_19521,N_19178);
nor U21672 (N_21672,N_17843,N_17995);
and U21673 (N_21673,N_19019,N_18697);
nand U21674 (N_21674,N_19867,N_19689);
and U21675 (N_21675,N_18198,N_19583);
and U21676 (N_21676,N_19936,N_17675);
or U21677 (N_21677,N_17887,N_19299);
or U21678 (N_21678,N_18676,N_18806);
and U21679 (N_21679,N_17928,N_18254);
or U21680 (N_21680,N_17777,N_19878);
nand U21681 (N_21681,N_17963,N_19933);
nand U21682 (N_21682,N_18291,N_18563);
and U21683 (N_21683,N_18231,N_18386);
xor U21684 (N_21684,N_18289,N_19938);
and U21685 (N_21685,N_19850,N_19547);
and U21686 (N_21686,N_19026,N_18867);
xnor U21687 (N_21687,N_19089,N_19380);
xnor U21688 (N_21688,N_18711,N_18381);
nor U21689 (N_21689,N_17690,N_18388);
and U21690 (N_21690,N_17598,N_17856);
and U21691 (N_21691,N_19560,N_18077);
nor U21692 (N_21692,N_18988,N_17917);
and U21693 (N_21693,N_17523,N_19761);
and U21694 (N_21694,N_19736,N_19689);
xor U21695 (N_21695,N_18425,N_19729);
xor U21696 (N_21696,N_17746,N_18657);
nor U21697 (N_21697,N_17833,N_17792);
and U21698 (N_21698,N_17610,N_19679);
nand U21699 (N_21699,N_18987,N_19961);
nand U21700 (N_21700,N_18002,N_17671);
or U21701 (N_21701,N_18004,N_18690);
nand U21702 (N_21702,N_17591,N_17638);
and U21703 (N_21703,N_18977,N_19556);
nor U21704 (N_21704,N_19422,N_18754);
and U21705 (N_21705,N_18177,N_19429);
or U21706 (N_21706,N_18186,N_18460);
or U21707 (N_21707,N_18056,N_19174);
or U21708 (N_21708,N_17544,N_17776);
or U21709 (N_21709,N_19144,N_18225);
nor U21710 (N_21710,N_17664,N_19529);
nor U21711 (N_21711,N_18805,N_19700);
xnor U21712 (N_21712,N_19705,N_19811);
or U21713 (N_21713,N_19929,N_17677);
nor U21714 (N_21714,N_17812,N_17849);
or U21715 (N_21715,N_18247,N_18309);
nor U21716 (N_21716,N_19158,N_19090);
and U21717 (N_21717,N_19561,N_18457);
or U21718 (N_21718,N_19466,N_18985);
nand U21719 (N_21719,N_19181,N_17558);
xnor U21720 (N_21720,N_18672,N_18461);
and U21721 (N_21721,N_19834,N_17865);
nand U21722 (N_21722,N_19091,N_18229);
and U21723 (N_21723,N_18196,N_19920);
nand U21724 (N_21724,N_19251,N_19717);
or U21725 (N_21725,N_18058,N_18994);
nor U21726 (N_21726,N_18036,N_19551);
and U21727 (N_21727,N_19429,N_17599);
and U21728 (N_21728,N_18621,N_19422);
nor U21729 (N_21729,N_18259,N_18300);
nand U21730 (N_21730,N_17587,N_19894);
nor U21731 (N_21731,N_18198,N_18982);
or U21732 (N_21732,N_18559,N_18687);
and U21733 (N_21733,N_17960,N_19307);
xnor U21734 (N_21734,N_17767,N_19892);
nand U21735 (N_21735,N_19171,N_19743);
nor U21736 (N_21736,N_19745,N_17922);
nor U21737 (N_21737,N_18570,N_17537);
nor U21738 (N_21738,N_18228,N_19133);
nand U21739 (N_21739,N_19905,N_17769);
and U21740 (N_21740,N_19599,N_18218);
nand U21741 (N_21741,N_19046,N_18654);
or U21742 (N_21742,N_19963,N_19006);
xnor U21743 (N_21743,N_18254,N_19091);
or U21744 (N_21744,N_19471,N_17968);
nand U21745 (N_21745,N_19737,N_19813);
nor U21746 (N_21746,N_18029,N_19376);
nand U21747 (N_21747,N_19526,N_18354);
nand U21748 (N_21748,N_19362,N_17663);
nand U21749 (N_21749,N_19984,N_18043);
and U21750 (N_21750,N_19375,N_19292);
nor U21751 (N_21751,N_17510,N_19179);
and U21752 (N_21752,N_19803,N_18022);
nand U21753 (N_21753,N_18516,N_17934);
nand U21754 (N_21754,N_17807,N_17541);
and U21755 (N_21755,N_19694,N_17890);
xor U21756 (N_21756,N_19730,N_19170);
nand U21757 (N_21757,N_18338,N_17552);
nand U21758 (N_21758,N_19482,N_18959);
and U21759 (N_21759,N_18261,N_18938);
xnor U21760 (N_21760,N_19032,N_17741);
and U21761 (N_21761,N_17637,N_18326);
xor U21762 (N_21762,N_18192,N_18429);
xor U21763 (N_21763,N_18088,N_18159);
xnor U21764 (N_21764,N_17816,N_19698);
nor U21765 (N_21765,N_17742,N_18228);
xor U21766 (N_21766,N_18724,N_18062);
xnor U21767 (N_21767,N_19318,N_19973);
nand U21768 (N_21768,N_19410,N_19843);
or U21769 (N_21769,N_17567,N_19650);
or U21770 (N_21770,N_19582,N_17530);
nand U21771 (N_21771,N_17886,N_19839);
or U21772 (N_21772,N_18161,N_17827);
xor U21773 (N_21773,N_18262,N_18079);
and U21774 (N_21774,N_19314,N_17989);
xor U21775 (N_21775,N_18381,N_17557);
nor U21776 (N_21776,N_18831,N_18772);
nor U21777 (N_21777,N_19330,N_19203);
nor U21778 (N_21778,N_19869,N_19213);
xor U21779 (N_21779,N_19735,N_19244);
nand U21780 (N_21780,N_19726,N_19885);
and U21781 (N_21781,N_18581,N_18313);
xnor U21782 (N_21782,N_17620,N_18567);
nor U21783 (N_21783,N_17667,N_19584);
xor U21784 (N_21784,N_19853,N_18091);
or U21785 (N_21785,N_19132,N_18086);
nor U21786 (N_21786,N_19390,N_18012);
nand U21787 (N_21787,N_18996,N_19854);
and U21788 (N_21788,N_18241,N_19919);
nor U21789 (N_21789,N_17951,N_18256);
or U21790 (N_21790,N_19393,N_19634);
nor U21791 (N_21791,N_18003,N_18636);
nand U21792 (N_21792,N_19410,N_17766);
nor U21793 (N_21793,N_19928,N_19363);
and U21794 (N_21794,N_18136,N_19792);
nor U21795 (N_21795,N_17948,N_19720);
xnor U21796 (N_21796,N_19609,N_18929);
and U21797 (N_21797,N_19621,N_17714);
nor U21798 (N_21798,N_18885,N_18832);
and U21799 (N_21799,N_17623,N_19703);
xnor U21800 (N_21800,N_17904,N_18891);
or U21801 (N_21801,N_18890,N_18210);
and U21802 (N_21802,N_18436,N_19404);
nor U21803 (N_21803,N_19220,N_18331);
nand U21804 (N_21804,N_18723,N_18295);
xor U21805 (N_21805,N_18961,N_18847);
nand U21806 (N_21806,N_17778,N_19672);
and U21807 (N_21807,N_18432,N_18247);
and U21808 (N_21808,N_19206,N_18659);
nor U21809 (N_21809,N_19692,N_19806);
nor U21810 (N_21810,N_18686,N_19191);
and U21811 (N_21811,N_18136,N_19133);
or U21812 (N_21812,N_17631,N_17594);
nor U21813 (N_21813,N_18003,N_17831);
and U21814 (N_21814,N_18904,N_18811);
nor U21815 (N_21815,N_17630,N_18379);
or U21816 (N_21816,N_19376,N_19464);
nand U21817 (N_21817,N_19308,N_18782);
nand U21818 (N_21818,N_19072,N_19612);
nor U21819 (N_21819,N_19017,N_19303);
or U21820 (N_21820,N_18249,N_18294);
nor U21821 (N_21821,N_19474,N_19029);
xnor U21822 (N_21822,N_18059,N_19745);
nand U21823 (N_21823,N_18039,N_18998);
or U21824 (N_21824,N_19609,N_18202);
and U21825 (N_21825,N_18362,N_18228);
nand U21826 (N_21826,N_19035,N_18038);
nor U21827 (N_21827,N_19745,N_18565);
or U21828 (N_21828,N_19591,N_17512);
nand U21829 (N_21829,N_19586,N_18777);
xor U21830 (N_21830,N_18465,N_19857);
xnor U21831 (N_21831,N_18898,N_19628);
or U21832 (N_21832,N_18122,N_19893);
and U21833 (N_21833,N_19974,N_18434);
and U21834 (N_21834,N_19891,N_19785);
or U21835 (N_21835,N_19265,N_19119);
nand U21836 (N_21836,N_18647,N_18308);
nor U21837 (N_21837,N_19299,N_19823);
or U21838 (N_21838,N_18216,N_18651);
or U21839 (N_21839,N_19631,N_18731);
and U21840 (N_21840,N_18242,N_17636);
xnor U21841 (N_21841,N_18653,N_17514);
xor U21842 (N_21842,N_18230,N_18363);
nand U21843 (N_21843,N_19612,N_19762);
nand U21844 (N_21844,N_18960,N_18111);
xnor U21845 (N_21845,N_18402,N_17752);
and U21846 (N_21846,N_17697,N_19946);
nor U21847 (N_21847,N_17792,N_18901);
nand U21848 (N_21848,N_19811,N_18923);
xor U21849 (N_21849,N_18512,N_19550);
xor U21850 (N_21850,N_19370,N_18023);
nor U21851 (N_21851,N_19411,N_18332);
nor U21852 (N_21852,N_18075,N_19295);
nand U21853 (N_21853,N_18151,N_19188);
or U21854 (N_21854,N_18201,N_18476);
and U21855 (N_21855,N_18547,N_18246);
xor U21856 (N_21856,N_19331,N_19007);
xor U21857 (N_21857,N_19759,N_18405);
nand U21858 (N_21858,N_19164,N_18592);
and U21859 (N_21859,N_18274,N_18985);
nor U21860 (N_21860,N_19293,N_19590);
or U21861 (N_21861,N_19866,N_19186);
and U21862 (N_21862,N_18971,N_18509);
nand U21863 (N_21863,N_18739,N_18201);
or U21864 (N_21864,N_18435,N_17830);
nor U21865 (N_21865,N_18043,N_18682);
xor U21866 (N_21866,N_18163,N_18779);
and U21867 (N_21867,N_18602,N_18134);
or U21868 (N_21868,N_18150,N_19525);
nand U21869 (N_21869,N_17854,N_18313);
xor U21870 (N_21870,N_19948,N_17528);
nor U21871 (N_21871,N_17932,N_18600);
nor U21872 (N_21872,N_18993,N_17929);
nor U21873 (N_21873,N_19798,N_19397);
nor U21874 (N_21874,N_19567,N_19748);
nand U21875 (N_21875,N_19516,N_18443);
nand U21876 (N_21876,N_18618,N_18273);
nor U21877 (N_21877,N_18968,N_18115);
or U21878 (N_21878,N_18893,N_17546);
xor U21879 (N_21879,N_18870,N_18086);
nor U21880 (N_21880,N_18468,N_19576);
and U21881 (N_21881,N_18983,N_18208);
nor U21882 (N_21882,N_18128,N_19443);
nand U21883 (N_21883,N_17966,N_19765);
and U21884 (N_21884,N_19914,N_18036);
or U21885 (N_21885,N_19494,N_17560);
nor U21886 (N_21886,N_17617,N_18221);
nand U21887 (N_21887,N_19530,N_19858);
nor U21888 (N_21888,N_18417,N_18334);
or U21889 (N_21889,N_19800,N_19271);
nor U21890 (N_21890,N_18667,N_18861);
or U21891 (N_21891,N_18640,N_19164);
nand U21892 (N_21892,N_18535,N_18145);
nand U21893 (N_21893,N_18194,N_17885);
or U21894 (N_21894,N_19857,N_17521);
nor U21895 (N_21895,N_18100,N_18925);
and U21896 (N_21896,N_17806,N_18282);
nor U21897 (N_21897,N_18814,N_18609);
nor U21898 (N_21898,N_19037,N_17659);
and U21899 (N_21899,N_18010,N_18264);
or U21900 (N_21900,N_19957,N_19012);
nand U21901 (N_21901,N_19928,N_18260);
or U21902 (N_21902,N_19346,N_19345);
xor U21903 (N_21903,N_18866,N_18952);
nor U21904 (N_21904,N_18390,N_19685);
xnor U21905 (N_21905,N_18111,N_18556);
nand U21906 (N_21906,N_18076,N_17691);
and U21907 (N_21907,N_17845,N_18811);
or U21908 (N_21908,N_19516,N_19340);
nor U21909 (N_21909,N_18213,N_18589);
nand U21910 (N_21910,N_17637,N_19004);
and U21911 (N_21911,N_18569,N_19527);
xnor U21912 (N_21912,N_18038,N_18370);
xor U21913 (N_21913,N_18466,N_18145);
or U21914 (N_21914,N_18636,N_19469);
and U21915 (N_21915,N_18742,N_18141);
or U21916 (N_21916,N_18038,N_18663);
or U21917 (N_21917,N_18252,N_18697);
xor U21918 (N_21918,N_19264,N_18226);
nor U21919 (N_21919,N_18883,N_19841);
and U21920 (N_21920,N_18614,N_19975);
nand U21921 (N_21921,N_19745,N_18238);
or U21922 (N_21922,N_19763,N_17526);
and U21923 (N_21923,N_19893,N_18300);
nor U21924 (N_21924,N_19312,N_19249);
or U21925 (N_21925,N_18738,N_18167);
and U21926 (N_21926,N_17989,N_19139);
xor U21927 (N_21927,N_17520,N_17690);
xnor U21928 (N_21928,N_17860,N_17746);
xnor U21929 (N_21929,N_18912,N_19944);
or U21930 (N_21930,N_18223,N_19346);
nand U21931 (N_21931,N_17500,N_18696);
xor U21932 (N_21932,N_18786,N_19472);
and U21933 (N_21933,N_17604,N_19555);
xnor U21934 (N_21934,N_18617,N_19029);
nor U21935 (N_21935,N_18241,N_17780);
nand U21936 (N_21936,N_18066,N_19432);
nor U21937 (N_21937,N_19988,N_18029);
nand U21938 (N_21938,N_19232,N_18202);
nor U21939 (N_21939,N_18344,N_19378);
and U21940 (N_21940,N_18901,N_19720);
nand U21941 (N_21941,N_19547,N_19001);
nor U21942 (N_21942,N_19794,N_18865);
or U21943 (N_21943,N_19793,N_18056);
or U21944 (N_21944,N_17733,N_18202);
and U21945 (N_21945,N_18084,N_18252);
or U21946 (N_21946,N_19858,N_19364);
nand U21947 (N_21947,N_19039,N_19050);
or U21948 (N_21948,N_17541,N_18644);
and U21949 (N_21949,N_19841,N_18209);
or U21950 (N_21950,N_17530,N_19991);
xnor U21951 (N_21951,N_18565,N_19408);
nor U21952 (N_21952,N_17977,N_18424);
nor U21953 (N_21953,N_19175,N_18952);
nor U21954 (N_21954,N_18559,N_18228);
nor U21955 (N_21955,N_17811,N_19305);
nor U21956 (N_21956,N_18638,N_18023);
nand U21957 (N_21957,N_19478,N_19371);
xnor U21958 (N_21958,N_17896,N_18028);
xnor U21959 (N_21959,N_17534,N_19124);
nor U21960 (N_21960,N_19656,N_18009);
xnor U21961 (N_21961,N_19409,N_17967);
xor U21962 (N_21962,N_17853,N_18085);
and U21963 (N_21963,N_17599,N_17771);
xor U21964 (N_21964,N_19163,N_18242);
nor U21965 (N_21965,N_19062,N_18965);
or U21966 (N_21966,N_19765,N_17674);
nand U21967 (N_21967,N_19516,N_17969);
xor U21968 (N_21968,N_19161,N_19526);
nor U21969 (N_21969,N_17588,N_18953);
xor U21970 (N_21970,N_18221,N_19335);
and U21971 (N_21971,N_19850,N_17534);
xnor U21972 (N_21972,N_18157,N_19063);
nand U21973 (N_21973,N_19406,N_19038);
or U21974 (N_21974,N_19599,N_18022);
or U21975 (N_21975,N_19226,N_17821);
nand U21976 (N_21976,N_19474,N_18856);
nand U21977 (N_21977,N_19649,N_19292);
and U21978 (N_21978,N_18063,N_18225);
or U21979 (N_21979,N_19204,N_18018);
xor U21980 (N_21980,N_19994,N_19410);
xor U21981 (N_21981,N_17792,N_17651);
nand U21982 (N_21982,N_17752,N_18074);
xnor U21983 (N_21983,N_19654,N_17783);
nor U21984 (N_21984,N_17921,N_18665);
or U21985 (N_21985,N_17816,N_17825);
and U21986 (N_21986,N_19292,N_19130);
nand U21987 (N_21987,N_19269,N_19899);
or U21988 (N_21988,N_19463,N_19574);
and U21989 (N_21989,N_18222,N_18103);
or U21990 (N_21990,N_19139,N_18526);
nand U21991 (N_21991,N_17737,N_18988);
nor U21992 (N_21992,N_19985,N_18015);
nand U21993 (N_21993,N_19969,N_19544);
nand U21994 (N_21994,N_19834,N_19857);
xor U21995 (N_21995,N_18941,N_19700);
nand U21996 (N_21996,N_18126,N_19372);
or U21997 (N_21997,N_18598,N_17797);
nand U21998 (N_21998,N_19599,N_17718);
nor U21999 (N_21999,N_19224,N_18003);
nor U22000 (N_22000,N_19226,N_18845);
and U22001 (N_22001,N_17566,N_19762);
or U22002 (N_22002,N_19381,N_19719);
nand U22003 (N_22003,N_19038,N_17931);
and U22004 (N_22004,N_19179,N_17624);
nand U22005 (N_22005,N_19548,N_19188);
or U22006 (N_22006,N_17914,N_19247);
or U22007 (N_22007,N_17671,N_17612);
xor U22008 (N_22008,N_18089,N_19171);
nor U22009 (N_22009,N_17677,N_19271);
nor U22010 (N_22010,N_19846,N_19753);
or U22011 (N_22011,N_17706,N_18953);
xnor U22012 (N_22012,N_19512,N_19608);
nand U22013 (N_22013,N_18709,N_18597);
xnor U22014 (N_22014,N_19114,N_18918);
nand U22015 (N_22015,N_19126,N_19884);
or U22016 (N_22016,N_17810,N_19655);
and U22017 (N_22017,N_19668,N_18701);
xnor U22018 (N_22018,N_18171,N_19963);
and U22019 (N_22019,N_17737,N_19192);
xor U22020 (N_22020,N_17547,N_19255);
and U22021 (N_22021,N_18412,N_17981);
nor U22022 (N_22022,N_19739,N_18801);
xnor U22023 (N_22023,N_18412,N_18486);
xnor U22024 (N_22024,N_19977,N_19750);
xor U22025 (N_22025,N_19760,N_18248);
xor U22026 (N_22026,N_18053,N_19854);
and U22027 (N_22027,N_19894,N_17907);
or U22028 (N_22028,N_17685,N_18775);
and U22029 (N_22029,N_19352,N_17545);
nor U22030 (N_22030,N_17921,N_18790);
or U22031 (N_22031,N_18194,N_18915);
or U22032 (N_22032,N_18805,N_19646);
xor U22033 (N_22033,N_18227,N_17878);
xor U22034 (N_22034,N_18875,N_19108);
nand U22035 (N_22035,N_18486,N_18005);
nand U22036 (N_22036,N_18643,N_19586);
nor U22037 (N_22037,N_19828,N_19921);
or U22038 (N_22038,N_18815,N_18928);
xnor U22039 (N_22039,N_19351,N_17606);
nor U22040 (N_22040,N_18631,N_18704);
nand U22041 (N_22041,N_19210,N_19170);
nor U22042 (N_22042,N_19004,N_19450);
xor U22043 (N_22043,N_18497,N_19403);
and U22044 (N_22044,N_19354,N_19941);
nor U22045 (N_22045,N_19139,N_19954);
nand U22046 (N_22046,N_17938,N_18309);
or U22047 (N_22047,N_19823,N_19571);
and U22048 (N_22048,N_18835,N_18939);
nand U22049 (N_22049,N_19447,N_19638);
nand U22050 (N_22050,N_19703,N_18571);
and U22051 (N_22051,N_17793,N_18701);
nand U22052 (N_22052,N_19202,N_19272);
xnor U22053 (N_22053,N_19797,N_19856);
nor U22054 (N_22054,N_19817,N_17691);
xor U22055 (N_22055,N_19960,N_17982);
nor U22056 (N_22056,N_17902,N_18412);
xnor U22057 (N_22057,N_19602,N_19666);
or U22058 (N_22058,N_17761,N_19384);
and U22059 (N_22059,N_18393,N_17660);
and U22060 (N_22060,N_17716,N_19736);
nand U22061 (N_22061,N_18399,N_18029);
nor U22062 (N_22062,N_17876,N_18812);
or U22063 (N_22063,N_19057,N_17881);
xnor U22064 (N_22064,N_18328,N_19565);
nor U22065 (N_22065,N_18350,N_17765);
xnor U22066 (N_22066,N_18202,N_18101);
or U22067 (N_22067,N_17501,N_17689);
or U22068 (N_22068,N_18858,N_19775);
xnor U22069 (N_22069,N_17839,N_17793);
nor U22070 (N_22070,N_18636,N_18891);
nand U22071 (N_22071,N_17910,N_17923);
or U22072 (N_22072,N_18294,N_18490);
nor U22073 (N_22073,N_17627,N_17653);
xnor U22074 (N_22074,N_18815,N_18723);
nand U22075 (N_22075,N_18924,N_18685);
xor U22076 (N_22076,N_18411,N_18845);
nand U22077 (N_22077,N_18038,N_19341);
and U22078 (N_22078,N_19560,N_19273);
xor U22079 (N_22079,N_19366,N_19796);
and U22080 (N_22080,N_18722,N_19724);
and U22081 (N_22081,N_17862,N_19526);
nand U22082 (N_22082,N_17960,N_19471);
xnor U22083 (N_22083,N_17881,N_18276);
nor U22084 (N_22084,N_18140,N_18064);
xnor U22085 (N_22085,N_18646,N_19499);
nand U22086 (N_22086,N_19139,N_19987);
xor U22087 (N_22087,N_18300,N_17961);
or U22088 (N_22088,N_17858,N_18117);
xnor U22089 (N_22089,N_19663,N_19686);
xor U22090 (N_22090,N_19542,N_18029);
xor U22091 (N_22091,N_19145,N_17912);
xor U22092 (N_22092,N_19081,N_19303);
nand U22093 (N_22093,N_18841,N_18481);
nand U22094 (N_22094,N_18659,N_19967);
xnor U22095 (N_22095,N_19434,N_19980);
nor U22096 (N_22096,N_19424,N_19325);
nor U22097 (N_22097,N_17822,N_19172);
and U22098 (N_22098,N_18195,N_18252);
nand U22099 (N_22099,N_19331,N_18279);
xnor U22100 (N_22100,N_17733,N_18233);
nor U22101 (N_22101,N_19806,N_17820);
or U22102 (N_22102,N_18974,N_17586);
or U22103 (N_22103,N_19154,N_18381);
and U22104 (N_22104,N_19341,N_19694);
and U22105 (N_22105,N_18842,N_17726);
and U22106 (N_22106,N_17885,N_18577);
nand U22107 (N_22107,N_18871,N_18994);
nor U22108 (N_22108,N_18535,N_17649);
and U22109 (N_22109,N_18495,N_18761);
xor U22110 (N_22110,N_18119,N_18974);
or U22111 (N_22111,N_19620,N_18880);
xnor U22112 (N_22112,N_19363,N_17550);
nand U22113 (N_22113,N_19477,N_19002);
xnor U22114 (N_22114,N_18693,N_19900);
or U22115 (N_22115,N_19222,N_19602);
nand U22116 (N_22116,N_19229,N_19966);
nand U22117 (N_22117,N_18486,N_17763);
nand U22118 (N_22118,N_18254,N_19578);
xor U22119 (N_22119,N_18190,N_19337);
and U22120 (N_22120,N_18253,N_18635);
or U22121 (N_22121,N_18143,N_18775);
or U22122 (N_22122,N_19962,N_19177);
xor U22123 (N_22123,N_17894,N_18923);
nand U22124 (N_22124,N_17523,N_19016);
nand U22125 (N_22125,N_18021,N_19195);
or U22126 (N_22126,N_19282,N_19702);
nand U22127 (N_22127,N_18235,N_17792);
or U22128 (N_22128,N_19149,N_19444);
and U22129 (N_22129,N_17914,N_19847);
nand U22130 (N_22130,N_19837,N_17966);
nand U22131 (N_22131,N_19547,N_18746);
and U22132 (N_22132,N_19594,N_19482);
nor U22133 (N_22133,N_18741,N_18998);
xnor U22134 (N_22134,N_19978,N_18974);
nand U22135 (N_22135,N_19310,N_18654);
and U22136 (N_22136,N_19667,N_18298);
nand U22137 (N_22137,N_19513,N_19977);
and U22138 (N_22138,N_19933,N_19754);
and U22139 (N_22139,N_18897,N_17826);
xor U22140 (N_22140,N_19433,N_18631);
and U22141 (N_22141,N_17863,N_19466);
or U22142 (N_22142,N_18278,N_17698);
or U22143 (N_22143,N_17907,N_18772);
xnor U22144 (N_22144,N_18244,N_17931);
or U22145 (N_22145,N_18136,N_19909);
and U22146 (N_22146,N_19417,N_19485);
or U22147 (N_22147,N_18173,N_17578);
and U22148 (N_22148,N_18173,N_19355);
xor U22149 (N_22149,N_18073,N_19827);
or U22150 (N_22150,N_18830,N_19432);
or U22151 (N_22151,N_18166,N_18996);
and U22152 (N_22152,N_18560,N_18957);
xor U22153 (N_22153,N_17668,N_18323);
nor U22154 (N_22154,N_18766,N_18862);
and U22155 (N_22155,N_18861,N_19760);
and U22156 (N_22156,N_18300,N_18331);
or U22157 (N_22157,N_19200,N_19921);
nand U22158 (N_22158,N_17678,N_18532);
xnor U22159 (N_22159,N_19048,N_18823);
xnor U22160 (N_22160,N_19176,N_18493);
xnor U22161 (N_22161,N_19346,N_18693);
nor U22162 (N_22162,N_18484,N_19247);
and U22163 (N_22163,N_18100,N_19028);
or U22164 (N_22164,N_19669,N_18084);
and U22165 (N_22165,N_19008,N_18292);
and U22166 (N_22166,N_18476,N_18916);
xnor U22167 (N_22167,N_17756,N_19337);
xnor U22168 (N_22168,N_18158,N_19521);
nand U22169 (N_22169,N_19137,N_19436);
xor U22170 (N_22170,N_17884,N_19230);
xor U22171 (N_22171,N_18527,N_19291);
nor U22172 (N_22172,N_19509,N_19207);
and U22173 (N_22173,N_18351,N_19427);
or U22174 (N_22174,N_18674,N_19215);
nor U22175 (N_22175,N_19117,N_19576);
nand U22176 (N_22176,N_18395,N_19127);
and U22177 (N_22177,N_19787,N_19474);
and U22178 (N_22178,N_19211,N_17833);
or U22179 (N_22179,N_18858,N_18188);
nand U22180 (N_22180,N_18494,N_19979);
nand U22181 (N_22181,N_19437,N_19511);
and U22182 (N_22182,N_19536,N_17818);
nor U22183 (N_22183,N_19080,N_19325);
nor U22184 (N_22184,N_19652,N_19012);
or U22185 (N_22185,N_18505,N_17810);
nor U22186 (N_22186,N_18732,N_19351);
or U22187 (N_22187,N_19401,N_19099);
nor U22188 (N_22188,N_19123,N_18748);
or U22189 (N_22189,N_18080,N_17520);
nor U22190 (N_22190,N_19249,N_18022);
xor U22191 (N_22191,N_19379,N_18873);
xnor U22192 (N_22192,N_19433,N_18149);
or U22193 (N_22193,N_19605,N_19750);
and U22194 (N_22194,N_19190,N_19024);
nand U22195 (N_22195,N_18560,N_19321);
nor U22196 (N_22196,N_19462,N_18385);
or U22197 (N_22197,N_19510,N_19544);
nand U22198 (N_22198,N_18449,N_18370);
and U22199 (N_22199,N_19054,N_17513);
xor U22200 (N_22200,N_17919,N_17869);
nand U22201 (N_22201,N_19861,N_19953);
xnor U22202 (N_22202,N_18090,N_19174);
xor U22203 (N_22203,N_19315,N_19422);
xnor U22204 (N_22204,N_19724,N_18779);
nand U22205 (N_22205,N_18604,N_17630);
or U22206 (N_22206,N_19295,N_18378);
xor U22207 (N_22207,N_18764,N_17960);
or U22208 (N_22208,N_18857,N_18573);
or U22209 (N_22209,N_18165,N_18652);
and U22210 (N_22210,N_19261,N_19440);
or U22211 (N_22211,N_18267,N_18845);
nand U22212 (N_22212,N_19450,N_19144);
or U22213 (N_22213,N_19208,N_18317);
nor U22214 (N_22214,N_19235,N_18862);
nand U22215 (N_22215,N_18509,N_19666);
and U22216 (N_22216,N_17763,N_18622);
xnor U22217 (N_22217,N_18823,N_17616);
nand U22218 (N_22218,N_18643,N_19222);
and U22219 (N_22219,N_19841,N_18749);
and U22220 (N_22220,N_18697,N_17761);
and U22221 (N_22221,N_17681,N_19205);
and U22222 (N_22222,N_18065,N_19580);
nor U22223 (N_22223,N_19170,N_19077);
nor U22224 (N_22224,N_19231,N_18634);
nor U22225 (N_22225,N_18078,N_18881);
nand U22226 (N_22226,N_19554,N_18259);
and U22227 (N_22227,N_18012,N_19724);
nand U22228 (N_22228,N_17630,N_19914);
nand U22229 (N_22229,N_19220,N_19193);
and U22230 (N_22230,N_19630,N_18108);
nand U22231 (N_22231,N_18886,N_18423);
and U22232 (N_22232,N_19903,N_18576);
or U22233 (N_22233,N_18669,N_19009);
and U22234 (N_22234,N_17778,N_19259);
xnor U22235 (N_22235,N_18785,N_17840);
nand U22236 (N_22236,N_17993,N_18362);
xor U22237 (N_22237,N_18280,N_18215);
or U22238 (N_22238,N_19290,N_18214);
nand U22239 (N_22239,N_17565,N_17896);
nor U22240 (N_22240,N_18163,N_19657);
nand U22241 (N_22241,N_19184,N_17907);
xnor U22242 (N_22242,N_19059,N_18468);
or U22243 (N_22243,N_19017,N_18768);
xnor U22244 (N_22244,N_19306,N_19001);
or U22245 (N_22245,N_18572,N_18131);
nor U22246 (N_22246,N_18772,N_18920);
and U22247 (N_22247,N_18334,N_19591);
and U22248 (N_22248,N_19650,N_18469);
nor U22249 (N_22249,N_18407,N_17908);
nor U22250 (N_22250,N_19160,N_19880);
or U22251 (N_22251,N_19932,N_19794);
and U22252 (N_22252,N_18068,N_19633);
and U22253 (N_22253,N_17604,N_17981);
nor U22254 (N_22254,N_19067,N_18957);
nor U22255 (N_22255,N_19782,N_18089);
nand U22256 (N_22256,N_19543,N_17756);
and U22257 (N_22257,N_18952,N_19602);
nor U22258 (N_22258,N_18453,N_19527);
nand U22259 (N_22259,N_18779,N_18614);
and U22260 (N_22260,N_19054,N_19855);
and U22261 (N_22261,N_18551,N_18775);
nand U22262 (N_22262,N_19402,N_18870);
nand U22263 (N_22263,N_19285,N_18293);
and U22264 (N_22264,N_18457,N_19063);
or U22265 (N_22265,N_19365,N_18671);
and U22266 (N_22266,N_18729,N_19600);
nor U22267 (N_22267,N_19216,N_17978);
and U22268 (N_22268,N_19790,N_19997);
nand U22269 (N_22269,N_19622,N_17902);
nor U22270 (N_22270,N_18668,N_18334);
and U22271 (N_22271,N_17728,N_17805);
nor U22272 (N_22272,N_19042,N_19490);
nand U22273 (N_22273,N_17814,N_17653);
and U22274 (N_22274,N_19023,N_18549);
nand U22275 (N_22275,N_17884,N_19239);
xnor U22276 (N_22276,N_19863,N_19274);
nand U22277 (N_22277,N_19264,N_17758);
nand U22278 (N_22278,N_19400,N_18111);
and U22279 (N_22279,N_19370,N_18391);
and U22280 (N_22280,N_17608,N_19234);
xnor U22281 (N_22281,N_18513,N_17861);
and U22282 (N_22282,N_17575,N_17865);
nand U22283 (N_22283,N_17766,N_19306);
nor U22284 (N_22284,N_19487,N_19826);
and U22285 (N_22285,N_18804,N_17569);
nor U22286 (N_22286,N_19605,N_17933);
nor U22287 (N_22287,N_19106,N_18843);
or U22288 (N_22288,N_18625,N_17791);
nand U22289 (N_22289,N_17922,N_18551);
and U22290 (N_22290,N_18468,N_18389);
xnor U22291 (N_22291,N_18268,N_19491);
xor U22292 (N_22292,N_19045,N_18967);
nand U22293 (N_22293,N_18063,N_17845);
xnor U22294 (N_22294,N_18280,N_19531);
nor U22295 (N_22295,N_19942,N_18718);
and U22296 (N_22296,N_19531,N_18767);
and U22297 (N_22297,N_18397,N_18900);
nor U22298 (N_22298,N_18204,N_18715);
or U22299 (N_22299,N_19109,N_18645);
and U22300 (N_22300,N_18684,N_17727);
nand U22301 (N_22301,N_19568,N_17729);
and U22302 (N_22302,N_18270,N_19706);
nand U22303 (N_22303,N_18786,N_19814);
or U22304 (N_22304,N_18738,N_19649);
or U22305 (N_22305,N_18140,N_18243);
or U22306 (N_22306,N_19126,N_19253);
or U22307 (N_22307,N_17697,N_17561);
and U22308 (N_22308,N_18477,N_19844);
nor U22309 (N_22309,N_19602,N_18248);
xor U22310 (N_22310,N_19415,N_17940);
and U22311 (N_22311,N_17574,N_19951);
nor U22312 (N_22312,N_19910,N_17998);
nor U22313 (N_22313,N_19304,N_19982);
or U22314 (N_22314,N_17723,N_19649);
nand U22315 (N_22315,N_18406,N_18567);
or U22316 (N_22316,N_19991,N_19406);
nand U22317 (N_22317,N_19649,N_18249);
nand U22318 (N_22318,N_18738,N_17553);
xor U22319 (N_22319,N_18917,N_17733);
nor U22320 (N_22320,N_17872,N_19486);
xnor U22321 (N_22321,N_18854,N_19966);
nand U22322 (N_22322,N_17760,N_18243);
nor U22323 (N_22323,N_17725,N_19006);
nand U22324 (N_22324,N_19600,N_17700);
and U22325 (N_22325,N_19266,N_18383);
nor U22326 (N_22326,N_19341,N_18912);
nor U22327 (N_22327,N_18819,N_19360);
and U22328 (N_22328,N_17997,N_18344);
or U22329 (N_22329,N_18378,N_18776);
nand U22330 (N_22330,N_18261,N_17505);
and U22331 (N_22331,N_18508,N_17964);
nand U22332 (N_22332,N_19926,N_19754);
nand U22333 (N_22333,N_19593,N_19386);
nand U22334 (N_22334,N_18796,N_17640);
nand U22335 (N_22335,N_18156,N_17951);
nand U22336 (N_22336,N_18579,N_18766);
nor U22337 (N_22337,N_17923,N_19482);
and U22338 (N_22338,N_18251,N_19427);
xor U22339 (N_22339,N_18380,N_19690);
nand U22340 (N_22340,N_19802,N_19878);
xor U22341 (N_22341,N_19060,N_17990);
nand U22342 (N_22342,N_19839,N_18816);
nor U22343 (N_22343,N_19628,N_19685);
nand U22344 (N_22344,N_19133,N_19937);
and U22345 (N_22345,N_18984,N_19903);
nand U22346 (N_22346,N_18054,N_17804);
or U22347 (N_22347,N_18665,N_19658);
nor U22348 (N_22348,N_19567,N_19976);
nor U22349 (N_22349,N_19291,N_19926);
and U22350 (N_22350,N_17984,N_19906);
or U22351 (N_22351,N_18608,N_18240);
or U22352 (N_22352,N_17552,N_19436);
and U22353 (N_22353,N_18682,N_19970);
nor U22354 (N_22354,N_19053,N_19798);
or U22355 (N_22355,N_19671,N_18638);
nand U22356 (N_22356,N_17829,N_19379);
nand U22357 (N_22357,N_17836,N_19133);
and U22358 (N_22358,N_19770,N_18365);
nand U22359 (N_22359,N_18615,N_17651);
or U22360 (N_22360,N_18002,N_19354);
nor U22361 (N_22361,N_19208,N_19682);
or U22362 (N_22362,N_19709,N_18940);
and U22363 (N_22363,N_18807,N_18070);
or U22364 (N_22364,N_18136,N_18494);
or U22365 (N_22365,N_18300,N_18898);
or U22366 (N_22366,N_19501,N_18840);
and U22367 (N_22367,N_18115,N_18760);
nor U22368 (N_22368,N_19676,N_18420);
nand U22369 (N_22369,N_17820,N_18576);
and U22370 (N_22370,N_19414,N_19586);
or U22371 (N_22371,N_17530,N_19741);
nand U22372 (N_22372,N_19330,N_19112);
and U22373 (N_22373,N_17550,N_18008);
nand U22374 (N_22374,N_18200,N_19273);
xor U22375 (N_22375,N_17771,N_19494);
or U22376 (N_22376,N_17984,N_18528);
nor U22377 (N_22377,N_18703,N_18014);
or U22378 (N_22378,N_18425,N_19120);
xor U22379 (N_22379,N_18124,N_18645);
nand U22380 (N_22380,N_19979,N_19852);
nand U22381 (N_22381,N_19858,N_19614);
or U22382 (N_22382,N_19782,N_18486);
nor U22383 (N_22383,N_19066,N_18496);
and U22384 (N_22384,N_18809,N_18934);
or U22385 (N_22385,N_18622,N_18095);
or U22386 (N_22386,N_19341,N_18562);
or U22387 (N_22387,N_19785,N_18321);
or U22388 (N_22388,N_17560,N_17738);
xor U22389 (N_22389,N_19466,N_18152);
nand U22390 (N_22390,N_19299,N_18601);
and U22391 (N_22391,N_18852,N_19689);
xor U22392 (N_22392,N_18322,N_19508);
nor U22393 (N_22393,N_18296,N_18254);
nor U22394 (N_22394,N_19959,N_19643);
and U22395 (N_22395,N_19499,N_17734);
nand U22396 (N_22396,N_17764,N_18365);
or U22397 (N_22397,N_19296,N_19154);
xor U22398 (N_22398,N_17953,N_19870);
xor U22399 (N_22399,N_18987,N_18625);
or U22400 (N_22400,N_19082,N_18322);
nor U22401 (N_22401,N_18022,N_18767);
nand U22402 (N_22402,N_18828,N_19083);
xnor U22403 (N_22403,N_17804,N_18273);
xor U22404 (N_22404,N_18634,N_19021);
and U22405 (N_22405,N_19702,N_17737);
nand U22406 (N_22406,N_19395,N_19432);
nand U22407 (N_22407,N_17678,N_19501);
or U22408 (N_22408,N_17952,N_19640);
nor U22409 (N_22409,N_19164,N_18170);
nand U22410 (N_22410,N_19395,N_18050);
xor U22411 (N_22411,N_18102,N_18292);
nor U22412 (N_22412,N_18743,N_18358);
or U22413 (N_22413,N_18071,N_17855);
nand U22414 (N_22414,N_19925,N_19049);
nand U22415 (N_22415,N_19813,N_17837);
nor U22416 (N_22416,N_18140,N_19062);
nand U22417 (N_22417,N_19271,N_19016);
nor U22418 (N_22418,N_17595,N_19821);
nor U22419 (N_22419,N_18585,N_19430);
and U22420 (N_22420,N_18254,N_18419);
and U22421 (N_22421,N_18034,N_18421);
nand U22422 (N_22422,N_17674,N_19094);
and U22423 (N_22423,N_19302,N_17963);
nor U22424 (N_22424,N_19058,N_18488);
nor U22425 (N_22425,N_17916,N_19084);
xor U22426 (N_22426,N_18389,N_18571);
nand U22427 (N_22427,N_17974,N_18575);
and U22428 (N_22428,N_17672,N_19992);
xor U22429 (N_22429,N_18298,N_19747);
xnor U22430 (N_22430,N_19456,N_19035);
and U22431 (N_22431,N_18194,N_19461);
or U22432 (N_22432,N_18923,N_19458);
and U22433 (N_22433,N_18555,N_18110);
xnor U22434 (N_22434,N_19065,N_19831);
or U22435 (N_22435,N_18808,N_19497);
nand U22436 (N_22436,N_19595,N_17665);
nor U22437 (N_22437,N_19875,N_17520);
nand U22438 (N_22438,N_17674,N_19997);
xnor U22439 (N_22439,N_19407,N_19470);
or U22440 (N_22440,N_19012,N_18695);
or U22441 (N_22441,N_18892,N_18283);
nor U22442 (N_22442,N_18908,N_19066);
and U22443 (N_22443,N_18691,N_18259);
nand U22444 (N_22444,N_18105,N_18741);
nand U22445 (N_22445,N_19051,N_17734);
xnor U22446 (N_22446,N_19722,N_18901);
nand U22447 (N_22447,N_17731,N_18996);
or U22448 (N_22448,N_17630,N_17661);
and U22449 (N_22449,N_19887,N_19770);
nand U22450 (N_22450,N_19601,N_18060);
nor U22451 (N_22451,N_19616,N_18099);
nor U22452 (N_22452,N_18525,N_17530);
nor U22453 (N_22453,N_18888,N_18272);
nand U22454 (N_22454,N_19301,N_17909);
nand U22455 (N_22455,N_18066,N_18205);
and U22456 (N_22456,N_18233,N_18733);
nor U22457 (N_22457,N_17718,N_18474);
nor U22458 (N_22458,N_18478,N_18642);
or U22459 (N_22459,N_19091,N_19864);
or U22460 (N_22460,N_19306,N_18832);
nor U22461 (N_22461,N_18975,N_17708);
nand U22462 (N_22462,N_17871,N_19250);
or U22463 (N_22463,N_19252,N_19957);
nand U22464 (N_22464,N_18612,N_17751);
nor U22465 (N_22465,N_18952,N_19193);
or U22466 (N_22466,N_17806,N_18921);
nor U22467 (N_22467,N_19331,N_19826);
and U22468 (N_22468,N_17883,N_19895);
nand U22469 (N_22469,N_19871,N_19617);
nand U22470 (N_22470,N_19380,N_18817);
and U22471 (N_22471,N_19421,N_17679);
or U22472 (N_22472,N_17601,N_18814);
or U22473 (N_22473,N_18006,N_19862);
xnor U22474 (N_22474,N_19079,N_18313);
nand U22475 (N_22475,N_17695,N_18434);
nor U22476 (N_22476,N_19392,N_18053);
nand U22477 (N_22477,N_18651,N_18680);
nand U22478 (N_22478,N_19574,N_18636);
nand U22479 (N_22479,N_19427,N_17744);
xnor U22480 (N_22480,N_19031,N_18320);
or U22481 (N_22481,N_19879,N_19069);
or U22482 (N_22482,N_18056,N_17804);
and U22483 (N_22483,N_19180,N_18767);
and U22484 (N_22484,N_18299,N_18490);
nand U22485 (N_22485,N_18047,N_17704);
or U22486 (N_22486,N_17829,N_17860);
xnor U22487 (N_22487,N_19575,N_19452);
nor U22488 (N_22488,N_19234,N_18308);
xor U22489 (N_22489,N_19135,N_18765);
xnor U22490 (N_22490,N_17639,N_18926);
or U22491 (N_22491,N_17995,N_19095);
nor U22492 (N_22492,N_18680,N_17983);
nand U22493 (N_22493,N_18642,N_19762);
and U22494 (N_22494,N_18897,N_19354);
xor U22495 (N_22495,N_19541,N_17875);
xnor U22496 (N_22496,N_19440,N_18545);
nor U22497 (N_22497,N_18698,N_19978);
nor U22498 (N_22498,N_19049,N_19165);
and U22499 (N_22499,N_18687,N_18056);
and U22500 (N_22500,N_21968,N_20470);
xnor U22501 (N_22501,N_20829,N_21955);
nor U22502 (N_22502,N_21610,N_22136);
nand U22503 (N_22503,N_20720,N_20451);
nand U22504 (N_22504,N_20343,N_21650);
xnor U22505 (N_22505,N_22192,N_21326);
nand U22506 (N_22506,N_20770,N_20597);
xnor U22507 (N_22507,N_22279,N_21864);
and U22508 (N_22508,N_20792,N_20203);
or U22509 (N_22509,N_21839,N_20010);
nand U22510 (N_22510,N_20989,N_22332);
and U22511 (N_22511,N_21708,N_21841);
nor U22512 (N_22512,N_20675,N_21299);
nand U22513 (N_22513,N_21428,N_22320);
nand U22514 (N_22514,N_21586,N_20944);
nand U22515 (N_22515,N_22411,N_22082);
nor U22516 (N_22516,N_20861,N_20196);
and U22517 (N_22517,N_22057,N_20623);
xnor U22518 (N_22518,N_20701,N_21571);
or U22519 (N_22519,N_22339,N_22424);
or U22520 (N_22520,N_20715,N_21157);
or U22521 (N_22521,N_20606,N_20580);
nor U22522 (N_22522,N_22297,N_21877);
and U22523 (N_22523,N_22414,N_20906);
or U22524 (N_22524,N_20333,N_21035);
nand U22525 (N_22525,N_22277,N_21859);
nor U22526 (N_22526,N_20639,N_20846);
or U22527 (N_22527,N_22209,N_22150);
xor U22528 (N_22528,N_20005,N_21582);
nor U22529 (N_22529,N_21774,N_21477);
xnor U22530 (N_22530,N_20960,N_20555);
nand U22531 (N_22531,N_21833,N_20516);
or U22532 (N_22532,N_20473,N_21129);
and U22533 (N_22533,N_21419,N_22013);
or U22534 (N_22534,N_20922,N_21899);
xor U22535 (N_22535,N_20129,N_22474);
nor U22536 (N_22536,N_21797,N_20457);
nor U22537 (N_22537,N_21584,N_20250);
and U22538 (N_22538,N_21113,N_20444);
xnor U22539 (N_22539,N_21607,N_21259);
nand U22540 (N_22540,N_21238,N_21048);
nor U22541 (N_22541,N_21889,N_21735);
nand U22542 (N_22542,N_21053,N_21004);
or U22543 (N_22543,N_21284,N_20283);
or U22544 (N_22544,N_21310,N_20383);
nand U22545 (N_22545,N_20756,N_20244);
or U22546 (N_22546,N_20560,N_20130);
or U22547 (N_22547,N_20318,N_21837);
nand U22548 (N_22548,N_21231,N_20181);
and U22549 (N_22549,N_22184,N_21036);
or U22550 (N_22550,N_22387,N_20569);
and U22551 (N_22551,N_20324,N_21423);
xor U22552 (N_22552,N_21921,N_20465);
xnor U22553 (N_22553,N_22287,N_21105);
nor U22554 (N_22554,N_21093,N_20706);
or U22555 (N_22555,N_20440,N_20267);
or U22556 (N_22556,N_20665,N_22173);
nand U22557 (N_22557,N_20587,N_20084);
xor U22558 (N_22558,N_22103,N_20995);
nor U22559 (N_22559,N_20657,N_21167);
xor U22560 (N_22560,N_20036,N_21963);
xor U22561 (N_22561,N_20046,N_20059);
nor U22562 (N_22562,N_22153,N_20771);
and U22563 (N_22563,N_20215,N_22161);
xor U22564 (N_22564,N_20864,N_20360);
xor U22565 (N_22565,N_21433,N_21830);
nor U22566 (N_22566,N_21999,N_22243);
or U22567 (N_22567,N_21456,N_20610);
nand U22568 (N_22568,N_21075,N_20040);
nand U22569 (N_22569,N_20228,N_20000);
or U22570 (N_22570,N_21849,N_20206);
and U22571 (N_22571,N_20656,N_21572);
xor U22572 (N_22572,N_21645,N_21401);
and U22573 (N_22573,N_20627,N_22453);
and U22574 (N_22574,N_21926,N_20474);
and U22575 (N_22575,N_22015,N_22374);
nand U22576 (N_22576,N_22205,N_20028);
xnor U22577 (N_22577,N_20734,N_21384);
or U22578 (N_22578,N_21871,N_20790);
nand U22579 (N_22579,N_21215,N_20817);
nand U22580 (N_22580,N_20220,N_22347);
nand U22581 (N_22581,N_20305,N_20872);
or U22582 (N_22582,N_20593,N_22206);
xor U22583 (N_22583,N_21365,N_20344);
nand U22584 (N_22584,N_20877,N_21249);
and U22585 (N_22585,N_22189,N_21620);
nor U22586 (N_22586,N_22346,N_22442);
xor U22587 (N_22587,N_20402,N_20594);
nand U22588 (N_22588,N_21756,N_20831);
and U22589 (N_22589,N_22405,N_20827);
and U22590 (N_22590,N_21187,N_20522);
xnor U22591 (N_22591,N_21531,N_22475);
and U22592 (N_22592,N_22469,N_21768);
nor U22593 (N_22593,N_20868,N_21228);
xnor U22594 (N_22594,N_21826,N_22149);
and U22595 (N_22595,N_21183,N_20353);
nor U22596 (N_22596,N_21244,N_21011);
and U22597 (N_22597,N_22264,N_22027);
and U22598 (N_22598,N_21415,N_21654);
xor U22599 (N_22599,N_21574,N_20096);
xnor U22600 (N_22600,N_21553,N_22385);
or U22601 (N_22601,N_20149,N_21406);
xnor U22602 (N_22602,N_21630,N_20018);
xor U22603 (N_22603,N_21915,N_21308);
nor U22604 (N_22604,N_20117,N_22140);
and U22605 (N_22605,N_21647,N_20534);
xnor U22606 (N_22606,N_20915,N_20556);
or U22607 (N_22607,N_22289,N_20184);
xnor U22608 (N_22608,N_20363,N_22102);
or U22609 (N_22609,N_22185,N_20559);
and U22610 (N_22610,N_20050,N_22056);
or U22611 (N_22611,N_22412,N_21573);
nor U22612 (N_22612,N_21490,N_20808);
xnor U22613 (N_22613,N_22317,N_20069);
nor U22614 (N_22614,N_22489,N_21264);
or U22615 (N_22615,N_20854,N_20509);
xor U22616 (N_22616,N_22284,N_21634);
nand U22617 (N_22617,N_21332,N_21865);
or U22618 (N_22618,N_20057,N_22298);
nand U22619 (N_22619,N_20904,N_20009);
xor U22620 (N_22620,N_20497,N_20286);
or U22621 (N_22621,N_21937,N_21085);
nand U22622 (N_22622,N_20273,N_20246);
xor U22623 (N_22623,N_20681,N_21175);
xor U22624 (N_22624,N_22128,N_20382);
or U22625 (N_22625,N_20385,N_20595);
and U22626 (N_22626,N_21588,N_20869);
nor U22627 (N_22627,N_21812,N_22214);
and U22628 (N_22628,N_22213,N_20322);
xnor U22629 (N_22629,N_21217,N_20055);
and U22630 (N_22630,N_21098,N_21972);
or U22631 (N_22631,N_21711,N_20733);
or U22632 (N_22632,N_22377,N_20553);
nor U22633 (N_22633,N_20899,N_22420);
nand U22634 (N_22634,N_20685,N_20260);
nor U22635 (N_22635,N_21883,N_21136);
nand U22636 (N_22636,N_20930,N_21118);
nor U22637 (N_22637,N_20186,N_20162);
and U22638 (N_22638,N_21543,N_21455);
or U22639 (N_22639,N_20094,N_20784);
or U22640 (N_22640,N_21227,N_21663);
or U22641 (N_22641,N_20970,N_21143);
and U22642 (N_22642,N_21243,N_21717);
nor U22643 (N_22643,N_21581,N_21764);
xor U22644 (N_22644,N_22367,N_21931);
nand U22645 (N_22645,N_21470,N_20153);
xnor U22646 (N_22646,N_20079,N_22302);
nor U22647 (N_22647,N_22038,N_22017);
nand U22648 (N_22648,N_20448,N_20530);
nor U22649 (N_22649,N_22250,N_21448);
and U22650 (N_22650,N_21392,N_21947);
or U22651 (N_22651,N_21715,N_20034);
and U22652 (N_22652,N_21418,N_20718);
nor U22653 (N_22653,N_22222,N_20416);
or U22654 (N_22654,N_22418,N_20622);
or U22655 (N_22655,N_20799,N_21771);
and U22656 (N_22656,N_20401,N_22491);
or U22657 (N_22657,N_20932,N_22360);
or U22658 (N_22658,N_21686,N_20889);
xor U22659 (N_22659,N_21593,N_21924);
or U22660 (N_22660,N_20966,N_21861);
or U22661 (N_22661,N_21305,N_21255);
xnor U22662 (N_22662,N_20807,N_22309);
and U22663 (N_22663,N_21638,N_22416);
or U22664 (N_22664,N_21631,N_20158);
nor U22665 (N_22665,N_20048,N_22037);
nand U22666 (N_22666,N_20145,N_21328);
or U22667 (N_22667,N_21148,N_21981);
xor U22668 (N_22668,N_21144,N_21576);
nand U22669 (N_22669,N_22174,N_21226);
nor U22670 (N_22670,N_22340,N_20662);
and U22671 (N_22671,N_21655,N_22018);
or U22672 (N_22672,N_20883,N_21950);
xor U22673 (N_22673,N_22392,N_20330);
xnor U22674 (N_22674,N_21885,N_20390);
xor U22675 (N_22675,N_20982,N_21132);
and U22676 (N_22676,N_20658,N_21585);
and U22677 (N_22677,N_20564,N_22242);
or U22678 (N_22678,N_20631,N_21427);
and U22679 (N_22679,N_22050,N_20230);
and U22680 (N_22680,N_22101,N_20881);
xor U22681 (N_22681,N_20703,N_21635);
xnor U22682 (N_22682,N_20408,N_20066);
nor U22683 (N_22683,N_20654,N_22458);
nor U22684 (N_22684,N_22246,N_22182);
or U22685 (N_22685,N_20418,N_21876);
and U22686 (N_22686,N_20480,N_22443);
nor U22687 (N_22687,N_20241,N_20753);
nor U22688 (N_22688,N_20858,N_21128);
nor U22689 (N_22689,N_21090,N_20815);
nor U22690 (N_22690,N_20052,N_20996);
nand U22691 (N_22691,N_20663,N_21589);
nor U22692 (N_22692,N_20882,N_21109);
and U22693 (N_22693,N_20315,N_22343);
nand U22694 (N_22694,N_20940,N_20271);
nand U22695 (N_22695,N_20852,N_22468);
xor U22696 (N_22696,N_21554,N_20615);
or U22697 (N_22697,N_20362,N_22471);
or U22698 (N_22698,N_22473,N_22430);
and U22699 (N_22699,N_20527,N_20667);
or U22700 (N_22700,N_20572,N_20788);
xor U22701 (N_22701,N_22413,N_22244);
and U22702 (N_22702,N_21856,N_21653);
xnor U22703 (N_22703,N_20929,N_22219);
nor U22704 (N_22704,N_20098,N_21835);
xnor U22705 (N_22705,N_20163,N_22338);
or U22706 (N_22706,N_22399,N_22479);
and U22707 (N_22707,N_20958,N_22472);
nor U22708 (N_22708,N_21346,N_20496);
and U22709 (N_22709,N_22019,N_21808);
or U22710 (N_22710,N_21194,N_21102);
xor U22711 (N_22711,N_20350,N_20060);
nand U22712 (N_22712,N_20201,N_21832);
nor U22713 (N_22713,N_21524,N_20430);
xnor U22714 (N_22714,N_21528,N_20452);
or U22715 (N_22715,N_22492,N_22373);
nand U22716 (N_22716,N_21665,N_20056);
nor U22717 (N_22717,N_20584,N_20987);
nand U22718 (N_22718,N_22076,N_20684);
xor U22719 (N_22719,N_20287,N_20219);
nor U22720 (N_22720,N_20289,N_21480);
xnor U22721 (N_22721,N_20863,N_21037);
xnor U22722 (N_22722,N_20873,N_20157);
and U22723 (N_22723,N_21141,N_20937);
xor U22724 (N_22724,N_20062,N_21056);
or U22725 (N_22725,N_21606,N_20367);
nand U22726 (N_22726,N_20732,N_20397);
or U22727 (N_22727,N_21938,N_20874);
and U22728 (N_22728,N_21140,N_22075);
xor U22729 (N_22729,N_20336,N_21759);
nor U22730 (N_22730,N_21472,N_22180);
nor U22731 (N_22731,N_22078,N_22423);
or U22732 (N_22732,N_22324,N_21953);
nand U22733 (N_22733,N_20074,N_21060);
xor U22734 (N_22734,N_20635,N_20304);
or U22735 (N_22735,N_20678,N_20189);
or U22736 (N_22736,N_21439,N_21942);
nor U22737 (N_22737,N_22276,N_21626);
or U22738 (N_22738,N_20380,N_20222);
or U22739 (N_22739,N_21349,N_21760);
nand U22740 (N_22740,N_22063,N_20979);
and U22741 (N_22741,N_22168,N_21032);
nand U22742 (N_22742,N_21133,N_22208);
xnor U22743 (N_22743,N_20110,N_21221);
xor U22744 (N_22744,N_20562,N_20781);
and U22745 (N_22745,N_20338,N_21730);
nor U22746 (N_22746,N_22084,N_21006);
or U22747 (N_22747,N_21996,N_21555);
nor U22748 (N_22748,N_21860,N_21829);
xor U22749 (N_22749,N_20400,N_22135);
and U22750 (N_22750,N_20511,N_21624);
xnor U22751 (N_22751,N_20772,N_21569);
xor U22752 (N_22752,N_21747,N_20694);
nand U22753 (N_22753,N_21903,N_20185);
and U22754 (N_22754,N_21919,N_21746);
or U22755 (N_22755,N_20747,N_22196);
or U22756 (N_22756,N_20752,N_22022);
xor U22757 (N_22757,N_20133,N_20032);
and U22758 (N_22758,N_21211,N_21193);
and U22759 (N_22759,N_22254,N_20956);
nor U22760 (N_22760,N_21946,N_20563);
xnor U22761 (N_22761,N_21088,N_21458);
or U22762 (N_22762,N_20298,N_22402);
nor U22763 (N_22763,N_21280,N_21256);
nand U22764 (N_22764,N_20568,N_20467);
and U22765 (N_22765,N_22398,N_22456);
nor U22766 (N_22766,N_20475,N_21978);
nand U22767 (N_22767,N_20755,N_20766);
and U22768 (N_22768,N_22032,N_20765);
nand U22769 (N_22769,N_20471,N_21754);
or U22770 (N_22770,N_20081,N_20977);
and U22771 (N_22771,N_20017,N_20460);
xor U22772 (N_22772,N_21799,N_21975);
xor U22773 (N_22773,N_20312,N_20967);
or U22774 (N_22774,N_22293,N_20319);
nand U22775 (N_22775,N_20719,N_20113);
xnor U22776 (N_22776,N_20642,N_20576);
nor U22777 (N_22777,N_21266,N_20986);
xor U22778 (N_22778,N_20943,N_22466);
nand U22779 (N_22779,N_20221,N_21965);
xnor U22780 (N_22780,N_22134,N_21302);
nor U22781 (N_22781,N_21107,N_22375);
nor U22782 (N_22782,N_20945,N_20969);
nand U22783 (N_22783,N_22039,N_20895);
and U22784 (N_22784,N_20754,N_21373);
or U22785 (N_22785,N_21867,N_20591);
and U22786 (N_22786,N_20603,N_20006);
xnor U22787 (N_22787,N_20368,N_20963);
or U22788 (N_22788,N_21805,N_22341);
or U22789 (N_22789,N_22047,N_21566);
and U22790 (N_22790,N_21870,N_22422);
or U22791 (N_22791,N_21063,N_20302);
nand U22792 (N_22792,N_22349,N_20019);
or U22793 (N_22793,N_21149,N_20742);
nand U22794 (N_22794,N_21013,N_20714);
or U22795 (N_22795,N_21468,N_20972);
or U22796 (N_22796,N_20263,N_21763);
or U22797 (N_22797,N_20962,N_21785);
nand U22798 (N_22798,N_22241,N_20599);
or U22799 (N_22799,N_22106,N_21740);
xor U22800 (N_22800,N_20101,N_20750);
and U22801 (N_22801,N_21753,N_21913);
nand U22802 (N_22802,N_22253,N_22162);
or U22803 (N_22803,N_21251,N_21030);
nand U22804 (N_22804,N_21929,N_21485);
xnor U22805 (N_22805,N_20649,N_21135);
and U22806 (N_22806,N_21278,N_21847);
and U22807 (N_22807,N_21031,N_21636);
nor U22808 (N_22808,N_20538,N_20692);
and U22809 (N_22809,N_20022,N_21277);
xnor U22810 (N_22810,N_21475,N_22081);
xnor U22811 (N_22811,N_21154,N_20609);
nand U22812 (N_22812,N_21390,N_21274);
xnor U22813 (N_22813,N_21241,N_21377);
xor U22814 (N_22814,N_21461,N_22487);
nand U22815 (N_22815,N_20494,N_22478);
or U22816 (N_22816,N_22490,N_21750);
nand U22817 (N_22817,N_20151,N_21073);
or U22818 (N_22818,N_20693,N_20510);
nor U22819 (N_22819,N_21214,N_22294);
nand U22820 (N_22820,N_20106,N_21659);
or U22821 (N_22821,N_21202,N_21998);
xor U22822 (N_22822,N_22021,N_21324);
or U22823 (N_22823,N_20023,N_20187);
xor U22824 (N_22824,N_21570,N_20920);
nor U22825 (N_22825,N_22459,N_21151);
or U22826 (N_22826,N_22465,N_22157);
nor U22827 (N_22827,N_21186,N_21961);
xor U22828 (N_22828,N_21446,N_20903);
or U22829 (N_22829,N_21820,N_20833);
and U22830 (N_22830,N_22427,N_21873);
xnor U22831 (N_22831,N_21904,N_20499);
nor U22832 (N_22832,N_21890,N_22499);
xor U22833 (N_22833,N_21666,N_21059);
xor U22834 (N_22834,N_21068,N_21552);
xnor U22835 (N_22835,N_20124,N_20073);
nor U22836 (N_22836,N_20688,N_20389);
or U22837 (N_22837,N_20211,N_22389);
or U22838 (N_22838,N_22220,N_21608);
nand U22839 (N_22839,N_20652,N_21233);
nor U22840 (N_22840,N_21467,N_21721);
nor U22841 (N_22841,N_21959,N_20851);
xor U22842 (N_22842,N_22381,N_21535);
and U22843 (N_22843,N_21207,N_22262);
nor U22844 (N_22844,N_20994,N_20998);
nor U22845 (N_22845,N_21858,N_20650);
and U22846 (N_22846,N_21253,N_20142);
nand U22847 (N_22847,N_20307,N_21731);
xor U22848 (N_22848,N_21245,N_20843);
nand U22849 (N_22849,N_20504,N_21117);
or U22850 (N_22850,N_21234,N_21558);
xnor U22851 (N_22851,N_21982,N_21337);
nor U22852 (N_22852,N_22433,N_21361);
xnor U22853 (N_22853,N_20661,N_21615);
nand U22854 (N_22854,N_22200,N_20825);
or U22855 (N_22855,N_20377,N_21103);
or U22856 (N_22856,N_21844,N_21375);
or U22857 (N_22857,N_20331,N_21122);
nor U22858 (N_22858,N_20893,N_20953);
nand U22859 (N_22859,N_21616,N_22143);
nand U22860 (N_22860,N_21967,N_20341);
nor U22861 (N_22861,N_21185,N_21920);
nand U22862 (N_22862,N_20823,N_22316);
or U22863 (N_22863,N_21242,N_21008);
nand U22864 (N_22864,N_21521,N_21462);
or U22865 (N_22865,N_20762,N_20632);
or U22866 (N_22866,N_22095,N_21729);
xor U22867 (N_22867,N_20498,N_22086);
xnor U22868 (N_22868,N_22269,N_22040);
or U22869 (N_22869,N_22226,N_22098);
nand U22870 (N_22870,N_20712,N_20466);
nor U22871 (N_22871,N_21413,N_21235);
nor U22872 (N_22872,N_21720,N_22003);
and U22873 (N_22873,N_22278,N_21065);
xor U22874 (N_22874,N_20916,N_20348);
nor U22875 (N_22875,N_21334,N_21246);
nand U22876 (N_22876,N_20704,N_20410);
or U22877 (N_22877,N_20166,N_22218);
xor U22878 (N_22878,N_20648,N_20109);
nand U22879 (N_22879,N_20118,N_21159);
or U22880 (N_22880,N_22495,N_21525);
and U22881 (N_22881,N_20923,N_22292);
xor U22882 (N_22882,N_20178,N_21957);
or U22883 (N_22883,N_20892,N_20573);
and U22884 (N_22884,N_21252,N_20108);
nand U22885 (N_22885,N_21518,N_21994);
or U22886 (N_22886,N_21536,N_20396);
xor U22887 (N_22887,N_20155,N_20699);
and U22888 (N_22888,N_21956,N_20218);
xor U22889 (N_22889,N_21044,N_22034);
xnor U22890 (N_22890,N_20042,N_20745);
xnor U22891 (N_22891,N_20002,N_21629);
and U22892 (N_22892,N_21681,N_20454);
and U22893 (N_22893,N_21514,N_21466);
nand U22894 (N_22894,N_20936,N_21643);
nor U22895 (N_22895,N_21471,N_21679);
and U22896 (N_22896,N_21041,N_20778);
and U22897 (N_22897,N_20976,N_22255);
nor U22898 (N_22898,N_20141,N_20281);
and U22899 (N_22899,N_20696,N_20992);
or U22900 (N_22900,N_20413,N_21696);
xnor U22901 (N_22901,N_22122,N_21597);
and U22902 (N_22902,N_21991,N_21265);
nor U22903 (N_22903,N_20700,N_22072);
and U22904 (N_22904,N_22096,N_20223);
xnor U22905 (N_22905,N_20909,N_22146);
or U22906 (N_22906,N_21208,N_20512);
nand U22907 (N_22907,N_21678,N_21739);
nand U22908 (N_22908,N_20860,N_20280);
or U22909 (N_22909,N_21984,N_21360);
xnor U22910 (N_22910,N_22147,N_22364);
xor U22911 (N_22911,N_21137,N_21275);
nand U22912 (N_22912,N_21622,N_21197);
and U22913 (N_22913,N_22175,N_22325);
xnor U22914 (N_22914,N_22438,N_21120);
and U22915 (N_22915,N_21911,N_20469);
or U22916 (N_22916,N_20214,N_21866);
and U22917 (N_22917,N_20303,N_21064);
or U22918 (N_22918,N_21713,N_22391);
xnor U22919 (N_22919,N_21209,N_21447);
xor U22920 (N_22920,N_21166,N_21807);
nor U22921 (N_22921,N_20763,N_21822);
or U22922 (N_22922,N_21047,N_22327);
or U22923 (N_22923,N_21449,N_20359);
or U22924 (N_22924,N_21281,N_22434);
and U22925 (N_22925,N_21339,N_21939);
and U22926 (N_22926,N_22178,N_20182);
xnor U22927 (N_22927,N_20557,N_21707);
and U22928 (N_22928,N_21726,N_21500);
nor U22929 (N_22929,N_20361,N_20240);
or U22930 (N_22930,N_21761,N_20154);
or U22931 (N_22931,N_20849,N_20870);
xor U22932 (N_22932,N_21765,N_22151);
xor U22933 (N_22933,N_21491,N_20802);
nand U22934 (N_22934,N_22238,N_22144);
nand U22935 (N_22935,N_20455,N_20671);
or U22936 (N_22936,N_20835,N_21941);
or U22937 (N_22937,N_22171,N_21250);
xnor U22938 (N_22938,N_20099,N_21441);
or U22939 (N_22939,N_22137,N_21321);
xor U22940 (N_22940,N_22055,N_22221);
xor U22941 (N_22941,N_21049,N_21817);
nor U22942 (N_22942,N_22415,N_20489);
nor U22943 (N_22943,N_20404,N_20347);
or U22944 (N_22944,N_22477,N_20116);
xnor U22945 (N_22945,N_20150,N_21189);
or U22946 (N_22946,N_20826,N_21960);
xnor U22947 (N_22947,N_22328,N_21298);
xnor U22948 (N_22948,N_21517,N_20256);
nor U22949 (N_22949,N_20607,N_22148);
nor U22950 (N_22950,N_20552,N_21095);
and U22951 (N_22951,N_21496,N_21072);
nor U22952 (N_22952,N_21970,N_20857);
nor U22953 (N_22953,N_21722,N_21066);
nor U22954 (N_22954,N_21201,N_22300);
nor U22955 (N_22955,N_21343,N_22061);
or U22956 (N_22956,N_20030,N_22382);
nor U22957 (N_22957,N_21879,N_22104);
nor U22958 (N_22958,N_21380,N_20299);
nor U22959 (N_22959,N_21505,N_21345);
nor U22960 (N_22960,N_21893,N_21824);
or U22961 (N_22961,N_22357,N_21983);
nor U22962 (N_22962,N_20456,N_20604);
nor U22963 (N_22963,N_22230,N_21409);
xnor U22964 (N_22964,N_20605,N_20713);
nor U22965 (N_22965,N_21078,N_21744);
and U22966 (N_22966,N_20537,N_20964);
and U22967 (N_22967,N_21675,N_21862);
nand U22968 (N_22968,N_20337,N_20041);
nand U22969 (N_22969,N_20917,N_21532);
and U22970 (N_22970,N_21762,N_22194);
nor U22971 (N_22971,N_21502,N_20613);
or U22972 (N_22972,N_20737,N_20476);
and U22973 (N_22973,N_20617,N_20549);
or U22974 (N_22974,N_20391,N_21749);
nor U22975 (N_22975,N_22070,N_22476);
xor U22976 (N_22976,N_22069,N_20645);
xor U22977 (N_22977,N_20634,N_22363);
nand U22978 (N_22978,N_21641,N_20047);
or U22979 (N_22979,N_21379,N_20314);
nand U22980 (N_22980,N_20126,N_21827);
and U22981 (N_22981,N_21506,N_22449);
nor U22982 (N_22982,N_21892,N_21442);
nand U22983 (N_22983,N_21512,N_20698);
xor U22984 (N_22984,N_21752,N_20035);
and U22985 (N_22985,N_20679,N_21261);
and U22986 (N_22986,N_20004,N_21618);
nor U22987 (N_22987,N_20636,N_22002);
xnor U22988 (N_22988,N_21464,N_22112);
xnor U22989 (N_22989,N_20545,N_20097);
or U22990 (N_22990,N_22181,N_20975);
and U22991 (N_22991,N_22097,N_20247);
and U22992 (N_22992,N_20135,N_21925);
nand U22993 (N_22993,N_21640,N_20585);
and U22994 (N_22994,N_22030,N_21604);
nand U22995 (N_22995,N_20103,N_21271);
or U22996 (N_22996,N_20345,N_20209);
and U22997 (N_22997,N_20172,N_20407);
nor U22998 (N_22998,N_20248,N_21800);
nand U22999 (N_22999,N_20072,N_20156);
xnor U23000 (N_23000,N_21385,N_21935);
and U23001 (N_23001,N_22115,N_21993);
or U23002 (N_23002,N_20646,N_20769);
xor U23003 (N_23003,N_20890,N_22348);
and U23004 (N_23004,N_21676,N_20296);
nor U23005 (N_23005,N_22306,N_22187);
nand U23006 (N_23006,N_20690,N_21725);
nor U23007 (N_23007,N_22190,N_20279);
and U23008 (N_23008,N_21815,N_20143);
and U23009 (N_23009,N_20641,N_21523);
xor U23010 (N_23010,N_20683,N_21705);
xor U23011 (N_23011,N_21778,N_20458);
xor U23012 (N_23012,N_21091,N_20723);
nor U23013 (N_23013,N_21089,N_20600);
and U23014 (N_23014,N_20759,N_21178);
nand U23015 (N_23015,N_21394,N_20011);
nand U23016 (N_23016,N_21486,N_21702);
nand U23017 (N_23017,N_22383,N_20625);
xor U23018 (N_23018,N_21045,N_21656);
nand U23019 (N_23019,N_22195,N_22053);
or U23020 (N_23020,N_20164,N_20459);
xor U23021 (N_23021,N_21594,N_20640);
nor U23022 (N_23022,N_20914,N_22011);
nand U23023 (N_23023,N_20207,N_20676);
nor U23024 (N_23024,N_20406,N_20095);
xor U23025 (N_23025,N_22345,N_21077);
xor U23026 (N_23026,N_20245,N_22179);
nor U23027 (N_23027,N_21387,N_22005);
nand U23028 (N_23028,N_20394,N_21819);
nand U23029 (N_23029,N_20515,N_22186);
nand U23030 (N_23030,N_21438,N_21367);
nand U23031 (N_23031,N_20811,N_22342);
or U23032 (N_23032,N_21445,N_21369);
and U23033 (N_23033,N_20886,N_20952);
nor U23034 (N_23034,N_22406,N_21192);
or U23035 (N_23035,N_21453,N_22308);
xnor U23036 (N_23036,N_20411,N_21303);
or U23037 (N_23037,N_22113,N_20818);
and U23038 (N_23038,N_21727,N_21478);
nor U23039 (N_23039,N_22049,N_20340);
and U23040 (N_23040,N_21262,N_21509);
nand U23041 (N_23041,N_20743,N_21488);
or U23042 (N_23042,N_20926,N_22080);
xor U23043 (N_23043,N_20900,N_20217);
nand U23044 (N_23044,N_21304,N_22066);
nand U23045 (N_23045,N_21457,N_21270);
or U23046 (N_23046,N_20810,N_21682);
nor U23047 (N_23047,N_20637,N_21687);
and U23048 (N_23048,N_21165,N_21029);
nand U23049 (N_23049,N_21596,N_20717);
or U23050 (N_23050,N_21383,N_22170);
and U23051 (N_23051,N_20935,N_21450);
xnor U23052 (N_23052,N_20523,N_20351);
and U23053 (N_23053,N_21174,N_22496);
or U23054 (N_23054,N_22009,N_20148);
nor U23055 (N_23055,N_20236,N_20127);
xor U23056 (N_23056,N_22467,N_20789);
or U23057 (N_23057,N_21796,N_21992);
xor U23058 (N_23058,N_20029,N_20785);
nor U23059 (N_23059,N_20983,N_21591);
xor U23060 (N_23060,N_20999,N_20179);
nand U23061 (N_23061,N_21114,N_20880);
nand U23062 (N_23062,N_22159,N_21501);
or U23063 (N_23063,N_20828,N_21590);
nor U23064 (N_23064,N_20169,N_20137);
or U23065 (N_23065,N_22087,N_22099);
and U23066 (N_23066,N_20837,N_22158);
nor U23067 (N_23067,N_21218,N_22270);
nand U23068 (N_23068,N_20268,N_21171);
or U23069 (N_23069,N_22118,N_22239);
and U23070 (N_23070,N_20339,N_20254);
nand U23071 (N_23071,N_20139,N_21838);
or U23072 (N_23072,N_22386,N_20520);
nor U23073 (N_23073,N_21495,N_20574);
xnor U23074 (N_23074,N_21203,N_21100);
and U23075 (N_23075,N_22429,N_20668);
or U23076 (N_23076,N_21319,N_20354);
or U23077 (N_23077,N_20529,N_22046);
nor U23078 (N_23078,N_21420,N_20779);
nand U23079 (N_23079,N_20957,N_20266);
nand U23080 (N_23080,N_20253,N_20213);
and U23081 (N_23081,N_22461,N_20102);
nand U23082 (N_23082,N_20532,N_20123);
nor U23083 (N_23083,N_20729,N_21121);
xnor U23084 (N_23084,N_20016,N_21776);
and U23085 (N_23085,N_22172,N_22119);
nor U23086 (N_23086,N_20934,N_22261);
and U23087 (N_23087,N_20370,N_20212);
or U23088 (N_23088,N_22060,N_21125);
nor U23089 (N_23089,N_21613,N_20434);
nand U23090 (N_23090,N_21811,N_20809);
nand U23091 (N_23091,N_21086,N_22071);
nand U23092 (N_23092,N_20037,N_20093);
or U23093 (N_23093,N_21225,N_21024);
nor U23094 (N_23094,N_21741,N_22370);
and U23095 (N_23095,N_22441,N_22463);
or U23096 (N_23096,N_21444,N_20891);
nand U23097 (N_23097,N_22132,N_20188);
or U23098 (N_23098,N_21522,N_21964);
xor U23099 (N_23099,N_20820,N_21191);
nor U23100 (N_23100,N_21150,N_22268);
xnor U23101 (N_23101,N_21301,N_20533);
or U23102 (N_23102,N_22142,N_21426);
xor U23103 (N_23103,N_20689,N_21546);
or U23104 (N_23104,N_20481,N_21300);
nor U23105 (N_23105,N_20195,N_21895);
xnor U23106 (N_23106,N_21980,N_21196);
or U23107 (N_23107,N_22454,N_22188);
or U23108 (N_23108,N_22355,N_22283);
or U23109 (N_23109,N_22212,N_21683);
nor U23110 (N_23110,N_21909,N_21540);
or U23111 (N_23111,N_20758,N_22323);
nor U23112 (N_23112,N_20077,N_22353);
nand U23113 (N_23113,N_21483,N_21314);
xor U23114 (N_23114,N_21212,N_21793);
and U23115 (N_23115,N_21079,N_22362);
nor U23116 (N_23116,N_21276,N_21944);
xnor U23117 (N_23117,N_21660,N_20705);
and U23118 (N_23118,N_20954,N_22154);
nand U23119 (N_23119,N_21697,N_20168);
nand U23120 (N_23120,N_20446,N_20647);
nand U23121 (N_23121,N_20087,N_22371);
xnor U23122 (N_23122,N_20373,N_20008);
nor U23123 (N_23123,N_21083,N_21504);
nand U23124 (N_23124,N_22252,N_21974);
and U23125 (N_23125,N_21061,N_20951);
or U23126 (N_23126,N_21498,N_21139);
nand U23127 (N_23127,N_21777,N_20990);
nand U23128 (N_23128,N_22435,N_20767);
nor U23129 (N_23129,N_21039,N_22207);
and U23130 (N_23130,N_22417,N_21318);
nor U23131 (N_23131,N_21602,N_21556);
nor U23132 (N_23132,N_21232,N_21476);
or U23133 (N_23133,N_21766,N_22237);
nand U23134 (N_23134,N_22227,N_21026);
nand U23135 (N_23135,N_22031,N_21434);
nor U23136 (N_23136,N_21547,N_20845);
nand U23137 (N_23137,N_21292,N_20061);
xnor U23138 (N_23138,N_20738,N_21745);
nor U23139 (N_23139,N_21916,N_20659);
nor U23140 (N_23140,N_21146,N_21734);
nand U23141 (N_23141,N_22322,N_22202);
nor U23142 (N_23142,N_20327,N_20746);
nand U23143 (N_23143,N_22074,N_21632);
or U23144 (N_23144,N_20797,N_20415);
xnor U23145 (N_23145,N_21359,N_21912);
xor U23146 (N_23146,N_21138,N_21987);
or U23147 (N_23147,N_20392,N_21131);
nor U23148 (N_23148,N_21648,N_21254);
nor U23149 (N_23149,N_22359,N_22068);
and U23150 (N_23150,N_20387,N_22311);
or U23151 (N_23151,N_21327,N_21979);
nor U23152 (N_23152,N_20782,N_20655);
nor U23153 (N_23153,N_20366,N_21863);
or U23154 (N_23154,N_22160,N_20501);
or U23155 (N_23155,N_21810,N_21000);
and U23156 (N_23156,N_21670,N_20760);
xnor U23157 (N_23157,N_20628,N_20170);
or U23158 (N_23158,N_20941,N_20071);
xor U23159 (N_23159,N_20120,N_20290);
nand U23160 (N_23160,N_22012,N_22281);
or U23161 (N_23161,N_21311,N_20971);
or U23162 (N_23162,N_21351,N_22033);
xor U23163 (N_23163,N_20378,N_22145);
nor U23164 (N_23164,N_20379,N_22067);
and U23165 (N_23165,N_22093,N_20836);
and U23166 (N_23166,N_20672,N_20089);
and U23167 (N_23167,N_20669,N_21995);
nand U23168 (N_23168,N_21633,N_22452);
nor U23169 (N_23169,N_21732,N_21548);
or U23170 (N_23170,N_20938,N_20426);
nand U23171 (N_23171,N_20748,N_21736);
nand U23172 (N_23172,N_20428,N_22282);
xnor U23173 (N_23173,N_20317,N_21484);
and U23174 (N_23174,N_20100,N_20138);
nand U23175 (N_23175,N_20695,N_20356);
nor U23176 (N_23176,N_21709,N_20258);
or U23177 (N_23177,N_22217,N_21551);
xor U23178 (N_23178,N_20259,N_21595);
nor U23179 (N_23179,N_20038,N_21775);
nor U23180 (N_23180,N_20357,N_21080);
nor U23181 (N_23181,N_20332,N_22042);
nor U23182 (N_23182,N_21184,N_20291);
or U23183 (N_23183,N_22307,N_20464);
or U23184 (N_23184,N_21350,N_20051);
nor U23185 (N_23185,N_20293,N_21070);
xor U23186 (N_23186,N_20284,N_21001);
or U23187 (N_23187,N_22120,N_22403);
nor U23188 (N_23188,N_22029,N_22265);
nor U23189 (N_23189,N_20269,N_21479);
xnor U23190 (N_23190,N_21087,N_21881);
xor U23191 (N_23191,N_20546,N_21286);
xnor U23192 (N_23192,N_20558,N_20535);
nand U23193 (N_23193,N_20461,N_22428);
or U23194 (N_23194,N_21043,N_22043);
nor U23195 (N_23195,N_20757,N_20136);
nand U23196 (N_23196,N_21003,N_21076);
xor U23197 (N_23197,N_20409,N_21598);
nor U23198 (N_23198,N_21742,N_21055);
nor U23199 (N_23199,N_21436,N_20014);
nor U23200 (N_23200,N_22274,N_20159);
xor U23201 (N_23201,N_22020,N_20911);
nor U23202 (N_23202,N_22024,N_21868);
and U23203 (N_23203,N_20592,N_21719);
nor U23204 (N_23204,N_21357,N_20794);
nor U23205 (N_23205,N_21850,N_20633);
nor U23206 (N_23206,N_21130,N_21407);
and U23207 (N_23207,N_22409,N_20208);
or U23208 (N_23208,N_20483,N_21333);
xor U23209 (N_23209,N_20618,N_21158);
nand U23210 (N_23210,N_21012,N_21789);
nor U23211 (N_23211,N_20544,N_21071);
xnor U23212 (N_23212,N_21580,N_21605);
and U23213 (N_23213,N_21758,N_21025);
nor U23214 (N_23214,N_20306,N_20866);
nor U23215 (N_23215,N_20887,N_20988);
xnor U23216 (N_23216,N_21344,N_20575);
nor U23217 (N_23217,N_21404,N_21529);
and U23218 (N_23218,N_20776,N_21239);
xnor U23219 (N_23219,N_20547,N_22026);
nor U23220 (N_23220,N_21698,N_20950);
nor U23221 (N_23221,N_21099,N_22198);
and U23222 (N_23222,N_22065,N_21544);
nor U23223 (N_23223,N_20565,N_20879);
xnor U23224 (N_23224,N_21923,N_20277);
nand U23225 (N_23225,N_20044,N_21127);
and U23226 (N_23226,N_20068,N_21537);
or U23227 (N_23227,N_22191,N_21156);
and U23228 (N_23228,N_21465,N_21403);
or U23229 (N_23229,N_22141,N_20482);
xnor U23230 (N_23230,N_21412,N_20165);
nor U23231 (N_23231,N_21397,N_20342);
nor U23232 (N_23232,N_21691,N_21028);
and U23233 (N_23233,N_20691,N_20805);
nand U23234 (N_23234,N_20134,N_20132);
nor U23235 (N_23235,N_20346,N_20980);
or U23236 (N_23236,N_20583,N_22138);
xnor U23237 (N_23237,N_21770,N_21482);
nand U23238 (N_23238,N_21293,N_21644);
xor U23239 (N_23239,N_20611,N_21493);
nor U23240 (N_23240,N_21354,N_20326);
and U23241 (N_23241,N_21353,N_21123);
xor U23242 (N_23242,N_20436,N_22169);
xor U23243 (N_23243,N_22044,N_22321);
nor U23244 (N_23244,N_22203,N_21587);
xnor U23245 (N_23245,N_21042,N_20783);
or U23246 (N_23246,N_20374,N_22299);
xnor U23247 (N_23247,N_21381,N_21692);
nand U23248 (N_23248,N_22133,N_20791);
or U23249 (N_23249,N_20525,N_21542);
xnor U23250 (N_23250,N_22152,N_21355);
nor U23251 (N_23251,N_20152,N_21283);
xnor U23252 (N_23252,N_20571,N_20442);
or U23253 (N_23253,N_20295,N_22290);
and U23254 (N_23254,N_21828,N_20644);
and U23255 (N_23255,N_21814,N_20075);
nor U23256 (N_23256,N_21519,N_20076);
or U23257 (N_23257,N_20997,N_20015);
nor U23258 (N_23258,N_20981,N_20842);
or U23259 (N_23259,N_22445,N_20910);
nand U23260 (N_23260,N_21115,N_20232);
nor U23261 (N_23261,N_22313,N_21481);
nand U23262 (N_23262,N_20619,N_21843);
xnor U23263 (N_23263,N_21907,N_20602);
and U23264 (N_23264,N_21034,N_22483);
and U23265 (N_23265,N_21152,N_21757);
xor U23266 (N_23266,N_21395,N_20550);
and U23267 (N_23267,N_20227,N_21393);
and U23268 (N_23268,N_22361,N_22197);
nor U23269 (N_23269,N_22028,N_21410);
or U23270 (N_23270,N_22114,N_20832);
xnor U23271 (N_23271,N_21282,N_21853);
nor U23272 (N_23272,N_22365,N_21795);
or U23273 (N_23273,N_20687,N_21172);
xor U23274 (N_23274,N_20567,N_21062);
and U23275 (N_23275,N_22085,N_22493);
and U23276 (N_23276,N_20581,N_21296);
and U23277 (N_23277,N_21336,N_22004);
nor U23278 (N_23278,N_21723,N_22352);
xnor U23279 (N_23279,N_21783,N_20310);
and U23280 (N_23280,N_21527,N_22240);
and U23281 (N_23281,N_21378,N_21142);
nor U23282 (N_23282,N_22092,N_20974);
and U23283 (N_23283,N_21804,N_20885);
xor U23284 (N_23284,N_22446,N_20848);
xor U23285 (N_23285,N_21857,N_22488);
or U23286 (N_23286,N_21917,N_22263);
or U23287 (N_23287,N_20243,N_20620);
and U23288 (N_23288,N_22390,N_20548);
and U23289 (N_23289,N_22223,N_21494);
xor U23290 (N_23290,N_21210,N_21908);
nand U23291 (N_23291,N_20224,N_22251);
nor U23292 (N_23292,N_21932,N_20147);
xnor U23293 (N_23293,N_22470,N_20536);
or U23294 (N_23294,N_22286,N_22394);
nand U23295 (N_23295,N_20205,N_21792);
nand U23296 (N_23296,N_22023,N_20173);
or U23297 (N_23297,N_20897,N_21780);
or U23298 (N_23298,N_20316,N_20335);
xor U23299 (N_23299,N_20420,N_20739);
nand U23300 (N_23300,N_20255,N_20526);
xnor U23301 (N_23301,N_21695,N_21342);
or U23302 (N_23302,N_22378,N_22494);
nand U23303 (N_23303,N_21190,N_21724);
xnor U23304 (N_23304,N_21347,N_21279);
xnor U23305 (N_23305,N_22272,N_21845);
and U23306 (N_23306,N_21704,N_21110);
xnor U23307 (N_23307,N_21652,N_22124);
nor U23308 (N_23308,N_20107,N_20463);
nand U23309 (N_23309,N_20122,N_21372);
and U23310 (N_23310,N_21575,N_21451);
xnor U23311 (N_23311,N_21545,N_22419);
and U23312 (N_23312,N_20865,N_20007);
or U23313 (N_23313,N_20183,N_20955);
or U23314 (N_23314,N_21674,N_20021);
or U23315 (N_23315,N_22183,N_20912);
xnor U23316 (N_23316,N_21429,N_21330);
xor U23317 (N_23317,N_22079,N_20856);
nor U23318 (N_23318,N_21943,N_20425);
and U23319 (N_23319,N_22457,N_20774);
nor U23320 (N_23320,N_22204,N_21313);
nor U23321 (N_23321,N_22330,N_20433);
xnor U23322 (N_23322,N_20626,N_21316);
nor U23323 (N_23323,N_20438,N_20517);
nand U23324 (N_23324,N_20670,N_21651);
or U23325 (N_23325,N_20736,N_21473);
or U23326 (N_23326,N_20450,N_20830);
xnor U23327 (N_23327,N_20894,N_22165);
and U23328 (N_23328,N_20519,N_22073);
and U23329 (N_23329,N_21699,N_21773);
nor U23330 (N_23330,N_21440,N_20128);
or U23331 (N_23331,N_22234,N_21153);
nand U23332 (N_23332,N_21818,N_21688);
xor U23333 (N_23333,N_20801,N_20834);
nor U23334 (N_23334,N_20878,N_20959);
and U23335 (N_23335,N_22455,N_22232);
xnor U23336 (N_23336,N_22088,N_21949);
nor U23337 (N_23337,N_20067,N_22090);
and U23338 (N_23338,N_21402,N_20086);
xor U23339 (N_23339,N_21834,N_20105);
xor U23340 (N_23340,N_20740,N_22314);
xor U23341 (N_23341,N_20787,N_22333);
nor U23342 (N_23342,N_21539,N_21728);
nor U23343 (N_23343,N_22376,N_20194);
and U23344 (N_23344,N_21204,N_21164);
or U23345 (N_23345,N_22109,N_21612);
nor U23346 (N_23346,N_21492,N_22125);
and U23347 (N_23347,N_21331,N_21672);
nor U23348 (N_23348,N_21195,N_22396);
and U23349 (N_23349,N_21469,N_20643);
xnor U23350 (N_23350,N_21269,N_21559);
xor U23351 (N_23351,N_20518,N_20764);
or U23352 (N_23352,N_21906,N_21668);
nand U23353 (N_23353,N_20479,N_22083);
or U23354 (N_23354,N_22064,N_21364);
nand U23355 (N_23355,N_20355,N_21182);
and U23356 (N_23356,N_22110,N_20506);
nand U23357 (N_23357,N_21971,N_22008);
nand U23358 (N_23358,N_20727,N_21294);
and U23359 (N_23359,N_21779,N_21329);
xnor U23360 (N_23360,N_21583,N_20908);
nand U23361 (N_23361,N_22285,N_20039);
nor U23362 (N_23362,N_20612,N_21291);
xnor U23363 (N_23363,N_21289,N_22010);
and U23364 (N_23364,N_21701,N_20447);
nor U23365 (N_23365,N_22210,N_21382);
nand U23366 (N_23366,N_20598,N_22448);
xnor U23367 (N_23367,N_21051,N_22177);
or U23368 (N_23368,N_20192,N_21989);
xnor U23369 (N_23369,N_20078,N_22315);
and U23370 (N_23370,N_20231,N_21119);
nand U23371 (N_23371,N_21169,N_21180);
nand U23372 (N_23372,N_22404,N_20238);
nand U23373 (N_23373,N_20608,N_22305);
nor U23374 (N_23374,N_21021,N_20708);
or U23375 (N_23375,N_21023,N_21541);
and U23376 (N_23376,N_20329,N_20973);
xor U23377 (N_23377,N_20309,N_21625);
or U23378 (N_23378,N_21934,N_21018);
nand U23379 (N_23379,N_22166,N_21199);
xor U23380 (N_23380,N_22215,N_21046);
xnor U23381 (N_23381,N_21463,N_21854);
xnor U23382 (N_23382,N_22266,N_21786);
and U23383 (N_23383,N_21703,N_22126);
nand U23384 (N_23384,N_20722,N_21669);
nand U23385 (N_23385,N_21813,N_20803);
or U23386 (N_23386,N_22048,N_20200);
xor U23387 (N_23387,N_20896,N_20091);
and U23388 (N_23388,N_20726,N_20931);
and U23389 (N_23389,N_21973,N_21966);
or U23390 (N_23390,N_21816,N_21787);
xnor U23391 (N_23391,N_20614,N_21206);
nand U23392 (N_23392,N_21599,N_20677);
nand U23393 (N_23393,N_21673,N_22498);
and U23394 (N_23394,N_20651,N_21295);
or U23395 (N_23395,N_22267,N_21335);
nor U23396 (N_23396,N_20796,N_22193);
and U23397 (N_23397,N_21014,N_20429);
or U23398 (N_23398,N_21664,N_20919);
nor U23399 (N_23399,N_20175,N_20539);
xnor U23400 (N_23400,N_21914,N_21052);
or U23401 (N_23401,N_21340,N_21533);
and U23402 (N_23402,N_21936,N_21508);
nand U23403 (N_23403,N_20445,N_21116);
nor U23404 (N_23404,N_21693,N_21323);
nand U23405 (N_23405,N_21416,N_21200);
nand U23406 (N_23406,N_20024,N_21155);
xor U23407 (N_23407,N_21106,N_20673);
nand U23408 (N_23408,N_20441,N_20844);
and U23409 (N_23409,N_20721,N_21905);
nand U23410 (N_23410,N_20616,N_20053);
and U23411 (N_23411,N_20800,N_21460);
nor U23412 (N_23412,N_20589,N_21884);
or U23413 (N_23413,N_21499,N_22105);
or U23414 (N_23414,N_21430,N_20088);
nand U23415 (N_23415,N_20140,N_22372);
or U23416 (N_23416,N_20570,N_21609);
nor U23417 (N_23417,N_21578,N_20949);
or U23418 (N_23418,N_20131,N_21662);
and U23419 (N_23419,N_22245,N_22224);
xor U23420 (N_23420,N_20798,N_20358);
nand U23421 (N_23421,N_20321,N_21038);
and U23422 (N_23422,N_20492,N_21160);
nor U23423 (N_23423,N_21623,N_21258);
nor U23424 (N_23424,N_20058,N_22089);
or U23425 (N_23425,N_21368,N_20507);
or U23426 (N_23426,N_20180,N_21325);
or U23427 (N_23427,N_20045,N_21922);
nand U23428 (N_23428,N_22007,N_21743);
nand U23429 (N_23429,N_21213,N_21179);
and U23430 (N_23430,N_20210,N_22393);
and U23431 (N_23431,N_21454,N_21869);
nand U23432 (N_23432,N_20928,N_22016);
nor U23433 (N_23433,N_22407,N_21806);
nand U23434 (N_23434,N_22248,N_21894);
or U23435 (N_23435,N_22337,N_21738);
nand U23436 (N_23436,N_20216,N_21755);
nand U23437 (N_23437,N_21082,N_21168);
nand U23438 (N_23438,N_20237,N_22397);
nor U23439 (N_23439,N_21802,N_22236);
and U23440 (N_23440,N_21712,N_21094);
nor U23441 (N_23441,N_20054,N_21287);
xnor U23442 (N_23442,N_20090,N_20064);
or U23443 (N_23443,N_21985,N_22091);
or U23444 (N_23444,N_21374,N_21538);
xor U23445 (N_23445,N_21366,N_20349);
nand U23446 (N_23446,N_20488,N_22130);
nor U23447 (N_23447,N_21408,N_20424);
or U23448 (N_23448,N_21005,N_20292);
nand U23449 (N_23449,N_21951,N_20543);
or U23450 (N_23450,N_21515,N_20898);
and U23451 (N_23451,N_21896,N_20741);
xnor U23452 (N_23452,N_21422,N_22041);
nand U23453 (N_23453,N_22384,N_20371);
nor U23454 (N_23454,N_20773,N_21952);
or U23455 (N_23455,N_20795,N_20235);
nand U23456 (N_23456,N_20502,N_21096);
or U23457 (N_23457,N_20566,N_21126);
xnor U23458 (N_23458,N_20422,N_21338);
nor U23459 (N_23459,N_20393,N_22395);
or U23460 (N_23460,N_21050,N_21163);
xor U23461 (N_23461,N_22129,N_21716);
nand U23462 (N_23462,N_21285,N_20775);
nand U23463 (N_23463,N_20398,N_20288);
and U23464 (N_23464,N_22410,N_20043);
xnor U23465 (N_23465,N_20751,N_20524);
xnor U23466 (N_23466,N_22288,N_20294);
nand U23467 (N_23467,N_21714,N_20432);
nor U23468 (N_23468,N_22350,N_20001);
nand U23469 (N_23469,N_21489,N_22062);
nor U23470 (N_23470,N_20697,N_21224);
or U23471 (N_23471,N_21878,N_21341);
xor U23472 (N_23472,N_22275,N_22054);
and U23473 (N_23473,N_20308,N_21677);
nor U23474 (N_23474,N_21297,N_21487);
and U23475 (N_23475,N_20487,N_22450);
nand U23476 (N_23476,N_21162,N_20323);
nor U23477 (N_23477,N_21791,N_21371);
nor U23478 (N_23478,N_22211,N_21809);
and U23479 (N_23479,N_21400,N_21557);
or U23480 (N_23480,N_21948,N_22045);
nand U23481 (N_23481,N_21986,N_21022);
nor U23482 (N_23482,N_21927,N_20257);
and U23483 (N_23483,N_20744,N_20629);
nand U23484 (N_23484,N_20435,N_20682);
xnor U23485 (N_23485,N_21511,N_21579);
or U23486 (N_23486,N_20768,N_20918);
xnor U23487 (N_23487,N_21352,N_20660);
nand U23488 (N_23488,N_20376,N_20710);
and U23489 (N_23489,N_20225,N_21425);
and U23490 (N_23490,N_20521,N_20161);
nor U23491 (N_23491,N_21642,N_20561);
or U23492 (N_23492,N_21619,N_22139);
nor U23493 (N_23493,N_21821,N_21836);
and U23494 (N_23494,N_21312,N_22426);
nor U23495 (N_23495,N_20160,N_20364);
or U23496 (N_23496,N_21534,N_21901);
xnor U23497 (N_23497,N_21309,N_20198);
or U23498 (N_23498,N_21432,N_21794);
nand U23499 (N_23499,N_20814,N_21851);
nand U23500 (N_23500,N_20125,N_20033);
and U23501 (N_23501,N_20477,N_20824);
and U23502 (N_23502,N_20369,N_20027);
nor U23503 (N_23503,N_22379,N_21017);
or U23504 (N_23504,N_20819,N_20111);
and U23505 (N_23505,N_21657,N_22356);
xor U23506 (N_23506,N_22001,N_21417);
nor U23507 (N_23507,N_21396,N_22199);
xor U23508 (N_23508,N_21737,N_22368);
or U23509 (N_23509,N_21263,N_20020);
or U23510 (N_23510,N_21886,N_21388);
nand U23511 (N_23511,N_20297,N_20541);
and U23512 (N_23512,N_21273,N_20114);
and U23513 (N_23513,N_21621,N_20199);
nor U23514 (N_23514,N_20531,N_21671);
or U23515 (N_23515,N_22431,N_22331);
xnor U23516 (N_23516,N_22006,N_21222);
and U23517 (N_23517,N_22167,N_21054);
nor U23518 (N_23518,N_22464,N_22231);
nor U23519 (N_23519,N_20300,N_22296);
and U23520 (N_23520,N_20841,N_21928);
and U23521 (N_23521,N_20403,N_21520);
xnor U23522 (N_23522,N_21081,N_21842);
and U23523 (N_23523,N_21474,N_21370);
xnor U23524 (N_23524,N_21628,N_20925);
xor U23525 (N_23525,N_21040,N_22485);
and U23526 (N_23526,N_21627,N_20012);
nor U23527 (N_23527,N_21399,N_21010);
xor U23528 (N_23528,N_21710,N_21198);
and U23529 (N_23529,N_21855,N_20204);
xor U23530 (N_23530,N_21846,N_21307);
nor U23531 (N_23531,N_21104,N_22077);
and U23532 (N_23532,N_20578,N_21782);
and U23533 (N_23533,N_22484,N_22051);
nand U23534 (N_23534,N_20702,N_22235);
xnor U23535 (N_23535,N_20514,N_20026);
or U23536 (N_23536,N_21825,N_20875);
nand U23537 (N_23537,N_20577,N_20709);
and U23538 (N_23538,N_20490,N_20850);
nor U23539 (N_23539,N_21831,N_21205);
nand U23540 (N_23540,N_21322,N_20313);
or U23541 (N_23541,N_20821,N_21389);
or U23542 (N_23542,N_21790,N_20554);
nor U23543 (N_23543,N_21058,N_20621);
nand U23544 (N_23544,N_21649,N_21611);
nand U23545 (N_23545,N_22369,N_22291);
nor U23546 (N_23546,N_21887,N_20901);
nand U23547 (N_23547,N_21639,N_21751);
and U23548 (N_23548,N_21358,N_21614);
and U23549 (N_23549,N_20624,N_21057);
xor U23550 (N_23550,N_22225,N_22000);
nand U23551 (N_23551,N_20242,N_22421);
xnor U23552 (N_23552,N_20725,N_22216);
nand U23553 (N_23553,N_22437,N_22273);
nand U23554 (N_23554,N_20716,N_22351);
or U23555 (N_23555,N_20806,N_22319);
nand U23556 (N_23556,N_21147,N_20190);
and U23557 (N_23557,N_20453,N_21240);
and U23558 (N_23558,N_21134,N_20638);
or U23559 (N_23559,N_21945,N_22059);
nand U23560 (N_23560,N_21236,N_20579);
nor U23561 (N_23561,N_22436,N_21067);
nor U23562 (N_23562,N_22100,N_22303);
xor U23563 (N_23563,N_20414,N_20063);
and U23564 (N_23564,N_20443,N_20395);
nand U23565 (N_23565,N_20888,N_20707);
and U23566 (N_23566,N_20735,N_20786);
and U23567 (N_23567,N_20484,N_22155);
or U23568 (N_23568,N_21997,N_22127);
nand U23569 (N_23569,N_20590,N_22366);
or U23570 (N_23570,N_22176,N_22481);
nor U23571 (N_23571,N_20666,N_20234);
and U23572 (N_23572,N_22334,N_20965);
and U23573 (N_23573,N_21097,N_21646);
xor U23574 (N_23574,N_22482,N_21497);
nor U23575 (N_23575,N_21220,N_22249);
nor U23576 (N_23576,N_22233,N_22486);
or U23577 (N_23577,N_20528,N_22304);
or U23578 (N_23578,N_20384,N_20859);
nor U23579 (N_23579,N_22121,N_20551);
or U23580 (N_23580,N_20121,N_21176);
or U23581 (N_23581,N_22036,N_22295);
nand U23582 (N_23582,N_21930,N_21181);
nor U23583 (N_23583,N_21803,N_20485);
nand U23584 (N_23584,N_20144,N_21526);
xor U23585 (N_23585,N_22408,N_22444);
or U23586 (N_23586,N_21700,N_20174);
and U23587 (N_23587,N_21562,N_20933);
or U23588 (N_23588,N_20381,N_21875);
or U23589 (N_23589,N_21007,N_21689);
xor U23590 (N_23590,N_21718,N_22480);
and U23591 (N_23591,N_21568,N_21684);
or U23592 (N_23592,N_20405,N_22257);
nand U23593 (N_23593,N_20462,N_22460);
or U23594 (N_23594,N_20822,N_21247);
nand U23595 (N_23595,N_22108,N_20274);
nand U23596 (N_23596,N_20686,N_22156);
and U23597 (N_23597,N_21317,N_20115);
nand U23598 (N_23598,N_21216,N_20275);
nand U23599 (N_23599,N_20664,N_21230);
nand U23600 (N_23600,N_20780,N_21564);
xor U23601 (N_23601,N_20839,N_20171);
or U23602 (N_23602,N_20399,N_20588);
and U23603 (N_23603,N_22025,N_22329);
nor U23604 (N_23604,N_21900,N_20813);
or U23605 (N_23605,N_20493,N_22388);
xnor U23606 (N_23606,N_21376,N_22094);
xor U23607 (N_23607,N_21990,N_21016);
nor U23608 (N_23608,N_20961,N_20838);
nor U23609 (N_23609,N_22123,N_20146);
or U23610 (N_23610,N_21902,N_20871);
and U23611 (N_23611,N_21706,N_21880);
or U23612 (N_23612,N_22201,N_21661);
and U23613 (N_23613,N_20229,N_21563);
nor U23614 (N_23614,N_20265,N_21027);
nand U23615 (N_23615,N_20191,N_20082);
or U23616 (N_23616,N_20749,N_21348);
nor U23617 (N_23617,N_20427,N_20486);
and U23618 (N_23618,N_20985,N_21788);
nand U23619 (N_23619,N_20262,N_21872);
nor U23620 (N_23620,N_20013,N_20948);
nand U23621 (N_23621,N_20386,N_22336);
nor U23622 (N_23622,N_20978,N_20468);
or U23623 (N_23623,N_20325,N_21002);
or U23624 (N_23624,N_21513,N_20984);
nand U23625 (N_23625,N_22462,N_21848);
xnor U23626 (N_23626,N_20421,N_20261);
and U23627 (N_23627,N_22014,N_20968);
and U23628 (N_23628,N_22425,N_22258);
nand U23629 (N_23629,N_21637,N_22439);
and U23630 (N_23630,N_21290,N_22052);
xor U23631 (N_23631,N_21229,N_20724);
nand U23632 (N_23632,N_21940,N_21781);
nor U23633 (N_23633,N_21219,N_22310);
nor U23634 (N_23634,N_21507,N_20372);
or U23635 (N_23635,N_21009,N_21101);
xor U23636 (N_23636,N_20902,N_20586);
xnor U23637 (N_23637,N_20177,N_20993);
and U23638 (N_23638,N_21840,N_20601);
or U23639 (N_23639,N_21424,N_20417);
xor U23640 (N_23640,N_21145,N_20491);
nand U23641 (N_23641,N_22058,N_21398);
or U23642 (N_23642,N_21414,N_21603);
nor U23643 (N_23643,N_21801,N_21320);
nand U23644 (N_23644,N_21601,N_21237);
and U23645 (N_23645,N_22326,N_21033);
xor U23646 (N_23646,N_22344,N_21510);
and U23647 (N_23647,N_20025,N_20761);
or U23648 (N_23648,N_20884,N_20542);
or U23649 (N_23649,N_20197,N_22318);
xor U23650 (N_23650,N_22400,N_20876);
nor U23651 (N_23651,N_20431,N_21272);
xnor U23652 (N_23652,N_20112,N_20711);
or U23653 (N_23653,N_21977,N_20328);
nand U23654 (N_23654,N_20419,N_20674);
and U23655 (N_23655,N_20334,N_21459);
nand U23656 (N_23656,N_21874,N_22107);
or U23657 (N_23657,N_22312,N_20924);
xnor U23658 (N_23658,N_21391,N_21356);
xor U23659 (N_23659,N_22229,N_20031);
nor U23660 (N_23660,N_21248,N_21411);
nand U23661 (N_23661,N_21910,N_21680);
nor U23662 (N_23662,N_21188,N_20065);
nand U23663 (N_23663,N_21567,N_20513);
and U23664 (N_23664,N_20202,N_20503);
nor U23665 (N_23665,N_20731,N_20840);
nand U23666 (N_23666,N_20003,N_21560);
and U23667 (N_23667,N_20104,N_22354);
xnor U23668 (N_23668,N_20921,N_20272);
xnor U23669 (N_23669,N_22247,N_21784);
or U23670 (N_23670,N_21962,N_22116);
nand U23671 (N_23671,N_22301,N_20423);
xnor U23672 (N_23672,N_21516,N_22358);
nand U23673 (N_23673,N_20495,N_21969);
and U23674 (N_23674,N_21577,N_21767);
xor U23675 (N_23675,N_21976,N_21363);
or U23676 (N_23676,N_21435,N_20540);
and U23677 (N_23677,N_21600,N_21074);
nand U23678 (N_23678,N_21421,N_21823);
xnor U23679 (N_23679,N_20239,N_21019);
and U23680 (N_23680,N_21111,N_20388);
or U23681 (N_23681,N_21170,N_21437);
nand U23682 (N_23682,N_21452,N_20167);
xnor U23683 (N_23683,N_22035,N_21315);
and U23684 (N_23684,N_20193,N_22432);
xor U23685 (N_23685,N_21549,N_20282);
nor U23686 (N_23686,N_21954,N_21561);
xor U23687 (N_23687,N_20927,N_21550);
xor U23688 (N_23688,N_21898,N_20311);
nor U23689 (N_23689,N_20508,N_20653);
nand U23690 (N_23690,N_21443,N_20285);
nor U23691 (N_23691,N_20847,N_21260);
nor U23692 (N_23692,N_21362,N_20070);
nand U23693 (N_23693,N_20375,N_22401);
nand U23694 (N_23694,N_21108,N_21020);
and U23695 (N_23695,N_21733,N_21897);
and U23696 (N_23696,N_21405,N_20437);
or U23697 (N_23697,N_21503,N_20816);
and U23698 (N_23698,N_20320,N_20083);
and U23699 (N_23699,N_20270,N_21888);
xnor U23700 (N_23700,N_20582,N_22131);
or U23701 (N_23701,N_20252,N_21267);
and U23702 (N_23702,N_20777,N_21223);
nand U23703 (N_23703,N_20913,N_21690);
nand U23704 (N_23704,N_20730,N_20630);
and U23705 (N_23705,N_20478,N_21958);
or U23706 (N_23706,N_20233,N_21852);
and U23707 (N_23707,N_21092,N_21882);
and U23708 (N_23708,N_20793,N_22447);
xnor U23709 (N_23709,N_21667,N_22451);
nor U23710 (N_23710,N_21748,N_21685);
or U23711 (N_23711,N_21658,N_20867);
nor U23712 (N_23712,N_22497,N_20680);
or U23713 (N_23713,N_21769,N_20278);
nor U23714 (N_23714,N_21112,N_20092);
xor U23715 (N_23715,N_20249,N_22260);
nor U23716 (N_23716,N_21177,N_20276);
and U23717 (N_23717,N_20862,N_21918);
xor U23718 (N_23718,N_21431,N_20264);
xor U23719 (N_23719,N_21015,N_21386);
and U23720 (N_23720,N_22271,N_22259);
nand U23721 (N_23721,N_20728,N_20080);
or U23722 (N_23722,N_20119,N_21268);
xnor U23723 (N_23723,N_22280,N_20472);
xor U23724 (N_23724,N_20049,N_20226);
xor U23725 (N_23725,N_21798,N_20905);
or U23726 (N_23726,N_22335,N_21069);
or U23727 (N_23727,N_20991,N_21257);
or U23728 (N_23728,N_21617,N_20907);
and U23729 (N_23729,N_20365,N_20085);
xnor U23730 (N_23730,N_20947,N_22117);
and U23731 (N_23731,N_21161,N_21933);
xor U23732 (N_23732,N_21530,N_20939);
or U23733 (N_23733,N_22380,N_21124);
and U23734 (N_23734,N_21288,N_22440);
nor U23735 (N_23735,N_22163,N_20812);
nand U23736 (N_23736,N_20804,N_20853);
nand U23737 (N_23737,N_20449,N_20301);
xnor U23738 (N_23738,N_22228,N_20500);
xnor U23739 (N_23739,N_20942,N_21891);
nor U23740 (N_23740,N_21988,N_21694);
and U23741 (N_23741,N_20946,N_20412);
or U23742 (N_23742,N_20176,N_22164);
xnor U23743 (N_23743,N_21306,N_21084);
or U23744 (N_23744,N_20439,N_22256);
nor U23745 (N_23745,N_20352,N_20596);
nand U23746 (N_23746,N_20251,N_21173);
xor U23747 (N_23747,N_22111,N_20855);
nand U23748 (N_23748,N_21592,N_20505);
xnor U23749 (N_23749,N_21565,N_21772);
nor U23750 (N_23750,N_20807,N_20597);
nor U23751 (N_23751,N_20027,N_20847);
nand U23752 (N_23752,N_21781,N_20789);
xor U23753 (N_23753,N_20189,N_20837);
nor U23754 (N_23754,N_20524,N_20590);
or U23755 (N_23755,N_21752,N_21619);
nand U23756 (N_23756,N_22253,N_20720);
or U23757 (N_23757,N_22395,N_22051);
nand U23758 (N_23758,N_22102,N_22362);
xnor U23759 (N_23759,N_20822,N_21314);
nand U23760 (N_23760,N_20839,N_20524);
and U23761 (N_23761,N_21787,N_22370);
nor U23762 (N_23762,N_22380,N_21518);
nor U23763 (N_23763,N_22006,N_20795);
nor U23764 (N_23764,N_21247,N_20856);
or U23765 (N_23765,N_21937,N_21852);
nor U23766 (N_23766,N_21782,N_20540);
and U23767 (N_23767,N_20598,N_20677);
nand U23768 (N_23768,N_20919,N_22357);
nor U23769 (N_23769,N_20412,N_20702);
or U23770 (N_23770,N_20343,N_21934);
nor U23771 (N_23771,N_20350,N_21912);
nand U23772 (N_23772,N_22208,N_21308);
xor U23773 (N_23773,N_21340,N_21211);
or U23774 (N_23774,N_21405,N_20627);
nor U23775 (N_23775,N_22472,N_22232);
or U23776 (N_23776,N_21892,N_21272);
nand U23777 (N_23777,N_21614,N_20707);
and U23778 (N_23778,N_21513,N_20800);
xnor U23779 (N_23779,N_21354,N_21137);
nand U23780 (N_23780,N_20251,N_22441);
nor U23781 (N_23781,N_20456,N_20374);
or U23782 (N_23782,N_21270,N_22024);
nor U23783 (N_23783,N_21196,N_21950);
nand U23784 (N_23784,N_20132,N_21156);
and U23785 (N_23785,N_20253,N_20182);
xor U23786 (N_23786,N_21948,N_21110);
or U23787 (N_23787,N_20258,N_20452);
or U23788 (N_23788,N_21551,N_21984);
nor U23789 (N_23789,N_20495,N_22441);
or U23790 (N_23790,N_21197,N_20420);
and U23791 (N_23791,N_21569,N_21965);
nor U23792 (N_23792,N_21318,N_22059);
nor U23793 (N_23793,N_20164,N_20458);
nor U23794 (N_23794,N_21518,N_20366);
nor U23795 (N_23795,N_22209,N_22282);
xor U23796 (N_23796,N_20731,N_21072);
nor U23797 (N_23797,N_21773,N_21831);
and U23798 (N_23798,N_20826,N_20918);
nand U23799 (N_23799,N_20984,N_20122);
nor U23800 (N_23800,N_20224,N_21140);
xor U23801 (N_23801,N_22133,N_21487);
xor U23802 (N_23802,N_20257,N_22459);
nor U23803 (N_23803,N_21880,N_20756);
or U23804 (N_23804,N_20763,N_21118);
nor U23805 (N_23805,N_21928,N_21193);
nand U23806 (N_23806,N_21999,N_21301);
nor U23807 (N_23807,N_21714,N_21883);
xor U23808 (N_23808,N_22313,N_22132);
nand U23809 (N_23809,N_20204,N_21574);
and U23810 (N_23810,N_20003,N_21824);
xnor U23811 (N_23811,N_21523,N_21524);
nand U23812 (N_23812,N_20998,N_21789);
and U23813 (N_23813,N_20672,N_20720);
xnor U23814 (N_23814,N_20172,N_20580);
and U23815 (N_23815,N_20737,N_20373);
nor U23816 (N_23816,N_21167,N_21521);
nand U23817 (N_23817,N_20521,N_20049);
nand U23818 (N_23818,N_21787,N_20233);
or U23819 (N_23819,N_21080,N_21237);
nand U23820 (N_23820,N_21945,N_20152);
or U23821 (N_23821,N_20259,N_22325);
xor U23822 (N_23822,N_20654,N_22420);
nor U23823 (N_23823,N_20651,N_20893);
nand U23824 (N_23824,N_21367,N_21897);
and U23825 (N_23825,N_21186,N_21520);
xor U23826 (N_23826,N_21610,N_20108);
nand U23827 (N_23827,N_20264,N_21140);
nand U23828 (N_23828,N_21546,N_21830);
nor U23829 (N_23829,N_21719,N_20127);
nand U23830 (N_23830,N_21881,N_20753);
nor U23831 (N_23831,N_20100,N_20460);
nand U23832 (N_23832,N_22025,N_20860);
xnor U23833 (N_23833,N_21372,N_20999);
nor U23834 (N_23834,N_22152,N_21729);
or U23835 (N_23835,N_20672,N_20024);
nor U23836 (N_23836,N_21390,N_20985);
xnor U23837 (N_23837,N_22268,N_22381);
or U23838 (N_23838,N_21338,N_20721);
nand U23839 (N_23839,N_20554,N_21282);
and U23840 (N_23840,N_20704,N_20807);
xnor U23841 (N_23841,N_20247,N_22201);
nor U23842 (N_23842,N_21411,N_20358);
xnor U23843 (N_23843,N_21433,N_20106);
nor U23844 (N_23844,N_21066,N_20738);
xnor U23845 (N_23845,N_21956,N_20415);
xnor U23846 (N_23846,N_20450,N_22177);
nand U23847 (N_23847,N_21987,N_22195);
nor U23848 (N_23848,N_21397,N_21150);
nor U23849 (N_23849,N_20072,N_22483);
xor U23850 (N_23850,N_21575,N_21294);
and U23851 (N_23851,N_20178,N_21662);
nor U23852 (N_23852,N_22158,N_22093);
xor U23853 (N_23853,N_22438,N_21909);
nor U23854 (N_23854,N_21248,N_22154);
xor U23855 (N_23855,N_22326,N_22090);
nor U23856 (N_23856,N_20830,N_21917);
or U23857 (N_23857,N_22121,N_22028);
nor U23858 (N_23858,N_20432,N_22217);
nand U23859 (N_23859,N_20222,N_22160);
or U23860 (N_23860,N_22180,N_21009);
nand U23861 (N_23861,N_22104,N_21252);
or U23862 (N_23862,N_21902,N_21625);
nor U23863 (N_23863,N_21735,N_22105);
or U23864 (N_23864,N_22472,N_20887);
nor U23865 (N_23865,N_21034,N_22418);
nand U23866 (N_23866,N_22294,N_20258);
or U23867 (N_23867,N_22357,N_20875);
and U23868 (N_23868,N_21322,N_22313);
nand U23869 (N_23869,N_20086,N_22240);
nor U23870 (N_23870,N_21503,N_21321);
nor U23871 (N_23871,N_22409,N_20765);
xnor U23872 (N_23872,N_21505,N_21670);
nor U23873 (N_23873,N_22487,N_20460);
nand U23874 (N_23874,N_21500,N_20449);
and U23875 (N_23875,N_21951,N_20257);
or U23876 (N_23876,N_20927,N_21749);
and U23877 (N_23877,N_21816,N_21018);
nor U23878 (N_23878,N_20768,N_20324);
or U23879 (N_23879,N_21266,N_20233);
nor U23880 (N_23880,N_22472,N_21947);
and U23881 (N_23881,N_21087,N_20922);
xor U23882 (N_23882,N_20200,N_20637);
nand U23883 (N_23883,N_21046,N_20702);
nor U23884 (N_23884,N_22305,N_20901);
nor U23885 (N_23885,N_21990,N_21867);
xnor U23886 (N_23886,N_22180,N_21972);
and U23887 (N_23887,N_21667,N_21191);
nor U23888 (N_23888,N_22294,N_21816);
or U23889 (N_23889,N_20106,N_21612);
nor U23890 (N_23890,N_22006,N_21461);
xor U23891 (N_23891,N_21800,N_20034);
or U23892 (N_23892,N_21282,N_20695);
xor U23893 (N_23893,N_21390,N_22312);
nor U23894 (N_23894,N_22224,N_21351);
nand U23895 (N_23895,N_20938,N_21786);
xnor U23896 (N_23896,N_21544,N_20079);
and U23897 (N_23897,N_20396,N_20549);
xnor U23898 (N_23898,N_22279,N_22047);
xor U23899 (N_23899,N_21921,N_22126);
and U23900 (N_23900,N_20801,N_21065);
xor U23901 (N_23901,N_21242,N_20597);
xnor U23902 (N_23902,N_21398,N_20257);
xnor U23903 (N_23903,N_21682,N_21499);
and U23904 (N_23904,N_20630,N_21639);
nor U23905 (N_23905,N_22025,N_20369);
xor U23906 (N_23906,N_20202,N_22095);
nor U23907 (N_23907,N_21687,N_22316);
xor U23908 (N_23908,N_22054,N_22123);
or U23909 (N_23909,N_21549,N_20796);
or U23910 (N_23910,N_20734,N_22291);
xor U23911 (N_23911,N_22372,N_20134);
nor U23912 (N_23912,N_20890,N_21813);
nor U23913 (N_23913,N_21553,N_20281);
xor U23914 (N_23914,N_21438,N_22085);
or U23915 (N_23915,N_21113,N_20807);
xor U23916 (N_23916,N_21366,N_21573);
or U23917 (N_23917,N_20699,N_20050);
nand U23918 (N_23918,N_22233,N_20561);
nand U23919 (N_23919,N_20685,N_20507);
and U23920 (N_23920,N_21095,N_21468);
xor U23921 (N_23921,N_22225,N_20582);
or U23922 (N_23922,N_20169,N_21548);
xor U23923 (N_23923,N_21356,N_21115);
nand U23924 (N_23924,N_21991,N_22277);
nor U23925 (N_23925,N_20963,N_20204);
and U23926 (N_23926,N_20504,N_20290);
and U23927 (N_23927,N_22400,N_22464);
nand U23928 (N_23928,N_20133,N_20153);
xnor U23929 (N_23929,N_21452,N_21487);
nand U23930 (N_23930,N_21660,N_20226);
xor U23931 (N_23931,N_21065,N_22120);
xor U23932 (N_23932,N_21580,N_21501);
or U23933 (N_23933,N_22135,N_20997);
nor U23934 (N_23934,N_20428,N_20769);
xnor U23935 (N_23935,N_20671,N_21950);
xor U23936 (N_23936,N_20079,N_21133);
nor U23937 (N_23937,N_22301,N_21199);
or U23938 (N_23938,N_20483,N_21069);
and U23939 (N_23939,N_20268,N_22461);
or U23940 (N_23940,N_20383,N_20995);
or U23941 (N_23941,N_20938,N_22022);
nor U23942 (N_23942,N_20337,N_20702);
nand U23943 (N_23943,N_20779,N_20805);
nand U23944 (N_23944,N_20579,N_20102);
and U23945 (N_23945,N_20479,N_20817);
nand U23946 (N_23946,N_21836,N_21204);
xor U23947 (N_23947,N_21333,N_22032);
and U23948 (N_23948,N_22190,N_21623);
xor U23949 (N_23949,N_22439,N_20458);
xnor U23950 (N_23950,N_21319,N_20732);
and U23951 (N_23951,N_21704,N_20955);
xor U23952 (N_23952,N_21092,N_20483);
or U23953 (N_23953,N_21498,N_21779);
and U23954 (N_23954,N_21292,N_22489);
nor U23955 (N_23955,N_20212,N_22430);
and U23956 (N_23956,N_20053,N_20110);
and U23957 (N_23957,N_20794,N_21920);
nor U23958 (N_23958,N_20364,N_20842);
nor U23959 (N_23959,N_21505,N_22005);
nand U23960 (N_23960,N_21285,N_20879);
nand U23961 (N_23961,N_20858,N_21766);
and U23962 (N_23962,N_20694,N_21646);
xnor U23963 (N_23963,N_20627,N_21890);
nand U23964 (N_23964,N_20596,N_21433);
nand U23965 (N_23965,N_22473,N_20475);
xor U23966 (N_23966,N_21143,N_20155);
xnor U23967 (N_23967,N_21116,N_22179);
xnor U23968 (N_23968,N_20027,N_21997);
xnor U23969 (N_23969,N_21938,N_21901);
xnor U23970 (N_23970,N_21836,N_21807);
or U23971 (N_23971,N_22255,N_20898);
nor U23972 (N_23972,N_22357,N_20934);
nor U23973 (N_23973,N_22256,N_20522);
nand U23974 (N_23974,N_20972,N_21223);
nor U23975 (N_23975,N_21075,N_21527);
or U23976 (N_23976,N_21411,N_20605);
and U23977 (N_23977,N_20720,N_21419);
nor U23978 (N_23978,N_22467,N_20884);
xnor U23979 (N_23979,N_21304,N_20418);
or U23980 (N_23980,N_20901,N_22291);
and U23981 (N_23981,N_20472,N_21387);
and U23982 (N_23982,N_20389,N_21442);
xnor U23983 (N_23983,N_22172,N_22173);
xnor U23984 (N_23984,N_22004,N_21894);
or U23985 (N_23985,N_20847,N_20913);
nor U23986 (N_23986,N_21004,N_22032);
or U23987 (N_23987,N_21270,N_21561);
or U23988 (N_23988,N_20072,N_20294);
nand U23989 (N_23989,N_21901,N_20859);
xnor U23990 (N_23990,N_20582,N_22209);
and U23991 (N_23991,N_21157,N_20992);
nor U23992 (N_23992,N_20100,N_21407);
or U23993 (N_23993,N_20231,N_20538);
or U23994 (N_23994,N_21254,N_20050);
or U23995 (N_23995,N_22184,N_21587);
or U23996 (N_23996,N_21315,N_20791);
xor U23997 (N_23997,N_21377,N_20530);
or U23998 (N_23998,N_20865,N_20254);
and U23999 (N_23999,N_20567,N_21966);
nor U24000 (N_24000,N_20025,N_21434);
nor U24001 (N_24001,N_22249,N_21562);
xnor U24002 (N_24002,N_20397,N_20561);
xor U24003 (N_24003,N_20922,N_21739);
or U24004 (N_24004,N_22136,N_22122);
and U24005 (N_24005,N_20971,N_21430);
nand U24006 (N_24006,N_21049,N_21740);
nand U24007 (N_24007,N_20695,N_22077);
or U24008 (N_24008,N_20996,N_20909);
nor U24009 (N_24009,N_22143,N_20819);
or U24010 (N_24010,N_20617,N_21946);
nand U24011 (N_24011,N_22037,N_21373);
xor U24012 (N_24012,N_20623,N_21477);
nor U24013 (N_24013,N_21488,N_21403);
nor U24014 (N_24014,N_21625,N_20383);
or U24015 (N_24015,N_22130,N_21785);
or U24016 (N_24016,N_22471,N_20428);
nor U24017 (N_24017,N_21243,N_21087);
xor U24018 (N_24018,N_20210,N_21899);
nand U24019 (N_24019,N_21189,N_21705);
and U24020 (N_24020,N_21886,N_20769);
nand U24021 (N_24021,N_22364,N_22210);
and U24022 (N_24022,N_21867,N_20554);
nand U24023 (N_24023,N_20797,N_21108);
nor U24024 (N_24024,N_21976,N_21734);
nor U24025 (N_24025,N_21895,N_20580);
and U24026 (N_24026,N_20978,N_20680);
and U24027 (N_24027,N_21605,N_20856);
nand U24028 (N_24028,N_20288,N_22470);
nand U24029 (N_24029,N_22092,N_21681);
xor U24030 (N_24030,N_20882,N_22083);
and U24031 (N_24031,N_22277,N_20256);
nor U24032 (N_24032,N_20464,N_22316);
nor U24033 (N_24033,N_22112,N_21588);
and U24034 (N_24034,N_21529,N_20419);
nand U24035 (N_24035,N_21232,N_21133);
nand U24036 (N_24036,N_20607,N_21115);
or U24037 (N_24037,N_21843,N_20764);
nand U24038 (N_24038,N_21930,N_21904);
or U24039 (N_24039,N_20632,N_21242);
nand U24040 (N_24040,N_20122,N_20346);
nand U24041 (N_24041,N_21823,N_21334);
nor U24042 (N_24042,N_21272,N_21945);
nor U24043 (N_24043,N_21838,N_20575);
nand U24044 (N_24044,N_20708,N_20139);
xnor U24045 (N_24045,N_21370,N_21935);
or U24046 (N_24046,N_22441,N_22435);
or U24047 (N_24047,N_21009,N_20649);
xor U24048 (N_24048,N_21639,N_20960);
nand U24049 (N_24049,N_22154,N_20450);
and U24050 (N_24050,N_21885,N_20045);
nor U24051 (N_24051,N_22299,N_20774);
xnor U24052 (N_24052,N_21577,N_20157);
nor U24053 (N_24053,N_20491,N_22060);
or U24054 (N_24054,N_21304,N_20745);
and U24055 (N_24055,N_22286,N_20072);
nor U24056 (N_24056,N_20747,N_21534);
nand U24057 (N_24057,N_21121,N_20739);
nand U24058 (N_24058,N_20022,N_20794);
xor U24059 (N_24059,N_20175,N_21470);
nor U24060 (N_24060,N_21248,N_20105);
xor U24061 (N_24061,N_20794,N_21559);
xor U24062 (N_24062,N_22195,N_21885);
xnor U24063 (N_24063,N_21234,N_20135);
nand U24064 (N_24064,N_20534,N_21756);
or U24065 (N_24065,N_22159,N_22320);
nor U24066 (N_24066,N_21007,N_21717);
or U24067 (N_24067,N_20483,N_21521);
or U24068 (N_24068,N_20365,N_21786);
or U24069 (N_24069,N_22153,N_21663);
nand U24070 (N_24070,N_22442,N_22374);
or U24071 (N_24071,N_21546,N_20369);
and U24072 (N_24072,N_21498,N_21094);
and U24073 (N_24073,N_21103,N_20265);
nor U24074 (N_24074,N_20793,N_21035);
and U24075 (N_24075,N_21650,N_20380);
xnor U24076 (N_24076,N_22233,N_20667);
and U24077 (N_24077,N_20293,N_21067);
or U24078 (N_24078,N_20819,N_20085);
and U24079 (N_24079,N_20754,N_20507);
nor U24080 (N_24080,N_21149,N_20474);
nand U24081 (N_24081,N_22049,N_20902);
nor U24082 (N_24082,N_20234,N_20107);
xor U24083 (N_24083,N_21684,N_21552);
nor U24084 (N_24084,N_21011,N_22084);
nand U24085 (N_24085,N_20692,N_21167);
xnor U24086 (N_24086,N_20394,N_21532);
nor U24087 (N_24087,N_22203,N_21961);
xnor U24088 (N_24088,N_20014,N_21307);
nor U24089 (N_24089,N_20988,N_20633);
and U24090 (N_24090,N_21891,N_22097);
and U24091 (N_24091,N_21640,N_21685);
nand U24092 (N_24092,N_22329,N_22119);
or U24093 (N_24093,N_21031,N_21609);
or U24094 (N_24094,N_20480,N_21093);
or U24095 (N_24095,N_22031,N_20040);
and U24096 (N_24096,N_20274,N_21047);
nand U24097 (N_24097,N_21611,N_21001);
or U24098 (N_24098,N_21081,N_20954);
nand U24099 (N_24099,N_20438,N_20078);
nor U24100 (N_24100,N_21312,N_21745);
or U24101 (N_24101,N_21051,N_20520);
nor U24102 (N_24102,N_20871,N_21526);
nand U24103 (N_24103,N_22194,N_22307);
xnor U24104 (N_24104,N_21056,N_22317);
and U24105 (N_24105,N_20385,N_20480);
xnor U24106 (N_24106,N_21936,N_21876);
nand U24107 (N_24107,N_20952,N_20327);
xor U24108 (N_24108,N_20523,N_20978);
nor U24109 (N_24109,N_20669,N_21622);
nand U24110 (N_24110,N_21970,N_21148);
and U24111 (N_24111,N_21429,N_20060);
nor U24112 (N_24112,N_22495,N_21466);
or U24113 (N_24113,N_21331,N_22251);
nand U24114 (N_24114,N_20854,N_22428);
xnor U24115 (N_24115,N_20979,N_20200);
or U24116 (N_24116,N_22321,N_20210);
nand U24117 (N_24117,N_20231,N_21590);
and U24118 (N_24118,N_21830,N_21331);
nand U24119 (N_24119,N_20004,N_21787);
or U24120 (N_24120,N_20537,N_22052);
nor U24121 (N_24121,N_20231,N_22436);
or U24122 (N_24122,N_21732,N_20090);
xor U24123 (N_24123,N_22388,N_21174);
nor U24124 (N_24124,N_20531,N_20017);
and U24125 (N_24125,N_20013,N_21374);
or U24126 (N_24126,N_21582,N_21569);
or U24127 (N_24127,N_21716,N_20723);
nor U24128 (N_24128,N_20209,N_21781);
nor U24129 (N_24129,N_20176,N_22055);
or U24130 (N_24130,N_22433,N_20052);
nor U24131 (N_24131,N_22057,N_22047);
and U24132 (N_24132,N_22163,N_20783);
and U24133 (N_24133,N_20082,N_20236);
and U24134 (N_24134,N_21757,N_21977);
or U24135 (N_24135,N_22330,N_21376);
xor U24136 (N_24136,N_22466,N_20087);
and U24137 (N_24137,N_20416,N_22161);
nor U24138 (N_24138,N_21996,N_20008);
xnor U24139 (N_24139,N_20531,N_22264);
and U24140 (N_24140,N_20898,N_20386);
and U24141 (N_24141,N_20059,N_22189);
xnor U24142 (N_24142,N_21603,N_20913);
and U24143 (N_24143,N_21975,N_22416);
xor U24144 (N_24144,N_21842,N_20453);
and U24145 (N_24145,N_21639,N_21618);
nand U24146 (N_24146,N_21840,N_20865);
nand U24147 (N_24147,N_20817,N_20720);
nand U24148 (N_24148,N_21400,N_20440);
or U24149 (N_24149,N_21699,N_20734);
xnor U24150 (N_24150,N_21333,N_21077);
nor U24151 (N_24151,N_21662,N_21818);
or U24152 (N_24152,N_20321,N_21406);
nand U24153 (N_24153,N_20684,N_21705);
nand U24154 (N_24154,N_20153,N_21514);
nor U24155 (N_24155,N_22329,N_21042);
nand U24156 (N_24156,N_21535,N_21670);
xnor U24157 (N_24157,N_20812,N_20076);
and U24158 (N_24158,N_21338,N_20852);
xor U24159 (N_24159,N_20570,N_22004);
xor U24160 (N_24160,N_21293,N_22090);
nor U24161 (N_24161,N_22363,N_20639);
and U24162 (N_24162,N_21994,N_22267);
nand U24163 (N_24163,N_20355,N_21173);
or U24164 (N_24164,N_20700,N_22295);
and U24165 (N_24165,N_22211,N_20594);
xnor U24166 (N_24166,N_22495,N_20774);
and U24167 (N_24167,N_21345,N_21237);
nor U24168 (N_24168,N_22153,N_20130);
and U24169 (N_24169,N_20038,N_21043);
and U24170 (N_24170,N_21576,N_20710);
nand U24171 (N_24171,N_20123,N_21232);
nor U24172 (N_24172,N_21183,N_20201);
nand U24173 (N_24173,N_21698,N_20477);
xor U24174 (N_24174,N_21316,N_22098);
nand U24175 (N_24175,N_21117,N_21745);
nor U24176 (N_24176,N_22194,N_21915);
nor U24177 (N_24177,N_21577,N_20210);
nor U24178 (N_24178,N_20674,N_20101);
nor U24179 (N_24179,N_20986,N_21854);
nor U24180 (N_24180,N_22252,N_22296);
nor U24181 (N_24181,N_21347,N_20950);
xnor U24182 (N_24182,N_20929,N_21356);
xnor U24183 (N_24183,N_20062,N_22040);
xor U24184 (N_24184,N_20247,N_21734);
or U24185 (N_24185,N_21473,N_21480);
nand U24186 (N_24186,N_21817,N_20546);
and U24187 (N_24187,N_21854,N_21688);
or U24188 (N_24188,N_21039,N_20718);
or U24189 (N_24189,N_22126,N_20094);
or U24190 (N_24190,N_21561,N_20426);
nand U24191 (N_24191,N_21142,N_22404);
nor U24192 (N_24192,N_20960,N_20956);
and U24193 (N_24193,N_21456,N_21735);
nand U24194 (N_24194,N_20967,N_21516);
nand U24195 (N_24195,N_21369,N_21273);
and U24196 (N_24196,N_21760,N_20866);
or U24197 (N_24197,N_22051,N_21860);
and U24198 (N_24198,N_21210,N_22043);
nand U24199 (N_24199,N_21252,N_21439);
nor U24200 (N_24200,N_21040,N_21358);
nand U24201 (N_24201,N_20938,N_22260);
or U24202 (N_24202,N_20971,N_20544);
or U24203 (N_24203,N_20457,N_22171);
nor U24204 (N_24204,N_21320,N_22005);
or U24205 (N_24205,N_21198,N_22433);
nand U24206 (N_24206,N_22026,N_20121);
xnor U24207 (N_24207,N_20477,N_21369);
nor U24208 (N_24208,N_22253,N_21170);
or U24209 (N_24209,N_20627,N_20596);
nand U24210 (N_24210,N_21211,N_21299);
nand U24211 (N_24211,N_20267,N_20016);
nand U24212 (N_24212,N_20389,N_20598);
or U24213 (N_24213,N_22100,N_21886);
and U24214 (N_24214,N_22066,N_21023);
nand U24215 (N_24215,N_20889,N_21377);
and U24216 (N_24216,N_20837,N_21017);
or U24217 (N_24217,N_20665,N_22247);
nor U24218 (N_24218,N_22109,N_20355);
nor U24219 (N_24219,N_22145,N_20604);
xnor U24220 (N_24220,N_21341,N_20757);
nor U24221 (N_24221,N_22021,N_21973);
nor U24222 (N_24222,N_20938,N_21592);
nor U24223 (N_24223,N_20039,N_21409);
or U24224 (N_24224,N_21889,N_20192);
and U24225 (N_24225,N_21788,N_20174);
xor U24226 (N_24226,N_21132,N_20317);
or U24227 (N_24227,N_21181,N_21464);
xnor U24228 (N_24228,N_21307,N_20021);
or U24229 (N_24229,N_22301,N_21703);
nand U24230 (N_24230,N_20892,N_22361);
or U24231 (N_24231,N_21505,N_20838);
nor U24232 (N_24232,N_21577,N_20516);
nor U24233 (N_24233,N_20230,N_20283);
and U24234 (N_24234,N_20396,N_20558);
and U24235 (N_24235,N_20888,N_20213);
xor U24236 (N_24236,N_22439,N_22149);
nor U24237 (N_24237,N_21108,N_20261);
or U24238 (N_24238,N_21943,N_20414);
and U24239 (N_24239,N_21040,N_20734);
nor U24240 (N_24240,N_22075,N_20734);
and U24241 (N_24241,N_21641,N_21331);
nor U24242 (N_24242,N_21587,N_21204);
and U24243 (N_24243,N_21070,N_20995);
and U24244 (N_24244,N_21855,N_21880);
xor U24245 (N_24245,N_21362,N_20724);
nor U24246 (N_24246,N_22342,N_21467);
and U24247 (N_24247,N_21463,N_20570);
nor U24248 (N_24248,N_21874,N_20998);
and U24249 (N_24249,N_21412,N_21275);
nand U24250 (N_24250,N_20889,N_21004);
xor U24251 (N_24251,N_21122,N_20345);
nand U24252 (N_24252,N_22334,N_20024);
or U24253 (N_24253,N_21158,N_21297);
and U24254 (N_24254,N_20729,N_22048);
nor U24255 (N_24255,N_21661,N_20770);
nor U24256 (N_24256,N_21934,N_22141);
and U24257 (N_24257,N_21501,N_21363);
nand U24258 (N_24258,N_21809,N_21882);
nor U24259 (N_24259,N_21164,N_21641);
and U24260 (N_24260,N_21796,N_20885);
or U24261 (N_24261,N_22472,N_20053);
or U24262 (N_24262,N_20840,N_20054);
nand U24263 (N_24263,N_21286,N_21452);
xor U24264 (N_24264,N_21907,N_21310);
nand U24265 (N_24265,N_22070,N_21798);
nor U24266 (N_24266,N_20057,N_21586);
and U24267 (N_24267,N_22337,N_22001);
xor U24268 (N_24268,N_21877,N_21353);
or U24269 (N_24269,N_20831,N_20353);
xor U24270 (N_24270,N_21614,N_20833);
nor U24271 (N_24271,N_20860,N_21160);
nand U24272 (N_24272,N_20228,N_22476);
xnor U24273 (N_24273,N_21274,N_20072);
and U24274 (N_24274,N_20751,N_21597);
nor U24275 (N_24275,N_20835,N_21618);
or U24276 (N_24276,N_20620,N_21103);
or U24277 (N_24277,N_21261,N_20459);
nor U24278 (N_24278,N_20320,N_20297);
nand U24279 (N_24279,N_21419,N_21031);
nor U24280 (N_24280,N_20983,N_21729);
nor U24281 (N_24281,N_20592,N_20958);
and U24282 (N_24282,N_22405,N_22193);
or U24283 (N_24283,N_21518,N_20305);
nor U24284 (N_24284,N_20717,N_21558);
and U24285 (N_24285,N_20494,N_20651);
nor U24286 (N_24286,N_21326,N_20784);
xor U24287 (N_24287,N_21890,N_20089);
xor U24288 (N_24288,N_21241,N_20776);
or U24289 (N_24289,N_20570,N_20325);
nand U24290 (N_24290,N_22184,N_21824);
or U24291 (N_24291,N_21261,N_20566);
or U24292 (N_24292,N_21555,N_20574);
or U24293 (N_24293,N_20962,N_21816);
xor U24294 (N_24294,N_21423,N_20810);
xnor U24295 (N_24295,N_20749,N_20727);
nor U24296 (N_24296,N_21626,N_21597);
or U24297 (N_24297,N_21866,N_20338);
and U24298 (N_24298,N_20606,N_22252);
or U24299 (N_24299,N_20688,N_20250);
xnor U24300 (N_24300,N_20886,N_21146);
or U24301 (N_24301,N_21451,N_21569);
or U24302 (N_24302,N_20188,N_22182);
and U24303 (N_24303,N_22116,N_20198);
and U24304 (N_24304,N_21495,N_21858);
nand U24305 (N_24305,N_21458,N_20450);
or U24306 (N_24306,N_21825,N_20894);
nand U24307 (N_24307,N_20655,N_20279);
xor U24308 (N_24308,N_22191,N_20964);
and U24309 (N_24309,N_21832,N_21304);
or U24310 (N_24310,N_21506,N_21441);
and U24311 (N_24311,N_21881,N_21888);
and U24312 (N_24312,N_20602,N_21249);
or U24313 (N_24313,N_22047,N_21581);
nand U24314 (N_24314,N_22071,N_20010);
nor U24315 (N_24315,N_21887,N_21241);
xor U24316 (N_24316,N_20431,N_20561);
or U24317 (N_24317,N_20348,N_21307);
or U24318 (N_24318,N_22361,N_21651);
nor U24319 (N_24319,N_22136,N_22036);
or U24320 (N_24320,N_22293,N_20326);
xnor U24321 (N_24321,N_20570,N_20158);
xor U24322 (N_24322,N_20918,N_21448);
nand U24323 (N_24323,N_22188,N_22053);
and U24324 (N_24324,N_20850,N_21738);
nor U24325 (N_24325,N_21157,N_22488);
nand U24326 (N_24326,N_21569,N_21135);
and U24327 (N_24327,N_21169,N_21731);
and U24328 (N_24328,N_21938,N_20523);
nand U24329 (N_24329,N_20381,N_21176);
nand U24330 (N_24330,N_21079,N_21086);
xor U24331 (N_24331,N_21480,N_20925);
xor U24332 (N_24332,N_20183,N_22097);
or U24333 (N_24333,N_21943,N_20343);
nand U24334 (N_24334,N_20009,N_20938);
and U24335 (N_24335,N_21797,N_22357);
nor U24336 (N_24336,N_22037,N_20855);
xor U24337 (N_24337,N_20509,N_20374);
nand U24338 (N_24338,N_21737,N_20047);
nand U24339 (N_24339,N_22391,N_21925);
xor U24340 (N_24340,N_21173,N_20386);
nor U24341 (N_24341,N_20386,N_20153);
and U24342 (N_24342,N_20621,N_22169);
or U24343 (N_24343,N_21166,N_20121);
xor U24344 (N_24344,N_20642,N_21029);
nor U24345 (N_24345,N_21791,N_20146);
nand U24346 (N_24346,N_22377,N_20373);
or U24347 (N_24347,N_20506,N_20914);
or U24348 (N_24348,N_22192,N_20425);
nor U24349 (N_24349,N_21180,N_21076);
xor U24350 (N_24350,N_20359,N_22105);
or U24351 (N_24351,N_22081,N_21736);
nand U24352 (N_24352,N_21081,N_22080);
or U24353 (N_24353,N_21271,N_20801);
xor U24354 (N_24354,N_21560,N_20574);
nand U24355 (N_24355,N_21404,N_21013);
nor U24356 (N_24356,N_22000,N_20846);
and U24357 (N_24357,N_21028,N_21227);
xor U24358 (N_24358,N_20288,N_20137);
nand U24359 (N_24359,N_21387,N_21110);
nand U24360 (N_24360,N_21307,N_21761);
nand U24361 (N_24361,N_22307,N_21602);
xor U24362 (N_24362,N_20247,N_22296);
nand U24363 (N_24363,N_20399,N_22456);
or U24364 (N_24364,N_21973,N_21852);
xnor U24365 (N_24365,N_21522,N_20892);
or U24366 (N_24366,N_20027,N_20421);
nand U24367 (N_24367,N_21834,N_21123);
or U24368 (N_24368,N_20855,N_20486);
nor U24369 (N_24369,N_21181,N_21355);
xor U24370 (N_24370,N_22409,N_22365);
nor U24371 (N_24371,N_21746,N_21949);
nand U24372 (N_24372,N_20659,N_20455);
nor U24373 (N_24373,N_21276,N_21509);
or U24374 (N_24374,N_20752,N_21907);
nor U24375 (N_24375,N_21945,N_22461);
nor U24376 (N_24376,N_21470,N_20090);
xor U24377 (N_24377,N_22110,N_21154);
or U24378 (N_24378,N_20534,N_20297);
xnor U24379 (N_24379,N_20436,N_20748);
or U24380 (N_24380,N_20339,N_20092);
nand U24381 (N_24381,N_21573,N_21182);
nor U24382 (N_24382,N_21671,N_20194);
nor U24383 (N_24383,N_20905,N_22197);
xnor U24384 (N_24384,N_20170,N_20543);
nand U24385 (N_24385,N_22331,N_20486);
nand U24386 (N_24386,N_21662,N_20273);
nor U24387 (N_24387,N_20106,N_21104);
xor U24388 (N_24388,N_21981,N_21815);
and U24389 (N_24389,N_20368,N_22320);
nor U24390 (N_24390,N_21947,N_21479);
nand U24391 (N_24391,N_22413,N_20977);
and U24392 (N_24392,N_20104,N_20749);
or U24393 (N_24393,N_22149,N_20578);
nand U24394 (N_24394,N_21886,N_20842);
xor U24395 (N_24395,N_21126,N_20506);
xnor U24396 (N_24396,N_21540,N_20212);
and U24397 (N_24397,N_21316,N_22065);
nand U24398 (N_24398,N_20632,N_21073);
nor U24399 (N_24399,N_21892,N_21964);
nand U24400 (N_24400,N_21417,N_21592);
or U24401 (N_24401,N_21357,N_20461);
nor U24402 (N_24402,N_21708,N_20037);
xor U24403 (N_24403,N_20265,N_21466);
or U24404 (N_24404,N_20763,N_21498);
or U24405 (N_24405,N_21683,N_21947);
xnor U24406 (N_24406,N_21698,N_20192);
and U24407 (N_24407,N_21687,N_20802);
and U24408 (N_24408,N_22270,N_21409);
nor U24409 (N_24409,N_20260,N_20916);
nor U24410 (N_24410,N_22306,N_21311);
nor U24411 (N_24411,N_22012,N_21736);
and U24412 (N_24412,N_20733,N_22102);
and U24413 (N_24413,N_22031,N_20463);
nor U24414 (N_24414,N_20436,N_20933);
xnor U24415 (N_24415,N_21145,N_20490);
or U24416 (N_24416,N_22302,N_20295);
xnor U24417 (N_24417,N_21679,N_21697);
or U24418 (N_24418,N_20194,N_21254);
nand U24419 (N_24419,N_20402,N_20567);
xor U24420 (N_24420,N_21823,N_21989);
xor U24421 (N_24421,N_20945,N_22288);
and U24422 (N_24422,N_20980,N_20530);
or U24423 (N_24423,N_22061,N_20501);
or U24424 (N_24424,N_22247,N_21419);
nand U24425 (N_24425,N_20557,N_21063);
nor U24426 (N_24426,N_21049,N_21117);
or U24427 (N_24427,N_20998,N_21451);
and U24428 (N_24428,N_22463,N_20384);
or U24429 (N_24429,N_20445,N_21160);
nand U24430 (N_24430,N_20621,N_20584);
xor U24431 (N_24431,N_20965,N_20411);
or U24432 (N_24432,N_21521,N_22409);
or U24433 (N_24433,N_20784,N_20257);
nand U24434 (N_24434,N_21835,N_20102);
xnor U24435 (N_24435,N_20169,N_21322);
nand U24436 (N_24436,N_20209,N_22489);
xor U24437 (N_24437,N_20327,N_20772);
and U24438 (N_24438,N_22340,N_20894);
and U24439 (N_24439,N_21728,N_21231);
or U24440 (N_24440,N_21591,N_22473);
nand U24441 (N_24441,N_22053,N_21308);
nor U24442 (N_24442,N_20681,N_21980);
nand U24443 (N_24443,N_22451,N_21327);
or U24444 (N_24444,N_20186,N_21731);
and U24445 (N_24445,N_21815,N_20619);
and U24446 (N_24446,N_21022,N_22303);
nor U24447 (N_24447,N_20843,N_20969);
and U24448 (N_24448,N_20029,N_20583);
and U24449 (N_24449,N_21352,N_21076);
xor U24450 (N_24450,N_21056,N_21713);
nand U24451 (N_24451,N_21802,N_22409);
xor U24452 (N_24452,N_21197,N_21758);
and U24453 (N_24453,N_20142,N_21585);
nor U24454 (N_24454,N_21770,N_22210);
xnor U24455 (N_24455,N_21523,N_22137);
or U24456 (N_24456,N_21032,N_20489);
and U24457 (N_24457,N_21858,N_22497);
nand U24458 (N_24458,N_21544,N_20178);
nand U24459 (N_24459,N_22423,N_21276);
or U24460 (N_24460,N_20096,N_20493);
or U24461 (N_24461,N_21046,N_20028);
nand U24462 (N_24462,N_21536,N_21903);
or U24463 (N_24463,N_21655,N_21780);
nor U24464 (N_24464,N_22238,N_21065);
or U24465 (N_24465,N_22170,N_22464);
and U24466 (N_24466,N_21977,N_21874);
nor U24467 (N_24467,N_21270,N_20987);
xor U24468 (N_24468,N_20700,N_21826);
or U24469 (N_24469,N_22117,N_21518);
nand U24470 (N_24470,N_21955,N_20464);
and U24471 (N_24471,N_21823,N_21228);
xnor U24472 (N_24472,N_22027,N_20613);
or U24473 (N_24473,N_21280,N_20268);
nand U24474 (N_24474,N_22492,N_21527);
and U24475 (N_24475,N_20238,N_20032);
nand U24476 (N_24476,N_20041,N_22287);
xor U24477 (N_24477,N_20451,N_20714);
or U24478 (N_24478,N_21454,N_21512);
and U24479 (N_24479,N_21132,N_21497);
xnor U24480 (N_24480,N_21661,N_21132);
nor U24481 (N_24481,N_20323,N_20538);
xor U24482 (N_24482,N_20835,N_22311);
nand U24483 (N_24483,N_20310,N_20872);
and U24484 (N_24484,N_21189,N_21237);
xnor U24485 (N_24485,N_20347,N_22089);
nand U24486 (N_24486,N_21619,N_21325);
nand U24487 (N_24487,N_22153,N_22122);
nor U24488 (N_24488,N_20870,N_20726);
xnor U24489 (N_24489,N_22246,N_21438);
and U24490 (N_24490,N_21768,N_21032);
nor U24491 (N_24491,N_21883,N_21784);
nor U24492 (N_24492,N_21482,N_21585);
and U24493 (N_24493,N_21563,N_20015);
xor U24494 (N_24494,N_20019,N_20320);
or U24495 (N_24495,N_21311,N_20217);
xor U24496 (N_24496,N_20653,N_21552);
or U24497 (N_24497,N_20271,N_20274);
or U24498 (N_24498,N_20022,N_21312);
and U24499 (N_24499,N_20163,N_20764);
nand U24500 (N_24500,N_20660,N_21388);
or U24501 (N_24501,N_20254,N_20348);
or U24502 (N_24502,N_20744,N_22166);
or U24503 (N_24503,N_21442,N_22407);
or U24504 (N_24504,N_20633,N_20852);
and U24505 (N_24505,N_20439,N_21643);
xor U24506 (N_24506,N_20214,N_21872);
nand U24507 (N_24507,N_21282,N_20195);
nor U24508 (N_24508,N_20687,N_21372);
and U24509 (N_24509,N_21898,N_20736);
nand U24510 (N_24510,N_20940,N_20871);
and U24511 (N_24511,N_21896,N_20212);
or U24512 (N_24512,N_21434,N_21810);
or U24513 (N_24513,N_20760,N_21558);
or U24514 (N_24514,N_21710,N_20755);
or U24515 (N_24515,N_21812,N_20001);
nor U24516 (N_24516,N_21516,N_20720);
and U24517 (N_24517,N_20402,N_20758);
xor U24518 (N_24518,N_21511,N_20657);
nor U24519 (N_24519,N_21678,N_20220);
xnor U24520 (N_24520,N_20578,N_22023);
or U24521 (N_24521,N_20738,N_21757);
and U24522 (N_24522,N_20953,N_22425);
nor U24523 (N_24523,N_21708,N_20819);
or U24524 (N_24524,N_20907,N_20112);
and U24525 (N_24525,N_22451,N_20508);
xnor U24526 (N_24526,N_22167,N_20418);
nand U24527 (N_24527,N_21500,N_22116);
nor U24528 (N_24528,N_20127,N_20747);
xnor U24529 (N_24529,N_22329,N_20885);
or U24530 (N_24530,N_21983,N_20887);
xor U24531 (N_24531,N_21771,N_21737);
or U24532 (N_24532,N_22187,N_20371);
nand U24533 (N_24533,N_20561,N_20094);
or U24534 (N_24534,N_21016,N_20994);
nor U24535 (N_24535,N_20139,N_20220);
nand U24536 (N_24536,N_20015,N_20719);
nand U24537 (N_24537,N_21363,N_20666);
nand U24538 (N_24538,N_21488,N_22260);
or U24539 (N_24539,N_21840,N_21244);
nand U24540 (N_24540,N_20751,N_22481);
nor U24541 (N_24541,N_21862,N_20968);
and U24542 (N_24542,N_21676,N_21406);
and U24543 (N_24543,N_21972,N_20343);
or U24544 (N_24544,N_22211,N_21297);
and U24545 (N_24545,N_20802,N_21267);
nor U24546 (N_24546,N_20852,N_21270);
nand U24547 (N_24547,N_20838,N_20688);
xnor U24548 (N_24548,N_22156,N_21212);
and U24549 (N_24549,N_20256,N_20914);
nand U24550 (N_24550,N_22190,N_20076);
and U24551 (N_24551,N_21078,N_21982);
nor U24552 (N_24552,N_20370,N_22242);
nand U24553 (N_24553,N_20287,N_20630);
or U24554 (N_24554,N_20009,N_22206);
nand U24555 (N_24555,N_20609,N_21409);
nand U24556 (N_24556,N_21558,N_22157);
nand U24557 (N_24557,N_21652,N_22468);
nor U24558 (N_24558,N_20402,N_21488);
and U24559 (N_24559,N_20765,N_21627);
and U24560 (N_24560,N_21238,N_20099);
nand U24561 (N_24561,N_20725,N_20077);
or U24562 (N_24562,N_22069,N_21492);
or U24563 (N_24563,N_20258,N_21512);
xor U24564 (N_24564,N_20278,N_21285);
and U24565 (N_24565,N_20587,N_20445);
nand U24566 (N_24566,N_20163,N_20303);
and U24567 (N_24567,N_21570,N_21898);
nor U24568 (N_24568,N_21689,N_22233);
and U24569 (N_24569,N_21622,N_21052);
nand U24570 (N_24570,N_20792,N_21161);
xnor U24571 (N_24571,N_22269,N_21495);
xor U24572 (N_24572,N_20781,N_20704);
or U24573 (N_24573,N_20845,N_21011);
and U24574 (N_24574,N_21207,N_20643);
nand U24575 (N_24575,N_20187,N_21758);
and U24576 (N_24576,N_20674,N_21220);
or U24577 (N_24577,N_20459,N_22384);
and U24578 (N_24578,N_20303,N_21208);
or U24579 (N_24579,N_20912,N_20180);
nor U24580 (N_24580,N_21995,N_20705);
or U24581 (N_24581,N_20928,N_22369);
xnor U24582 (N_24582,N_22404,N_21866);
and U24583 (N_24583,N_20218,N_20144);
and U24584 (N_24584,N_21394,N_20233);
nor U24585 (N_24585,N_21908,N_22423);
and U24586 (N_24586,N_22312,N_21858);
xnor U24587 (N_24587,N_22160,N_20164);
or U24588 (N_24588,N_21694,N_22264);
nand U24589 (N_24589,N_21489,N_21994);
or U24590 (N_24590,N_20002,N_21519);
and U24591 (N_24591,N_20056,N_21489);
xor U24592 (N_24592,N_22353,N_21980);
and U24593 (N_24593,N_22385,N_21087);
nand U24594 (N_24594,N_21371,N_20504);
nor U24595 (N_24595,N_20907,N_22440);
or U24596 (N_24596,N_21737,N_20781);
xnor U24597 (N_24597,N_20798,N_21917);
or U24598 (N_24598,N_20353,N_20238);
and U24599 (N_24599,N_20016,N_21072);
and U24600 (N_24600,N_20523,N_21381);
nand U24601 (N_24601,N_21880,N_22072);
and U24602 (N_24602,N_21831,N_20548);
and U24603 (N_24603,N_22315,N_20955);
and U24604 (N_24604,N_21492,N_21309);
and U24605 (N_24605,N_21848,N_21411);
nand U24606 (N_24606,N_21759,N_20114);
nor U24607 (N_24607,N_20729,N_21401);
xnor U24608 (N_24608,N_21099,N_21860);
and U24609 (N_24609,N_20559,N_21465);
and U24610 (N_24610,N_21682,N_21441);
nand U24611 (N_24611,N_21332,N_21110);
nor U24612 (N_24612,N_21603,N_20667);
nand U24613 (N_24613,N_22069,N_20365);
nor U24614 (N_24614,N_20993,N_20709);
and U24615 (N_24615,N_20541,N_20640);
or U24616 (N_24616,N_20026,N_21558);
and U24617 (N_24617,N_22275,N_20532);
and U24618 (N_24618,N_20193,N_20308);
xnor U24619 (N_24619,N_21034,N_22157);
and U24620 (N_24620,N_20993,N_22236);
nand U24621 (N_24621,N_21789,N_20177);
and U24622 (N_24622,N_20609,N_20829);
nand U24623 (N_24623,N_20107,N_21666);
nor U24624 (N_24624,N_20443,N_22260);
nand U24625 (N_24625,N_21414,N_21816);
nand U24626 (N_24626,N_21259,N_21397);
and U24627 (N_24627,N_22216,N_21417);
and U24628 (N_24628,N_22420,N_20690);
and U24629 (N_24629,N_22020,N_20269);
xor U24630 (N_24630,N_20965,N_21972);
nor U24631 (N_24631,N_21777,N_21502);
and U24632 (N_24632,N_20346,N_20492);
nand U24633 (N_24633,N_21477,N_22096);
or U24634 (N_24634,N_20913,N_22000);
and U24635 (N_24635,N_20524,N_21050);
nor U24636 (N_24636,N_21216,N_21500);
nand U24637 (N_24637,N_22288,N_21824);
nand U24638 (N_24638,N_21863,N_21789);
xnor U24639 (N_24639,N_20413,N_22131);
nand U24640 (N_24640,N_22204,N_21651);
nor U24641 (N_24641,N_20233,N_20136);
or U24642 (N_24642,N_21391,N_20281);
nor U24643 (N_24643,N_20979,N_20521);
and U24644 (N_24644,N_20779,N_20809);
nor U24645 (N_24645,N_21455,N_20714);
nor U24646 (N_24646,N_21392,N_22341);
nor U24647 (N_24647,N_20505,N_20470);
xor U24648 (N_24648,N_20214,N_21394);
and U24649 (N_24649,N_21348,N_20019);
and U24650 (N_24650,N_21584,N_21342);
and U24651 (N_24651,N_22235,N_22166);
or U24652 (N_24652,N_20649,N_20347);
or U24653 (N_24653,N_22235,N_21038);
nand U24654 (N_24654,N_20315,N_22244);
xor U24655 (N_24655,N_20198,N_20601);
nor U24656 (N_24656,N_20694,N_20515);
and U24657 (N_24657,N_20662,N_20463);
xor U24658 (N_24658,N_20820,N_21945);
nor U24659 (N_24659,N_22197,N_22429);
xor U24660 (N_24660,N_21340,N_21770);
nand U24661 (N_24661,N_20828,N_20280);
nor U24662 (N_24662,N_22251,N_20791);
and U24663 (N_24663,N_20410,N_21561);
nand U24664 (N_24664,N_20881,N_21170);
nor U24665 (N_24665,N_20183,N_22243);
and U24666 (N_24666,N_21000,N_20435);
nor U24667 (N_24667,N_20759,N_20908);
xnor U24668 (N_24668,N_22499,N_20332);
xor U24669 (N_24669,N_21840,N_22035);
nor U24670 (N_24670,N_22239,N_21681);
nor U24671 (N_24671,N_20074,N_21246);
nor U24672 (N_24672,N_22493,N_20418);
and U24673 (N_24673,N_21059,N_21073);
or U24674 (N_24674,N_21674,N_21439);
and U24675 (N_24675,N_22491,N_22018);
xor U24676 (N_24676,N_22268,N_20335);
or U24677 (N_24677,N_21193,N_21591);
xnor U24678 (N_24678,N_22109,N_21870);
and U24679 (N_24679,N_22049,N_21543);
xnor U24680 (N_24680,N_20655,N_21463);
or U24681 (N_24681,N_20340,N_21695);
and U24682 (N_24682,N_20931,N_21284);
nand U24683 (N_24683,N_20779,N_21782);
and U24684 (N_24684,N_22282,N_20256);
nor U24685 (N_24685,N_20188,N_21454);
or U24686 (N_24686,N_21243,N_21360);
nand U24687 (N_24687,N_21262,N_21084);
xnor U24688 (N_24688,N_21164,N_21729);
nor U24689 (N_24689,N_22338,N_21523);
nor U24690 (N_24690,N_20875,N_22044);
nor U24691 (N_24691,N_21830,N_21157);
xnor U24692 (N_24692,N_20880,N_21835);
xnor U24693 (N_24693,N_21564,N_21076);
nand U24694 (N_24694,N_22077,N_21656);
and U24695 (N_24695,N_20112,N_22102);
or U24696 (N_24696,N_20504,N_21985);
nor U24697 (N_24697,N_20368,N_21186);
or U24698 (N_24698,N_20708,N_21443);
or U24699 (N_24699,N_20892,N_20585);
nor U24700 (N_24700,N_21349,N_22270);
nor U24701 (N_24701,N_21224,N_21814);
nand U24702 (N_24702,N_22099,N_20161);
nor U24703 (N_24703,N_20579,N_21150);
and U24704 (N_24704,N_22337,N_20800);
xor U24705 (N_24705,N_22111,N_21799);
nor U24706 (N_24706,N_21949,N_22198);
and U24707 (N_24707,N_20589,N_20558);
nor U24708 (N_24708,N_20652,N_20695);
nor U24709 (N_24709,N_20553,N_20209);
or U24710 (N_24710,N_20877,N_21195);
or U24711 (N_24711,N_22103,N_20787);
nand U24712 (N_24712,N_20230,N_21437);
nor U24713 (N_24713,N_21581,N_20798);
and U24714 (N_24714,N_21506,N_20675);
or U24715 (N_24715,N_20167,N_20275);
nand U24716 (N_24716,N_21006,N_22113);
xor U24717 (N_24717,N_21623,N_22141);
nand U24718 (N_24718,N_20418,N_20022);
or U24719 (N_24719,N_22399,N_21679);
and U24720 (N_24720,N_21158,N_20126);
xor U24721 (N_24721,N_21954,N_20713);
and U24722 (N_24722,N_21805,N_22076);
nand U24723 (N_24723,N_22475,N_21416);
nor U24724 (N_24724,N_21341,N_21838);
or U24725 (N_24725,N_22072,N_21023);
and U24726 (N_24726,N_20087,N_20375);
or U24727 (N_24727,N_22176,N_21777);
nand U24728 (N_24728,N_21883,N_21803);
xnor U24729 (N_24729,N_21144,N_22254);
or U24730 (N_24730,N_20197,N_22275);
or U24731 (N_24731,N_20928,N_20795);
or U24732 (N_24732,N_20183,N_20249);
xor U24733 (N_24733,N_21529,N_21213);
or U24734 (N_24734,N_20564,N_21472);
nand U24735 (N_24735,N_21210,N_20634);
xnor U24736 (N_24736,N_21842,N_21355);
or U24737 (N_24737,N_20553,N_20773);
or U24738 (N_24738,N_20622,N_20426);
nor U24739 (N_24739,N_21453,N_21085);
and U24740 (N_24740,N_21894,N_20252);
or U24741 (N_24741,N_22122,N_21473);
nand U24742 (N_24742,N_21480,N_20667);
nor U24743 (N_24743,N_21094,N_21738);
and U24744 (N_24744,N_22090,N_21653);
xor U24745 (N_24745,N_21289,N_22005);
or U24746 (N_24746,N_21295,N_20912);
nor U24747 (N_24747,N_21105,N_22094);
or U24748 (N_24748,N_20412,N_21474);
nand U24749 (N_24749,N_21931,N_22473);
xnor U24750 (N_24750,N_20926,N_20439);
or U24751 (N_24751,N_20896,N_20985);
xnor U24752 (N_24752,N_22077,N_20645);
or U24753 (N_24753,N_21903,N_20706);
xnor U24754 (N_24754,N_21188,N_20496);
nor U24755 (N_24755,N_20536,N_21033);
xor U24756 (N_24756,N_22124,N_21390);
or U24757 (N_24757,N_20480,N_21390);
nor U24758 (N_24758,N_20024,N_21091);
nand U24759 (N_24759,N_21515,N_22043);
nor U24760 (N_24760,N_21659,N_22348);
nor U24761 (N_24761,N_20053,N_22186);
xnor U24762 (N_24762,N_20805,N_22229);
xnor U24763 (N_24763,N_20006,N_21399);
or U24764 (N_24764,N_21474,N_22339);
xor U24765 (N_24765,N_20203,N_20699);
and U24766 (N_24766,N_20843,N_20084);
and U24767 (N_24767,N_20281,N_21068);
nor U24768 (N_24768,N_20298,N_20485);
xor U24769 (N_24769,N_21824,N_21723);
and U24770 (N_24770,N_22440,N_20193);
and U24771 (N_24771,N_20225,N_21628);
or U24772 (N_24772,N_21602,N_20808);
nand U24773 (N_24773,N_21406,N_20296);
nor U24774 (N_24774,N_20662,N_21435);
nand U24775 (N_24775,N_21549,N_21353);
and U24776 (N_24776,N_20989,N_21170);
xnor U24777 (N_24777,N_21703,N_21686);
xnor U24778 (N_24778,N_22464,N_20930);
and U24779 (N_24779,N_22060,N_21033);
or U24780 (N_24780,N_21406,N_22129);
nand U24781 (N_24781,N_21114,N_20349);
and U24782 (N_24782,N_21607,N_21139);
xnor U24783 (N_24783,N_20742,N_20223);
xor U24784 (N_24784,N_21641,N_21648);
nand U24785 (N_24785,N_20804,N_21568);
or U24786 (N_24786,N_20424,N_20478);
nor U24787 (N_24787,N_20744,N_20262);
nor U24788 (N_24788,N_21198,N_22232);
nand U24789 (N_24789,N_21553,N_20407);
or U24790 (N_24790,N_21637,N_22401);
xnor U24791 (N_24791,N_22301,N_21544);
xor U24792 (N_24792,N_22413,N_22240);
nor U24793 (N_24793,N_22094,N_22292);
xor U24794 (N_24794,N_20940,N_21940);
and U24795 (N_24795,N_20117,N_21443);
or U24796 (N_24796,N_20977,N_21433);
and U24797 (N_24797,N_22237,N_20569);
and U24798 (N_24798,N_20194,N_20219);
and U24799 (N_24799,N_22165,N_20239);
nand U24800 (N_24800,N_21483,N_22464);
nor U24801 (N_24801,N_22028,N_21944);
nand U24802 (N_24802,N_22202,N_20625);
and U24803 (N_24803,N_21247,N_22157);
or U24804 (N_24804,N_20138,N_20270);
nand U24805 (N_24805,N_21229,N_22497);
nor U24806 (N_24806,N_20224,N_21930);
nor U24807 (N_24807,N_20165,N_21500);
or U24808 (N_24808,N_21253,N_20726);
and U24809 (N_24809,N_22161,N_21719);
nand U24810 (N_24810,N_20450,N_20811);
xor U24811 (N_24811,N_20912,N_20752);
or U24812 (N_24812,N_21985,N_21195);
nand U24813 (N_24813,N_22409,N_21900);
and U24814 (N_24814,N_20531,N_21057);
nor U24815 (N_24815,N_21740,N_20317);
nor U24816 (N_24816,N_22073,N_21932);
nor U24817 (N_24817,N_21289,N_20378);
or U24818 (N_24818,N_20988,N_22123);
nor U24819 (N_24819,N_20968,N_20254);
or U24820 (N_24820,N_22302,N_21727);
or U24821 (N_24821,N_20112,N_21879);
or U24822 (N_24822,N_21184,N_20182);
nand U24823 (N_24823,N_20155,N_21590);
or U24824 (N_24824,N_21525,N_21069);
nand U24825 (N_24825,N_21982,N_20892);
and U24826 (N_24826,N_21793,N_20643);
xnor U24827 (N_24827,N_21205,N_21311);
and U24828 (N_24828,N_21763,N_21067);
xor U24829 (N_24829,N_21940,N_22167);
or U24830 (N_24830,N_20853,N_20028);
nor U24831 (N_24831,N_20960,N_20223);
and U24832 (N_24832,N_20515,N_22487);
xor U24833 (N_24833,N_20179,N_21256);
or U24834 (N_24834,N_21847,N_20775);
or U24835 (N_24835,N_20635,N_22051);
xor U24836 (N_24836,N_20884,N_20848);
nand U24837 (N_24837,N_22423,N_21167);
xor U24838 (N_24838,N_21861,N_20803);
xor U24839 (N_24839,N_21601,N_22130);
xnor U24840 (N_24840,N_20364,N_22488);
nor U24841 (N_24841,N_20506,N_21240);
nor U24842 (N_24842,N_22060,N_22133);
nor U24843 (N_24843,N_21371,N_21777);
and U24844 (N_24844,N_20701,N_21188);
nand U24845 (N_24845,N_20165,N_20302);
nor U24846 (N_24846,N_21707,N_20852);
xnor U24847 (N_24847,N_20102,N_21747);
nand U24848 (N_24848,N_21848,N_20079);
and U24849 (N_24849,N_20662,N_21264);
nor U24850 (N_24850,N_20653,N_21574);
and U24851 (N_24851,N_22458,N_21374);
or U24852 (N_24852,N_20071,N_20081);
nor U24853 (N_24853,N_22371,N_20678);
nor U24854 (N_24854,N_20970,N_21348);
nand U24855 (N_24855,N_21857,N_21296);
and U24856 (N_24856,N_20837,N_21647);
nand U24857 (N_24857,N_20872,N_21378);
xor U24858 (N_24858,N_21173,N_20604);
xnor U24859 (N_24859,N_21963,N_21356);
nand U24860 (N_24860,N_22368,N_20838);
and U24861 (N_24861,N_21785,N_20521);
xnor U24862 (N_24862,N_20750,N_22069);
xnor U24863 (N_24863,N_21012,N_21030);
nand U24864 (N_24864,N_22268,N_20140);
xnor U24865 (N_24865,N_20906,N_20128);
or U24866 (N_24866,N_20957,N_20436);
and U24867 (N_24867,N_21995,N_20957);
nand U24868 (N_24868,N_20745,N_20101);
and U24869 (N_24869,N_21830,N_22228);
nor U24870 (N_24870,N_21672,N_21206);
xnor U24871 (N_24871,N_21361,N_20884);
nor U24872 (N_24872,N_20494,N_22032);
and U24873 (N_24873,N_21708,N_21386);
nor U24874 (N_24874,N_20666,N_20999);
xnor U24875 (N_24875,N_20272,N_21979);
xnor U24876 (N_24876,N_21685,N_22266);
or U24877 (N_24877,N_20523,N_20801);
nand U24878 (N_24878,N_20555,N_22221);
xnor U24879 (N_24879,N_21361,N_20443);
xnor U24880 (N_24880,N_20437,N_20446);
xor U24881 (N_24881,N_21748,N_21686);
nor U24882 (N_24882,N_20400,N_21231);
nand U24883 (N_24883,N_20649,N_20118);
nor U24884 (N_24884,N_20021,N_21572);
and U24885 (N_24885,N_21010,N_21816);
or U24886 (N_24886,N_21998,N_21069);
and U24887 (N_24887,N_21429,N_21393);
nand U24888 (N_24888,N_20734,N_21590);
nand U24889 (N_24889,N_21609,N_21524);
nor U24890 (N_24890,N_21341,N_20479);
or U24891 (N_24891,N_21797,N_22414);
or U24892 (N_24892,N_20049,N_21906);
or U24893 (N_24893,N_21713,N_21118);
and U24894 (N_24894,N_22107,N_21227);
or U24895 (N_24895,N_21659,N_21426);
or U24896 (N_24896,N_21200,N_21948);
nand U24897 (N_24897,N_22304,N_21142);
and U24898 (N_24898,N_21378,N_21127);
nor U24899 (N_24899,N_20784,N_20745);
nor U24900 (N_24900,N_22286,N_21761);
nand U24901 (N_24901,N_20746,N_22330);
nor U24902 (N_24902,N_20729,N_20744);
nor U24903 (N_24903,N_20474,N_21133);
or U24904 (N_24904,N_20244,N_21374);
nand U24905 (N_24905,N_20263,N_22330);
nor U24906 (N_24906,N_20496,N_21738);
and U24907 (N_24907,N_21829,N_22379);
xor U24908 (N_24908,N_21765,N_20936);
nor U24909 (N_24909,N_20069,N_22243);
or U24910 (N_24910,N_20607,N_22186);
xor U24911 (N_24911,N_21484,N_21255);
and U24912 (N_24912,N_21884,N_21669);
nor U24913 (N_24913,N_21354,N_20590);
and U24914 (N_24914,N_20471,N_20741);
and U24915 (N_24915,N_20109,N_21212);
nor U24916 (N_24916,N_21959,N_21004);
xnor U24917 (N_24917,N_22108,N_22124);
and U24918 (N_24918,N_22190,N_22400);
xor U24919 (N_24919,N_20026,N_21872);
nand U24920 (N_24920,N_20804,N_21676);
nand U24921 (N_24921,N_20052,N_20962);
nor U24922 (N_24922,N_20991,N_21195);
nor U24923 (N_24923,N_20127,N_20343);
xnor U24924 (N_24924,N_20402,N_20066);
or U24925 (N_24925,N_21507,N_22392);
xor U24926 (N_24926,N_22362,N_21732);
and U24927 (N_24927,N_22118,N_21139);
or U24928 (N_24928,N_21216,N_20583);
nor U24929 (N_24929,N_22398,N_20230);
xor U24930 (N_24930,N_20826,N_20436);
or U24931 (N_24931,N_20081,N_20511);
nand U24932 (N_24932,N_22137,N_20561);
or U24933 (N_24933,N_20081,N_22374);
nor U24934 (N_24934,N_20359,N_21262);
nor U24935 (N_24935,N_20710,N_21111);
and U24936 (N_24936,N_20696,N_21891);
nor U24937 (N_24937,N_20174,N_20009);
nand U24938 (N_24938,N_21376,N_22106);
or U24939 (N_24939,N_21573,N_20516);
and U24940 (N_24940,N_20459,N_22408);
nor U24941 (N_24941,N_21985,N_22163);
nand U24942 (N_24942,N_20343,N_20876);
xor U24943 (N_24943,N_21470,N_20522);
xnor U24944 (N_24944,N_20571,N_20693);
nand U24945 (N_24945,N_20871,N_20017);
or U24946 (N_24946,N_20692,N_21919);
and U24947 (N_24947,N_20987,N_21113);
and U24948 (N_24948,N_21356,N_20544);
nor U24949 (N_24949,N_20446,N_22302);
xnor U24950 (N_24950,N_22073,N_20067);
or U24951 (N_24951,N_21132,N_20237);
xnor U24952 (N_24952,N_20819,N_21237);
xnor U24953 (N_24953,N_22237,N_21897);
or U24954 (N_24954,N_22346,N_20483);
nand U24955 (N_24955,N_21144,N_21469);
nor U24956 (N_24956,N_20555,N_20440);
and U24957 (N_24957,N_20778,N_22141);
xnor U24958 (N_24958,N_22488,N_20122);
or U24959 (N_24959,N_22240,N_20746);
nand U24960 (N_24960,N_20276,N_20447);
nor U24961 (N_24961,N_21883,N_21196);
and U24962 (N_24962,N_20101,N_20395);
and U24963 (N_24963,N_20445,N_22332);
and U24964 (N_24964,N_20653,N_22079);
or U24965 (N_24965,N_22200,N_21340);
or U24966 (N_24966,N_20738,N_21575);
nor U24967 (N_24967,N_21781,N_20655);
xor U24968 (N_24968,N_22088,N_20844);
nor U24969 (N_24969,N_21835,N_21075);
xor U24970 (N_24970,N_21934,N_21297);
nand U24971 (N_24971,N_21223,N_21981);
nand U24972 (N_24972,N_21089,N_21794);
or U24973 (N_24973,N_22034,N_22018);
xor U24974 (N_24974,N_22499,N_21979);
xnor U24975 (N_24975,N_20113,N_20593);
and U24976 (N_24976,N_20636,N_22427);
and U24977 (N_24977,N_21616,N_20540);
nor U24978 (N_24978,N_21690,N_21262);
nand U24979 (N_24979,N_21069,N_21357);
nand U24980 (N_24980,N_22462,N_21838);
nand U24981 (N_24981,N_20562,N_20451);
or U24982 (N_24982,N_22043,N_20427);
or U24983 (N_24983,N_21494,N_22228);
and U24984 (N_24984,N_21020,N_22406);
xor U24985 (N_24985,N_20880,N_22245);
and U24986 (N_24986,N_20833,N_21566);
nand U24987 (N_24987,N_21891,N_21870);
xnor U24988 (N_24988,N_22203,N_20125);
nand U24989 (N_24989,N_20110,N_20160);
nor U24990 (N_24990,N_20929,N_20683);
nor U24991 (N_24991,N_20136,N_20808);
nand U24992 (N_24992,N_21824,N_22071);
nor U24993 (N_24993,N_20019,N_20127);
nand U24994 (N_24994,N_20133,N_21271);
nor U24995 (N_24995,N_20298,N_21218);
or U24996 (N_24996,N_20349,N_21505);
xor U24997 (N_24997,N_20734,N_21884);
nand U24998 (N_24998,N_22074,N_21069);
and U24999 (N_24999,N_21791,N_21363);
or U25000 (N_25000,N_24527,N_23540);
and U25001 (N_25001,N_23880,N_23508);
nand U25002 (N_25002,N_22621,N_24694);
nor U25003 (N_25003,N_23626,N_23425);
nor U25004 (N_25004,N_24646,N_23891);
nand U25005 (N_25005,N_22995,N_24530);
nand U25006 (N_25006,N_23906,N_23661);
and U25007 (N_25007,N_23590,N_23799);
and U25008 (N_25008,N_24259,N_24939);
nand U25009 (N_25009,N_22737,N_23336);
nor U25010 (N_25010,N_24962,N_23472);
nor U25011 (N_25011,N_22680,N_24461);
nor U25012 (N_25012,N_22665,N_23178);
nor U25013 (N_25013,N_24675,N_24546);
xnor U25014 (N_25014,N_24520,N_23379);
or U25015 (N_25015,N_23409,N_23471);
or U25016 (N_25016,N_23618,N_24576);
xor U25017 (N_25017,N_22856,N_23610);
nand U25018 (N_25018,N_22527,N_24777);
or U25019 (N_25019,N_23196,N_23313);
and U25020 (N_25020,N_23845,N_24519);
nor U25021 (N_25021,N_24674,N_23652);
and U25022 (N_25022,N_23459,N_23375);
xnor U25023 (N_25023,N_24376,N_23838);
nand U25024 (N_25024,N_23867,N_22566);
and U25025 (N_25025,N_23453,N_23953);
nand U25026 (N_25026,N_23023,N_24008);
xnor U25027 (N_25027,N_24426,N_23837);
xnor U25028 (N_25028,N_23377,N_24915);
nor U25029 (N_25029,N_22874,N_23355);
nand U25030 (N_25030,N_24014,N_22689);
nor U25031 (N_25031,N_24507,N_24806);
or U25032 (N_25032,N_22518,N_23172);
nor U25033 (N_25033,N_23272,N_24936);
xnor U25034 (N_25034,N_22637,N_23300);
and U25035 (N_25035,N_24400,N_22557);
xnor U25036 (N_25036,N_22952,N_23089);
or U25037 (N_25037,N_24882,N_24130);
nor U25038 (N_25038,N_24528,N_24811);
nor U25039 (N_25039,N_23018,N_23996);
nor U25040 (N_25040,N_24825,N_24748);
nor U25041 (N_25041,N_24625,N_23246);
xor U25042 (N_25042,N_23124,N_24132);
nand U25043 (N_25043,N_22533,N_24518);
or U25044 (N_25044,N_24542,N_23116);
nor U25045 (N_25045,N_23117,N_23285);
nand U25046 (N_25046,N_24592,N_24558);
nor U25047 (N_25047,N_23636,N_24954);
nor U25048 (N_25048,N_23668,N_24328);
xnor U25049 (N_25049,N_24466,N_24891);
xor U25050 (N_25050,N_23020,N_24900);
nand U25051 (N_25051,N_23977,N_23734);
nor U25052 (N_25052,N_24185,N_22537);
nand U25053 (N_25053,N_23176,N_22605);
xor U25054 (N_25054,N_23782,N_24499);
nand U25055 (N_25055,N_24651,N_22751);
and U25056 (N_25056,N_23105,N_22649);
or U25057 (N_25057,N_24738,N_23950);
xnor U25058 (N_25058,N_23119,N_23936);
xnor U25059 (N_25059,N_23536,N_24683);
or U25060 (N_25060,N_23726,N_24015);
and U25061 (N_25061,N_22611,N_23570);
nor U25062 (N_25062,N_23710,N_24053);
and U25063 (N_25063,N_24199,N_24335);
nor U25064 (N_25064,N_24222,N_24492);
and U25065 (N_25065,N_23299,N_22642);
and U25066 (N_25066,N_24813,N_23824);
xnor U25067 (N_25067,N_23964,N_23476);
and U25068 (N_25068,N_24575,N_24975);
or U25069 (N_25069,N_23433,N_22812);
xnor U25070 (N_25070,N_23639,N_23650);
nor U25071 (N_25071,N_23582,N_24427);
nand U25072 (N_25072,N_23421,N_24039);
or U25073 (N_25073,N_24658,N_23467);
or U25074 (N_25074,N_23776,N_22943);
xnor U25075 (N_25075,N_23888,N_23623);
or U25076 (N_25076,N_22722,N_23963);
nand U25077 (N_25077,N_24458,N_22937);
xor U25078 (N_25078,N_22854,N_23737);
or U25079 (N_25079,N_24317,N_23941);
nand U25080 (N_25080,N_23656,N_23644);
or U25081 (N_25081,N_24456,N_23454);
nand U25082 (N_25082,N_24380,N_24161);
nor U25083 (N_25083,N_23307,N_23199);
nor U25084 (N_25084,N_23609,N_22789);
and U25085 (N_25085,N_23957,N_24559);
or U25086 (N_25086,N_23431,N_24513);
or U25087 (N_25087,N_23037,N_24122);
and U25088 (N_25088,N_22626,N_23062);
nor U25089 (N_25089,N_23429,N_24163);
nor U25090 (N_25090,N_22852,N_24739);
xor U25091 (N_25091,N_24701,N_24260);
xor U25092 (N_25092,N_23797,N_22643);
nor U25093 (N_25093,N_22652,N_24961);
xnor U25094 (N_25094,N_23702,N_23632);
nor U25095 (N_25095,N_24733,N_22586);
xor U25096 (N_25096,N_24171,N_23000);
nand U25097 (N_25097,N_24393,N_23095);
and U25098 (N_25098,N_24689,N_24460);
nand U25099 (N_25099,N_24843,N_24211);
nand U25100 (N_25100,N_22926,N_23059);
nor U25101 (N_25101,N_23374,N_24996);
and U25102 (N_25102,N_24781,N_22880);
nor U25103 (N_25103,N_22699,N_24440);
nand U25104 (N_25104,N_24055,N_23600);
nor U25105 (N_25105,N_24106,N_24157);
xnor U25106 (N_25106,N_23149,N_23744);
and U25107 (N_25107,N_24602,N_22738);
nand U25108 (N_25108,N_22734,N_24190);
nor U25109 (N_25109,N_23677,N_24343);
or U25110 (N_25110,N_23088,N_22500);
or U25111 (N_25111,N_23629,N_23279);
nor U25112 (N_25112,N_24668,N_23860);
or U25113 (N_25113,N_22771,N_23542);
xnor U25114 (N_25114,N_24946,N_24833);
nor U25115 (N_25115,N_23039,N_22976);
xor U25116 (N_25116,N_23514,N_23318);
nand U25117 (N_25117,N_22992,N_22598);
nand U25118 (N_25118,N_24150,N_22645);
and U25119 (N_25119,N_23794,N_24858);
or U25120 (N_25120,N_24917,N_23589);
nor U25121 (N_25121,N_24242,N_24956);
nor U25122 (N_25122,N_23356,N_23158);
nand U25123 (N_25123,N_24792,N_23614);
and U25124 (N_25124,N_23993,N_22530);
nand U25125 (N_25125,N_23877,N_22761);
nand U25126 (N_25126,N_24567,N_23136);
nand U25127 (N_25127,N_23143,N_23491);
xor U25128 (N_25128,N_24787,N_24444);
nand U25129 (N_25129,N_24824,N_22668);
nand U25130 (N_25130,N_24045,N_24652);
nand U25131 (N_25131,N_24056,N_23649);
or U25132 (N_25132,N_23730,N_23451);
nand U25133 (N_25133,N_23883,N_24860);
nor U25134 (N_25134,N_24820,N_22932);
or U25135 (N_25135,N_23813,N_22818);
xor U25136 (N_25136,N_23593,N_23319);
xor U25137 (N_25137,N_23567,N_23364);
and U25138 (N_25138,N_23897,N_23351);
nand U25139 (N_25139,N_22661,N_24449);
nand U25140 (N_25140,N_24502,N_23282);
xor U25141 (N_25141,N_23306,N_23248);
nor U25142 (N_25142,N_22747,N_23738);
and U25143 (N_25143,N_23648,N_24310);
nor U25144 (N_25144,N_24435,N_22785);
nor U25145 (N_25145,N_24959,N_22938);
or U25146 (N_25146,N_23865,N_23495);
or U25147 (N_25147,N_22563,N_23752);
xor U25148 (N_25148,N_23747,N_24623);
and U25149 (N_25149,N_24578,N_23006);
nand U25150 (N_25150,N_23297,N_24639);
and U25151 (N_25151,N_24062,N_22630);
or U25152 (N_25152,N_23750,N_24415);
nor U25153 (N_25153,N_24454,N_24491);
xnor U25154 (N_25154,N_24475,N_22646);
nand U25155 (N_25155,N_24005,N_22591);
nand U25156 (N_25156,N_24077,N_22855);
or U25157 (N_25157,N_23305,N_23569);
nor U25158 (N_25158,N_24798,N_23893);
xor U25159 (N_25159,N_24043,N_22617);
xnor U25160 (N_25160,N_22982,N_23790);
xnor U25161 (N_25161,N_24702,N_24712);
nand U25162 (N_25162,N_24284,N_23541);
or U25163 (N_25163,N_23532,N_23826);
nand U25164 (N_25164,N_22569,N_23952);
and U25165 (N_25165,N_24918,N_24387);
and U25166 (N_25166,N_23742,N_24204);
and U25167 (N_25167,N_23915,N_24133);
xnor U25168 (N_25168,N_22583,N_23245);
xnor U25169 (N_25169,N_22987,N_23024);
or U25170 (N_25170,N_22956,N_23271);
nor U25171 (N_25171,N_24590,N_24110);
nand U25172 (N_25172,N_23159,N_22687);
and U25173 (N_25173,N_23327,N_23256);
or U25174 (N_25174,N_23916,N_24238);
nor U25175 (N_25175,N_24921,N_24670);
nand U25176 (N_25176,N_22748,N_23662);
or U25177 (N_25177,N_23718,N_24898);
xor U25178 (N_25178,N_23751,N_23745);
nor U25179 (N_25179,N_24972,N_22593);
nand U25180 (N_25180,N_24753,N_24883);
nand U25181 (N_25181,N_23690,N_23320);
or U25182 (N_25182,N_22596,N_24448);
or U25183 (N_25183,N_22715,N_22823);
xor U25184 (N_25184,N_22554,N_24589);
xor U25185 (N_25185,N_22623,N_22775);
nand U25186 (N_25186,N_23337,N_24455);
nor U25187 (N_25187,N_22931,N_22669);
xnor U25188 (N_25188,N_22870,N_24124);
or U25189 (N_25189,N_24246,N_23721);
nand U25190 (N_25190,N_24060,N_23693);
nand U25191 (N_25191,N_23554,N_24805);
nor U25192 (N_25192,N_24141,N_22894);
and U25193 (N_25193,N_24618,N_23414);
or U25194 (N_25194,N_23910,N_24919);
xor U25195 (N_25195,N_24731,N_23348);
nand U25196 (N_25196,N_24913,N_24275);
nor U25197 (N_25197,N_23358,N_22519);
xnor U25198 (N_25198,N_23383,N_22769);
and U25199 (N_25199,N_22824,N_22595);
or U25200 (N_25200,N_24501,N_23251);
or U25201 (N_25201,N_22825,N_22887);
nor U25202 (N_25202,N_24566,N_23907);
and U25203 (N_25203,N_24756,N_24930);
or U25204 (N_25204,N_23148,N_24600);
nand U25205 (N_25205,N_22736,N_24561);
or U25206 (N_25206,N_23455,N_22845);
nor U25207 (N_25207,N_23968,N_24299);
nor U25208 (N_25208,N_24363,N_23654);
or U25209 (N_25209,N_24245,N_24247);
or U25210 (N_25210,N_23268,N_23970);
and U25211 (N_25211,N_24102,N_24904);
and U25212 (N_25212,N_22828,N_24421);
nand U25213 (N_25213,N_23557,N_23233);
and U25214 (N_25214,N_22838,N_23505);
and U25215 (N_25215,N_22857,N_22817);
nor U25216 (N_25216,N_22889,N_24484);
nor U25217 (N_25217,N_22872,N_23868);
and U25218 (N_25218,N_24337,N_23349);
nand U25219 (N_25219,N_24306,N_24654);
nand U25220 (N_25220,N_22905,N_24752);
xor U25221 (N_25221,N_24321,N_23887);
nand U25222 (N_25222,N_22981,N_24661);
and U25223 (N_25223,N_23174,N_23703);
or U25224 (N_25224,N_24438,N_23100);
xnor U25225 (N_25225,N_24534,N_24793);
nor U25226 (N_25226,N_23956,N_24944);
nand U25227 (N_25227,N_23154,N_22978);
xor U25228 (N_25228,N_24740,N_24927);
and U25229 (N_25229,N_23722,N_24751);
nor U25230 (N_25230,N_23852,N_23680);
or U25231 (N_25231,N_24319,N_22890);
xnor U25232 (N_25232,N_24660,N_23736);
nor U25233 (N_25233,N_23983,N_24829);
xor U25234 (N_25234,N_24872,N_23958);
nor U25235 (N_25235,N_24974,N_24804);
nor U25236 (N_25236,N_24399,N_24617);
nor U25237 (N_25237,N_22560,N_23461);
nor U25238 (N_25238,N_24932,N_24963);
nand U25239 (N_25239,N_22899,N_23520);
xnor U25240 (N_25240,N_24003,N_24548);
nand U25241 (N_25241,N_23660,N_23369);
nor U25242 (N_25242,N_24532,N_24431);
and U25243 (N_25243,N_23820,N_24164);
xor U25244 (N_25244,N_24552,N_24386);
and U25245 (N_25245,N_24298,N_23978);
xnor U25246 (N_25246,N_23030,N_23942);
xnor U25247 (N_25247,N_23014,N_22962);
nand U25248 (N_25248,N_24291,N_23008);
xor U25249 (N_25249,N_24403,N_23114);
xor U25250 (N_25250,N_24925,N_23683);
nor U25251 (N_25251,N_24826,N_23805);
or U25252 (N_25252,N_23216,N_23640);
xor U25253 (N_25253,N_24671,N_23457);
or U25254 (N_25254,N_22509,N_23102);
nor U25255 (N_25255,N_23269,N_24865);
xnor U25256 (N_25256,N_23490,N_23164);
xor U25257 (N_25257,N_22575,N_23743);
or U25258 (N_25258,N_23903,N_22850);
or U25259 (N_25259,N_23049,N_23599);
or U25260 (N_25260,N_22994,N_23118);
nor U25261 (N_25261,N_22524,N_24195);
nand U25262 (N_25262,N_24314,N_23316);
xnor U25263 (N_25263,N_22757,N_22879);
or U25264 (N_25264,N_24550,N_24420);
nor U25265 (N_25265,N_23277,N_24188);
or U25266 (N_25266,N_22777,N_24911);
or U25267 (N_25267,N_24994,N_23894);
or U25268 (N_25268,N_22572,N_23998);
nand U25269 (N_25269,N_24116,N_24182);
nor U25270 (N_25270,N_22989,N_23366);
xor U25271 (N_25271,N_22939,N_22638);
or U25272 (N_25272,N_24707,N_24286);
nand U25273 (N_25273,N_24516,N_24572);
or U25274 (N_25274,N_23577,N_22927);
nor U25275 (N_25275,N_24030,N_23005);
nor U25276 (N_25276,N_23129,N_24842);
xnor U25277 (N_25277,N_24236,N_24086);
or U25278 (N_25278,N_24628,N_24569);
xor U25279 (N_25279,N_23892,N_22664);
xnor U25280 (N_25280,N_22766,N_24416);
xnor U25281 (N_25281,N_23244,N_24907);
or U25282 (N_25282,N_24690,N_24470);
xnor U25283 (N_25283,N_22547,N_22505);
xnor U25284 (N_25284,N_22656,N_24451);
xor U25285 (N_25285,N_23912,N_24296);
and U25286 (N_25286,N_24814,N_24774);
nand U25287 (N_25287,N_24794,N_24396);
xnor U25288 (N_25288,N_22716,N_22561);
nor U25289 (N_25289,N_23575,N_23552);
nand U25290 (N_25290,N_24277,N_24153);
nor U25291 (N_25291,N_23029,N_23111);
and U25292 (N_25292,N_23036,N_22641);
xor U25293 (N_25293,N_23937,N_24682);
or U25294 (N_25294,N_24007,N_24425);
and U25295 (N_25295,N_23449,N_22644);
nand U25296 (N_25296,N_23047,N_24656);
and U25297 (N_25297,N_23754,N_24160);
xnor U25298 (N_25298,N_23482,N_22562);
nor U25299 (N_25299,N_22941,N_24640);
nand U25300 (N_25300,N_22750,N_22888);
nor U25301 (N_25301,N_22658,N_24010);
or U25302 (N_25302,N_24067,N_24997);
or U25303 (N_25303,N_22867,N_23243);
and U25304 (N_25304,N_23917,N_24032);
or U25305 (N_25305,N_24713,N_23723);
xnor U25306 (N_25306,N_22871,N_22820);
and U25307 (N_25307,N_24174,N_23359);
and U25308 (N_25308,N_23427,N_23238);
or U25309 (N_25309,N_23478,N_24268);
xnor U25310 (N_25310,N_22729,N_24487);
nand U25311 (N_25311,N_23671,N_23064);
or U25312 (N_25312,N_24221,N_24311);
nor U25313 (N_25313,N_24018,N_24358);
nand U25314 (N_25314,N_24676,N_23878);
nor U25315 (N_25315,N_23619,N_23769);
nand U25316 (N_25316,N_24844,N_22773);
and U25317 (N_25317,N_22615,N_24031);
or U25318 (N_25318,N_23240,N_23714);
xnor U25319 (N_25319,N_24285,N_24379);
and U25320 (N_25320,N_22674,N_22712);
nand U25321 (N_25321,N_23727,N_24338);
xnor U25322 (N_25322,N_23441,N_23195);
nor U25323 (N_25323,N_23222,N_24743);
or U25324 (N_25324,N_24822,N_23716);
nand U25325 (N_25325,N_23010,N_23697);
or U25326 (N_25326,N_23571,N_23767);
xnor U25327 (N_25327,N_22673,N_24192);
nor U25328 (N_25328,N_22904,N_22677);
xor U25329 (N_25329,N_23361,N_23909);
nor U25330 (N_25330,N_23132,N_24278);
nand U25331 (N_25331,N_24845,N_24347);
nor U25332 (N_25332,N_22835,N_24782);
xnor U25333 (N_25333,N_23885,N_22807);
and U25334 (N_25334,N_24888,N_23462);
or U25335 (N_25335,N_22912,N_22698);
nand U25336 (N_25336,N_24257,N_23463);
nor U25337 (N_25337,N_23920,N_24802);
and U25338 (N_25338,N_22805,N_23704);
nand U25339 (N_25339,N_23989,N_22759);
xnor U25340 (N_25340,N_23994,N_23753);
and U25341 (N_25341,N_23218,N_23230);
xor U25342 (N_25342,N_24026,N_24280);
nand U25343 (N_25343,N_24721,N_24933);
nor U25344 (N_25344,N_22834,N_22787);
or U25345 (N_25345,N_23389,N_24821);
nor U25346 (N_25346,N_22684,N_22708);
nor U25347 (N_25347,N_23202,N_23328);
or U25348 (N_25348,N_23849,N_24212);
nand U25349 (N_25349,N_24406,N_24672);
or U25350 (N_25350,N_22551,N_24765);
and U25351 (N_25351,N_23211,N_24044);
nor U25352 (N_25352,N_24706,N_22616);
or U25353 (N_25353,N_23060,N_24331);
nand U25354 (N_25354,N_23353,N_24992);
xor U25355 (N_25355,N_22842,N_23384);
and U25356 (N_25356,N_24905,N_24129);
and U25357 (N_25357,N_23875,N_24186);
xor U25358 (N_25358,N_23071,N_23363);
or U25359 (N_25359,N_23289,N_23701);
xor U25360 (N_25360,N_23576,N_24784);
or U25361 (N_25361,N_24279,N_23940);
nor U25362 (N_25362,N_24375,N_23857);
or U25363 (N_25363,N_22686,N_23053);
and U25364 (N_25364,N_24295,N_23262);
nor U25365 (N_25365,N_23665,N_24899);
and U25366 (N_25366,N_24866,N_24716);
nand U25367 (N_25367,N_22650,N_23259);
nand U25368 (N_25368,N_24092,N_22696);
nand U25369 (N_25369,N_23628,N_24162);
or U25370 (N_25370,N_23063,N_24854);
and U25371 (N_25371,N_24579,N_22826);
and U25372 (N_25372,N_24622,N_24679);
nand U25373 (N_25373,N_23266,N_24201);
and U25374 (N_25374,N_23666,N_23263);
and U25375 (N_25375,N_24385,N_24093);
and U25376 (N_25376,N_24341,N_22848);
nand U25377 (N_25377,N_24645,N_23960);
nor U25378 (N_25378,N_22951,N_22977);
xor U25379 (N_25379,N_23988,N_23584);
xor U25380 (N_25380,N_23967,N_23712);
and U25381 (N_25381,N_23929,N_23775);
nor U25382 (N_25382,N_24271,N_23191);
xor U25383 (N_25383,N_23624,N_24024);
or U25384 (N_25384,N_22587,N_22797);
and U25385 (N_25385,N_23247,N_24950);
nor U25386 (N_25386,N_23226,N_24471);
and U25387 (N_25387,N_23608,N_22570);
nor U25388 (N_25388,N_22749,N_23217);
nand U25389 (N_25389,N_23905,N_22881);
and U25390 (N_25390,N_22831,N_22997);
xor U25391 (N_25391,N_23533,N_24282);
or U25392 (N_25392,N_24789,N_22517);
nand U25393 (N_25393,N_22740,N_22909);
nor U25394 (N_25394,N_23413,N_24483);
xnor U25395 (N_25395,N_23434,N_23464);
nor U25396 (N_25396,N_23756,N_24349);
xnor U25397 (N_25397,N_24993,N_24588);
xor U25398 (N_25398,N_23382,N_24662);
and U25399 (N_25399,N_23080,N_22830);
xor U25400 (N_25400,N_23859,N_24434);
and U25401 (N_25401,N_22922,N_23368);
nor U25402 (N_25402,N_24839,N_23167);
xor U25403 (N_25403,N_24796,N_24868);
nand U25404 (N_25404,N_23234,N_23796);
xor U25405 (N_25405,N_22752,N_24462);
and U25406 (N_25406,N_23543,N_24924);
xor U25407 (N_25407,N_24232,N_24515);
nor U25408 (N_25408,N_23257,N_22612);
nor U25409 (N_25409,N_22863,N_23264);
or U25410 (N_25410,N_24903,N_23655);
and U25411 (N_25411,N_23294,N_23523);
or U25412 (N_25412,N_23679,N_23840);
nand U25413 (N_25413,N_22627,N_23419);
or U25414 (N_25414,N_24935,N_24759);
nor U25415 (N_25415,N_23345,N_23653);
or U25416 (N_25416,N_24313,N_24990);
nand U25417 (N_25417,N_24973,N_23831);
xor U25418 (N_25418,N_23955,N_24859);
xnor U25419 (N_25419,N_22703,N_24995);
nor U25420 (N_25420,N_22629,N_23651);
or U25421 (N_25421,N_24202,N_24424);
nand U25422 (N_25422,N_22883,N_22942);
or U25423 (N_25423,N_24037,N_22782);
nor U25424 (N_25424,N_24745,N_23094);
xnor U25425 (N_25425,N_22849,N_23007);
nor U25426 (N_25426,N_23192,N_24480);
or U25427 (N_25427,N_23919,N_22685);
and U25428 (N_25428,N_24976,N_23293);
or U25429 (N_25429,N_24433,N_24079);
or U25430 (N_25430,N_24841,N_23889);
nor U25431 (N_25431,N_23979,N_24808);
nand U25432 (N_25432,N_24078,N_24439);
xor U25433 (N_25433,N_23207,N_23739);
nor U25434 (N_25434,N_22815,N_24971);
and U25435 (N_25435,N_22774,N_22914);
or U25436 (N_25436,N_22514,N_22767);
nor U25437 (N_25437,N_23706,N_22676);
or U25438 (N_25438,N_22675,N_23862);
nand U25439 (N_25439,N_22793,N_24766);
nor U25440 (N_25440,N_23339,N_24922);
nand U25441 (N_25441,N_23846,N_23951);
and U25442 (N_25442,N_23732,N_22860);
nand U25443 (N_25443,N_23051,N_23685);
nor U25444 (N_25444,N_23475,N_24040);
nor U25445 (N_25445,N_23034,N_22670);
xor U25446 (N_25446,N_24340,N_24013);
or U25447 (N_25447,N_23711,N_24580);
or U25448 (N_25448,N_24850,N_22634);
nand U25449 (N_25449,N_23984,N_24583);
nor U25450 (N_25450,N_22965,N_23138);
nor U25451 (N_25451,N_24730,N_23276);
nand U25452 (N_25452,N_22756,N_23344);
or U25453 (N_25453,N_22843,N_23808);
xor U25454 (N_25454,N_23692,N_23500);
nor U25455 (N_25455,N_23439,N_23343);
nor U25456 (N_25456,N_22606,N_24429);
or U25457 (N_25457,N_23828,N_24256);
nor U25458 (N_25458,N_24705,N_23255);
or U25459 (N_25459,N_23232,N_22884);
nor U25460 (N_25460,N_23515,N_23426);
or U25461 (N_25461,N_24633,N_22633);
or U25462 (N_25462,N_24562,N_23510);
nor U25463 (N_25463,N_22810,N_23107);
nor U25464 (N_25464,N_22996,N_23545);
nor U25465 (N_25465,N_23698,N_22919);
nor U25466 (N_25466,N_23976,N_23511);
nand U25467 (N_25467,N_24364,N_23870);
nor U25468 (N_25468,N_24147,N_23474);
nor U25469 (N_25469,N_23959,N_24497);
and U25470 (N_25470,N_24704,N_22796);
and U25471 (N_25471,N_24354,N_24582);
nand U25472 (N_25472,N_23003,N_22917);
or U25473 (N_25473,N_24595,N_22955);
or U25474 (N_25474,N_24938,N_23851);
nor U25475 (N_25475,N_23904,N_24407);
nor U25476 (N_25476,N_23335,N_23249);
or U25477 (N_25477,N_22930,N_22559);
xnor U25478 (N_25478,N_24504,N_23031);
and U25479 (N_25479,N_22553,N_23686);
nor U25480 (N_25480,N_22556,N_23310);
xor U25481 (N_25481,N_23659,N_24952);
and U25482 (N_25482,N_23770,N_23798);
or U25483 (N_25483,N_23076,N_24521);
and U25484 (N_25484,N_24596,N_24964);
nor U25485 (N_25485,N_24333,N_24624);
or U25486 (N_25486,N_23139,N_23325);
nor U25487 (N_25487,N_24890,N_23157);
and U25488 (N_25488,N_23017,N_24968);
and U25489 (N_25489,N_23595,N_23026);
xnor U25490 (N_25490,N_24012,N_24000);
or U25491 (N_25491,N_23657,N_22585);
and U25492 (N_25492,N_24361,N_23179);
nand U25493 (N_25493,N_24412,N_23801);
or U25494 (N_25494,N_23911,N_24818);
xor U25495 (N_25495,N_23321,N_24776);
nand U25496 (N_25496,N_24746,N_23333);
xor U25497 (N_25497,N_23365,N_23378);
xnor U25498 (N_25498,N_24118,N_24217);
and U25499 (N_25499,N_23109,N_23806);
or U25500 (N_25500,N_22502,N_24302);
and U25501 (N_25501,N_24308,N_23267);
and U25502 (N_25502,N_24960,N_23284);
nor U25503 (N_25503,N_24446,N_24500);
nand U25504 (N_25504,N_24414,N_24011);
and U25505 (N_25505,N_24666,N_23700);
nor U25506 (N_25506,N_23578,N_24248);
xor U25507 (N_25507,N_22535,N_23611);
or U25508 (N_25508,N_23522,N_23987);
xor U25509 (N_25509,N_24540,N_24761);
xor U25510 (N_25510,N_23772,N_23633);
or U25511 (N_25511,N_23220,N_24958);
nor U25512 (N_25512,N_22730,N_24653);
nor U25513 (N_25513,N_23546,N_23881);
nand U25514 (N_25514,N_23676,N_23357);
and U25515 (N_25515,N_24063,N_24443);
xnor U25516 (N_25516,N_23253,N_23923);
nand U25517 (N_25517,N_22795,N_23513);
nand U25518 (N_25518,N_24360,N_24342);
or U25519 (N_25519,N_24665,N_24638);
xor U25520 (N_25520,N_23544,N_23572);
xor U25521 (N_25521,N_22967,N_23819);
nor U25522 (N_25522,N_24072,N_22907);
xor U25523 (N_25523,N_24880,N_23181);
nand U25524 (N_25524,N_24365,N_23352);
nor U25525 (N_25525,N_24134,N_23033);
or U25526 (N_25526,N_23748,N_23151);
xnor U25527 (N_25527,N_23879,N_22577);
or U25528 (N_25528,N_24737,N_23497);
nand U25529 (N_25529,N_22525,N_23688);
xor U25530 (N_25530,N_24531,N_22924);
nand U25531 (N_25531,N_23021,N_24539);
or U25532 (N_25532,N_24912,N_22655);
and U25533 (N_25533,N_23807,N_23961);
and U25534 (N_25534,N_22589,N_23205);
and U25535 (N_25535,N_23163,N_24897);
and U25536 (N_25536,N_22571,N_23396);
or U25537 (N_25537,N_23091,N_24098);
or U25538 (N_25538,N_24445,N_24215);
or U25539 (N_25539,N_24876,N_24695);
and U25540 (N_25540,N_23501,N_23759);
nor U25541 (N_25541,N_23286,N_24862);
nand U25542 (N_25542,N_22503,N_23972);
nor U25543 (N_25543,N_22568,N_23965);
or U25544 (N_25544,N_24169,N_22546);
nor U25545 (N_25545,N_22806,N_24476);
nand U25546 (N_25546,N_23928,N_23563);
or U25547 (N_25547,N_24718,N_23720);
and U25548 (N_25548,N_24076,N_23612);
and U25549 (N_25549,N_23592,N_22803);
and U25550 (N_25550,N_22719,N_22692);
nor U25551 (N_25551,N_22564,N_23598);
xor U25552 (N_25552,N_23499,N_23043);
xnor U25553 (N_25553,N_23673,N_24612);
and U25554 (N_25554,N_23850,N_23643);
nand U25555 (N_25555,N_24353,N_24332);
and U25556 (N_25556,N_22822,N_24554);
nand U25557 (N_25557,N_22590,N_23966);
or U25558 (N_25558,N_23044,N_24411);
nand U25559 (N_25559,N_24848,N_22839);
or U25560 (N_25560,N_24722,N_24249);
xor U25561 (N_25561,N_24832,N_23123);
and U25562 (N_25562,N_24755,N_22833);
nand U25563 (N_25563,N_23058,N_24538);
and U25564 (N_25564,N_22682,N_23466);
nand U25565 (N_25565,N_23038,N_24227);
xnor U25566 (N_25566,N_24346,N_24301);
nand U25567 (N_25567,N_22538,N_22631);
or U25568 (N_25568,N_24783,N_23678);
or U25569 (N_25569,N_23771,N_24329);
nand U25570 (N_25570,N_22970,N_24189);
or U25571 (N_25571,N_23487,N_24173);
xnor U25572 (N_25572,N_24209,N_24352);
xor U25573 (N_25573,N_24535,N_24144);
or U25574 (N_25574,N_23789,N_24565);
xnor U25575 (N_25575,N_24657,N_23606);
or U25576 (N_25576,N_24131,N_22973);
xor U25577 (N_25577,N_24288,N_23314);
or U25578 (N_25578,N_24887,N_22814);
nand U25579 (N_25579,N_24490,N_23934);
nor U25580 (N_25580,N_22920,N_22647);
and U25581 (N_25581,N_24152,N_22521);
xnor U25582 (N_25582,N_22772,N_23990);
or U25583 (N_25583,N_23625,N_22993);
nor U25584 (N_25584,N_24937,N_24336);
or U25585 (N_25585,N_23601,N_23301);
or U25586 (N_25586,N_22552,N_24405);
nand U25587 (N_25587,N_22733,N_24191);
nor U25588 (N_25588,N_24442,N_23634);
nand U25589 (N_25589,N_24294,N_23596);
xor U25590 (N_25590,N_24213,N_23969);
or U25591 (N_25591,N_23933,N_24757);
nand U25592 (N_25592,N_22578,N_24736);
xnor U25593 (N_25593,N_23908,N_22574);
and U25594 (N_25594,N_22602,N_24693);
xnor U25595 (N_25595,N_24664,N_24395);
and U25596 (N_25596,N_24075,N_23093);
xnor U25597 (N_25597,N_24253,N_23827);
nand U25598 (N_25598,N_22542,N_24474);
xnor U25599 (N_25599,N_23669,N_24488);
and U25600 (N_25600,N_23664,N_22697);
xor U25601 (N_25601,N_23392,N_24762);
nor U25602 (N_25602,N_23183,N_24083);
nand U25603 (N_25603,N_24940,N_24574);
nor U25604 (N_25604,N_22758,N_24070);
nor U25605 (N_25605,N_22679,N_22743);
or U25606 (N_25606,N_24316,N_22934);
or U25607 (N_25607,N_24764,N_24196);
and U25608 (N_25608,N_23112,N_23586);
and U25609 (N_25609,N_23142,N_24610);
nor U25610 (N_25610,N_24851,N_24001);
and U25611 (N_25611,N_23512,N_24727);
nand U25612 (N_25612,N_24069,N_24647);
nand U25613 (N_25613,N_22548,N_24351);
nand U25614 (N_25614,N_24593,N_24111);
and U25615 (N_25615,N_23408,N_24481);
and U25616 (N_25616,N_24557,N_24510);
or U25617 (N_25617,N_23428,N_23156);
and U25618 (N_25618,N_23537,N_23274);
nor U25619 (N_25619,N_23731,N_22770);
nor U25620 (N_25620,N_24413,N_24947);
nor U25621 (N_25621,N_24472,N_24051);
xor U25622 (N_25622,N_22711,N_24629);
xor U25623 (N_25623,N_23896,N_23445);
and U25624 (N_25624,N_23914,N_23086);
nor U25625 (N_25625,N_23312,N_23558);
or U25626 (N_25626,N_23555,N_23681);
nor U25627 (N_25627,N_23134,N_23786);
or U25628 (N_25628,N_24023,N_22721);
and U25629 (N_25629,N_24780,N_24095);
nor U25630 (N_25630,N_23550,N_24485);
or U25631 (N_25631,N_23504,N_23214);
or U25632 (N_25632,N_24505,N_24601);
or U25633 (N_25633,N_24942,N_22877);
xnor U25634 (N_25634,N_24526,N_24120);
nand U25635 (N_25635,N_22508,N_23607);
and U25636 (N_25636,N_24495,N_24315);
xnor U25637 (N_25637,N_23663,N_23390);
or U25638 (N_25638,N_24828,N_22691);
nand U25639 (N_25639,N_24983,N_22714);
or U25640 (N_25640,N_22923,N_24100);
or U25641 (N_25641,N_23061,N_24464);
xnor U25642 (N_25642,N_22958,N_24436);
nand U25643 (N_25643,N_23140,N_23525);
and U25644 (N_25644,N_24909,N_24348);
and U25645 (N_25645,N_23646,N_23417);
or U25646 (N_25646,N_24320,N_24357);
or U25647 (N_25647,N_23535,N_24183);
nand U25648 (N_25648,N_24585,N_23376);
nand U25649 (N_25649,N_23347,N_23647);
nor U25650 (N_25650,N_23573,N_24791);
xor U25651 (N_25651,N_23208,N_23362);
nor U25652 (N_25652,N_22710,N_24231);
nand U25653 (N_25653,N_24725,N_24849);
and U25654 (N_25654,N_23579,N_23925);
xor U25655 (N_25655,N_23999,N_24630);
nand U25656 (N_25656,N_23804,N_22901);
nand U25657 (N_25657,N_23350,N_24795);
and U25658 (N_25658,N_23551,N_23932);
or U25659 (N_25659,N_22983,N_22895);
xor U25660 (N_25660,N_23144,N_24059);
nand U25661 (N_25661,N_24224,N_23691);
and U25662 (N_25662,N_24986,N_22704);
nand U25663 (N_25663,N_23715,N_23631);
nand U25664 (N_25664,N_23054,N_23388);
and U25665 (N_25665,N_23458,N_24167);
and U25666 (N_25666,N_23843,N_23075);
nand U25667 (N_25667,N_24303,N_22829);
and U25668 (N_25668,N_23153,N_22727);
xor U25669 (N_25669,N_23225,N_23854);
xor U25670 (N_25670,N_24606,N_23591);
xor U25671 (N_25671,N_23346,N_23106);
nand U25672 (N_25672,N_22853,N_22801);
or U25673 (N_25673,N_24482,N_24807);
nor U25674 (N_25674,N_22975,N_23638);
nand U25675 (N_25675,N_22800,N_22876);
nor U25676 (N_25676,N_22897,N_24097);
nand U25677 (N_25677,N_24478,N_23184);
nand U25678 (N_25678,N_22990,N_24139);
nand U25679 (N_25679,N_24856,N_24388);
and U25680 (N_25680,N_24955,N_22522);
or U25681 (N_25681,N_24714,N_24035);
nor U25682 (N_25682,N_23371,N_23126);
or U25683 (N_25683,N_24636,N_22588);
nand U25684 (N_25684,N_23165,N_24803);
nor U25685 (N_25685,N_24878,N_24957);
or U25686 (N_25686,N_24117,N_23025);
xnor U25687 (N_25687,N_23340,N_23997);
nor U25688 (N_25688,N_22663,N_23423);
nand U25689 (N_25689,N_24096,N_24409);
nor U25690 (N_25690,N_23186,N_22671);
and U25691 (N_25691,N_23072,N_23489);
xor U25692 (N_25692,N_24071,N_22667);
nor U25693 (N_25693,N_23783,N_23568);
nor U25694 (N_25694,N_23170,N_24769);
and U25695 (N_25695,N_22678,N_23019);
xor U25696 (N_25696,N_24326,N_23108);
xnor U25697 (N_25697,N_24494,N_24673);
nand U25698 (N_25698,N_23538,N_24194);
nand U25699 (N_25699,N_22725,N_22804);
or U25700 (N_25700,N_23130,N_23939);
or U25701 (N_25701,N_23341,N_24127);
or U25702 (N_25702,N_24881,N_22555);
and U25703 (N_25703,N_23503,N_24469);
nand U25704 (N_25704,N_24325,N_24547);
nor U25705 (N_25705,N_23231,N_23309);
xor U25706 (N_25706,N_23667,N_24094);
xor U25707 (N_25707,N_22582,N_23201);
xnor U25708 (N_25708,N_23781,N_24050);
xor U25709 (N_25709,N_22573,N_24669);
xnor U25710 (N_25710,N_22544,N_22510);
nor U25711 (N_25711,N_24747,N_23065);
and U25712 (N_25712,N_24571,N_24819);
and U25713 (N_25713,N_24985,N_22746);
nor U25714 (N_25714,N_23288,N_24467);
and U25715 (N_25715,N_24945,N_22906);
nor U25716 (N_25716,N_24724,N_24879);
xnor U25717 (N_25717,N_24863,N_23864);
nand U25718 (N_25718,N_23099,N_23684);
xor U25719 (N_25719,N_23381,N_22507);
and U25720 (N_25720,N_24943,N_23326);
nand U25721 (N_25721,N_24428,N_23616);
xnor U25722 (N_25722,N_22868,N_24345);
nor U25723 (N_25723,N_22558,N_23066);
or U25724 (N_25724,N_23699,N_24074);
nand U25725 (N_25725,N_24457,N_24667);
nand U25726 (N_25726,N_24322,N_24929);
nor U25727 (N_25727,N_22614,N_24563);
nand U25728 (N_25728,N_23809,N_24970);
nand U25729 (N_25729,N_24644,N_23954);
nand U25730 (N_25730,N_23169,N_23562);
or U25731 (N_25731,N_23935,N_23564);
and U25732 (N_25732,N_23872,N_24377);
and U25733 (N_25733,N_24800,N_23871);
nand U25734 (N_25734,N_23986,N_22529);
or U25735 (N_25735,N_24892,N_22504);
nor U25736 (N_25736,N_23260,N_22511);
or U25737 (N_25737,N_23841,N_24577);
nor U25738 (N_25738,N_24216,N_24512);
nor U25739 (N_25739,N_24696,N_22765);
or U25740 (N_25740,N_23788,N_24853);
nand U25741 (N_25741,N_23194,N_24597);
nand U25742 (N_25742,N_23135,N_24068);
nand U25743 (N_25743,N_24978,N_23121);
nor U25744 (N_25744,N_24002,N_24889);
nor U25745 (N_25745,N_23443,N_24966);
nand U25746 (N_25746,N_24896,N_24229);
or U25747 (N_25747,N_24057,N_24272);
xnor U25748 (N_25748,N_22742,N_22660);
and U25749 (N_25749,N_24218,N_24090);
nand U25750 (N_25750,N_22755,N_24401);
xor U25751 (N_25751,N_22784,N_22693);
or U25752 (N_25752,N_23531,N_23483);
or U25753 (N_25753,N_23780,N_24522);
and U25754 (N_25754,N_22832,N_24545);
and U25755 (N_25755,N_23587,N_23834);
xor U25756 (N_25756,N_24750,N_24087);
or U25757 (N_25757,N_24991,N_22902);
xnor U25758 (N_25758,N_23332,N_23473);
or U25759 (N_25759,N_23479,N_23411);
and U25760 (N_25760,N_24166,N_24728);
xor U25761 (N_25761,N_24533,N_23237);
or U25762 (N_25762,N_24168,N_24857);
or U25763 (N_25763,N_23811,N_24041);
nor U25764 (N_25764,N_24430,N_22918);
nor U25765 (N_25765,N_24620,N_24681);
and U25766 (N_25766,N_24143,N_23492);
nand U25767 (N_25767,N_23948,N_23412);
and U25768 (N_25768,N_22601,N_23735);
and U25769 (N_25769,N_22864,N_23162);
or U25770 (N_25770,N_23415,N_24549);
nor U25771 (N_25771,N_23407,N_23778);
nor U25772 (N_25772,N_24362,N_22780);
and U25773 (N_25773,N_22528,N_23604);
xor U25774 (N_25774,N_22813,N_24877);
xnor U25775 (N_25775,N_23757,N_24176);
or U25776 (N_25776,N_24239,N_24551);
or U25777 (N_25777,N_22713,N_22683);
nand U25778 (N_25778,N_22960,N_22513);
and U25779 (N_25779,N_22954,N_23283);
nor U25780 (N_25780,N_24121,N_24251);
nor U25781 (N_25781,N_22847,N_24758);
nor U25782 (N_25782,N_22783,N_23553);
nand U25783 (N_25783,N_24046,N_23975);
and U25784 (N_25784,N_22600,N_23518);
nand U25785 (N_25785,N_22622,N_23791);
or U25786 (N_25786,N_24165,N_24498);
or U25787 (N_25787,N_22886,N_24243);
xnor U25788 (N_25788,N_24207,N_24148);
xnor U25789 (N_25789,N_24626,N_23465);
or U25790 (N_25790,N_24698,N_23866);
nand U25791 (N_25791,N_22549,N_24381);
nand U25792 (N_25792,N_24276,N_23187);
nand U25793 (N_25793,N_23096,N_23708);
and U25794 (N_25794,N_23224,N_24408);
and U25795 (N_25795,N_22717,N_23009);
nor U25796 (N_25796,N_24107,N_24187);
or U25797 (N_25797,N_23406,N_23242);
or U25798 (N_25798,N_24969,N_23016);
nor U25799 (N_25799,N_24514,N_23090);
and U25800 (N_25800,N_23450,N_24269);
and U25801 (N_25801,N_22964,N_24369);
and U25802 (N_25802,N_23833,N_23768);
or U25803 (N_25803,N_22968,N_23874);
xnor U25804 (N_25804,N_22651,N_24006);
nor U25805 (N_25805,N_23250,N_24586);
and U25806 (N_25806,N_24297,N_23168);
nor U25807 (N_25807,N_22581,N_23223);
and U25808 (N_25808,N_24149,N_22827);
or U25809 (N_25809,N_24267,N_22618);
xnor U25810 (N_25810,N_24591,N_22980);
or U25811 (N_25811,N_22536,N_22739);
or U25812 (N_25812,N_22966,N_23594);
nor U25813 (N_25813,N_22709,N_23635);
xor U25814 (N_25814,N_24184,N_22690);
and U25815 (N_25815,N_22636,N_24754);
nand U25816 (N_25816,N_24109,N_24370);
and U25817 (N_25817,N_24650,N_23295);
or U25818 (N_25818,N_23821,N_23946);
and U25819 (N_25819,N_23814,N_24613);
nor U25820 (N_25820,N_24895,N_23070);
or U25821 (N_25821,N_23401,N_24873);
nand U25822 (N_25822,N_24114,N_22635);
xnor U25823 (N_25823,N_24786,N_23817);
and U25824 (N_25824,N_23869,N_23395);
or U25825 (N_25825,N_23530,N_24125);
xnor U25826 (N_25826,N_23842,N_24817);
xnor U25827 (N_25827,N_24729,N_24923);
xor U25828 (N_25828,N_24197,N_22620);
nor U25829 (N_25829,N_22836,N_22816);
nand U25830 (N_25830,N_22565,N_24208);
and U25831 (N_25831,N_24261,N_23098);
and U25832 (N_25832,N_24274,N_23055);
nor U25833 (N_25833,N_23052,N_23210);
and U25834 (N_25834,N_24901,N_22506);
and U25835 (N_25835,N_24835,N_22594);
xor U25836 (N_25836,N_23486,N_23762);
xor U25837 (N_25837,N_24140,N_23035);
nor U25838 (N_25838,N_23995,N_24344);
xnor U25839 (N_25839,N_24371,N_23810);
and U25840 (N_25840,N_22632,N_24717);
nor U25841 (N_25841,N_24735,N_24508);
and U25842 (N_25842,N_23944,N_24523);
nor U25843 (N_25843,N_23630,N_23204);
nor U25844 (N_25844,N_23469,N_22526);
and U25845 (N_25845,N_23620,N_23839);
or U25846 (N_25846,N_24760,N_24270);
xnor U25847 (N_25847,N_24214,N_23613);
and U25848 (N_25848,N_24447,N_22720);
nand U25849 (N_25849,N_24749,N_23882);
xor U25850 (N_25850,N_23040,N_22788);
xor U25851 (N_25851,N_24205,N_23484);
xnor U25852 (N_25852,N_22985,N_22776);
nand U25853 (N_25853,N_23815,N_24869);
nor U25854 (N_25854,N_24418,N_23331);
xor U25855 (N_25855,N_24948,N_23161);
or U25856 (N_25856,N_24038,N_23193);
nor U25857 (N_25857,N_23292,N_23329);
nor U25858 (N_25858,N_24643,N_22802);
and U25859 (N_25859,N_22986,N_24984);
xnor U25860 (N_25860,N_24812,N_23835);
xnor U25861 (N_25861,N_24708,N_24350);
xor U25862 (N_25862,N_23398,N_23281);
nand U25863 (N_25863,N_22532,N_24493);
or U25864 (N_25864,N_23185,N_24179);
xor U25865 (N_25865,N_23323,N_24719);
xnor U25866 (N_25866,N_24228,N_23435);
nand U25867 (N_25867,N_24867,N_24181);
nand U25868 (N_25868,N_22961,N_24374);
nor U25869 (N_25869,N_23856,N_24809);
nor U25870 (N_25870,N_22523,N_23707);
nand U25871 (N_25871,N_24142,N_23981);
or U25872 (N_25872,N_24170,N_23324);
or U25873 (N_25873,N_23836,N_24137);
nand U25874 (N_25874,N_23087,N_22603);
nand U25875 (N_25875,N_24916,N_23832);
nor U25876 (N_25876,N_23991,N_22837);
nand U25877 (N_25877,N_23372,N_23470);
xnor U25878 (N_25878,N_23861,N_23004);
nand U25879 (N_25879,N_24115,N_23393);
xnor U25880 (N_25880,N_24477,N_23101);
or U25881 (N_25881,N_22869,N_22896);
nand U25882 (N_25882,N_24655,N_23494);
nand U25883 (N_25883,N_24237,N_22607);
nor U25884 (N_25884,N_23580,N_23046);
nand U25885 (N_25885,N_23436,N_22979);
xor U25886 (N_25886,N_24621,N_22798);
nor U25887 (N_25887,N_24126,N_22781);
and U25888 (N_25888,N_24723,N_22949);
nor U25889 (N_25889,N_24544,N_23206);
nor U25890 (N_25890,N_23083,N_24790);
nor U25891 (N_25891,N_24861,N_24771);
nor U25892 (N_25892,N_24608,N_24419);
nor U25893 (N_25893,N_23078,N_24138);
nor U25894 (N_25894,N_24967,N_24744);
xnor U25895 (N_25895,N_23002,N_22921);
xor U25896 (N_25896,N_23173,N_23155);
xor U25897 (N_25897,N_23045,N_23784);
nand U25898 (N_25898,N_23615,N_23645);
or U25899 (N_25899,N_23974,N_22779);
xnor U25900 (N_25900,N_24830,N_22628);
and U25901 (N_25901,N_23012,N_24570);
and U25902 (N_25902,N_23719,N_24977);
or U25903 (N_25903,N_24886,N_22539);
nand U25904 (N_25904,N_23641,N_23493);
xnor U25905 (N_25905,N_24537,N_23709);
and U25906 (N_25906,N_23658,N_23588);
nor U25907 (N_25907,N_23145,N_23795);
and U25908 (N_25908,N_24846,N_23670);
nand U25909 (N_25909,N_23521,N_22648);
xnor U25910 (N_25910,N_23280,N_23304);
or U25911 (N_25911,N_22540,N_22768);
nor U25912 (N_25912,N_23873,N_22604);
nor U25913 (N_25913,N_22724,N_23913);
xnor U25914 (N_25914,N_24404,N_23565);
nor U25915 (N_25915,N_24703,N_22873);
nor U25916 (N_25916,N_24450,N_24265);
nand U25917 (N_25917,N_22543,N_24034);
nor U25918 (N_25918,N_24058,N_24290);
nor U25919 (N_25919,N_22694,N_24312);
nand U25920 (N_25920,N_24200,N_24452);
or U25921 (N_25921,N_23787,N_23696);
nand U25922 (N_25922,N_24465,N_24392);
nand U25923 (N_25923,N_23561,N_22723);
nand U25924 (N_25924,N_24368,N_23330);
nand U25925 (N_25925,N_23812,N_24402);
nand U25926 (N_25926,N_24893,N_23085);
and U25927 (N_25927,N_23236,N_24080);
and U25928 (N_25928,N_22851,N_24536);
nor U25929 (N_25929,N_24517,N_23104);
or U25930 (N_25930,N_24390,N_22910);
nor U25931 (N_25931,N_23938,N_23803);
or U25932 (N_25932,N_24979,N_22550);
nor U25933 (N_25933,N_22597,N_22925);
nand U25934 (N_25934,N_24611,N_23705);
nand U25935 (N_25935,N_24009,N_23338);
or U25936 (N_25936,N_23298,N_23853);
xnor U25937 (N_25937,N_24047,N_22999);
or U25938 (N_25938,N_23830,N_22946);
nor U25939 (N_25939,N_24827,N_24324);
xor U25940 (N_25940,N_23050,N_22799);
nor U25941 (N_25941,N_24101,N_22681);
nor U25942 (N_25942,N_24838,N_23197);
xnor U25943 (N_25943,N_23103,N_23985);
or U25944 (N_25944,N_23410,N_22875);
nor U25945 (N_25945,N_23215,N_22659);
and U25946 (N_25946,N_22662,N_22726);
nand U25947 (N_25947,N_22745,N_23068);
xor U25948 (N_25948,N_23733,N_24631);
xor U25949 (N_25949,N_23180,N_24128);
xnor U25950 (N_25950,N_23446,N_24941);
nor U25951 (N_25951,N_22688,N_23717);
or U25952 (N_25952,N_24263,N_24105);
nand U25953 (N_25953,N_23422,N_23380);
xnor U25954 (N_25954,N_24234,N_23498);
or U25955 (N_25955,N_24641,N_23027);
nand U25956 (N_25956,N_23802,N_23848);
and U25957 (N_25957,N_24219,N_23822);
xnor U25958 (N_25958,N_23924,N_24145);
nand U25959 (N_25959,N_23519,N_24022);
xor U25960 (N_25960,N_22935,N_23175);
and U25961 (N_25961,N_23273,N_23947);
or U25962 (N_25962,N_24875,N_23403);
and U25963 (N_25963,N_23404,N_22882);
xnor U25964 (N_25964,N_24711,N_24052);
xor U25965 (N_25965,N_23416,N_24091);
nor U25966 (N_25966,N_22753,N_24604);
and U25967 (N_25967,N_23227,N_23092);
xor U25968 (N_25968,N_24616,N_23602);
and U25969 (N_25969,N_24677,N_23200);
nor U25970 (N_25970,N_22567,N_22878);
xnor U25971 (N_25971,N_22794,N_22584);
or U25972 (N_25972,N_24250,N_24953);
nand U25973 (N_25973,N_24339,N_22512);
nand U25974 (N_25974,N_23115,N_24028);
and U25975 (N_25975,N_23334,N_24573);
nor U25976 (N_25976,N_24178,N_24797);
or U25977 (N_25977,N_23120,N_23127);
nor U25978 (N_25978,N_22613,N_22731);
or U25979 (N_25979,N_24061,N_23597);
nand U25980 (N_25980,N_22790,N_23015);
or U25981 (N_25981,N_24463,N_23270);
nand U25982 (N_25982,N_24437,N_23481);
or U25983 (N_25983,N_22705,N_24356);
nor U25984 (N_25984,N_23774,N_23922);
nand U25985 (N_25985,N_23930,N_22695);
or U25986 (N_25986,N_23931,N_24678);
xnor U25987 (N_25987,N_24788,N_24732);
xnor U25988 (N_25988,N_23182,N_24359);
and U25989 (N_25989,N_23890,N_24225);
or U25990 (N_25990,N_22718,N_24389);
or U25991 (N_25991,N_23898,N_24323);
and U25992 (N_25992,N_23278,N_22786);
and U25993 (N_25993,N_22984,N_24823);
xor U25994 (N_25994,N_23477,N_22501);
xor U25995 (N_25995,N_23258,N_23528);
and U25996 (N_25996,N_23980,N_24815);
xor U25997 (N_25997,N_24529,N_24598);
or U25998 (N_25998,N_23150,N_22859);
nand U25999 (N_25999,N_23391,N_23488);
nand U26000 (N_26000,N_23147,N_24697);
xnor U26001 (N_26001,N_23468,N_24999);
xnor U26002 (N_26002,N_24742,N_23069);
or U26003 (N_26003,N_23146,N_24734);
or U26004 (N_26004,N_23943,N_24479);
nand U26005 (N_26005,N_24685,N_24235);
nand U26006 (N_26006,N_23420,N_24175);
nand U26007 (N_26007,N_24366,N_24085);
or U26008 (N_26008,N_24382,N_24441);
and U26009 (N_26009,N_22969,N_22861);
nand U26010 (N_26010,N_22928,N_24203);
and U26011 (N_26011,N_23763,N_23605);
and U26012 (N_26012,N_23438,N_22702);
nor U26013 (N_26013,N_24556,N_24486);
and U26014 (N_26014,N_23360,N_24642);
or U26015 (N_26015,N_23125,N_24373);
or U26016 (N_26016,N_23755,N_22892);
xor U26017 (N_26017,N_23079,N_24240);
nand U26018 (N_26018,N_24607,N_24309);
nor U26019 (N_26019,N_23177,N_24663);
and U26020 (N_26020,N_24564,N_23622);
nor U26021 (N_26021,N_24609,N_22657);
and U26022 (N_26022,N_23212,N_24054);
xor U26023 (N_26023,N_23549,N_22609);
xnor U26024 (N_26024,N_23261,N_24258);
nor U26025 (N_26025,N_23041,N_24560);
nor U26026 (N_26026,N_22516,N_24770);
nand U26027 (N_26027,N_24155,N_23315);
and U26028 (N_26028,N_24779,N_22808);
or U26029 (N_26029,N_22610,N_22974);
or U26030 (N_26030,N_23800,N_24928);
nor U26031 (N_26031,N_23171,N_24084);
nor U26032 (N_26032,N_23825,N_24135);
or U26033 (N_26033,N_24680,N_23728);
or U26034 (N_26034,N_24987,N_24926);
nor U26035 (N_26035,N_23621,N_24158);
or U26036 (N_26036,N_23863,N_23818);
and U26037 (N_26037,N_24210,N_22624);
nor U26038 (N_26038,N_23229,N_22957);
nand U26039 (N_26039,N_22913,N_23342);
xor U26040 (N_26040,N_23221,N_23527);
and U26041 (N_26041,N_24151,N_24064);
or U26042 (N_26042,N_23617,N_23529);
nor U26043 (N_26043,N_22762,N_23516);
and U26044 (N_26044,N_24159,N_23001);
nand U26045 (N_26045,N_23895,N_23901);
nor U26046 (N_26046,N_23816,N_22971);
xor U26047 (N_26047,N_23448,N_22706);
or U26048 (N_26048,N_23440,N_23792);
nor U26049 (N_26049,N_22819,N_23311);
or U26050 (N_26050,N_23447,N_24112);
or U26051 (N_26051,N_24949,N_24951);
xor U26052 (N_26052,N_23682,N_23581);
nor U26053 (N_26053,N_22866,N_23097);
nand U26054 (N_26054,N_22541,N_24099);
or U26055 (N_26055,N_23689,N_24017);
nor U26056 (N_26056,N_23067,N_23241);
xor U26057 (N_26057,N_23637,N_23131);
nand U26058 (N_26058,N_24773,N_24635);
nand U26059 (N_26059,N_24220,N_22900);
or U26060 (N_26060,N_24367,N_22592);
nand U26061 (N_26061,N_24741,N_23785);
and U26062 (N_26062,N_24489,N_23603);
nand U26063 (N_26063,N_23048,N_23548);
nor U26064 (N_26064,N_22515,N_24767);
and U26065 (N_26065,N_22950,N_24496);
nand U26066 (N_26066,N_23190,N_24541);
nor U26067 (N_26067,N_24410,N_24686);
nor U26068 (N_26068,N_24304,N_24836);
nor U26069 (N_26069,N_24553,N_23496);
or U26070 (N_26070,N_24506,N_24965);
nand U26071 (N_26071,N_24029,N_23764);
and U26072 (N_26072,N_23900,N_24394);
or U26073 (N_26073,N_23113,N_24511);
xnor U26074 (N_26074,N_22579,N_23082);
or U26075 (N_26075,N_24193,N_23290);
xnor U26076 (N_26076,N_22963,N_22911);
nor U26077 (N_26077,N_22840,N_24989);
or U26078 (N_26078,N_24908,N_24587);
nand U26079 (N_26079,N_23354,N_24581);
nor U26080 (N_26080,N_23057,N_24874);
or U26081 (N_26081,N_23729,N_23982);
nor U26082 (N_26082,N_24831,N_23884);
nor U26083 (N_26083,N_23452,N_23110);
and U26084 (N_26084,N_24383,N_22948);
or U26085 (N_26085,N_24154,N_24637);
nor U26086 (N_26086,N_23265,N_22811);
nand U26087 (N_26087,N_24834,N_24931);
xor U26088 (N_26088,N_24775,N_23534);
xnor U26089 (N_26089,N_24119,N_24327);
and U26090 (N_26090,N_24266,N_24605);
nand U26091 (N_26091,N_24398,N_23133);
or U26092 (N_26092,N_23308,N_23444);
nand U26093 (N_26093,N_22707,N_23927);
nor U26094 (N_26094,N_23291,N_24021);
or U26095 (N_26095,N_24104,N_23627);
xnor U26096 (N_26096,N_22741,N_24709);
xor U26097 (N_26097,N_23921,N_22858);
and U26098 (N_26098,N_22791,N_24146);
nand U26099 (N_26099,N_23585,N_24810);
nand U26100 (N_26100,N_23517,N_23213);
and U26101 (N_26101,N_24334,N_23188);
or U26102 (N_26102,N_24049,N_22846);
nand U26103 (N_26103,N_24906,N_23793);
and U26104 (N_26104,N_23876,N_24254);
nor U26105 (N_26105,N_22764,N_24840);
and U26106 (N_26106,N_24330,N_24648);
or U26107 (N_26107,N_23042,N_23855);
nand U26108 (N_26108,N_24198,N_22908);
and U26109 (N_26109,N_23672,N_24649);
or U26110 (N_26110,N_23296,N_24287);
nand U26111 (N_26111,N_23945,N_23725);
nand U26112 (N_26112,N_23137,N_22792);
and U26113 (N_26113,N_24293,N_24632);
and U26114 (N_26114,N_22929,N_24088);
and U26115 (N_26115,N_22534,N_24871);
xnor U26116 (N_26116,N_22972,N_22844);
nor U26117 (N_26117,N_22885,N_23317);
or U26118 (N_26118,N_24688,N_23509);
nand U26119 (N_26119,N_23405,N_23022);
nor U26120 (N_26120,N_24016,N_24720);
xnor U26121 (N_26121,N_22778,N_24066);
nand U26122 (N_26122,N_23418,N_23926);
xor U26123 (N_26123,N_22893,N_24615);
nand U26124 (N_26124,N_23209,N_23560);
and U26125 (N_26125,N_24422,N_24432);
xnor U26126 (N_26126,N_23219,N_23399);
nor U26127 (N_26127,N_23687,N_23373);
and U26128 (N_26128,N_24503,N_24252);
and U26129 (N_26129,N_24816,N_22891);
xnor U26130 (N_26130,N_22998,N_23198);
nand U26131 (N_26131,N_24156,N_23740);
or U26132 (N_26132,N_23506,N_22576);
nand U26133 (N_26133,N_22903,N_23400);
xor U26134 (N_26134,N_24894,N_24283);
and U26135 (N_26135,N_22654,N_24847);
nand U26136 (N_26136,N_24568,N_22944);
and U26137 (N_26137,N_22862,N_23583);
or U26138 (N_26138,N_23675,N_24108);
nand U26139 (N_26139,N_24073,N_24281);
xor U26140 (N_26140,N_24355,N_23394);
nor U26141 (N_26141,N_23303,N_23252);
or U26142 (N_26142,N_23074,N_24692);
or U26143 (N_26143,N_24772,N_24384);
or U26144 (N_26144,N_24036,N_23502);
and U26145 (N_26145,N_23228,N_24292);
or U26146 (N_26146,N_23430,N_24391);
nand U26147 (N_26147,N_24423,N_23642);
nor U26148 (N_26148,N_22625,N_23275);
and U26149 (N_26149,N_23674,N_24910);
nand U26150 (N_26150,N_24172,N_24659);
xor U26151 (N_26151,N_24255,N_24318);
nor U26152 (N_26152,N_23724,N_24785);
and U26153 (N_26153,N_23695,N_23056);
nand U26154 (N_26154,N_23918,N_23765);
and U26155 (N_26155,N_23949,N_22988);
nor U26156 (N_26156,N_22915,N_23084);
xnor U26157 (N_26157,N_24980,N_22728);
nand U26158 (N_26158,N_23011,N_23886);
and U26159 (N_26159,N_22821,N_23287);
xor U26160 (N_26160,N_23128,N_24300);
xnor U26161 (N_26161,N_23032,N_22700);
and U26162 (N_26162,N_24837,N_24524);
nor U26163 (N_26163,N_24988,N_24223);
nand U26164 (N_26164,N_24019,N_24687);
or U26165 (N_26165,N_24042,N_23239);
xnor U26166 (N_26166,N_24799,N_24206);
or U26167 (N_26167,N_24264,N_24934);
xor U26168 (N_26168,N_23973,N_23460);
or U26169 (N_26169,N_24684,N_22580);
nand U26170 (N_26170,N_24982,N_23847);
and U26171 (N_26171,N_24273,N_22936);
and U26172 (N_26172,N_24417,N_23402);
nand U26173 (N_26173,N_24870,N_23971);
xor U26174 (N_26174,N_24289,N_23302);
nor U26175 (N_26175,N_23858,N_24555);
and U26176 (N_26176,N_24103,N_23013);
or U26177 (N_26177,N_24902,N_24230);
or U26178 (N_26178,N_24262,N_23437);
nor U26179 (N_26179,N_23081,N_23387);
nand U26180 (N_26180,N_23507,N_23758);
xor U26181 (N_26181,N_24700,N_24113);
nand U26182 (N_26182,N_23844,N_24180);
or U26183 (N_26183,N_23189,N_22640);
nor U26184 (N_26184,N_24614,N_23485);
nand U26185 (N_26185,N_24864,N_23761);
and U26186 (N_26186,N_23777,N_24543);
nor U26187 (N_26187,N_22959,N_24634);
and U26188 (N_26188,N_22865,N_23203);
nand U26189 (N_26189,N_24855,N_23432);
xor U26190 (N_26190,N_23962,N_22744);
or U26191 (N_26191,N_23370,N_23713);
xor U26192 (N_26192,N_23773,N_22898);
nor U26193 (N_26193,N_24726,N_24710);
nand U26194 (N_26194,N_24397,N_24459);
or U26195 (N_26195,N_23442,N_22701);
or U26196 (N_26196,N_23122,N_23779);
and U26197 (N_26197,N_23397,N_23456);
and U26198 (N_26198,N_22763,N_24778);
or U26199 (N_26199,N_24233,N_23385);
nand U26200 (N_26200,N_22809,N_23694);
nand U26201 (N_26201,N_23829,N_24004);
xnor U26202 (N_26202,N_24244,N_24619);
xor U26203 (N_26203,N_23574,N_24914);
and U26204 (N_26204,N_23899,N_23322);
or U26205 (N_26205,N_23028,N_22619);
xor U26206 (N_26206,N_23746,N_22653);
xor U26207 (N_26207,N_24378,N_24048);
nand U26208 (N_26208,N_24372,N_24998);
and U26209 (N_26209,N_23073,N_22754);
and U26210 (N_26210,N_22841,N_24307);
xor U26211 (N_26211,N_22933,N_23254);
and U26212 (N_26212,N_24136,N_23559);
nand U26213 (N_26213,N_23823,N_24920);
nand U26214 (N_26214,N_22520,N_24763);
nand U26215 (N_26215,N_24627,N_24699);
and U26216 (N_26216,N_22940,N_23526);
xnor U26217 (N_26217,N_23160,N_23992);
or U26218 (N_26218,N_23386,N_23766);
or U26219 (N_26219,N_22760,N_23547);
and U26220 (N_26220,N_22735,N_24603);
or U26221 (N_26221,N_22916,N_22945);
nor U26222 (N_26222,N_23741,N_23760);
nor U26223 (N_26223,N_24801,N_24033);
nor U26224 (N_26224,N_23566,N_24025);
xor U26225 (N_26225,N_24082,N_24089);
or U26226 (N_26226,N_24468,N_23152);
nor U26227 (N_26227,N_24305,N_23524);
nand U26228 (N_26228,N_24123,N_22947);
or U26229 (N_26229,N_23235,N_22599);
xnor U26230 (N_26230,N_23424,N_23480);
and U26231 (N_26231,N_24884,N_24027);
or U26232 (N_26232,N_24981,N_22666);
or U26233 (N_26233,N_22531,N_24594);
or U26234 (N_26234,N_22672,N_24584);
xor U26235 (N_26235,N_22545,N_24768);
nor U26236 (N_26236,N_23141,N_22732);
nand U26237 (N_26237,N_23367,N_23556);
or U26238 (N_26238,N_22608,N_23166);
xnor U26239 (N_26239,N_24852,N_24241);
xor U26240 (N_26240,N_23902,N_24509);
nor U26241 (N_26241,N_24177,N_22953);
or U26242 (N_26242,N_24081,N_24885);
and U26243 (N_26243,N_23539,N_23077);
xor U26244 (N_26244,N_24525,N_24715);
xor U26245 (N_26245,N_24065,N_24599);
nand U26246 (N_26246,N_24020,N_22991);
or U26247 (N_26247,N_24226,N_22639);
and U26248 (N_26248,N_24691,N_23749);
nor U26249 (N_26249,N_24473,N_24453);
and U26250 (N_26250,N_23543,N_24093);
or U26251 (N_26251,N_23104,N_22715);
or U26252 (N_26252,N_23003,N_24513);
and U26253 (N_26253,N_23400,N_23110);
nand U26254 (N_26254,N_23081,N_23114);
nor U26255 (N_26255,N_23664,N_24427);
and U26256 (N_26256,N_24973,N_22605);
xor U26257 (N_26257,N_23478,N_24878);
or U26258 (N_26258,N_24131,N_23191);
and U26259 (N_26259,N_23397,N_22926);
xnor U26260 (N_26260,N_23373,N_23823);
nor U26261 (N_26261,N_22808,N_23103);
or U26262 (N_26262,N_24938,N_23435);
nor U26263 (N_26263,N_22715,N_24699);
nor U26264 (N_26264,N_22571,N_22948);
nand U26265 (N_26265,N_23812,N_24419);
xor U26266 (N_26266,N_23890,N_24843);
or U26267 (N_26267,N_24478,N_24120);
nor U26268 (N_26268,N_22993,N_24683);
nor U26269 (N_26269,N_23098,N_24192);
and U26270 (N_26270,N_24534,N_22945);
and U26271 (N_26271,N_24578,N_23886);
xnor U26272 (N_26272,N_22805,N_23411);
or U26273 (N_26273,N_23798,N_24520);
xnor U26274 (N_26274,N_24355,N_24922);
and U26275 (N_26275,N_24374,N_22622);
nor U26276 (N_26276,N_24743,N_22877);
xor U26277 (N_26277,N_23087,N_22735);
nor U26278 (N_26278,N_23988,N_23978);
and U26279 (N_26279,N_23657,N_24937);
nor U26280 (N_26280,N_23032,N_24925);
xnor U26281 (N_26281,N_23166,N_23920);
nor U26282 (N_26282,N_24704,N_23927);
nand U26283 (N_26283,N_24611,N_23601);
or U26284 (N_26284,N_23574,N_23827);
or U26285 (N_26285,N_24813,N_24308);
nand U26286 (N_26286,N_24407,N_24960);
xnor U26287 (N_26287,N_22824,N_24896);
nand U26288 (N_26288,N_23860,N_24004);
or U26289 (N_26289,N_23514,N_22755);
and U26290 (N_26290,N_23316,N_22911);
and U26291 (N_26291,N_23169,N_23998);
and U26292 (N_26292,N_24949,N_23162);
xor U26293 (N_26293,N_23317,N_23150);
or U26294 (N_26294,N_24213,N_22527);
xnor U26295 (N_26295,N_23573,N_23634);
xor U26296 (N_26296,N_22596,N_24141);
or U26297 (N_26297,N_24740,N_24182);
xor U26298 (N_26298,N_22559,N_24327);
nor U26299 (N_26299,N_22737,N_22662);
and U26300 (N_26300,N_24772,N_22558);
or U26301 (N_26301,N_24206,N_23575);
nor U26302 (N_26302,N_23207,N_22969);
or U26303 (N_26303,N_22880,N_23883);
xnor U26304 (N_26304,N_22788,N_23748);
nor U26305 (N_26305,N_22605,N_24783);
and U26306 (N_26306,N_23524,N_23364);
or U26307 (N_26307,N_24924,N_24228);
xnor U26308 (N_26308,N_24032,N_23911);
or U26309 (N_26309,N_24563,N_24187);
nand U26310 (N_26310,N_24186,N_23426);
and U26311 (N_26311,N_22913,N_24554);
and U26312 (N_26312,N_23962,N_22933);
xor U26313 (N_26313,N_24252,N_23458);
nand U26314 (N_26314,N_23700,N_24963);
and U26315 (N_26315,N_24330,N_23600);
nor U26316 (N_26316,N_23983,N_23496);
xor U26317 (N_26317,N_23133,N_24161);
nor U26318 (N_26318,N_24056,N_23335);
and U26319 (N_26319,N_23897,N_22730);
xnor U26320 (N_26320,N_24526,N_24199);
and U26321 (N_26321,N_22639,N_24731);
nand U26322 (N_26322,N_23799,N_23886);
xnor U26323 (N_26323,N_24249,N_23293);
nand U26324 (N_26324,N_23219,N_24582);
and U26325 (N_26325,N_24958,N_22908);
nor U26326 (N_26326,N_22985,N_23669);
nand U26327 (N_26327,N_22516,N_23667);
xor U26328 (N_26328,N_23432,N_23505);
nand U26329 (N_26329,N_23780,N_23455);
or U26330 (N_26330,N_24293,N_24882);
or U26331 (N_26331,N_22823,N_24722);
nor U26332 (N_26332,N_23552,N_22854);
nand U26333 (N_26333,N_23089,N_22563);
or U26334 (N_26334,N_22567,N_23102);
or U26335 (N_26335,N_23006,N_23898);
xor U26336 (N_26336,N_23963,N_24345);
nor U26337 (N_26337,N_22575,N_22720);
xor U26338 (N_26338,N_24715,N_23999);
nand U26339 (N_26339,N_24030,N_24481);
and U26340 (N_26340,N_23419,N_23208);
nand U26341 (N_26341,N_22601,N_22506);
nor U26342 (N_26342,N_23387,N_24650);
xor U26343 (N_26343,N_23295,N_23163);
and U26344 (N_26344,N_22965,N_23889);
nor U26345 (N_26345,N_24825,N_24966);
nand U26346 (N_26346,N_24702,N_22885);
xor U26347 (N_26347,N_24087,N_24188);
or U26348 (N_26348,N_23608,N_24802);
and U26349 (N_26349,N_23444,N_24137);
nand U26350 (N_26350,N_24857,N_24203);
and U26351 (N_26351,N_24403,N_23186);
nand U26352 (N_26352,N_23359,N_24931);
xor U26353 (N_26353,N_22689,N_22626);
and U26354 (N_26354,N_24813,N_23253);
and U26355 (N_26355,N_23766,N_24100);
nor U26356 (N_26356,N_23173,N_24586);
and U26357 (N_26357,N_24533,N_23912);
or U26358 (N_26358,N_22554,N_24166);
and U26359 (N_26359,N_24226,N_24380);
or U26360 (N_26360,N_23532,N_24874);
or U26361 (N_26361,N_23213,N_24207);
or U26362 (N_26362,N_24177,N_24957);
and U26363 (N_26363,N_24094,N_24592);
xor U26364 (N_26364,N_23932,N_23534);
nand U26365 (N_26365,N_23275,N_23715);
nand U26366 (N_26366,N_23677,N_23474);
nor U26367 (N_26367,N_22791,N_24718);
or U26368 (N_26368,N_24417,N_23894);
xnor U26369 (N_26369,N_24281,N_23242);
nor U26370 (N_26370,N_22780,N_24768);
or U26371 (N_26371,N_24895,N_22988);
or U26372 (N_26372,N_24077,N_23260);
nor U26373 (N_26373,N_24046,N_23919);
xor U26374 (N_26374,N_23048,N_23708);
or U26375 (N_26375,N_22715,N_24720);
nor U26376 (N_26376,N_23165,N_24613);
xor U26377 (N_26377,N_23576,N_23619);
and U26378 (N_26378,N_22942,N_23020);
nor U26379 (N_26379,N_23913,N_23094);
nand U26380 (N_26380,N_23051,N_23663);
xnor U26381 (N_26381,N_24617,N_24041);
nand U26382 (N_26382,N_23439,N_24024);
and U26383 (N_26383,N_22972,N_23584);
or U26384 (N_26384,N_24142,N_24139);
nor U26385 (N_26385,N_24745,N_22817);
or U26386 (N_26386,N_24647,N_23837);
nand U26387 (N_26387,N_24749,N_24553);
xor U26388 (N_26388,N_24111,N_24626);
or U26389 (N_26389,N_23254,N_22753);
or U26390 (N_26390,N_24107,N_23904);
xnor U26391 (N_26391,N_23848,N_23245);
nand U26392 (N_26392,N_23704,N_23981);
nand U26393 (N_26393,N_24008,N_23267);
nor U26394 (N_26394,N_23989,N_22640);
or U26395 (N_26395,N_22781,N_23805);
and U26396 (N_26396,N_24116,N_24026);
xor U26397 (N_26397,N_23065,N_24116);
xor U26398 (N_26398,N_24013,N_23392);
nor U26399 (N_26399,N_23437,N_24584);
nand U26400 (N_26400,N_22950,N_23253);
nor U26401 (N_26401,N_24542,N_23162);
nor U26402 (N_26402,N_23456,N_24269);
nand U26403 (N_26403,N_24622,N_24477);
xor U26404 (N_26404,N_22579,N_24814);
xnor U26405 (N_26405,N_23852,N_24317);
and U26406 (N_26406,N_23364,N_24621);
xor U26407 (N_26407,N_24256,N_23372);
nor U26408 (N_26408,N_22951,N_24711);
nor U26409 (N_26409,N_23447,N_24592);
nand U26410 (N_26410,N_23927,N_22698);
and U26411 (N_26411,N_23801,N_23984);
xor U26412 (N_26412,N_23258,N_24006);
and U26413 (N_26413,N_24561,N_23989);
nand U26414 (N_26414,N_23840,N_24983);
nand U26415 (N_26415,N_23543,N_24715);
nand U26416 (N_26416,N_23118,N_23488);
nand U26417 (N_26417,N_23573,N_24231);
nor U26418 (N_26418,N_23017,N_24643);
or U26419 (N_26419,N_24678,N_23313);
and U26420 (N_26420,N_24981,N_24024);
xor U26421 (N_26421,N_23303,N_22985);
nor U26422 (N_26422,N_23493,N_23432);
nand U26423 (N_26423,N_24310,N_23579);
nor U26424 (N_26424,N_24575,N_23038);
nor U26425 (N_26425,N_24518,N_22878);
xor U26426 (N_26426,N_23978,N_24222);
nand U26427 (N_26427,N_24182,N_24432);
nand U26428 (N_26428,N_22694,N_22537);
nand U26429 (N_26429,N_24006,N_23606);
nor U26430 (N_26430,N_24948,N_23634);
xnor U26431 (N_26431,N_23703,N_23371);
nand U26432 (N_26432,N_23249,N_24747);
or U26433 (N_26433,N_23510,N_23628);
and U26434 (N_26434,N_24708,N_23131);
nand U26435 (N_26435,N_24217,N_23089);
and U26436 (N_26436,N_22613,N_24504);
nand U26437 (N_26437,N_24045,N_24248);
and U26438 (N_26438,N_23633,N_23279);
nor U26439 (N_26439,N_23795,N_24730);
and U26440 (N_26440,N_22537,N_24687);
or U26441 (N_26441,N_24145,N_24255);
nand U26442 (N_26442,N_23869,N_23849);
xnor U26443 (N_26443,N_23260,N_24994);
nor U26444 (N_26444,N_24955,N_24935);
or U26445 (N_26445,N_23975,N_22544);
xor U26446 (N_26446,N_23069,N_22613);
or U26447 (N_26447,N_23734,N_23385);
nand U26448 (N_26448,N_24679,N_23577);
or U26449 (N_26449,N_23056,N_24522);
nand U26450 (N_26450,N_22611,N_24313);
nand U26451 (N_26451,N_24065,N_22734);
xnor U26452 (N_26452,N_22664,N_23617);
xor U26453 (N_26453,N_22804,N_24539);
nand U26454 (N_26454,N_22620,N_23715);
xor U26455 (N_26455,N_23006,N_23467);
nor U26456 (N_26456,N_22940,N_24181);
or U26457 (N_26457,N_23806,N_23399);
or U26458 (N_26458,N_24119,N_24933);
nor U26459 (N_26459,N_23815,N_24571);
nand U26460 (N_26460,N_24849,N_24967);
nand U26461 (N_26461,N_24164,N_22889);
nor U26462 (N_26462,N_23665,N_24045);
nand U26463 (N_26463,N_24660,N_24348);
xnor U26464 (N_26464,N_22755,N_24082);
nand U26465 (N_26465,N_23154,N_23567);
xor U26466 (N_26466,N_23159,N_24551);
and U26467 (N_26467,N_23180,N_24719);
and U26468 (N_26468,N_23664,N_23428);
or U26469 (N_26469,N_23433,N_24233);
nor U26470 (N_26470,N_23348,N_24291);
nor U26471 (N_26471,N_23499,N_23502);
xnor U26472 (N_26472,N_23172,N_23851);
xnor U26473 (N_26473,N_24074,N_23147);
or U26474 (N_26474,N_22577,N_23880);
nor U26475 (N_26475,N_24478,N_23340);
xor U26476 (N_26476,N_23745,N_23444);
or U26477 (N_26477,N_24676,N_24734);
nand U26478 (N_26478,N_24164,N_23005);
nor U26479 (N_26479,N_22784,N_22755);
nand U26480 (N_26480,N_23768,N_24677);
or U26481 (N_26481,N_24181,N_24476);
nor U26482 (N_26482,N_24594,N_23969);
or U26483 (N_26483,N_23306,N_24759);
xnor U26484 (N_26484,N_22650,N_22588);
nand U26485 (N_26485,N_24357,N_22939);
xnor U26486 (N_26486,N_24531,N_23921);
nand U26487 (N_26487,N_24215,N_24814);
and U26488 (N_26488,N_22860,N_22943);
xnor U26489 (N_26489,N_24216,N_24841);
nor U26490 (N_26490,N_23520,N_24348);
and U26491 (N_26491,N_24625,N_24483);
and U26492 (N_26492,N_23625,N_23177);
nor U26493 (N_26493,N_23586,N_23121);
nand U26494 (N_26494,N_24726,N_23080);
nor U26495 (N_26495,N_23600,N_24180);
nor U26496 (N_26496,N_24435,N_24206);
and U26497 (N_26497,N_23322,N_24004);
or U26498 (N_26498,N_22537,N_22957);
and U26499 (N_26499,N_24679,N_24236);
and U26500 (N_26500,N_24312,N_23477);
xnor U26501 (N_26501,N_23180,N_22877);
and U26502 (N_26502,N_22859,N_23475);
nor U26503 (N_26503,N_23126,N_22936);
xnor U26504 (N_26504,N_23249,N_22594);
nor U26505 (N_26505,N_23540,N_24197);
nor U26506 (N_26506,N_24335,N_24272);
and U26507 (N_26507,N_23487,N_23169);
nor U26508 (N_26508,N_24881,N_23466);
xor U26509 (N_26509,N_22707,N_22567);
nand U26510 (N_26510,N_24655,N_24151);
or U26511 (N_26511,N_22743,N_24893);
nor U26512 (N_26512,N_23179,N_24565);
and U26513 (N_26513,N_24604,N_22946);
and U26514 (N_26514,N_23541,N_24186);
nand U26515 (N_26515,N_23710,N_24354);
nand U26516 (N_26516,N_23821,N_23672);
or U26517 (N_26517,N_24877,N_24821);
and U26518 (N_26518,N_23554,N_24535);
nor U26519 (N_26519,N_24071,N_23908);
nor U26520 (N_26520,N_23999,N_23481);
and U26521 (N_26521,N_22554,N_22854);
xor U26522 (N_26522,N_24000,N_24400);
and U26523 (N_26523,N_22800,N_23627);
nor U26524 (N_26524,N_23679,N_23727);
nor U26525 (N_26525,N_23483,N_24264);
and U26526 (N_26526,N_24995,N_24537);
or U26527 (N_26527,N_23874,N_24042);
and U26528 (N_26528,N_22986,N_23653);
and U26529 (N_26529,N_22926,N_23579);
xor U26530 (N_26530,N_24303,N_23976);
and U26531 (N_26531,N_24770,N_23171);
and U26532 (N_26532,N_22844,N_22654);
nor U26533 (N_26533,N_23478,N_24258);
and U26534 (N_26534,N_23619,N_23530);
nand U26535 (N_26535,N_23882,N_23002);
or U26536 (N_26536,N_23710,N_24979);
nor U26537 (N_26537,N_24956,N_23814);
xnor U26538 (N_26538,N_24966,N_23653);
and U26539 (N_26539,N_24208,N_24402);
nor U26540 (N_26540,N_22939,N_24333);
or U26541 (N_26541,N_23677,N_23263);
nor U26542 (N_26542,N_24009,N_23797);
xnor U26543 (N_26543,N_22766,N_22836);
and U26544 (N_26544,N_24822,N_24650);
xnor U26545 (N_26545,N_22977,N_23130);
and U26546 (N_26546,N_24818,N_24883);
nor U26547 (N_26547,N_22759,N_24265);
and U26548 (N_26548,N_24544,N_23745);
xor U26549 (N_26549,N_23691,N_24575);
or U26550 (N_26550,N_24246,N_23294);
or U26551 (N_26551,N_22641,N_24953);
or U26552 (N_26552,N_24540,N_24489);
or U26553 (N_26553,N_24545,N_22570);
and U26554 (N_26554,N_23775,N_24776);
nor U26555 (N_26555,N_22918,N_24451);
xor U26556 (N_26556,N_22600,N_24955);
xor U26557 (N_26557,N_24621,N_24677);
or U26558 (N_26558,N_24183,N_23078);
and U26559 (N_26559,N_23201,N_23134);
nand U26560 (N_26560,N_22539,N_24248);
nor U26561 (N_26561,N_24692,N_22710);
xor U26562 (N_26562,N_23540,N_24956);
nor U26563 (N_26563,N_23194,N_23727);
xor U26564 (N_26564,N_24055,N_23258);
nor U26565 (N_26565,N_23729,N_24802);
nand U26566 (N_26566,N_24044,N_22688);
nand U26567 (N_26567,N_24981,N_22729);
and U26568 (N_26568,N_23299,N_24680);
and U26569 (N_26569,N_23612,N_24737);
and U26570 (N_26570,N_22568,N_22875);
nor U26571 (N_26571,N_23990,N_23776);
and U26572 (N_26572,N_24821,N_23057);
xnor U26573 (N_26573,N_22671,N_23805);
and U26574 (N_26574,N_23155,N_24186);
and U26575 (N_26575,N_23148,N_23026);
or U26576 (N_26576,N_23675,N_24115);
or U26577 (N_26577,N_24100,N_23173);
nand U26578 (N_26578,N_24517,N_22672);
or U26579 (N_26579,N_23650,N_24902);
and U26580 (N_26580,N_22586,N_24698);
nand U26581 (N_26581,N_23705,N_23058);
or U26582 (N_26582,N_24594,N_23541);
or U26583 (N_26583,N_24918,N_23373);
nand U26584 (N_26584,N_23957,N_22905);
xnor U26585 (N_26585,N_24206,N_24716);
xor U26586 (N_26586,N_24679,N_24809);
xor U26587 (N_26587,N_22988,N_23606);
nand U26588 (N_26588,N_23704,N_24066);
nand U26589 (N_26589,N_24970,N_24808);
nand U26590 (N_26590,N_22556,N_23150);
or U26591 (N_26591,N_24796,N_24591);
or U26592 (N_26592,N_22582,N_22674);
nand U26593 (N_26593,N_24233,N_23882);
or U26594 (N_26594,N_23825,N_24574);
nand U26595 (N_26595,N_23676,N_23831);
nand U26596 (N_26596,N_22714,N_24637);
and U26597 (N_26597,N_23272,N_23535);
nor U26598 (N_26598,N_24815,N_24146);
or U26599 (N_26599,N_23885,N_24714);
xnor U26600 (N_26600,N_24179,N_22567);
nor U26601 (N_26601,N_22750,N_23250);
and U26602 (N_26602,N_23547,N_22635);
and U26603 (N_26603,N_23343,N_23797);
xnor U26604 (N_26604,N_22844,N_23767);
nor U26605 (N_26605,N_24925,N_24432);
nor U26606 (N_26606,N_22803,N_22529);
or U26607 (N_26607,N_22534,N_22845);
or U26608 (N_26608,N_24972,N_24377);
or U26609 (N_26609,N_24920,N_24226);
nor U26610 (N_26610,N_24696,N_24675);
or U26611 (N_26611,N_23824,N_23671);
xor U26612 (N_26612,N_24947,N_22606);
xnor U26613 (N_26613,N_24702,N_22922);
xor U26614 (N_26614,N_22772,N_23339);
and U26615 (N_26615,N_23176,N_22734);
xnor U26616 (N_26616,N_24416,N_22947);
nor U26617 (N_26617,N_23234,N_24471);
xnor U26618 (N_26618,N_22937,N_23030);
xor U26619 (N_26619,N_24128,N_24356);
or U26620 (N_26620,N_23109,N_24783);
and U26621 (N_26621,N_22722,N_23504);
or U26622 (N_26622,N_24393,N_24945);
nor U26623 (N_26623,N_22561,N_23606);
and U26624 (N_26624,N_24707,N_23838);
or U26625 (N_26625,N_23955,N_22610);
nand U26626 (N_26626,N_24090,N_24490);
nand U26627 (N_26627,N_22979,N_24112);
or U26628 (N_26628,N_23366,N_23007);
xor U26629 (N_26629,N_24369,N_24845);
and U26630 (N_26630,N_23396,N_24692);
or U26631 (N_26631,N_24581,N_24215);
xnor U26632 (N_26632,N_24961,N_24682);
and U26633 (N_26633,N_24472,N_23121);
nand U26634 (N_26634,N_23517,N_22930);
and U26635 (N_26635,N_24522,N_22533);
or U26636 (N_26636,N_24340,N_23868);
or U26637 (N_26637,N_23202,N_23045);
xor U26638 (N_26638,N_24234,N_24601);
and U26639 (N_26639,N_23291,N_24223);
nand U26640 (N_26640,N_23051,N_24603);
nand U26641 (N_26641,N_22917,N_22579);
nand U26642 (N_26642,N_23640,N_24324);
or U26643 (N_26643,N_23316,N_23483);
and U26644 (N_26644,N_24623,N_24450);
or U26645 (N_26645,N_23510,N_24590);
xnor U26646 (N_26646,N_22558,N_22733);
nor U26647 (N_26647,N_24141,N_22708);
and U26648 (N_26648,N_22534,N_23353);
and U26649 (N_26649,N_24092,N_23052);
and U26650 (N_26650,N_22566,N_24453);
xor U26651 (N_26651,N_23665,N_23077);
nand U26652 (N_26652,N_23922,N_24219);
or U26653 (N_26653,N_24677,N_24150);
nor U26654 (N_26654,N_23956,N_22776);
nor U26655 (N_26655,N_24527,N_23480);
nor U26656 (N_26656,N_22875,N_24901);
xor U26657 (N_26657,N_24341,N_24133);
xor U26658 (N_26658,N_24800,N_24992);
nor U26659 (N_26659,N_23205,N_24859);
or U26660 (N_26660,N_22878,N_23882);
or U26661 (N_26661,N_23929,N_23928);
xnor U26662 (N_26662,N_24557,N_24653);
xnor U26663 (N_26663,N_23942,N_24298);
or U26664 (N_26664,N_22949,N_23834);
and U26665 (N_26665,N_24110,N_24980);
nand U26666 (N_26666,N_23784,N_23540);
and U26667 (N_26667,N_24639,N_23462);
xor U26668 (N_26668,N_23942,N_22609);
nand U26669 (N_26669,N_24013,N_24432);
xnor U26670 (N_26670,N_23712,N_23606);
or U26671 (N_26671,N_23849,N_24851);
nor U26672 (N_26672,N_24492,N_24323);
nor U26673 (N_26673,N_24621,N_24292);
and U26674 (N_26674,N_23862,N_23665);
or U26675 (N_26675,N_24165,N_24955);
or U26676 (N_26676,N_24982,N_22671);
and U26677 (N_26677,N_24770,N_23232);
xor U26678 (N_26678,N_23318,N_22615);
nand U26679 (N_26679,N_24135,N_22578);
nor U26680 (N_26680,N_23052,N_22671);
nor U26681 (N_26681,N_24693,N_22672);
xor U26682 (N_26682,N_23121,N_22734);
or U26683 (N_26683,N_24382,N_24220);
or U26684 (N_26684,N_24546,N_24523);
xor U26685 (N_26685,N_23635,N_22738);
nor U26686 (N_26686,N_24753,N_24268);
or U26687 (N_26687,N_22701,N_24940);
xnor U26688 (N_26688,N_24283,N_22959);
and U26689 (N_26689,N_23301,N_22801);
xnor U26690 (N_26690,N_22824,N_23713);
or U26691 (N_26691,N_22915,N_24673);
nor U26692 (N_26692,N_24332,N_24766);
and U26693 (N_26693,N_23812,N_22715);
or U26694 (N_26694,N_23420,N_23064);
nand U26695 (N_26695,N_24798,N_23878);
nand U26696 (N_26696,N_22797,N_22851);
and U26697 (N_26697,N_23582,N_24108);
nor U26698 (N_26698,N_23117,N_24311);
nor U26699 (N_26699,N_23167,N_23829);
xor U26700 (N_26700,N_22857,N_23145);
xnor U26701 (N_26701,N_24231,N_22616);
xnor U26702 (N_26702,N_24016,N_23964);
and U26703 (N_26703,N_23060,N_23711);
nor U26704 (N_26704,N_23177,N_23987);
nand U26705 (N_26705,N_22679,N_22954);
and U26706 (N_26706,N_23621,N_23676);
nand U26707 (N_26707,N_23863,N_22817);
or U26708 (N_26708,N_23575,N_24308);
nor U26709 (N_26709,N_23344,N_24491);
or U26710 (N_26710,N_23797,N_23286);
nand U26711 (N_26711,N_22647,N_24098);
xnor U26712 (N_26712,N_23150,N_23924);
xor U26713 (N_26713,N_23803,N_24690);
or U26714 (N_26714,N_24883,N_22592);
nand U26715 (N_26715,N_24117,N_24375);
or U26716 (N_26716,N_23198,N_23993);
nand U26717 (N_26717,N_24830,N_24119);
and U26718 (N_26718,N_23489,N_23176);
nand U26719 (N_26719,N_22897,N_24241);
nand U26720 (N_26720,N_23269,N_24736);
or U26721 (N_26721,N_24111,N_24773);
nand U26722 (N_26722,N_22925,N_23422);
or U26723 (N_26723,N_24648,N_24375);
nor U26724 (N_26724,N_23245,N_22975);
xnor U26725 (N_26725,N_24932,N_23140);
xnor U26726 (N_26726,N_24266,N_24404);
nand U26727 (N_26727,N_23873,N_24049);
nand U26728 (N_26728,N_24666,N_24161);
and U26729 (N_26729,N_23086,N_22663);
and U26730 (N_26730,N_24339,N_24479);
or U26731 (N_26731,N_23545,N_23054);
nor U26732 (N_26732,N_24381,N_23152);
xor U26733 (N_26733,N_23398,N_23251);
nand U26734 (N_26734,N_24269,N_22566);
xnor U26735 (N_26735,N_24350,N_22758);
nor U26736 (N_26736,N_22514,N_24756);
and U26737 (N_26737,N_24834,N_22513);
nor U26738 (N_26738,N_24420,N_23211);
nand U26739 (N_26739,N_22748,N_23283);
or U26740 (N_26740,N_23479,N_23174);
xnor U26741 (N_26741,N_22502,N_24502);
and U26742 (N_26742,N_24364,N_24655);
xor U26743 (N_26743,N_24952,N_22598);
and U26744 (N_26744,N_22686,N_24370);
xnor U26745 (N_26745,N_24438,N_23878);
nor U26746 (N_26746,N_23982,N_23603);
nor U26747 (N_26747,N_23586,N_24792);
nand U26748 (N_26748,N_23546,N_22862);
xor U26749 (N_26749,N_24696,N_23095);
nand U26750 (N_26750,N_23577,N_24961);
nand U26751 (N_26751,N_24630,N_23354);
nand U26752 (N_26752,N_24411,N_24707);
nand U26753 (N_26753,N_24761,N_23665);
and U26754 (N_26754,N_23274,N_24198);
nand U26755 (N_26755,N_22867,N_24753);
or U26756 (N_26756,N_23942,N_24685);
xnor U26757 (N_26757,N_24855,N_23635);
nor U26758 (N_26758,N_24959,N_23765);
nand U26759 (N_26759,N_23624,N_24023);
or U26760 (N_26760,N_24305,N_23869);
xor U26761 (N_26761,N_23311,N_24751);
nor U26762 (N_26762,N_22993,N_22919);
xnor U26763 (N_26763,N_24636,N_23014);
or U26764 (N_26764,N_24771,N_23669);
and U26765 (N_26765,N_22739,N_24618);
and U26766 (N_26766,N_24257,N_24141);
nor U26767 (N_26767,N_23324,N_23270);
and U26768 (N_26768,N_24534,N_24375);
nand U26769 (N_26769,N_24949,N_23807);
nand U26770 (N_26770,N_22790,N_22901);
and U26771 (N_26771,N_23529,N_22860);
xor U26772 (N_26772,N_23653,N_23495);
nand U26773 (N_26773,N_23679,N_24788);
nand U26774 (N_26774,N_23818,N_22831);
nand U26775 (N_26775,N_23375,N_23679);
xnor U26776 (N_26776,N_22661,N_23834);
and U26777 (N_26777,N_24058,N_24046);
or U26778 (N_26778,N_23124,N_23296);
or U26779 (N_26779,N_23286,N_24750);
or U26780 (N_26780,N_23278,N_24818);
or U26781 (N_26781,N_23473,N_24928);
nand U26782 (N_26782,N_24704,N_22725);
xor U26783 (N_26783,N_23104,N_22976);
xnor U26784 (N_26784,N_24077,N_24133);
xor U26785 (N_26785,N_24656,N_22570);
and U26786 (N_26786,N_24706,N_23256);
nand U26787 (N_26787,N_24032,N_24019);
nor U26788 (N_26788,N_23285,N_23781);
xnor U26789 (N_26789,N_24724,N_24839);
nor U26790 (N_26790,N_23500,N_24155);
nand U26791 (N_26791,N_24328,N_23946);
nand U26792 (N_26792,N_23469,N_24653);
or U26793 (N_26793,N_23636,N_23934);
and U26794 (N_26794,N_24131,N_24741);
nor U26795 (N_26795,N_24302,N_22594);
and U26796 (N_26796,N_24878,N_24859);
and U26797 (N_26797,N_24459,N_23340);
nand U26798 (N_26798,N_24958,N_23894);
xnor U26799 (N_26799,N_23000,N_23673);
nor U26800 (N_26800,N_23103,N_23244);
xnor U26801 (N_26801,N_24501,N_24130);
and U26802 (N_26802,N_23378,N_24435);
nor U26803 (N_26803,N_24734,N_24163);
nor U26804 (N_26804,N_23606,N_24424);
nor U26805 (N_26805,N_23958,N_22530);
or U26806 (N_26806,N_23919,N_24744);
and U26807 (N_26807,N_23193,N_24020);
nand U26808 (N_26808,N_23034,N_23569);
xor U26809 (N_26809,N_23350,N_24081);
and U26810 (N_26810,N_23680,N_23110);
xnor U26811 (N_26811,N_23677,N_23442);
nand U26812 (N_26812,N_23753,N_24401);
xnor U26813 (N_26813,N_24235,N_23567);
or U26814 (N_26814,N_22750,N_22869);
nand U26815 (N_26815,N_22755,N_24528);
and U26816 (N_26816,N_24582,N_22648);
or U26817 (N_26817,N_22535,N_23946);
nand U26818 (N_26818,N_23924,N_23980);
nand U26819 (N_26819,N_24742,N_24716);
and U26820 (N_26820,N_22704,N_24076);
xor U26821 (N_26821,N_24034,N_24268);
nand U26822 (N_26822,N_24986,N_23754);
nor U26823 (N_26823,N_24121,N_23282);
or U26824 (N_26824,N_23995,N_23587);
xor U26825 (N_26825,N_22711,N_23229);
nor U26826 (N_26826,N_23465,N_24697);
nand U26827 (N_26827,N_23330,N_23045);
xnor U26828 (N_26828,N_23149,N_24904);
xnor U26829 (N_26829,N_24124,N_23075);
or U26830 (N_26830,N_24877,N_22858);
nor U26831 (N_26831,N_22773,N_24955);
xnor U26832 (N_26832,N_24420,N_23390);
or U26833 (N_26833,N_24182,N_24984);
xor U26834 (N_26834,N_23718,N_24322);
and U26835 (N_26835,N_23297,N_24102);
nand U26836 (N_26836,N_23708,N_23083);
or U26837 (N_26837,N_24985,N_23176);
xor U26838 (N_26838,N_24011,N_24830);
nor U26839 (N_26839,N_23747,N_22871);
nor U26840 (N_26840,N_23335,N_24489);
or U26841 (N_26841,N_23940,N_24073);
and U26842 (N_26842,N_23191,N_24692);
xnor U26843 (N_26843,N_23408,N_24673);
nand U26844 (N_26844,N_23790,N_22879);
xor U26845 (N_26845,N_24312,N_23362);
and U26846 (N_26846,N_23673,N_24453);
nor U26847 (N_26847,N_23213,N_23935);
xor U26848 (N_26848,N_23612,N_23981);
nor U26849 (N_26849,N_22949,N_24179);
nand U26850 (N_26850,N_23231,N_24298);
nand U26851 (N_26851,N_24201,N_23416);
nor U26852 (N_26852,N_22523,N_24887);
and U26853 (N_26853,N_24320,N_23042);
or U26854 (N_26854,N_22969,N_24831);
nand U26855 (N_26855,N_23701,N_24192);
nor U26856 (N_26856,N_23154,N_24821);
or U26857 (N_26857,N_23031,N_23798);
xnor U26858 (N_26858,N_23300,N_22803);
nand U26859 (N_26859,N_24872,N_23366);
nand U26860 (N_26860,N_22695,N_24173);
xnor U26861 (N_26861,N_24655,N_24832);
xnor U26862 (N_26862,N_24213,N_23451);
nand U26863 (N_26863,N_24126,N_24569);
xor U26864 (N_26864,N_24902,N_22642);
xnor U26865 (N_26865,N_23071,N_24524);
nand U26866 (N_26866,N_23972,N_23375);
and U26867 (N_26867,N_23721,N_22797);
xnor U26868 (N_26868,N_22941,N_24587);
xnor U26869 (N_26869,N_23937,N_23503);
or U26870 (N_26870,N_24672,N_24671);
nor U26871 (N_26871,N_23555,N_23480);
nor U26872 (N_26872,N_22910,N_24641);
and U26873 (N_26873,N_23854,N_22638);
nand U26874 (N_26874,N_24434,N_22604);
nand U26875 (N_26875,N_24091,N_23484);
nor U26876 (N_26876,N_24894,N_23357);
and U26877 (N_26877,N_22535,N_24886);
or U26878 (N_26878,N_22526,N_23041);
nor U26879 (N_26879,N_23862,N_24794);
xor U26880 (N_26880,N_24821,N_23704);
nand U26881 (N_26881,N_22674,N_23964);
nor U26882 (N_26882,N_24162,N_24597);
xnor U26883 (N_26883,N_23283,N_23049);
or U26884 (N_26884,N_24634,N_23882);
nor U26885 (N_26885,N_23780,N_22572);
nand U26886 (N_26886,N_23133,N_23126);
xor U26887 (N_26887,N_24523,N_23508);
and U26888 (N_26888,N_24247,N_24655);
xnor U26889 (N_26889,N_24410,N_22741);
and U26890 (N_26890,N_23862,N_24264);
or U26891 (N_26891,N_23422,N_22871);
nand U26892 (N_26892,N_23025,N_23705);
xor U26893 (N_26893,N_24435,N_24800);
and U26894 (N_26894,N_23287,N_23091);
nand U26895 (N_26895,N_24434,N_24312);
or U26896 (N_26896,N_23066,N_23725);
or U26897 (N_26897,N_24759,N_24975);
or U26898 (N_26898,N_24066,N_24086);
xnor U26899 (N_26899,N_24863,N_22576);
and U26900 (N_26900,N_22666,N_22507);
xnor U26901 (N_26901,N_24173,N_24178);
and U26902 (N_26902,N_24291,N_24938);
and U26903 (N_26903,N_23194,N_24688);
or U26904 (N_26904,N_23197,N_24815);
and U26905 (N_26905,N_23881,N_23694);
nor U26906 (N_26906,N_22974,N_24033);
nor U26907 (N_26907,N_23886,N_22793);
or U26908 (N_26908,N_22718,N_23415);
xnor U26909 (N_26909,N_22677,N_23928);
nand U26910 (N_26910,N_22722,N_24914);
and U26911 (N_26911,N_23977,N_22708);
or U26912 (N_26912,N_23509,N_23281);
xnor U26913 (N_26913,N_24223,N_23085);
and U26914 (N_26914,N_23440,N_24106);
xnor U26915 (N_26915,N_23530,N_24197);
and U26916 (N_26916,N_24337,N_22891);
nor U26917 (N_26917,N_24895,N_23559);
xor U26918 (N_26918,N_24335,N_23179);
nand U26919 (N_26919,N_24051,N_23946);
nand U26920 (N_26920,N_24588,N_24869);
nor U26921 (N_26921,N_24647,N_23195);
nand U26922 (N_26922,N_22627,N_23230);
xor U26923 (N_26923,N_22987,N_24002);
or U26924 (N_26924,N_23766,N_24224);
xnor U26925 (N_26925,N_23409,N_22974);
nand U26926 (N_26926,N_24569,N_23647);
nand U26927 (N_26927,N_23627,N_23342);
xor U26928 (N_26928,N_23807,N_23971);
nand U26929 (N_26929,N_23490,N_24139);
nor U26930 (N_26930,N_24529,N_24421);
and U26931 (N_26931,N_23795,N_24959);
nand U26932 (N_26932,N_22795,N_24550);
nand U26933 (N_26933,N_22948,N_22983);
and U26934 (N_26934,N_24282,N_23629);
or U26935 (N_26935,N_22689,N_22758);
nand U26936 (N_26936,N_24864,N_24461);
xor U26937 (N_26937,N_23627,N_24832);
xnor U26938 (N_26938,N_24967,N_24213);
or U26939 (N_26939,N_23600,N_23355);
and U26940 (N_26940,N_23904,N_23214);
nand U26941 (N_26941,N_24283,N_24311);
nand U26942 (N_26942,N_24623,N_22940);
nand U26943 (N_26943,N_22587,N_24506);
or U26944 (N_26944,N_23170,N_22969);
nor U26945 (N_26945,N_24817,N_23849);
xnor U26946 (N_26946,N_23130,N_23728);
nand U26947 (N_26947,N_24259,N_23363);
nor U26948 (N_26948,N_23423,N_23710);
xor U26949 (N_26949,N_24176,N_24458);
xor U26950 (N_26950,N_24908,N_22911);
nor U26951 (N_26951,N_23952,N_23786);
and U26952 (N_26952,N_24187,N_22852);
xor U26953 (N_26953,N_22938,N_23652);
nor U26954 (N_26954,N_23598,N_23148);
and U26955 (N_26955,N_24174,N_22755);
nor U26956 (N_26956,N_22764,N_23632);
xnor U26957 (N_26957,N_22747,N_24416);
xor U26958 (N_26958,N_22965,N_22895);
nand U26959 (N_26959,N_24513,N_22949);
nand U26960 (N_26960,N_23572,N_24489);
xnor U26961 (N_26961,N_24893,N_24855);
xnor U26962 (N_26962,N_23565,N_22839);
nand U26963 (N_26963,N_24436,N_22935);
xnor U26964 (N_26964,N_22552,N_24766);
nor U26965 (N_26965,N_24035,N_23859);
nand U26966 (N_26966,N_24288,N_23603);
xor U26967 (N_26967,N_23213,N_24976);
nor U26968 (N_26968,N_23114,N_24721);
xor U26969 (N_26969,N_23485,N_23362);
nand U26970 (N_26970,N_23515,N_23565);
nand U26971 (N_26971,N_23414,N_24089);
nor U26972 (N_26972,N_23097,N_24093);
nand U26973 (N_26973,N_23045,N_23091);
or U26974 (N_26974,N_24462,N_23938);
nor U26975 (N_26975,N_23928,N_24429);
nand U26976 (N_26976,N_23416,N_24170);
nor U26977 (N_26977,N_23188,N_22977);
xor U26978 (N_26978,N_23331,N_23666);
or U26979 (N_26979,N_23519,N_22961);
nand U26980 (N_26980,N_23089,N_24373);
nor U26981 (N_26981,N_24342,N_22968);
nor U26982 (N_26982,N_24932,N_24174);
nand U26983 (N_26983,N_23228,N_23530);
and U26984 (N_26984,N_23726,N_23677);
nand U26985 (N_26985,N_23215,N_24801);
nand U26986 (N_26986,N_24773,N_24594);
nand U26987 (N_26987,N_22996,N_24192);
nand U26988 (N_26988,N_23297,N_24119);
nor U26989 (N_26989,N_24743,N_24267);
or U26990 (N_26990,N_23957,N_23552);
or U26991 (N_26991,N_23857,N_23898);
xor U26992 (N_26992,N_23602,N_24229);
nor U26993 (N_26993,N_22767,N_24888);
xnor U26994 (N_26994,N_22808,N_23868);
nor U26995 (N_26995,N_23772,N_23946);
nor U26996 (N_26996,N_22859,N_24671);
or U26997 (N_26997,N_24213,N_22503);
nand U26998 (N_26998,N_22555,N_24321);
or U26999 (N_26999,N_24154,N_24500);
and U27000 (N_27000,N_23164,N_24140);
or U27001 (N_27001,N_23609,N_23591);
nand U27002 (N_27002,N_23670,N_24164);
and U27003 (N_27003,N_22504,N_24873);
or U27004 (N_27004,N_24914,N_23342);
or U27005 (N_27005,N_23343,N_23746);
nand U27006 (N_27006,N_24446,N_24836);
nand U27007 (N_27007,N_22964,N_23491);
xor U27008 (N_27008,N_24415,N_23486);
nor U27009 (N_27009,N_23634,N_23088);
xor U27010 (N_27010,N_24889,N_24760);
xor U27011 (N_27011,N_22560,N_23749);
nor U27012 (N_27012,N_23840,N_24261);
nor U27013 (N_27013,N_24206,N_23067);
and U27014 (N_27014,N_22873,N_23154);
xnor U27015 (N_27015,N_24986,N_24315);
nand U27016 (N_27016,N_24496,N_23463);
xor U27017 (N_27017,N_22930,N_23190);
nand U27018 (N_27018,N_22888,N_24208);
or U27019 (N_27019,N_24666,N_23945);
or U27020 (N_27020,N_23966,N_23933);
and U27021 (N_27021,N_24320,N_24269);
nand U27022 (N_27022,N_23828,N_22964);
xor U27023 (N_27023,N_23605,N_24822);
nor U27024 (N_27024,N_23181,N_24592);
or U27025 (N_27025,N_23985,N_23053);
and U27026 (N_27026,N_23227,N_24950);
nand U27027 (N_27027,N_22578,N_22712);
nor U27028 (N_27028,N_23664,N_24902);
nor U27029 (N_27029,N_24102,N_24120);
xor U27030 (N_27030,N_23805,N_22884);
nand U27031 (N_27031,N_23724,N_23736);
or U27032 (N_27032,N_24917,N_24105);
and U27033 (N_27033,N_23355,N_23227);
nor U27034 (N_27034,N_23665,N_23791);
xnor U27035 (N_27035,N_22968,N_23022);
xor U27036 (N_27036,N_24998,N_22897);
nor U27037 (N_27037,N_24841,N_24160);
or U27038 (N_27038,N_23323,N_23620);
and U27039 (N_27039,N_24236,N_23241);
nand U27040 (N_27040,N_23340,N_22728);
or U27041 (N_27041,N_22934,N_22936);
and U27042 (N_27042,N_24017,N_22819);
nor U27043 (N_27043,N_24517,N_23887);
and U27044 (N_27044,N_24041,N_22620);
nor U27045 (N_27045,N_24493,N_24785);
nand U27046 (N_27046,N_24955,N_23487);
nand U27047 (N_27047,N_22994,N_23470);
xor U27048 (N_27048,N_24407,N_24380);
nor U27049 (N_27049,N_22624,N_23237);
nor U27050 (N_27050,N_23781,N_23300);
nand U27051 (N_27051,N_22619,N_24571);
and U27052 (N_27052,N_22887,N_23064);
or U27053 (N_27053,N_23268,N_22789);
and U27054 (N_27054,N_24738,N_22648);
nor U27055 (N_27055,N_22914,N_24171);
xnor U27056 (N_27056,N_23763,N_24592);
or U27057 (N_27057,N_23136,N_24131);
xor U27058 (N_27058,N_24614,N_23737);
and U27059 (N_27059,N_24909,N_23545);
or U27060 (N_27060,N_24638,N_22985);
or U27061 (N_27061,N_24808,N_23525);
nand U27062 (N_27062,N_23676,N_24642);
and U27063 (N_27063,N_24744,N_22851);
or U27064 (N_27064,N_23283,N_23985);
or U27065 (N_27065,N_22809,N_23592);
and U27066 (N_27066,N_22624,N_23467);
and U27067 (N_27067,N_22685,N_24509);
and U27068 (N_27068,N_24553,N_23215);
or U27069 (N_27069,N_23693,N_22823);
and U27070 (N_27070,N_24899,N_22511);
and U27071 (N_27071,N_23474,N_24193);
xor U27072 (N_27072,N_22895,N_24289);
nand U27073 (N_27073,N_24127,N_23731);
or U27074 (N_27074,N_23267,N_24876);
nand U27075 (N_27075,N_24749,N_24148);
or U27076 (N_27076,N_23364,N_24736);
xnor U27077 (N_27077,N_22797,N_22567);
nand U27078 (N_27078,N_23212,N_23517);
and U27079 (N_27079,N_22627,N_24804);
xor U27080 (N_27080,N_24743,N_24871);
and U27081 (N_27081,N_23305,N_24087);
nor U27082 (N_27082,N_24440,N_23657);
nor U27083 (N_27083,N_24481,N_23356);
or U27084 (N_27084,N_23454,N_23654);
nor U27085 (N_27085,N_22708,N_23953);
xnor U27086 (N_27086,N_23112,N_24051);
nor U27087 (N_27087,N_23332,N_24475);
or U27088 (N_27088,N_24770,N_22602);
or U27089 (N_27089,N_24876,N_24885);
or U27090 (N_27090,N_23498,N_24365);
and U27091 (N_27091,N_23511,N_23246);
or U27092 (N_27092,N_24985,N_22827);
and U27093 (N_27093,N_23687,N_24986);
nor U27094 (N_27094,N_24178,N_24342);
and U27095 (N_27095,N_23237,N_24017);
nor U27096 (N_27096,N_22720,N_24615);
xnor U27097 (N_27097,N_23025,N_22676);
and U27098 (N_27098,N_23316,N_22904);
and U27099 (N_27099,N_23526,N_23429);
and U27100 (N_27100,N_23653,N_23469);
nor U27101 (N_27101,N_22764,N_24511);
or U27102 (N_27102,N_23538,N_22902);
nor U27103 (N_27103,N_24293,N_22618);
xnor U27104 (N_27104,N_22881,N_22925);
nand U27105 (N_27105,N_24688,N_24944);
nand U27106 (N_27106,N_24902,N_23543);
nand U27107 (N_27107,N_24149,N_22667);
nand U27108 (N_27108,N_23060,N_23061);
nor U27109 (N_27109,N_24101,N_24924);
nor U27110 (N_27110,N_24136,N_23024);
and U27111 (N_27111,N_24213,N_22582);
or U27112 (N_27112,N_23205,N_24153);
nand U27113 (N_27113,N_24147,N_24363);
nand U27114 (N_27114,N_23649,N_24879);
xor U27115 (N_27115,N_24237,N_22754);
nand U27116 (N_27116,N_23931,N_23465);
xor U27117 (N_27117,N_23750,N_24783);
nor U27118 (N_27118,N_23720,N_23868);
and U27119 (N_27119,N_24623,N_23227);
nand U27120 (N_27120,N_23345,N_24616);
and U27121 (N_27121,N_22738,N_22739);
or U27122 (N_27122,N_24388,N_22825);
or U27123 (N_27123,N_22581,N_22527);
xor U27124 (N_27124,N_23254,N_23709);
nor U27125 (N_27125,N_24627,N_23646);
xor U27126 (N_27126,N_22958,N_23222);
nor U27127 (N_27127,N_23611,N_23382);
nor U27128 (N_27128,N_23899,N_24509);
and U27129 (N_27129,N_23518,N_23691);
nor U27130 (N_27130,N_24361,N_23851);
and U27131 (N_27131,N_22852,N_22669);
xnor U27132 (N_27132,N_24988,N_24476);
nand U27133 (N_27133,N_24185,N_23727);
nor U27134 (N_27134,N_22523,N_24119);
xnor U27135 (N_27135,N_23291,N_23320);
nor U27136 (N_27136,N_23225,N_24321);
xnor U27137 (N_27137,N_23567,N_23839);
and U27138 (N_27138,N_24863,N_24511);
or U27139 (N_27139,N_22557,N_23120);
nand U27140 (N_27140,N_24768,N_23589);
and U27141 (N_27141,N_22675,N_23165);
nor U27142 (N_27142,N_24564,N_23782);
and U27143 (N_27143,N_23691,N_22665);
nor U27144 (N_27144,N_24124,N_23308);
or U27145 (N_27145,N_22707,N_22574);
nor U27146 (N_27146,N_24246,N_23510);
nand U27147 (N_27147,N_22916,N_22925);
and U27148 (N_27148,N_22603,N_23515);
and U27149 (N_27149,N_23568,N_24462);
nor U27150 (N_27150,N_22879,N_22784);
and U27151 (N_27151,N_23254,N_24598);
nor U27152 (N_27152,N_24633,N_24702);
or U27153 (N_27153,N_23008,N_23782);
and U27154 (N_27154,N_24599,N_23551);
or U27155 (N_27155,N_23635,N_24785);
nand U27156 (N_27156,N_22788,N_23611);
nand U27157 (N_27157,N_24877,N_23304);
and U27158 (N_27158,N_22527,N_23242);
and U27159 (N_27159,N_24851,N_23519);
or U27160 (N_27160,N_23688,N_24157);
nand U27161 (N_27161,N_24374,N_24233);
nor U27162 (N_27162,N_24260,N_23803);
nor U27163 (N_27163,N_23212,N_23046);
nand U27164 (N_27164,N_24916,N_23740);
and U27165 (N_27165,N_24883,N_22575);
nor U27166 (N_27166,N_24994,N_23512);
or U27167 (N_27167,N_24040,N_22741);
or U27168 (N_27168,N_23403,N_23095);
nor U27169 (N_27169,N_22688,N_24021);
nor U27170 (N_27170,N_24937,N_23112);
xor U27171 (N_27171,N_24525,N_24382);
nand U27172 (N_27172,N_23563,N_23454);
nand U27173 (N_27173,N_23019,N_24924);
or U27174 (N_27174,N_23639,N_24675);
xor U27175 (N_27175,N_24430,N_22584);
or U27176 (N_27176,N_23426,N_23090);
or U27177 (N_27177,N_24047,N_22786);
xor U27178 (N_27178,N_24727,N_22982);
nor U27179 (N_27179,N_23900,N_22939);
and U27180 (N_27180,N_22812,N_23565);
nor U27181 (N_27181,N_24992,N_24747);
nand U27182 (N_27182,N_24905,N_22908);
xor U27183 (N_27183,N_23430,N_24238);
or U27184 (N_27184,N_23240,N_22574);
nand U27185 (N_27185,N_22774,N_23184);
or U27186 (N_27186,N_24453,N_23181);
and U27187 (N_27187,N_24372,N_23078);
nand U27188 (N_27188,N_23495,N_24102);
xor U27189 (N_27189,N_24844,N_24450);
nand U27190 (N_27190,N_23358,N_23691);
nor U27191 (N_27191,N_24125,N_23724);
and U27192 (N_27192,N_23901,N_23380);
nand U27193 (N_27193,N_24376,N_24450);
or U27194 (N_27194,N_24717,N_23811);
and U27195 (N_27195,N_22585,N_24701);
and U27196 (N_27196,N_23586,N_23789);
nand U27197 (N_27197,N_24683,N_24332);
xnor U27198 (N_27198,N_22952,N_23733);
nand U27199 (N_27199,N_22707,N_23363);
xnor U27200 (N_27200,N_23912,N_24366);
nor U27201 (N_27201,N_24239,N_22507);
or U27202 (N_27202,N_22975,N_24732);
and U27203 (N_27203,N_24033,N_22840);
xnor U27204 (N_27204,N_24533,N_22882);
nand U27205 (N_27205,N_23850,N_24870);
nand U27206 (N_27206,N_24589,N_23346);
nand U27207 (N_27207,N_24761,N_23624);
or U27208 (N_27208,N_22925,N_22740);
nor U27209 (N_27209,N_24145,N_23719);
nand U27210 (N_27210,N_22849,N_23765);
nand U27211 (N_27211,N_23189,N_24092);
or U27212 (N_27212,N_23108,N_24324);
nor U27213 (N_27213,N_23550,N_23763);
xnor U27214 (N_27214,N_24595,N_24776);
nor U27215 (N_27215,N_23078,N_24406);
nor U27216 (N_27216,N_22829,N_24600);
and U27217 (N_27217,N_24784,N_22842);
xor U27218 (N_27218,N_23430,N_23978);
nor U27219 (N_27219,N_23247,N_24467);
nand U27220 (N_27220,N_23137,N_23562);
or U27221 (N_27221,N_22666,N_23710);
or U27222 (N_27222,N_22891,N_23887);
xnor U27223 (N_27223,N_23636,N_24585);
and U27224 (N_27224,N_24461,N_23216);
xor U27225 (N_27225,N_23606,N_23674);
nand U27226 (N_27226,N_22756,N_23477);
or U27227 (N_27227,N_22986,N_24845);
nor U27228 (N_27228,N_23963,N_24728);
and U27229 (N_27229,N_24457,N_24579);
nand U27230 (N_27230,N_22683,N_24786);
nor U27231 (N_27231,N_22910,N_22702);
or U27232 (N_27232,N_23900,N_22888);
xor U27233 (N_27233,N_23949,N_24542);
nand U27234 (N_27234,N_24690,N_24358);
nor U27235 (N_27235,N_24138,N_22560);
nand U27236 (N_27236,N_24165,N_24789);
or U27237 (N_27237,N_24297,N_23398);
or U27238 (N_27238,N_22736,N_22919);
nand U27239 (N_27239,N_23235,N_23883);
and U27240 (N_27240,N_24822,N_23811);
or U27241 (N_27241,N_23435,N_23727);
xnor U27242 (N_27242,N_22798,N_23337);
and U27243 (N_27243,N_24148,N_22922);
nand U27244 (N_27244,N_23238,N_23110);
and U27245 (N_27245,N_23372,N_22825);
xnor U27246 (N_27246,N_22965,N_24885);
or U27247 (N_27247,N_23272,N_24175);
nor U27248 (N_27248,N_23067,N_24007);
and U27249 (N_27249,N_23047,N_23566);
xnor U27250 (N_27250,N_24397,N_24370);
nor U27251 (N_27251,N_24125,N_23735);
nand U27252 (N_27252,N_22704,N_24954);
nand U27253 (N_27253,N_22702,N_24345);
or U27254 (N_27254,N_22955,N_24388);
nor U27255 (N_27255,N_23134,N_23813);
and U27256 (N_27256,N_23883,N_23990);
nor U27257 (N_27257,N_24090,N_23455);
nor U27258 (N_27258,N_22608,N_23896);
nor U27259 (N_27259,N_23872,N_22798);
xnor U27260 (N_27260,N_22508,N_23136);
nor U27261 (N_27261,N_24936,N_24922);
nor U27262 (N_27262,N_24272,N_23105);
xnor U27263 (N_27263,N_22825,N_22642);
nor U27264 (N_27264,N_23016,N_24106);
xnor U27265 (N_27265,N_24647,N_22706);
nand U27266 (N_27266,N_24753,N_23381);
and U27267 (N_27267,N_24351,N_23326);
or U27268 (N_27268,N_23995,N_24251);
xor U27269 (N_27269,N_23209,N_24182);
nand U27270 (N_27270,N_23489,N_24320);
nand U27271 (N_27271,N_22660,N_22630);
xor U27272 (N_27272,N_23302,N_24074);
or U27273 (N_27273,N_23395,N_24575);
nor U27274 (N_27274,N_22532,N_23857);
and U27275 (N_27275,N_24256,N_24072);
or U27276 (N_27276,N_23522,N_24906);
nand U27277 (N_27277,N_23264,N_23133);
nor U27278 (N_27278,N_23964,N_24675);
nor U27279 (N_27279,N_22914,N_22730);
nor U27280 (N_27280,N_23077,N_24769);
nor U27281 (N_27281,N_23838,N_23283);
xnor U27282 (N_27282,N_23735,N_24811);
nor U27283 (N_27283,N_24631,N_23093);
nor U27284 (N_27284,N_23651,N_23611);
xnor U27285 (N_27285,N_24295,N_24976);
and U27286 (N_27286,N_23148,N_23316);
xnor U27287 (N_27287,N_23798,N_24722);
or U27288 (N_27288,N_23660,N_24831);
and U27289 (N_27289,N_23214,N_23590);
and U27290 (N_27290,N_24448,N_24446);
and U27291 (N_27291,N_23577,N_24736);
and U27292 (N_27292,N_24447,N_24436);
and U27293 (N_27293,N_22832,N_23120);
or U27294 (N_27294,N_23398,N_23453);
xor U27295 (N_27295,N_24689,N_22823);
xor U27296 (N_27296,N_22626,N_23835);
xnor U27297 (N_27297,N_23713,N_23193);
nand U27298 (N_27298,N_23799,N_24211);
and U27299 (N_27299,N_22912,N_22753);
xnor U27300 (N_27300,N_23993,N_23128);
nand U27301 (N_27301,N_23561,N_23529);
xor U27302 (N_27302,N_24737,N_24148);
xor U27303 (N_27303,N_24563,N_24626);
nor U27304 (N_27304,N_22666,N_24709);
nor U27305 (N_27305,N_24407,N_24421);
or U27306 (N_27306,N_23480,N_23487);
and U27307 (N_27307,N_23412,N_23303);
nand U27308 (N_27308,N_24319,N_22867);
nand U27309 (N_27309,N_23292,N_22890);
nor U27310 (N_27310,N_23418,N_24757);
or U27311 (N_27311,N_24355,N_23862);
nand U27312 (N_27312,N_23039,N_23037);
nand U27313 (N_27313,N_24819,N_24203);
nand U27314 (N_27314,N_24048,N_22936);
nand U27315 (N_27315,N_22922,N_23460);
nand U27316 (N_27316,N_24540,N_24001);
xnor U27317 (N_27317,N_22609,N_23442);
xor U27318 (N_27318,N_23300,N_23661);
or U27319 (N_27319,N_23940,N_24865);
xnor U27320 (N_27320,N_23261,N_23327);
nand U27321 (N_27321,N_24140,N_22734);
and U27322 (N_27322,N_24052,N_23406);
xor U27323 (N_27323,N_24257,N_24596);
nor U27324 (N_27324,N_24547,N_24758);
xnor U27325 (N_27325,N_22791,N_23629);
nor U27326 (N_27326,N_24790,N_24024);
and U27327 (N_27327,N_24233,N_23618);
or U27328 (N_27328,N_24247,N_23380);
and U27329 (N_27329,N_23808,N_23001);
or U27330 (N_27330,N_23346,N_24940);
nand U27331 (N_27331,N_23672,N_24364);
nand U27332 (N_27332,N_22662,N_23312);
nor U27333 (N_27333,N_24165,N_24213);
nor U27334 (N_27334,N_24845,N_24744);
nor U27335 (N_27335,N_23330,N_24707);
xor U27336 (N_27336,N_24559,N_23207);
nand U27337 (N_27337,N_22581,N_24847);
nand U27338 (N_27338,N_22738,N_23399);
and U27339 (N_27339,N_24641,N_23482);
or U27340 (N_27340,N_23045,N_22897);
nor U27341 (N_27341,N_23104,N_23389);
xnor U27342 (N_27342,N_22985,N_22543);
nor U27343 (N_27343,N_23366,N_23934);
nor U27344 (N_27344,N_22986,N_24910);
nor U27345 (N_27345,N_22952,N_24536);
nand U27346 (N_27346,N_23895,N_24164);
or U27347 (N_27347,N_22531,N_24556);
xnor U27348 (N_27348,N_24044,N_23838);
or U27349 (N_27349,N_22907,N_24775);
nor U27350 (N_27350,N_24111,N_23962);
nor U27351 (N_27351,N_24948,N_24041);
nand U27352 (N_27352,N_23186,N_23339);
xnor U27353 (N_27353,N_23083,N_24123);
xor U27354 (N_27354,N_23488,N_23791);
nor U27355 (N_27355,N_24319,N_22976);
nand U27356 (N_27356,N_24983,N_23632);
xor U27357 (N_27357,N_22539,N_23129);
nor U27358 (N_27358,N_24691,N_23357);
and U27359 (N_27359,N_22896,N_24594);
and U27360 (N_27360,N_23641,N_23317);
nor U27361 (N_27361,N_22977,N_23664);
xnor U27362 (N_27362,N_23335,N_24269);
or U27363 (N_27363,N_24774,N_24812);
xnor U27364 (N_27364,N_24375,N_24175);
nand U27365 (N_27365,N_24022,N_22550);
or U27366 (N_27366,N_24977,N_22614);
nor U27367 (N_27367,N_22755,N_24276);
or U27368 (N_27368,N_23047,N_22744);
nand U27369 (N_27369,N_22605,N_22785);
nand U27370 (N_27370,N_22525,N_24668);
nor U27371 (N_27371,N_24920,N_22801);
nor U27372 (N_27372,N_24060,N_22763);
nand U27373 (N_27373,N_24034,N_24735);
xnor U27374 (N_27374,N_23186,N_24118);
and U27375 (N_27375,N_24944,N_23356);
nor U27376 (N_27376,N_24592,N_23190);
nor U27377 (N_27377,N_23786,N_24321);
nor U27378 (N_27378,N_23731,N_22869);
xor U27379 (N_27379,N_24342,N_23572);
nor U27380 (N_27380,N_23098,N_24444);
xnor U27381 (N_27381,N_23380,N_23198);
or U27382 (N_27382,N_24508,N_24908);
nand U27383 (N_27383,N_24335,N_24995);
nor U27384 (N_27384,N_23081,N_23934);
nor U27385 (N_27385,N_24232,N_24625);
xor U27386 (N_27386,N_24049,N_24517);
xor U27387 (N_27387,N_24778,N_24080);
xnor U27388 (N_27388,N_24211,N_23441);
xnor U27389 (N_27389,N_22821,N_24609);
and U27390 (N_27390,N_22897,N_24424);
xnor U27391 (N_27391,N_24586,N_23885);
nor U27392 (N_27392,N_22817,N_24691);
nand U27393 (N_27393,N_24233,N_24181);
and U27394 (N_27394,N_23085,N_24777);
nor U27395 (N_27395,N_24142,N_24493);
and U27396 (N_27396,N_24498,N_22902);
or U27397 (N_27397,N_23182,N_24455);
nand U27398 (N_27398,N_23433,N_24486);
and U27399 (N_27399,N_23377,N_23429);
xor U27400 (N_27400,N_23072,N_23184);
nor U27401 (N_27401,N_22524,N_23790);
nor U27402 (N_27402,N_24880,N_24661);
xor U27403 (N_27403,N_23224,N_22679);
xnor U27404 (N_27404,N_24641,N_23460);
or U27405 (N_27405,N_22779,N_22501);
nand U27406 (N_27406,N_23225,N_23035);
xnor U27407 (N_27407,N_24283,N_24260);
nor U27408 (N_27408,N_24156,N_22733);
nand U27409 (N_27409,N_23550,N_23823);
and U27410 (N_27410,N_24414,N_24522);
and U27411 (N_27411,N_23272,N_24354);
xnor U27412 (N_27412,N_23754,N_22802);
and U27413 (N_27413,N_23978,N_24649);
nor U27414 (N_27414,N_23570,N_23199);
nor U27415 (N_27415,N_24268,N_23770);
and U27416 (N_27416,N_24259,N_23512);
xnor U27417 (N_27417,N_24143,N_24972);
xnor U27418 (N_27418,N_23390,N_23001);
and U27419 (N_27419,N_24045,N_22800);
nor U27420 (N_27420,N_23698,N_24831);
xor U27421 (N_27421,N_23097,N_23289);
nand U27422 (N_27422,N_24080,N_24453);
nor U27423 (N_27423,N_23411,N_24642);
xor U27424 (N_27424,N_24209,N_24962);
xnor U27425 (N_27425,N_24804,N_22871);
nand U27426 (N_27426,N_24289,N_24341);
nand U27427 (N_27427,N_22916,N_24525);
or U27428 (N_27428,N_23311,N_24817);
nand U27429 (N_27429,N_24518,N_24900);
xor U27430 (N_27430,N_23325,N_24658);
xnor U27431 (N_27431,N_22908,N_23037);
and U27432 (N_27432,N_23472,N_23188);
or U27433 (N_27433,N_22507,N_24209);
and U27434 (N_27434,N_22533,N_22556);
xor U27435 (N_27435,N_23293,N_22653);
xnor U27436 (N_27436,N_24235,N_24846);
xnor U27437 (N_27437,N_24981,N_24135);
nand U27438 (N_27438,N_22634,N_22507);
nor U27439 (N_27439,N_24299,N_23455);
or U27440 (N_27440,N_23845,N_23861);
nor U27441 (N_27441,N_22981,N_23782);
nand U27442 (N_27442,N_22849,N_23304);
or U27443 (N_27443,N_24909,N_23263);
and U27444 (N_27444,N_23781,N_24155);
nand U27445 (N_27445,N_22509,N_24444);
or U27446 (N_27446,N_23902,N_24646);
nor U27447 (N_27447,N_23536,N_22692);
nand U27448 (N_27448,N_24926,N_24978);
and U27449 (N_27449,N_23608,N_22875);
nor U27450 (N_27450,N_23122,N_24996);
nor U27451 (N_27451,N_24285,N_24412);
and U27452 (N_27452,N_23240,N_22609);
nor U27453 (N_27453,N_23343,N_24208);
or U27454 (N_27454,N_23418,N_23835);
and U27455 (N_27455,N_22562,N_24989);
nand U27456 (N_27456,N_23639,N_24960);
nand U27457 (N_27457,N_24386,N_23729);
and U27458 (N_27458,N_23999,N_23540);
nand U27459 (N_27459,N_23085,N_23391);
nor U27460 (N_27460,N_23185,N_23878);
and U27461 (N_27461,N_23287,N_23020);
nand U27462 (N_27462,N_23329,N_23692);
nand U27463 (N_27463,N_24345,N_24750);
nand U27464 (N_27464,N_23963,N_23160);
nand U27465 (N_27465,N_22840,N_22627);
and U27466 (N_27466,N_23385,N_23281);
and U27467 (N_27467,N_23726,N_24313);
xor U27468 (N_27468,N_23084,N_22739);
nand U27469 (N_27469,N_23033,N_23657);
xor U27470 (N_27470,N_22967,N_23108);
and U27471 (N_27471,N_24376,N_22958);
or U27472 (N_27472,N_24011,N_23219);
or U27473 (N_27473,N_24014,N_24028);
nand U27474 (N_27474,N_23592,N_24147);
nand U27475 (N_27475,N_24939,N_22528);
nor U27476 (N_27476,N_24882,N_23827);
xor U27477 (N_27477,N_23361,N_24502);
nand U27478 (N_27478,N_24220,N_23912);
and U27479 (N_27479,N_22732,N_22503);
nor U27480 (N_27480,N_23932,N_23842);
xnor U27481 (N_27481,N_24546,N_23935);
and U27482 (N_27482,N_24558,N_22811);
nor U27483 (N_27483,N_23972,N_23501);
nand U27484 (N_27484,N_23014,N_23787);
nand U27485 (N_27485,N_24962,N_24665);
and U27486 (N_27486,N_22757,N_23623);
nor U27487 (N_27487,N_23571,N_24973);
and U27488 (N_27488,N_22924,N_22579);
or U27489 (N_27489,N_23759,N_24340);
or U27490 (N_27490,N_23186,N_23912);
nand U27491 (N_27491,N_24218,N_22547);
or U27492 (N_27492,N_23556,N_23009);
nand U27493 (N_27493,N_23868,N_23373);
and U27494 (N_27494,N_24055,N_22691);
nor U27495 (N_27495,N_23972,N_23317);
or U27496 (N_27496,N_24775,N_23045);
or U27497 (N_27497,N_24862,N_23394);
or U27498 (N_27498,N_24747,N_24241);
or U27499 (N_27499,N_23359,N_23916);
or U27500 (N_27500,N_27222,N_25830);
and U27501 (N_27501,N_26403,N_27030);
or U27502 (N_27502,N_27016,N_26861);
xor U27503 (N_27503,N_27138,N_27190);
nand U27504 (N_27504,N_27461,N_26082);
xor U27505 (N_27505,N_26895,N_26996);
nand U27506 (N_27506,N_26104,N_25583);
or U27507 (N_27507,N_26840,N_25113);
or U27508 (N_27508,N_27313,N_25204);
nand U27509 (N_27509,N_26411,N_26136);
nor U27510 (N_27510,N_27234,N_26149);
xor U27511 (N_27511,N_27272,N_26657);
or U27512 (N_27512,N_25897,N_27176);
nand U27513 (N_27513,N_25304,N_25868);
or U27514 (N_27514,N_27162,N_25738);
xor U27515 (N_27515,N_26547,N_26659);
and U27516 (N_27516,N_25071,N_26365);
nor U27517 (N_27517,N_26542,N_27246);
nor U27518 (N_27518,N_25865,N_26930);
and U27519 (N_27519,N_25674,N_25112);
and U27520 (N_27520,N_26453,N_25266);
and U27521 (N_27521,N_27207,N_26604);
nand U27522 (N_27522,N_26218,N_25318);
and U27523 (N_27523,N_25426,N_27035);
and U27524 (N_27524,N_25351,N_26451);
and U27525 (N_27525,N_27054,N_26828);
xor U27526 (N_27526,N_27331,N_25983);
nand U27527 (N_27527,N_25264,N_27482);
and U27528 (N_27528,N_26617,N_27282);
and U27529 (N_27529,N_25160,N_26631);
and U27530 (N_27530,N_25591,N_26535);
nand U27531 (N_27531,N_25746,N_26327);
nand U27532 (N_27532,N_25059,N_25612);
xnor U27533 (N_27533,N_25507,N_26269);
or U27534 (N_27534,N_25791,N_27367);
and U27535 (N_27535,N_25793,N_26837);
or U27536 (N_27536,N_26129,N_25068);
xor U27537 (N_27537,N_27354,N_25963);
and U27538 (N_27538,N_25989,N_26879);
xnor U27539 (N_27539,N_25907,N_25012);
xnor U27540 (N_27540,N_27368,N_26097);
and U27541 (N_27541,N_27450,N_26958);
xnor U27542 (N_27542,N_26199,N_25713);
and U27543 (N_27543,N_26198,N_25592);
xor U27544 (N_27544,N_25052,N_25329);
and U27545 (N_27545,N_26810,N_25905);
xor U27546 (N_27546,N_26039,N_25536);
or U27547 (N_27547,N_27244,N_26668);
and U27548 (N_27548,N_25586,N_25107);
xnor U27549 (N_27549,N_26170,N_26557);
xor U27550 (N_27550,N_26138,N_26296);
nand U27551 (N_27551,N_26119,N_27305);
xnor U27552 (N_27552,N_25640,N_26417);
nor U27553 (N_27553,N_25566,N_26941);
nand U27554 (N_27554,N_25794,N_27494);
and U27555 (N_27555,N_26144,N_25152);
or U27556 (N_27556,N_25171,N_26445);
nand U27557 (N_27557,N_26421,N_25360);
and U27558 (N_27558,N_25365,N_26181);
nand U27559 (N_27559,N_26666,N_26654);
xor U27560 (N_27560,N_26456,N_27416);
and U27561 (N_27561,N_25981,N_25325);
xnor U27562 (N_27562,N_25652,N_25655);
nor U27563 (N_27563,N_25557,N_27084);
xor U27564 (N_27564,N_26917,N_25946);
nor U27565 (N_27565,N_26044,N_27134);
nand U27566 (N_27566,N_25486,N_25632);
or U27567 (N_27567,N_25103,N_26795);
or U27568 (N_27568,N_26592,N_25386);
nor U27569 (N_27569,N_27019,N_25142);
nand U27570 (N_27570,N_26527,N_27100);
and U27571 (N_27571,N_27433,N_26863);
xor U27572 (N_27572,N_26574,N_26802);
or U27573 (N_27573,N_25747,N_25589);
and U27574 (N_27574,N_25378,N_26094);
xnor U27575 (N_27575,N_26134,N_25022);
and U27576 (N_27576,N_26771,N_25416);
and U27577 (N_27577,N_25229,N_26823);
or U27578 (N_27578,N_25331,N_26226);
nor U27579 (N_27579,N_25526,N_26706);
and U27580 (N_27580,N_26115,N_27146);
or U27581 (N_27581,N_26680,N_25452);
or U27582 (N_27582,N_25125,N_25273);
xor U27583 (N_27583,N_26105,N_25294);
and U27584 (N_27584,N_25228,N_25305);
or U27585 (N_27585,N_25222,N_25484);
or U27586 (N_27586,N_25197,N_27298);
or U27587 (N_27587,N_26686,N_25493);
xnor U27588 (N_27588,N_25104,N_27475);
or U27589 (N_27589,N_25036,N_25182);
nand U27590 (N_27590,N_27017,N_26948);
or U27591 (N_27591,N_25827,N_26068);
and U27592 (N_27592,N_26896,N_26767);
nor U27593 (N_27593,N_25672,N_26600);
nor U27594 (N_27594,N_26845,N_26041);
and U27595 (N_27595,N_25205,N_26818);
nor U27596 (N_27596,N_25710,N_26153);
and U27597 (N_27597,N_25853,N_27446);
nor U27598 (N_27598,N_25997,N_25321);
nand U27599 (N_27599,N_25395,N_26834);
or U27600 (N_27600,N_26781,N_26057);
or U27601 (N_27601,N_27068,N_25418);
xnor U27602 (N_27602,N_26311,N_25720);
and U27603 (N_27603,N_26211,N_25976);
xnor U27604 (N_27604,N_25780,N_25906);
nand U27605 (N_27605,N_26185,N_26467);
and U27606 (N_27606,N_25616,N_26983);
and U27607 (N_27607,N_26869,N_26559);
nor U27608 (N_27608,N_26333,N_25006);
and U27609 (N_27609,N_25163,N_25024);
and U27610 (N_27610,N_26491,N_26926);
or U27611 (N_27611,N_26335,N_25538);
xnor U27612 (N_27612,N_25885,N_26258);
nand U27613 (N_27613,N_26384,N_26867);
nor U27614 (N_27614,N_25080,N_26699);
xor U27615 (N_27615,N_27193,N_26914);
nor U27616 (N_27616,N_26748,N_26871);
xnor U27617 (N_27617,N_26239,N_26159);
and U27618 (N_27618,N_25792,N_27008);
nand U27619 (N_27619,N_26415,N_27290);
or U27620 (N_27620,N_25096,N_27071);
nor U27621 (N_27621,N_25320,N_27294);
or U27622 (N_27622,N_25604,N_27439);
nand U27623 (N_27623,N_26088,N_25563);
or U27624 (N_27624,N_25813,N_26570);
and U27625 (N_27625,N_26851,N_25137);
and U27626 (N_27626,N_26233,N_27140);
nor U27627 (N_27627,N_27306,N_27277);
xor U27628 (N_27628,N_25520,N_26207);
nor U27629 (N_27629,N_26644,N_25786);
nor U27630 (N_27630,N_25013,N_27063);
and U27631 (N_27631,N_27281,N_25300);
xor U27632 (N_27632,N_26897,N_25157);
nor U27633 (N_27633,N_27179,N_26430);
or U27634 (N_27634,N_27120,N_27421);
nand U27635 (N_27635,N_26911,N_25268);
and U27636 (N_27636,N_25644,N_26681);
nand U27637 (N_27637,N_26006,N_25773);
nand U27638 (N_27638,N_26555,N_26909);
nand U27639 (N_27639,N_26302,N_26540);
nand U27640 (N_27640,N_26908,N_25761);
xor U27641 (N_27641,N_25457,N_25169);
xor U27642 (N_27642,N_25111,N_25755);
nand U27643 (N_27643,N_26792,N_26982);
xor U27644 (N_27644,N_25174,N_25630);
xor U27645 (N_27645,N_27142,N_25777);
xnor U27646 (N_27646,N_25002,N_26987);
and U27647 (N_27647,N_25722,N_26313);
xor U27648 (N_27648,N_27411,N_25145);
nand U27649 (N_27649,N_26721,N_26541);
and U27650 (N_27650,N_25986,N_26562);
xor U27651 (N_27651,N_25399,N_27260);
or U27652 (N_27652,N_25719,N_26368);
or U27653 (N_27653,N_27208,N_27403);
or U27654 (N_27654,N_26326,N_25122);
nor U27655 (N_27655,N_26986,N_26569);
and U27656 (N_27656,N_27401,N_27221);
and U27657 (N_27657,N_26319,N_25432);
nor U27658 (N_27658,N_25322,N_26378);
and U27659 (N_27659,N_26949,N_25134);
nand U27660 (N_27660,N_26977,N_25725);
nand U27661 (N_27661,N_26847,N_25129);
nand U27662 (N_27662,N_27216,N_26798);
nand U27663 (N_27663,N_27099,N_26003);
xnor U27664 (N_27664,N_25186,N_27187);
and U27665 (N_27665,N_25991,N_27286);
or U27666 (N_27666,N_26675,N_26599);
and U27667 (N_27667,N_26971,N_25588);
nand U27668 (N_27668,N_27212,N_25394);
nand U27669 (N_27669,N_26161,N_27022);
and U27670 (N_27670,N_25420,N_25866);
nor U27671 (N_27671,N_26838,N_27192);
and U27672 (N_27672,N_26393,N_26900);
and U27673 (N_27673,N_25825,N_25503);
or U27674 (N_27674,N_25500,N_27449);
or U27675 (N_27675,N_26475,N_25442);
nand U27676 (N_27676,N_27161,N_25642);
nor U27677 (N_27677,N_25849,N_25425);
or U27678 (N_27678,N_26815,N_26640);
nand U27679 (N_27679,N_25224,N_25847);
xor U27680 (N_27680,N_27414,N_27040);
and U27681 (N_27681,N_25451,N_27145);
or U27682 (N_27682,N_25481,N_27078);
or U27683 (N_27683,N_27122,N_25025);
nand U27684 (N_27684,N_25028,N_26292);
or U27685 (N_27685,N_26012,N_25930);
nand U27686 (N_27686,N_27443,N_25390);
nand U27687 (N_27687,N_26274,N_25975);
and U27688 (N_27688,N_25691,N_26270);
nand U27689 (N_27689,N_26860,N_26040);
xor U27690 (N_27690,N_25996,N_27010);
xnor U27691 (N_27691,N_25806,N_27339);
or U27692 (N_27692,N_25745,N_25203);
or U27693 (N_27693,N_25212,N_25048);
xor U27694 (N_27694,N_25307,N_25605);
or U27695 (N_27695,N_26615,N_25333);
nand U27696 (N_27696,N_25367,N_26704);
nand U27697 (N_27697,N_26947,N_26713);
nand U27698 (N_27698,N_25141,N_25686);
or U27699 (N_27699,N_25637,N_25077);
xor U27700 (N_27700,N_26868,N_27188);
and U27701 (N_27701,N_25402,N_25443);
xor U27702 (N_27702,N_26469,N_27185);
nand U27703 (N_27703,N_26217,N_27196);
xnor U27704 (N_27704,N_25090,N_26512);
and U27705 (N_27705,N_26441,N_26755);
xor U27706 (N_27706,N_26758,N_25291);
and U27707 (N_27707,N_26091,N_25415);
or U27708 (N_27708,N_27295,N_26206);
xor U27709 (N_27709,N_26405,N_26854);
xnor U27710 (N_27710,N_26037,N_27168);
nor U27711 (N_27711,N_26817,N_27249);
nor U27712 (N_27712,N_25471,N_26718);
xor U27713 (N_27713,N_27287,N_25032);
xnor U27714 (N_27714,N_26122,N_25593);
or U27715 (N_27715,N_26901,N_26009);
and U27716 (N_27716,N_25492,N_25454);
nand U27717 (N_27717,N_26757,N_25594);
xnor U27718 (N_27718,N_26248,N_26740);
nand U27719 (N_27719,N_26359,N_25364);
or U27720 (N_27720,N_27480,N_25230);
and U27721 (N_27721,N_26919,N_25377);
nor U27722 (N_27722,N_25990,N_26228);
nand U27723 (N_27723,N_26503,N_26090);
nand U27724 (N_27724,N_27156,N_26752);
nand U27725 (N_27725,N_26320,N_26673);
nor U27726 (N_27726,N_27147,N_25184);
xor U27727 (N_27727,N_27173,N_26447);
xnor U27728 (N_27728,N_27311,N_25857);
nand U27729 (N_27729,N_25355,N_26608);
nor U27730 (N_27730,N_25067,N_26197);
nor U27731 (N_27731,N_25833,N_26408);
nor U27732 (N_27732,N_25759,N_26960);
nor U27733 (N_27733,N_27058,N_26306);
or U27734 (N_27734,N_26893,N_26150);
and U27735 (N_27735,N_25623,N_26525);
nand U27736 (N_27736,N_25276,N_26820);
and U27737 (N_27737,N_26321,N_26396);
and U27738 (N_27738,N_26031,N_27137);
or U27739 (N_27739,N_27316,N_26663);
and U27740 (N_27740,N_26598,N_26959);
and U27741 (N_27741,N_27003,N_26450);
xor U27742 (N_27742,N_25105,N_25498);
or U27743 (N_27743,N_25701,N_25347);
and U27744 (N_27744,N_26448,N_25466);
nor U27745 (N_27745,N_26444,N_27301);
nand U27746 (N_27746,N_26052,N_26011);
nor U27747 (N_27747,N_25380,N_26166);
or U27748 (N_27748,N_27130,N_27096);
nand U27749 (N_27749,N_26826,N_25008);
and U27750 (N_27750,N_25949,N_26374);
nand U27751 (N_27751,N_26109,N_27308);
xor U27752 (N_27752,N_26358,N_25290);
nor U27753 (N_27753,N_27189,N_26618);
or U27754 (N_27754,N_27001,N_26912);
and U27755 (N_27755,N_27288,N_27033);
xnor U27756 (N_27756,N_27167,N_27252);
nand U27757 (N_27757,N_27299,N_25660);
or U27758 (N_27758,N_26784,N_27110);
and U27759 (N_27759,N_27093,N_26624);
xnor U27760 (N_27760,N_25735,N_25288);
or U27761 (N_27761,N_26293,N_27293);
nand U27762 (N_27762,N_26202,N_27228);
nor U27763 (N_27763,N_25435,N_26566);
or U27764 (N_27764,N_26312,N_27257);
xor U27765 (N_27765,N_27013,N_26521);
xor U27766 (N_27766,N_26209,N_26392);
and U27767 (N_27767,N_25577,N_26219);
nor U27768 (N_27768,N_27459,N_26332);
or U27769 (N_27769,N_25982,N_25888);
nand U27770 (N_27770,N_26126,N_25317);
xnor U27771 (N_27771,N_25165,N_26377);
and U27772 (N_27772,N_26730,N_26436);
nor U27773 (N_27773,N_25246,N_27029);
nor U27774 (N_27774,N_25037,N_26004);
nor U27775 (N_27775,N_26807,N_26831);
nand U27776 (N_27776,N_27314,N_26371);
nand U27777 (N_27777,N_25734,N_27326);
xor U27778 (N_27778,N_26194,N_26251);
xnor U27779 (N_27779,N_26250,N_26880);
or U27780 (N_27780,N_26936,N_25940);
xor U27781 (N_27781,N_25544,N_27180);
and U27782 (N_27782,N_27210,N_25003);
and U27783 (N_27783,N_26518,N_25584);
or U27784 (N_27784,N_26140,N_26882);
and U27785 (N_27785,N_25543,N_26687);
nand U27786 (N_27786,N_26697,N_25966);
nand U27787 (N_27787,N_27423,N_25688);
nand U27788 (N_27788,N_25094,N_25207);
xor U27789 (N_27789,N_27055,N_25571);
xnor U27790 (N_27790,N_27358,N_25408);
xor U27791 (N_27791,N_26339,N_27342);
nand U27792 (N_27792,N_26746,N_25501);
nand U27793 (N_27793,N_25334,N_27322);
and U27794 (N_27794,N_25121,N_26106);
nor U27795 (N_27795,N_26702,N_27119);
nand U27796 (N_27796,N_26859,N_25699);
nor U27797 (N_27797,N_25869,N_27081);
and U27798 (N_27798,N_25219,N_25533);
and U27799 (N_27799,N_27259,N_25915);
or U27800 (N_27800,N_25608,N_26289);
xnor U27801 (N_27801,N_25014,N_26285);
or U27802 (N_27802,N_25658,N_26772);
and U27803 (N_27803,N_25423,N_26788);
or U27804 (N_27804,N_26264,N_25412);
or U27805 (N_27805,N_26856,N_25265);
and U27806 (N_27806,N_25877,N_25834);
nor U27807 (N_27807,N_25668,N_26790);
xnor U27808 (N_27808,N_25373,N_25895);
and U27809 (N_27809,N_25622,N_26055);
nor U27810 (N_27810,N_27409,N_25808);
nand U27811 (N_27811,N_25928,N_27102);
nor U27812 (N_27812,N_27429,N_26002);
xor U27813 (N_27813,N_25757,N_26343);
or U27814 (N_27814,N_27061,N_26969);
or U27815 (N_27815,N_25569,N_25570);
and U27816 (N_27816,N_26414,N_26634);
nand U27817 (N_27817,N_27083,N_26483);
xor U27818 (N_27818,N_25170,N_26186);
or U27819 (N_27819,N_25731,N_25948);
nand U27820 (N_27820,N_26988,N_26331);
nor U27821 (N_27821,N_25234,N_25958);
nand U27822 (N_27822,N_26999,N_26520);
and U27823 (N_27823,N_25448,N_25695);
nand U27824 (N_27824,N_26210,N_27417);
nand U27825 (N_27825,N_26892,N_27452);
and U27826 (N_27826,N_26545,N_26329);
nor U27827 (N_27827,N_25034,N_25220);
and U27828 (N_27828,N_25771,N_25039);
or U27829 (N_27829,N_27390,N_27031);
and U27830 (N_27830,N_26994,N_27283);
nand U27831 (N_27831,N_26297,N_25397);
xor U27832 (N_27832,N_27225,N_27097);
xor U27833 (N_27833,N_25639,N_25261);
xor U27834 (N_27834,N_27280,N_26388);
or U27835 (N_27835,N_26180,N_26990);
and U27836 (N_27836,N_25098,N_25896);
and U27837 (N_27837,N_25474,N_25467);
nor U27838 (N_27838,N_27114,N_26183);
xnor U27839 (N_27839,N_25078,N_25535);
nor U27840 (N_27840,N_25231,N_25767);
xnor U27841 (N_27841,N_26147,N_25086);
xor U27842 (N_27842,N_26007,N_27402);
nand U27843 (N_27843,N_26498,N_27497);
nand U27844 (N_27844,N_25393,N_26972);
xor U27845 (N_27845,N_25944,N_26310);
xnor U27846 (N_27846,N_25741,N_26092);
nand U27847 (N_27847,N_26220,N_25283);
nand U27848 (N_27848,N_25029,N_25066);
nor U27849 (N_27849,N_26067,N_26418);
or U27850 (N_27850,N_25957,N_25657);
xor U27851 (N_27851,N_27255,N_26072);
and U27852 (N_27852,N_25585,N_26424);
or U27853 (N_27853,N_26811,N_25891);
or U27854 (N_27854,N_25760,N_25770);
xnor U27855 (N_27855,N_25539,N_26693);
and U27856 (N_27856,N_26533,N_25260);
and U27857 (N_27857,N_26030,N_25215);
nand U27858 (N_27858,N_25109,N_25597);
nor U27859 (N_27859,N_25118,N_25095);
and U27860 (N_27860,N_26458,N_26381);
xor U27861 (N_27861,N_27256,N_26279);
nand U27862 (N_27862,N_26244,N_25776);
nor U27863 (N_27863,N_26102,N_25602);
or U27864 (N_27864,N_25050,N_25634);
nand U27865 (N_27865,N_26957,N_26410);
or U27866 (N_27866,N_25476,N_26048);
xnor U27867 (N_27867,N_26212,N_25398);
xnor U27868 (N_27868,N_26674,N_25758);
nand U27869 (N_27869,N_25076,N_25097);
nand U27870 (N_27870,N_26490,N_25817);
nand U27871 (N_27871,N_26862,N_27405);
nand U27872 (N_27872,N_27074,N_26446);
nor U27873 (N_27873,N_26605,N_27465);
or U27874 (N_27874,N_25609,N_26968);
or U27875 (N_27875,N_26502,N_25580);
nor U27876 (N_27876,N_25925,N_25952);
and U27877 (N_27877,N_27343,N_25647);
and U27878 (N_27878,N_27148,N_26137);
xor U27879 (N_27879,N_26222,N_26685);
xnor U27880 (N_27880,N_25936,N_27300);
nor U27881 (N_27881,N_26736,N_25433);
or U27882 (N_27882,N_26355,N_25559);
and U27883 (N_27883,N_25206,N_26084);
nor U27884 (N_27884,N_25703,N_26178);
and U27885 (N_27885,N_26791,N_26386);
and U27886 (N_27886,N_26695,N_25514);
and U27887 (N_27887,N_25807,N_25324);
and U27888 (N_27888,N_27067,N_25766);
or U27889 (N_27889,N_26648,N_25178);
xnor U27890 (N_27890,N_26103,N_26962);
xnor U27891 (N_27891,N_26400,N_25960);
and U27892 (N_27892,N_26769,N_27113);
xnor U27893 (N_27893,N_27387,N_27470);
or U27894 (N_27894,N_26806,N_27165);
and U27895 (N_27895,N_25298,N_26976);
and U27896 (N_27896,N_25370,N_26889);
xnor U27897 (N_27897,N_25621,N_25831);
nor U27898 (N_27898,N_26283,N_25274);
nor U27899 (N_27899,N_26461,N_26543);
xnor U27900 (N_27900,N_25384,N_27455);
nor U27901 (N_27901,N_25601,N_25253);
xnor U27902 (N_27902,N_26708,N_25924);
xor U27903 (N_27903,N_26184,N_26964);
or U27904 (N_27904,N_27117,N_27374);
nand U27905 (N_27905,N_25664,N_25388);
nor U27906 (N_27906,N_25579,N_26073);
nor U27907 (N_27907,N_27404,N_27007);
nor U27908 (N_27908,N_27200,N_26841);
nand U27909 (N_27909,N_25489,N_25117);
nand U27910 (N_27910,N_26412,N_26382);
or U27911 (N_27911,N_25482,N_25185);
and U27912 (N_27912,N_25614,N_26829);
and U27913 (N_27913,N_25669,N_26191);
nor U27914 (N_27914,N_25363,N_25042);
xor U27915 (N_27915,N_27353,N_27247);
and U27916 (N_27916,N_25653,N_27098);
and U27917 (N_27917,N_25239,N_26146);
and U27918 (N_27918,N_26782,N_26937);
and U27919 (N_27919,N_27383,N_25009);
xor U27920 (N_27920,N_25315,N_26492);
nand U27921 (N_27921,N_26588,N_26872);
nor U27922 (N_27922,N_26086,N_25439);
nand U27923 (N_27923,N_25369,N_25843);
and U27924 (N_27924,N_25043,N_25023);
xnor U27925 (N_27925,N_26164,N_25598);
or U27926 (N_27926,N_27408,N_27385);
nor U27927 (N_27927,N_26855,N_25954);
nor U27928 (N_27928,N_26593,N_25774);
or U27929 (N_27929,N_27276,N_25560);
and U27930 (N_27930,N_27079,N_25516);
xnor U27931 (N_27931,N_26954,N_25040);
and U27932 (N_27932,N_26452,N_25547);
xor U27933 (N_27933,N_26553,N_25651);
or U27934 (N_27934,N_25153,N_27062);
nor U27935 (N_27935,N_26071,N_26070);
and U27936 (N_27936,N_26078,N_25342);
nand U27937 (N_27937,N_27462,N_26225);
nand U27938 (N_27938,N_25998,N_26076);
nor U27939 (N_27939,N_26581,N_25323);
or U27940 (N_27940,N_25041,N_27178);
nand U27941 (N_27941,N_26981,N_25821);
xor U27942 (N_27942,N_25422,N_25407);
xnor U27943 (N_27943,N_25978,N_27359);
and U27944 (N_27944,N_27005,N_26108);
and U27945 (N_27945,N_25419,N_26305);
xor U27946 (N_27946,N_26677,N_25309);
xor U27947 (N_27947,N_26989,N_25870);
nand U27948 (N_27948,N_26653,N_26347);
and U27949 (N_27949,N_25082,N_26658);
xnor U27950 (N_27950,N_25555,N_26208);
nor U27951 (N_27951,N_27418,N_26891);
xor U27952 (N_27952,N_25581,N_25387);
xnor U27953 (N_27953,N_25081,N_26822);
nor U27954 (N_27954,N_27080,N_27279);
nand U27955 (N_27955,N_26028,N_25546);
or U27956 (N_27956,N_25567,N_27307);
nor U27957 (N_27957,N_25939,N_26931);
or U27958 (N_27958,N_26703,N_25742);
and U27959 (N_27959,N_25470,N_25465);
nor U27960 (N_27960,N_25804,N_25763);
nor U27961 (N_27961,N_25729,N_27262);
or U27962 (N_27962,N_25973,N_25271);
and U27963 (N_27963,N_26732,N_26852);
or U27964 (N_27964,N_27199,N_26021);
and U27965 (N_27965,N_26918,N_27324);
and U27966 (N_27966,N_27400,N_27194);
xor U27967 (N_27967,N_25385,N_25162);
nor U27968 (N_27968,N_26464,N_26130);
xnor U27969 (N_27969,N_27415,N_26171);
xor U27970 (N_27970,N_26603,N_25438);
nor U27971 (N_27971,N_25826,N_27434);
nand U27972 (N_27972,N_27183,N_26380);
and U27973 (N_27973,N_26563,N_26027);
nand U27974 (N_27974,N_27395,N_25379);
or U27975 (N_27975,N_27496,N_25818);
nand U27976 (N_27976,N_25607,N_26589);
and U27977 (N_27977,N_25556,N_25374);
nor U27978 (N_27978,N_26783,N_25964);
and U27979 (N_27979,N_27251,N_25992);
or U27980 (N_27980,N_26776,N_25837);
nor U27981 (N_27981,N_25856,N_26728);
nor U27982 (N_27982,N_26951,N_25862);
and U27983 (N_27983,N_27352,N_25968);
nor U27984 (N_27984,N_26511,N_26013);
and U27985 (N_27985,N_26158,N_26584);
or U27986 (N_27986,N_25959,N_25988);
nor U27987 (N_27987,N_25781,N_27292);
or U27988 (N_27988,N_26607,N_26291);
xnor U27989 (N_27989,N_25328,N_27164);
nand U27990 (N_27990,N_25819,N_25472);
nand U27991 (N_27991,N_25070,N_26998);
nand U27992 (N_27992,N_25183,N_25822);
xnor U27993 (N_27993,N_26187,N_26360);
xnor U27994 (N_27994,N_27369,N_26515);
nand U27995 (N_27995,N_27492,N_26804);
and U27996 (N_27996,N_26572,N_26029);
xnor U27997 (N_27997,N_25911,N_26707);
nand U27998 (N_27998,N_25226,N_26985);
nand U27999 (N_27999,N_27202,N_26571);
xnor U28000 (N_28000,N_25828,N_25670);
xnor U28001 (N_28001,N_25020,N_25515);
and U28002 (N_28002,N_27493,N_25396);
and U28003 (N_28003,N_25573,N_25680);
nand U28004 (N_28004,N_27386,N_26404);
nor U28005 (N_28005,N_26356,N_26284);
and U28006 (N_28006,N_27357,N_25967);
and U28007 (N_28007,N_26204,N_25613);
xor U28008 (N_28008,N_25899,N_27472);
nand U28009 (N_28009,N_25214,N_25548);
nand U28010 (N_28010,N_26978,N_25461);
and U28011 (N_28011,N_26652,N_26878);
nor U28012 (N_28012,N_25343,N_27253);
nand U28013 (N_28013,N_25285,N_26223);
nand U28014 (N_28014,N_25678,N_27270);
xnor U28015 (N_28015,N_25252,N_27366);
nor U28016 (N_28016,N_26398,N_25269);
nor U28017 (N_28017,N_25576,N_25628);
xnor U28018 (N_28018,N_25417,N_27000);
and U28019 (N_28019,N_26929,N_26338);
nand U28020 (N_28020,N_25277,N_27065);
and U28021 (N_28021,N_25596,N_26500);
and U28022 (N_28022,N_26849,N_26952);
or U28023 (N_28023,N_25236,N_27388);
nand U28024 (N_28024,N_25832,N_25884);
nand U28025 (N_28025,N_26399,N_25803);
nor U28026 (N_28026,N_25509,N_27154);
xor U28027 (N_28027,N_26630,N_25044);
nor U28028 (N_28028,N_26812,N_26672);
nor U28029 (N_28029,N_27424,N_26061);
and U28030 (N_28030,N_27092,N_27360);
or U28031 (N_28031,N_26145,N_26459);
or U28032 (N_28032,N_25666,N_27266);
and U28033 (N_28033,N_26486,N_26286);
or U28034 (N_28034,N_26489,N_25733);
and U28035 (N_28035,N_26480,N_25019);
and U28036 (N_28036,N_25513,N_26616);
nor U28037 (N_28037,N_27048,N_26364);
or U28038 (N_28038,N_27126,N_26117);
and U28039 (N_28039,N_26317,N_27491);
nor U28040 (N_28040,N_26249,N_26036);
nor U28041 (N_28041,N_26636,N_27323);
and U28042 (N_28042,N_25357,N_27315);
or U28043 (N_28043,N_26953,N_26934);
or U28044 (N_28044,N_25031,N_26925);
nand U28045 (N_28045,N_26025,N_26583);
nor U28046 (N_28046,N_25213,N_27489);
nand U28047 (N_28047,N_26100,N_27041);
nand U28048 (N_28048,N_25158,N_27477);
nor U28049 (N_28049,N_25456,N_27442);
or U28050 (N_28050,N_26698,N_25961);
or U28051 (N_28051,N_25434,N_25615);
nand U28052 (N_28052,N_25146,N_26888);
or U28053 (N_28053,N_26449,N_25428);
nor U28054 (N_28054,N_25262,N_25392);
nand U28055 (N_28055,N_26316,N_26830);
and U28056 (N_28056,N_27312,N_26422);
nand U28057 (N_28057,N_27046,N_25698);
or U28058 (N_28058,N_27478,N_26465);
xnor U28059 (N_28059,N_25128,N_27069);
and U28060 (N_28060,N_25886,N_27004);
nor U28061 (N_28061,N_26610,N_25942);
nor U28062 (N_28062,N_27125,N_25123);
nand U28063 (N_28063,N_27471,N_25916);
xnor U28064 (N_28064,N_25690,N_26254);
and U28065 (N_28065,N_25625,N_26282);
nand U28066 (N_28066,N_25716,N_25154);
and U28067 (N_28067,N_25468,N_26843);
nor U28068 (N_28068,N_25053,N_26546);
xnor U28069 (N_28069,N_26263,N_25430);
xnor U28070 (N_28070,N_26290,N_27011);
xnor U28071 (N_28071,N_27483,N_26252);
nand U28072 (N_28072,N_25227,N_27044);
and U28073 (N_28073,N_26114,N_25233);
xnor U28074 (N_28074,N_25180,N_26334);
or U28075 (N_28075,N_25389,N_25823);
nor U28076 (N_28076,N_26932,N_26945);
nor U28077 (N_28077,N_26215,N_27198);
or U28078 (N_28078,N_26363,N_25314);
nand U28079 (N_28079,N_25863,N_26629);
nand U28080 (N_28080,N_27220,N_25049);
nand U28081 (N_28081,N_27009,N_25119);
xor U28082 (N_28082,N_26315,N_27435);
nand U28083 (N_28083,N_25488,N_25292);
or U28084 (N_28084,N_25312,N_26156);
xnor U28085 (N_28085,N_25835,N_27106);
xor U28086 (N_28086,N_26638,N_26743);
nor U28087 (N_28087,N_27393,N_25565);
and U28088 (N_28088,N_25947,N_26438);
nor U28089 (N_28089,N_26715,N_26261);
xnor U28090 (N_28090,N_25383,N_25918);
and U28091 (N_28091,N_25935,N_26729);
xor U28092 (N_28092,N_25270,N_25984);
and U28093 (N_28093,N_25772,N_26858);
nand U28094 (N_28094,N_25648,N_26579);
xnor U28095 (N_28095,N_27376,N_25143);
or U28096 (N_28096,N_25258,N_26670);
and U28097 (N_28097,N_26484,N_26079);
xnor U28098 (N_28098,N_25861,N_26839);
and U28099 (N_28099,N_27318,N_27155);
xor U28100 (N_28100,N_27337,N_27420);
nor U28101 (N_28101,N_25499,N_25809);
and U28102 (N_28102,N_26742,N_25892);
nor U28103 (N_28103,N_26887,N_25120);
or U28104 (N_28104,N_25521,N_26299);
nand U28105 (N_28105,N_25491,N_26789);
or U28106 (N_28106,N_26272,N_26035);
nand U28107 (N_28107,N_25980,N_26726);
or U28108 (N_28108,N_25882,N_26001);
and U28109 (N_28109,N_26397,N_26457);
nor U28110 (N_28110,N_25685,N_26069);
or U28111 (N_28111,N_26833,N_27050);
or U28112 (N_28112,N_25797,N_25524);
and U28113 (N_28113,N_27015,N_25511);
xnor U28114 (N_28114,N_26245,N_25898);
xor U28115 (N_28115,N_25330,N_26975);
nor U28116 (N_28116,N_25700,N_25479);
xor U28117 (N_28117,N_25149,N_26237);
or U28118 (N_28118,N_25871,N_27365);
or U28119 (N_28119,N_27380,N_26288);
nand U28120 (N_28120,N_26779,N_25512);
nand U28121 (N_28121,N_27191,N_26620);
and U28122 (N_28122,N_27370,N_25293);
nand U28123 (N_28123,N_25718,N_26534);
xnor U28124 (N_28124,N_27051,N_26309);
or U28125 (N_28125,N_27135,N_27448);
nand U28126 (N_28126,N_26694,N_26064);
nand U28127 (N_28127,N_25873,N_26560);
or U28128 (N_28128,N_27158,N_26690);
nand U28129 (N_28129,N_26760,N_25661);
nand U28130 (N_28130,N_25730,N_26294);
xor U28131 (N_28131,N_25344,N_26301);
nand U28132 (N_28132,N_25179,N_26622);
nor U28133 (N_28133,N_25744,N_26005);
and U28134 (N_28134,N_26231,N_27344);
nand U28135 (N_28135,N_27021,N_26565);
nand U28136 (N_28136,N_27319,N_25483);
and U28137 (N_28137,N_26850,N_25057);
and U28138 (N_28138,N_26065,N_25775);
or U28139 (N_28139,N_25768,N_25502);
xor U28140 (N_28140,N_26785,N_26967);
and U28141 (N_28141,N_25065,N_25072);
nor U28142 (N_28142,N_26966,N_25173);
or U28143 (N_28143,N_26621,N_27467);
or U28144 (N_28144,N_25166,N_26714);
nor U28145 (N_28145,N_26548,N_26174);
and U28146 (N_28146,N_26481,N_26455);
xnor U28147 (N_28147,N_26902,N_26842);
xor U28148 (N_28148,N_25679,N_26367);
and U28149 (N_28149,N_26213,N_26300);
xnor U28150 (N_28150,N_26409,N_26023);
xnor U28151 (N_28151,N_26907,N_27371);
nand U28152 (N_28152,N_27039,N_25540);
nor U28153 (N_28153,N_26361,N_26734);
and U28154 (N_28154,N_27018,N_26944);
xor U28155 (N_28155,N_26665,N_25189);
nor U28156 (N_28156,N_25812,N_26468);
or U28157 (N_28157,N_27116,N_26087);
and U28158 (N_28158,N_27437,N_25723);
and U28159 (N_28159,N_27042,N_27133);
and U28160 (N_28160,N_27350,N_27232);
xnor U28161 (N_28161,N_25950,N_27310);
nand U28162 (N_28162,N_26575,N_26391);
nor U28163 (N_28163,N_25726,N_26667);
or U28164 (N_28164,N_27238,N_27129);
or U28165 (N_28165,N_25138,N_27087);
and U28166 (N_28166,N_26786,N_26711);
and U28167 (N_28167,N_27499,N_27181);
xor U28168 (N_28168,N_25890,N_27085);
or U28169 (N_28169,N_25092,N_26577);
or U28170 (N_28170,N_27070,N_27101);
nand U28171 (N_28171,N_25427,N_26857);
and U28172 (N_28172,N_26205,N_25549);
nand U28173 (N_28173,N_25671,N_26885);
nor U28174 (N_28174,N_25284,N_26051);
or U28175 (N_28175,N_25574,N_25301);
and U28176 (N_28176,N_26429,N_27153);
and U28177 (N_28177,N_27095,N_25682);
xnor U28178 (N_28178,N_25414,N_27303);
and U28179 (N_28179,N_25450,N_26691);
nand U28180 (N_28180,N_26591,N_25603);
nand U28181 (N_28181,N_26514,N_26096);
nor U28182 (N_28182,N_25839,N_26425);
xor U28183 (N_28183,N_27278,N_25218);
or U28184 (N_28184,N_26123,N_26224);
nor U28185 (N_28185,N_26664,N_27056);
nand U28186 (N_28186,N_25282,N_26303);
or U28187 (N_28187,N_26234,N_26488);
nand U28188 (N_28188,N_26168,N_26257);
nor U28189 (N_28189,N_25693,N_27243);
nor U28190 (N_28190,N_25858,N_27143);
xor U28191 (N_28191,N_27052,N_27254);
or U28192 (N_28192,N_26645,N_27327);
xnor U28193 (N_28193,N_27274,N_26435);
xnor U28194 (N_28194,N_26246,N_26531);
and U28195 (N_28195,N_26336,N_26683);
xor U28196 (N_28196,N_26020,N_25938);
nand U28197 (N_28197,N_25970,N_26649);
xnor U28198 (N_28198,N_27139,N_27269);
and U28199 (N_28199,N_26345,N_27211);
xnor U28200 (N_28200,N_25202,N_27227);
nand U28201 (N_28201,N_27451,N_27127);
xnor U28202 (N_28202,N_25429,N_25665);
nor U28203 (N_28203,N_27267,N_25194);
or U28204 (N_28204,N_26522,N_25455);
xnor U28205 (N_28205,N_26099,N_27291);
nand U28206 (N_28206,N_26827,N_26110);
or U28207 (N_28207,N_25192,N_25552);
nand U28208 (N_28208,N_25217,N_25851);
and U28209 (N_28209,N_25130,N_25056);
xor U28210 (N_28210,N_26942,N_26337);
nor U28211 (N_28211,N_25311,N_27245);
nor U28212 (N_28212,N_27223,N_25287);
and U28213 (N_28213,N_26125,N_25148);
or U28214 (N_28214,N_26524,N_25453);
and U28215 (N_28215,N_26120,N_25626);
nor U28216 (N_28216,N_26406,N_26516);
and U28217 (N_28217,N_26582,N_25063);
xor U28218 (N_28218,N_26075,N_25382);
nor U28219 (N_28219,N_25345,N_26260);
xnor U28220 (N_28220,N_25505,N_25168);
and U28221 (N_28221,N_25133,N_25855);
and U28222 (N_28222,N_26974,N_25475);
or U28223 (N_28223,N_26720,N_26081);
or U28224 (N_28224,N_26463,N_25550);
nand U28225 (N_28225,N_26454,N_25606);
or U28226 (N_28226,N_26189,N_26881);
or U28227 (N_28227,N_25150,N_26506);
nand U28228 (N_28228,N_26754,N_25534);
and U28229 (N_28229,N_27195,N_26780);
xor U28230 (N_28230,N_26701,N_25662);
and U28231 (N_28231,N_25075,N_25656);
xor U28232 (N_28232,N_25993,N_26913);
xnor U28233 (N_28233,N_26716,N_27057);
and U28234 (N_28234,N_26899,N_25542);
and U28235 (N_28235,N_27151,N_27355);
or U28236 (N_28236,N_26609,N_27378);
and U28237 (N_28237,N_26325,N_26836);
or U28238 (N_28238,N_26046,N_27111);
xnor U28239 (N_28239,N_26160,N_27094);
nand U28240 (N_28240,N_25530,N_26808);
xnor U28241 (N_28241,N_25972,N_26154);
or U28242 (N_28242,N_25241,N_25198);
and U28243 (N_28243,N_25316,N_25815);
nand U28244 (N_28244,N_27265,N_25572);
and U28245 (N_28245,N_26495,N_26544);
or U28246 (N_28246,N_25297,N_27108);
nor U28247 (N_28247,N_26426,N_25361);
or U28248 (N_28248,N_26496,N_25977);
nand U28249 (N_28249,N_26401,N_26737);
or U28250 (N_28250,N_26201,N_26373);
xnor U28251 (N_28251,N_25106,N_25244);
or U28252 (N_28252,N_26835,N_26280);
and U28253 (N_28253,N_25820,N_26389);
nand U28254 (N_28254,N_25485,N_25965);
xnor U28255 (N_28255,N_26370,N_26487);
nor U28256 (N_28256,N_25551,N_26256);
or U28257 (N_28257,N_25302,N_25463);
nand U28258 (N_28258,N_25523,N_26602);
xnor U28259 (N_28259,N_26530,N_25411);
and U28260 (N_28260,N_26376,N_27422);
nand U28261 (N_28261,N_25629,N_27406);
and U28262 (N_28262,N_26731,N_26709);
xor U28263 (N_28263,N_25979,N_27436);
or U28264 (N_28264,N_26432,N_26298);
or U28265 (N_28265,N_26877,N_27239);
and U28266 (N_28266,N_26650,N_26362);
and U28267 (N_28267,N_25405,N_26884);
and U28268 (N_28268,N_25272,N_25814);
nand U28269 (N_28269,N_25962,N_26240);
xnor U28270 (N_28270,N_25295,N_26042);
xor U28271 (N_28271,N_26816,N_25156);
nand U28272 (N_28272,N_26273,N_26763);
nor U28273 (N_28273,N_25558,N_26923);
or U28274 (N_28274,N_26764,N_25289);
nand U28275 (N_28275,N_27476,N_26870);
xnor U28276 (N_28276,N_27384,N_26753);
xor U28277 (N_28277,N_26550,N_25881);
xnor U28278 (N_28278,N_26385,N_25590);
xnor U28279 (N_28279,N_25689,N_27128);
nand U28280 (N_28280,N_25490,N_25164);
or U28281 (N_28281,N_27163,N_25635);
nand U28282 (N_28282,N_26034,N_27250);
xor U28283 (N_28283,N_25506,N_25015);
xor U28284 (N_28284,N_25115,N_26676);
or U28285 (N_28285,N_26916,N_27351);
or U28286 (N_28286,N_27285,N_26727);
nand U28287 (N_28287,N_26330,N_25974);
or U28288 (N_28288,N_25683,N_27399);
nor U28289 (N_28289,N_27486,N_26832);
nor U28290 (N_28290,N_25303,N_25721);
xor U28291 (N_28291,N_26482,N_25223);
nand U28292 (N_28292,N_25100,N_26402);
xor U28293 (N_28293,N_26353,N_25889);
or U28294 (N_28294,N_26056,N_27348);
or U28295 (N_28295,N_25714,N_27432);
nand U28296 (N_28296,N_26344,N_25751);
and U28297 (N_28297,N_26060,N_26906);
nand U28298 (N_28298,N_27440,N_26710);
xor U28299 (N_28299,N_25522,N_26573);
xor U28300 (N_28300,N_25595,N_26744);
or U28301 (N_28301,N_27248,N_26749);
xnor U28302 (N_28302,N_26188,N_27217);
nor U28303 (N_28303,N_26564,N_26558);
nor U28304 (N_28304,N_26323,N_27186);
or U28305 (N_28305,N_25238,N_26167);
nor U28306 (N_28306,N_26437,N_26232);
or U28307 (N_28307,N_25709,N_25069);
or U28308 (N_28308,N_25880,N_26152);
and U28309 (N_28309,N_25306,N_26689);
nor U28310 (N_28310,N_25811,N_26793);
nor U28311 (N_28311,N_25199,N_27488);
or U28312 (N_28312,N_25654,N_25692);
nor U28313 (N_28313,N_26955,N_26262);
nand U28314 (N_28314,N_26568,N_26597);
xnor U28315 (N_28315,N_25917,N_26538);
nor U28316 (N_28316,N_26063,N_27224);
nor U28317 (N_28317,N_25201,N_26058);
xnor U28318 (N_28318,N_25800,N_27468);
xnor U28319 (N_28319,N_25887,N_26623);
nand U28320 (N_28320,N_26095,N_25210);
xor U28321 (N_28321,N_25335,N_25788);
xnor U28322 (N_28322,N_27204,N_25181);
and U28323 (N_28323,N_26628,N_26505);
nand U28324 (N_28324,N_25446,N_26537);
xor U28325 (N_28325,N_27118,N_25737);
and U28326 (N_28326,N_26163,N_26304);
nand U28327 (N_28327,N_25836,N_26390);
or U28328 (N_28328,N_25391,N_25286);
xnor U28329 (N_28329,N_27398,N_26950);
nor U28330 (N_28330,N_26474,N_27329);
nand U28331 (N_28331,N_27381,N_26032);
xor U28332 (N_28332,N_25010,N_26281);
xor U28333 (N_28333,N_25528,N_27361);
and U28334 (N_28334,N_25151,N_26349);
or U28335 (N_28335,N_25913,N_25371);
or U28336 (N_28336,N_25167,N_27456);
and U28337 (N_28337,N_26278,N_25144);
and U28338 (N_28338,N_27184,N_27469);
nor U28339 (N_28339,N_25254,N_25702);
xnor U28340 (N_28340,N_26723,N_26601);
xor U28341 (N_28341,N_27082,N_26148);
nand U28342 (N_28342,N_27066,N_25931);
nand U28343 (N_28343,N_25749,N_26651);
nand U28344 (N_28344,N_26443,N_26965);
nor U28345 (N_28345,N_26357,N_26824);
nand U28346 (N_28346,N_25611,N_26118);
and U28347 (N_28347,N_25732,N_27049);
and U28348 (N_28348,N_25064,N_25175);
nand U28349 (N_28349,N_25087,N_25728);
nand U28350 (N_28350,N_26719,N_26765);
and U28351 (N_28351,N_27273,N_26626);
nand U28352 (N_28352,N_27172,N_25431);
xor U28353 (N_28353,N_26595,N_26910);
nand U28354 (N_28354,N_25257,N_27258);
xor U28355 (N_28355,N_25496,N_27175);
xnor U28356 (N_28356,N_27036,N_25061);
or U28357 (N_28357,N_25136,N_27218);
nand U28358 (N_28358,N_26646,N_25840);
nor U28359 (N_28359,N_26738,N_26705);
nor U28360 (N_28360,N_25263,N_26266);
and U28361 (N_28361,N_27333,N_27321);
xnor U28362 (N_28362,N_25102,N_27372);
or U28363 (N_28363,N_26314,N_25883);
nor U28364 (N_28364,N_25469,N_25681);
xnor U28365 (N_28365,N_26229,N_25313);
nand U28366 (N_28366,N_27349,N_26688);
nand U28367 (N_28367,N_25441,N_25578);
xnor U28368 (N_28368,N_25910,N_25932);
nor U28369 (N_28369,N_25641,N_26059);
or U28370 (N_28370,N_25999,N_27325);
nor U28371 (N_28371,N_27012,N_25409);
and U28372 (N_28372,N_26801,N_25955);
nor U28373 (N_28373,N_26038,N_25449);
nor U28374 (N_28374,N_25278,N_25099);
nand U28375 (N_28375,N_26093,N_27141);
and U28376 (N_28376,N_26662,N_25617);
nand U28377 (N_28377,N_25705,N_27064);
xnor U28378 (N_28378,N_26641,N_27261);
xor U28379 (N_28379,N_26018,N_26242);
and U28380 (N_28380,N_26797,N_26554);
xnor U28381 (N_28381,N_25211,N_26318);
nor U28382 (N_28382,N_25406,N_26354);
and U28383 (N_28383,N_25011,N_25712);
and U28384 (N_28384,N_25554,N_25445);
nor U28385 (N_28385,N_26221,N_26045);
nor U28386 (N_28386,N_25348,N_27473);
or U28387 (N_28387,N_25953,N_26759);
or U28388 (N_28388,N_27330,N_26678);
nor U28389 (N_28389,N_25779,N_26271);
xnor U28390 (N_28390,N_25256,N_27028);
nand U28391 (N_28391,N_25659,N_27169);
nand U28392 (N_28392,N_26128,N_25752);
nor U28393 (N_28393,N_26348,N_25875);
xor U28394 (N_28394,N_25908,N_26519);
xor U28395 (N_28395,N_26172,N_25846);
or U28396 (N_28396,N_25872,N_25582);
nand U28397 (N_28397,N_25929,N_26656);
nand U28398 (N_28398,N_25187,N_26848);
nand U28399 (N_28399,N_25242,N_27076);
nand U28400 (N_28400,N_25058,N_26898);
and U28401 (N_28401,N_26241,N_26920);
nor U28402 (N_28402,N_27072,N_26509);
nand U28403 (N_28403,N_25900,N_25945);
xor U28404 (N_28404,N_25684,N_25956);
or U28405 (N_28405,N_26460,N_25829);
nand U28406 (N_28406,N_26745,N_25275);
nor U28407 (N_28407,N_25675,N_26085);
xnor U28408 (N_28408,N_25919,N_27457);
nand U28409 (N_28409,N_25750,N_27485);
xnor U28410 (N_28410,N_26739,N_26642);
and U28411 (N_28411,N_26342,N_25844);
nor U28412 (N_28412,N_26513,N_25352);
or U28413 (N_28413,N_27131,N_27209);
nor U28414 (N_28414,N_25627,N_25553);
nand U28415 (N_28415,N_26876,N_26308);
nor U28416 (N_28416,N_26054,N_25132);
nand U28417 (N_28417,N_26904,N_25677);
nand U28418 (N_28418,N_26922,N_26661);
and U28419 (N_28419,N_27197,N_26875);
or U28420 (N_28420,N_26938,N_26473);
or U28421 (N_28421,N_26053,N_25864);
xor U28422 (N_28422,N_27498,N_25901);
xor U28423 (N_28423,N_26761,N_25349);
xor U28424 (N_28424,N_26322,N_26596);
nor U28425 (N_28425,N_26000,N_25805);
and U28426 (N_28426,N_25867,N_25816);
and U28427 (N_28427,N_25047,N_27086);
or U28428 (N_28428,N_25912,N_26594);
nor U28429 (N_28429,N_26627,N_25245);
xor U28430 (N_28430,N_25250,N_27091);
or U28431 (N_28431,N_26434,N_25473);
and U28432 (N_28432,N_26111,N_27271);
or U28433 (N_28433,N_25083,N_26203);
nor U28434 (N_28434,N_27043,N_27375);
or U28435 (N_28435,N_27284,N_27235);
nand U28436 (N_28436,N_25727,N_26176);
and U28437 (N_28437,N_25842,N_26499);
xor U28438 (N_28438,N_26192,N_26074);
xnor U28439 (N_28439,N_25209,N_27023);
and U28440 (N_28440,N_27152,N_27396);
and U28441 (N_28441,N_27340,N_25914);
and U28442 (N_28442,N_27341,N_25060);
nor U28443 (N_28443,N_27236,N_26508);
nor U28444 (N_28444,N_26995,N_26517);
and U28445 (N_28445,N_25336,N_25706);
nand U28446 (N_28446,N_25249,N_25778);
xnor U28447 (N_28447,N_26476,N_25225);
nor U28448 (N_28448,N_27242,N_25007);
nor U28449 (N_28449,N_26019,N_25281);
nand U28450 (N_28450,N_27159,N_26259);
nand U28451 (N_28451,N_27206,N_26431);
nand U28452 (N_28452,N_25495,N_26940);
or U28453 (N_28453,N_25062,N_25208);
nand U28454 (N_28454,N_26049,N_26733);
xnor U28455 (N_28455,N_26155,N_25161);
and U28456 (N_28456,N_25147,N_25089);
xnor U28457 (N_28457,N_26894,N_27032);
or U28458 (N_28458,N_27150,N_25909);
xnor U28459 (N_28459,N_25850,N_27170);
xnor U28460 (N_28460,N_25798,N_25401);
or U28461 (N_28461,N_25810,N_25005);
and U28462 (N_28462,N_27037,N_27157);
or U28463 (N_28463,N_27373,N_26124);
nand U28464 (N_28464,N_25480,N_27215);
and U28465 (N_28465,N_25127,N_25694);
nand U28466 (N_28466,N_26015,N_27177);
or U28467 (N_28467,N_27481,N_25994);
xnor U28468 (N_28468,N_26633,N_25618);
nor U28469 (N_28469,N_27026,N_25926);
and U28470 (N_28470,N_26905,N_26794);
nand U28471 (N_28471,N_27345,N_26956);
xor U28472 (N_28472,N_25893,N_26295);
xor U28473 (N_28473,N_25073,N_26010);
or U28474 (N_28474,N_25561,N_25624);
and U28475 (N_28475,N_26350,N_26387);
nor U28476 (N_28476,N_25903,N_25190);
and U28477 (N_28477,N_26750,N_26787);
or U28478 (N_28478,N_27302,N_26696);
and U28479 (N_28479,N_26433,N_25934);
nor U28480 (N_28480,N_25018,N_25460);
nor U28481 (N_28481,N_25462,N_27002);
nand U28482 (N_28482,N_25410,N_25280);
xnor U28483 (N_28483,N_26022,N_25400);
or U28484 (N_28484,N_26236,N_26643);
nand U28485 (N_28485,N_26157,N_25748);
xor U28486 (N_28486,N_25299,N_26235);
or U28487 (N_28487,N_26924,N_26427);
or U28488 (N_28488,N_26865,N_25327);
or U28489 (N_28489,N_25240,N_25575);
nand U28490 (N_28490,N_27025,N_25782);
or U28491 (N_28491,N_27419,N_27226);
or U28492 (N_28492,N_25717,N_26494);
nor U28493 (N_28493,N_26523,N_25375);
xor U28494 (N_28494,N_25487,N_26700);
or U28495 (N_28495,N_27289,N_26416);
nor U28496 (N_28496,N_27105,N_25447);
or U28497 (N_28497,N_25568,N_26992);
nand U28498 (N_28498,N_26372,N_25004);
xor U28499 (N_28499,N_27174,N_25436);
and U28500 (N_28500,N_25159,N_27038);
nor U28501 (N_28501,N_26268,N_25027);
or U28502 (N_28502,N_25845,N_25518);
and U28503 (N_28503,N_26324,N_26864);
and U28504 (N_28504,N_26712,N_27407);
and U28505 (N_28505,N_25785,N_25051);
xnor U28506 (N_28506,N_25527,N_25055);
nor U28507 (N_28507,N_26774,N_25196);
and U28508 (N_28508,N_26632,N_27335);
nand U28509 (N_28509,N_26684,N_25902);
xor U28510 (N_28510,N_25216,N_26614);
nand U28511 (N_28511,N_26419,N_26169);
and U28512 (N_28512,N_27332,N_26647);
nor U28513 (N_28513,N_26200,N_26466);
nor U28514 (N_28514,N_25638,N_27182);
xor U28515 (N_28515,N_25789,N_26805);
or U28516 (N_28516,N_25085,N_27410);
nor U28517 (N_28517,N_25587,N_25687);
xnor U28518 (N_28518,N_27463,N_26024);
or U28519 (N_28519,N_25079,N_26796);
nor U28520 (N_28520,N_26722,N_26873);
and U28521 (N_28521,N_25356,N_26008);
nor U28522 (N_28522,N_26590,N_25368);
nand U28523 (N_28523,N_26552,N_27479);
nand U28524 (N_28524,N_26340,N_25874);
xnor U28525 (N_28525,N_26612,N_26139);
or U28526 (N_28526,N_25743,N_26671);
xnor U28527 (N_28527,N_27060,N_26267);
nor U28528 (N_28528,N_26395,N_26098);
or U28529 (N_28529,N_27427,N_26504);
or U28530 (N_28530,N_26510,N_26497);
xor U28531 (N_28531,N_26886,N_27304);
nor U28532 (N_28532,N_26980,N_25339);
nand U28533 (N_28533,N_26407,N_26619);
and U28534 (N_28534,N_26143,N_25927);
or U28535 (N_28535,N_26939,N_26946);
nand U28536 (N_28536,N_25177,N_25708);
and U28537 (N_28537,N_27347,N_27201);
nand U28538 (N_28538,N_27426,N_26131);
xnor U28539 (N_28539,N_26501,N_25787);
nor U28540 (N_28540,N_26903,N_27205);
or U28541 (N_28541,N_25000,N_25620);
xor U28542 (N_28542,N_25824,N_25038);
nand U28543 (N_28543,N_26874,N_25131);
and U28544 (N_28544,N_25232,N_26735);
xnor U28545 (N_28545,N_26413,N_25545);
and U28546 (N_28546,N_26844,N_26277);
nand U28547 (N_28547,N_25852,N_25221);
nor U28548 (N_28548,N_27444,N_26539);
nor U28549 (N_28549,N_26341,N_26825);
or U28550 (N_28550,N_25404,N_27006);
nor U28551 (N_28551,N_26984,N_25319);
and U28552 (N_28552,N_26062,N_26083);
or U28553 (N_28553,N_27394,N_25259);
nor U28554 (N_28554,N_27219,N_25764);
nor U28555 (N_28555,N_25971,N_27338);
xnor U28556 (N_28556,N_27309,N_26660);
nor U28557 (N_28557,N_25878,N_27073);
xor U28558 (N_28558,N_25017,N_25599);
xnor U28559 (N_28559,N_27241,N_27090);
nand U28560 (N_28560,N_27460,N_25337);
nor U28561 (N_28561,N_25904,N_26526);
or U28562 (N_28562,N_26756,N_25403);
nand U28563 (N_28563,N_27109,N_27296);
or U28564 (N_28564,N_27297,N_27123);
nor U28565 (N_28565,N_25711,N_25045);
nand U28566 (N_28566,N_25799,N_26179);
and U28567 (N_28567,N_25848,N_25673);
and U28568 (N_28568,N_26846,N_26439);
nor U28569 (N_28569,N_25537,N_26287);
nor U28570 (N_28570,N_26352,N_26047);
nand U28571 (N_28571,N_25646,N_26692);
or U28572 (N_28572,N_27382,N_27447);
xnor U28573 (N_28573,N_26190,N_25894);
or U28574 (N_28574,N_26255,N_25021);
nand U28575 (N_28575,N_25643,N_26773);
nand U28576 (N_28576,N_26230,N_25619);
xor U28577 (N_28577,N_27454,N_26586);
or U28578 (N_28578,N_26135,N_27213);
xor U28579 (N_28579,N_25541,N_26635);
nor U28580 (N_28580,N_27495,N_27045);
nand U28581 (N_28581,N_25155,N_26116);
nor U28582 (N_28582,N_27263,N_25969);
xnor U28583 (N_28583,N_26462,N_25531);
nor U28584 (N_28584,N_26253,N_26679);
xor U28585 (N_28585,N_25235,N_26121);
xnor U28586 (N_28586,N_25697,N_27379);
nor U28587 (N_28587,N_26747,N_26033);
nor U28588 (N_28588,N_27453,N_27024);
nand U28589 (N_28589,N_25200,N_25354);
and U28590 (N_28590,N_25631,N_26637);
or U28591 (N_28591,N_25116,N_25923);
and U28592 (N_28592,N_26227,N_26766);
nand U28593 (N_28593,N_26493,N_26307);
nand U28594 (N_28594,N_26440,N_25093);
or U28595 (N_28595,N_27425,N_26813);
xnor U28596 (N_28596,N_26077,N_26379);
or U28597 (N_28597,N_27112,N_25564);
and U28598 (N_28598,N_26800,N_25676);
or U28599 (N_28599,N_26238,N_25922);
or U28600 (N_28600,N_27132,N_27144);
and U28601 (N_28601,N_25172,N_26549);
and U28602 (N_28602,N_26276,N_27428);
xor U28603 (N_28603,N_25255,N_26762);
xor U28604 (N_28604,N_25477,N_26970);
nand U28605 (N_28605,N_25332,N_25783);
nor U28606 (N_28606,N_26717,N_27412);
xor U28607 (N_28607,N_25437,N_27160);
nor U28608 (N_28608,N_26265,N_26214);
nor U28609 (N_28609,N_26375,N_26141);
and U28610 (N_28610,N_26529,N_26112);
xnor U28611 (N_28611,N_25987,N_25921);
nand U28612 (N_28612,N_26470,N_25667);
or U28613 (N_28613,N_26613,N_26195);
nor U28614 (N_28614,N_26080,N_26611);
and U28615 (N_28615,N_26921,N_27458);
nand U28616 (N_28616,N_25381,N_27230);
nor U28617 (N_28617,N_25372,N_25995);
xor U28618 (N_28618,N_25529,N_25016);
nand U28619 (N_28619,N_26173,N_27136);
nor U28620 (N_28620,N_25510,N_25879);
or U28621 (N_28621,N_27027,N_25633);
xnor U28622 (N_28622,N_26127,N_27077);
xor U28623 (N_28623,N_26883,N_26420);
or U28624 (N_28624,N_27430,N_26346);
and U28625 (N_28625,N_25026,N_26803);
nand U28626 (N_28626,N_26193,N_27431);
xnor U28627 (N_28627,N_25600,N_26979);
xor U28628 (N_28628,N_25636,N_27356);
and U28629 (N_28629,N_25517,N_26561);
xor U28630 (N_28630,N_27264,N_25243);
nor U28631 (N_28631,N_27088,N_25933);
nor U28632 (N_28632,N_26578,N_25353);
and U28633 (N_28633,N_25362,N_25413);
or U28634 (N_28634,N_26814,N_25139);
xnor U28635 (N_28635,N_26528,N_26567);
nand U28636 (N_28636,N_27121,N_26133);
and U28637 (N_28637,N_26963,N_25796);
nand U28638 (N_28638,N_26132,N_26866);
xor U28639 (N_28639,N_26625,N_26066);
nor U28640 (N_28640,N_27474,N_27377);
nand U28641 (N_28641,N_27171,N_25346);
nand U28642 (N_28642,N_25784,N_26991);
and U28643 (N_28643,N_25650,N_27104);
and U28644 (N_28644,N_25478,N_25088);
nand U28645 (N_28645,N_26536,N_27336);
nor U28646 (N_28646,N_26383,N_26669);
and U28647 (N_28647,N_26050,N_25444);
nand U28648 (N_28648,N_25458,N_27115);
xor U28649 (N_28649,N_27392,N_26655);
nand U28650 (N_28650,N_25951,N_25860);
or U28651 (N_28651,N_26935,N_25497);
and U28652 (N_28652,N_26724,N_25341);
nand U28653 (N_28653,N_26961,N_25795);
or U28654 (N_28654,N_25440,N_25841);
nand U28655 (N_28655,N_25108,N_25696);
or U28656 (N_28656,N_26606,N_26477);
nand U28657 (N_28657,N_25248,N_25802);
or U28658 (N_28658,N_26775,N_26196);
nand U28659 (N_28659,N_26369,N_26142);
and U28660 (N_28660,N_27166,N_26423);
nor U28661 (N_28661,N_25376,N_25237);
and U28662 (N_28662,N_25084,N_26017);
or U28663 (N_28663,N_27075,N_25110);
xor U28664 (N_28664,N_27089,N_26101);
and U28665 (N_28665,N_25114,N_26243);
xor U28666 (N_28666,N_25326,N_26973);
nor U28667 (N_28667,N_26151,N_25740);
or U28668 (N_28668,N_27413,N_26428);
xnor U28669 (N_28669,N_26725,N_26182);
or U28670 (N_28670,N_27328,N_25046);
nor U28671 (N_28671,N_27047,N_26682);
or U28672 (N_28672,N_25790,N_26997);
nor U28673 (N_28673,N_25193,N_25769);
nor U28674 (N_28674,N_26275,N_26026);
nor U28675 (N_28675,N_25247,N_25765);
nand U28676 (N_28676,N_26113,N_27203);
nand U28677 (N_28677,N_26165,N_26351);
and U28678 (N_28678,N_25532,N_27229);
and U28679 (N_28679,N_27124,N_26933);
and U28680 (N_28680,N_26819,N_25876);
or U28681 (N_28681,N_27490,N_26532);
or U28682 (N_28682,N_26915,N_25267);
and U28683 (N_28683,N_25508,N_26043);
nor U28684 (N_28684,N_25424,N_25358);
and U28685 (N_28685,N_25663,N_26741);
and U28686 (N_28686,N_25762,N_27320);
nand U28687 (N_28687,N_27484,N_27441);
nand U28688 (N_28688,N_26328,N_26507);
xor U28689 (N_28689,N_27053,N_26809);
nand U28690 (N_28690,N_27317,N_27034);
nand U28691 (N_28691,N_25054,N_27275);
or U28692 (N_28692,N_27149,N_26853);
or U28693 (N_28693,N_25519,N_26778);
or U28694 (N_28694,N_25859,N_27237);
and U28695 (N_28695,N_25251,N_27445);
or U28696 (N_28696,N_26014,N_26751);
nand U28697 (N_28697,N_26768,N_25754);
and U28698 (N_28698,N_25739,N_27268);
nor U28699 (N_28699,N_26472,N_27363);
or U28700 (N_28700,N_25279,N_26770);
and U28701 (N_28701,N_25296,N_26366);
and U28702 (N_28702,N_25135,N_26580);
xor U28703 (N_28703,N_25854,N_25308);
xnor U28704 (N_28704,N_26551,N_26890);
xor U28705 (N_28705,N_25464,N_26928);
nor U28706 (N_28706,N_27466,N_27438);
or U28707 (N_28707,N_25366,N_25001);
xnor U28708 (N_28708,N_26107,N_25753);
nand U28709 (N_28709,N_25504,N_25359);
xnor U28710 (N_28710,N_25649,N_27103);
nor U28711 (N_28711,N_27233,N_25030);
xnor U28712 (N_28712,N_25941,N_25074);
or U28713 (N_28713,N_26471,N_25338);
nor U28714 (N_28714,N_26216,N_25191);
nor U28715 (N_28715,N_27362,N_26639);
nand U28716 (N_28716,N_25195,N_25838);
nand U28717 (N_28717,N_25562,N_25140);
nor U28718 (N_28718,N_26943,N_25707);
nand U28719 (N_28719,N_27487,N_25124);
or U28720 (N_28720,N_25715,N_25310);
nand U28721 (N_28721,N_26927,N_25724);
nor U28722 (N_28722,N_26478,N_26394);
xnor U28723 (N_28723,N_26442,N_26162);
or U28724 (N_28724,N_27389,N_26777);
or U28725 (N_28725,N_27364,N_26479);
and U28726 (N_28726,N_25101,N_27240);
and U28727 (N_28727,N_25350,N_26089);
and U28728 (N_28728,N_26247,N_26587);
xnor U28729 (N_28729,N_26485,N_25736);
nand U28730 (N_28730,N_27107,N_27231);
nor U28731 (N_28731,N_26585,N_27214);
nor U28732 (N_28732,N_27020,N_25035);
nand U28733 (N_28733,N_27059,N_26576);
nand U28734 (N_28734,N_25459,N_26799);
xor U28735 (N_28735,N_26175,N_25645);
nor U28736 (N_28736,N_26821,N_25704);
or U28737 (N_28737,N_25188,N_25126);
or U28738 (N_28738,N_25610,N_26177);
xnor U28739 (N_28739,N_27334,N_25937);
or U28740 (N_28740,N_25340,N_25756);
nor U28741 (N_28741,N_25525,N_25176);
xor U28742 (N_28742,N_27346,N_27014);
nand U28743 (N_28743,N_25033,N_25943);
or U28744 (N_28744,N_25985,N_27391);
nand U28745 (N_28745,N_26556,N_27464);
and U28746 (N_28746,N_25421,N_25801);
xor U28747 (N_28747,N_25920,N_25494);
or U28748 (N_28748,N_27397,N_25091);
or U28749 (N_28749,N_26993,N_26016);
or U28750 (N_28750,N_26988,N_26015);
and U28751 (N_28751,N_25639,N_25859);
or U28752 (N_28752,N_25630,N_25868);
nor U28753 (N_28753,N_25695,N_27089);
and U28754 (N_28754,N_25998,N_27357);
nand U28755 (N_28755,N_27110,N_27011);
nor U28756 (N_28756,N_26328,N_27323);
xnor U28757 (N_28757,N_25741,N_25363);
xor U28758 (N_28758,N_26589,N_26463);
or U28759 (N_28759,N_25247,N_27312);
xor U28760 (N_28760,N_25902,N_27366);
xor U28761 (N_28761,N_26356,N_25527);
nand U28762 (N_28762,N_27129,N_25596);
xnor U28763 (N_28763,N_25515,N_26928);
and U28764 (N_28764,N_27353,N_25640);
and U28765 (N_28765,N_26660,N_25151);
nor U28766 (N_28766,N_27155,N_26260);
xor U28767 (N_28767,N_26732,N_25002);
nor U28768 (N_28768,N_26071,N_25023);
and U28769 (N_28769,N_25293,N_25423);
or U28770 (N_28770,N_27478,N_26641);
nor U28771 (N_28771,N_26725,N_25829);
nor U28772 (N_28772,N_27438,N_26228);
xor U28773 (N_28773,N_26521,N_27499);
xor U28774 (N_28774,N_25809,N_27247);
xor U28775 (N_28775,N_25657,N_25845);
or U28776 (N_28776,N_26633,N_26868);
nor U28777 (N_28777,N_26181,N_25752);
nand U28778 (N_28778,N_26485,N_25817);
xnor U28779 (N_28779,N_25103,N_26951);
nand U28780 (N_28780,N_25265,N_25828);
nand U28781 (N_28781,N_25826,N_26833);
nor U28782 (N_28782,N_27036,N_25555);
xnor U28783 (N_28783,N_26216,N_25697);
or U28784 (N_28784,N_26311,N_27109);
xor U28785 (N_28785,N_27238,N_25334);
nand U28786 (N_28786,N_25020,N_26478);
nor U28787 (N_28787,N_26695,N_27448);
or U28788 (N_28788,N_26418,N_26015);
or U28789 (N_28789,N_25989,N_26604);
nor U28790 (N_28790,N_27311,N_25854);
nand U28791 (N_28791,N_26098,N_27286);
xnor U28792 (N_28792,N_26314,N_26456);
nand U28793 (N_28793,N_25566,N_27148);
or U28794 (N_28794,N_26143,N_25718);
nand U28795 (N_28795,N_25367,N_27166);
and U28796 (N_28796,N_25432,N_25010);
nand U28797 (N_28797,N_27274,N_26917);
and U28798 (N_28798,N_25295,N_27023);
and U28799 (N_28799,N_26075,N_25801);
and U28800 (N_28800,N_27019,N_27469);
or U28801 (N_28801,N_26507,N_25394);
or U28802 (N_28802,N_27150,N_26403);
and U28803 (N_28803,N_27364,N_27008);
nor U28804 (N_28804,N_26959,N_27054);
or U28805 (N_28805,N_25281,N_25870);
nor U28806 (N_28806,N_25149,N_27254);
and U28807 (N_28807,N_25274,N_25641);
nor U28808 (N_28808,N_27092,N_26247);
or U28809 (N_28809,N_26369,N_26751);
and U28810 (N_28810,N_25100,N_26369);
or U28811 (N_28811,N_25973,N_25775);
or U28812 (N_28812,N_26528,N_26780);
nand U28813 (N_28813,N_25764,N_25954);
xnor U28814 (N_28814,N_26963,N_25457);
xor U28815 (N_28815,N_26705,N_25930);
or U28816 (N_28816,N_27418,N_25489);
xor U28817 (N_28817,N_26425,N_26103);
and U28818 (N_28818,N_25623,N_26492);
nand U28819 (N_28819,N_25627,N_25882);
xor U28820 (N_28820,N_25393,N_25205);
and U28821 (N_28821,N_25731,N_26306);
and U28822 (N_28822,N_25337,N_27249);
or U28823 (N_28823,N_27460,N_26493);
nor U28824 (N_28824,N_25500,N_25588);
nor U28825 (N_28825,N_26624,N_27371);
nor U28826 (N_28826,N_27432,N_26949);
and U28827 (N_28827,N_25401,N_25999);
or U28828 (N_28828,N_25801,N_25470);
xnor U28829 (N_28829,N_27068,N_26121);
and U28830 (N_28830,N_25531,N_25654);
nand U28831 (N_28831,N_26460,N_26006);
nor U28832 (N_28832,N_27162,N_27120);
nand U28833 (N_28833,N_26456,N_27289);
or U28834 (N_28834,N_27027,N_26009);
nor U28835 (N_28835,N_27139,N_26516);
nor U28836 (N_28836,N_25624,N_25712);
or U28837 (N_28837,N_26082,N_25606);
and U28838 (N_28838,N_25954,N_25127);
nand U28839 (N_28839,N_25665,N_27394);
nand U28840 (N_28840,N_25719,N_25817);
and U28841 (N_28841,N_26848,N_25936);
or U28842 (N_28842,N_26415,N_26259);
xnor U28843 (N_28843,N_25468,N_27270);
nand U28844 (N_28844,N_27177,N_27121);
nand U28845 (N_28845,N_27282,N_27107);
or U28846 (N_28846,N_26677,N_25911);
or U28847 (N_28847,N_25314,N_25731);
xor U28848 (N_28848,N_25205,N_26505);
xnor U28849 (N_28849,N_27002,N_25171);
xnor U28850 (N_28850,N_26176,N_26720);
and U28851 (N_28851,N_25292,N_26036);
and U28852 (N_28852,N_25425,N_25250);
xor U28853 (N_28853,N_26257,N_25581);
nor U28854 (N_28854,N_26003,N_25479);
and U28855 (N_28855,N_25771,N_27341);
xor U28856 (N_28856,N_25725,N_26688);
nand U28857 (N_28857,N_26309,N_27148);
nand U28858 (N_28858,N_26022,N_25101);
or U28859 (N_28859,N_25872,N_26985);
and U28860 (N_28860,N_26279,N_26177);
or U28861 (N_28861,N_25623,N_26974);
and U28862 (N_28862,N_26188,N_25429);
nor U28863 (N_28863,N_25947,N_26881);
or U28864 (N_28864,N_27314,N_25461);
and U28865 (N_28865,N_27363,N_26270);
and U28866 (N_28866,N_27271,N_26902);
nor U28867 (N_28867,N_25978,N_25666);
or U28868 (N_28868,N_25303,N_26527);
and U28869 (N_28869,N_26011,N_26783);
and U28870 (N_28870,N_27267,N_27329);
xor U28871 (N_28871,N_26700,N_25238);
or U28872 (N_28872,N_26163,N_26948);
xor U28873 (N_28873,N_27005,N_27294);
nand U28874 (N_28874,N_27475,N_25821);
nand U28875 (N_28875,N_27395,N_25369);
and U28876 (N_28876,N_27127,N_25392);
nor U28877 (N_28877,N_26977,N_27364);
or U28878 (N_28878,N_25400,N_26379);
nor U28879 (N_28879,N_25222,N_27056);
xnor U28880 (N_28880,N_26011,N_27451);
and U28881 (N_28881,N_25151,N_25587);
or U28882 (N_28882,N_26250,N_27167);
or U28883 (N_28883,N_26440,N_25489);
nor U28884 (N_28884,N_26063,N_26815);
and U28885 (N_28885,N_25354,N_26321);
or U28886 (N_28886,N_26525,N_26166);
nand U28887 (N_28887,N_25228,N_26404);
nor U28888 (N_28888,N_26921,N_26102);
or U28889 (N_28889,N_26887,N_26970);
or U28890 (N_28890,N_27246,N_25263);
and U28891 (N_28891,N_25356,N_25267);
nor U28892 (N_28892,N_25683,N_25413);
xnor U28893 (N_28893,N_26733,N_25186);
or U28894 (N_28894,N_25860,N_26331);
xnor U28895 (N_28895,N_26194,N_25373);
nand U28896 (N_28896,N_26114,N_27153);
nand U28897 (N_28897,N_26779,N_25907);
nand U28898 (N_28898,N_27348,N_25284);
or U28899 (N_28899,N_25909,N_25965);
and U28900 (N_28900,N_25375,N_26526);
and U28901 (N_28901,N_25401,N_25815);
nand U28902 (N_28902,N_26500,N_26012);
nor U28903 (N_28903,N_25128,N_25415);
and U28904 (N_28904,N_25667,N_26749);
and U28905 (N_28905,N_25694,N_25586);
xor U28906 (N_28906,N_26826,N_25766);
or U28907 (N_28907,N_26065,N_26133);
xnor U28908 (N_28908,N_26902,N_26925);
or U28909 (N_28909,N_25611,N_26990);
xor U28910 (N_28910,N_26880,N_25776);
and U28911 (N_28911,N_26788,N_25617);
xor U28912 (N_28912,N_26051,N_25481);
and U28913 (N_28913,N_26884,N_27008);
nor U28914 (N_28914,N_25601,N_26809);
nor U28915 (N_28915,N_25641,N_26071);
or U28916 (N_28916,N_27094,N_26257);
and U28917 (N_28917,N_27421,N_25075);
or U28918 (N_28918,N_25645,N_25640);
nand U28919 (N_28919,N_26341,N_27244);
and U28920 (N_28920,N_26745,N_26102);
and U28921 (N_28921,N_26966,N_25143);
and U28922 (N_28922,N_26681,N_26413);
or U28923 (N_28923,N_26646,N_26865);
or U28924 (N_28924,N_25527,N_26236);
and U28925 (N_28925,N_25881,N_26224);
nor U28926 (N_28926,N_27482,N_26249);
xor U28927 (N_28927,N_25526,N_26511);
nor U28928 (N_28928,N_26967,N_25807);
xor U28929 (N_28929,N_25553,N_25208);
nand U28930 (N_28930,N_25350,N_26818);
or U28931 (N_28931,N_26888,N_27080);
or U28932 (N_28932,N_26508,N_25190);
nor U28933 (N_28933,N_26587,N_25181);
or U28934 (N_28934,N_25204,N_26515);
nor U28935 (N_28935,N_26273,N_25159);
nor U28936 (N_28936,N_27375,N_26668);
xnor U28937 (N_28937,N_27188,N_26165);
or U28938 (N_28938,N_26919,N_26929);
xnor U28939 (N_28939,N_26999,N_25852);
nor U28940 (N_28940,N_26422,N_25613);
nand U28941 (N_28941,N_25738,N_25793);
xor U28942 (N_28942,N_25539,N_26189);
nand U28943 (N_28943,N_27262,N_26015);
or U28944 (N_28944,N_25623,N_26742);
xnor U28945 (N_28945,N_25413,N_27447);
nand U28946 (N_28946,N_27270,N_27326);
nor U28947 (N_28947,N_26549,N_27175);
nand U28948 (N_28948,N_26055,N_26390);
xnor U28949 (N_28949,N_26638,N_26916);
nand U28950 (N_28950,N_26135,N_25928);
or U28951 (N_28951,N_25473,N_26331);
nor U28952 (N_28952,N_26913,N_25052);
nor U28953 (N_28953,N_25118,N_26559);
or U28954 (N_28954,N_26639,N_27115);
nand U28955 (N_28955,N_25554,N_27494);
xnor U28956 (N_28956,N_26166,N_27363);
or U28957 (N_28957,N_27445,N_26642);
xnor U28958 (N_28958,N_26998,N_25150);
nor U28959 (N_28959,N_26325,N_27488);
nand U28960 (N_28960,N_26546,N_27408);
nand U28961 (N_28961,N_26464,N_26803);
nor U28962 (N_28962,N_26608,N_27124);
nand U28963 (N_28963,N_27383,N_27001);
nand U28964 (N_28964,N_26513,N_26792);
or U28965 (N_28965,N_26829,N_27341);
or U28966 (N_28966,N_26368,N_26629);
or U28967 (N_28967,N_25926,N_25568);
xor U28968 (N_28968,N_25223,N_25109);
xnor U28969 (N_28969,N_25641,N_26103);
or U28970 (N_28970,N_26776,N_25626);
nor U28971 (N_28971,N_26634,N_25350);
or U28972 (N_28972,N_25600,N_25340);
or U28973 (N_28973,N_26748,N_25851);
or U28974 (N_28974,N_26444,N_26816);
xnor U28975 (N_28975,N_25105,N_25544);
or U28976 (N_28976,N_25242,N_25521);
xnor U28977 (N_28977,N_26603,N_25147);
and U28978 (N_28978,N_25255,N_26769);
nor U28979 (N_28979,N_25134,N_25626);
or U28980 (N_28980,N_25228,N_26362);
or U28981 (N_28981,N_26289,N_27021);
nor U28982 (N_28982,N_27193,N_25775);
xor U28983 (N_28983,N_27153,N_27468);
nor U28984 (N_28984,N_25282,N_26319);
or U28985 (N_28985,N_26667,N_26906);
and U28986 (N_28986,N_26192,N_26827);
xnor U28987 (N_28987,N_26854,N_27118);
xnor U28988 (N_28988,N_25533,N_26865);
nor U28989 (N_28989,N_26207,N_26024);
and U28990 (N_28990,N_25980,N_26848);
nor U28991 (N_28991,N_27170,N_27427);
nor U28992 (N_28992,N_27405,N_26171);
or U28993 (N_28993,N_25223,N_26167);
xor U28994 (N_28994,N_25417,N_25097);
xnor U28995 (N_28995,N_27184,N_25652);
and U28996 (N_28996,N_25187,N_26075);
or U28997 (N_28997,N_26048,N_25204);
or U28998 (N_28998,N_25497,N_26257);
and U28999 (N_28999,N_25774,N_27473);
nor U29000 (N_29000,N_25253,N_26524);
xnor U29001 (N_29001,N_25387,N_25973);
xnor U29002 (N_29002,N_26546,N_27372);
nor U29003 (N_29003,N_27238,N_26777);
xnor U29004 (N_29004,N_27379,N_26392);
nor U29005 (N_29005,N_25640,N_25111);
nand U29006 (N_29006,N_26262,N_27064);
and U29007 (N_29007,N_25752,N_27124);
and U29008 (N_29008,N_27060,N_26547);
nor U29009 (N_29009,N_25126,N_25809);
nor U29010 (N_29010,N_25800,N_26477);
xnor U29011 (N_29011,N_25133,N_26815);
and U29012 (N_29012,N_26786,N_26261);
nor U29013 (N_29013,N_25669,N_26808);
and U29014 (N_29014,N_26417,N_25565);
nand U29015 (N_29015,N_25167,N_26403);
nor U29016 (N_29016,N_27309,N_25274);
and U29017 (N_29017,N_26395,N_26352);
nand U29018 (N_29018,N_25498,N_26191);
or U29019 (N_29019,N_27086,N_25138);
xor U29020 (N_29020,N_25277,N_27053);
and U29021 (N_29021,N_25255,N_25150);
nand U29022 (N_29022,N_25949,N_26835);
or U29023 (N_29023,N_26442,N_26268);
nor U29024 (N_29024,N_26498,N_25406);
and U29025 (N_29025,N_27143,N_25937);
nand U29026 (N_29026,N_27406,N_26993);
xor U29027 (N_29027,N_25289,N_27127);
nor U29028 (N_29028,N_27123,N_25413);
and U29029 (N_29029,N_25664,N_25160);
xor U29030 (N_29030,N_26723,N_26896);
nor U29031 (N_29031,N_27088,N_26053);
nor U29032 (N_29032,N_27411,N_25223);
or U29033 (N_29033,N_26842,N_27436);
nor U29034 (N_29034,N_26629,N_26091);
and U29035 (N_29035,N_26571,N_26220);
xnor U29036 (N_29036,N_27065,N_27283);
nor U29037 (N_29037,N_25568,N_25804);
or U29038 (N_29038,N_25817,N_27264);
and U29039 (N_29039,N_27499,N_25476);
xor U29040 (N_29040,N_27428,N_25119);
nand U29041 (N_29041,N_27326,N_25180);
nor U29042 (N_29042,N_25320,N_25939);
xnor U29043 (N_29043,N_25270,N_26164);
and U29044 (N_29044,N_25266,N_26964);
nand U29045 (N_29045,N_26551,N_26610);
nor U29046 (N_29046,N_25727,N_25830);
and U29047 (N_29047,N_26597,N_26452);
and U29048 (N_29048,N_26163,N_27427);
or U29049 (N_29049,N_25094,N_25237);
nand U29050 (N_29050,N_26884,N_25410);
nor U29051 (N_29051,N_25168,N_26085);
nand U29052 (N_29052,N_25829,N_26193);
nor U29053 (N_29053,N_27210,N_26684);
nand U29054 (N_29054,N_26850,N_26216);
xor U29055 (N_29055,N_25338,N_25085);
nor U29056 (N_29056,N_26137,N_25518);
or U29057 (N_29057,N_25588,N_26375);
or U29058 (N_29058,N_27025,N_25926);
xor U29059 (N_29059,N_27376,N_27051);
nand U29060 (N_29060,N_26199,N_25390);
xor U29061 (N_29061,N_25322,N_27458);
nand U29062 (N_29062,N_25382,N_26530);
nor U29063 (N_29063,N_25567,N_25598);
nand U29064 (N_29064,N_26436,N_25544);
or U29065 (N_29065,N_26432,N_26737);
nor U29066 (N_29066,N_25029,N_25543);
or U29067 (N_29067,N_26893,N_26298);
nand U29068 (N_29068,N_27171,N_26701);
nand U29069 (N_29069,N_25237,N_25284);
and U29070 (N_29070,N_25525,N_26905);
xor U29071 (N_29071,N_26687,N_27059);
and U29072 (N_29072,N_25249,N_25666);
xnor U29073 (N_29073,N_25020,N_26553);
or U29074 (N_29074,N_26405,N_25114);
and U29075 (N_29075,N_25449,N_26526);
and U29076 (N_29076,N_27443,N_26239);
nor U29077 (N_29077,N_25743,N_25284);
nand U29078 (N_29078,N_26668,N_26184);
xnor U29079 (N_29079,N_27424,N_26089);
xnor U29080 (N_29080,N_25740,N_26611);
or U29081 (N_29081,N_25925,N_25269);
nor U29082 (N_29082,N_25937,N_27154);
and U29083 (N_29083,N_26715,N_25582);
nor U29084 (N_29084,N_26738,N_27014);
nand U29085 (N_29085,N_25263,N_25863);
xnor U29086 (N_29086,N_25699,N_27181);
nor U29087 (N_29087,N_26999,N_25769);
xnor U29088 (N_29088,N_26277,N_25195);
and U29089 (N_29089,N_27391,N_27173);
or U29090 (N_29090,N_25844,N_26127);
xnor U29091 (N_29091,N_26831,N_26400);
nand U29092 (N_29092,N_26100,N_27312);
and U29093 (N_29093,N_26843,N_26641);
nand U29094 (N_29094,N_25865,N_25352);
nor U29095 (N_29095,N_25952,N_27253);
nor U29096 (N_29096,N_25940,N_26796);
xnor U29097 (N_29097,N_27179,N_27395);
xor U29098 (N_29098,N_26461,N_26156);
and U29099 (N_29099,N_27270,N_25822);
and U29100 (N_29100,N_26283,N_26152);
nand U29101 (N_29101,N_26174,N_26502);
and U29102 (N_29102,N_26454,N_25878);
and U29103 (N_29103,N_25522,N_26879);
nand U29104 (N_29104,N_27046,N_25588);
nand U29105 (N_29105,N_25032,N_27044);
nor U29106 (N_29106,N_25426,N_27193);
nand U29107 (N_29107,N_26907,N_26836);
and U29108 (N_29108,N_25505,N_26769);
nand U29109 (N_29109,N_27288,N_25097);
or U29110 (N_29110,N_25329,N_27347);
and U29111 (N_29111,N_26639,N_25868);
xnor U29112 (N_29112,N_25044,N_25813);
nor U29113 (N_29113,N_26277,N_27365);
nand U29114 (N_29114,N_26568,N_25411);
nor U29115 (N_29115,N_27224,N_27339);
nor U29116 (N_29116,N_26517,N_26685);
xnor U29117 (N_29117,N_25138,N_26240);
nand U29118 (N_29118,N_26756,N_26036);
or U29119 (N_29119,N_27226,N_26844);
nand U29120 (N_29120,N_27303,N_25759);
nor U29121 (N_29121,N_27221,N_26744);
and U29122 (N_29122,N_25300,N_27036);
or U29123 (N_29123,N_25665,N_25932);
nand U29124 (N_29124,N_25820,N_25933);
xor U29125 (N_29125,N_26926,N_27246);
nand U29126 (N_29126,N_26118,N_26716);
xnor U29127 (N_29127,N_27350,N_25588);
nand U29128 (N_29128,N_26934,N_27003);
and U29129 (N_29129,N_26202,N_25429);
xnor U29130 (N_29130,N_27163,N_25334);
or U29131 (N_29131,N_25019,N_26879);
and U29132 (N_29132,N_26518,N_26334);
xor U29133 (N_29133,N_27082,N_25707);
xor U29134 (N_29134,N_26342,N_26083);
or U29135 (N_29135,N_26879,N_26356);
nand U29136 (N_29136,N_25353,N_25202);
nand U29137 (N_29137,N_25158,N_25952);
nand U29138 (N_29138,N_26961,N_26779);
or U29139 (N_29139,N_25604,N_25987);
or U29140 (N_29140,N_26228,N_25864);
and U29141 (N_29141,N_26693,N_27104);
nand U29142 (N_29142,N_26649,N_25124);
nand U29143 (N_29143,N_25397,N_26113);
or U29144 (N_29144,N_25231,N_25152);
xor U29145 (N_29145,N_25748,N_27489);
nor U29146 (N_29146,N_26189,N_26712);
and U29147 (N_29147,N_25321,N_26770);
or U29148 (N_29148,N_26759,N_25918);
nand U29149 (N_29149,N_25842,N_27309);
nand U29150 (N_29150,N_25941,N_26036);
nand U29151 (N_29151,N_25557,N_26040);
nand U29152 (N_29152,N_26947,N_26688);
or U29153 (N_29153,N_26726,N_26388);
nand U29154 (N_29154,N_26546,N_25890);
and U29155 (N_29155,N_25752,N_25101);
xor U29156 (N_29156,N_25182,N_26404);
or U29157 (N_29157,N_27005,N_27213);
and U29158 (N_29158,N_27484,N_27376);
or U29159 (N_29159,N_27310,N_27232);
and U29160 (N_29160,N_26245,N_27227);
nor U29161 (N_29161,N_26259,N_27123);
and U29162 (N_29162,N_25257,N_27342);
xnor U29163 (N_29163,N_25133,N_27413);
nand U29164 (N_29164,N_25825,N_26600);
nor U29165 (N_29165,N_26218,N_27163);
or U29166 (N_29166,N_25973,N_26549);
and U29167 (N_29167,N_25776,N_25801);
xor U29168 (N_29168,N_27302,N_26197);
nand U29169 (N_29169,N_26655,N_26401);
nor U29170 (N_29170,N_26525,N_27219);
and U29171 (N_29171,N_25402,N_26579);
xnor U29172 (N_29172,N_25869,N_25867);
nand U29173 (N_29173,N_25460,N_27043);
and U29174 (N_29174,N_25458,N_25479);
nor U29175 (N_29175,N_25279,N_27471);
and U29176 (N_29176,N_25210,N_27206);
nand U29177 (N_29177,N_25804,N_25034);
xnor U29178 (N_29178,N_27362,N_25019);
xor U29179 (N_29179,N_27476,N_25309);
or U29180 (N_29180,N_25445,N_26465);
or U29181 (N_29181,N_27400,N_27432);
nand U29182 (N_29182,N_26817,N_26724);
nand U29183 (N_29183,N_25233,N_25742);
xnor U29184 (N_29184,N_25589,N_26419);
nor U29185 (N_29185,N_26055,N_27141);
nor U29186 (N_29186,N_26616,N_25683);
and U29187 (N_29187,N_27198,N_26708);
and U29188 (N_29188,N_26998,N_25919);
nor U29189 (N_29189,N_26667,N_25339);
or U29190 (N_29190,N_25133,N_26381);
or U29191 (N_29191,N_26227,N_25583);
or U29192 (N_29192,N_27030,N_25690);
xor U29193 (N_29193,N_25100,N_25178);
or U29194 (N_29194,N_26694,N_26710);
and U29195 (N_29195,N_25260,N_27242);
xor U29196 (N_29196,N_25979,N_26469);
or U29197 (N_29197,N_25750,N_27236);
nand U29198 (N_29198,N_25602,N_26662);
nand U29199 (N_29199,N_25828,N_25277);
or U29200 (N_29200,N_26341,N_26676);
or U29201 (N_29201,N_27420,N_26109);
nand U29202 (N_29202,N_26450,N_25847);
xnor U29203 (N_29203,N_26208,N_25419);
and U29204 (N_29204,N_25144,N_25954);
and U29205 (N_29205,N_27348,N_25781);
or U29206 (N_29206,N_26868,N_26549);
nor U29207 (N_29207,N_26623,N_25056);
xor U29208 (N_29208,N_25988,N_27301);
nor U29209 (N_29209,N_26404,N_26021);
nand U29210 (N_29210,N_27260,N_26334);
nand U29211 (N_29211,N_26470,N_25759);
xnor U29212 (N_29212,N_27242,N_25175);
xnor U29213 (N_29213,N_25019,N_25514);
nor U29214 (N_29214,N_25918,N_27302);
and U29215 (N_29215,N_25625,N_25059);
or U29216 (N_29216,N_25158,N_25805);
nor U29217 (N_29217,N_26605,N_26478);
and U29218 (N_29218,N_27083,N_26980);
nand U29219 (N_29219,N_25160,N_25796);
xor U29220 (N_29220,N_26058,N_25739);
nor U29221 (N_29221,N_26590,N_25109);
xnor U29222 (N_29222,N_25740,N_25793);
xor U29223 (N_29223,N_25255,N_26044);
nand U29224 (N_29224,N_27152,N_25909);
or U29225 (N_29225,N_25770,N_27177);
xor U29226 (N_29226,N_27279,N_25000);
nor U29227 (N_29227,N_25028,N_26325);
or U29228 (N_29228,N_27258,N_25810);
xor U29229 (N_29229,N_25762,N_25495);
or U29230 (N_29230,N_25421,N_26317);
nor U29231 (N_29231,N_27229,N_25691);
or U29232 (N_29232,N_27316,N_27260);
nor U29233 (N_29233,N_25728,N_25317);
or U29234 (N_29234,N_26148,N_27287);
xnor U29235 (N_29235,N_26820,N_25775);
xnor U29236 (N_29236,N_25881,N_26396);
or U29237 (N_29237,N_25848,N_26932);
and U29238 (N_29238,N_25076,N_25570);
xor U29239 (N_29239,N_27210,N_25811);
nor U29240 (N_29240,N_27456,N_26525);
xnor U29241 (N_29241,N_27264,N_26165);
nor U29242 (N_29242,N_25852,N_25751);
nor U29243 (N_29243,N_27151,N_27270);
and U29244 (N_29244,N_26310,N_27444);
and U29245 (N_29245,N_25554,N_27387);
xor U29246 (N_29246,N_26363,N_25408);
or U29247 (N_29247,N_26191,N_26963);
xor U29248 (N_29248,N_27298,N_26894);
and U29249 (N_29249,N_26948,N_25002);
nand U29250 (N_29250,N_25795,N_26095);
nor U29251 (N_29251,N_25512,N_25447);
nand U29252 (N_29252,N_26183,N_26173);
nand U29253 (N_29253,N_27311,N_27475);
nand U29254 (N_29254,N_25450,N_26108);
xnor U29255 (N_29255,N_25326,N_25044);
nand U29256 (N_29256,N_25394,N_26494);
or U29257 (N_29257,N_25426,N_25638);
or U29258 (N_29258,N_26861,N_26741);
xnor U29259 (N_29259,N_25428,N_25505);
nor U29260 (N_29260,N_25816,N_25958);
and U29261 (N_29261,N_26761,N_25898);
or U29262 (N_29262,N_26438,N_25761);
nor U29263 (N_29263,N_25298,N_26690);
or U29264 (N_29264,N_26541,N_26080);
or U29265 (N_29265,N_26275,N_26713);
and U29266 (N_29266,N_26259,N_25155);
nand U29267 (N_29267,N_25437,N_26988);
and U29268 (N_29268,N_27357,N_25317);
nor U29269 (N_29269,N_25238,N_26523);
nor U29270 (N_29270,N_26839,N_26892);
nand U29271 (N_29271,N_25519,N_25434);
nor U29272 (N_29272,N_27421,N_26764);
or U29273 (N_29273,N_26669,N_26716);
nand U29274 (N_29274,N_26175,N_25109);
or U29275 (N_29275,N_27371,N_27281);
nand U29276 (N_29276,N_25839,N_26450);
and U29277 (N_29277,N_25309,N_27211);
xnor U29278 (N_29278,N_25014,N_25883);
and U29279 (N_29279,N_26381,N_25571);
nand U29280 (N_29280,N_26698,N_27237);
or U29281 (N_29281,N_25843,N_26474);
nor U29282 (N_29282,N_25963,N_27345);
and U29283 (N_29283,N_25161,N_26558);
or U29284 (N_29284,N_25496,N_27110);
nand U29285 (N_29285,N_25373,N_25500);
nor U29286 (N_29286,N_25423,N_26053);
or U29287 (N_29287,N_27143,N_27356);
and U29288 (N_29288,N_26966,N_26015);
xor U29289 (N_29289,N_25850,N_25563);
nor U29290 (N_29290,N_27450,N_25729);
or U29291 (N_29291,N_27253,N_26818);
xnor U29292 (N_29292,N_26154,N_25831);
or U29293 (N_29293,N_26653,N_25705);
and U29294 (N_29294,N_26488,N_25494);
or U29295 (N_29295,N_26596,N_26542);
xnor U29296 (N_29296,N_25220,N_27302);
nor U29297 (N_29297,N_25918,N_26197);
nor U29298 (N_29298,N_25200,N_27435);
and U29299 (N_29299,N_26034,N_25504);
nand U29300 (N_29300,N_27380,N_27429);
or U29301 (N_29301,N_25116,N_25013);
nand U29302 (N_29302,N_25403,N_25542);
nor U29303 (N_29303,N_27038,N_26236);
nand U29304 (N_29304,N_25897,N_25423);
or U29305 (N_29305,N_25292,N_26450);
and U29306 (N_29306,N_26660,N_25612);
and U29307 (N_29307,N_25214,N_25977);
xnor U29308 (N_29308,N_25562,N_27405);
or U29309 (N_29309,N_26459,N_25180);
nand U29310 (N_29310,N_26357,N_26935);
and U29311 (N_29311,N_25965,N_26628);
and U29312 (N_29312,N_26606,N_25816);
or U29313 (N_29313,N_26568,N_26194);
xor U29314 (N_29314,N_27410,N_26191);
and U29315 (N_29315,N_25376,N_27061);
or U29316 (N_29316,N_26836,N_25942);
nand U29317 (N_29317,N_25482,N_26711);
or U29318 (N_29318,N_25813,N_26658);
and U29319 (N_29319,N_26273,N_25490);
or U29320 (N_29320,N_27120,N_25603);
xor U29321 (N_29321,N_25947,N_26352);
nand U29322 (N_29322,N_27174,N_26635);
and U29323 (N_29323,N_26434,N_25586);
nand U29324 (N_29324,N_26008,N_27360);
or U29325 (N_29325,N_25168,N_25281);
and U29326 (N_29326,N_25273,N_26183);
or U29327 (N_29327,N_27020,N_25423);
xor U29328 (N_29328,N_25235,N_25803);
and U29329 (N_29329,N_25424,N_25211);
and U29330 (N_29330,N_27302,N_25423);
nand U29331 (N_29331,N_26329,N_25151);
and U29332 (N_29332,N_25533,N_25420);
xnor U29333 (N_29333,N_25996,N_25647);
and U29334 (N_29334,N_26233,N_26381);
nor U29335 (N_29335,N_26562,N_26037);
nand U29336 (N_29336,N_25139,N_27080);
xor U29337 (N_29337,N_27349,N_26264);
xor U29338 (N_29338,N_25312,N_26383);
xor U29339 (N_29339,N_26644,N_26548);
xor U29340 (N_29340,N_25318,N_25753);
xnor U29341 (N_29341,N_25586,N_26944);
or U29342 (N_29342,N_25722,N_25297);
xor U29343 (N_29343,N_25623,N_25387);
nor U29344 (N_29344,N_25771,N_25155);
xor U29345 (N_29345,N_27232,N_25276);
nor U29346 (N_29346,N_25357,N_25706);
xnor U29347 (N_29347,N_25118,N_26753);
xnor U29348 (N_29348,N_25215,N_26874);
xnor U29349 (N_29349,N_25376,N_26564);
nand U29350 (N_29350,N_25477,N_25966);
nor U29351 (N_29351,N_25461,N_26261);
nand U29352 (N_29352,N_25046,N_27397);
nor U29353 (N_29353,N_26492,N_25966);
nand U29354 (N_29354,N_26310,N_26222);
and U29355 (N_29355,N_25547,N_26273);
nor U29356 (N_29356,N_27100,N_26732);
or U29357 (N_29357,N_26931,N_26352);
or U29358 (N_29358,N_26518,N_26806);
or U29359 (N_29359,N_25245,N_25741);
nor U29360 (N_29360,N_26820,N_26387);
nor U29361 (N_29361,N_26408,N_27486);
nor U29362 (N_29362,N_27275,N_25970);
nand U29363 (N_29363,N_25997,N_25258);
nand U29364 (N_29364,N_27134,N_26933);
and U29365 (N_29365,N_25805,N_27073);
nand U29366 (N_29366,N_26420,N_26596);
nor U29367 (N_29367,N_25586,N_26021);
xnor U29368 (N_29368,N_26891,N_27048);
or U29369 (N_29369,N_25818,N_25180);
xor U29370 (N_29370,N_26590,N_26347);
and U29371 (N_29371,N_26610,N_25770);
or U29372 (N_29372,N_25412,N_25360);
xnor U29373 (N_29373,N_25996,N_25843);
nand U29374 (N_29374,N_27484,N_25765);
nor U29375 (N_29375,N_25718,N_25466);
nor U29376 (N_29376,N_25215,N_25235);
xnor U29377 (N_29377,N_26797,N_26770);
nor U29378 (N_29378,N_25734,N_25949);
or U29379 (N_29379,N_26111,N_26225);
and U29380 (N_29380,N_27117,N_26025);
nand U29381 (N_29381,N_27378,N_26459);
or U29382 (N_29382,N_26468,N_26012);
and U29383 (N_29383,N_25870,N_25421);
or U29384 (N_29384,N_25806,N_27268);
or U29385 (N_29385,N_25541,N_26089);
nor U29386 (N_29386,N_27093,N_26362);
or U29387 (N_29387,N_26611,N_26581);
nand U29388 (N_29388,N_27086,N_25542);
and U29389 (N_29389,N_25480,N_26988);
and U29390 (N_29390,N_26074,N_25702);
xor U29391 (N_29391,N_25002,N_25966);
or U29392 (N_29392,N_26489,N_26437);
and U29393 (N_29393,N_26057,N_26295);
xor U29394 (N_29394,N_26917,N_27016);
and U29395 (N_29395,N_25262,N_25319);
xor U29396 (N_29396,N_26564,N_25318);
xnor U29397 (N_29397,N_26905,N_27484);
xnor U29398 (N_29398,N_26789,N_25019);
xor U29399 (N_29399,N_27409,N_27292);
and U29400 (N_29400,N_26282,N_26751);
nand U29401 (N_29401,N_25766,N_25068);
and U29402 (N_29402,N_25662,N_26258);
and U29403 (N_29403,N_26907,N_26760);
xnor U29404 (N_29404,N_27441,N_25880);
and U29405 (N_29405,N_26266,N_25223);
or U29406 (N_29406,N_26734,N_25813);
nand U29407 (N_29407,N_25636,N_27138);
or U29408 (N_29408,N_26886,N_25548);
and U29409 (N_29409,N_27012,N_26058);
xor U29410 (N_29410,N_25978,N_26422);
and U29411 (N_29411,N_27052,N_26171);
nor U29412 (N_29412,N_25474,N_26298);
nor U29413 (N_29413,N_27479,N_25931);
or U29414 (N_29414,N_26303,N_25643);
xnor U29415 (N_29415,N_27080,N_25954);
nor U29416 (N_29416,N_26603,N_26231);
and U29417 (N_29417,N_26422,N_27323);
and U29418 (N_29418,N_25728,N_25307);
nand U29419 (N_29419,N_25924,N_25298);
nor U29420 (N_29420,N_27406,N_26018);
xnor U29421 (N_29421,N_26909,N_26840);
nor U29422 (N_29422,N_25443,N_26291);
nand U29423 (N_29423,N_26024,N_25013);
and U29424 (N_29424,N_25248,N_25236);
nand U29425 (N_29425,N_26254,N_25080);
xor U29426 (N_29426,N_26364,N_26269);
xnor U29427 (N_29427,N_27461,N_27002);
xnor U29428 (N_29428,N_26370,N_25993);
nor U29429 (N_29429,N_26633,N_25023);
or U29430 (N_29430,N_26655,N_27325);
or U29431 (N_29431,N_25925,N_25903);
nand U29432 (N_29432,N_25715,N_26266);
or U29433 (N_29433,N_26669,N_25012);
nor U29434 (N_29434,N_26285,N_25709);
nand U29435 (N_29435,N_25971,N_26643);
and U29436 (N_29436,N_26180,N_27028);
nor U29437 (N_29437,N_27066,N_25281);
xor U29438 (N_29438,N_25284,N_27481);
xor U29439 (N_29439,N_26952,N_25458);
nand U29440 (N_29440,N_26340,N_25560);
and U29441 (N_29441,N_25159,N_25434);
nand U29442 (N_29442,N_27456,N_26015);
xor U29443 (N_29443,N_27448,N_25041);
xnor U29444 (N_29444,N_27275,N_26077);
and U29445 (N_29445,N_26611,N_27437);
nand U29446 (N_29446,N_26666,N_27426);
and U29447 (N_29447,N_25828,N_26674);
nand U29448 (N_29448,N_27417,N_25629);
nor U29449 (N_29449,N_25318,N_26052);
or U29450 (N_29450,N_26077,N_26043);
and U29451 (N_29451,N_25369,N_25749);
xnor U29452 (N_29452,N_27313,N_26662);
nand U29453 (N_29453,N_25814,N_25652);
or U29454 (N_29454,N_25902,N_26652);
and U29455 (N_29455,N_25108,N_27390);
xnor U29456 (N_29456,N_26686,N_26482);
and U29457 (N_29457,N_27459,N_27150);
xor U29458 (N_29458,N_25332,N_25969);
or U29459 (N_29459,N_25888,N_25878);
nor U29460 (N_29460,N_25019,N_26507);
or U29461 (N_29461,N_25797,N_25906);
xnor U29462 (N_29462,N_26276,N_25725);
or U29463 (N_29463,N_26669,N_25986);
and U29464 (N_29464,N_26386,N_25316);
or U29465 (N_29465,N_27256,N_25324);
xor U29466 (N_29466,N_25799,N_25578);
and U29467 (N_29467,N_25099,N_26666);
xnor U29468 (N_29468,N_27420,N_25184);
and U29469 (N_29469,N_25572,N_25154);
or U29470 (N_29470,N_26986,N_26482);
nand U29471 (N_29471,N_26366,N_26036);
or U29472 (N_29472,N_26432,N_25945);
or U29473 (N_29473,N_25751,N_25666);
or U29474 (N_29474,N_25821,N_27236);
nor U29475 (N_29475,N_25977,N_26982);
nand U29476 (N_29476,N_26844,N_26930);
or U29477 (N_29477,N_27386,N_27160);
nor U29478 (N_29478,N_26000,N_25909);
xor U29479 (N_29479,N_27139,N_26210);
nor U29480 (N_29480,N_26200,N_27395);
xor U29481 (N_29481,N_26947,N_26062);
or U29482 (N_29482,N_25162,N_27408);
xor U29483 (N_29483,N_27444,N_26245);
xor U29484 (N_29484,N_25019,N_27408);
nor U29485 (N_29485,N_25559,N_26772);
nor U29486 (N_29486,N_26884,N_26931);
nand U29487 (N_29487,N_25927,N_27360);
and U29488 (N_29488,N_25299,N_26649);
or U29489 (N_29489,N_26955,N_25600);
nor U29490 (N_29490,N_25001,N_25567);
nor U29491 (N_29491,N_25775,N_25630);
or U29492 (N_29492,N_25156,N_27136);
and U29493 (N_29493,N_25795,N_25384);
nor U29494 (N_29494,N_25555,N_26735);
nor U29495 (N_29495,N_26991,N_26986);
or U29496 (N_29496,N_27223,N_26711);
nor U29497 (N_29497,N_27063,N_25959);
nor U29498 (N_29498,N_25728,N_25953);
nor U29499 (N_29499,N_25926,N_25240);
nor U29500 (N_29500,N_26119,N_26738);
nand U29501 (N_29501,N_25612,N_27109);
xnor U29502 (N_29502,N_26532,N_25684);
nand U29503 (N_29503,N_26698,N_25554);
nor U29504 (N_29504,N_27263,N_27365);
or U29505 (N_29505,N_25516,N_25622);
nand U29506 (N_29506,N_27050,N_25416);
and U29507 (N_29507,N_27226,N_25614);
or U29508 (N_29508,N_26305,N_25856);
or U29509 (N_29509,N_26534,N_25710);
nand U29510 (N_29510,N_26122,N_26225);
and U29511 (N_29511,N_27249,N_26542);
or U29512 (N_29512,N_25349,N_27419);
xor U29513 (N_29513,N_26896,N_25363);
and U29514 (N_29514,N_25496,N_25837);
nand U29515 (N_29515,N_25398,N_25071);
or U29516 (N_29516,N_26630,N_25036);
or U29517 (N_29517,N_26776,N_25836);
xor U29518 (N_29518,N_25766,N_26010);
nand U29519 (N_29519,N_26665,N_25947);
nand U29520 (N_29520,N_25499,N_25201);
or U29521 (N_29521,N_25449,N_26884);
nand U29522 (N_29522,N_27081,N_26008);
nor U29523 (N_29523,N_26264,N_26405);
and U29524 (N_29524,N_26648,N_26844);
xor U29525 (N_29525,N_26159,N_25630);
and U29526 (N_29526,N_26688,N_25500);
nand U29527 (N_29527,N_25986,N_27271);
xor U29528 (N_29528,N_26394,N_26060);
and U29529 (N_29529,N_27373,N_25894);
nor U29530 (N_29530,N_25830,N_27296);
and U29531 (N_29531,N_26152,N_25076);
nor U29532 (N_29532,N_25957,N_25653);
nand U29533 (N_29533,N_27256,N_25563);
or U29534 (N_29534,N_26103,N_25598);
nand U29535 (N_29535,N_25916,N_26301);
and U29536 (N_29536,N_26881,N_27130);
nand U29537 (N_29537,N_25214,N_27198);
nor U29538 (N_29538,N_25183,N_26785);
or U29539 (N_29539,N_26441,N_25005);
or U29540 (N_29540,N_27007,N_26425);
or U29541 (N_29541,N_25730,N_26586);
nand U29542 (N_29542,N_26575,N_26074);
or U29543 (N_29543,N_26168,N_25225);
nor U29544 (N_29544,N_26715,N_26527);
nand U29545 (N_29545,N_27385,N_27400);
nand U29546 (N_29546,N_25537,N_25612);
nand U29547 (N_29547,N_25544,N_25512);
or U29548 (N_29548,N_26184,N_26559);
and U29549 (N_29549,N_25353,N_25667);
nor U29550 (N_29550,N_26683,N_26645);
xnor U29551 (N_29551,N_26161,N_27045);
or U29552 (N_29552,N_27153,N_25276);
xor U29553 (N_29553,N_26383,N_26712);
and U29554 (N_29554,N_26603,N_25257);
and U29555 (N_29555,N_25226,N_25591);
and U29556 (N_29556,N_26897,N_25844);
nand U29557 (N_29557,N_26571,N_26841);
nor U29558 (N_29558,N_26766,N_26810);
xor U29559 (N_29559,N_26971,N_26285);
xnor U29560 (N_29560,N_27149,N_26299);
xnor U29561 (N_29561,N_27428,N_25306);
and U29562 (N_29562,N_25000,N_26958);
and U29563 (N_29563,N_25274,N_26233);
or U29564 (N_29564,N_25670,N_26228);
or U29565 (N_29565,N_26330,N_26737);
or U29566 (N_29566,N_26471,N_25429);
or U29567 (N_29567,N_25501,N_26562);
or U29568 (N_29568,N_25245,N_27380);
and U29569 (N_29569,N_26812,N_26693);
and U29570 (N_29570,N_26228,N_25398);
and U29571 (N_29571,N_26806,N_25893);
or U29572 (N_29572,N_25449,N_25188);
and U29573 (N_29573,N_26160,N_25496);
xnor U29574 (N_29574,N_26395,N_26945);
and U29575 (N_29575,N_27040,N_25332);
xnor U29576 (N_29576,N_27194,N_26188);
or U29577 (N_29577,N_25196,N_25226);
or U29578 (N_29578,N_25579,N_27328);
or U29579 (N_29579,N_25778,N_26062);
or U29580 (N_29580,N_25512,N_26965);
nor U29581 (N_29581,N_27357,N_26842);
and U29582 (N_29582,N_25388,N_26412);
nand U29583 (N_29583,N_25443,N_26813);
nor U29584 (N_29584,N_26561,N_27054);
xor U29585 (N_29585,N_27345,N_26882);
nor U29586 (N_29586,N_26074,N_26002);
nand U29587 (N_29587,N_25189,N_25487);
and U29588 (N_29588,N_25716,N_26916);
nand U29589 (N_29589,N_26700,N_26146);
or U29590 (N_29590,N_26698,N_25986);
nor U29591 (N_29591,N_26418,N_25515);
and U29592 (N_29592,N_25813,N_25391);
or U29593 (N_29593,N_26085,N_27299);
nor U29594 (N_29594,N_25409,N_25280);
nor U29595 (N_29595,N_25138,N_25200);
and U29596 (N_29596,N_25646,N_27000);
nand U29597 (N_29597,N_27068,N_25306);
xor U29598 (N_29598,N_25381,N_26535);
nor U29599 (N_29599,N_26973,N_26235);
xor U29600 (N_29600,N_27108,N_25491);
xnor U29601 (N_29601,N_25054,N_26040);
xnor U29602 (N_29602,N_26502,N_27338);
xnor U29603 (N_29603,N_26431,N_25003);
or U29604 (N_29604,N_26859,N_25986);
nand U29605 (N_29605,N_25556,N_25610);
nor U29606 (N_29606,N_25302,N_26238);
and U29607 (N_29607,N_26975,N_27226);
or U29608 (N_29608,N_25417,N_27277);
or U29609 (N_29609,N_25485,N_25488);
nor U29610 (N_29610,N_26305,N_25848);
nor U29611 (N_29611,N_25192,N_26901);
nand U29612 (N_29612,N_27469,N_26091);
xor U29613 (N_29613,N_26613,N_26989);
and U29614 (N_29614,N_26228,N_26662);
nand U29615 (N_29615,N_27115,N_25071);
nor U29616 (N_29616,N_25280,N_26745);
xnor U29617 (N_29617,N_26983,N_25375);
nand U29618 (N_29618,N_25373,N_25600);
xor U29619 (N_29619,N_26304,N_25221);
nor U29620 (N_29620,N_26807,N_26475);
and U29621 (N_29621,N_26379,N_26880);
nand U29622 (N_29622,N_26205,N_27183);
and U29623 (N_29623,N_25161,N_26892);
nor U29624 (N_29624,N_26830,N_27028);
nand U29625 (N_29625,N_25639,N_25148);
or U29626 (N_29626,N_26328,N_26417);
nand U29627 (N_29627,N_27376,N_27350);
and U29628 (N_29628,N_27139,N_26510);
or U29629 (N_29629,N_25083,N_26930);
and U29630 (N_29630,N_25075,N_27258);
nand U29631 (N_29631,N_25797,N_25398);
xnor U29632 (N_29632,N_25366,N_26198);
or U29633 (N_29633,N_25678,N_26890);
nand U29634 (N_29634,N_26289,N_26464);
or U29635 (N_29635,N_26462,N_25828);
xnor U29636 (N_29636,N_25635,N_26796);
nand U29637 (N_29637,N_26600,N_27028);
xnor U29638 (N_29638,N_26610,N_27094);
or U29639 (N_29639,N_25924,N_26396);
xnor U29640 (N_29640,N_25409,N_27029);
nor U29641 (N_29641,N_25939,N_26945);
nand U29642 (N_29642,N_26533,N_25630);
nand U29643 (N_29643,N_27223,N_25548);
nand U29644 (N_29644,N_25799,N_26453);
nand U29645 (N_29645,N_26482,N_26999);
xor U29646 (N_29646,N_26071,N_26613);
nor U29647 (N_29647,N_25821,N_26020);
or U29648 (N_29648,N_25281,N_25278);
nand U29649 (N_29649,N_25253,N_26896);
or U29650 (N_29650,N_26619,N_27132);
nor U29651 (N_29651,N_25087,N_26514);
xnor U29652 (N_29652,N_26346,N_25062);
xor U29653 (N_29653,N_27258,N_27159);
and U29654 (N_29654,N_25896,N_27159);
and U29655 (N_29655,N_27030,N_26590);
xnor U29656 (N_29656,N_26653,N_25915);
xor U29657 (N_29657,N_25899,N_27187);
nor U29658 (N_29658,N_27329,N_27404);
nor U29659 (N_29659,N_25296,N_27140);
nand U29660 (N_29660,N_25307,N_26250);
nand U29661 (N_29661,N_25397,N_25780);
xnor U29662 (N_29662,N_27335,N_26861);
nor U29663 (N_29663,N_25886,N_25833);
nor U29664 (N_29664,N_27054,N_25847);
or U29665 (N_29665,N_26493,N_26819);
or U29666 (N_29666,N_25239,N_26458);
xor U29667 (N_29667,N_25789,N_25589);
nor U29668 (N_29668,N_27295,N_26365);
nand U29669 (N_29669,N_26309,N_26085);
nand U29670 (N_29670,N_27199,N_26396);
nor U29671 (N_29671,N_25812,N_25579);
nor U29672 (N_29672,N_27400,N_26904);
xor U29673 (N_29673,N_26629,N_26776);
and U29674 (N_29674,N_25846,N_27005);
or U29675 (N_29675,N_25909,N_26832);
nand U29676 (N_29676,N_26498,N_25561);
nor U29677 (N_29677,N_27374,N_25501);
xnor U29678 (N_29678,N_27214,N_25483);
or U29679 (N_29679,N_27030,N_25022);
and U29680 (N_29680,N_26258,N_27208);
nor U29681 (N_29681,N_27271,N_27315);
nand U29682 (N_29682,N_26743,N_25259);
or U29683 (N_29683,N_27382,N_27021);
or U29684 (N_29684,N_26970,N_25843);
or U29685 (N_29685,N_26205,N_26235);
and U29686 (N_29686,N_25719,N_26180);
nor U29687 (N_29687,N_26882,N_27021);
and U29688 (N_29688,N_25287,N_26093);
or U29689 (N_29689,N_27203,N_25255);
xnor U29690 (N_29690,N_25909,N_25022);
and U29691 (N_29691,N_27291,N_25179);
or U29692 (N_29692,N_25787,N_25132);
and U29693 (N_29693,N_26646,N_26821);
nor U29694 (N_29694,N_25478,N_26593);
and U29695 (N_29695,N_25705,N_27411);
nand U29696 (N_29696,N_25785,N_26646);
or U29697 (N_29697,N_27147,N_26473);
nor U29698 (N_29698,N_26908,N_25412);
nand U29699 (N_29699,N_26522,N_25990);
nand U29700 (N_29700,N_26066,N_25329);
xnor U29701 (N_29701,N_26699,N_26777);
nor U29702 (N_29702,N_26836,N_27495);
xor U29703 (N_29703,N_25713,N_26011);
or U29704 (N_29704,N_26089,N_25548);
nand U29705 (N_29705,N_26344,N_25421);
nor U29706 (N_29706,N_26555,N_26107);
and U29707 (N_29707,N_26846,N_25675);
xor U29708 (N_29708,N_25009,N_25649);
and U29709 (N_29709,N_26708,N_26384);
and U29710 (N_29710,N_27122,N_25202);
xor U29711 (N_29711,N_26985,N_26896);
xnor U29712 (N_29712,N_26670,N_26724);
and U29713 (N_29713,N_25582,N_26386);
nand U29714 (N_29714,N_26949,N_25116);
nand U29715 (N_29715,N_27127,N_27036);
nor U29716 (N_29716,N_25542,N_25084);
nand U29717 (N_29717,N_26541,N_26737);
nor U29718 (N_29718,N_27191,N_26802);
nor U29719 (N_29719,N_26097,N_25653);
nor U29720 (N_29720,N_27376,N_25410);
nor U29721 (N_29721,N_25805,N_25248);
nand U29722 (N_29722,N_27368,N_25930);
nor U29723 (N_29723,N_25778,N_25195);
or U29724 (N_29724,N_27000,N_26753);
xnor U29725 (N_29725,N_25279,N_27285);
nor U29726 (N_29726,N_27250,N_25266);
nor U29727 (N_29727,N_25485,N_27315);
xnor U29728 (N_29728,N_26884,N_25333);
and U29729 (N_29729,N_26705,N_25035);
and U29730 (N_29730,N_26844,N_27469);
xnor U29731 (N_29731,N_27016,N_25082);
or U29732 (N_29732,N_27378,N_27223);
nor U29733 (N_29733,N_27475,N_26183);
nand U29734 (N_29734,N_25112,N_25827);
nor U29735 (N_29735,N_26361,N_26632);
xor U29736 (N_29736,N_25697,N_27115);
xor U29737 (N_29737,N_26962,N_26840);
xnor U29738 (N_29738,N_27312,N_26697);
xnor U29739 (N_29739,N_27343,N_25861);
nand U29740 (N_29740,N_25645,N_25989);
nor U29741 (N_29741,N_25571,N_27090);
nand U29742 (N_29742,N_26473,N_26618);
and U29743 (N_29743,N_27076,N_26718);
xnor U29744 (N_29744,N_25272,N_27427);
or U29745 (N_29745,N_25128,N_27375);
nor U29746 (N_29746,N_25012,N_27014);
or U29747 (N_29747,N_25417,N_26734);
nor U29748 (N_29748,N_27425,N_26974);
or U29749 (N_29749,N_27228,N_27455);
nor U29750 (N_29750,N_25944,N_25333);
nand U29751 (N_29751,N_25484,N_26223);
nor U29752 (N_29752,N_25983,N_27231);
nor U29753 (N_29753,N_25556,N_25140);
nand U29754 (N_29754,N_26967,N_26835);
and U29755 (N_29755,N_26884,N_27291);
nor U29756 (N_29756,N_25476,N_26654);
nor U29757 (N_29757,N_25212,N_26972);
or U29758 (N_29758,N_25954,N_25357);
nor U29759 (N_29759,N_25964,N_26779);
or U29760 (N_29760,N_25544,N_26753);
nand U29761 (N_29761,N_25672,N_26973);
and U29762 (N_29762,N_27327,N_25270);
xnor U29763 (N_29763,N_25843,N_27339);
xnor U29764 (N_29764,N_25439,N_25211);
or U29765 (N_29765,N_27350,N_26246);
nor U29766 (N_29766,N_27232,N_25452);
xor U29767 (N_29767,N_26834,N_26146);
or U29768 (N_29768,N_25869,N_26291);
xor U29769 (N_29769,N_25508,N_25875);
nor U29770 (N_29770,N_27114,N_25502);
or U29771 (N_29771,N_25310,N_25969);
nor U29772 (N_29772,N_26133,N_25503);
xor U29773 (N_29773,N_26675,N_25634);
and U29774 (N_29774,N_26177,N_27021);
and U29775 (N_29775,N_26065,N_26462);
and U29776 (N_29776,N_25097,N_25483);
and U29777 (N_29777,N_25681,N_25542);
and U29778 (N_29778,N_26269,N_25587);
xor U29779 (N_29779,N_26602,N_26168);
nor U29780 (N_29780,N_26081,N_27068);
xor U29781 (N_29781,N_26019,N_25354);
nor U29782 (N_29782,N_26277,N_25181);
nand U29783 (N_29783,N_26923,N_27375);
nand U29784 (N_29784,N_25020,N_25659);
and U29785 (N_29785,N_25673,N_26817);
nor U29786 (N_29786,N_26821,N_26279);
or U29787 (N_29787,N_26347,N_26217);
nor U29788 (N_29788,N_27330,N_26628);
and U29789 (N_29789,N_26655,N_26635);
or U29790 (N_29790,N_26115,N_25372);
xor U29791 (N_29791,N_26340,N_25837);
and U29792 (N_29792,N_25618,N_26926);
xnor U29793 (N_29793,N_27160,N_25525);
and U29794 (N_29794,N_25960,N_25501);
xnor U29795 (N_29795,N_25950,N_25547);
and U29796 (N_29796,N_27195,N_25023);
xnor U29797 (N_29797,N_27163,N_27085);
or U29798 (N_29798,N_26714,N_26009);
or U29799 (N_29799,N_27336,N_25800);
xnor U29800 (N_29800,N_25128,N_26046);
nand U29801 (N_29801,N_25208,N_25986);
or U29802 (N_29802,N_25480,N_25408);
nand U29803 (N_29803,N_25811,N_25507);
nand U29804 (N_29804,N_26402,N_26766);
nand U29805 (N_29805,N_25020,N_27087);
or U29806 (N_29806,N_25548,N_25413);
or U29807 (N_29807,N_25232,N_25216);
nor U29808 (N_29808,N_25062,N_25154);
and U29809 (N_29809,N_25800,N_27328);
nor U29810 (N_29810,N_25479,N_25420);
and U29811 (N_29811,N_25389,N_25390);
nand U29812 (N_29812,N_25031,N_27447);
nor U29813 (N_29813,N_27147,N_25897);
xor U29814 (N_29814,N_26658,N_26817);
and U29815 (N_29815,N_25872,N_26987);
or U29816 (N_29816,N_26716,N_26667);
nor U29817 (N_29817,N_26819,N_27121);
xnor U29818 (N_29818,N_25555,N_26813);
or U29819 (N_29819,N_25408,N_26456);
and U29820 (N_29820,N_26484,N_25598);
or U29821 (N_29821,N_26781,N_26691);
nand U29822 (N_29822,N_26200,N_25206);
nor U29823 (N_29823,N_27188,N_25081);
and U29824 (N_29824,N_25450,N_27280);
xor U29825 (N_29825,N_26477,N_25922);
nor U29826 (N_29826,N_26480,N_27116);
xnor U29827 (N_29827,N_26738,N_25623);
xnor U29828 (N_29828,N_25078,N_26586);
nor U29829 (N_29829,N_25728,N_25383);
or U29830 (N_29830,N_26919,N_26450);
nor U29831 (N_29831,N_27351,N_26980);
and U29832 (N_29832,N_25345,N_26927);
and U29833 (N_29833,N_26675,N_26705);
nor U29834 (N_29834,N_25887,N_25559);
nand U29835 (N_29835,N_25082,N_26979);
and U29836 (N_29836,N_26819,N_26704);
xnor U29837 (N_29837,N_25800,N_25795);
nor U29838 (N_29838,N_26531,N_26217);
and U29839 (N_29839,N_26449,N_26457);
or U29840 (N_29840,N_25057,N_25109);
and U29841 (N_29841,N_26076,N_25493);
nor U29842 (N_29842,N_25168,N_25705);
and U29843 (N_29843,N_27376,N_26399);
nor U29844 (N_29844,N_26612,N_25633);
xor U29845 (N_29845,N_26567,N_25202);
nand U29846 (N_29846,N_26033,N_25180);
or U29847 (N_29847,N_25596,N_26912);
nand U29848 (N_29848,N_25007,N_27287);
or U29849 (N_29849,N_25258,N_25013);
and U29850 (N_29850,N_27414,N_26743);
xnor U29851 (N_29851,N_26891,N_25598);
nor U29852 (N_29852,N_26824,N_26847);
or U29853 (N_29853,N_27357,N_26415);
and U29854 (N_29854,N_25134,N_27080);
or U29855 (N_29855,N_25519,N_26504);
or U29856 (N_29856,N_25272,N_26162);
or U29857 (N_29857,N_27247,N_27447);
xor U29858 (N_29858,N_27134,N_25428);
nand U29859 (N_29859,N_25922,N_27378);
nand U29860 (N_29860,N_26710,N_25607);
nor U29861 (N_29861,N_26527,N_26470);
nor U29862 (N_29862,N_26193,N_26710);
xnor U29863 (N_29863,N_25680,N_27371);
or U29864 (N_29864,N_25795,N_25269);
nor U29865 (N_29865,N_27459,N_26520);
and U29866 (N_29866,N_25124,N_25120);
nand U29867 (N_29867,N_25525,N_25860);
and U29868 (N_29868,N_25828,N_26777);
nor U29869 (N_29869,N_25848,N_27430);
nand U29870 (N_29870,N_25671,N_25901);
and U29871 (N_29871,N_25058,N_25717);
and U29872 (N_29872,N_26377,N_25005);
nand U29873 (N_29873,N_27105,N_25952);
nor U29874 (N_29874,N_27139,N_25169);
or U29875 (N_29875,N_26671,N_27242);
nand U29876 (N_29876,N_26526,N_25377);
xor U29877 (N_29877,N_26746,N_26757);
nor U29878 (N_29878,N_26561,N_26256);
and U29879 (N_29879,N_25215,N_25069);
nor U29880 (N_29880,N_26220,N_25906);
nor U29881 (N_29881,N_26311,N_27355);
xor U29882 (N_29882,N_26393,N_25852);
and U29883 (N_29883,N_26296,N_25626);
or U29884 (N_29884,N_27402,N_25921);
or U29885 (N_29885,N_27448,N_27137);
nor U29886 (N_29886,N_25058,N_26201);
nand U29887 (N_29887,N_25949,N_26053);
nor U29888 (N_29888,N_27189,N_25579);
xor U29889 (N_29889,N_25051,N_26307);
or U29890 (N_29890,N_25731,N_26263);
xor U29891 (N_29891,N_25312,N_26375);
nor U29892 (N_29892,N_25531,N_26263);
or U29893 (N_29893,N_25454,N_26084);
nand U29894 (N_29894,N_25011,N_26370);
nor U29895 (N_29895,N_25090,N_25251);
xor U29896 (N_29896,N_26118,N_25231);
xnor U29897 (N_29897,N_26793,N_27267);
nor U29898 (N_29898,N_27321,N_25913);
and U29899 (N_29899,N_25380,N_26950);
nor U29900 (N_29900,N_26135,N_25343);
nand U29901 (N_29901,N_25384,N_26631);
xnor U29902 (N_29902,N_27217,N_25043);
nor U29903 (N_29903,N_25300,N_25192);
or U29904 (N_29904,N_26495,N_25128);
xor U29905 (N_29905,N_25195,N_25445);
xor U29906 (N_29906,N_27255,N_25995);
nor U29907 (N_29907,N_26959,N_25153);
nand U29908 (N_29908,N_25966,N_27115);
xnor U29909 (N_29909,N_26801,N_26066);
xnor U29910 (N_29910,N_25589,N_25948);
nor U29911 (N_29911,N_25742,N_26601);
xnor U29912 (N_29912,N_25232,N_27200);
nand U29913 (N_29913,N_25259,N_26684);
xnor U29914 (N_29914,N_26709,N_26522);
xnor U29915 (N_29915,N_27330,N_25913);
xor U29916 (N_29916,N_25174,N_25102);
or U29917 (N_29917,N_26764,N_26311);
and U29918 (N_29918,N_25790,N_25022);
or U29919 (N_29919,N_27130,N_26703);
nand U29920 (N_29920,N_25234,N_27420);
or U29921 (N_29921,N_27484,N_26477);
xor U29922 (N_29922,N_26136,N_25517);
xnor U29923 (N_29923,N_26146,N_26049);
and U29924 (N_29924,N_26008,N_25550);
or U29925 (N_29925,N_26084,N_26342);
nor U29926 (N_29926,N_25938,N_25183);
and U29927 (N_29927,N_25885,N_25271);
nor U29928 (N_29928,N_27477,N_25494);
and U29929 (N_29929,N_26769,N_27133);
xnor U29930 (N_29930,N_25553,N_27236);
nor U29931 (N_29931,N_26167,N_25264);
or U29932 (N_29932,N_26110,N_25788);
xor U29933 (N_29933,N_25435,N_26781);
xnor U29934 (N_29934,N_25966,N_27015);
xnor U29935 (N_29935,N_26841,N_26717);
or U29936 (N_29936,N_26048,N_25609);
nand U29937 (N_29937,N_25101,N_27489);
or U29938 (N_29938,N_26718,N_27443);
nor U29939 (N_29939,N_26634,N_25100);
xnor U29940 (N_29940,N_27338,N_26697);
and U29941 (N_29941,N_25898,N_26929);
nand U29942 (N_29942,N_25881,N_25058);
and U29943 (N_29943,N_25845,N_25817);
xor U29944 (N_29944,N_25348,N_26016);
xor U29945 (N_29945,N_26867,N_25017);
or U29946 (N_29946,N_26418,N_26415);
and U29947 (N_29947,N_26463,N_26433);
and U29948 (N_29948,N_26678,N_27410);
nand U29949 (N_29949,N_25404,N_26398);
nor U29950 (N_29950,N_25344,N_25011);
nand U29951 (N_29951,N_26072,N_27322);
and U29952 (N_29952,N_27142,N_25177);
xnor U29953 (N_29953,N_25247,N_25073);
or U29954 (N_29954,N_26158,N_25302);
or U29955 (N_29955,N_26846,N_26206);
nand U29956 (N_29956,N_25456,N_26088);
and U29957 (N_29957,N_25347,N_26108);
xnor U29958 (N_29958,N_26120,N_25807);
xnor U29959 (N_29959,N_26332,N_27221);
or U29960 (N_29960,N_27498,N_26079);
xor U29961 (N_29961,N_26477,N_25681);
and U29962 (N_29962,N_25260,N_27363);
xor U29963 (N_29963,N_25621,N_25053);
nor U29964 (N_29964,N_27464,N_25336);
nand U29965 (N_29965,N_26651,N_26102);
or U29966 (N_29966,N_27039,N_25216);
and U29967 (N_29967,N_27163,N_25004);
nand U29968 (N_29968,N_27025,N_25313);
or U29969 (N_29969,N_26733,N_26115);
nand U29970 (N_29970,N_25504,N_27359);
and U29971 (N_29971,N_26964,N_25392);
nor U29972 (N_29972,N_26129,N_25435);
nor U29973 (N_29973,N_26251,N_26662);
xnor U29974 (N_29974,N_27456,N_26825);
nand U29975 (N_29975,N_25174,N_26545);
nor U29976 (N_29976,N_26676,N_25908);
nor U29977 (N_29977,N_25861,N_26181);
nor U29978 (N_29978,N_27273,N_26179);
nor U29979 (N_29979,N_25072,N_25138);
nand U29980 (N_29980,N_25117,N_25932);
nand U29981 (N_29981,N_27474,N_26495);
or U29982 (N_29982,N_25912,N_26296);
and U29983 (N_29983,N_27233,N_25780);
or U29984 (N_29984,N_25175,N_26774);
or U29985 (N_29985,N_26903,N_25778);
nor U29986 (N_29986,N_25664,N_26742);
and U29987 (N_29987,N_26939,N_27246);
xor U29988 (N_29988,N_25745,N_27306);
and U29989 (N_29989,N_25825,N_26818);
and U29990 (N_29990,N_27058,N_26917);
or U29991 (N_29991,N_26757,N_26875);
or U29992 (N_29992,N_26925,N_26941);
nand U29993 (N_29993,N_26151,N_27252);
nor U29994 (N_29994,N_26288,N_27202);
or U29995 (N_29995,N_27015,N_26081);
or U29996 (N_29996,N_27177,N_26513);
nor U29997 (N_29997,N_27170,N_26673);
xnor U29998 (N_29998,N_25328,N_26783);
nand U29999 (N_29999,N_27035,N_26291);
and U30000 (N_30000,N_28205,N_29648);
or U30001 (N_30001,N_28127,N_28091);
nand U30002 (N_30002,N_28490,N_29180);
xor U30003 (N_30003,N_29152,N_29317);
xnor U30004 (N_30004,N_28526,N_28022);
xnor U30005 (N_30005,N_28906,N_29594);
xor U30006 (N_30006,N_29685,N_28465);
nor U30007 (N_30007,N_29121,N_27520);
nor U30008 (N_30008,N_29170,N_27733);
nand U30009 (N_30009,N_27833,N_29944);
xor U30010 (N_30010,N_27646,N_28655);
and U30011 (N_30011,N_29559,N_28606);
nor U30012 (N_30012,N_29676,N_28397);
nor U30013 (N_30013,N_28569,N_28550);
or U30014 (N_30014,N_29848,N_29887);
or U30015 (N_30015,N_27991,N_29083);
nand U30016 (N_30016,N_28133,N_29591);
and U30017 (N_30017,N_29181,N_29896);
or U30018 (N_30018,N_29245,N_28568);
and U30019 (N_30019,N_29773,N_29712);
and U30020 (N_30020,N_28846,N_29455);
xnor U30021 (N_30021,N_29932,N_27870);
xor U30022 (N_30022,N_27570,N_27948);
nor U30023 (N_30023,N_27543,N_29775);
nand U30024 (N_30024,N_29207,N_28839);
nor U30025 (N_30025,N_28722,N_29383);
nor U30026 (N_30026,N_29628,N_28631);
xnor U30027 (N_30027,N_28105,N_28380);
and U30028 (N_30028,N_29939,N_29184);
xor U30029 (N_30029,N_27697,N_28688);
or U30030 (N_30030,N_28888,N_28609);
xnor U30031 (N_30031,N_28618,N_27686);
nor U30032 (N_30032,N_27512,N_27625);
nor U30033 (N_30033,N_29321,N_28795);
xnor U30034 (N_30034,N_28059,N_27746);
and U30035 (N_30035,N_29988,N_28416);
or U30036 (N_30036,N_28774,N_28851);
or U30037 (N_30037,N_28295,N_28373);
nand U30038 (N_30038,N_29414,N_27700);
or U30039 (N_30039,N_28979,N_28641);
and U30040 (N_30040,N_28927,N_28701);
nor U30041 (N_30041,N_28312,N_29835);
nor U30042 (N_30042,N_28625,N_27590);
nor U30043 (N_30043,N_28650,N_29711);
or U30044 (N_30044,N_29030,N_28990);
nor U30045 (N_30045,N_29094,N_29829);
xnor U30046 (N_30046,N_28462,N_29570);
nand U30047 (N_30047,N_29440,N_28532);
nor U30048 (N_30048,N_28323,N_29022);
and U30049 (N_30049,N_27943,N_28995);
nand U30050 (N_30050,N_29123,N_29320);
nor U30051 (N_30051,N_27663,N_27676);
or U30052 (N_30052,N_28772,N_29436);
xor U30053 (N_30053,N_28900,N_29062);
or U30054 (N_30054,N_29113,N_29484);
nor U30055 (N_30055,N_29836,N_28659);
xor U30056 (N_30056,N_29762,N_29754);
or U30057 (N_30057,N_27995,N_28125);
nand U30058 (N_30058,N_29086,N_29212);
nor U30059 (N_30059,N_29681,N_27982);
and U30060 (N_30060,N_27783,N_29778);
xnor U30061 (N_30061,N_29707,N_29980);
xnor U30062 (N_30062,N_28752,N_27990);
and U30063 (N_30063,N_27566,N_28513);
nor U30064 (N_30064,N_27758,N_28949);
nor U30065 (N_30065,N_28369,N_29911);
nand U30066 (N_30066,N_27537,N_29553);
or U30067 (N_30067,N_29817,N_27550);
xor U30068 (N_30068,N_27913,N_28595);
xnor U30069 (N_30069,N_27722,N_28744);
or U30070 (N_30070,N_29112,N_28703);
nor U30071 (N_30071,N_28959,N_28824);
xor U30072 (N_30072,N_27750,N_27919);
nor U30073 (N_30073,N_28756,N_28845);
nor U30074 (N_30074,N_29515,N_28931);
xnor U30075 (N_30075,N_29563,N_27630);
and U30076 (N_30076,N_28668,N_28518);
or U30077 (N_30077,N_27953,N_28149);
nor U30078 (N_30078,N_27893,N_29169);
nor U30079 (N_30079,N_28068,N_27992);
and U30080 (N_30080,N_29106,N_27578);
nand U30081 (N_30081,N_28685,N_28634);
or U30082 (N_30082,N_28502,N_27954);
nand U30083 (N_30083,N_28539,N_28183);
nor U30084 (N_30084,N_29091,N_29095);
nand U30085 (N_30085,N_28515,N_29937);
and U30086 (N_30086,N_27639,N_29781);
and U30087 (N_30087,N_29313,N_27659);
or U30088 (N_30088,N_27669,N_29950);
and U30089 (N_30089,N_29286,N_29085);
and U30090 (N_30090,N_29623,N_29649);
xor U30091 (N_30091,N_28600,N_27863);
nand U30092 (N_30092,N_28519,N_28691);
nand U30093 (N_30093,N_27635,N_29331);
and U30094 (N_30094,N_29878,N_29441);
and U30095 (N_30095,N_28135,N_28801);
xnor U30096 (N_30096,N_29188,N_28467);
and U30097 (N_30097,N_28507,N_27989);
nand U30098 (N_30098,N_28277,N_28197);
nand U30099 (N_30099,N_29010,N_28039);
nor U30100 (N_30100,N_28976,N_28769);
nor U30101 (N_30101,N_28543,N_29466);
and U30102 (N_30102,N_28740,N_29396);
nor U30103 (N_30103,N_29630,N_29415);
and U30104 (N_30104,N_29801,N_27579);
or U30105 (N_30105,N_27629,N_28709);
and U30106 (N_30106,N_27602,N_29105);
nand U30107 (N_30107,N_28436,N_29742);
xor U30108 (N_30108,N_29907,N_29229);
xor U30109 (N_30109,N_29869,N_28363);
nand U30110 (N_30110,N_29490,N_28758);
or U30111 (N_30111,N_29584,N_29716);
or U30112 (N_30112,N_28870,N_29266);
xor U30113 (N_30113,N_29476,N_29823);
nand U30114 (N_30114,N_28713,N_29862);
xor U30115 (N_30115,N_27553,N_28842);
xnor U30116 (N_30116,N_29462,N_29028);
nand U30117 (N_30117,N_29997,N_29066);
or U30118 (N_30118,N_29251,N_28360);
nand U30119 (N_30119,N_28573,N_28372);
and U30120 (N_30120,N_29400,N_28861);
nor U30121 (N_30121,N_29351,N_27946);
and U30122 (N_30122,N_29325,N_28386);
xnor U30123 (N_30123,N_29209,N_27988);
nand U30124 (N_30124,N_29362,N_28643);
and U30125 (N_30125,N_28476,N_28917);
and U30126 (N_30126,N_29644,N_28348);
nor U30127 (N_30127,N_28055,N_28245);
and U30128 (N_30128,N_29177,N_27776);
nand U30129 (N_30129,N_27816,N_28563);
or U30130 (N_30130,N_27771,N_28435);
nand U30131 (N_30131,N_27614,N_27793);
or U30132 (N_30132,N_27586,N_28002);
and U30133 (N_30133,N_29332,N_28460);
nand U30134 (N_30134,N_29468,N_29909);
nand U30135 (N_30135,N_29612,N_29750);
xnor U30136 (N_30136,N_28376,N_27956);
nand U30137 (N_30137,N_29731,N_29079);
or U30138 (N_30138,N_27661,N_28154);
nor U30139 (N_30139,N_28445,N_29984);
or U30140 (N_30140,N_27707,N_27647);
nor U30141 (N_30141,N_28297,N_28594);
and U30142 (N_30142,N_28893,N_28096);
or U30143 (N_30143,N_29689,N_27949);
nand U30144 (N_30144,N_27641,N_29956);
or U30145 (N_30145,N_29934,N_28863);
or U30146 (N_30146,N_28905,N_29507);
xnor U30147 (N_30147,N_28212,N_28967);
xnor U30148 (N_30148,N_29784,N_29398);
nand U30149 (N_30149,N_29561,N_29339);
xor U30150 (N_30150,N_28768,N_28102);
xor U30151 (N_30151,N_28880,N_28305);
nand U30152 (N_30152,N_29892,N_29970);
or U30153 (N_30153,N_28424,N_29337);
or U30154 (N_30154,N_29926,N_28596);
and U30155 (N_30155,N_29061,N_27662);
and U30156 (N_30156,N_28895,N_29993);
nor U30157 (N_30157,N_29874,N_29602);
xnor U30158 (N_30158,N_28255,N_28199);
or U30159 (N_30159,N_29885,N_28850);
nand U30160 (N_30160,N_28017,N_29705);
or U30161 (N_30161,N_28874,N_29960);
and U30162 (N_30162,N_28510,N_29994);
and U30163 (N_30163,N_28062,N_29995);
nand U30164 (N_30164,N_29147,N_29135);
nor U30165 (N_30165,N_29356,N_29726);
or U30166 (N_30166,N_27552,N_28494);
nor U30167 (N_30167,N_27908,N_29016);
and U30168 (N_30168,N_28737,N_29033);
and U30169 (N_30169,N_29524,N_28444);
xnor U30170 (N_30170,N_28064,N_28559);
and U30171 (N_30171,N_28124,N_28937);
nor U30172 (N_30172,N_28731,N_27778);
nand U30173 (N_30173,N_28030,N_27889);
nand U30174 (N_30174,N_28815,N_28457);
xor U30175 (N_30175,N_29388,N_27885);
nand U30176 (N_30176,N_28894,N_27828);
nor U30177 (N_30177,N_29223,N_29650);
xnor U30178 (N_30178,N_28946,N_29381);
or U30179 (N_30179,N_28987,N_28213);
xor U30180 (N_30180,N_28763,N_28304);
nand U30181 (N_30181,N_27767,N_28018);
nor U30182 (N_30182,N_28583,N_28551);
nor U30183 (N_30183,N_29420,N_29914);
nor U30184 (N_30184,N_29306,N_28919);
nor U30185 (N_30185,N_28443,N_27762);
or U30186 (N_30186,N_27900,N_29148);
or U30187 (N_30187,N_29897,N_29355);
or U30188 (N_30188,N_28089,N_28056);
xnor U30189 (N_30189,N_29497,N_28391);
nand U30190 (N_30190,N_29378,N_27924);
nor U30191 (N_30191,N_28252,N_29270);
xnor U30192 (N_30192,N_27691,N_28697);
nand U30193 (N_30193,N_28735,N_29670);
xnor U30194 (N_30194,N_29483,N_29881);
nor U30195 (N_30195,N_28349,N_29904);
xnor U30196 (N_30196,N_29192,N_29958);
and U30197 (N_30197,N_28470,N_28387);
nor U30198 (N_30198,N_27959,N_28725);
or U30199 (N_30199,N_29189,N_28031);
xnor U30200 (N_30200,N_29875,N_29452);
nand U30201 (N_30201,N_28378,N_29770);
nor U30202 (N_30202,N_29432,N_27677);
nor U30203 (N_30203,N_29617,N_29654);
nand U30204 (N_30204,N_27987,N_28854);
xnor U30205 (N_30205,N_27564,N_29735);
nand U30206 (N_30206,N_29384,N_28202);
xor U30207 (N_30207,N_28791,N_29424);
xnor U30208 (N_30208,N_29791,N_28804);
nand U30209 (N_30209,N_28274,N_28317);
nand U30210 (N_30210,N_27575,N_27742);
and U30211 (N_30211,N_29009,N_28482);
and U30212 (N_30212,N_28481,N_28066);
nand U30213 (N_30213,N_28817,N_29849);
and U30214 (N_30214,N_27905,N_29866);
xor U30215 (N_30215,N_27935,N_29074);
nand U30216 (N_30216,N_27560,N_28294);
nand U30217 (N_30217,N_29990,N_28965);
and U30218 (N_30218,N_28747,N_27612);
nand U30219 (N_30219,N_27916,N_28548);
or U30220 (N_30220,N_29333,N_29783);
and U30221 (N_30221,N_29653,N_27626);
nor U30222 (N_30222,N_28652,N_27645);
xor U30223 (N_30223,N_27842,N_29191);
nand U30224 (N_30224,N_29289,N_28517);
nand U30225 (N_30225,N_27653,N_29380);
nor U30226 (N_30226,N_28765,N_28131);
xnor U30227 (N_30227,N_28982,N_28330);
or U30228 (N_30228,N_29480,N_28157);
xnor U30229 (N_30229,N_29419,N_29643);
or U30230 (N_30230,N_27734,N_28816);
nand U30231 (N_30231,N_29311,N_28279);
or U30232 (N_30232,N_27985,N_28434);
nand U30233 (N_30233,N_29239,N_28867);
nor U30234 (N_30234,N_29763,N_29719);
xor U30235 (N_30235,N_27814,N_28624);
and U30236 (N_30236,N_29813,N_27631);
nor U30237 (N_30237,N_29099,N_27821);
nand U30238 (N_30238,N_29305,N_27844);
nand U30239 (N_30239,N_29855,N_29733);
or U30240 (N_30240,N_29989,N_29903);
nand U30241 (N_30241,N_27832,N_28429);
nand U30242 (N_30242,N_29609,N_28052);
nor U30243 (N_30243,N_29743,N_27593);
and U30244 (N_30244,N_29277,N_28075);
xor U30245 (N_30245,N_29512,N_27955);
nor U30246 (N_30246,N_28628,N_28243);
and U30247 (N_30247,N_28333,N_27873);
xnor U30248 (N_30248,N_29403,N_27972);
nand U30249 (N_30249,N_29021,N_28239);
nor U30250 (N_30250,N_29555,N_29366);
nor U30251 (N_30251,N_27940,N_27654);
or U30252 (N_30252,N_28500,N_27779);
or U30253 (N_30253,N_28399,N_29749);
nand U30254 (N_30254,N_27915,N_29746);
xor U30255 (N_30255,N_28367,N_27968);
nor U30256 (N_30256,N_27848,N_27652);
xnor U30257 (N_30257,N_28637,N_27978);
and U30258 (N_30258,N_29071,N_27636);
nor U30259 (N_30259,N_29371,N_28407);
nor U30260 (N_30260,N_27791,N_28474);
or U30261 (N_30261,N_27557,N_28217);
and U30262 (N_30262,N_29842,N_28253);
nor U30263 (N_30263,N_29411,N_29870);
nand U30264 (N_30264,N_29470,N_28222);
xor U30265 (N_30265,N_29531,N_27650);
nand U30266 (N_30266,N_28076,N_28060);
or U30267 (N_30267,N_28950,N_29395);
nand U30268 (N_30268,N_27737,N_28834);
nor U30269 (N_30269,N_29494,N_28947);
nor U30270 (N_30270,N_29126,N_28547);
nor U30271 (N_30271,N_29274,N_27899);
or U30272 (N_30272,N_27501,N_28148);
and U30273 (N_30273,N_29730,N_29882);
nand U30274 (N_30274,N_28475,N_27613);
nor U30275 (N_30275,N_29652,N_28352);
nor U30276 (N_30276,N_27966,N_27581);
nand U30277 (N_30277,N_29109,N_28869);
nand U30278 (N_30278,N_29698,N_29634);
nand U30279 (N_30279,N_29727,N_29089);
or U30280 (N_30280,N_28622,N_29341);
nor U30281 (N_30281,N_29430,N_28356);
and U30282 (N_30282,N_29361,N_28669);
and U30283 (N_30283,N_27514,N_28238);
and U30284 (N_30284,N_28891,N_28695);
nand U30285 (N_30285,N_28777,N_28359);
nand U30286 (N_30286,N_28726,N_27684);
or U30287 (N_30287,N_28383,N_28026);
nand U30288 (N_30288,N_28412,N_28484);
nor U30289 (N_30289,N_28389,N_27807);
nor U30290 (N_30290,N_28263,N_29544);
xnor U30291 (N_30291,N_29768,N_27588);
nand U30292 (N_30292,N_29607,N_28261);
nand U30293 (N_30293,N_28049,N_27694);
xnor U30294 (N_30294,N_28000,N_29164);
nand U30295 (N_30295,N_29661,N_28406);
nand U30296 (N_30296,N_29292,N_27508);
or U30297 (N_30297,N_29151,N_29521);
nor U30298 (N_30298,N_28511,N_28322);
and U30299 (N_30299,N_28454,N_27752);
nor U30300 (N_30300,N_29790,N_29160);
xnor U30301 (N_30301,N_28366,N_28401);
nand U30302 (N_30302,N_27739,N_29758);
xor U30303 (N_30303,N_29613,N_29172);
and U30304 (N_30304,N_28907,N_29263);
nor U30305 (N_30305,N_28073,N_28408);
or U30306 (N_30306,N_29895,N_29502);
nand U30307 (N_30307,N_28087,N_28311);
or U30308 (N_30308,N_28301,N_29008);
or U30309 (N_30309,N_29693,N_27721);
nand U30310 (N_30310,N_28398,N_28866);
nor U30311 (N_30311,N_28598,N_28796);
xnor U30312 (N_30312,N_28123,N_29663);
nor U30313 (N_30313,N_28307,N_29679);
xnor U30314 (N_30314,N_29050,N_29611);
and U30315 (N_30315,N_28902,N_29443);
nor U30316 (N_30316,N_27788,N_29640);
nand U30317 (N_30317,N_28471,N_29966);
nor U30318 (N_30318,N_29873,N_28119);
xnor U30319 (N_30319,N_28847,N_29872);
xnor U30320 (N_30320,N_29214,N_28298);
nand U30321 (N_30321,N_28542,N_29969);
or U30322 (N_30322,N_27751,N_28313);
nand U30323 (N_30323,N_29827,N_28745);
xor U30324 (N_30324,N_29401,N_28878);
and U30325 (N_30325,N_28844,N_29821);
and U30326 (N_30326,N_28792,N_28572);
xnor U30327 (N_30327,N_29883,N_28897);
or U30328 (N_30328,N_28325,N_29668);
and U30329 (N_30329,N_28964,N_28343);
xor U30330 (N_30330,N_29275,N_29672);
nor U30331 (N_30331,N_28240,N_29481);
nand U30332 (N_30332,N_28955,N_27584);
nand U30333 (N_30333,N_28440,N_29520);
or U30334 (N_30334,N_29692,N_28636);
and U30335 (N_30335,N_29459,N_28021);
xnor U30336 (N_30336,N_29863,N_28589);
nor U30337 (N_30337,N_27608,N_29360);
or U30338 (N_30338,N_28775,N_27774);
nand U30339 (N_30339,N_28530,N_29504);
and U30340 (N_30340,N_27549,N_29831);
and U30341 (N_30341,N_29788,N_29639);
xnor U30342 (N_30342,N_29684,N_27740);
nand U30343 (N_30343,N_29084,N_29811);
xor U30344 (N_30344,N_29636,N_27786);
xor U30345 (N_30345,N_27538,N_27583);
and U30346 (N_30346,N_29986,N_29945);
nand U30347 (N_30347,N_27554,N_29868);
nand U30348 (N_30348,N_29696,N_27904);
or U30349 (N_30349,N_28742,N_28078);
or U30350 (N_30350,N_29081,N_28784);
nor U30351 (N_30351,N_28938,N_28853);
nand U30352 (N_30352,N_28206,N_29282);
or U30353 (N_30353,N_28394,N_29856);
or U30354 (N_30354,N_29961,N_28933);
nor U30355 (N_30355,N_27713,N_28771);
xnor U30356 (N_30356,N_27879,N_29865);
xnor U30357 (N_30357,N_28464,N_29421);
or U30358 (N_30358,N_28005,N_29655);
or U30359 (N_30359,N_27815,N_29677);
and U30360 (N_30360,N_28557,N_28523);
nand U30361 (N_30361,N_29427,N_29955);
nor U30362 (N_30362,N_29018,N_29382);
nor U30363 (N_30363,N_29413,N_28065);
and U30364 (N_30364,N_28170,N_28054);
or U30365 (N_30365,N_29031,N_28006);
or U30366 (N_30366,N_29621,N_28182);
xnor U30367 (N_30367,N_29837,N_27527);
nor U30368 (N_30368,N_29198,N_29530);
and U30369 (N_30369,N_28259,N_29307);
nor U30370 (N_30370,N_29514,N_28001);
xor U30371 (N_30371,N_28686,N_28751);
and U30372 (N_30372,N_27886,N_28338);
or U30373 (N_30373,N_29254,N_28402);
and U30374 (N_30374,N_29771,N_28421);
or U30375 (N_30375,N_29314,N_27753);
and U30376 (N_30376,N_29547,N_29220);
nor U30377 (N_30377,N_28449,N_29417);
nor U30378 (N_30378,N_29833,N_28077);
or U30379 (N_30379,N_27719,N_29554);
nor U30380 (N_30380,N_27769,N_27569);
and U30381 (N_30381,N_28101,N_28176);
xor U30382 (N_30382,N_28043,N_29488);
xnor U30383 (N_30383,N_29486,N_29464);
nor U30384 (N_30384,N_27822,N_28582);
nor U30385 (N_30385,N_29088,N_28080);
or U30386 (N_30386,N_28578,N_28284);
xnor U30387 (N_30387,N_29060,N_28909);
nor U30388 (N_30388,N_28061,N_29626);
nand U30389 (N_30389,N_28674,N_27632);
and U30390 (N_30390,N_29278,N_29844);
and U30391 (N_30391,N_27922,N_27624);
and U30392 (N_30392,N_29316,N_28809);
and U30393 (N_30393,N_29824,N_29034);
nor U30394 (N_30394,N_28365,N_27745);
xnor U30395 (N_30395,N_29035,N_28447);
xor U30396 (N_30396,N_28008,N_28109);
nand U30397 (N_30397,N_28174,N_29943);
and U30398 (N_30398,N_28836,N_29739);
nor U30399 (N_30399,N_29949,N_28452);
nor U30400 (N_30400,N_27932,N_27568);
xnor U30401 (N_30401,N_29635,N_27880);
or U30402 (N_30402,N_28201,N_29595);
xnor U30403 (N_30403,N_29761,N_27921);
or U30404 (N_30404,N_29326,N_28881);
or U30405 (N_30405,N_28914,N_29216);
xnor U30406 (N_30406,N_27709,N_28940);
nand U30407 (N_30407,N_28945,N_29450);
nand U30408 (N_30408,N_29938,N_29281);
nand U30409 (N_30409,N_29962,N_28374);
nand U30410 (N_30410,N_28220,N_29052);
nand U30411 (N_30411,N_29581,N_27835);
xnor U30412 (N_30412,N_29877,N_29087);
nand U30413 (N_30413,N_28354,N_27507);
and U30414 (N_30414,N_28698,N_29116);
nor U30415 (N_30415,N_29900,N_27898);
or U30416 (N_30416,N_29012,N_28848);
xnor U30417 (N_30417,N_29537,N_29246);
xor U30418 (N_30418,N_28608,N_28985);
nand U30419 (N_30419,N_28993,N_29171);
xor U30420 (N_30420,N_28288,N_29797);
xor U30421 (N_30421,N_29119,N_28610);
nand U30422 (N_30422,N_29100,N_28468);
xnor U30423 (N_30423,N_28983,N_27618);
and U30424 (N_30424,N_29072,N_28282);
nor U30425 (N_30425,N_27730,N_27690);
nand U30426 (N_30426,N_29227,N_28728);
and U30427 (N_30427,N_28292,N_29338);
xnor U30428 (N_30428,N_29335,N_27874);
nor U30429 (N_30429,N_28739,N_27577);
nand U30430 (N_30430,N_28699,N_28302);
nor U30431 (N_30431,N_28051,N_28336);
nand U30432 (N_30432,N_27944,N_29551);
or U30433 (N_30433,N_29533,N_28720);
nand U30434 (N_30434,N_28678,N_29998);
nand U30435 (N_30435,N_27958,N_29871);
xnor U30436 (N_30436,N_28528,N_29006);
xnor U30437 (N_30437,N_29342,N_28276);
and U30438 (N_30438,N_27696,N_29077);
nand U30439 (N_30439,N_29558,N_27670);
or U30440 (N_30440,N_29579,N_29605);
nor U30441 (N_30441,N_27765,N_29629);
nand U30442 (N_30442,N_29287,N_27759);
nor U30443 (N_30443,N_29428,N_29182);
nand U30444 (N_30444,N_28689,N_29447);
nand U30445 (N_30445,N_27910,N_29936);
nand U30446 (N_30446,N_29359,N_28296);
or U30447 (N_30447,N_27976,N_27615);
nand U30448 (N_30448,N_29691,N_27803);
nand U30449 (N_30449,N_29747,N_28023);
xor U30450 (N_30450,N_27542,N_29027);
xnor U30451 (N_30451,N_27931,N_28944);
nand U30452 (N_30452,N_29120,N_28972);
or U30453 (N_30453,N_28546,N_27547);
and U30454 (N_30454,N_28829,N_29700);
nor U30455 (N_30455,N_28045,N_29260);
and U30456 (N_30456,N_27726,N_29701);
nand U30457 (N_30457,N_28450,N_29429);
nand U30458 (N_30458,N_28347,N_29917);
or U30459 (N_30459,N_28267,N_29454);
and U30460 (N_30460,N_28048,N_28841);
and U30461 (N_30461,N_27573,N_28375);
or U30462 (N_30462,N_29153,N_28262);
nor U30463 (N_30463,N_29353,N_29408);
nor U30464 (N_30464,N_29614,N_28009);
and U30465 (N_30465,N_27971,N_28549);
or U30466 (N_30466,N_27876,N_27911);
xnor U30467 (N_30467,N_27858,N_29981);
xor U30468 (N_30468,N_28015,N_28868);
nand U30469 (N_30469,N_28651,N_29645);
nor U30470 (N_30470,N_28409,N_29678);
or U30471 (N_30471,N_28524,N_27843);
nor U30472 (N_30472,N_27888,N_29310);
and U30473 (N_30473,N_28319,N_28177);
nand U30474 (N_30474,N_27772,N_28272);
or U30475 (N_30475,N_28029,N_27506);
xor U30476 (N_30476,N_29902,N_28633);
or U30477 (N_30477,N_28033,N_29777);
xor U30478 (N_30478,N_28478,N_28704);
nor U30479 (N_30479,N_29688,N_27525);
xor U30480 (N_30480,N_29186,N_27790);
or U30481 (N_30481,N_28607,N_29036);
xor U30482 (N_30482,N_29924,N_29840);
or U30483 (N_30483,N_27831,N_29196);
nand U30484 (N_30484,N_29439,N_28453);
and U30485 (N_30485,N_28831,N_28107);
nor U30486 (N_30486,N_29832,N_27545);
and U30487 (N_30487,N_29667,N_29983);
and U30488 (N_30488,N_28423,N_28193);
and U30489 (N_30489,N_27969,N_27882);
nand U30490 (N_30490,N_28901,N_29959);
or U30491 (N_30491,N_29638,N_28658);
and U30492 (N_30492,N_29143,N_27559);
nor U30493 (N_30493,N_29841,N_28418);
and U30494 (N_30494,N_28156,N_28216);
nor U30495 (N_30495,N_29880,N_28761);
and U30496 (N_30496,N_27897,N_28936);
nand U30497 (N_30497,N_28283,N_27729);
or U30498 (N_30498,N_27727,N_29390);
nor U30499 (N_30499,N_28430,N_29243);
or U30500 (N_30500,N_29987,N_29556);
nand U30501 (N_30501,N_28859,N_27728);
nand U30502 (N_30502,N_28112,N_28326);
or U30503 (N_30503,N_29293,N_27823);
and U30504 (N_30504,N_27682,N_29787);
nor U30505 (N_30505,N_28040,N_29766);
xor U30506 (N_30506,N_28957,N_27675);
or U30507 (N_30507,N_28111,N_28024);
or U30508 (N_30508,N_28339,N_27920);
nand U30509 (N_30509,N_28910,N_29272);
nor U30510 (N_30510,N_28254,N_28103);
and U30511 (N_30511,N_29409,N_29503);
nor U30512 (N_30512,N_27768,N_29003);
nand U30513 (N_30513,N_29516,N_29423);
and U30514 (N_30514,N_27500,N_28186);
or U30515 (N_30515,N_27595,N_29200);
or U30516 (N_30516,N_27836,N_29925);
and U30517 (N_30517,N_29552,N_28181);
xor U30518 (N_30518,N_29673,N_29593);
nor U30519 (N_30519,N_27780,N_27896);
and U30520 (N_30520,N_28014,N_27957);
nand U30521 (N_30521,N_27587,N_27698);
nor U30522 (N_30522,N_28309,N_29368);
or U30523 (N_30523,N_29218,N_28579);
nor U30524 (N_30524,N_29912,N_29322);
nor U30525 (N_30525,N_29472,N_29846);
nand U30526 (N_30526,N_27642,N_28431);
or U30527 (N_30527,N_29358,N_29202);
nor U30528 (N_30528,N_29205,N_29662);
and U30529 (N_30529,N_27679,N_29363);
or U30530 (N_30530,N_28889,N_28599);
and U30531 (N_30531,N_27633,N_28802);
or U30532 (N_30532,N_29808,N_28257);
and U30533 (N_30533,N_28224,N_29578);
xor U30534 (N_30534,N_28136,N_28635);
nor U30535 (N_30535,N_29604,N_28876);
nand U30536 (N_30536,N_29922,N_29461);
xnor U30537 (N_30537,N_28069,N_27883);
and U30538 (N_30538,N_27928,N_29175);
nor U30539 (N_30539,N_27980,N_28422);
nand U30540 (N_30540,N_29590,N_29387);
nand U30541 (N_30541,N_28923,N_29279);
nor U30542 (N_30542,N_28800,N_27846);
nand U30543 (N_30543,N_29803,N_29405);
nand U30544 (N_30544,N_29145,N_28738);
or U30545 (N_30545,N_29487,N_29457);
xor U30546 (N_30546,N_28782,N_27761);
nand U30547 (N_30547,N_27975,N_29001);
xor U30548 (N_30548,N_27787,N_29804);
nand U30549 (N_30549,N_27718,N_29920);
or U30550 (N_30550,N_27865,N_29114);
xor U30551 (N_30551,N_28192,N_28675);
or U30552 (N_30552,N_28939,N_29178);
xor U30553 (N_30553,N_29906,N_27884);
or U30554 (N_30554,N_28390,N_27755);
or U30555 (N_30555,N_29910,N_28459);
nor U30556 (N_30556,N_29250,N_28036);
xor U30557 (N_30557,N_29796,N_29142);
nor U30558 (N_30558,N_29807,N_29467);
and U30559 (N_30559,N_28175,N_29686);
or U30560 (N_30560,N_27917,N_29794);
and U30561 (N_30561,N_29703,N_29789);
and U30562 (N_30562,N_29343,N_29641);
and U30563 (N_30563,N_27658,N_28591);
nand U30564 (N_30564,N_28050,N_29864);
nand U30565 (N_30565,N_28639,N_28151);
xnor U30566 (N_30566,N_27594,N_29659);
nor U30567 (N_30567,N_28797,N_28593);
or U30568 (N_30568,N_29345,N_29809);
nor U30569 (N_30569,N_28746,N_28654);
and U30570 (N_30570,N_28099,N_27655);
nand U30571 (N_30571,N_28653,N_28256);
nand U30572 (N_30572,N_28705,N_29379);
xnor U30573 (N_30573,N_28168,N_28673);
nor U30574 (N_30574,N_28585,N_27712);
nand U30575 (N_30575,N_28491,N_28395);
and U30576 (N_30576,N_28114,N_28743);
or U30577 (N_30577,N_28013,N_27941);
nand U30578 (N_30578,N_28364,N_28554);
nand U30579 (N_30579,N_29536,N_28280);
xor U30580 (N_30580,N_28617,N_29073);
nand U30581 (N_30581,N_28512,N_28499);
and U30582 (N_30582,N_29709,N_28196);
nand U30583 (N_30583,N_28823,N_28753);
and U30584 (N_30584,N_27604,N_29426);
nand U30585 (N_30585,N_28053,N_29968);
nand U30586 (N_30586,N_27637,N_28954);
nor U30587 (N_30587,N_27834,N_27591);
xnor U30588 (N_30588,N_29585,N_29348);
nand U30589 (N_30589,N_27857,N_27974);
nor U30590 (N_30590,N_27801,N_28749);
and U30591 (N_30591,N_27860,N_28072);
and U30592 (N_30592,N_28027,N_28178);
nor U30593 (N_30593,N_29682,N_27785);
or U30594 (N_30594,N_28680,N_28315);
xnor U30595 (N_30595,N_29527,N_28988);
and U30596 (N_30596,N_29724,N_29150);
nand U30597 (N_30597,N_27854,N_27531);
nand U30598 (N_30598,N_29041,N_28318);
xnor U30599 (N_30599,N_29601,N_29103);
or U30600 (N_30600,N_29295,N_28779);
or U30601 (N_30601,N_29315,N_28037);
nand U30602 (N_30602,N_28095,N_27620);
nor U30603 (N_30603,N_29460,N_29933);
nor U30604 (N_30604,N_27563,N_29549);
and U30605 (N_30605,N_29133,N_27802);
or U30606 (N_30606,N_27530,N_27509);
nor U30607 (N_30607,N_27671,N_27961);
or U30608 (N_30608,N_28211,N_27706);
nand U30609 (N_30609,N_27819,N_29894);
nand U30610 (N_30610,N_28890,N_27692);
or U30611 (N_30611,N_28719,N_28533);
or U30612 (N_30612,N_29510,N_28975);
and U30613 (N_30613,N_29194,N_27796);
and U30614 (N_30614,N_29434,N_28584);
and U30615 (N_30615,N_29818,N_28144);
and U30616 (N_30616,N_28714,N_29023);
nor U30617 (N_30617,N_27812,N_28980);
xnor U30618 (N_30618,N_29049,N_28538);
and U30619 (N_30619,N_27930,N_28835);
xor U30620 (N_30620,N_28085,N_29139);
xnor U30621 (N_30621,N_29965,N_27789);
nor U30622 (N_30622,N_28852,N_28540);
or U30623 (N_30623,N_28190,N_27979);
nand U30624 (N_30624,N_29232,N_29620);
or U30625 (N_30625,N_29158,N_29323);
or U30626 (N_30626,N_28962,N_29999);
or U30627 (N_30627,N_27619,N_29513);
xnor U30628 (N_30628,N_28371,N_28229);
or U30629 (N_30629,N_28231,N_28566);
nor U30630 (N_30630,N_28143,N_29535);
and U30631 (N_30631,N_28345,N_29451);
xnor U30632 (N_30632,N_29656,N_29058);
and U30633 (N_30633,N_29258,N_28368);
and U30634 (N_30634,N_28953,N_29853);
xor U30635 (N_30635,N_28644,N_29159);
nor U30636 (N_30636,N_28419,N_29587);
nand U30637 (N_30637,N_28828,N_29101);
nor U30638 (N_30638,N_28748,N_29283);
and U30639 (N_30639,N_29422,N_29324);
and U30640 (N_30640,N_27699,N_29717);
or U30641 (N_30641,N_27562,N_29543);
nand U30642 (N_30642,N_27513,N_29674);
or U30643 (N_30643,N_28766,N_29954);
and U30644 (N_30644,N_28516,N_28268);
nor U30645 (N_30645,N_28388,N_27516);
xor U30646 (N_30646,N_28620,N_28134);
or U30647 (N_30647,N_29996,N_27963);
xor U30648 (N_30648,N_29410,N_29541);
nor U30649 (N_30649,N_29666,N_29308);
nor U30650 (N_30650,N_29573,N_29118);
nand U30651 (N_30651,N_29301,N_29328);
and U30652 (N_30652,N_28382,N_28187);
or U30653 (N_30653,N_29802,N_29525);
and U30654 (N_30654,N_29154,N_27536);
nand U30655 (N_30655,N_28721,N_28787);
nand U30656 (N_30656,N_28812,N_27845);
xnor U30657 (N_30657,N_29608,N_29564);
or U30658 (N_30658,N_28727,N_27680);
xor U30659 (N_30659,N_29571,N_27875);
and U30660 (N_30660,N_29026,N_29505);
xor U30661 (N_30661,N_27580,N_27853);
or U30662 (N_30662,N_27711,N_28420);
nand U30663 (N_30663,N_28716,N_27518);
xnor U30664 (N_30664,N_29599,N_27555);
nand U30665 (N_30665,N_29374,N_29642);
xor U30666 (N_30666,N_27681,N_28035);
and U30667 (N_30667,N_29473,N_29888);
xor U30668 (N_30668,N_28493,N_29588);
or U30669 (N_30669,N_28291,N_28996);
or U30670 (N_30670,N_29572,N_27973);
and U30671 (N_30671,N_28989,N_27638);
xnor U30672 (N_30672,N_28958,N_28562);
and U30673 (N_30673,N_28079,N_29610);
xor U30674 (N_30674,N_27799,N_28762);
xor U30675 (N_30675,N_27627,N_28236);
nand U30676 (N_30676,N_29859,N_28355);
nand U30677 (N_30677,N_29637,N_29442);
xnor U30678 (N_30678,N_29946,N_27757);
xnor U30679 (N_30679,N_28687,N_29372);
nand U30680 (N_30680,N_28501,N_28041);
xnor U30681 (N_30681,N_28113,N_29115);
nor U30682 (N_30682,N_27634,N_28882);
xnor U30683 (N_30683,N_29500,N_28115);
or U30684 (N_30684,N_28392,N_29951);
nand U30685 (N_30685,N_27524,N_27617);
and U30686 (N_30686,N_28623,N_29418);
and U30687 (N_30687,N_28665,N_28969);
xor U30688 (N_30688,N_28071,N_28473);
nor U30689 (N_30689,N_29671,N_27649);
nand U30690 (N_30690,N_27592,N_28555);
nand U30691 (N_30691,N_28403,N_29539);
nor U30692 (N_30692,N_29257,N_27732);
nand U30693 (N_30693,N_27610,N_29916);
nand U30694 (N_30694,N_29456,N_28167);
and U30695 (N_30695,N_28911,N_28715);
and U30696 (N_30696,N_29199,N_29948);
nand U30697 (N_30697,N_28503,N_28790);
and U30698 (N_30698,N_27872,N_28586);
and U30699 (N_30699,N_29755,N_29819);
and U30700 (N_30700,N_27775,N_28084);
nor U30701 (N_30701,N_28656,N_28604);
nor U30702 (N_30702,N_29493,N_29013);
nand U30703 (N_30703,N_29972,N_27825);
nand U30704 (N_30704,N_28184,N_29127);
and U30705 (N_30705,N_29276,N_28601);
nand U30706 (N_30706,N_28320,N_28759);
nand U30707 (N_30707,N_29631,N_29518);
nor U30708 (N_30708,N_27582,N_27738);
nor U30709 (N_30709,N_29000,N_29858);
or U30710 (N_30710,N_29176,N_28871);
nor U30711 (N_30711,N_28487,N_27585);
nand U30712 (N_30712,N_28463,N_29195);
nand U30713 (N_30713,N_28660,N_27942);
or U30714 (N_30714,N_28918,N_29165);
or U30715 (N_30715,N_27502,N_28693);
nand U30716 (N_30716,N_29660,N_28781);
xor U30717 (N_30717,N_28963,N_29208);
nor U30718 (N_30718,N_27522,N_27710);
or U30719 (N_30719,N_29728,N_28233);
nor U30720 (N_30720,N_29122,N_29190);
and U30721 (N_30721,N_29695,N_28750);
xor U30722 (N_30722,N_27660,N_28657);
nand U30723 (N_30723,N_28495,N_29294);
or U30724 (N_30724,N_29370,N_28926);
xnor U30725 (N_30725,N_28706,N_27598);
or U30726 (N_30726,N_28251,N_28153);
nor U30727 (N_30727,N_29529,N_27945);
nor U30728 (N_30728,N_28147,N_28614);
and U30729 (N_30729,N_28241,N_27741);
nor U30730 (N_30730,N_27589,N_29453);
or U30731 (N_30731,N_28138,N_28786);
nand U30732 (N_30732,N_29063,N_28616);
nand U30733 (N_30733,N_28619,N_27950);
nand U30734 (N_30734,N_28760,N_27744);
nand U30735 (N_30735,N_28860,N_28342);
or U30736 (N_30736,N_29974,N_28671);
nand U30737 (N_30737,N_27511,N_29567);
nor U30738 (N_30738,N_28819,N_28864);
and U30739 (N_30739,N_29369,N_29162);
or U30740 (N_30740,N_28558,N_27622);
nor U30741 (N_30741,N_28729,N_28158);
or U30742 (N_30742,N_27998,N_28358);
xor U30743 (N_30743,N_28208,N_28247);
and U30744 (N_30744,N_28708,N_28767);
xor U30745 (N_30745,N_27850,N_28249);
nor U30746 (N_30746,N_28132,N_27505);
xor U30747 (N_30747,N_28898,N_27841);
xor U30748 (N_30748,N_29665,N_28226);
nand U30749 (N_30749,N_28011,N_28696);
or U30750 (N_30750,N_29273,N_28044);
and U30751 (N_30751,N_27864,N_28108);
or U30752 (N_30752,N_27984,N_27605);
and U30753 (N_30753,N_28522,N_28690);
and U30754 (N_30754,N_29446,N_27777);
nand U30755 (N_30755,N_29759,N_29586);
xnor U30756 (N_30756,N_28271,N_28700);
nand U30757 (N_30757,N_27809,N_29545);
nand U30758 (N_30758,N_27999,N_28717);
and U30759 (N_30759,N_29201,N_29879);
nor U30760 (N_30760,N_29540,N_28808);
nand U30761 (N_30761,N_27576,N_28520);
and U30762 (N_30762,N_29805,N_29210);
or U30763 (N_30763,N_27869,N_27702);
and U30764 (N_30764,N_29708,N_28334);
xnor U30765 (N_30765,N_28754,N_29173);
nor U30766 (N_30766,N_29622,N_28612);
nand U30767 (N_30767,N_28986,N_29769);
nor U30768 (N_30768,N_28129,N_27644);
nand U30769 (N_30769,N_27544,N_28611);
nand U30770 (N_30770,N_29284,N_29489);
or U30771 (N_30771,N_29354,N_29104);
xor U30772 (N_30772,N_29580,N_29007);
and U30773 (N_30773,N_29825,N_29785);
and U30774 (N_30774,N_29857,N_27668);
and U30775 (N_30775,N_28603,N_28090);
or U30776 (N_30776,N_29141,N_28935);
or U30777 (N_30777,N_29475,N_29592);
nand U30778 (N_30778,N_29235,N_29269);
or U30779 (N_30779,N_27926,N_28521);
and U30780 (N_30780,N_29262,N_29522);
and U30781 (N_30781,N_29806,N_29402);
or U30782 (N_30782,N_29445,N_29256);
or U30783 (N_30783,N_28117,N_28883);
nand U30784 (N_30784,N_29219,N_29694);
nor U30785 (N_30785,N_29780,N_28592);
or U30786 (N_30786,N_29108,N_28570);
nand U30787 (N_30787,N_29506,N_29437);
and U30788 (N_30788,N_29291,N_29830);
or U30789 (N_30789,N_28100,N_27546);
nand U30790 (N_30790,N_27714,N_27616);
nor U30791 (N_30791,N_28142,N_29921);
xor U30792 (N_30792,N_29155,N_29357);
nor U30793 (N_30793,N_29534,N_27705);
xnor U30794 (N_30794,N_28377,N_28414);
or U30795 (N_30795,N_28813,N_28278);
xor U30796 (N_30796,N_28120,N_28264);
xor U30797 (N_30797,N_29815,N_28640);
nor U30798 (N_30798,N_29737,N_28970);
and U30799 (N_30799,N_28544,N_29632);
nand U30800 (N_30800,N_29538,N_28541);
and U30801 (N_30801,N_28188,N_27890);
and U30802 (N_30802,N_28605,N_27918);
nand U30803 (N_30803,N_27804,N_28016);
and U30804 (N_30804,N_28577,N_28046);
nor U30805 (N_30805,N_29977,N_29240);
xnor U30806 (N_30806,N_29923,N_28627);
nand U30807 (N_30807,N_29252,N_28666);
nand U30808 (N_30808,N_29854,N_29076);
nand U30809 (N_30809,N_28455,N_28682);
nand U30810 (N_30810,N_27565,N_29048);
nor U30811 (N_30811,N_27781,N_27723);
and U30812 (N_30812,N_27795,N_28012);
and U30813 (N_30813,N_29606,N_29704);
nor U30814 (N_30814,N_27735,N_29548);
nand U30815 (N_30815,N_29285,N_28999);
nand U30816 (N_30816,N_28514,N_27811);
and U30817 (N_30817,N_28929,N_29930);
and U30818 (N_30818,N_29583,N_27993);
and U30819 (N_30819,N_29017,N_29891);
nor U30820 (N_30820,N_29664,N_28496);
or U30821 (N_30821,N_28877,N_29044);
xnor U30822 (N_30822,N_27664,N_29020);
and U30823 (N_30823,N_27866,N_27611);
nor U30824 (N_30824,N_29051,N_29090);
nor U30825 (N_30825,N_29928,N_27724);
and U30826 (N_30826,N_28093,N_29043);
or U30827 (N_30827,N_27529,N_29391);
and U30828 (N_30828,N_28180,N_27651);
nand U30829 (N_30829,N_29991,N_28971);
and U30830 (N_30830,N_28679,N_29498);
xnor U30831 (N_30831,N_28140,N_28130);
nor U30832 (N_30832,N_29059,N_27962);
xnor U30833 (N_30833,N_28741,N_28221);
nor U30834 (N_30834,N_28028,N_29680);
nor U30835 (N_30835,N_28152,N_27965);
or U30836 (N_30836,N_29448,N_29732);
nand U30837 (N_30837,N_29399,N_29627);
xor U30838 (N_30838,N_28081,N_28472);
or U30839 (N_30839,N_28350,N_28613);
nor U30840 (N_30840,N_29373,N_29463);
nor U30841 (N_30841,N_27797,N_29756);
and U30842 (N_30842,N_29330,N_28545);
nand U30843 (N_30843,N_29757,N_28321);
xor U30844 (N_30844,N_29298,N_28576);
or U30845 (N_30845,N_29197,N_28314);
nor U30846 (N_30846,N_28432,N_27534);
xnor U30847 (N_30847,N_29265,N_28564);
nand U30848 (N_30848,N_28025,N_28385);
xnor U30849 (N_30849,N_28733,N_28924);
nand U30850 (N_30850,N_28505,N_28337);
nand U30851 (N_30851,N_29166,N_27994);
nand U30852 (N_30852,N_29068,N_27665);
and U30853 (N_30853,N_29929,N_29334);
or U30854 (N_30854,N_27667,N_29065);
xnor U30855 (N_30855,N_29024,N_28811);
xor U30856 (N_30856,N_29947,N_27903);
or U30857 (N_30857,N_28920,N_29255);
or U30858 (N_30858,N_29327,N_29776);
nor U30859 (N_30859,N_29312,N_28857);
or U30860 (N_30860,N_27674,N_27503);
nor U30861 (N_30861,N_28948,N_29217);
and U30862 (N_30862,N_29075,N_28626);
nand U30863 (N_30863,N_28961,N_27909);
nand U30864 (N_30864,N_29025,N_29057);
and U30865 (N_30865,N_28218,N_29376);
nor U30866 (N_30866,N_28968,N_29568);
or U30867 (N_30867,N_27673,N_29569);
nor U30868 (N_30868,N_28232,N_27964);
or U30869 (N_30869,N_29528,N_27600);
xnor U30870 (N_30870,N_28172,N_29230);
and U30871 (N_30871,N_29847,N_27720);
xor U30872 (N_30872,N_28200,N_29798);
xnor U30873 (N_30873,N_29225,N_27937);
nor U30874 (N_30874,N_29814,N_28351);
xnor U30875 (N_30875,N_29117,N_28299);
xnor U30876 (N_30876,N_28285,N_28410);
and U30877 (N_30877,N_28966,N_29918);
nor U30878 (N_30878,N_29288,N_29386);
nand U30879 (N_30879,N_29745,N_28778);
nand U30880 (N_30880,N_29098,N_29236);
nor U30881 (N_30881,N_28396,N_27808);
xnor U30882 (N_30882,N_28286,N_27881);
and U30883 (N_30883,N_28265,N_27725);
and U30884 (N_30884,N_28858,N_28266);
or U30885 (N_30885,N_29318,N_28362);
or U30886 (N_30886,N_29161,N_29953);
xor U30887 (N_30887,N_28250,N_27852);
and U30888 (N_30888,N_29134,N_27887);
nor U30889 (N_30889,N_28903,N_27731);
nor U30890 (N_30890,N_28998,N_29416);
or U30891 (N_30891,N_28799,N_29002);
or U30892 (N_30892,N_28189,N_27601);
xor U30893 (N_30893,N_27628,N_27515);
xor U30894 (N_30894,N_28258,N_28974);
and U30895 (N_30895,N_27701,N_29253);
and U30896 (N_30896,N_29465,N_29319);
xor U30897 (N_30897,N_27599,N_27561);
or U30898 (N_30898,N_28486,N_28820);
nand U30899 (N_30899,N_29206,N_28862);
nor U30900 (N_30900,N_27894,N_28466);
or U30901 (N_30901,N_29485,N_29876);
nand U30902 (N_30902,N_27861,N_27798);
nor U30903 (N_30903,N_27532,N_29392);
or U30904 (N_30904,N_28357,N_28483);
nand U30905 (N_30905,N_27766,N_29786);
nor U30906 (N_30906,N_29346,N_29053);
nor U30907 (N_30907,N_27859,N_29149);
xnor U30908 (N_30908,N_29744,N_27986);
nand U30909 (N_30909,N_29940,N_29377);
xor U30910 (N_30910,N_28683,N_29344);
xnor U30911 (N_30911,N_27939,N_27952);
or U30912 (N_30912,N_29340,N_28128);
xor U30913 (N_30913,N_29042,N_29560);
xnor U30914 (N_30914,N_29137,N_29615);
nand U30915 (N_30915,N_28155,N_28438);
xnor U30916 (N_30916,N_29710,N_27818);
and U30917 (N_30917,N_29658,N_29812);
nand U30918 (N_30918,N_28942,N_29509);
nor U30919 (N_30919,N_28581,N_28451);
and U30920 (N_30920,N_28928,N_28209);
and U30921 (N_30921,N_29751,N_28597);
or U30922 (N_30922,N_29575,N_27540);
or U30923 (N_30923,N_29303,N_28814);
nand U30924 (N_30924,N_28150,N_29729);
and U30925 (N_30925,N_29193,N_29941);
nand U30926 (N_30926,N_29736,N_27708);
nand U30927 (N_30927,N_28332,N_27830);
nor U30928 (N_30928,N_28379,N_29714);
xor U30929 (N_30929,N_27997,N_28145);
or U30930 (N_30930,N_29203,N_28228);
nand U30931 (N_30931,N_29385,N_28649);
xor U30932 (N_30932,N_29110,N_28978);
nand U30933 (N_30933,N_27983,N_29542);
nand U30934 (N_30934,N_29890,N_28925);
xnor U30935 (N_30935,N_28019,N_29973);
and U30936 (N_30936,N_28477,N_28160);
xor U30937 (N_30937,N_29055,N_29299);
or U30938 (N_30938,N_27747,N_28489);
xor U30939 (N_30939,N_29082,N_28003);
or U30940 (N_30940,N_28843,N_28082);
nand U30941 (N_30941,N_28899,N_29479);
or U30942 (N_30942,N_29971,N_27657);
xor U30943 (N_30943,N_29302,N_27892);
xnor U30944 (N_30944,N_29839,N_27749);
xnor U30945 (N_30945,N_29435,N_28270);
or U30946 (N_30946,N_29760,N_27541);
and U30947 (N_30947,N_27933,N_28057);
xnor U30948 (N_30948,N_28973,N_27960);
or U30949 (N_30949,N_29268,N_28734);
nand U30950 (N_30950,N_28244,N_28694);
xor U30951 (N_30951,N_28856,N_27754);
and U30952 (N_30952,N_29248,N_27743);
and U30953 (N_30953,N_28104,N_29054);
and U30954 (N_30954,N_28219,N_28997);
nor U30955 (N_30955,N_28855,N_28896);
xnor U30956 (N_30956,N_29576,N_29029);
xnor U30957 (N_30957,N_28506,N_29474);
nand U30958 (N_30958,N_29096,N_29397);
or U30959 (N_30959,N_27504,N_28684);
xnor U30960 (N_30960,N_28875,N_27829);
nor U30961 (N_30961,N_28571,N_28711);
nand U30962 (N_30962,N_28393,N_29845);
nor U30963 (N_30963,N_29107,N_28230);
and U30964 (N_30964,N_28662,N_28807);
xor U30965 (N_30965,N_28642,N_29039);
or U30966 (N_30966,N_29124,N_29603);
or U30967 (N_30967,N_28324,N_29886);
nor U30968 (N_30968,N_28428,N_28020);
xor U30969 (N_30969,N_27763,N_27678);
and U30970 (N_30970,N_28553,N_29347);
xor U30971 (N_30971,N_28004,N_28329);
or U30972 (N_30972,N_28010,N_28892);
nor U30973 (N_30973,N_29215,N_28615);
nand U30974 (N_30974,N_29975,N_29247);
and U30975 (N_30975,N_29492,N_29404);
nor U30976 (N_30976,N_28648,N_28485);
nor U30977 (N_30977,N_29860,N_28461);
nand U30978 (N_30978,N_28736,N_29725);
xor U30979 (N_30979,N_29764,N_28764);
nor U30980 (N_30980,N_28504,N_29720);
nand U30981 (N_30981,N_28810,N_28793);
or U30982 (N_30982,N_28492,N_28237);
and U30983 (N_30983,N_28780,N_29241);
xnor U30984 (N_30984,N_29280,N_27571);
and U30985 (N_30985,N_28621,N_27839);
or U30986 (N_30986,N_29651,N_28798);
or U30987 (N_30987,N_29297,N_28672);
nor U30988 (N_30988,N_29174,N_28915);
nor U30989 (N_30989,N_27717,N_27817);
and U30990 (N_30990,N_29070,N_28300);
nand U30991 (N_30991,N_28508,N_29080);
or U30992 (N_30992,N_29131,N_29130);
nor U30993 (N_30993,N_27824,N_28565);
xnor U30994 (N_30994,N_28960,N_29721);
xor U30995 (N_30995,N_28785,N_27947);
and U30996 (N_30996,N_27574,N_28702);
nand U30997 (N_30997,N_27981,N_29838);
xor U30998 (N_30998,N_28934,N_27596);
xor U30999 (N_30999,N_27837,N_28163);
nand U31000 (N_31000,N_28803,N_29913);
nor U31001 (N_31001,N_28198,N_28047);
and U31002 (N_31002,N_29767,N_27996);
nand U31003 (N_31003,N_28645,N_27517);
nor U31004 (N_31004,N_29523,N_29412);
nand U31005 (N_31005,N_27539,N_29931);
and U31006 (N_31006,N_29718,N_29244);
xor U31007 (N_31007,N_28308,N_28248);
and U31008 (N_31008,N_27688,N_28346);
nand U31009 (N_31009,N_29985,N_29893);
nor U31010 (N_31010,N_27867,N_28913);
xor U31011 (N_31011,N_29367,N_28951);
nand U31012 (N_31012,N_29495,N_27849);
nor U31013 (N_31013,N_27906,N_28498);
nand U31014 (N_31014,N_28331,N_28400);
and U31015 (N_31015,N_29526,N_29156);
nor U31016 (N_31016,N_29624,N_28981);
xor U31017 (N_31017,N_27683,N_29296);
nor U31018 (N_31018,N_28204,N_29738);
nand U31019 (N_31019,N_27907,N_27929);
or U31020 (N_31020,N_28437,N_28580);
nor U31021 (N_31021,N_29828,N_28681);
nand U31022 (N_31022,N_29889,N_28723);
or U31023 (N_31023,N_29167,N_29935);
and U31024 (N_31024,N_29967,N_29146);
and U31025 (N_31025,N_28732,N_28067);
nor U31026 (N_31026,N_29224,N_28849);
or U31027 (N_31027,N_28441,N_29519);
nand U31028 (N_31028,N_27704,N_28126);
nand U31029 (N_31029,N_29478,N_28724);
and U31030 (N_31030,N_28977,N_29905);
nor U31031 (N_31031,N_27794,N_28290);
or U31032 (N_31032,N_29300,N_28074);
or U31033 (N_31033,N_29577,N_27609);
or U31034 (N_31034,N_27851,N_28908);
xor U31035 (N_31035,N_29799,N_29431);
nor U31036 (N_31036,N_28164,N_28647);
nand U31037 (N_31037,N_28886,N_27597);
nand U31038 (N_31038,N_28872,N_27826);
or U31039 (N_31039,N_28007,N_28275);
nor U31040 (N_31040,N_27572,N_28904);
and U31041 (N_31041,N_28783,N_28991);
and U31042 (N_31042,N_28509,N_29616);
and U31043 (N_31043,N_27685,N_29820);
xnor U31044 (N_31044,N_27967,N_29565);
nor U31045 (N_31045,N_29582,N_29963);
nand U31046 (N_31046,N_29259,N_27607);
or U31047 (N_31047,N_27891,N_29657);
and U31048 (N_31048,N_29019,N_29093);
xnor U31049 (N_31049,N_29697,N_28529);
or U31050 (N_31050,N_29772,N_27695);
nor U31051 (N_31051,N_28425,N_29015);
nand U31052 (N_31052,N_28235,N_28994);
xor U31053 (N_31053,N_29144,N_28446);
or U31054 (N_31054,N_28488,N_28141);
nor U31055 (N_31055,N_27556,N_29425);
and U31056 (N_31056,N_28676,N_27548);
or U31057 (N_31057,N_29713,N_28191);
nand U31058 (N_31058,N_27533,N_28667);
or U31059 (N_31059,N_29005,N_28776);
nand U31060 (N_31060,N_29752,N_28316);
nand U31061 (N_31061,N_27648,N_27773);
xor U31062 (N_31062,N_29329,N_29779);
nor U31063 (N_31063,N_29125,N_28832);
xnor U31064 (N_31064,N_29211,N_28534);
or U31065 (N_31065,N_28110,N_29765);
and U31066 (N_31066,N_27925,N_27535);
nor U31067 (N_31067,N_28335,N_28531);
nand U31068 (N_31068,N_29011,N_29699);
nor U31069 (N_31069,N_29092,N_29861);
or U31070 (N_31070,N_28873,N_28770);
xor U31071 (N_31071,N_29600,N_29597);
nor U31072 (N_31072,N_27847,N_28840);
or U31073 (N_31073,N_28806,N_28203);
nor U31074 (N_31074,N_29740,N_27643);
xnor U31075 (N_31075,N_29826,N_29982);
or U31076 (N_31076,N_28405,N_29349);
and U31077 (N_31077,N_28185,N_28941);
and U31078 (N_31078,N_28661,N_28826);
nor U31079 (N_31079,N_29249,N_27760);
and U31080 (N_31080,N_29037,N_28536);
nor U31081 (N_31081,N_28034,N_28789);
and U31082 (N_31082,N_28556,N_28930);
xnor U31083 (N_31083,N_28943,N_28439);
and U31084 (N_31084,N_28602,N_29690);
xnor U31085 (N_31085,N_27912,N_29365);
or U31086 (N_31086,N_29469,N_28575);
or U31087 (N_31087,N_28773,N_28088);
nor U31088 (N_31088,N_28214,N_29433);
and U31089 (N_31089,N_29619,N_29843);
nand U31090 (N_31090,N_28638,N_29625);
xor U31091 (N_31091,N_29915,N_28269);
and U31092 (N_31092,N_28146,N_29675);
or U31093 (N_31093,N_28227,N_29647);
and U31094 (N_31094,N_28223,N_29793);
xor U31095 (N_31095,N_28293,N_27977);
and U31096 (N_31096,N_27603,N_29187);
or U31097 (N_31097,N_28306,N_29014);
xor U31098 (N_31098,N_28932,N_27868);
nor U31099 (N_31099,N_28588,N_29491);
xor U31100 (N_31100,N_27687,N_29067);
nand U31101 (N_31101,N_29901,N_29562);
or U31102 (N_31102,N_29238,N_29111);
xnor U31103 (N_31103,N_29389,N_29908);
and U31104 (N_31104,N_29852,N_28822);
and U31105 (N_31105,N_29884,N_29508);
nor U31106 (N_31106,N_29267,N_29040);
and U31107 (N_31107,N_28281,N_28415);
and U31108 (N_31108,N_28646,N_28712);
xor U31109 (N_31109,N_28710,N_29702);
nor U31110 (N_31110,N_28404,N_28121);
nand U31111 (N_31111,N_28063,N_29898);
nand U31112 (N_31112,N_29136,N_27792);
nor U31113 (N_31113,N_27693,N_29979);
xnor U31114 (N_31114,N_28755,N_29589);
nor U31115 (N_31115,N_29976,N_28169);
xnor U31116 (N_31116,N_29782,N_29221);
or U31117 (N_31117,N_29032,N_28137);
and U31118 (N_31118,N_29501,N_29517);
or U31119 (N_31119,N_28480,N_27782);
and U31120 (N_31120,N_27800,N_29618);
or U31121 (N_31121,N_28179,N_27521);
nor U31122 (N_31122,N_29226,N_29179);
nor U31123 (N_31123,N_28032,N_28458);
nand U31124 (N_31124,N_28118,N_28567);
xor U31125 (N_31125,N_27938,N_28885);
nor U31126 (N_31126,N_28479,N_27526);
xnor U31127 (N_31127,N_28381,N_27703);
xnor U31128 (N_31128,N_28038,N_29557);
nand U31129 (N_31129,N_29598,N_28992);
or U31130 (N_31130,N_28830,N_28097);
nand U31131 (N_31131,N_28384,N_27715);
nor U31132 (N_31132,N_28225,N_28273);
or U31133 (N_31133,N_28165,N_28879);
xnor U31134 (N_31134,N_29496,N_27936);
xnor U31135 (N_31135,N_29393,N_27923);
and U31136 (N_31136,N_28411,N_27810);
nor U31137 (N_31137,N_28677,N_29138);
and U31138 (N_31138,N_28794,N_27558);
nand U31139 (N_31139,N_28287,N_29004);
nand U31140 (N_31140,N_28730,N_28663);
xnor U31141 (N_31141,N_27838,N_28083);
xnor U31142 (N_31142,N_28070,N_29183);
or U31143 (N_31143,N_28707,N_28833);
and U31144 (N_31144,N_28370,N_27951);
xnor U31145 (N_31145,N_29056,N_28215);
nor U31146 (N_31146,N_29038,N_29078);
nand U31147 (N_31147,N_27689,N_29444);
or U31148 (N_31148,N_29482,N_29407);
nor U31149 (N_31149,N_29237,N_29499);
or U31150 (N_31150,N_27805,N_29304);
and U31151 (N_31151,N_27827,N_29045);
nor U31152 (N_31152,N_29157,N_29834);
nor U31153 (N_31153,N_28827,N_27856);
and U31154 (N_31154,N_29477,N_29867);
or U31155 (N_31155,N_29532,N_28805);
and U31156 (N_31156,N_29722,N_28092);
nor U31157 (N_31157,N_27927,N_27656);
or U31158 (N_31158,N_29290,N_27813);
xnor U31159 (N_31159,N_28361,N_29129);
nor U31160 (N_31160,N_29795,N_28162);
xnor U31161 (N_31161,N_29222,N_28098);
and U31162 (N_31162,N_29438,N_28821);
nand U31163 (N_31163,N_28884,N_28442);
xor U31164 (N_31164,N_29816,N_29228);
nor U31165 (N_31165,N_28094,N_27806);
nand U31166 (N_31166,N_28289,N_28427);
nand U31167 (N_31167,N_28058,N_29132);
nand U31168 (N_31168,N_28433,N_27840);
and U31169 (N_31169,N_29375,N_27551);
nor U31170 (N_31170,N_28456,N_29774);
nor U31171 (N_31171,N_27606,N_29992);
nand U31172 (N_31172,N_28417,N_28340);
and U31173 (N_31173,N_28328,N_29669);
and U31174 (N_31174,N_27901,N_28664);
nand U31175 (N_31175,N_29264,N_28171);
nand U31176 (N_31176,N_27666,N_27877);
nor U31177 (N_31177,N_27756,N_29899);
and U31178 (N_31178,N_29406,N_28207);
xor U31179 (N_31179,N_29511,N_29792);
and U31180 (N_31180,N_29458,N_28552);
nand U31181 (N_31181,N_27621,N_27784);
and U31182 (N_31182,N_28195,N_28922);
nand U31183 (N_31183,N_27820,N_28692);
or U31184 (N_31184,N_28561,N_29957);
and U31185 (N_31185,N_29046,N_27878);
and U31186 (N_31186,N_27871,N_28310);
and U31187 (N_31187,N_28788,N_28159);
nand U31188 (N_31188,N_27640,N_29140);
and U31189 (N_31189,N_28260,N_28242);
nand U31190 (N_31190,N_28497,N_28413);
or U31191 (N_31191,N_29047,N_27914);
nand U31192 (N_31192,N_28341,N_27748);
nor U31193 (N_31193,N_28535,N_29449);
nor U31194 (N_31194,N_28086,N_28116);
xor U31195 (N_31195,N_29213,N_29271);
and U31196 (N_31196,N_28838,N_28574);
or U31197 (N_31197,N_28194,N_29394);
nand U31198 (N_31198,N_28353,N_29102);
or U31199 (N_31199,N_29715,N_28837);
nor U31200 (N_31200,N_29850,N_29734);
xor U31201 (N_31201,N_29234,N_29242);
or U31202 (N_31202,N_29069,N_28344);
nor U31203 (N_31203,N_27672,N_28887);
nor U31204 (N_31204,N_29566,N_29851);
nand U31205 (N_31205,N_29550,N_29097);
xor U31206 (N_31206,N_28426,N_29748);
nor U31207 (N_31207,N_28166,N_29128);
nand U31208 (N_31208,N_28921,N_28106);
or U31209 (N_31209,N_28122,N_27510);
xnor U31210 (N_31210,N_27519,N_28632);
xnor U31211 (N_31211,N_28629,N_28757);
nand U31212 (N_31212,N_28587,N_28303);
nor U31213 (N_31213,N_27862,N_29741);
and U31214 (N_31214,N_27736,N_27623);
nand U31215 (N_31215,N_28525,N_27528);
xor U31216 (N_31216,N_29919,N_29927);
xor U31217 (N_31217,N_27716,N_29978);
or U31218 (N_31218,N_28818,N_29596);
nand U31219 (N_31219,N_29723,N_28527);
and U31220 (N_31220,N_29942,N_27523);
nand U31221 (N_31221,N_29261,N_27902);
or U31222 (N_31222,N_29471,N_29233);
and U31223 (N_31223,N_29687,N_29683);
xor U31224 (N_31224,N_28042,N_29350);
xor U31225 (N_31225,N_29753,N_28825);
nand U31226 (N_31226,N_28630,N_28327);
xor U31227 (N_31227,N_27770,N_28246);
and U31228 (N_31228,N_29646,N_29185);
nor U31229 (N_31229,N_28916,N_29168);
and U31230 (N_31230,N_27895,N_28234);
xor U31231 (N_31231,N_28173,N_28718);
and U31232 (N_31232,N_29706,N_28865);
and U31233 (N_31233,N_29352,N_27764);
nand U31234 (N_31234,N_28670,N_27855);
nand U31235 (N_31235,N_28590,N_27934);
or U31236 (N_31236,N_29574,N_29364);
or U31237 (N_31237,N_29633,N_29810);
or U31238 (N_31238,N_29336,N_29822);
and U31239 (N_31239,N_29204,N_28560);
nand U31240 (N_31240,N_28161,N_29800);
or U31241 (N_31241,N_28448,N_28139);
xnor U31242 (N_31242,N_28984,N_28537);
and U31243 (N_31243,N_29231,N_28469);
or U31244 (N_31244,N_28952,N_29952);
or U31245 (N_31245,N_27970,N_27567);
xor U31246 (N_31246,N_29064,N_29163);
or U31247 (N_31247,N_29964,N_29309);
xor U31248 (N_31248,N_28912,N_28956);
nor U31249 (N_31249,N_29546,N_28210);
nor U31250 (N_31250,N_29142,N_29881);
xnor U31251 (N_31251,N_27590,N_29441);
and U31252 (N_31252,N_28567,N_28622);
nand U31253 (N_31253,N_28767,N_27597);
nor U31254 (N_31254,N_28069,N_29673);
and U31255 (N_31255,N_27766,N_29356);
nand U31256 (N_31256,N_28305,N_28045);
and U31257 (N_31257,N_28298,N_29216);
nand U31258 (N_31258,N_29103,N_28868);
nor U31259 (N_31259,N_28539,N_29742);
and U31260 (N_31260,N_28862,N_28246);
nor U31261 (N_31261,N_27658,N_28036);
nor U31262 (N_31262,N_27642,N_29273);
nor U31263 (N_31263,N_28392,N_29803);
xor U31264 (N_31264,N_27945,N_27628);
or U31265 (N_31265,N_27951,N_28447);
xor U31266 (N_31266,N_27717,N_27853);
nand U31267 (N_31267,N_29184,N_27608);
and U31268 (N_31268,N_27855,N_29504);
or U31269 (N_31269,N_28679,N_27636);
and U31270 (N_31270,N_29758,N_28085);
or U31271 (N_31271,N_29086,N_29683);
nor U31272 (N_31272,N_29951,N_28735);
nor U31273 (N_31273,N_29861,N_27649);
and U31274 (N_31274,N_28442,N_28560);
nor U31275 (N_31275,N_29628,N_29614);
nand U31276 (N_31276,N_27702,N_29732);
and U31277 (N_31277,N_29201,N_27734);
or U31278 (N_31278,N_27822,N_28177);
or U31279 (N_31279,N_29852,N_28755);
and U31280 (N_31280,N_28466,N_29843);
nand U31281 (N_31281,N_28098,N_28825);
xnor U31282 (N_31282,N_28752,N_28475);
or U31283 (N_31283,N_29963,N_29024);
nand U31284 (N_31284,N_28844,N_27943);
xnor U31285 (N_31285,N_28309,N_29495);
and U31286 (N_31286,N_28742,N_27679);
nor U31287 (N_31287,N_29258,N_28776);
or U31288 (N_31288,N_29054,N_27969);
or U31289 (N_31289,N_27628,N_29634);
or U31290 (N_31290,N_29067,N_29496);
nor U31291 (N_31291,N_29869,N_27781);
nand U31292 (N_31292,N_28553,N_27841);
nand U31293 (N_31293,N_29812,N_28646);
nand U31294 (N_31294,N_29870,N_29470);
xnor U31295 (N_31295,N_29141,N_29323);
xor U31296 (N_31296,N_29094,N_29034);
and U31297 (N_31297,N_28892,N_28328);
or U31298 (N_31298,N_27994,N_27728);
nand U31299 (N_31299,N_29166,N_27979);
nand U31300 (N_31300,N_28631,N_29626);
nand U31301 (N_31301,N_28994,N_28473);
and U31302 (N_31302,N_28106,N_29691);
xnor U31303 (N_31303,N_29554,N_27863);
nand U31304 (N_31304,N_28967,N_28961);
and U31305 (N_31305,N_28536,N_29958);
nand U31306 (N_31306,N_27958,N_27819);
nor U31307 (N_31307,N_29271,N_28819);
nand U31308 (N_31308,N_28777,N_29243);
or U31309 (N_31309,N_27650,N_29267);
nor U31310 (N_31310,N_27821,N_27833);
xor U31311 (N_31311,N_27839,N_29432);
nand U31312 (N_31312,N_27707,N_29382);
and U31313 (N_31313,N_28378,N_29712);
xor U31314 (N_31314,N_27862,N_28433);
and U31315 (N_31315,N_28710,N_27903);
or U31316 (N_31316,N_29540,N_27707);
or U31317 (N_31317,N_29635,N_28792);
nor U31318 (N_31318,N_28446,N_27796);
or U31319 (N_31319,N_29278,N_29138);
or U31320 (N_31320,N_29300,N_29049);
or U31321 (N_31321,N_28464,N_27892);
nand U31322 (N_31322,N_29188,N_27844);
nand U31323 (N_31323,N_29038,N_28616);
nor U31324 (N_31324,N_27861,N_28817);
nor U31325 (N_31325,N_28314,N_29947);
xnor U31326 (N_31326,N_29056,N_29380);
xnor U31327 (N_31327,N_28275,N_28703);
xor U31328 (N_31328,N_28593,N_28551);
or U31329 (N_31329,N_29470,N_29150);
or U31330 (N_31330,N_29438,N_28877);
or U31331 (N_31331,N_27814,N_28173);
xor U31332 (N_31332,N_29202,N_29568);
or U31333 (N_31333,N_29529,N_29192);
nor U31334 (N_31334,N_29671,N_29349);
xor U31335 (N_31335,N_27890,N_28480);
xor U31336 (N_31336,N_29651,N_29202);
xor U31337 (N_31337,N_27844,N_28972);
nand U31338 (N_31338,N_29911,N_27998);
nor U31339 (N_31339,N_29884,N_29158);
nor U31340 (N_31340,N_27834,N_27760);
nor U31341 (N_31341,N_28655,N_28380);
or U31342 (N_31342,N_28523,N_29647);
nor U31343 (N_31343,N_27624,N_29601);
nand U31344 (N_31344,N_29897,N_28405);
xor U31345 (N_31345,N_28521,N_27998);
nor U31346 (N_31346,N_28301,N_27676);
xnor U31347 (N_31347,N_28215,N_29923);
and U31348 (N_31348,N_29751,N_29525);
xnor U31349 (N_31349,N_29269,N_27771);
and U31350 (N_31350,N_28808,N_29022);
nor U31351 (N_31351,N_27728,N_28198);
nand U31352 (N_31352,N_29802,N_28876);
xnor U31353 (N_31353,N_29873,N_27794);
and U31354 (N_31354,N_29595,N_29315);
nor U31355 (N_31355,N_27639,N_27634);
nand U31356 (N_31356,N_28488,N_28454);
nor U31357 (N_31357,N_27942,N_29273);
nor U31358 (N_31358,N_28797,N_29183);
and U31359 (N_31359,N_29527,N_29433);
xor U31360 (N_31360,N_28893,N_27725);
xnor U31361 (N_31361,N_29159,N_27547);
or U31362 (N_31362,N_29101,N_27598);
nor U31363 (N_31363,N_29313,N_29777);
xnor U31364 (N_31364,N_29887,N_28238);
and U31365 (N_31365,N_28349,N_29714);
or U31366 (N_31366,N_28199,N_27694);
or U31367 (N_31367,N_29563,N_29659);
or U31368 (N_31368,N_28260,N_28836);
nor U31369 (N_31369,N_28011,N_28098);
or U31370 (N_31370,N_29316,N_28097);
xnor U31371 (N_31371,N_27815,N_29660);
and U31372 (N_31372,N_29253,N_27695);
nand U31373 (N_31373,N_28665,N_28960);
nor U31374 (N_31374,N_29418,N_28485);
xnor U31375 (N_31375,N_27964,N_29405);
nand U31376 (N_31376,N_28560,N_27671);
xor U31377 (N_31377,N_28028,N_28563);
xnor U31378 (N_31378,N_29657,N_28693);
xnor U31379 (N_31379,N_29821,N_27781);
nor U31380 (N_31380,N_29985,N_27672);
nand U31381 (N_31381,N_28774,N_29883);
xnor U31382 (N_31382,N_29384,N_28246);
nor U31383 (N_31383,N_27601,N_27815);
xor U31384 (N_31384,N_29580,N_29821);
nor U31385 (N_31385,N_27840,N_29957);
nand U31386 (N_31386,N_28312,N_29273);
nand U31387 (N_31387,N_27507,N_27504);
nand U31388 (N_31388,N_28742,N_28007);
xnor U31389 (N_31389,N_29181,N_29619);
or U31390 (N_31390,N_28229,N_27870);
xnor U31391 (N_31391,N_27509,N_28944);
nor U31392 (N_31392,N_29825,N_29000);
and U31393 (N_31393,N_28653,N_28523);
or U31394 (N_31394,N_29953,N_29901);
xnor U31395 (N_31395,N_28786,N_29761);
nand U31396 (N_31396,N_27902,N_28174);
xor U31397 (N_31397,N_28935,N_29953);
and U31398 (N_31398,N_28116,N_29615);
nand U31399 (N_31399,N_29572,N_29454);
xnor U31400 (N_31400,N_27944,N_28981);
xnor U31401 (N_31401,N_27880,N_28075);
nand U31402 (N_31402,N_27776,N_28013);
nand U31403 (N_31403,N_28344,N_29829);
nand U31404 (N_31404,N_28622,N_28539);
nor U31405 (N_31405,N_29812,N_27889);
xnor U31406 (N_31406,N_28532,N_28744);
or U31407 (N_31407,N_28248,N_29075);
xnor U31408 (N_31408,N_28072,N_27882);
or U31409 (N_31409,N_29108,N_28440);
xnor U31410 (N_31410,N_28803,N_29904);
or U31411 (N_31411,N_27505,N_27668);
nand U31412 (N_31412,N_27911,N_27788);
nand U31413 (N_31413,N_27886,N_29914);
or U31414 (N_31414,N_27848,N_28143);
nor U31415 (N_31415,N_28784,N_29129);
or U31416 (N_31416,N_29602,N_29250);
nor U31417 (N_31417,N_29467,N_27968);
and U31418 (N_31418,N_29635,N_28310);
nor U31419 (N_31419,N_28057,N_28317);
xnor U31420 (N_31420,N_28640,N_28423);
nor U31421 (N_31421,N_28675,N_28687);
nor U31422 (N_31422,N_27990,N_29787);
xnor U31423 (N_31423,N_29612,N_27512);
nand U31424 (N_31424,N_27650,N_28758);
or U31425 (N_31425,N_28290,N_29604);
nand U31426 (N_31426,N_27551,N_28386);
xor U31427 (N_31427,N_28214,N_28529);
nor U31428 (N_31428,N_29315,N_28631);
nand U31429 (N_31429,N_28036,N_28721);
nand U31430 (N_31430,N_29011,N_29955);
and U31431 (N_31431,N_28539,N_29484);
or U31432 (N_31432,N_28740,N_28350);
and U31433 (N_31433,N_29534,N_29444);
nor U31434 (N_31434,N_29590,N_29580);
and U31435 (N_31435,N_29465,N_29949);
or U31436 (N_31436,N_27762,N_28714);
and U31437 (N_31437,N_28081,N_29494);
nor U31438 (N_31438,N_29206,N_29530);
and U31439 (N_31439,N_29444,N_29242);
nor U31440 (N_31440,N_28715,N_27757);
nor U31441 (N_31441,N_28448,N_29310);
xnor U31442 (N_31442,N_29271,N_27663);
or U31443 (N_31443,N_27628,N_27898);
nand U31444 (N_31444,N_29943,N_29650);
nand U31445 (N_31445,N_29479,N_29355);
and U31446 (N_31446,N_29022,N_28800);
or U31447 (N_31447,N_29790,N_29158);
nor U31448 (N_31448,N_28557,N_28142);
and U31449 (N_31449,N_29063,N_28022);
nand U31450 (N_31450,N_28464,N_27934);
xnor U31451 (N_31451,N_29926,N_27638);
nor U31452 (N_31452,N_28758,N_29764);
xnor U31453 (N_31453,N_29745,N_29167);
xnor U31454 (N_31454,N_27857,N_28338);
nand U31455 (N_31455,N_28246,N_28192);
or U31456 (N_31456,N_28469,N_29804);
xnor U31457 (N_31457,N_29790,N_28628);
xor U31458 (N_31458,N_28941,N_29989);
or U31459 (N_31459,N_28652,N_29219);
or U31460 (N_31460,N_29797,N_28868);
and U31461 (N_31461,N_28323,N_27994);
nor U31462 (N_31462,N_28242,N_28075);
xor U31463 (N_31463,N_28816,N_27910);
nor U31464 (N_31464,N_28457,N_27600);
nand U31465 (N_31465,N_29256,N_27558);
and U31466 (N_31466,N_29189,N_29814);
and U31467 (N_31467,N_27781,N_28547);
or U31468 (N_31468,N_29015,N_29260);
xnor U31469 (N_31469,N_27670,N_28669);
and U31470 (N_31470,N_28470,N_29103);
and U31471 (N_31471,N_29209,N_29163);
xnor U31472 (N_31472,N_27647,N_28714);
nor U31473 (N_31473,N_27725,N_29851);
and U31474 (N_31474,N_29874,N_29508);
xnor U31475 (N_31475,N_29541,N_29078);
xor U31476 (N_31476,N_28522,N_28195);
nand U31477 (N_31477,N_29145,N_28853);
nor U31478 (N_31478,N_27641,N_28000);
xnor U31479 (N_31479,N_29116,N_27964);
nand U31480 (N_31480,N_28009,N_28766);
xnor U31481 (N_31481,N_28248,N_27941);
xor U31482 (N_31482,N_28737,N_29754);
nand U31483 (N_31483,N_27955,N_29240);
nand U31484 (N_31484,N_29851,N_27566);
nand U31485 (N_31485,N_29791,N_29817);
or U31486 (N_31486,N_28482,N_29398);
and U31487 (N_31487,N_29281,N_29544);
xor U31488 (N_31488,N_29672,N_29894);
or U31489 (N_31489,N_29122,N_27777);
and U31490 (N_31490,N_29239,N_27983);
xnor U31491 (N_31491,N_28280,N_28656);
nor U31492 (N_31492,N_28245,N_28007);
or U31493 (N_31493,N_28150,N_29738);
nand U31494 (N_31494,N_28692,N_28270);
and U31495 (N_31495,N_29219,N_28935);
and U31496 (N_31496,N_27919,N_28500);
nor U31497 (N_31497,N_29905,N_28286);
and U31498 (N_31498,N_28192,N_29806);
and U31499 (N_31499,N_29431,N_29403);
nand U31500 (N_31500,N_28908,N_29680);
or U31501 (N_31501,N_28023,N_28004);
and U31502 (N_31502,N_28463,N_29446);
xnor U31503 (N_31503,N_29481,N_28096);
nor U31504 (N_31504,N_29516,N_29632);
nand U31505 (N_31505,N_28998,N_28634);
or U31506 (N_31506,N_28256,N_28962);
xor U31507 (N_31507,N_28713,N_27663);
xor U31508 (N_31508,N_28001,N_29405);
and U31509 (N_31509,N_27808,N_28029);
xor U31510 (N_31510,N_29802,N_28822);
xnor U31511 (N_31511,N_28423,N_29232);
or U31512 (N_31512,N_29894,N_28264);
and U31513 (N_31513,N_28801,N_27556);
nand U31514 (N_31514,N_28665,N_28326);
and U31515 (N_31515,N_27683,N_27800);
nand U31516 (N_31516,N_29899,N_29282);
and U31517 (N_31517,N_29251,N_27776);
nand U31518 (N_31518,N_29686,N_29775);
or U31519 (N_31519,N_29727,N_29102);
and U31520 (N_31520,N_29692,N_28235);
nor U31521 (N_31521,N_28410,N_28812);
or U31522 (N_31522,N_29001,N_28030);
and U31523 (N_31523,N_28480,N_29132);
nand U31524 (N_31524,N_29282,N_28867);
xor U31525 (N_31525,N_28159,N_28059);
nand U31526 (N_31526,N_27708,N_27961);
and U31527 (N_31527,N_28414,N_28892);
nand U31528 (N_31528,N_28426,N_29019);
xor U31529 (N_31529,N_28081,N_29469);
and U31530 (N_31530,N_28516,N_28812);
nor U31531 (N_31531,N_29660,N_28181);
nand U31532 (N_31532,N_27574,N_28522);
and U31533 (N_31533,N_28793,N_29373);
nand U31534 (N_31534,N_29503,N_29697);
xnor U31535 (N_31535,N_28974,N_28176);
xor U31536 (N_31536,N_28123,N_28217);
xnor U31537 (N_31537,N_27529,N_27579);
and U31538 (N_31538,N_29140,N_28717);
and U31539 (N_31539,N_29375,N_29066);
xor U31540 (N_31540,N_28291,N_28710);
or U31541 (N_31541,N_29036,N_29280);
and U31542 (N_31542,N_27986,N_29203);
or U31543 (N_31543,N_28094,N_28866);
nor U31544 (N_31544,N_28044,N_28794);
nor U31545 (N_31545,N_29834,N_29407);
nand U31546 (N_31546,N_29655,N_28531);
and U31547 (N_31547,N_28955,N_28075);
and U31548 (N_31548,N_28943,N_29756);
nand U31549 (N_31549,N_28822,N_28738);
nor U31550 (N_31550,N_28460,N_28517);
or U31551 (N_31551,N_28677,N_28590);
xnor U31552 (N_31552,N_28743,N_27646);
xnor U31553 (N_31553,N_29727,N_28704);
xor U31554 (N_31554,N_27891,N_29084);
nand U31555 (N_31555,N_29045,N_28746);
xnor U31556 (N_31556,N_29883,N_27568);
or U31557 (N_31557,N_27770,N_28898);
nor U31558 (N_31558,N_27541,N_28658);
nor U31559 (N_31559,N_29376,N_28157);
nand U31560 (N_31560,N_28842,N_28026);
and U31561 (N_31561,N_27926,N_29962);
and U31562 (N_31562,N_27758,N_29833);
nand U31563 (N_31563,N_28252,N_29944);
nand U31564 (N_31564,N_27616,N_28667);
nand U31565 (N_31565,N_28360,N_29223);
and U31566 (N_31566,N_28722,N_28740);
nor U31567 (N_31567,N_29397,N_28109);
nand U31568 (N_31568,N_28271,N_28633);
or U31569 (N_31569,N_28339,N_29202);
nand U31570 (N_31570,N_29700,N_28871);
or U31571 (N_31571,N_29992,N_28994);
nand U31572 (N_31572,N_29147,N_29934);
nand U31573 (N_31573,N_28425,N_27539);
nand U31574 (N_31574,N_29784,N_27721);
nor U31575 (N_31575,N_28585,N_28374);
or U31576 (N_31576,N_29964,N_27738);
or U31577 (N_31577,N_28652,N_29138);
xnor U31578 (N_31578,N_28804,N_28700);
xor U31579 (N_31579,N_28592,N_29407);
and U31580 (N_31580,N_28744,N_28598);
or U31581 (N_31581,N_28426,N_29582);
xor U31582 (N_31582,N_29564,N_27847);
or U31583 (N_31583,N_29682,N_27829);
xor U31584 (N_31584,N_29535,N_29426);
nor U31585 (N_31585,N_28752,N_27730);
xnor U31586 (N_31586,N_28491,N_28894);
and U31587 (N_31587,N_29742,N_27561);
or U31588 (N_31588,N_28970,N_28769);
and U31589 (N_31589,N_29245,N_28884);
xor U31590 (N_31590,N_27873,N_29244);
xnor U31591 (N_31591,N_28076,N_28367);
xnor U31592 (N_31592,N_29189,N_28786);
nand U31593 (N_31593,N_29077,N_27586);
and U31594 (N_31594,N_28550,N_27695);
nand U31595 (N_31595,N_29767,N_28927);
or U31596 (N_31596,N_28825,N_28221);
and U31597 (N_31597,N_29062,N_28232);
or U31598 (N_31598,N_28239,N_29282);
xor U31599 (N_31599,N_28087,N_29520);
or U31600 (N_31600,N_27847,N_28540);
xor U31601 (N_31601,N_29119,N_27963);
xnor U31602 (N_31602,N_28115,N_29835);
or U31603 (N_31603,N_28385,N_29796);
nor U31604 (N_31604,N_28626,N_27763);
nor U31605 (N_31605,N_27576,N_29678);
nor U31606 (N_31606,N_28245,N_28483);
nor U31607 (N_31607,N_27876,N_28333);
xnor U31608 (N_31608,N_27626,N_28959);
and U31609 (N_31609,N_29414,N_27675);
and U31610 (N_31610,N_28533,N_28857);
or U31611 (N_31611,N_29567,N_29465);
and U31612 (N_31612,N_29121,N_29734);
nor U31613 (N_31613,N_29603,N_29905);
xor U31614 (N_31614,N_29006,N_28354);
or U31615 (N_31615,N_29216,N_28257);
and U31616 (N_31616,N_28336,N_28335);
nor U31617 (N_31617,N_28804,N_27861);
and U31618 (N_31618,N_28724,N_29765);
xnor U31619 (N_31619,N_27742,N_28332);
nand U31620 (N_31620,N_28317,N_29416);
nor U31621 (N_31621,N_29018,N_29023);
nand U31622 (N_31622,N_29413,N_28973);
nand U31623 (N_31623,N_29658,N_28785);
and U31624 (N_31624,N_28277,N_27547);
or U31625 (N_31625,N_29717,N_28942);
xnor U31626 (N_31626,N_28807,N_28758);
and U31627 (N_31627,N_28970,N_28036);
nand U31628 (N_31628,N_29692,N_28732);
xnor U31629 (N_31629,N_28459,N_29603);
xor U31630 (N_31630,N_28858,N_27693);
xnor U31631 (N_31631,N_28009,N_27850);
nand U31632 (N_31632,N_28666,N_29137);
or U31633 (N_31633,N_29450,N_27887);
nor U31634 (N_31634,N_29557,N_28587);
xor U31635 (N_31635,N_28994,N_28260);
xor U31636 (N_31636,N_27816,N_28834);
nand U31637 (N_31637,N_28867,N_28053);
nor U31638 (N_31638,N_29726,N_29325);
nor U31639 (N_31639,N_29651,N_29616);
and U31640 (N_31640,N_28241,N_28771);
and U31641 (N_31641,N_28907,N_29769);
nand U31642 (N_31642,N_28276,N_28416);
xnor U31643 (N_31643,N_28224,N_28220);
and U31644 (N_31644,N_29889,N_28825);
nor U31645 (N_31645,N_27766,N_28441);
nand U31646 (N_31646,N_29070,N_29781);
nand U31647 (N_31647,N_28199,N_27836);
nor U31648 (N_31648,N_27633,N_28554);
nor U31649 (N_31649,N_28705,N_28939);
nor U31650 (N_31650,N_29407,N_29158);
and U31651 (N_31651,N_29155,N_29902);
xor U31652 (N_31652,N_29450,N_28824);
nor U31653 (N_31653,N_29932,N_28755);
and U31654 (N_31654,N_29308,N_27663);
and U31655 (N_31655,N_28071,N_29929);
or U31656 (N_31656,N_27646,N_29657);
xor U31657 (N_31657,N_28611,N_29485);
nor U31658 (N_31658,N_29193,N_27667);
and U31659 (N_31659,N_28509,N_29203);
nor U31660 (N_31660,N_29140,N_28260);
nor U31661 (N_31661,N_29578,N_28346);
and U31662 (N_31662,N_27781,N_28132);
nor U31663 (N_31663,N_29782,N_29512);
or U31664 (N_31664,N_29736,N_29937);
nor U31665 (N_31665,N_28573,N_29601);
nand U31666 (N_31666,N_29822,N_27756);
xor U31667 (N_31667,N_28104,N_29311);
or U31668 (N_31668,N_28286,N_29278);
nand U31669 (N_31669,N_29804,N_28581);
or U31670 (N_31670,N_29619,N_28850);
or U31671 (N_31671,N_27973,N_27917);
nand U31672 (N_31672,N_29852,N_28297);
nand U31673 (N_31673,N_29768,N_27896);
xnor U31674 (N_31674,N_28915,N_29239);
or U31675 (N_31675,N_28809,N_28666);
or U31676 (N_31676,N_28957,N_28511);
or U31677 (N_31677,N_28636,N_28021);
nand U31678 (N_31678,N_28058,N_28639);
and U31679 (N_31679,N_28744,N_29315);
nor U31680 (N_31680,N_29821,N_28248);
nand U31681 (N_31681,N_28857,N_28879);
xor U31682 (N_31682,N_27798,N_27932);
xnor U31683 (N_31683,N_29383,N_27971);
xnor U31684 (N_31684,N_29936,N_27553);
or U31685 (N_31685,N_28621,N_27955);
or U31686 (N_31686,N_28236,N_28952);
or U31687 (N_31687,N_29985,N_29551);
and U31688 (N_31688,N_29376,N_28434);
nand U31689 (N_31689,N_28583,N_28955);
nor U31690 (N_31690,N_29256,N_27842);
or U31691 (N_31691,N_29497,N_28020);
xnor U31692 (N_31692,N_27623,N_28504);
and U31693 (N_31693,N_29137,N_28167);
nand U31694 (N_31694,N_28765,N_29136);
nor U31695 (N_31695,N_27872,N_28048);
nor U31696 (N_31696,N_28144,N_27779);
or U31697 (N_31697,N_27919,N_29180);
and U31698 (N_31698,N_27734,N_29142);
nor U31699 (N_31699,N_29696,N_29047);
and U31700 (N_31700,N_28098,N_28326);
xnor U31701 (N_31701,N_29472,N_28304);
or U31702 (N_31702,N_28685,N_28966);
nor U31703 (N_31703,N_29492,N_27857);
nand U31704 (N_31704,N_27916,N_28534);
or U31705 (N_31705,N_29308,N_29193);
and U31706 (N_31706,N_29239,N_28979);
and U31707 (N_31707,N_28517,N_28656);
nand U31708 (N_31708,N_29604,N_28224);
or U31709 (N_31709,N_27866,N_29526);
xnor U31710 (N_31710,N_29637,N_27612);
nor U31711 (N_31711,N_28436,N_27974);
and U31712 (N_31712,N_28767,N_27595);
and U31713 (N_31713,N_27685,N_29587);
xor U31714 (N_31714,N_27783,N_28411);
nand U31715 (N_31715,N_28132,N_27992);
and U31716 (N_31716,N_28461,N_27672);
or U31717 (N_31717,N_29419,N_29171);
nor U31718 (N_31718,N_27801,N_29129);
xnor U31719 (N_31719,N_29059,N_28110);
nor U31720 (N_31720,N_28912,N_28114);
nor U31721 (N_31721,N_27810,N_29662);
nand U31722 (N_31722,N_29457,N_27787);
or U31723 (N_31723,N_28894,N_28013);
and U31724 (N_31724,N_29039,N_29214);
or U31725 (N_31725,N_29352,N_28377);
nor U31726 (N_31726,N_27720,N_29605);
nand U31727 (N_31727,N_28321,N_29925);
nand U31728 (N_31728,N_28546,N_28674);
nand U31729 (N_31729,N_28332,N_28011);
and U31730 (N_31730,N_28483,N_29833);
nand U31731 (N_31731,N_29956,N_29986);
xor U31732 (N_31732,N_28287,N_27781);
nor U31733 (N_31733,N_28827,N_28878);
or U31734 (N_31734,N_27523,N_28916);
or U31735 (N_31735,N_27977,N_29577);
nor U31736 (N_31736,N_28197,N_29726);
xor U31737 (N_31737,N_29568,N_27828);
and U31738 (N_31738,N_29436,N_29618);
xor U31739 (N_31739,N_28948,N_27762);
and U31740 (N_31740,N_28769,N_29230);
nand U31741 (N_31741,N_29330,N_28765);
nor U31742 (N_31742,N_28764,N_29983);
and U31743 (N_31743,N_28024,N_28274);
xnor U31744 (N_31744,N_27609,N_27823);
nor U31745 (N_31745,N_27670,N_29165);
or U31746 (N_31746,N_27752,N_29228);
xnor U31747 (N_31747,N_29666,N_29060);
xor U31748 (N_31748,N_27639,N_29408);
or U31749 (N_31749,N_28011,N_28376);
nand U31750 (N_31750,N_27801,N_29374);
and U31751 (N_31751,N_29338,N_28049);
nor U31752 (N_31752,N_27818,N_28647);
or U31753 (N_31753,N_28218,N_28224);
nand U31754 (N_31754,N_29717,N_28278);
nand U31755 (N_31755,N_27900,N_28978);
and U31756 (N_31756,N_28636,N_28352);
nor U31757 (N_31757,N_28290,N_27640);
nand U31758 (N_31758,N_27827,N_27577);
and U31759 (N_31759,N_28609,N_28371);
nand U31760 (N_31760,N_28572,N_28447);
or U31761 (N_31761,N_28267,N_27552);
xor U31762 (N_31762,N_29354,N_29250);
nor U31763 (N_31763,N_28496,N_28595);
nor U31764 (N_31764,N_29385,N_29460);
or U31765 (N_31765,N_28534,N_29336);
and U31766 (N_31766,N_28628,N_27869);
or U31767 (N_31767,N_29826,N_28062);
or U31768 (N_31768,N_29872,N_29891);
xor U31769 (N_31769,N_29652,N_27724);
nand U31770 (N_31770,N_27556,N_28611);
and U31771 (N_31771,N_27848,N_28795);
and U31772 (N_31772,N_28681,N_28939);
or U31773 (N_31773,N_29708,N_28121);
and U31774 (N_31774,N_27821,N_29905);
or U31775 (N_31775,N_27969,N_29281);
and U31776 (N_31776,N_29480,N_29825);
nand U31777 (N_31777,N_29355,N_29516);
and U31778 (N_31778,N_27887,N_28295);
or U31779 (N_31779,N_27517,N_27557);
nor U31780 (N_31780,N_27612,N_29283);
and U31781 (N_31781,N_27838,N_29123);
xnor U31782 (N_31782,N_28427,N_29239);
nand U31783 (N_31783,N_27640,N_29645);
nand U31784 (N_31784,N_29905,N_29654);
nand U31785 (N_31785,N_29254,N_28711);
and U31786 (N_31786,N_29692,N_29627);
nor U31787 (N_31787,N_28983,N_28678);
xor U31788 (N_31788,N_29481,N_28741);
xnor U31789 (N_31789,N_28326,N_27919);
nand U31790 (N_31790,N_27660,N_27858);
or U31791 (N_31791,N_28606,N_28105);
or U31792 (N_31792,N_28388,N_28672);
nand U31793 (N_31793,N_29324,N_27895);
nor U31794 (N_31794,N_29215,N_29098);
or U31795 (N_31795,N_29421,N_29924);
nand U31796 (N_31796,N_29651,N_28723);
or U31797 (N_31797,N_28918,N_29243);
nand U31798 (N_31798,N_29550,N_28766);
and U31799 (N_31799,N_29625,N_28272);
or U31800 (N_31800,N_28392,N_28627);
and U31801 (N_31801,N_29188,N_27555);
nor U31802 (N_31802,N_29716,N_28471);
and U31803 (N_31803,N_28643,N_29377);
nand U31804 (N_31804,N_27776,N_29555);
nand U31805 (N_31805,N_28961,N_29534);
and U31806 (N_31806,N_27586,N_28394);
and U31807 (N_31807,N_28768,N_29555);
or U31808 (N_31808,N_27830,N_29838);
and U31809 (N_31809,N_28807,N_28441);
xnor U31810 (N_31810,N_28556,N_28417);
or U31811 (N_31811,N_27886,N_28186);
or U31812 (N_31812,N_29803,N_29676);
xor U31813 (N_31813,N_27679,N_28985);
xor U31814 (N_31814,N_27543,N_27836);
nor U31815 (N_31815,N_28013,N_28196);
and U31816 (N_31816,N_27875,N_28832);
nand U31817 (N_31817,N_27710,N_27806);
and U31818 (N_31818,N_29172,N_28683);
nand U31819 (N_31819,N_27750,N_28456);
or U31820 (N_31820,N_28489,N_28026);
xnor U31821 (N_31821,N_29404,N_29082);
or U31822 (N_31822,N_28933,N_27904);
nand U31823 (N_31823,N_28541,N_28723);
nor U31824 (N_31824,N_28113,N_28303);
and U31825 (N_31825,N_29692,N_29830);
xnor U31826 (N_31826,N_28973,N_29842);
xor U31827 (N_31827,N_29968,N_28004);
and U31828 (N_31828,N_28685,N_27936);
nand U31829 (N_31829,N_28503,N_27606);
or U31830 (N_31830,N_29460,N_29849);
nor U31831 (N_31831,N_29005,N_27953);
nand U31832 (N_31832,N_29289,N_28026);
nand U31833 (N_31833,N_29568,N_27539);
and U31834 (N_31834,N_27682,N_29021);
or U31835 (N_31835,N_28089,N_28208);
xor U31836 (N_31836,N_28147,N_29717);
nand U31837 (N_31837,N_29095,N_28843);
or U31838 (N_31838,N_28056,N_27843);
nor U31839 (N_31839,N_27571,N_29042);
and U31840 (N_31840,N_29627,N_28339);
xnor U31841 (N_31841,N_29723,N_27777);
xnor U31842 (N_31842,N_29286,N_29281);
xor U31843 (N_31843,N_27743,N_29148);
nand U31844 (N_31844,N_27775,N_29097);
nor U31845 (N_31845,N_27555,N_29414);
nor U31846 (N_31846,N_29012,N_27711);
and U31847 (N_31847,N_29261,N_28328);
xor U31848 (N_31848,N_27904,N_27707);
xor U31849 (N_31849,N_28461,N_29815);
or U31850 (N_31850,N_29923,N_29952);
xnor U31851 (N_31851,N_27522,N_29998);
nor U31852 (N_31852,N_29520,N_28716);
xnor U31853 (N_31853,N_29463,N_27590);
nor U31854 (N_31854,N_28017,N_28966);
nor U31855 (N_31855,N_29838,N_28789);
nor U31856 (N_31856,N_28588,N_28637);
and U31857 (N_31857,N_27599,N_29243);
and U31858 (N_31858,N_28867,N_29717);
xor U31859 (N_31859,N_29363,N_27894);
and U31860 (N_31860,N_29412,N_29066);
or U31861 (N_31861,N_28229,N_29067);
and U31862 (N_31862,N_29438,N_29597);
and U31863 (N_31863,N_28404,N_29361);
xor U31864 (N_31864,N_27613,N_28446);
xor U31865 (N_31865,N_28537,N_29382);
and U31866 (N_31866,N_29754,N_28795);
and U31867 (N_31867,N_27858,N_28734);
xnor U31868 (N_31868,N_29151,N_28368);
and U31869 (N_31869,N_28400,N_29952);
or U31870 (N_31870,N_28040,N_29293);
xor U31871 (N_31871,N_29026,N_29387);
xnor U31872 (N_31872,N_29985,N_29292);
nor U31873 (N_31873,N_29074,N_27646);
and U31874 (N_31874,N_28064,N_29828);
xnor U31875 (N_31875,N_28772,N_27664);
nor U31876 (N_31876,N_27701,N_29388);
nor U31877 (N_31877,N_27658,N_28504);
nand U31878 (N_31878,N_28991,N_29350);
nand U31879 (N_31879,N_27977,N_27961);
and U31880 (N_31880,N_27933,N_27938);
nand U31881 (N_31881,N_28659,N_29121);
and U31882 (N_31882,N_29143,N_28796);
or U31883 (N_31883,N_29095,N_29704);
xor U31884 (N_31884,N_29596,N_28379);
or U31885 (N_31885,N_29850,N_29980);
xnor U31886 (N_31886,N_29775,N_29804);
xor U31887 (N_31887,N_29442,N_29499);
nand U31888 (N_31888,N_27771,N_28683);
xnor U31889 (N_31889,N_28304,N_29798);
and U31890 (N_31890,N_28093,N_28575);
or U31891 (N_31891,N_27970,N_28356);
or U31892 (N_31892,N_29437,N_29405);
nor U31893 (N_31893,N_29428,N_28949);
nor U31894 (N_31894,N_28265,N_29785);
or U31895 (N_31895,N_28832,N_28926);
or U31896 (N_31896,N_28309,N_27935);
and U31897 (N_31897,N_28686,N_27749);
xnor U31898 (N_31898,N_28790,N_28464);
xnor U31899 (N_31899,N_29666,N_29442);
or U31900 (N_31900,N_27528,N_28094);
and U31901 (N_31901,N_28961,N_29029);
or U31902 (N_31902,N_29293,N_28816);
and U31903 (N_31903,N_29501,N_29344);
xnor U31904 (N_31904,N_28541,N_28557);
nor U31905 (N_31905,N_27696,N_29131);
nor U31906 (N_31906,N_28903,N_28098);
xnor U31907 (N_31907,N_29085,N_28892);
and U31908 (N_31908,N_29051,N_28107);
nand U31909 (N_31909,N_28096,N_28077);
xor U31910 (N_31910,N_27913,N_29562);
nor U31911 (N_31911,N_29182,N_28656);
xnor U31912 (N_31912,N_29411,N_29453);
xor U31913 (N_31913,N_29288,N_28847);
nand U31914 (N_31914,N_27591,N_28161);
xor U31915 (N_31915,N_28957,N_28656);
or U31916 (N_31916,N_27719,N_27706);
and U31917 (N_31917,N_27552,N_28508);
xor U31918 (N_31918,N_28384,N_28906);
and U31919 (N_31919,N_28354,N_28752);
and U31920 (N_31920,N_27806,N_28315);
or U31921 (N_31921,N_28539,N_28542);
or U31922 (N_31922,N_28943,N_28588);
or U31923 (N_31923,N_28795,N_28522);
nor U31924 (N_31924,N_27930,N_28148);
or U31925 (N_31925,N_28260,N_29692);
or U31926 (N_31926,N_27818,N_27779);
nor U31927 (N_31927,N_28624,N_29630);
and U31928 (N_31928,N_28649,N_29450);
xor U31929 (N_31929,N_29137,N_28047);
xor U31930 (N_31930,N_29781,N_29260);
or U31931 (N_31931,N_28031,N_28320);
nor U31932 (N_31932,N_28033,N_29327);
or U31933 (N_31933,N_27859,N_29244);
nand U31934 (N_31934,N_28678,N_28885);
xnor U31935 (N_31935,N_29852,N_27757);
nand U31936 (N_31936,N_28878,N_27732);
xnor U31937 (N_31937,N_29298,N_29143);
xor U31938 (N_31938,N_27501,N_27811);
and U31939 (N_31939,N_28651,N_28184);
or U31940 (N_31940,N_27676,N_29508);
xnor U31941 (N_31941,N_27879,N_29238);
nor U31942 (N_31942,N_28440,N_27586);
xor U31943 (N_31943,N_28728,N_28140);
nor U31944 (N_31944,N_27816,N_28853);
nor U31945 (N_31945,N_29857,N_27574);
nand U31946 (N_31946,N_28716,N_28165);
and U31947 (N_31947,N_28988,N_29055);
or U31948 (N_31948,N_27623,N_29102);
and U31949 (N_31949,N_29363,N_28632);
nand U31950 (N_31950,N_29586,N_27810);
nor U31951 (N_31951,N_27819,N_28180);
nand U31952 (N_31952,N_27891,N_29197);
xor U31953 (N_31953,N_28561,N_28611);
xor U31954 (N_31954,N_29820,N_28523);
and U31955 (N_31955,N_28548,N_28962);
or U31956 (N_31956,N_29234,N_28262);
nand U31957 (N_31957,N_29293,N_27742);
nor U31958 (N_31958,N_28705,N_27995);
xor U31959 (N_31959,N_29611,N_28398);
xor U31960 (N_31960,N_29264,N_27907);
nor U31961 (N_31961,N_28412,N_28234);
nor U31962 (N_31962,N_29061,N_28032);
or U31963 (N_31963,N_28003,N_28180);
nor U31964 (N_31964,N_27608,N_28548);
and U31965 (N_31965,N_28928,N_27823);
nand U31966 (N_31966,N_29617,N_29859);
or U31967 (N_31967,N_28566,N_28723);
nor U31968 (N_31968,N_28620,N_28544);
nor U31969 (N_31969,N_29103,N_28919);
nor U31970 (N_31970,N_29398,N_28874);
nand U31971 (N_31971,N_27659,N_28208);
and U31972 (N_31972,N_27980,N_29125);
nand U31973 (N_31973,N_28723,N_29968);
xor U31974 (N_31974,N_29805,N_27694);
nand U31975 (N_31975,N_29328,N_27950);
xnor U31976 (N_31976,N_27583,N_29325);
xor U31977 (N_31977,N_29917,N_29516);
xnor U31978 (N_31978,N_28142,N_29324);
and U31979 (N_31979,N_29638,N_27575);
nor U31980 (N_31980,N_29830,N_28906);
or U31981 (N_31981,N_27695,N_29255);
or U31982 (N_31982,N_28650,N_27838);
xor U31983 (N_31983,N_29457,N_29936);
xor U31984 (N_31984,N_27580,N_28075);
xnor U31985 (N_31985,N_29305,N_28199);
nor U31986 (N_31986,N_28311,N_28976);
and U31987 (N_31987,N_29370,N_29642);
or U31988 (N_31988,N_29664,N_29907);
nand U31989 (N_31989,N_27913,N_28756);
nor U31990 (N_31990,N_28420,N_28456);
nand U31991 (N_31991,N_29944,N_28586);
or U31992 (N_31992,N_27601,N_29954);
or U31993 (N_31993,N_29758,N_29983);
nand U31994 (N_31994,N_28277,N_29047);
and U31995 (N_31995,N_29313,N_28068);
and U31996 (N_31996,N_29979,N_28632);
nor U31997 (N_31997,N_29840,N_28899);
nand U31998 (N_31998,N_29149,N_28343);
nand U31999 (N_31999,N_29613,N_28468);
or U32000 (N_32000,N_28119,N_29570);
and U32001 (N_32001,N_29923,N_28970);
nor U32002 (N_32002,N_29624,N_29692);
xnor U32003 (N_32003,N_28858,N_27593);
xor U32004 (N_32004,N_28438,N_27638);
and U32005 (N_32005,N_27945,N_29445);
and U32006 (N_32006,N_29746,N_28895);
and U32007 (N_32007,N_27636,N_29049);
nor U32008 (N_32008,N_27726,N_29333);
nand U32009 (N_32009,N_28080,N_28272);
nand U32010 (N_32010,N_27831,N_28841);
xor U32011 (N_32011,N_29920,N_27723);
or U32012 (N_32012,N_27902,N_29691);
nor U32013 (N_32013,N_28850,N_29523);
xor U32014 (N_32014,N_29833,N_29056);
nand U32015 (N_32015,N_29199,N_27592);
nor U32016 (N_32016,N_29283,N_28581);
and U32017 (N_32017,N_28706,N_29542);
and U32018 (N_32018,N_27529,N_29475);
xor U32019 (N_32019,N_27798,N_29703);
and U32020 (N_32020,N_28430,N_28563);
or U32021 (N_32021,N_29827,N_29604);
nor U32022 (N_32022,N_29097,N_27711);
or U32023 (N_32023,N_28111,N_29387);
or U32024 (N_32024,N_29917,N_28805);
or U32025 (N_32025,N_29143,N_29144);
or U32026 (N_32026,N_28423,N_28248);
nand U32027 (N_32027,N_29434,N_28254);
xnor U32028 (N_32028,N_29803,N_29324);
nor U32029 (N_32029,N_29102,N_28070);
xnor U32030 (N_32030,N_27740,N_27957);
or U32031 (N_32031,N_29426,N_29505);
nor U32032 (N_32032,N_28462,N_29122);
xor U32033 (N_32033,N_29239,N_29994);
nand U32034 (N_32034,N_28752,N_29363);
nand U32035 (N_32035,N_27841,N_27913);
xor U32036 (N_32036,N_27998,N_28044);
nor U32037 (N_32037,N_28696,N_27660);
nand U32038 (N_32038,N_28431,N_28443);
nor U32039 (N_32039,N_28501,N_27683);
nand U32040 (N_32040,N_27557,N_29430);
xnor U32041 (N_32041,N_27814,N_27548);
xnor U32042 (N_32042,N_29123,N_29153);
or U32043 (N_32043,N_29224,N_28144);
xor U32044 (N_32044,N_29035,N_27668);
nor U32045 (N_32045,N_28220,N_29729);
and U32046 (N_32046,N_29395,N_29323);
nand U32047 (N_32047,N_28467,N_29416);
xnor U32048 (N_32048,N_28696,N_29015);
nor U32049 (N_32049,N_28618,N_27855);
and U32050 (N_32050,N_29236,N_28116);
or U32051 (N_32051,N_28607,N_28346);
xor U32052 (N_32052,N_29545,N_29489);
nor U32053 (N_32053,N_28428,N_29476);
nand U32054 (N_32054,N_29419,N_29249);
and U32055 (N_32055,N_29379,N_29070);
nor U32056 (N_32056,N_28649,N_28417);
or U32057 (N_32057,N_28930,N_28883);
nor U32058 (N_32058,N_28915,N_29374);
nor U32059 (N_32059,N_29840,N_29479);
xor U32060 (N_32060,N_28112,N_28013);
nand U32061 (N_32061,N_29599,N_28135);
xnor U32062 (N_32062,N_29062,N_27609);
or U32063 (N_32063,N_28134,N_28344);
xnor U32064 (N_32064,N_29810,N_27662);
nor U32065 (N_32065,N_28203,N_27892);
and U32066 (N_32066,N_28016,N_27821);
nor U32067 (N_32067,N_29765,N_29790);
nor U32068 (N_32068,N_28409,N_29249);
nand U32069 (N_32069,N_27765,N_29810);
or U32070 (N_32070,N_28440,N_27529);
and U32071 (N_32071,N_28410,N_29544);
nor U32072 (N_32072,N_29137,N_28753);
or U32073 (N_32073,N_28761,N_28643);
or U32074 (N_32074,N_29332,N_28416);
or U32075 (N_32075,N_29762,N_27740);
nand U32076 (N_32076,N_28539,N_28627);
or U32077 (N_32077,N_28136,N_29238);
nor U32078 (N_32078,N_28204,N_28211);
nor U32079 (N_32079,N_28052,N_29987);
xnor U32080 (N_32080,N_29967,N_27657);
nand U32081 (N_32081,N_28424,N_28724);
and U32082 (N_32082,N_29097,N_28185);
and U32083 (N_32083,N_28958,N_27927);
nand U32084 (N_32084,N_29604,N_29239);
or U32085 (N_32085,N_27682,N_29124);
xor U32086 (N_32086,N_27985,N_28919);
nor U32087 (N_32087,N_29907,N_29593);
nand U32088 (N_32088,N_28545,N_28086);
nand U32089 (N_32089,N_27560,N_28718);
nand U32090 (N_32090,N_27748,N_29657);
or U32091 (N_32091,N_27599,N_27551);
xor U32092 (N_32092,N_28085,N_29739);
xor U32093 (N_32093,N_29618,N_29784);
or U32094 (N_32094,N_29035,N_29840);
nand U32095 (N_32095,N_29185,N_27504);
and U32096 (N_32096,N_27515,N_28211);
xnor U32097 (N_32097,N_29703,N_29771);
and U32098 (N_32098,N_28772,N_27698);
xor U32099 (N_32099,N_27882,N_27862);
xnor U32100 (N_32100,N_29748,N_28576);
or U32101 (N_32101,N_29132,N_28774);
or U32102 (N_32102,N_28572,N_28079);
xnor U32103 (N_32103,N_29114,N_28252);
or U32104 (N_32104,N_28521,N_29648);
and U32105 (N_32105,N_28874,N_29076);
and U32106 (N_32106,N_29318,N_27508);
or U32107 (N_32107,N_29479,N_28087);
nand U32108 (N_32108,N_27607,N_29239);
or U32109 (N_32109,N_29828,N_27713);
or U32110 (N_32110,N_27958,N_28182);
nor U32111 (N_32111,N_29569,N_27593);
nor U32112 (N_32112,N_29311,N_29993);
xnor U32113 (N_32113,N_28122,N_29511);
and U32114 (N_32114,N_27563,N_29501);
and U32115 (N_32115,N_28292,N_27608);
nor U32116 (N_32116,N_29862,N_29152);
and U32117 (N_32117,N_28849,N_29346);
and U32118 (N_32118,N_29446,N_29449);
nand U32119 (N_32119,N_29580,N_28869);
nor U32120 (N_32120,N_27922,N_27787);
or U32121 (N_32121,N_29443,N_29090);
and U32122 (N_32122,N_28181,N_29248);
and U32123 (N_32123,N_28481,N_28960);
or U32124 (N_32124,N_28595,N_29985);
nor U32125 (N_32125,N_29364,N_28551);
nand U32126 (N_32126,N_27964,N_28095);
or U32127 (N_32127,N_29838,N_28066);
xnor U32128 (N_32128,N_28557,N_27702);
xor U32129 (N_32129,N_28304,N_29453);
or U32130 (N_32130,N_27942,N_29726);
or U32131 (N_32131,N_29300,N_29267);
or U32132 (N_32132,N_29050,N_28032);
xnor U32133 (N_32133,N_27853,N_28854);
or U32134 (N_32134,N_28554,N_29043);
nor U32135 (N_32135,N_28440,N_27753);
or U32136 (N_32136,N_29647,N_27537);
and U32137 (N_32137,N_29108,N_29299);
nand U32138 (N_32138,N_29646,N_28565);
xnor U32139 (N_32139,N_29702,N_27863);
and U32140 (N_32140,N_29119,N_28148);
xnor U32141 (N_32141,N_28053,N_28690);
or U32142 (N_32142,N_28064,N_29898);
or U32143 (N_32143,N_28633,N_29444);
or U32144 (N_32144,N_29782,N_28007);
nand U32145 (N_32145,N_29116,N_28953);
nand U32146 (N_32146,N_27849,N_27594);
or U32147 (N_32147,N_27627,N_28850);
xor U32148 (N_32148,N_29360,N_27610);
or U32149 (N_32149,N_28095,N_29354);
nand U32150 (N_32150,N_29716,N_28825);
xor U32151 (N_32151,N_27755,N_28626);
or U32152 (N_32152,N_29300,N_29880);
nand U32153 (N_32153,N_28980,N_28101);
nand U32154 (N_32154,N_27840,N_27852);
xnor U32155 (N_32155,N_28135,N_29240);
or U32156 (N_32156,N_29465,N_28978);
nand U32157 (N_32157,N_28992,N_29146);
nor U32158 (N_32158,N_29095,N_27759);
nor U32159 (N_32159,N_28817,N_28694);
nor U32160 (N_32160,N_28483,N_27636);
nand U32161 (N_32161,N_27913,N_27813);
nand U32162 (N_32162,N_27636,N_29130);
xnor U32163 (N_32163,N_29879,N_27864);
nand U32164 (N_32164,N_29449,N_29102);
and U32165 (N_32165,N_28888,N_27833);
and U32166 (N_32166,N_29933,N_28969);
nor U32167 (N_32167,N_29129,N_29195);
xor U32168 (N_32168,N_28233,N_28500);
and U32169 (N_32169,N_27765,N_29313);
nor U32170 (N_32170,N_28585,N_28447);
nor U32171 (N_32171,N_28870,N_27911);
and U32172 (N_32172,N_28315,N_28707);
nor U32173 (N_32173,N_29308,N_29068);
or U32174 (N_32174,N_27541,N_27843);
nand U32175 (N_32175,N_27540,N_29512);
xor U32176 (N_32176,N_28856,N_28813);
nor U32177 (N_32177,N_28376,N_27774);
or U32178 (N_32178,N_27963,N_28520);
or U32179 (N_32179,N_28960,N_29194);
or U32180 (N_32180,N_28358,N_28027);
nor U32181 (N_32181,N_29597,N_29372);
nand U32182 (N_32182,N_28676,N_28334);
and U32183 (N_32183,N_29367,N_29890);
nor U32184 (N_32184,N_28392,N_28738);
and U32185 (N_32185,N_28630,N_27655);
and U32186 (N_32186,N_29212,N_27590);
or U32187 (N_32187,N_28955,N_29547);
and U32188 (N_32188,N_27529,N_29376);
nor U32189 (N_32189,N_29005,N_27671);
and U32190 (N_32190,N_28392,N_29473);
nand U32191 (N_32191,N_28719,N_28459);
or U32192 (N_32192,N_27685,N_29968);
xnor U32193 (N_32193,N_27530,N_28277);
nand U32194 (N_32194,N_29285,N_29014);
nor U32195 (N_32195,N_28034,N_29379);
nor U32196 (N_32196,N_29189,N_29231);
nand U32197 (N_32197,N_29792,N_28021);
nand U32198 (N_32198,N_28471,N_29288);
and U32199 (N_32199,N_27681,N_29501);
and U32200 (N_32200,N_28443,N_29408);
xnor U32201 (N_32201,N_27910,N_28821);
and U32202 (N_32202,N_29300,N_27789);
and U32203 (N_32203,N_27798,N_29003);
or U32204 (N_32204,N_27717,N_27939);
nor U32205 (N_32205,N_28318,N_29660);
nor U32206 (N_32206,N_29794,N_28270);
or U32207 (N_32207,N_29790,N_29470);
and U32208 (N_32208,N_29717,N_28725);
nand U32209 (N_32209,N_27898,N_28854);
xnor U32210 (N_32210,N_28397,N_27529);
xor U32211 (N_32211,N_29069,N_29627);
or U32212 (N_32212,N_27964,N_28056);
or U32213 (N_32213,N_28717,N_29157);
nand U32214 (N_32214,N_27962,N_28990);
xnor U32215 (N_32215,N_28579,N_28222);
or U32216 (N_32216,N_27530,N_29284);
nand U32217 (N_32217,N_29026,N_27899);
nor U32218 (N_32218,N_28641,N_28763);
nand U32219 (N_32219,N_29666,N_27717);
nand U32220 (N_32220,N_27698,N_29157);
xor U32221 (N_32221,N_28301,N_27893);
and U32222 (N_32222,N_29991,N_28796);
xnor U32223 (N_32223,N_29081,N_28506);
or U32224 (N_32224,N_29182,N_27750);
or U32225 (N_32225,N_29689,N_29293);
or U32226 (N_32226,N_29799,N_28697);
nand U32227 (N_32227,N_27800,N_29156);
nor U32228 (N_32228,N_28810,N_28650);
nand U32229 (N_32229,N_29356,N_27700);
or U32230 (N_32230,N_29499,N_28032);
nand U32231 (N_32231,N_29509,N_27823);
or U32232 (N_32232,N_29292,N_29570);
xor U32233 (N_32233,N_29318,N_29988);
nor U32234 (N_32234,N_28584,N_28341);
nor U32235 (N_32235,N_29791,N_29810);
or U32236 (N_32236,N_29725,N_27873);
xor U32237 (N_32237,N_29829,N_28820);
nand U32238 (N_32238,N_28313,N_28636);
and U32239 (N_32239,N_29080,N_28065);
nor U32240 (N_32240,N_29012,N_29993);
nand U32241 (N_32241,N_27716,N_28515);
nand U32242 (N_32242,N_27676,N_28077);
nor U32243 (N_32243,N_29152,N_28163);
nand U32244 (N_32244,N_29834,N_29510);
and U32245 (N_32245,N_29654,N_28370);
nand U32246 (N_32246,N_27500,N_28368);
nor U32247 (N_32247,N_28395,N_29424);
nor U32248 (N_32248,N_29320,N_28370);
and U32249 (N_32249,N_27893,N_27754);
nor U32250 (N_32250,N_27677,N_28544);
nor U32251 (N_32251,N_28423,N_27799);
nor U32252 (N_32252,N_28688,N_29497);
xnor U32253 (N_32253,N_28557,N_28488);
or U32254 (N_32254,N_29650,N_29807);
nor U32255 (N_32255,N_28435,N_28295);
nor U32256 (N_32256,N_28271,N_28485);
or U32257 (N_32257,N_28658,N_28126);
xnor U32258 (N_32258,N_29356,N_29470);
xor U32259 (N_32259,N_28730,N_28553);
xor U32260 (N_32260,N_27745,N_28551);
nor U32261 (N_32261,N_28566,N_29324);
xor U32262 (N_32262,N_28051,N_29991);
or U32263 (N_32263,N_28249,N_29046);
or U32264 (N_32264,N_27974,N_29338);
nor U32265 (N_32265,N_28395,N_28614);
or U32266 (N_32266,N_29990,N_28166);
xor U32267 (N_32267,N_29549,N_28218);
nor U32268 (N_32268,N_29677,N_29690);
and U32269 (N_32269,N_27860,N_27539);
nor U32270 (N_32270,N_27997,N_28391);
nand U32271 (N_32271,N_28036,N_27552);
or U32272 (N_32272,N_29192,N_29623);
nand U32273 (N_32273,N_28516,N_29072);
xor U32274 (N_32274,N_28269,N_29047);
nor U32275 (N_32275,N_28633,N_29962);
nor U32276 (N_32276,N_29927,N_27951);
xor U32277 (N_32277,N_29393,N_28750);
nand U32278 (N_32278,N_28355,N_28618);
xnor U32279 (N_32279,N_28061,N_28714);
or U32280 (N_32280,N_28873,N_27825);
or U32281 (N_32281,N_27800,N_29565);
nor U32282 (N_32282,N_27819,N_29762);
xor U32283 (N_32283,N_28101,N_27975);
or U32284 (N_32284,N_27971,N_28156);
nor U32285 (N_32285,N_27838,N_29475);
nand U32286 (N_32286,N_28754,N_29479);
nand U32287 (N_32287,N_28397,N_29764);
nor U32288 (N_32288,N_29045,N_28011);
nor U32289 (N_32289,N_28564,N_29773);
and U32290 (N_32290,N_29819,N_27758);
xnor U32291 (N_32291,N_28264,N_28792);
xor U32292 (N_32292,N_29899,N_29372);
or U32293 (N_32293,N_28841,N_28069);
or U32294 (N_32294,N_29116,N_29500);
or U32295 (N_32295,N_29629,N_29835);
or U32296 (N_32296,N_28165,N_28876);
and U32297 (N_32297,N_29215,N_29903);
xnor U32298 (N_32298,N_29241,N_27720);
nand U32299 (N_32299,N_29645,N_29308);
nor U32300 (N_32300,N_27831,N_27635);
and U32301 (N_32301,N_29655,N_28940);
xnor U32302 (N_32302,N_27804,N_27656);
or U32303 (N_32303,N_28980,N_28601);
nor U32304 (N_32304,N_29660,N_28394);
xor U32305 (N_32305,N_28325,N_28823);
nand U32306 (N_32306,N_29744,N_28265);
nand U32307 (N_32307,N_29726,N_27814);
xor U32308 (N_32308,N_29433,N_29008);
nand U32309 (N_32309,N_28062,N_27722);
or U32310 (N_32310,N_27847,N_28837);
nor U32311 (N_32311,N_29884,N_28764);
or U32312 (N_32312,N_28332,N_29200);
xnor U32313 (N_32313,N_29725,N_28941);
nor U32314 (N_32314,N_29350,N_29949);
and U32315 (N_32315,N_29459,N_28891);
xor U32316 (N_32316,N_28699,N_27897);
and U32317 (N_32317,N_29410,N_29394);
and U32318 (N_32318,N_29053,N_29702);
and U32319 (N_32319,N_29802,N_27654);
xnor U32320 (N_32320,N_29769,N_27811);
xnor U32321 (N_32321,N_28926,N_27807);
xor U32322 (N_32322,N_29912,N_28134);
or U32323 (N_32323,N_29512,N_29582);
xnor U32324 (N_32324,N_28314,N_29124);
nor U32325 (N_32325,N_27950,N_28788);
nand U32326 (N_32326,N_27741,N_27716);
nor U32327 (N_32327,N_29501,N_29393);
nor U32328 (N_32328,N_29237,N_28842);
nor U32329 (N_32329,N_28106,N_28452);
nand U32330 (N_32330,N_27718,N_28319);
nor U32331 (N_32331,N_29789,N_28234);
xor U32332 (N_32332,N_27812,N_28382);
nand U32333 (N_32333,N_28337,N_29109);
and U32334 (N_32334,N_29599,N_28040);
xor U32335 (N_32335,N_28798,N_29321);
and U32336 (N_32336,N_29084,N_28286);
and U32337 (N_32337,N_29045,N_28487);
and U32338 (N_32338,N_29305,N_27915);
nor U32339 (N_32339,N_29879,N_28777);
and U32340 (N_32340,N_29147,N_29556);
or U32341 (N_32341,N_28018,N_29104);
xnor U32342 (N_32342,N_28190,N_28583);
and U32343 (N_32343,N_28497,N_28117);
nor U32344 (N_32344,N_29052,N_27984);
nor U32345 (N_32345,N_28347,N_28783);
nand U32346 (N_32346,N_28116,N_29069);
xnor U32347 (N_32347,N_29116,N_29123);
nor U32348 (N_32348,N_28399,N_28640);
xor U32349 (N_32349,N_28600,N_28175);
nor U32350 (N_32350,N_29265,N_29805);
or U32351 (N_32351,N_28131,N_28305);
nand U32352 (N_32352,N_28612,N_27635);
nor U32353 (N_32353,N_29985,N_29327);
xor U32354 (N_32354,N_29066,N_29612);
nand U32355 (N_32355,N_27939,N_29355);
xor U32356 (N_32356,N_29207,N_29442);
nand U32357 (N_32357,N_27591,N_27541);
nand U32358 (N_32358,N_27769,N_28408);
xnor U32359 (N_32359,N_29199,N_28923);
and U32360 (N_32360,N_27601,N_29402);
or U32361 (N_32361,N_28071,N_28558);
or U32362 (N_32362,N_28511,N_29393);
or U32363 (N_32363,N_27839,N_29181);
and U32364 (N_32364,N_28735,N_27784);
and U32365 (N_32365,N_27664,N_28835);
xnor U32366 (N_32366,N_27707,N_27919);
or U32367 (N_32367,N_29024,N_29607);
nand U32368 (N_32368,N_29682,N_28996);
and U32369 (N_32369,N_29666,N_29709);
nor U32370 (N_32370,N_28013,N_28309);
xor U32371 (N_32371,N_27961,N_29870);
nand U32372 (N_32372,N_29273,N_27639);
and U32373 (N_32373,N_28793,N_29963);
or U32374 (N_32374,N_28994,N_29293);
or U32375 (N_32375,N_27583,N_28839);
xor U32376 (N_32376,N_27786,N_29881);
nand U32377 (N_32377,N_29153,N_29294);
and U32378 (N_32378,N_29293,N_28590);
and U32379 (N_32379,N_28094,N_29557);
xnor U32380 (N_32380,N_29797,N_29889);
xor U32381 (N_32381,N_29183,N_28732);
nand U32382 (N_32382,N_29100,N_28685);
or U32383 (N_32383,N_27506,N_28534);
xnor U32384 (N_32384,N_28299,N_28217);
xnor U32385 (N_32385,N_28993,N_28780);
nand U32386 (N_32386,N_28816,N_27859);
or U32387 (N_32387,N_28783,N_28374);
and U32388 (N_32388,N_28079,N_29017);
and U32389 (N_32389,N_27993,N_28387);
nor U32390 (N_32390,N_28777,N_28140);
xor U32391 (N_32391,N_27867,N_29657);
nor U32392 (N_32392,N_29439,N_29506);
nor U32393 (N_32393,N_29126,N_27501);
and U32394 (N_32394,N_28952,N_27883);
or U32395 (N_32395,N_29453,N_29674);
nor U32396 (N_32396,N_28416,N_27913);
nand U32397 (N_32397,N_28192,N_27542);
xnor U32398 (N_32398,N_29902,N_29790);
nand U32399 (N_32399,N_28986,N_29353);
xor U32400 (N_32400,N_28182,N_29962);
xnor U32401 (N_32401,N_27862,N_29216);
nand U32402 (N_32402,N_28163,N_28732);
and U32403 (N_32403,N_29380,N_28300);
xor U32404 (N_32404,N_28846,N_29465);
and U32405 (N_32405,N_28341,N_27876);
nand U32406 (N_32406,N_29483,N_28461);
nor U32407 (N_32407,N_28801,N_28380);
nand U32408 (N_32408,N_27764,N_28575);
nand U32409 (N_32409,N_29500,N_28064);
and U32410 (N_32410,N_29822,N_27901);
and U32411 (N_32411,N_29939,N_28402);
nand U32412 (N_32412,N_28842,N_29618);
xor U32413 (N_32413,N_29425,N_27687);
nand U32414 (N_32414,N_27870,N_28524);
and U32415 (N_32415,N_27651,N_28146);
or U32416 (N_32416,N_27728,N_27838);
or U32417 (N_32417,N_29849,N_27565);
or U32418 (N_32418,N_28089,N_29294);
nand U32419 (N_32419,N_29793,N_29326);
nor U32420 (N_32420,N_28313,N_28270);
xnor U32421 (N_32421,N_27560,N_28142);
or U32422 (N_32422,N_27520,N_29601);
xor U32423 (N_32423,N_27680,N_29420);
and U32424 (N_32424,N_28719,N_28938);
nor U32425 (N_32425,N_28487,N_27551);
xnor U32426 (N_32426,N_29286,N_27900);
nand U32427 (N_32427,N_29264,N_29822);
nor U32428 (N_32428,N_28305,N_28983);
xnor U32429 (N_32429,N_29865,N_28934);
xnor U32430 (N_32430,N_29381,N_29130);
and U32431 (N_32431,N_29767,N_28953);
nor U32432 (N_32432,N_29754,N_27995);
and U32433 (N_32433,N_28294,N_27754);
nor U32434 (N_32434,N_29454,N_28345);
nand U32435 (N_32435,N_29407,N_28907);
xor U32436 (N_32436,N_29991,N_29786);
or U32437 (N_32437,N_28916,N_28353);
or U32438 (N_32438,N_28833,N_29009);
and U32439 (N_32439,N_28676,N_27708);
nand U32440 (N_32440,N_28697,N_29749);
nand U32441 (N_32441,N_29080,N_28546);
or U32442 (N_32442,N_29842,N_29759);
xor U32443 (N_32443,N_28124,N_27568);
xnor U32444 (N_32444,N_29872,N_29674);
nor U32445 (N_32445,N_29445,N_29887);
and U32446 (N_32446,N_27596,N_28672);
nor U32447 (N_32447,N_27848,N_29858);
nand U32448 (N_32448,N_27771,N_28702);
xor U32449 (N_32449,N_29007,N_29287);
or U32450 (N_32450,N_28475,N_27810);
xnor U32451 (N_32451,N_27767,N_29859);
xor U32452 (N_32452,N_29986,N_29676);
nand U32453 (N_32453,N_29414,N_27979);
nor U32454 (N_32454,N_27751,N_28650);
and U32455 (N_32455,N_29536,N_27995);
nor U32456 (N_32456,N_28510,N_29789);
xor U32457 (N_32457,N_29891,N_29687);
nor U32458 (N_32458,N_28988,N_28604);
and U32459 (N_32459,N_29286,N_29104);
nor U32460 (N_32460,N_29819,N_27538);
xnor U32461 (N_32461,N_28278,N_29250);
nor U32462 (N_32462,N_28832,N_27817);
xor U32463 (N_32463,N_28531,N_28416);
xnor U32464 (N_32464,N_28372,N_27887);
and U32465 (N_32465,N_28788,N_28575);
and U32466 (N_32466,N_29175,N_28842);
nor U32467 (N_32467,N_29168,N_29681);
xor U32468 (N_32468,N_27600,N_29252);
nand U32469 (N_32469,N_29072,N_29473);
xnor U32470 (N_32470,N_28331,N_28579);
or U32471 (N_32471,N_29339,N_28534);
or U32472 (N_32472,N_27925,N_28854);
nand U32473 (N_32473,N_28505,N_29351);
or U32474 (N_32474,N_27819,N_28307);
nand U32475 (N_32475,N_27697,N_27853);
nor U32476 (N_32476,N_29921,N_27529);
nand U32477 (N_32477,N_29909,N_29578);
and U32478 (N_32478,N_28631,N_28933);
nor U32479 (N_32479,N_27813,N_28996);
or U32480 (N_32480,N_27756,N_29400);
nor U32481 (N_32481,N_29752,N_28831);
or U32482 (N_32482,N_27919,N_27837);
and U32483 (N_32483,N_27940,N_29934);
and U32484 (N_32484,N_27778,N_28403);
or U32485 (N_32485,N_28979,N_28503);
nor U32486 (N_32486,N_28358,N_28240);
and U32487 (N_32487,N_28946,N_29365);
or U32488 (N_32488,N_28077,N_29383);
nand U32489 (N_32489,N_28287,N_28590);
nand U32490 (N_32490,N_27776,N_28292);
xor U32491 (N_32491,N_28520,N_27829);
and U32492 (N_32492,N_28778,N_28207);
and U32493 (N_32493,N_28022,N_28145);
nor U32494 (N_32494,N_29552,N_28501);
xor U32495 (N_32495,N_29677,N_28730);
and U32496 (N_32496,N_29697,N_29098);
nor U32497 (N_32497,N_29227,N_28156);
or U32498 (N_32498,N_28563,N_28148);
or U32499 (N_32499,N_29508,N_28605);
xnor U32500 (N_32500,N_31193,N_30570);
and U32501 (N_32501,N_30696,N_32202);
nor U32502 (N_32502,N_30568,N_31178);
or U32503 (N_32503,N_31712,N_32006);
or U32504 (N_32504,N_30463,N_31394);
and U32505 (N_32505,N_30864,N_30227);
nand U32506 (N_32506,N_31256,N_30824);
xor U32507 (N_32507,N_30911,N_31058);
or U32508 (N_32508,N_30338,N_31095);
nor U32509 (N_32509,N_30341,N_30523);
or U32510 (N_32510,N_31552,N_30237);
nor U32511 (N_32511,N_30575,N_32444);
or U32512 (N_32512,N_31540,N_32253);
or U32513 (N_32513,N_31233,N_31406);
nor U32514 (N_32514,N_30711,N_31044);
and U32515 (N_32515,N_31805,N_30176);
or U32516 (N_32516,N_31150,N_32486);
or U32517 (N_32517,N_31449,N_30037);
xnor U32518 (N_32518,N_31462,N_32381);
xnor U32519 (N_32519,N_31688,N_32452);
nand U32520 (N_32520,N_30404,N_30287);
or U32521 (N_32521,N_30811,N_30397);
xor U32522 (N_32522,N_31781,N_31112);
nand U32523 (N_32523,N_30332,N_32179);
xnor U32524 (N_32524,N_31590,N_31851);
and U32525 (N_32525,N_32364,N_30647);
and U32526 (N_32526,N_30008,N_31436);
xnor U32527 (N_32527,N_31732,N_30145);
nor U32528 (N_32528,N_32127,N_31988);
xnor U32529 (N_32529,N_30874,N_31513);
nand U32530 (N_32530,N_30866,N_31853);
or U32531 (N_32531,N_30152,N_32245);
and U32532 (N_32532,N_30887,N_30094);
or U32533 (N_32533,N_31611,N_30858);
nor U32534 (N_32534,N_31629,N_32476);
and U32535 (N_32535,N_31765,N_32488);
nand U32536 (N_32536,N_31990,N_31183);
or U32537 (N_32537,N_30444,N_30848);
nand U32538 (N_32538,N_31268,N_31745);
nand U32539 (N_32539,N_30067,N_30788);
nor U32540 (N_32540,N_30372,N_31922);
nand U32541 (N_32541,N_31530,N_30052);
and U32542 (N_32542,N_30106,N_30307);
or U32543 (N_32543,N_30311,N_31751);
and U32544 (N_32544,N_30506,N_31868);
and U32545 (N_32545,N_31921,N_30770);
or U32546 (N_32546,N_30177,N_32300);
and U32547 (N_32547,N_32081,N_30620);
xor U32548 (N_32548,N_31184,N_31027);
nand U32549 (N_32549,N_31148,N_31844);
and U32550 (N_32550,N_30481,N_30772);
nor U32551 (N_32551,N_31848,N_32330);
or U32552 (N_32552,N_30465,N_31188);
nor U32553 (N_32553,N_30740,N_30718);
xor U32554 (N_32554,N_31738,N_31906);
nand U32555 (N_32555,N_30756,N_30112);
nand U32556 (N_32556,N_31799,N_32413);
nor U32557 (N_32557,N_31963,N_31594);
nor U32558 (N_32558,N_31203,N_32361);
nand U32559 (N_32559,N_31077,N_30579);
or U32560 (N_32560,N_32449,N_30862);
or U32561 (N_32561,N_30605,N_31155);
or U32562 (N_32562,N_30498,N_31826);
or U32563 (N_32563,N_31156,N_31979);
xor U32564 (N_32564,N_31453,N_31473);
and U32565 (N_32565,N_30651,N_31201);
nor U32566 (N_32566,N_32148,N_30019);
xor U32567 (N_32567,N_31776,N_31763);
or U32568 (N_32568,N_30365,N_31429);
nor U32569 (N_32569,N_31424,N_31866);
nand U32570 (N_32570,N_31820,N_30680);
xnor U32571 (N_32571,N_30108,N_32184);
nand U32572 (N_32572,N_32320,N_30169);
or U32573 (N_32573,N_31172,N_30441);
or U32574 (N_32574,N_31981,N_32029);
nand U32575 (N_32575,N_30072,N_30088);
and U32576 (N_32576,N_30946,N_30692);
and U32577 (N_32577,N_31091,N_31630);
nor U32578 (N_32578,N_32333,N_30985);
and U32579 (N_32579,N_30412,N_30903);
xor U32580 (N_32580,N_30741,N_32086);
nor U32581 (N_32581,N_30980,N_31067);
nor U32582 (N_32582,N_32387,N_32058);
and U32583 (N_32583,N_32312,N_32067);
xor U32584 (N_32584,N_30725,N_30458);
xor U32585 (N_32585,N_31499,N_32464);
or U32586 (N_32586,N_31541,N_30846);
or U32587 (N_32587,N_31220,N_30077);
xnor U32588 (N_32588,N_30834,N_31497);
xor U32589 (N_32589,N_30793,N_30295);
xor U32590 (N_32590,N_30906,N_31551);
nor U32591 (N_32591,N_32323,N_31599);
nand U32592 (N_32592,N_32338,N_30863);
nor U32593 (N_32593,N_30713,N_31415);
nor U32594 (N_32594,N_31525,N_31152);
xnor U32595 (N_32595,N_30670,N_30061);
nand U32596 (N_32596,N_31408,N_30432);
nand U32597 (N_32597,N_30102,N_31287);
nor U32598 (N_32598,N_32351,N_30005);
or U32599 (N_32599,N_31364,N_30800);
nand U32600 (N_32600,N_31089,N_30784);
or U32601 (N_32601,N_30403,N_31855);
nor U32602 (N_32602,N_30258,N_31359);
and U32603 (N_32603,N_30248,N_31617);
nor U32604 (N_32604,N_31674,N_30484);
and U32605 (N_32605,N_32360,N_30136);
and U32606 (N_32606,N_30244,N_31167);
nand U32607 (N_32607,N_30831,N_31157);
xor U32608 (N_32608,N_30766,N_32378);
or U32609 (N_32609,N_30998,N_30600);
xnor U32610 (N_32610,N_31775,N_30556);
xnor U32611 (N_32611,N_31725,N_30423);
nor U32612 (N_32612,N_32078,N_31812);
nand U32613 (N_32613,N_31622,N_30908);
or U32614 (N_32614,N_31883,N_31686);
xnor U32615 (N_32615,N_30485,N_32170);
xor U32616 (N_32616,N_30271,N_31894);
xor U32617 (N_32617,N_31191,N_32064);
nor U32618 (N_32618,N_30918,N_32383);
or U32619 (N_32619,N_31567,N_30167);
nand U32620 (N_32620,N_30893,N_30532);
or U32621 (N_32621,N_32372,N_30511);
nor U32622 (N_32622,N_30882,N_30489);
or U32623 (N_32623,N_32395,N_30666);
nand U32624 (N_32624,N_31949,N_31915);
nor U32625 (N_32625,N_31495,N_32454);
and U32626 (N_32626,N_30209,N_32283);
and U32627 (N_32627,N_32374,N_31888);
and U32628 (N_32628,N_31041,N_31318);
and U32629 (N_32629,N_31299,N_30901);
nor U32630 (N_32630,N_30815,N_32479);
or U32631 (N_32631,N_30122,N_30510);
nor U32632 (N_32632,N_30440,N_32328);
xor U32633 (N_32633,N_31115,N_31940);
or U32634 (N_32634,N_30038,N_31623);
nand U32635 (N_32635,N_31864,N_30936);
xnor U32636 (N_32636,N_30656,N_31478);
nor U32637 (N_32637,N_30141,N_30071);
nor U32638 (N_32638,N_30306,N_32377);
xor U32639 (N_32639,N_31312,N_31746);
and U32640 (N_32640,N_31218,N_31856);
or U32641 (N_32641,N_30431,N_30852);
or U32642 (N_32642,N_31321,N_32324);
nand U32643 (N_32643,N_31254,N_31279);
nand U32644 (N_32644,N_31263,N_31253);
and U32645 (N_32645,N_32132,N_31802);
xnor U32646 (N_32646,N_31367,N_32494);
nand U32647 (N_32647,N_30009,N_31224);
or U32648 (N_32648,N_31953,N_31438);
xor U32649 (N_32649,N_30947,N_30616);
and U32650 (N_32650,N_32062,N_30551);
nand U32651 (N_32651,N_32362,N_32302);
nor U32652 (N_32652,N_30368,N_30667);
nor U32653 (N_32653,N_32366,N_31422);
nand U32654 (N_32654,N_32273,N_32082);
xnor U32655 (N_32655,N_30123,N_32472);
and U32656 (N_32656,N_31837,N_30631);
nor U32657 (N_32657,N_32435,N_30508);
or U32658 (N_32658,N_32329,N_31040);
or U32659 (N_32659,N_30538,N_30157);
xor U32660 (N_32660,N_31399,N_31428);
xnor U32661 (N_32661,N_31669,N_31015);
nor U32662 (N_32662,N_31212,N_31801);
and U32663 (N_32663,N_32389,N_31616);
xor U32664 (N_32664,N_31199,N_30950);
nor U32665 (N_32665,N_32487,N_31941);
or U32666 (N_32666,N_32332,N_31356);
xor U32667 (N_32667,N_32033,N_31282);
nor U32668 (N_32668,N_30087,N_31580);
nor U32669 (N_32669,N_30388,N_31595);
and U32670 (N_32670,N_31681,N_31929);
or U32671 (N_32671,N_32077,N_31579);
or U32672 (N_32672,N_31235,N_31443);
nor U32673 (N_32673,N_31790,N_30888);
xnor U32674 (N_32674,N_32246,N_30607);
nand U32675 (N_32675,N_30709,N_31717);
nand U32676 (N_32676,N_30066,N_32255);
nand U32677 (N_32677,N_30348,N_31510);
or U32678 (N_32678,N_31392,N_30154);
or U32679 (N_32679,N_30319,N_31146);
or U32680 (N_32680,N_31186,N_30124);
nor U32681 (N_32681,N_31144,N_32261);
and U32682 (N_32682,N_32186,N_30924);
nand U32683 (N_32683,N_32438,N_30585);
and U32684 (N_32684,N_31306,N_30612);
and U32685 (N_32685,N_31578,N_30878);
nand U32686 (N_32686,N_31369,N_31419);
xor U32687 (N_32687,N_32160,N_30199);
nor U32688 (N_32688,N_30584,N_30004);
nor U32689 (N_32689,N_30531,N_31161);
nor U32690 (N_32690,N_32201,N_30305);
or U32691 (N_32691,N_31691,N_30398);
xnor U32692 (N_32692,N_31154,N_31999);
nand U32693 (N_32693,N_30957,N_31412);
and U32694 (N_32694,N_32157,N_32133);
nor U32695 (N_32695,N_31085,N_30638);
xor U32696 (N_32696,N_30405,N_32140);
and U32697 (N_32697,N_30650,N_32365);
and U32698 (N_32698,N_30483,N_32489);
xnor U32699 (N_32699,N_32232,N_32341);
nor U32700 (N_32700,N_31606,N_32244);
and U32701 (N_32701,N_31023,N_31522);
or U32702 (N_32702,N_31272,N_30640);
nor U32703 (N_32703,N_30128,N_31749);
xnor U32704 (N_32704,N_32084,N_30768);
or U32705 (N_32705,N_31679,N_30466);
nor U32706 (N_32706,N_30146,N_30502);
nor U32707 (N_32707,N_30062,N_32423);
nand U32708 (N_32708,N_32288,N_32197);
nand U32709 (N_32709,N_31469,N_31944);
and U32710 (N_32710,N_31434,N_31409);
and U32711 (N_32711,N_30972,N_30528);
nor U32712 (N_32712,N_31936,N_32420);
xor U32713 (N_32713,N_31343,N_30479);
xnor U32714 (N_32714,N_32400,N_31713);
nand U32715 (N_32715,N_30421,N_30748);
nor U32716 (N_32716,N_32214,N_30525);
and U32717 (N_32717,N_30581,N_31302);
nor U32718 (N_32718,N_31685,N_31333);
or U32719 (N_32719,N_31440,N_31954);
nand U32720 (N_32720,N_30468,N_31741);
nor U32721 (N_32721,N_31116,N_30917);
nor U32722 (N_32722,N_31330,N_31692);
nor U32723 (N_32723,N_31643,N_32355);
nand U32724 (N_32724,N_32146,N_31229);
or U32725 (N_32725,N_30153,N_31536);
xor U32726 (N_32726,N_32308,N_32385);
or U32727 (N_32727,N_31391,N_31886);
nor U32728 (N_32728,N_31106,N_30657);
nor U32729 (N_32729,N_32155,N_30053);
or U32730 (N_32730,N_31834,N_31896);
or U32731 (N_32731,N_30833,N_30030);
nor U32732 (N_32732,N_31935,N_31633);
or U32733 (N_32733,N_31709,N_30691);
or U32734 (N_32734,N_31774,N_30084);
nor U32735 (N_32735,N_32168,N_30313);
nor U32736 (N_32736,N_30642,N_31880);
xor U32737 (N_32737,N_32159,N_31083);
and U32738 (N_32738,N_31032,N_31511);
nand U32739 (N_32739,N_30475,N_30595);
xor U32740 (N_32740,N_32022,N_31123);
nand U32741 (N_32741,N_31304,N_31624);
and U32742 (N_32742,N_32139,N_31948);
and U32743 (N_32743,N_30907,N_32128);
nor U32744 (N_32744,N_31170,N_30242);
nor U32745 (N_32745,N_30637,N_30817);
and U32746 (N_32746,N_32290,N_31099);
xor U32747 (N_32747,N_31727,N_30586);
xnor U32748 (N_32748,N_32490,N_31753);
or U32749 (N_32749,N_32286,N_32258);
and U32750 (N_32750,N_30762,N_30745);
xnor U32751 (N_32751,N_30672,N_30433);
nand U32752 (N_32752,N_31262,N_31223);
nand U32753 (N_32753,N_31494,N_30239);
or U32754 (N_32754,N_30247,N_31997);
nand U32755 (N_32755,N_31822,N_32226);
or U32756 (N_32756,N_31601,N_31528);
nand U32757 (N_32757,N_32450,N_30422);
nor U32758 (N_32758,N_31597,N_30899);
and U32759 (N_32759,N_32335,N_30916);
nor U32760 (N_32760,N_31145,N_32008);
or U32761 (N_32761,N_30288,N_30493);
nand U32762 (N_32762,N_30447,N_31159);
xor U32763 (N_32763,N_30386,N_30003);
nor U32764 (N_32764,N_30794,N_32259);
nor U32765 (N_32765,N_32265,N_30265);
nand U32766 (N_32766,N_31800,N_31082);
nor U32767 (N_32767,N_31577,N_31336);
nor U32768 (N_32768,N_31003,N_30114);
and U32769 (N_32769,N_31714,N_31750);
or U32770 (N_32770,N_32072,N_30455);
and U32771 (N_32771,N_30266,N_31240);
nor U32772 (N_32772,N_30369,N_32178);
or U32773 (N_32773,N_30792,N_30540);
or U32774 (N_32774,N_32024,N_30370);
or U32775 (N_32775,N_31852,N_31195);
nor U32776 (N_32776,N_31779,N_30801);
nor U32777 (N_32777,N_31034,N_31784);
nor U32778 (N_32778,N_30320,N_30276);
nand U32779 (N_32779,N_31381,N_30393);
xnor U32780 (N_32780,N_30041,N_31715);
and U32781 (N_32781,N_31484,N_30842);
nor U32782 (N_32782,N_30803,N_30739);
nand U32783 (N_32783,N_31919,N_31442);
or U32784 (N_32784,N_30501,N_32434);
xor U32785 (N_32785,N_32268,N_30614);
xor U32786 (N_32786,N_30996,N_30827);
xnor U32787 (N_32787,N_31134,N_30492);
and U32788 (N_32788,N_31891,N_32037);
nor U32789 (N_32789,N_30715,N_32020);
or U32790 (N_32790,N_30719,N_31995);
nor U32791 (N_32791,N_30353,N_31829);
xnor U32792 (N_32792,N_31242,N_31390);
nand U32793 (N_32793,N_30563,N_30336);
xor U32794 (N_32794,N_30749,N_30582);
and U32795 (N_32795,N_30042,N_31723);
nand U32796 (N_32796,N_30580,N_32195);
nand U32797 (N_32797,N_30300,N_30340);
nor U32798 (N_32798,N_30686,N_30951);
nand U32799 (N_32799,N_31393,N_32189);
or U32800 (N_32800,N_31311,N_31383);
nor U32801 (N_32801,N_31592,N_32291);
or U32802 (N_32802,N_32073,N_31678);
nand U32803 (N_32803,N_30158,N_30663);
or U32804 (N_32804,N_31734,N_32461);
and U32805 (N_32805,N_30357,N_31724);
xnor U32806 (N_32806,N_31185,N_32236);
nand U32807 (N_32807,N_31008,N_30814);
nor U32808 (N_32808,N_30659,N_31052);
or U32809 (N_32809,N_30829,N_30889);
nand U32810 (N_32810,N_30012,N_31210);
nor U32811 (N_32811,N_32309,N_32122);
and U32812 (N_32812,N_30210,N_31910);
or U32813 (N_32813,N_31503,N_32388);
and U32814 (N_32814,N_30362,N_31363);
and U32815 (N_32815,N_31895,N_30944);
xor U32816 (N_32816,N_30389,N_31360);
nand U32817 (N_32817,N_31490,N_31942);
and U32818 (N_32818,N_30683,N_32028);
xnor U32819 (N_32819,N_30188,N_32359);
nor U32820 (N_32820,N_30738,N_31729);
and U32821 (N_32821,N_32102,N_32121);
xor U32822 (N_32822,N_30920,N_32013);
nor U32823 (N_32823,N_30931,N_32241);
xnor U32824 (N_32824,N_31987,N_31487);
nor U32825 (N_32825,N_30127,N_32433);
or U32826 (N_32826,N_32293,N_31926);
xor U32827 (N_32827,N_30354,N_30063);
nor U32828 (N_32828,N_31591,N_30168);
and U32829 (N_32829,N_30660,N_31500);
and U32830 (N_32830,N_30940,N_30180);
or U32831 (N_32831,N_30818,N_31584);
or U32832 (N_32832,N_30669,N_32198);
nor U32833 (N_32833,N_30661,N_31973);
nand U32834 (N_32834,N_31897,N_32042);
xnor U32835 (N_32835,N_32411,N_30997);
nand U32836 (N_32836,N_32275,N_30625);
xnor U32837 (N_32837,N_30658,N_30791);
xor U32838 (N_32838,N_32453,N_31350);
or U32839 (N_32839,N_30594,N_32223);
nor U32840 (N_32840,N_31632,N_32422);
xor U32841 (N_32841,N_30643,N_30844);
and U32842 (N_32842,N_30943,N_32369);
nor U32843 (N_32843,N_31783,N_30927);
nand U32844 (N_32844,N_30407,N_32326);
or U32845 (N_32845,N_32262,N_30499);
nand U32846 (N_32846,N_31445,N_30111);
and U32847 (N_32847,N_31761,N_30759);
xor U32848 (N_32848,N_30790,N_30641);
xnor U32849 (N_32849,N_30774,N_30549);
or U32850 (N_32850,N_31328,N_30017);
xor U32851 (N_32851,N_31276,N_30095);
nand U32852 (N_32852,N_30876,N_31731);
xor U32853 (N_32853,N_31474,N_32243);
and U32854 (N_32854,N_31230,N_31559);
and U32855 (N_32855,N_30026,N_31792);
nand U32856 (N_32856,N_31056,N_32440);
or U32857 (N_32857,N_30476,N_31832);
xnor U32858 (N_32858,N_30304,N_30161);
nand U32859 (N_32859,N_32458,N_31012);
nand U32860 (N_32860,N_31575,N_32390);
xnor U32861 (N_32861,N_31573,N_30080);
xor U32862 (N_32862,N_30135,N_30032);
nor U32863 (N_32863,N_32207,N_32027);
xor U32864 (N_32864,N_31017,N_31952);
nor U32865 (N_32865,N_32206,N_31947);
xnor U32866 (N_32866,N_31726,N_30820);
nand U32867 (N_32867,N_30934,N_30333);
or U32868 (N_32868,N_30546,N_30207);
nor U32869 (N_32869,N_30065,N_32023);
xor U32870 (N_32870,N_32141,N_30622);
or U32871 (N_32871,N_31102,N_30232);
xnor U32872 (N_32872,N_31411,N_30376);
xnor U32873 (N_32873,N_31859,N_32004);
nand U32874 (N_32874,N_32240,N_30254);
nand U32875 (N_32875,N_30314,N_30092);
and U32876 (N_32876,N_31329,N_31209);
nand U32877 (N_32877,N_32439,N_31720);
or U32878 (N_32878,N_32176,N_30777);
or U32879 (N_32879,N_30821,N_30277);
nor U32880 (N_32880,N_31650,N_31704);
nor U32881 (N_32881,N_31554,N_31379);
nand U32882 (N_32882,N_32250,N_32498);
nand U32883 (N_32883,N_30263,N_31342);
nand U32884 (N_32884,N_30560,N_30543);
or U32885 (N_32885,N_31872,N_30832);
or U32886 (N_32886,N_32052,N_32147);
or U32887 (N_32887,N_31006,N_31817);
nor U32888 (N_32888,N_31718,N_30513);
nand U32889 (N_32889,N_32040,N_31526);
nand U32890 (N_32890,N_30262,N_32301);
nand U32891 (N_32891,N_31250,N_31389);
or U32892 (N_32892,N_31966,N_30608);
and U32893 (N_32893,N_32091,N_32169);
xor U32894 (N_32894,N_30202,N_32281);
nand U32895 (N_32895,N_31400,N_30259);
nand U32896 (N_32896,N_32032,N_31609);
nor U32897 (N_32897,N_30225,N_31004);
or U32898 (N_32898,N_30805,N_32491);
or U32899 (N_32899,N_32235,N_30861);
or U32900 (N_32900,N_30325,N_30869);
or U32901 (N_32901,N_31671,N_30173);
and U32902 (N_32902,N_30897,N_31217);
and U32903 (N_32903,N_31730,N_30720);
xor U32904 (N_32904,N_31496,N_31539);
or U32905 (N_32905,N_31892,N_32282);
nor U32906 (N_32906,N_31327,N_30408);
xnor U32907 (N_32907,N_31171,N_31523);
or U32908 (N_32908,N_31347,N_31192);
xor U32909 (N_32909,N_31702,N_30016);
nor U32910 (N_32910,N_30545,N_31989);
xnor U32911 (N_32911,N_32099,N_31770);
nor U32912 (N_32912,N_30597,N_32321);
nor U32913 (N_32913,N_30281,N_32229);
nand U32914 (N_32914,N_30134,N_31768);
and U32915 (N_32915,N_31060,N_32145);
and U32916 (N_32916,N_31326,N_30836);
and U32917 (N_32917,N_30414,N_31149);
nand U32918 (N_32918,N_30138,N_30434);
and U32919 (N_32919,N_30609,N_31252);
nor U32920 (N_32920,N_30646,N_31021);
nand U32921 (N_32921,N_32230,N_30081);
nor U32922 (N_32922,N_30881,N_31543);
or U32923 (N_32923,N_32209,N_32167);
nand U32924 (N_32924,N_30875,N_30070);
or U32925 (N_32925,N_31065,N_32474);
and U32926 (N_32926,N_31736,N_31387);
or U32927 (N_32927,N_31324,N_31045);
xnor U32928 (N_32928,N_30912,N_31945);
and U32929 (N_32929,N_31520,N_31244);
nand U32930 (N_32930,N_30257,N_31804);
xnor U32931 (N_32931,N_30895,N_31396);
nand U32932 (N_32932,N_32292,N_32484);
nand U32933 (N_32933,N_32213,N_31862);
nand U32934 (N_32934,N_30192,N_32459);
xor U32935 (N_32935,N_30537,N_31794);
xnor U32936 (N_32936,N_31431,N_30160);
xnor U32937 (N_32937,N_30877,N_31423);
and U32938 (N_32938,N_30558,N_32113);
nor U32939 (N_32939,N_30260,N_30044);
nor U32940 (N_32940,N_30904,N_31069);
nor U32941 (N_32941,N_30671,N_32313);
nor U32942 (N_32942,N_31547,N_30025);
nand U32943 (N_32943,N_31457,N_30054);
and U32944 (N_32944,N_31833,N_30522);
xnor U32945 (N_32945,N_31904,N_32192);
xor U32946 (N_32946,N_31984,N_30747);
or U32947 (N_32947,N_30505,N_31808);
and U32948 (N_32948,N_32218,N_30089);
xnor U32949 (N_32949,N_31177,N_32347);
or U32950 (N_32950,N_31103,N_30964);
xor U32951 (N_32951,N_30515,N_30883);
and U32952 (N_32952,N_31917,N_30182);
nand U32953 (N_32953,N_30022,N_32063);
and U32954 (N_32954,N_32203,N_30981);
nor U32955 (N_32955,N_32120,N_30456);
xor U32956 (N_32956,N_30668,N_31035);
nand U32957 (N_32957,N_30027,N_31777);
and U32958 (N_32958,N_32083,N_30486);
xor U32959 (N_32959,N_31977,N_32228);
or U32960 (N_32960,N_30624,N_31197);
or U32961 (N_32961,N_32447,N_31168);
nand U32962 (N_32962,N_31066,N_30955);
nor U32963 (N_32963,N_30885,N_32087);
xnor U32964 (N_32964,N_31135,N_31690);
and U32965 (N_32965,N_32256,N_31682);
or U32966 (N_32966,N_31114,N_31030);
nor U32967 (N_32967,N_30564,N_31076);
xor U32968 (N_32968,N_30710,N_32357);
xor U32969 (N_32969,N_30589,N_31410);
nand U32970 (N_32970,N_30378,N_32429);
nor U32971 (N_32971,N_30097,N_31301);
or U32972 (N_32972,N_31908,N_30665);
or U32973 (N_32973,N_32248,N_31345);
nand U32974 (N_32974,N_30184,N_30343);
or U32975 (N_32975,N_31695,N_30855);
or U32976 (N_32976,N_31126,N_30807);
xor U32977 (N_32977,N_32493,N_32456);
xor U32978 (N_32978,N_31010,N_30409);
xor U32979 (N_32979,N_30377,N_30541);
and U32980 (N_32980,N_31960,N_30406);
xnor U32981 (N_32981,N_31346,N_31213);
xor U32982 (N_32982,N_32125,N_30473);
nand U32983 (N_32983,N_32068,N_30935);
or U32984 (N_32984,N_30808,N_31059);
xor U32985 (N_32985,N_32278,N_31827);
or U32986 (N_32986,N_30131,N_30384);
nor U32987 (N_32987,N_31286,N_31788);
or U32988 (N_32988,N_32174,N_30282);
or U32989 (N_32989,N_30096,N_30023);
nor U32990 (N_32990,N_31874,N_31502);
xnor U32991 (N_32991,N_31506,N_30561);
and U32992 (N_32992,N_32462,N_30076);
or U32993 (N_32993,N_31053,N_30334);
xnor U32994 (N_32994,N_32003,N_30171);
and U32995 (N_32995,N_30395,N_32049);
and U32996 (N_32996,N_31444,N_30769);
nor U32997 (N_32997,N_32346,N_31641);
and U32998 (N_32998,N_31703,N_32473);
nand U32999 (N_32999,N_30373,N_30949);
xor U33000 (N_33000,N_30879,N_30069);
nor U33001 (N_33001,N_31850,N_32134);
xor U33002 (N_33002,N_30648,N_32172);
or U33003 (N_33003,N_31460,N_31375);
xnor U33004 (N_33004,N_32109,N_31081);
nand U33005 (N_33005,N_31631,N_32354);
or U33006 (N_33006,N_30559,N_32118);
nand U33007 (N_33007,N_32270,N_30816);
xnor U33008 (N_33008,N_30318,N_30714);
and U33009 (N_33009,N_31672,N_32343);
nor U33010 (N_33010,N_30841,N_31418);
xor U33011 (N_33011,N_31867,N_32151);
nand U33012 (N_33012,N_31176,N_30635);
nor U33013 (N_33013,N_31884,N_31358);
nand U33014 (N_33014,N_32191,N_30236);
and U33015 (N_33015,N_31839,N_31181);
nand U33016 (N_33016,N_30825,N_31627);
nor U33017 (N_33017,N_30707,N_30965);
and U33018 (N_33018,N_31138,N_30352);
nand U33019 (N_33019,N_30402,N_31659);
and U33020 (N_33020,N_30929,N_31507);
nor U33021 (N_33021,N_31493,N_30233);
xnor U33022 (N_33022,N_31907,N_30891);
and U33023 (N_33023,N_32051,N_32363);
nor U33024 (N_33024,N_32257,N_32043);
nand U33025 (N_33025,N_32430,N_32272);
or U33026 (N_33026,N_31923,N_31297);
xor U33027 (N_33027,N_30487,N_32123);
or U33028 (N_33028,N_30645,N_31937);
and U33029 (N_33029,N_30555,N_30630);
or U33030 (N_33030,N_30235,N_31823);
nor U33031 (N_33031,N_30420,N_30284);
and U33032 (N_33032,N_31124,N_31401);
and U33033 (N_33033,N_31600,N_30988);
and U33034 (N_33034,N_30048,N_31214);
xnor U33035 (N_33035,N_31437,N_32010);
nor U33036 (N_33036,N_30569,N_31615);
and U33037 (N_33037,N_31227,N_31673);
nand U33038 (N_33038,N_32164,N_31310);
nand U33039 (N_33039,N_30435,N_30349);
nand U33040 (N_33040,N_30982,N_30383);
nand U33041 (N_33041,N_31563,N_30215);
nor U33042 (N_33042,N_31382,N_30494);
nor U33043 (N_33043,N_31221,N_31051);
nor U33044 (N_33044,N_30787,N_31613);
nand U33045 (N_33045,N_32352,N_30598);
nor U33046 (N_33046,N_30928,N_31569);
or U33047 (N_33047,N_30746,N_31470);
or U33048 (N_33048,N_32220,N_32342);
nor U33049 (N_33049,N_30149,N_31639);
nor U33050 (N_33050,N_30228,N_32138);
or U33051 (N_33051,N_30413,N_30117);
nor U33052 (N_33052,N_30221,N_32093);
and U33053 (N_33053,N_30722,N_31468);
nand U33054 (N_33054,N_31555,N_31560);
and U33055 (N_33055,N_30046,N_30159);
nor U33056 (N_33056,N_30850,N_30871);
nor U33057 (N_33057,N_31648,N_31258);
or U33058 (N_33058,N_31911,N_31598);
or U33059 (N_33059,N_30410,N_30457);
nand U33060 (N_33060,N_30922,N_30033);
nand U33061 (N_33061,N_30542,N_32090);
or U33062 (N_33062,N_30178,N_31341);
xnor U33063 (N_33063,N_30391,N_30778);
nand U33064 (N_33064,N_30557,N_30051);
nor U33065 (N_33065,N_30632,N_31972);
or U33066 (N_33066,N_31634,N_30674);
xor U33067 (N_33067,N_30971,N_31386);
xnor U33068 (N_33068,N_30098,N_30302);
nor U33069 (N_33069,N_31467,N_32469);
nand U33070 (N_33070,N_30035,N_32380);
xor U33071 (N_33071,N_31975,N_32391);
xor U33072 (N_33072,N_31780,N_32451);
or U33073 (N_33073,N_31247,N_30448);
and U33074 (N_33074,N_30723,N_31939);
nor U33075 (N_33075,N_31090,N_30984);
nand U33076 (N_33076,N_31706,N_32358);
nor U33077 (N_33077,N_31038,N_31372);
and U33078 (N_33078,N_31614,N_32216);
xor U33079 (N_33079,N_30703,N_32368);
nand U33080 (N_33080,N_32016,N_31019);
nor U33081 (N_33081,N_32421,N_30367);
and U33082 (N_33082,N_32379,N_30454);
nand U33083 (N_33083,N_31477,N_32219);
nor U33084 (N_33084,N_30593,N_32314);
or U33085 (N_33085,N_30133,N_31657);
nor U33086 (N_33086,N_31446,N_31707);
nor U33087 (N_33087,N_30308,N_31086);
nand U33088 (N_33088,N_32470,N_31315);
nor U33089 (N_33089,N_32480,N_31451);
and U33090 (N_33090,N_30424,N_30926);
nor U33091 (N_33091,N_32317,N_30382);
nor U33092 (N_33092,N_31970,N_31441);
xnor U33093 (N_33093,N_30213,N_30429);
nor U33094 (N_33094,N_32419,N_30512);
nand U33095 (N_33095,N_30195,N_32348);
xnor U33096 (N_33096,N_32396,N_32339);
xor U33097 (N_33097,N_30798,N_30385);
nand U33098 (N_33098,N_30342,N_31142);
xnor U33099 (N_33099,N_30544,N_30056);
nand U33100 (N_33100,N_30865,N_31546);
nor U33101 (N_33101,N_30143,N_30450);
nor U33102 (N_33102,N_32011,N_31986);
xnor U33103 (N_33103,N_32034,N_30702);
xor U33104 (N_33104,N_31307,N_31900);
and U33105 (N_33105,N_31913,N_31666);
and U33106 (N_33106,N_30074,N_32080);
nor U33107 (N_33107,N_30064,N_32035);
and U33108 (N_33108,N_32089,N_30990);
xor U33109 (N_33109,N_31976,N_30572);
nand U33110 (N_33110,N_30400,N_31593);
xnor U33111 (N_33111,N_32153,N_30203);
xnor U33112 (N_33112,N_31479,N_31132);
xnor U33113 (N_33113,N_32106,N_31352);
nand U33114 (N_33114,N_30101,N_30268);
xnor U33115 (N_33115,N_30329,N_31325);
nor U33116 (N_33116,N_30480,N_32427);
nor U33117 (N_33117,N_31959,N_31687);
xor U33118 (N_33118,N_30654,N_31196);
xor U33119 (N_33119,N_30204,N_31334);
nor U33120 (N_33120,N_31699,N_31049);
nor U33121 (N_33121,N_31028,N_31385);
nand U33122 (N_33122,N_30283,N_30488);
and U33123 (N_33123,N_30442,N_30509);
nand U33124 (N_33124,N_30913,N_30993);
nor U33125 (N_33125,N_30839,N_31384);
and U33126 (N_33126,N_30142,N_30419);
xor U33127 (N_33127,N_30571,N_31332);
and U33128 (N_33128,N_30565,N_31162);
xor U33129 (N_33129,N_31863,N_32416);
nand U33130 (N_33130,N_31280,N_32047);
or U33131 (N_33131,N_32404,N_32175);
nand U33132 (N_33132,N_32116,N_30472);
and U33133 (N_33133,N_31791,N_31043);
nand U33134 (N_33134,N_32224,N_31814);
xor U33135 (N_33135,N_32110,N_30819);
nand U33136 (N_33136,N_30930,N_31151);
nor U33137 (N_33137,N_32009,N_32193);
xor U33138 (N_33138,N_30452,N_31637);
nand U33139 (N_33139,N_30681,N_31876);
or U33140 (N_33140,N_32238,N_31362);
nor U33141 (N_33141,N_30968,N_31016);
nor U33142 (N_33142,N_32295,N_31903);
nor U33143 (N_33143,N_32039,N_31642);
nand U33144 (N_33144,N_30884,N_30155);
nand U33145 (N_33145,N_32371,N_31951);
nor U33146 (N_33146,N_30554,N_31845);
nor U33147 (N_33147,N_31645,N_31005);
nor U33148 (N_33148,N_31819,N_31251);
or U33149 (N_33149,N_30933,N_30860);
and U33150 (N_33150,N_32111,N_31587);
nand U33151 (N_33151,N_31946,N_32254);
or U33152 (N_33152,N_32467,N_31248);
nor U33153 (N_33153,N_32376,N_32196);
xor U33154 (N_33154,N_31757,N_30055);
or U33155 (N_33155,N_31816,N_30075);
and U33156 (N_33156,N_30539,N_31225);
nor U33157 (N_33157,N_31458,N_30166);
or U33158 (N_33158,N_30776,N_31098);
and U33159 (N_33159,N_30970,N_32200);
and U33160 (N_33160,N_30216,N_31289);
and U33161 (N_33161,N_31243,N_32038);
nand U33162 (N_33162,N_31656,N_30948);
or U33163 (N_33163,N_31216,N_30297);
xnor U33164 (N_33164,N_32417,N_30049);
or U33165 (N_33165,N_30469,N_30752);
and U33166 (N_33166,N_30925,N_31798);
xnor U33167 (N_33167,N_31448,N_30795);
and U33168 (N_33168,N_31957,N_31700);
nor U33169 (N_33169,N_32492,N_30576);
xnor U33170 (N_33170,N_30764,N_32231);
nand U33171 (N_33171,N_31958,N_30664);
xor U33172 (N_33172,N_30147,N_32412);
xor U33173 (N_33173,N_31463,N_32337);
nand U33174 (N_33174,N_30973,N_32107);
or U33175 (N_33175,N_30760,N_31968);
xnor U33176 (N_33176,N_30396,N_30673);
nand U33177 (N_33177,N_32296,N_30437);
or U33178 (N_33178,N_30685,N_30191);
and U33179 (N_33179,N_32129,N_30896);
nor U33180 (N_33180,N_30574,N_30708);
and U33181 (N_33181,N_31284,N_30701);
nor U33182 (N_33182,N_30107,N_32304);
xnor U33183 (N_33183,N_30073,N_30034);
and U33184 (N_33184,N_30436,N_30417);
or U33185 (N_33185,N_30761,N_30953);
and U33186 (N_33186,N_30196,N_32059);
nor U33187 (N_33187,N_31646,N_30662);
or U33188 (N_33188,N_31064,N_30245);
xnor U33189 (N_33189,N_31677,N_30326);
xor U33190 (N_33190,N_31371,N_30446);
xnor U33191 (N_33191,N_31492,N_30678);
and U33192 (N_33192,N_31165,N_31074);
nand U33193 (N_33193,N_32446,N_32410);
or U33194 (N_33194,N_31353,N_30520);
and U33195 (N_33195,N_31239,N_32375);
nor U33196 (N_33196,N_31320,N_31048);
or U33197 (N_33197,N_31841,N_30737);
nand U33198 (N_33198,N_31160,N_32233);
xnor U33199 (N_33199,N_30536,N_30240);
and U33200 (N_33200,N_30754,N_30278);
nand U33201 (N_33201,N_31107,N_31100);
and U33202 (N_33202,N_30286,N_30036);
xnor U33203 (N_33203,N_31485,N_30115);
nor U33204 (N_33204,N_30639,N_30838);
and U33205 (N_33205,N_32001,N_32199);
or U33206 (N_33206,N_31793,N_31335);
xor U33207 (N_33207,N_32264,N_31909);
or U33208 (N_33208,N_30653,N_30782);
nor U33209 (N_33209,N_32418,N_31842);
nand U33210 (N_33210,N_31414,N_31202);
nor U33211 (N_33211,N_32050,N_30148);
nand U33212 (N_33212,N_30535,N_30381);
xor U33213 (N_33213,N_30193,N_31854);
nor U33214 (N_33214,N_30453,N_30744);
xnor U33215 (N_33215,N_30992,N_31654);
xor U33216 (N_33216,N_30068,N_31498);
nor U33217 (N_33217,N_32239,N_30351);
and U33218 (N_33218,N_30285,N_30932);
nor U33219 (N_33219,N_31902,N_30356);
nor U33220 (N_33220,N_31698,N_30165);
xnor U33221 (N_33221,N_30214,N_31427);
nor U33222 (N_33222,N_30886,N_30958);
or U33223 (N_33223,N_30301,N_30802);
or U33224 (N_33224,N_30374,N_31121);
and U33225 (N_33225,N_31621,N_30529);
nor U33226 (N_33226,N_32267,N_31838);
nand U33227 (N_33227,N_31517,N_31670);
or U33228 (N_33228,N_31542,N_31501);
and U33229 (N_33229,N_31787,N_31885);
xor U33230 (N_33230,N_30577,N_30534);
nor U33231 (N_33231,N_32070,N_32382);
and U33232 (N_33232,N_30938,N_32455);
xor U33233 (N_33233,N_31047,N_30716);
and U33234 (N_33234,N_30013,N_30804);
xnor U33235 (N_33235,N_30704,N_30757);
or U33236 (N_33236,N_31882,N_31605);
nor U33237 (N_33237,N_30057,N_32163);
or U33238 (N_33238,N_31752,N_31298);
nand U33239 (N_33239,N_30905,N_30694);
nor U33240 (N_33240,N_30700,N_31811);
nand U33241 (N_33241,N_30002,N_30272);
xnor U33242 (N_33242,N_31129,N_30241);
xnor U33243 (N_33243,N_31836,N_31020);
xor U33244 (N_33244,N_30679,N_30179);
nor U33245 (N_33245,N_30394,N_30854);
nand U33246 (N_33246,N_31265,N_31604);
nor U33247 (N_33247,N_30482,N_32161);
nor U33248 (N_33248,N_30977,N_30758);
and U33249 (N_33249,N_30024,N_31550);
xor U33250 (N_33250,N_31620,N_32299);
and U33251 (N_33251,N_31277,N_31153);
or U33252 (N_33252,N_30507,N_32018);
or U33253 (N_33253,N_30592,N_31796);
or U33254 (N_33254,N_32242,N_31464);
and U33255 (N_33255,N_30618,N_30733);
xnor U33256 (N_33256,N_31636,N_30443);
xnor U33257 (N_33257,N_32386,N_32401);
xor U33258 (N_33258,N_30379,N_30578);
or U33259 (N_33259,N_31245,N_30986);
or U33260 (N_33260,N_31398,N_31574);
nand U33261 (N_33261,N_32392,N_31529);
nor U33262 (N_33262,N_31967,N_31649);
nor U33263 (N_33263,N_32260,N_31179);
nor U33264 (N_33264,N_31610,N_32289);
and U33265 (N_33265,N_32096,N_31553);
or U33266 (N_33266,N_32497,N_30937);
and U33267 (N_33267,N_32234,N_30438);
nor U33268 (N_33268,N_32056,N_31532);
and U33269 (N_33269,N_31377,N_30550);
nand U33270 (N_33270,N_30474,N_32331);
or U33271 (N_33271,N_30231,N_31810);
nand U33272 (N_33272,N_30857,N_31288);
nand U33273 (N_33273,N_32025,N_30208);
nor U33274 (N_33274,N_30613,N_31537);
nand U33275 (N_33275,N_30812,N_32445);
or U33276 (N_33276,N_31232,N_31618);
and U33277 (N_33277,N_32431,N_30461);
and U33278 (N_33278,N_30830,N_31241);
or U33279 (N_33279,N_31626,N_31846);
and U33280 (N_33280,N_32173,N_30902);
or U33281 (N_33281,N_31924,N_31481);
nor U33282 (N_33282,N_31435,N_31403);
nor U33283 (N_33283,N_30610,N_31519);
nor U33284 (N_33284,N_30845,N_31355);
and U33285 (N_33285,N_31365,N_32334);
or U33286 (N_33286,N_30294,N_31175);
or U33287 (N_33287,N_30234,N_30144);
nor U33288 (N_33288,N_32075,N_31285);
nor U33289 (N_33289,N_32399,N_31190);
xor U33290 (N_33290,N_31564,N_31466);
or U33291 (N_33291,N_32097,N_31504);
xnor U33292 (N_33292,N_31300,N_30590);
nor U33293 (N_33293,N_30775,N_31782);
nand U33294 (N_33294,N_31237,N_31405);
xor U33295 (N_33295,N_32215,N_30425);
nor U33296 (N_33296,N_31665,N_30428);
nand U33297 (N_33297,N_31865,N_31139);
nand U33298 (N_33298,N_32166,N_30851);
nor U33299 (N_33299,N_31119,N_30705);
nor U33300 (N_33300,N_32092,N_30478);
nor U33301 (N_33301,N_30132,N_32393);
nand U33302 (N_33302,N_32307,N_30358);
nor U33303 (N_33303,N_32398,N_31612);
or U33304 (N_33304,N_31433,N_30224);
nand U33305 (N_33305,N_31789,N_31675);
xor U33306 (N_33306,N_31374,N_32208);
nand U33307 (N_33307,N_31914,N_31465);
nor U33308 (N_33308,N_31680,N_31538);
and U33309 (N_33309,N_30514,N_31025);
nand U33310 (N_33310,N_31073,N_31849);
xnor U33311 (N_33311,N_32171,N_30321);
nand U33312 (N_33312,N_31291,N_31571);
or U33313 (N_33313,N_31029,N_30172);
and U33314 (N_33314,N_31261,N_32482);
xor U33315 (N_33315,N_31147,N_30059);
nand U33316 (N_33316,N_31728,N_32266);
nand U33317 (N_33317,N_31840,N_32311);
nand U33318 (N_33318,N_30020,N_31912);
or U33319 (N_33319,N_30961,N_31475);
nand U33320 (N_33320,N_32021,N_32017);
nor U33321 (N_33321,N_30731,N_32306);
and U33322 (N_33322,N_31771,N_31255);
or U33323 (N_33323,N_30411,N_31483);
nor U33324 (N_33324,N_30243,N_32319);
xnor U33325 (N_33325,N_30728,N_30611);
xor U33326 (N_33326,N_32182,N_31024);
nand U33327 (N_33327,N_31772,N_30344);
nand U33328 (N_33328,N_32428,N_30303);
xor U33329 (N_33329,N_32066,N_31965);
and U33330 (N_33330,N_30217,N_31136);
and U33331 (N_33331,N_31557,N_30083);
and U33332 (N_33332,N_31417,N_30898);
nor U33333 (N_33333,N_31996,N_30604);
xnor U33334 (N_33334,N_31535,N_32327);
nor U33335 (N_33335,N_30497,N_30500);
or U33336 (N_33336,N_30491,N_31821);
xnor U33337 (N_33337,N_32158,N_31635);
xnor U33338 (N_33338,N_31721,N_31660);
nand U33339 (N_33339,N_31194,N_30014);
nand U33340 (N_33340,N_31602,N_32005);
nand U33341 (N_33341,N_31296,N_31133);
xor U33342 (N_33342,N_32279,N_31290);
or U33343 (N_33343,N_30983,N_31031);
and U33344 (N_33344,N_30729,N_31668);
or U33345 (N_33345,N_32356,N_31072);
or U33346 (N_33346,N_30270,N_30799);
nor U33347 (N_33347,N_32105,N_31269);
xnor U33348 (N_33348,N_30293,N_32285);
nand U33349 (N_33349,N_30296,N_31589);
xor U33350 (N_33350,N_30090,N_31455);
nand U33351 (N_33351,N_30445,N_31565);
nand U33352 (N_33352,N_31421,N_30335);
xor U33353 (N_33353,N_31174,N_30698);
or U33354 (N_33354,N_32124,N_31835);
and U33355 (N_33355,N_31608,N_32442);
or U33356 (N_33356,N_32126,N_31011);
xor U33357 (N_33357,N_30626,N_32349);
nand U33358 (N_33358,N_30999,N_31653);
or U33359 (N_33359,N_31625,N_30118);
xnor U33360 (N_33360,N_31313,N_30212);
or U33361 (N_33361,N_31111,N_31825);
xor U33362 (N_33362,N_31858,N_31655);
and U33363 (N_33363,N_31857,N_31556);
and U33364 (N_33364,N_31071,N_30712);
nand U33365 (N_33365,N_31180,N_30636);
xor U33366 (N_33366,N_32112,N_30366);
xnor U33367 (N_33367,N_30163,N_32000);
or U33368 (N_33368,N_31766,N_31486);
or U33369 (N_33369,N_30783,N_31701);
xor U33370 (N_33370,N_30346,N_31323);
xnor U33371 (N_33371,N_30470,N_32053);
xnor U33372 (N_33372,N_30109,N_30859);
or U33373 (N_33373,N_31969,N_31693);
nand U33374 (N_33374,N_31303,N_31380);
and U33375 (N_33375,N_32054,N_30919);
nor U33376 (N_33376,N_30093,N_31860);
and U33377 (N_33377,N_31426,N_30548);
and U33378 (N_33378,N_30347,N_30085);
or U33379 (N_33379,N_32277,N_31236);
nor U33380 (N_33380,N_32152,N_30330);
or U33381 (N_33381,N_31182,N_31628);
xnor U33382 (N_33382,N_30843,N_31402);
xnor U33383 (N_33383,N_31893,N_30130);
and U33384 (N_33384,N_31022,N_31773);
xor U33385 (N_33385,N_30915,N_30399);
nor U33386 (N_33386,N_32397,N_30767);
or U33387 (N_33387,N_31505,N_32448);
or U33388 (N_33388,N_30310,N_30292);
and U33389 (N_33389,N_30994,N_31222);
nor U33390 (N_33390,N_31831,N_31271);
and U33391 (N_33391,N_31813,N_30987);
nor U33392 (N_33392,N_30518,N_30058);
nor U33393 (N_33393,N_30249,N_30945);
or U33394 (N_33394,N_31204,N_31566);
nand U33395 (N_33395,N_31314,N_31962);
and U33396 (N_33396,N_31260,N_30894);
or U33397 (N_33397,N_31760,N_32303);
or U33398 (N_33398,N_30104,N_31515);
nand U33399 (N_33399,N_30279,N_30763);
xor U33400 (N_33400,N_32154,N_31733);
or U33401 (N_33401,N_32468,N_30868);
and U33402 (N_33402,N_31588,N_31104);
nand U33403 (N_33403,N_31582,N_30495);
nand U33404 (N_33404,N_30079,N_32350);
or U33405 (N_33405,N_31322,N_31742);
and U33406 (N_33406,N_30187,N_31603);
nor U33407 (N_33407,N_32443,N_30521);
nand U33408 (N_33408,N_32069,N_30361);
nand U33409 (N_33409,N_32101,N_31747);
and U33410 (N_33410,N_31219,N_31785);
nand U33411 (N_33411,N_30164,N_32217);
xor U33412 (N_33412,N_32384,N_31961);
nand U33413 (N_33413,N_31430,N_30290);
or U33414 (N_33414,N_31452,N_30837);
and U33415 (N_33415,N_31432,N_31361);
nor U33416 (N_33416,N_31166,N_30039);
and U33417 (N_33417,N_30941,N_30269);
or U33418 (N_33418,N_32150,N_31927);
and U33419 (N_33419,N_30126,N_31545);
and U33420 (N_33420,N_31125,N_30299);
or U33421 (N_33421,N_31309,N_31093);
or U33422 (N_33422,N_30298,N_30552);
and U33423 (N_33423,N_32181,N_32162);
nor U33424 (N_33424,N_31778,N_30099);
xnor U33425 (N_33425,N_32143,N_30001);
xor U33426 (N_33426,N_32041,N_30350);
nor U33427 (N_33427,N_30596,N_31141);
nor U33428 (N_33428,N_31508,N_30416);
xor U33429 (N_33429,N_30649,N_30676);
xor U33430 (N_33430,N_31249,N_31764);
xor U33431 (N_33431,N_30464,N_31994);
or U33432 (N_33432,N_32194,N_30755);
and U33433 (N_33433,N_31338,N_30909);
nand U33434 (N_33434,N_31875,N_32104);
nand U33435 (N_33435,N_31109,N_31471);
xnor U33436 (N_33436,N_30205,N_32019);
and U33437 (N_33437,N_32322,N_31743);
or U33438 (N_33438,N_30113,N_30533);
nand U33439 (N_33439,N_30750,N_32031);
and U33440 (N_33440,N_30634,N_30519);
and U33441 (N_33441,N_30390,N_31113);
nor U33442 (N_33442,N_31404,N_31316);
and U33443 (N_33443,N_30220,N_31658);
nor U33444 (N_33444,N_30567,N_30355);
and U33445 (N_33445,N_30960,N_30317);
xnor U33446 (N_33446,N_31815,N_31955);
nand U33447 (N_33447,N_32222,N_32085);
xnor U33448 (N_33448,N_31534,N_32117);
or U33449 (N_33449,N_31294,N_30451);
nand U33450 (N_33450,N_31274,N_31980);
xor U33451 (N_33451,N_31762,N_31596);
nor U33452 (N_33452,N_30121,N_30629);
and U33453 (N_33453,N_31735,N_31514);
or U33454 (N_33454,N_30726,N_32294);
nor U33455 (N_33455,N_32119,N_32475);
nand U33456 (N_33456,N_30006,N_32144);
and U33457 (N_33457,N_31000,N_31647);
nand U33458 (N_33458,N_32227,N_30602);
nor U33459 (N_33459,N_30503,N_31663);
nor U33460 (N_33460,N_31964,N_30847);
xor U33461 (N_33461,N_30337,N_32251);
xor U33462 (N_33462,N_30900,N_32100);
and U33463 (N_33463,N_30974,N_30890);
nand U33464 (N_33464,N_32061,N_30189);
or U33465 (N_33465,N_31871,N_31512);
nor U33466 (N_33466,N_31898,N_30823);
nor U33467 (N_33467,N_31055,N_31267);
nand U33468 (N_33468,N_31078,N_32340);
and U33469 (N_33469,N_30867,N_30785);
or U33470 (N_33470,N_31956,N_31806);
nand U33471 (N_33471,N_31454,N_30872);
and U33472 (N_33472,N_31281,N_31037);
nand U33473 (N_33473,N_31039,N_31054);
nand U33474 (N_33474,N_32187,N_31667);
xnor U33475 (N_33475,N_31638,N_31711);
xnor U33476 (N_33476,N_30000,N_32247);
nand U33477 (N_33477,N_31009,N_30942);
nor U33478 (N_33478,N_30078,N_31548);
nor U33479 (N_33479,N_31524,N_32088);
and U33480 (N_33480,N_30690,N_31283);
xnor U33481 (N_33481,N_32002,N_32344);
xor U33482 (N_33482,N_30426,N_30151);
nor U33483 (N_33483,N_30677,N_31158);
or U33484 (N_33484,N_30954,N_30796);
nand U33485 (N_33485,N_31561,N_30185);
xor U33486 (N_33486,N_30174,N_32402);
or U33487 (N_33487,N_30050,N_30810);
xnor U33488 (N_33488,N_30695,N_30813);
and U33489 (N_33489,N_31036,N_31163);
or U33490 (N_33490,N_32131,N_32408);
and U33491 (N_33491,N_30345,N_30439);
xor U33492 (N_33492,N_30806,N_31873);
nand U33493 (N_33493,N_32403,N_31373);
nor U33494 (N_33494,N_32485,N_31585);
and U33495 (N_33495,N_30910,N_30255);
xnor U33496 (N_33496,N_31337,N_30652);
or U33497 (N_33497,N_31140,N_32046);
or U33498 (N_33498,N_32310,N_32185);
nor U33499 (N_33499,N_32460,N_30250);
nand U33500 (N_33500,N_31607,N_30732);
xor U33501 (N_33501,N_32345,N_31246);
xnor U33502 (N_33502,N_31094,N_31950);
nor U33503 (N_33503,N_30892,N_31050);
nand U33504 (N_33504,N_31769,N_31084);
nor U33505 (N_33505,N_32045,N_31974);
xnor U33506 (N_33506,N_31407,N_30206);
or U33507 (N_33507,N_32115,N_30724);
nand U33508 (N_33508,N_30392,N_30706);
and U33509 (N_33509,N_30621,N_31719);
nor U33510 (N_33510,N_31818,N_31619);
or U33511 (N_33511,N_30742,N_31544);
nand U33512 (N_33512,N_31349,N_30880);
nor U33513 (N_33513,N_30315,N_31018);
nor U33514 (N_33514,N_31087,N_31108);
or U33515 (N_33515,N_30956,N_32325);
and U33516 (N_33516,N_30119,N_31881);
nor U33517 (N_33517,N_32477,N_31847);
and U33518 (N_33518,N_30967,N_31344);
or U33519 (N_33519,N_30140,N_31002);
or U33520 (N_33520,N_32405,N_32204);
or U33521 (N_33521,N_30223,N_31943);
or U33522 (N_33522,N_32297,N_31013);
or U33523 (N_33523,N_32026,N_31130);
nand U33524 (N_33524,N_32336,N_30978);
nand U33525 (N_33525,N_31809,N_31710);
nor U33526 (N_33526,N_31376,N_32076);
and U33527 (N_33527,N_30273,N_30327);
or U33528 (N_33528,N_30007,N_32287);
and U33529 (N_33529,N_30328,N_30995);
or U33530 (N_33530,N_30617,N_31014);
nor U33531 (N_33531,N_30959,N_31292);
nor U33532 (N_33532,N_31993,N_31127);
or U33533 (N_33533,N_31131,N_31744);
nand U33534 (N_33534,N_30280,N_30991);
xnor U33535 (N_33535,N_32457,N_31985);
nand U33536 (N_33536,N_30781,N_30360);
nand U33537 (N_33537,N_31472,N_32298);
nand U33538 (N_33538,N_30129,N_31890);
or U33539 (N_33539,N_31531,N_31568);
nor U33540 (N_33540,N_31739,N_32074);
nand U33541 (N_33541,N_31694,N_32135);
xor U33542 (N_33542,N_31143,N_30043);
nor U33543 (N_33543,N_32481,N_32414);
nor U33544 (N_33544,N_30939,N_31057);
or U33545 (N_33545,N_31348,N_30504);
and U33546 (N_33546,N_31070,N_32432);
xnor U33547 (N_33547,N_30186,N_31518);
or U33548 (N_33548,N_31368,N_30246);
and U33549 (N_33549,N_31079,N_31878);
nor U33550 (N_33550,N_32211,N_30467);
and U33551 (N_33551,N_30606,N_31767);
nor U33552 (N_33552,N_31562,N_30322);
and U33553 (N_33553,N_30721,N_30962);
nor U33554 (N_33554,N_32495,N_31339);
and U33555 (N_33555,N_30267,N_30359);
and U33556 (N_33556,N_31696,N_30031);
xor U33557 (N_33557,N_31092,N_32406);
nand U33558 (N_33558,N_32057,N_31270);
xnor U33559 (N_33559,N_30251,N_31932);
nand U33560 (N_33560,N_30603,N_31905);
nand U33561 (N_33561,N_32014,N_31491);
or U33562 (N_33562,N_30363,N_32188);
xor U33563 (N_33563,N_32094,N_31319);
nor U33564 (N_33564,N_32071,N_30139);
nand U33565 (N_33565,N_30387,N_30753);
nand U33566 (N_33566,N_32165,N_30312);
and U33567 (N_33567,N_30309,N_30418);
nor U33568 (N_33568,N_31527,N_30091);
xnor U33569 (N_33569,N_31576,N_30110);
and U33570 (N_33570,N_30856,N_30120);
nand U33571 (N_33571,N_30125,N_31459);
nand U33572 (N_33572,N_32130,N_31476);
and U33573 (N_33573,N_31901,N_31830);
and U33574 (N_33574,N_31916,N_31164);
nor U33575 (N_33575,N_32180,N_31795);
xor U33576 (N_33576,N_31689,N_32463);
nor U33577 (N_33577,N_32249,N_31169);
nor U33578 (N_33578,N_32036,N_30222);
or U33579 (N_33579,N_31740,N_30230);
xor U33580 (N_33580,N_31128,N_32466);
nor U33581 (N_33581,N_30524,N_31208);
and U33582 (N_33582,N_32007,N_30289);
nand U33583 (N_33583,N_30826,N_30274);
nand U33584 (N_33584,N_30923,N_30211);
xor U33585 (N_33585,N_31533,N_31934);
nand U33586 (N_33586,N_31697,N_31521);
xnor U33587 (N_33587,N_31925,N_30162);
nor U33588 (N_33588,N_30979,N_32221);
nor U33589 (N_33589,N_32103,N_31080);
and U33590 (N_33590,N_31549,N_30375);
xor U33591 (N_33591,N_30116,N_32394);
or U33592 (N_33592,N_31351,N_31378);
or U33593 (N_33593,N_32441,N_31061);
xnor U33594 (N_33594,N_32190,N_30697);
nor U33595 (N_33595,N_31226,N_32276);
xor U33596 (N_33596,N_32280,N_30045);
and U33597 (N_33597,N_30364,N_31938);
and U33598 (N_33598,N_31992,N_31231);
or U33599 (N_33599,N_32183,N_30219);
and U33600 (N_33600,N_30969,N_31295);
or U33601 (N_33601,N_32407,N_31206);
and U33602 (N_33602,N_30218,N_30623);
nand U33603 (N_33603,N_30018,N_31096);
xor U33604 (N_33604,N_30797,N_31413);
or U33605 (N_33605,N_30952,N_30736);
xor U33606 (N_33606,N_32499,N_31187);
xnor U33607 (N_33607,N_31869,N_31877);
and U33608 (N_33608,N_31118,N_31489);
nand U33609 (N_33609,N_31676,N_32048);
xnor U33610 (N_33610,N_32274,N_30835);
or U33611 (N_33611,N_30516,N_31207);
or U33612 (N_33612,N_30082,N_31211);
and U33613 (N_33613,N_31662,N_31644);
and U33614 (N_33614,N_30264,N_32252);
nand U33615 (N_33615,N_30734,N_31887);
nor U33616 (N_33616,N_31683,N_30021);
and U33617 (N_33617,N_31920,N_30779);
or U33618 (N_33618,N_30870,N_32370);
nor U33619 (N_33619,N_30430,N_30226);
nor U33620 (N_33620,N_32496,N_30765);
nand U33621 (N_33621,N_32269,N_30459);
xnor U33622 (N_33622,N_30324,N_30809);
nor U33623 (N_33623,N_31516,N_31305);
nor U33624 (N_33624,N_30975,N_30040);
and U33625 (N_33625,N_32426,N_30771);
or U33626 (N_33626,N_31278,N_32367);
nor U33627 (N_33627,N_31456,N_31238);
xnor U33628 (N_33628,N_31722,N_31737);
nand U33629 (N_33629,N_32114,N_30687);
nor U33630 (N_33630,N_30194,N_31117);
or U33631 (N_33631,N_31308,N_30490);
xor U33632 (N_33632,N_30526,N_30462);
xor U33633 (N_33633,N_30371,N_30699);
xor U33634 (N_33634,N_31828,N_31509);
xor U33635 (N_33635,N_32060,N_31397);
nor U33636 (N_33636,N_30727,N_31026);
xnor U33637 (N_33637,N_30644,N_30583);
nor U33638 (N_33638,N_30190,N_30183);
nand U33639 (N_33639,N_30316,N_30789);
xnor U33640 (N_33640,N_31370,N_31317);
nand U33641 (N_33641,N_31870,N_31661);
or U33642 (N_33642,N_31824,N_32142);
nor U33643 (N_33643,N_32055,N_31273);
nand U33644 (N_33644,N_31716,N_31664);
and U33645 (N_33645,N_31684,N_30047);
xnor U33646 (N_33646,N_31275,N_32284);
xnor U33647 (N_33647,N_32316,N_32149);
or U33648 (N_33648,N_31416,N_31420);
nand U33649 (N_33649,N_30840,N_30103);
nor U33650 (N_33650,N_31137,N_30015);
and U33651 (N_33651,N_31173,N_31928);
nand U33652 (N_33652,N_30914,N_30743);
xnor U33653 (N_33653,N_30717,N_31097);
or U33654 (N_33654,N_30275,N_30655);
or U33655 (N_33655,N_31652,N_32015);
and U33656 (N_33656,N_30682,N_31918);
nor U33657 (N_33657,N_30849,N_30460);
and U33658 (N_33658,N_31062,N_31266);
xnor U33659 (N_33659,N_31110,N_31120);
and U33660 (N_33660,N_31480,N_31357);
and U33661 (N_33661,N_31200,N_30619);
and U33662 (N_33662,N_30562,N_31759);
nor U33663 (N_33663,N_32353,N_30170);
or U33664 (N_33664,N_30323,N_30527);
nor U33665 (N_33665,N_31971,N_32136);
nand U33666 (N_33666,N_30427,N_32437);
nor U33667 (N_33667,N_30471,N_30181);
xor U33668 (N_33668,N_30449,N_31583);
or U33669 (N_33669,N_32415,N_32271);
or U33670 (N_33670,N_31807,N_30415);
and U33671 (N_33671,N_31293,N_32318);
or U33672 (N_33672,N_31075,N_30105);
and U33673 (N_33673,N_31930,N_32478);
or U33674 (N_33674,N_32012,N_30010);
xor U33675 (N_33675,N_31978,N_31843);
xnor U33676 (N_33676,N_30751,N_30566);
nand U33677 (N_33677,N_30086,N_31046);
nor U33678 (N_33678,N_32065,N_31991);
xnor U33679 (N_33679,N_30530,N_31101);
and U33680 (N_33680,N_32044,N_32095);
and U33681 (N_33681,N_31388,N_32177);
or U33682 (N_33682,N_30853,N_30339);
and U33683 (N_33683,N_31228,N_31756);
and U33684 (N_33684,N_30601,N_31797);
nor U33685 (N_33685,N_30291,N_31450);
and U33686 (N_33686,N_30477,N_30773);
or U33687 (N_33687,N_30573,N_30496);
and U33688 (N_33688,N_30011,N_31705);
xor U33689 (N_33689,N_31651,N_32409);
nor U33690 (N_33690,N_31105,N_30401);
nor U33691 (N_33691,N_31879,N_31198);
nor U33692 (N_33692,N_30060,N_31931);
or U33693 (N_33693,N_30730,N_30963);
and U33694 (N_33694,N_30633,N_31001);
or U33695 (N_33695,N_31803,N_31205);
nor U33696 (N_33696,N_30201,N_32471);
xor U33697 (N_33697,N_31331,N_30198);
and U33698 (N_33698,N_30517,N_31640);
xnor U33699 (N_33699,N_30553,N_31033);
xor U33700 (N_33700,N_32315,N_32305);
nand U33701 (N_33701,N_30780,N_32108);
or U33702 (N_33702,N_32465,N_30197);
or U33703 (N_33703,N_31354,N_32205);
xor U33704 (N_33704,N_30156,N_30100);
nor U33705 (N_33705,N_30627,N_30684);
xnor U33706 (N_33706,N_30591,N_31063);
nand U33707 (N_33707,N_32210,N_32156);
nand U33708 (N_33708,N_30689,N_30256);
xnor U33709 (N_33709,N_31708,N_31439);
and U33710 (N_33710,N_30238,N_31998);
or U33711 (N_33711,N_30873,N_31748);
nand U33712 (N_33712,N_30989,N_30029);
nand U33713 (N_33713,N_31395,N_30828);
nor U33714 (N_33714,N_30150,N_31899);
xnor U33715 (N_33715,N_31570,N_31215);
xnor U33716 (N_33716,N_31482,N_31581);
nor U33717 (N_33717,N_30693,N_31264);
nor U33718 (N_33718,N_31257,N_30547);
and U33719 (N_33719,N_31983,N_30735);
nand U33720 (N_33720,N_30261,N_30786);
nor U33721 (N_33721,N_31861,N_30175);
or U33722 (N_33722,N_32424,N_31786);
or U33723 (N_33723,N_30688,N_31586);
and U33724 (N_33724,N_32483,N_32263);
nand U33725 (N_33725,N_32137,N_30599);
nand U33726 (N_33726,N_32212,N_31425);
and U33727 (N_33727,N_31007,N_31758);
nand U33728 (N_33728,N_31189,N_31366);
xor U33729 (N_33729,N_31982,N_32098);
nand U33730 (N_33730,N_30615,N_31572);
nand U33731 (N_33731,N_31122,N_30380);
nor U33732 (N_33732,N_30200,N_32425);
nor U33733 (N_33733,N_31461,N_30588);
and U33734 (N_33734,N_30028,N_31068);
xor U33735 (N_33735,N_31234,N_30921);
nand U33736 (N_33736,N_30253,N_30587);
and U33737 (N_33737,N_31933,N_31558);
nand U33738 (N_33738,N_30966,N_31754);
nor U33739 (N_33739,N_32030,N_31088);
or U33740 (N_33740,N_32237,N_32225);
nor U33741 (N_33741,N_30331,N_30252);
and U33742 (N_33742,N_31340,N_30628);
or U33743 (N_33743,N_32079,N_30229);
nor U33744 (N_33744,N_31259,N_30137);
and U33745 (N_33745,N_31042,N_30822);
nor U33746 (N_33746,N_31755,N_32373);
and U33747 (N_33747,N_32436,N_31447);
xor U33748 (N_33748,N_31488,N_31889);
nor U33749 (N_33749,N_30675,N_30976);
nor U33750 (N_33750,N_32379,N_31996);
and U33751 (N_33751,N_30119,N_31390);
nor U33752 (N_33752,N_32167,N_32142);
xnor U33753 (N_33753,N_32470,N_31240);
nand U33754 (N_33754,N_30656,N_31075);
nor U33755 (N_33755,N_30339,N_32284);
or U33756 (N_33756,N_31674,N_31585);
or U33757 (N_33757,N_31320,N_31091);
nand U33758 (N_33758,N_30727,N_32111);
xor U33759 (N_33759,N_30492,N_31781);
or U33760 (N_33760,N_31768,N_31843);
nand U33761 (N_33761,N_30230,N_31929);
and U33762 (N_33762,N_31031,N_31040);
or U33763 (N_33763,N_32334,N_32003);
nor U33764 (N_33764,N_30526,N_30536);
nor U33765 (N_33765,N_31494,N_30659);
or U33766 (N_33766,N_30992,N_30125);
and U33767 (N_33767,N_32259,N_30551);
xnor U33768 (N_33768,N_31181,N_31144);
nor U33769 (N_33769,N_31271,N_30299);
xor U33770 (N_33770,N_31626,N_30188);
and U33771 (N_33771,N_32006,N_31052);
nor U33772 (N_33772,N_30256,N_30403);
or U33773 (N_33773,N_31886,N_30625);
nor U33774 (N_33774,N_31134,N_31859);
and U33775 (N_33775,N_30722,N_30509);
nand U33776 (N_33776,N_31995,N_30178);
xnor U33777 (N_33777,N_32334,N_32191);
nor U33778 (N_33778,N_30664,N_30602);
nor U33779 (N_33779,N_31669,N_31168);
xnor U33780 (N_33780,N_30665,N_31524);
and U33781 (N_33781,N_31885,N_31630);
xor U33782 (N_33782,N_30805,N_31588);
or U33783 (N_33783,N_30092,N_30279);
nor U33784 (N_33784,N_30918,N_30238);
xor U33785 (N_33785,N_32257,N_30988);
xor U33786 (N_33786,N_32065,N_32210);
nand U33787 (N_33787,N_32402,N_30598);
nor U33788 (N_33788,N_30562,N_30545);
xor U33789 (N_33789,N_30446,N_30653);
nor U33790 (N_33790,N_31524,N_30475);
nor U33791 (N_33791,N_31928,N_31963);
or U33792 (N_33792,N_31399,N_30439);
and U33793 (N_33793,N_30793,N_31687);
xor U33794 (N_33794,N_31600,N_30727);
nor U33795 (N_33795,N_30466,N_30333);
and U33796 (N_33796,N_30372,N_31238);
or U33797 (N_33797,N_31274,N_31104);
and U33798 (N_33798,N_31756,N_30987);
or U33799 (N_33799,N_30782,N_31867);
xor U33800 (N_33800,N_30428,N_30074);
and U33801 (N_33801,N_31444,N_31109);
nor U33802 (N_33802,N_32309,N_30310);
nor U33803 (N_33803,N_31063,N_32393);
nand U33804 (N_33804,N_30506,N_32167);
nor U33805 (N_33805,N_30897,N_31769);
nor U33806 (N_33806,N_31667,N_32038);
or U33807 (N_33807,N_30771,N_32496);
and U33808 (N_33808,N_30381,N_31506);
nand U33809 (N_33809,N_30848,N_31549);
or U33810 (N_33810,N_32293,N_31071);
nor U33811 (N_33811,N_30159,N_30261);
xnor U33812 (N_33812,N_31619,N_30312);
and U33813 (N_33813,N_31925,N_31691);
nand U33814 (N_33814,N_30353,N_31234);
or U33815 (N_33815,N_31218,N_31533);
xor U33816 (N_33816,N_32264,N_31083);
xnor U33817 (N_33817,N_30363,N_31630);
or U33818 (N_33818,N_32287,N_31051);
nor U33819 (N_33819,N_30301,N_31250);
xor U33820 (N_33820,N_30665,N_31384);
and U33821 (N_33821,N_31319,N_30986);
or U33822 (N_33822,N_32157,N_31867);
xnor U33823 (N_33823,N_32029,N_31191);
or U33824 (N_33824,N_31466,N_31101);
nand U33825 (N_33825,N_31241,N_32217);
xnor U33826 (N_33826,N_32079,N_31728);
nand U33827 (N_33827,N_31532,N_32264);
or U33828 (N_33828,N_31559,N_31772);
or U33829 (N_33829,N_32455,N_30620);
nand U33830 (N_33830,N_31846,N_30053);
xnor U33831 (N_33831,N_30353,N_31138);
nand U33832 (N_33832,N_31205,N_32053);
nor U33833 (N_33833,N_30346,N_32127);
xnor U33834 (N_33834,N_30947,N_30288);
nand U33835 (N_33835,N_32422,N_30508);
xnor U33836 (N_33836,N_31077,N_31944);
nor U33837 (N_33837,N_31527,N_32289);
nor U33838 (N_33838,N_31117,N_31279);
xor U33839 (N_33839,N_31958,N_31003);
nor U33840 (N_33840,N_30758,N_30170);
xnor U33841 (N_33841,N_30322,N_30825);
and U33842 (N_33842,N_32354,N_32201);
and U33843 (N_33843,N_32272,N_30815);
xor U33844 (N_33844,N_30268,N_31487);
xor U33845 (N_33845,N_31705,N_32027);
and U33846 (N_33846,N_31255,N_30889);
nor U33847 (N_33847,N_31812,N_30164);
nor U33848 (N_33848,N_30724,N_30578);
xor U33849 (N_33849,N_30905,N_30759);
nand U33850 (N_33850,N_31841,N_31432);
xnor U33851 (N_33851,N_31021,N_31706);
or U33852 (N_33852,N_30152,N_30075);
nor U33853 (N_33853,N_32475,N_30911);
nor U33854 (N_33854,N_31276,N_31345);
and U33855 (N_33855,N_30858,N_30634);
and U33856 (N_33856,N_31018,N_32189);
nor U33857 (N_33857,N_32032,N_31596);
xnor U33858 (N_33858,N_32302,N_31553);
and U33859 (N_33859,N_30302,N_30372);
or U33860 (N_33860,N_31794,N_30265);
or U33861 (N_33861,N_31020,N_31066);
and U33862 (N_33862,N_32364,N_31526);
or U33863 (N_33863,N_30299,N_30494);
nand U33864 (N_33864,N_30746,N_31264);
nor U33865 (N_33865,N_32000,N_30996);
xor U33866 (N_33866,N_30896,N_32396);
nand U33867 (N_33867,N_31422,N_31478);
or U33868 (N_33868,N_30331,N_30264);
xnor U33869 (N_33869,N_30447,N_32100);
and U33870 (N_33870,N_31889,N_31611);
xnor U33871 (N_33871,N_30548,N_30404);
or U33872 (N_33872,N_30435,N_31317);
xnor U33873 (N_33873,N_30362,N_32374);
nor U33874 (N_33874,N_30132,N_32084);
or U33875 (N_33875,N_30611,N_30145);
and U33876 (N_33876,N_31243,N_32212);
xor U33877 (N_33877,N_31905,N_30688);
nor U33878 (N_33878,N_31248,N_30335);
nor U33879 (N_33879,N_30270,N_31249);
nor U33880 (N_33880,N_32338,N_31577);
and U33881 (N_33881,N_31690,N_31915);
xnor U33882 (N_33882,N_30210,N_32144);
or U33883 (N_33883,N_32372,N_30385);
nand U33884 (N_33884,N_30595,N_31277);
xnor U33885 (N_33885,N_30493,N_30398);
and U33886 (N_33886,N_31464,N_30201);
xnor U33887 (N_33887,N_32124,N_30403);
nor U33888 (N_33888,N_32485,N_32191);
nand U33889 (N_33889,N_32027,N_30917);
nor U33890 (N_33890,N_31982,N_31882);
nor U33891 (N_33891,N_32466,N_31155);
nand U33892 (N_33892,N_31179,N_31200);
and U33893 (N_33893,N_31534,N_31514);
xor U33894 (N_33894,N_30290,N_30444);
xor U33895 (N_33895,N_31536,N_30924);
and U33896 (N_33896,N_31242,N_30658);
xnor U33897 (N_33897,N_32284,N_31798);
or U33898 (N_33898,N_31866,N_31783);
xnor U33899 (N_33899,N_31929,N_32149);
nand U33900 (N_33900,N_30553,N_31916);
nor U33901 (N_33901,N_32028,N_32021);
and U33902 (N_33902,N_30658,N_30691);
and U33903 (N_33903,N_30264,N_30779);
nor U33904 (N_33904,N_31903,N_30285);
nor U33905 (N_33905,N_30205,N_31107);
xnor U33906 (N_33906,N_30240,N_31267);
xnor U33907 (N_33907,N_31030,N_31193);
nor U33908 (N_33908,N_32447,N_31349);
or U33909 (N_33909,N_30315,N_31853);
nand U33910 (N_33910,N_30349,N_30072);
nor U33911 (N_33911,N_32050,N_31745);
and U33912 (N_33912,N_32226,N_30242);
xnor U33913 (N_33913,N_30762,N_32470);
and U33914 (N_33914,N_30031,N_31205);
nand U33915 (N_33915,N_30100,N_31298);
nand U33916 (N_33916,N_32307,N_31106);
xnor U33917 (N_33917,N_31419,N_30338);
nand U33918 (N_33918,N_31466,N_31235);
xnor U33919 (N_33919,N_30765,N_32326);
or U33920 (N_33920,N_31814,N_31476);
nor U33921 (N_33921,N_30780,N_30996);
or U33922 (N_33922,N_31031,N_30650);
and U33923 (N_33923,N_32243,N_31527);
nand U33924 (N_33924,N_31411,N_31227);
or U33925 (N_33925,N_31712,N_30690);
and U33926 (N_33926,N_30939,N_30234);
nor U33927 (N_33927,N_31113,N_32272);
xor U33928 (N_33928,N_30277,N_30131);
or U33929 (N_33929,N_32387,N_31162);
nand U33930 (N_33930,N_30648,N_30855);
nand U33931 (N_33931,N_31712,N_31163);
nor U33932 (N_33932,N_31220,N_31995);
xnor U33933 (N_33933,N_30057,N_30866);
or U33934 (N_33934,N_30048,N_32163);
nor U33935 (N_33935,N_30514,N_30168);
nor U33936 (N_33936,N_30263,N_32144);
or U33937 (N_33937,N_32207,N_30787);
nand U33938 (N_33938,N_30505,N_32407);
xnor U33939 (N_33939,N_32318,N_31212);
or U33940 (N_33940,N_30546,N_31739);
or U33941 (N_33941,N_30418,N_31484);
nor U33942 (N_33942,N_31397,N_32487);
and U33943 (N_33943,N_30989,N_30656);
and U33944 (N_33944,N_31504,N_30883);
nand U33945 (N_33945,N_30856,N_30837);
nor U33946 (N_33946,N_31909,N_31044);
xor U33947 (N_33947,N_30157,N_31154);
nand U33948 (N_33948,N_30921,N_31897);
and U33949 (N_33949,N_31757,N_31524);
xor U33950 (N_33950,N_31897,N_30375);
xor U33951 (N_33951,N_30361,N_30752);
and U33952 (N_33952,N_31743,N_30410);
nor U33953 (N_33953,N_30768,N_31343);
nor U33954 (N_33954,N_31767,N_31418);
nand U33955 (N_33955,N_30766,N_30053);
or U33956 (N_33956,N_31544,N_31564);
or U33957 (N_33957,N_31379,N_30279);
or U33958 (N_33958,N_32372,N_30318);
nand U33959 (N_33959,N_32030,N_31278);
and U33960 (N_33960,N_31841,N_30790);
xnor U33961 (N_33961,N_30544,N_30305);
nor U33962 (N_33962,N_31574,N_30137);
nor U33963 (N_33963,N_31178,N_30651);
and U33964 (N_33964,N_31488,N_30197);
or U33965 (N_33965,N_31584,N_31170);
nand U33966 (N_33966,N_32462,N_31738);
or U33967 (N_33967,N_32443,N_30425);
nor U33968 (N_33968,N_31776,N_31084);
nor U33969 (N_33969,N_31416,N_31729);
nand U33970 (N_33970,N_30747,N_31999);
nand U33971 (N_33971,N_30345,N_30639);
nand U33972 (N_33972,N_31708,N_32061);
and U33973 (N_33973,N_31251,N_30934);
nand U33974 (N_33974,N_31241,N_32197);
or U33975 (N_33975,N_30025,N_30841);
and U33976 (N_33976,N_31026,N_32417);
nand U33977 (N_33977,N_32477,N_32033);
or U33978 (N_33978,N_31274,N_31649);
nand U33979 (N_33979,N_30138,N_31324);
nand U33980 (N_33980,N_31226,N_30315);
nand U33981 (N_33981,N_30141,N_32218);
and U33982 (N_33982,N_31109,N_31402);
and U33983 (N_33983,N_31814,N_32174);
xor U33984 (N_33984,N_31340,N_30607);
xor U33985 (N_33985,N_30085,N_32185);
nand U33986 (N_33986,N_32058,N_31841);
nor U33987 (N_33987,N_31704,N_30982);
nand U33988 (N_33988,N_32208,N_31507);
xnor U33989 (N_33989,N_30391,N_30111);
or U33990 (N_33990,N_31536,N_30368);
nor U33991 (N_33991,N_31583,N_31484);
and U33992 (N_33992,N_30934,N_30761);
xnor U33993 (N_33993,N_30706,N_32402);
nor U33994 (N_33994,N_31862,N_30537);
nand U33995 (N_33995,N_30825,N_30932);
nand U33996 (N_33996,N_31527,N_31579);
nor U33997 (N_33997,N_30942,N_30491);
xnor U33998 (N_33998,N_32317,N_32226);
xnor U33999 (N_33999,N_31026,N_31930);
nand U34000 (N_34000,N_31524,N_30846);
or U34001 (N_34001,N_30987,N_30907);
xnor U34002 (N_34002,N_32290,N_32167);
or U34003 (N_34003,N_30409,N_32124);
xnor U34004 (N_34004,N_31109,N_31326);
xnor U34005 (N_34005,N_32106,N_32450);
and U34006 (N_34006,N_31257,N_30890);
nor U34007 (N_34007,N_30825,N_31260);
xnor U34008 (N_34008,N_30803,N_32492);
and U34009 (N_34009,N_32438,N_31707);
nand U34010 (N_34010,N_31925,N_31468);
or U34011 (N_34011,N_31988,N_30610);
nor U34012 (N_34012,N_31668,N_31054);
or U34013 (N_34013,N_32113,N_30526);
and U34014 (N_34014,N_32480,N_32422);
and U34015 (N_34015,N_32434,N_31811);
or U34016 (N_34016,N_30176,N_31903);
xor U34017 (N_34017,N_32481,N_31059);
nor U34018 (N_34018,N_30270,N_32086);
and U34019 (N_34019,N_30996,N_30435);
xor U34020 (N_34020,N_30627,N_30434);
xnor U34021 (N_34021,N_30263,N_31560);
xor U34022 (N_34022,N_31853,N_31204);
or U34023 (N_34023,N_31181,N_32048);
xnor U34024 (N_34024,N_30433,N_30456);
nand U34025 (N_34025,N_30715,N_30684);
and U34026 (N_34026,N_31737,N_32279);
nand U34027 (N_34027,N_31432,N_31304);
xnor U34028 (N_34028,N_32209,N_31228);
nand U34029 (N_34029,N_30243,N_30659);
nand U34030 (N_34030,N_31363,N_30575);
and U34031 (N_34031,N_32169,N_31810);
xnor U34032 (N_34032,N_30503,N_31835);
or U34033 (N_34033,N_32085,N_32061);
nor U34034 (N_34034,N_30473,N_32352);
nor U34035 (N_34035,N_32493,N_30514);
or U34036 (N_34036,N_32373,N_31729);
nor U34037 (N_34037,N_31910,N_30114);
nor U34038 (N_34038,N_32015,N_30285);
nor U34039 (N_34039,N_32050,N_31123);
or U34040 (N_34040,N_30451,N_30832);
nor U34041 (N_34041,N_31047,N_30076);
nor U34042 (N_34042,N_30155,N_30026);
or U34043 (N_34043,N_31756,N_30567);
xor U34044 (N_34044,N_32110,N_30598);
and U34045 (N_34045,N_30543,N_31267);
and U34046 (N_34046,N_30272,N_31283);
and U34047 (N_34047,N_31659,N_31732);
or U34048 (N_34048,N_32423,N_31249);
or U34049 (N_34049,N_32413,N_30001);
nor U34050 (N_34050,N_30460,N_31772);
or U34051 (N_34051,N_31993,N_30527);
nand U34052 (N_34052,N_31603,N_32021);
nand U34053 (N_34053,N_31853,N_31988);
and U34054 (N_34054,N_30965,N_31432);
nor U34055 (N_34055,N_32041,N_31813);
nor U34056 (N_34056,N_30334,N_32313);
nor U34057 (N_34057,N_31224,N_31162);
nand U34058 (N_34058,N_30075,N_31152);
nor U34059 (N_34059,N_32061,N_31794);
and U34060 (N_34060,N_32277,N_31072);
nand U34061 (N_34061,N_32039,N_31655);
xor U34062 (N_34062,N_31805,N_31507);
nor U34063 (N_34063,N_30763,N_30560);
nand U34064 (N_34064,N_31786,N_31865);
nand U34065 (N_34065,N_31560,N_31954);
nand U34066 (N_34066,N_31588,N_32013);
xor U34067 (N_34067,N_31227,N_31099);
or U34068 (N_34068,N_30447,N_30624);
or U34069 (N_34069,N_32446,N_30958);
nor U34070 (N_34070,N_31947,N_31639);
nand U34071 (N_34071,N_30655,N_31487);
nor U34072 (N_34072,N_30042,N_30889);
and U34073 (N_34073,N_31300,N_30681);
nor U34074 (N_34074,N_30196,N_31781);
nor U34075 (N_34075,N_32417,N_30626);
or U34076 (N_34076,N_30450,N_30050);
nand U34077 (N_34077,N_32093,N_31597);
nand U34078 (N_34078,N_30127,N_31086);
and U34079 (N_34079,N_31794,N_30311);
nor U34080 (N_34080,N_32214,N_32183);
or U34081 (N_34081,N_31623,N_32158);
xor U34082 (N_34082,N_30122,N_31687);
xnor U34083 (N_34083,N_31928,N_30082);
nor U34084 (N_34084,N_31528,N_30153);
nor U34085 (N_34085,N_31697,N_30579);
nand U34086 (N_34086,N_31830,N_32300);
nor U34087 (N_34087,N_31324,N_30558);
or U34088 (N_34088,N_30323,N_31302);
nor U34089 (N_34089,N_32103,N_31848);
xnor U34090 (N_34090,N_30228,N_30550);
nand U34091 (N_34091,N_32042,N_30001);
and U34092 (N_34092,N_31073,N_32125);
nor U34093 (N_34093,N_31769,N_30399);
and U34094 (N_34094,N_31729,N_30834);
nor U34095 (N_34095,N_32224,N_32152);
and U34096 (N_34096,N_31365,N_31497);
nand U34097 (N_34097,N_31190,N_30778);
and U34098 (N_34098,N_30856,N_30440);
and U34099 (N_34099,N_31535,N_31115);
nor U34100 (N_34100,N_30110,N_30528);
xnor U34101 (N_34101,N_32029,N_31180);
xor U34102 (N_34102,N_31761,N_30913);
and U34103 (N_34103,N_30859,N_32477);
xnor U34104 (N_34104,N_32216,N_31336);
and U34105 (N_34105,N_32014,N_31729);
nand U34106 (N_34106,N_30435,N_31343);
nor U34107 (N_34107,N_30758,N_30876);
or U34108 (N_34108,N_32212,N_30879);
or U34109 (N_34109,N_30280,N_30754);
or U34110 (N_34110,N_31774,N_30563);
nor U34111 (N_34111,N_30856,N_31082);
nor U34112 (N_34112,N_30984,N_32167);
xnor U34113 (N_34113,N_30325,N_31989);
or U34114 (N_34114,N_30454,N_31159);
xor U34115 (N_34115,N_31953,N_30416);
nor U34116 (N_34116,N_30125,N_31364);
xnor U34117 (N_34117,N_31624,N_30309);
nor U34118 (N_34118,N_31920,N_31727);
nand U34119 (N_34119,N_31753,N_30612);
xnor U34120 (N_34120,N_30355,N_30609);
nor U34121 (N_34121,N_30663,N_31468);
and U34122 (N_34122,N_32270,N_32401);
nor U34123 (N_34123,N_30903,N_31054);
xor U34124 (N_34124,N_31307,N_31995);
nand U34125 (N_34125,N_30445,N_30701);
and U34126 (N_34126,N_32456,N_32478);
or U34127 (N_34127,N_31777,N_32392);
xnor U34128 (N_34128,N_32270,N_31373);
and U34129 (N_34129,N_32486,N_31987);
nor U34130 (N_34130,N_32475,N_32270);
xor U34131 (N_34131,N_31775,N_31883);
or U34132 (N_34132,N_30154,N_31114);
or U34133 (N_34133,N_32002,N_31225);
and U34134 (N_34134,N_31192,N_30577);
nand U34135 (N_34135,N_30251,N_31017);
and U34136 (N_34136,N_30377,N_31620);
xnor U34137 (N_34137,N_30233,N_30929);
nand U34138 (N_34138,N_31987,N_31114);
xor U34139 (N_34139,N_31911,N_30169);
and U34140 (N_34140,N_30206,N_32419);
and U34141 (N_34141,N_30841,N_31035);
nand U34142 (N_34142,N_30465,N_31460);
or U34143 (N_34143,N_32382,N_30638);
xnor U34144 (N_34144,N_31124,N_31742);
nand U34145 (N_34145,N_32243,N_32180);
and U34146 (N_34146,N_30070,N_32445);
xor U34147 (N_34147,N_32429,N_31209);
or U34148 (N_34148,N_31659,N_30020);
and U34149 (N_34149,N_32004,N_31469);
nand U34150 (N_34150,N_30449,N_31253);
xor U34151 (N_34151,N_32044,N_31890);
nand U34152 (N_34152,N_30928,N_31086);
xor U34153 (N_34153,N_30026,N_30038);
xor U34154 (N_34154,N_32473,N_30357);
or U34155 (N_34155,N_30031,N_31000);
and U34156 (N_34156,N_30160,N_32372);
or U34157 (N_34157,N_30851,N_30158);
xnor U34158 (N_34158,N_30840,N_30356);
or U34159 (N_34159,N_30080,N_31526);
nor U34160 (N_34160,N_30574,N_30776);
or U34161 (N_34161,N_31454,N_30249);
xor U34162 (N_34162,N_30038,N_31843);
xnor U34163 (N_34163,N_30504,N_32292);
xnor U34164 (N_34164,N_32152,N_30176);
or U34165 (N_34165,N_30231,N_30529);
xnor U34166 (N_34166,N_31967,N_31454);
nor U34167 (N_34167,N_31917,N_31457);
xor U34168 (N_34168,N_30521,N_32370);
nor U34169 (N_34169,N_31871,N_31599);
xnor U34170 (N_34170,N_31887,N_31261);
xor U34171 (N_34171,N_31566,N_30447);
nor U34172 (N_34172,N_30256,N_31485);
and U34173 (N_34173,N_30931,N_30175);
nor U34174 (N_34174,N_30154,N_31269);
nand U34175 (N_34175,N_32106,N_32351);
nor U34176 (N_34176,N_30417,N_31785);
xor U34177 (N_34177,N_32268,N_30507);
and U34178 (N_34178,N_30483,N_31899);
nor U34179 (N_34179,N_31406,N_31062);
nor U34180 (N_34180,N_31491,N_30561);
and U34181 (N_34181,N_32158,N_30238);
xnor U34182 (N_34182,N_30661,N_32041);
or U34183 (N_34183,N_32139,N_31499);
xnor U34184 (N_34184,N_31737,N_30645);
nand U34185 (N_34185,N_30259,N_31449);
nand U34186 (N_34186,N_31843,N_30633);
and U34187 (N_34187,N_31295,N_30719);
nand U34188 (N_34188,N_30567,N_30500);
nand U34189 (N_34189,N_32488,N_30718);
and U34190 (N_34190,N_32196,N_31022);
nor U34191 (N_34191,N_30828,N_31437);
nand U34192 (N_34192,N_31333,N_31234);
or U34193 (N_34193,N_31482,N_30343);
xnor U34194 (N_34194,N_30538,N_32420);
nor U34195 (N_34195,N_30507,N_32356);
and U34196 (N_34196,N_30188,N_31800);
and U34197 (N_34197,N_30046,N_31878);
nor U34198 (N_34198,N_31649,N_30884);
nand U34199 (N_34199,N_30034,N_31885);
xor U34200 (N_34200,N_31700,N_31514);
xor U34201 (N_34201,N_31727,N_32393);
nor U34202 (N_34202,N_30685,N_30892);
nor U34203 (N_34203,N_30568,N_31694);
nand U34204 (N_34204,N_30361,N_32336);
and U34205 (N_34205,N_30996,N_30933);
and U34206 (N_34206,N_31911,N_31677);
or U34207 (N_34207,N_30992,N_31270);
xnor U34208 (N_34208,N_30290,N_31179);
or U34209 (N_34209,N_30161,N_31004);
nor U34210 (N_34210,N_30119,N_31961);
xnor U34211 (N_34211,N_31128,N_30756);
xor U34212 (N_34212,N_31007,N_32145);
and U34213 (N_34213,N_31471,N_30886);
nand U34214 (N_34214,N_32247,N_30510);
nand U34215 (N_34215,N_31021,N_31488);
or U34216 (N_34216,N_30022,N_32351);
or U34217 (N_34217,N_31270,N_30975);
or U34218 (N_34218,N_31267,N_31538);
nand U34219 (N_34219,N_30935,N_30527);
and U34220 (N_34220,N_30548,N_32225);
nand U34221 (N_34221,N_30177,N_30831);
nand U34222 (N_34222,N_31744,N_31635);
nand U34223 (N_34223,N_32379,N_30922);
or U34224 (N_34224,N_31617,N_30102);
and U34225 (N_34225,N_32370,N_31042);
or U34226 (N_34226,N_31854,N_31839);
xnor U34227 (N_34227,N_31065,N_30733);
nor U34228 (N_34228,N_31993,N_30696);
and U34229 (N_34229,N_31302,N_31409);
xor U34230 (N_34230,N_31475,N_31802);
nand U34231 (N_34231,N_32093,N_31169);
and U34232 (N_34232,N_32221,N_31520);
nor U34233 (N_34233,N_30577,N_30789);
nand U34234 (N_34234,N_32312,N_32382);
nor U34235 (N_34235,N_31463,N_30453);
xor U34236 (N_34236,N_30921,N_32178);
or U34237 (N_34237,N_32109,N_31203);
nor U34238 (N_34238,N_30332,N_31096);
nor U34239 (N_34239,N_32075,N_31199);
or U34240 (N_34240,N_30011,N_30417);
nor U34241 (N_34241,N_30069,N_31409);
nor U34242 (N_34242,N_30449,N_31333);
xor U34243 (N_34243,N_30911,N_30480);
xnor U34244 (N_34244,N_32081,N_31706);
nor U34245 (N_34245,N_31013,N_31971);
nor U34246 (N_34246,N_30956,N_31435);
nor U34247 (N_34247,N_31972,N_31425);
xnor U34248 (N_34248,N_30931,N_30325);
nor U34249 (N_34249,N_30364,N_30280);
and U34250 (N_34250,N_31728,N_31255);
nand U34251 (N_34251,N_31051,N_30974);
nand U34252 (N_34252,N_31032,N_31567);
or U34253 (N_34253,N_31522,N_31878);
or U34254 (N_34254,N_32243,N_31134);
nand U34255 (N_34255,N_31812,N_32194);
and U34256 (N_34256,N_31628,N_32069);
nor U34257 (N_34257,N_30317,N_32435);
nor U34258 (N_34258,N_30984,N_30024);
nor U34259 (N_34259,N_31640,N_30097);
or U34260 (N_34260,N_31592,N_32349);
and U34261 (N_34261,N_31662,N_30133);
or U34262 (N_34262,N_30829,N_31969);
xor U34263 (N_34263,N_30735,N_32150);
nand U34264 (N_34264,N_32434,N_32359);
or U34265 (N_34265,N_30450,N_30629);
or U34266 (N_34266,N_31934,N_31744);
nand U34267 (N_34267,N_32222,N_31217);
xnor U34268 (N_34268,N_31019,N_30489);
or U34269 (N_34269,N_30674,N_31172);
nor U34270 (N_34270,N_30371,N_31493);
and U34271 (N_34271,N_31624,N_30087);
xor U34272 (N_34272,N_31020,N_30893);
or U34273 (N_34273,N_31921,N_30929);
nand U34274 (N_34274,N_30438,N_32404);
xnor U34275 (N_34275,N_30001,N_30135);
nor U34276 (N_34276,N_30636,N_32187);
or U34277 (N_34277,N_31075,N_31451);
xnor U34278 (N_34278,N_30152,N_30355);
xor U34279 (N_34279,N_32248,N_32348);
nor U34280 (N_34280,N_30010,N_30794);
and U34281 (N_34281,N_30788,N_31143);
and U34282 (N_34282,N_32090,N_31603);
nor U34283 (N_34283,N_30517,N_30737);
xnor U34284 (N_34284,N_31789,N_30536);
or U34285 (N_34285,N_31342,N_31799);
nor U34286 (N_34286,N_31943,N_32103);
xnor U34287 (N_34287,N_30757,N_31939);
nand U34288 (N_34288,N_31926,N_31146);
or U34289 (N_34289,N_31615,N_30438);
or U34290 (N_34290,N_31608,N_31909);
xor U34291 (N_34291,N_31266,N_32422);
nand U34292 (N_34292,N_31523,N_30674);
and U34293 (N_34293,N_31773,N_31180);
or U34294 (N_34294,N_30125,N_31124);
and U34295 (N_34295,N_31278,N_32320);
nand U34296 (N_34296,N_30539,N_32220);
and U34297 (N_34297,N_30386,N_31309);
and U34298 (N_34298,N_31423,N_31091);
nand U34299 (N_34299,N_30634,N_30318);
nor U34300 (N_34300,N_30106,N_31029);
nor U34301 (N_34301,N_32368,N_30327);
or U34302 (N_34302,N_32023,N_30809);
nand U34303 (N_34303,N_32335,N_30286);
and U34304 (N_34304,N_31000,N_32495);
or U34305 (N_34305,N_30348,N_30072);
nand U34306 (N_34306,N_31075,N_30122);
nor U34307 (N_34307,N_32267,N_30727);
or U34308 (N_34308,N_30473,N_31729);
and U34309 (N_34309,N_31785,N_31671);
or U34310 (N_34310,N_32135,N_31078);
nand U34311 (N_34311,N_31390,N_31526);
or U34312 (N_34312,N_30356,N_32147);
and U34313 (N_34313,N_31093,N_31278);
xor U34314 (N_34314,N_31865,N_30231);
nor U34315 (N_34315,N_30465,N_32373);
or U34316 (N_34316,N_30713,N_31737);
or U34317 (N_34317,N_30804,N_32043);
or U34318 (N_34318,N_31109,N_31731);
and U34319 (N_34319,N_31991,N_31444);
or U34320 (N_34320,N_32239,N_30265);
and U34321 (N_34321,N_32428,N_30098);
or U34322 (N_34322,N_30798,N_31054);
nor U34323 (N_34323,N_30591,N_32499);
nor U34324 (N_34324,N_32226,N_32380);
nor U34325 (N_34325,N_31376,N_30155);
nor U34326 (N_34326,N_30618,N_32385);
and U34327 (N_34327,N_31270,N_31973);
and U34328 (N_34328,N_30312,N_31568);
nand U34329 (N_34329,N_30433,N_31928);
nand U34330 (N_34330,N_30026,N_30209);
or U34331 (N_34331,N_30388,N_30560);
or U34332 (N_34332,N_31134,N_30773);
and U34333 (N_34333,N_30356,N_30391);
nand U34334 (N_34334,N_30937,N_30761);
or U34335 (N_34335,N_32209,N_32372);
nor U34336 (N_34336,N_30015,N_30663);
or U34337 (N_34337,N_32422,N_30258);
or U34338 (N_34338,N_30183,N_30198);
nor U34339 (N_34339,N_32438,N_30474);
nand U34340 (N_34340,N_30547,N_31509);
nor U34341 (N_34341,N_32392,N_32137);
xor U34342 (N_34342,N_31844,N_30521);
nor U34343 (N_34343,N_31743,N_30674);
or U34344 (N_34344,N_30713,N_32095);
or U34345 (N_34345,N_32324,N_31828);
and U34346 (N_34346,N_30478,N_31894);
nand U34347 (N_34347,N_31626,N_30937);
nor U34348 (N_34348,N_32148,N_30269);
nor U34349 (N_34349,N_30448,N_32170);
xor U34350 (N_34350,N_31155,N_30217);
and U34351 (N_34351,N_30248,N_30731);
nand U34352 (N_34352,N_31112,N_30768);
or U34353 (N_34353,N_32097,N_32012);
or U34354 (N_34354,N_31044,N_30298);
xor U34355 (N_34355,N_30408,N_30701);
and U34356 (N_34356,N_31368,N_30649);
xor U34357 (N_34357,N_31655,N_31121);
nor U34358 (N_34358,N_30068,N_31290);
nand U34359 (N_34359,N_31977,N_31993);
nor U34360 (N_34360,N_30695,N_31705);
xor U34361 (N_34361,N_31238,N_30454);
and U34362 (N_34362,N_30845,N_31930);
and U34363 (N_34363,N_31193,N_30338);
nor U34364 (N_34364,N_30786,N_30102);
nor U34365 (N_34365,N_31586,N_30511);
xnor U34366 (N_34366,N_31294,N_30123);
and U34367 (N_34367,N_31770,N_32333);
nor U34368 (N_34368,N_31681,N_31776);
nand U34369 (N_34369,N_30741,N_30857);
and U34370 (N_34370,N_30939,N_32087);
and U34371 (N_34371,N_32398,N_32254);
nand U34372 (N_34372,N_31563,N_30867);
or U34373 (N_34373,N_30949,N_32224);
nand U34374 (N_34374,N_32323,N_31647);
nand U34375 (N_34375,N_31923,N_30904);
xnor U34376 (N_34376,N_31199,N_30219);
and U34377 (N_34377,N_30024,N_31467);
or U34378 (N_34378,N_30284,N_31928);
nor U34379 (N_34379,N_30005,N_32294);
nand U34380 (N_34380,N_30773,N_31566);
nand U34381 (N_34381,N_30289,N_32312);
nor U34382 (N_34382,N_32097,N_30136);
or U34383 (N_34383,N_32000,N_31452);
nor U34384 (N_34384,N_30811,N_32101);
xnor U34385 (N_34385,N_30961,N_30905);
and U34386 (N_34386,N_31149,N_32299);
or U34387 (N_34387,N_32170,N_31653);
xor U34388 (N_34388,N_30156,N_30340);
or U34389 (N_34389,N_32019,N_30587);
xor U34390 (N_34390,N_30825,N_32202);
or U34391 (N_34391,N_30526,N_32335);
or U34392 (N_34392,N_31093,N_31205);
nor U34393 (N_34393,N_30203,N_30266);
nand U34394 (N_34394,N_31362,N_31270);
nand U34395 (N_34395,N_30348,N_31631);
nand U34396 (N_34396,N_30696,N_32046);
or U34397 (N_34397,N_30305,N_31812);
xor U34398 (N_34398,N_30446,N_30057);
xnor U34399 (N_34399,N_30269,N_30077);
xor U34400 (N_34400,N_31852,N_31608);
nor U34401 (N_34401,N_30774,N_31260);
xnor U34402 (N_34402,N_32033,N_31362);
nor U34403 (N_34403,N_30752,N_31399);
or U34404 (N_34404,N_31889,N_31409);
nand U34405 (N_34405,N_31831,N_30808);
or U34406 (N_34406,N_32205,N_30552);
xnor U34407 (N_34407,N_31316,N_32313);
nand U34408 (N_34408,N_32279,N_30738);
and U34409 (N_34409,N_30062,N_31650);
xnor U34410 (N_34410,N_30097,N_31842);
and U34411 (N_34411,N_31304,N_31714);
and U34412 (N_34412,N_30219,N_31998);
xnor U34413 (N_34413,N_31360,N_31733);
nor U34414 (N_34414,N_30144,N_32080);
nor U34415 (N_34415,N_31274,N_31909);
nor U34416 (N_34416,N_32185,N_32437);
nor U34417 (N_34417,N_31943,N_31326);
and U34418 (N_34418,N_30031,N_32299);
xor U34419 (N_34419,N_32402,N_31200);
nand U34420 (N_34420,N_30872,N_30438);
nand U34421 (N_34421,N_31633,N_30391);
nor U34422 (N_34422,N_32439,N_31359);
or U34423 (N_34423,N_31250,N_31076);
xnor U34424 (N_34424,N_30108,N_31692);
and U34425 (N_34425,N_31135,N_30889);
or U34426 (N_34426,N_31810,N_30293);
xnor U34427 (N_34427,N_30462,N_31845);
or U34428 (N_34428,N_32231,N_30888);
nor U34429 (N_34429,N_30645,N_32059);
nor U34430 (N_34430,N_30864,N_31536);
nand U34431 (N_34431,N_30386,N_31654);
nand U34432 (N_34432,N_30229,N_30446);
nand U34433 (N_34433,N_31547,N_30790);
xnor U34434 (N_34434,N_31937,N_31295);
nand U34435 (N_34435,N_30378,N_30363);
and U34436 (N_34436,N_31633,N_30813);
nor U34437 (N_34437,N_32170,N_30351);
nand U34438 (N_34438,N_30011,N_31011);
nor U34439 (N_34439,N_32197,N_30061);
nand U34440 (N_34440,N_30510,N_32158);
xor U34441 (N_34441,N_30371,N_31268);
and U34442 (N_34442,N_31131,N_31006);
or U34443 (N_34443,N_30647,N_30549);
nor U34444 (N_34444,N_32404,N_31770);
nand U34445 (N_34445,N_31788,N_30345);
nand U34446 (N_34446,N_30085,N_30996);
and U34447 (N_34447,N_31864,N_30816);
xnor U34448 (N_34448,N_31053,N_30830);
nand U34449 (N_34449,N_31746,N_31181);
nand U34450 (N_34450,N_30739,N_31483);
nand U34451 (N_34451,N_30648,N_32139);
nand U34452 (N_34452,N_30659,N_32187);
or U34453 (N_34453,N_31271,N_30039);
nand U34454 (N_34454,N_32098,N_31289);
nand U34455 (N_34455,N_30170,N_31585);
xor U34456 (N_34456,N_32277,N_31131);
nor U34457 (N_34457,N_30734,N_30977);
nor U34458 (N_34458,N_30170,N_30047);
nor U34459 (N_34459,N_31604,N_32403);
or U34460 (N_34460,N_31928,N_31636);
and U34461 (N_34461,N_31681,N_32398);
nor U34462 (N_34462,N_31992,N_32012);
nor U34463 (N_34463,N_30686,N_30765);
nor U34464 (N_34464,N_31124,N_31665);
and U34465 (N_34465,N_30917,N_30024);
nand U34466 (N_34466,N_32294,N_31744);
nor U34467 (N_34467,N_30233,N_30376);
and U34468 (N_34468,N_31654,N_32016);
nor U34469 (N_34469,N_31064,N_32300);
nand U34470 (N_34470,N_30408,N_30078);
nor U34471 (N_34471,N_30949,N_30610);
or U34472 (N_34472,N_30865,N_31769);
nor U34473 (N_34473,N_31517,N_31742);
or U34474 (N_34474,N_32177,N_31737);
or U34475 (N_34475,N_30237,N_30822);
xnor U34476 (N_34476,N_30997,N_32138);
or U34477 (N_34477,N_31250,N_31681);
xor U34478 (N_34478,N_30165,N_31859);
or U34479 (N_34479,N_31407,N_30945);
or U34480 (N_34480,N_31501,N_32146);
and U34481 (N_34481,N_31166,N_31955);
xor U34482 (N_34482,N_32161,N_30336);
nor U34483 (N_34483,N_30443,N_32335);
and U34484 (N_34484,N_32063,N_32391);
and U34485 (N_34485,N_31166,N_30123);
nand U34486 (N_34486,N_31504,N_31770);
nand U34487 (N_34487,N_32032,N_31251);
or U34488 (N_34488,N_31871,N_31424);
xnor U34489 (N_34489,N_31867,N_32205);
or U34490 (N_34490,N_31662,N_30117);
xor U34491 (N_34491,N_30577,N_30086);
nand U34492 (N_34492,N_31601,N_30588);
or U34493 (N_34493,N_31793,N_31448);
or U34494 (N_34494,N_31804,N_30793);
or U34495 (N_34495,N_32263,N_31863);
nand U34496 (N_34496,N_31249,N_31178);
nand U34497 (N_34497,N_31702,N_30446);
or U34498 (N_34498,N_32301,N_31502);
nor U34499 (N_34499,N_32109,N_30476);
nand U34500 (N_34500,N_30826,N_31532);
nor U34501 (N_34501,N_31505,N_30287);
xnor U34502 (N_34502,N_30310,N_30573);
and U34503 (N_34503,N_30706,N_30141);
nor U34504 (N_34504,N_30987,N_31351);
or U34505 (N_34505,N_31908,N_32099);
or U34506 (N_34506,N_31845,N_32257);
nor U34507 (N_34507,N_31362,N_31096);
nand U34508 (N_34508,N_30191,N_30658);
xor U34509 (N_34509,N_31717,N_30362);
nor U34510 (N_34510,N_31650,N_32194);
xnor U34511 (N_34511,N_32086,N_31151);
or U34512 (N_34512,N_31274,N_31012);
xnor U34513 (N_34513,N_32317,N_32314);
xnor U34514 (N_34514,N_32443,N_31649);
xnor U34515 (N_34515,N_30228,N_31366);
or U34516 (N_34516,N_32354,N_31485);
nand U34517 (N_34517,N_31828,N_32160);
nor U34518 (N_34518,N_30532,N_30768);
nor U34519 (N_34519,N_32462,N_30275);
nand U34520 (N_34520,N_30404,N_30328);
nor U34521 (N_34521,N_31427,N_31248);
nand U34522 (N_34522,N_30130,N_31703);
xor U34523 (N_34523,N_30839,N_32393);
or U34524 (N_34524,N_31263,N_32298);
xor U34525 (N_34525,N_30985,N_31789);
nand U34526 (N_34526,N_31716,N_31799);
or U34527 (N_34527,N_31281,N_32208);
xnor U34528 (N_34528,N_31709,N_31138);
nor U34529 (N_34529,N_30992,N_32275);
and U34530 (N_34530,N_30134,N_30321);
or U34531 (N_34531,N_31957,N_32225);
xor U34532 (N_34532,N_31743,N_30706);
nand U34533 (N_34533,N_32221,N_32383);
and U34534 (N_34534,N_30862,N_31872);
or U34535 (N_34535,N_31218,N_31331);
nor U34536 (N_34536,N_32161,N_30315);
and U34537 (N_34537,N_30163,N_30073);
or U34538 (N_34538,N_31517,N_31427);
xnor U34539 (N_34539,N_30645,N_30132);
xnor U34540 (N_34540,N_30625,N_30546);
and U34541 (N_34541,N_30525,N_31515);
nand U34542 (N_34542,N_31193,N_31588);
nor U34543 (N_34543,N_31958,N_31145);
nor U34544 (N_34544,N_30339,N_30575);
xor U34545 (N_34545,N_31473,N_30272);
nand U34546 (N_34546,N_31898,N_30786);
or U34547 (N_34547,N_30259,N_30386);
nor U34548 (N_34548,N_31596,N_30850);
or U34549 (N_34549,N_30381,N_31960);
nand U34550 (N_34550,N_30795,N_30280);
or U34551 (N_34551,N_31802,N_32316);
and U34552 (N_34552,N_31118,N_31759);
and U34553 (N_34553,N_31284,N_30150);
nor U34554 (N_34554,N_30827,N_30293);
nor U34555 (N_34555,N_30002,N_31864);
and U34556 (N_34556,N_30048,N_32106);
nand U34557 (N_34557,N_30817,N_30188);
xor U34558 (N_34558,N_30914,N_30230);
nand U34559 (N_34559,N_31500,N_30962);
nand U34560 (N_34560,N_31754,N_30478);
and U34561 (N_34561,N_30540,N_30652);
nand U34562 (N_34562,N_31856,N_32391);
nand U34563 (N_34563,N_31569,N_31343);
and U34564 (N_34564,N_32291,N_30691);
and U34565 (N_34565,N_30455,N_30818);
xnor U34566 (N_34566,N_31679,N_32227);
nand U34567 (N_34567,N_30608,N_30609);
nor U34568 (N_34568,N_31888,N_30787);
xor U34569 (N_34569,N_32252,N_30535);
and U34570 (N_34570,N_32140,N_32200);
xnor U34571 (N_34571,N_32374,N_30635);
xor U34572 (N_34572,N_31265,N_32127);
nand U34573 (N_34573,N_32237,N_31564);
or U34574 (N_34574,N_30701,N_30639);
or U34575 (N_34575,N_30421,N_32468);
nand U34576 (N_34576,N_31012,N_31652);
xor U34577 (N_34577,N_31083,N_31898);
xor U34578 (N_34578,N_31001,N_32104);
xnor U34579 (N_34579,N_31375,N_30380);
xor U34580 (N_34580,N_30620,N_31536);
xnor U34581 (N_34581,N_31744,N_31281);
and U34582 (N_34582,N_30270,N_31753);
or U34583 (N_34583,N_32428,N_31727);
and U34584 (N_34584,N_30141,N_32471);
or U34585 (N_34585,N_31403,N_30959);
and U34586 (N_34586,N_32400,N_30647);
nand U34587 (N_34587,N_31697,N_32162);
nand U34588 (N_34588,N_32331,N_30130);
and U34589 (N_34589,N_32363,N_31577);
xnor U34590 (N_34590,N_32180,N_30596);
or U34591 (N_34591,N_32141,N_30949);
or U34592 (N_34592,N_32032,N_30658);
xor U34593 (N_34593,N_32001,N_30322);
or U34594 (N_34594,N_30903,N_32472);
nand U34595 (N_34595,N_32240,N_31568);
xnor U34596 (N_34596,N_31259,N_31540);
or U34597 (N_34597,N_30502,N_32156);
xor U34598 (N_34598,N_31133,N_31285);
nor U34599 (N_34599,N_30990,N_30214);
and U34600 (N_34600,N_31016,N_31971);
nor U34601 (N_34601,N_31897,N_32270);
or U34602 (N_34602,N_30447,N_31998);
xor U34603 (N_34603,N_31603,N_30824);
or U34604 (N_34604,N_32108,N_31462);
nand U34605 (N_34605,N_32261,N_32216);
or U34606 (N_34606,N_31771,N_31734);
or U34607 (N_34607,N_32379,N_31557);
nor U34608 (N_34608,N_31321,N_31393);
xnor U34609 (N_34609,N_30695,N_31526);
nand U34610 (N_34610,N_30239,N_30690);
nor U34611 (N_34611,N_31413,N_31982);
nor U34612 (N_34612,N_32010,N_32097);
xnor U34613 (N_34613,N_31935,N_31285);
and U34614 (N_34614,N_31700,N_32450);
or U34615 (N_34615,N_30877,N_32114);
and U34616 (N_34616,N_31040,N_30696);
nor U34617 (N_34617,N_30948,N_30518);
and U34618 (N_34618,N_30132,N_31854);
nor U34619 (N_34619,N_31484,N_30446);
nand U34620 (N_34620,N_31804,N_31224);
and U34621 (N_34621,N_32490,N_32231);
nand U34622 (N_34622,N_31514,N_30378);
nand U34623 (N_34623,N_31169,N_31614);
or U34624 (N_34624,N_30788,N_31384);
nand U34625 (N_34625,N_32421,N_30863);
xor U34626 (N_34626,N_31285,N_31353);
nand U34627 (N_34627,N_31102,N_31370);
and U34628 (N_34628,N_30132,N_31956);
nor U34629 (N_34629,N_30175,N_30430);
nand U34630 (N_34630,N_31284,N_30033);
xor U34631 (N_34631,N_30699,N_30471);
xnor U34632 (N_34632,N_31668,N_31514);
xnor U34633 (N_34633,N_31024,N_32354);
xor U34634 (N_34634,N_30620,N_30416);
or U34635 (N_34635,N_31069,N_31648);
or U34636 (N_34636,N_30658,N_32330);
xnor U34637 (N_34637,N_31448,N_31579);
nor U34638 (N_34638,N_31067,N_31989);
and U34639 (N_34639,N_31515,N_31952);
nand U34640 (N_34640,N_32266,N_32447);
and U34641 (N_34641,N_30819,N_32307);
and U34642 (N_34642,N_31266,N_30630);
nand U34643 (N_34643,N_30998,N_30578);
and U34644 (N_34644,N_30955,N_30509);
xor U34645 (N_34645,N_32307,N_30191);
and U34646 (N_34646,N_31154,N_31912);
nor U34647 (N_34647,N_31986,N_31925);
xnor U34648 (N_34648,N_32361,N_31365);
nand U34649 (N_34649,N_32107,N_31605);
or U34650 (N_34650,N_31940,N_30145);
xnor U34651 (N_34651,N_31189,N_31422);
xor U34652 (N_34652,N_31772,N_30989);
or U34653 (N_34653,N_31572,N_30500);
or U34654 (N_34654,N_31802,N_30119);
or U34655 (N_34655,N_30378,N_31594);
or U34656 (N_34656,N_32087,N_31712);
nand U34657 (N_34657,N_31924,N_32228);
or U34658 (N_34658,N_32311,N_30522);
nor U34659 (N_34659,N_30072,N_32435);
and U34660 (N_34660,N_30165,N_30726);
or U34661 (N_34661,N_32019,N_30495);
nand U34662 (N_34662,N_32134,N_30826);
nand U34663 (N_34663,N_31381,N_31535);
nand U34664 (N_34664,N_31927,N_31838);
nand U34665 (N_34665,N_30478,N_30697);
nand U34666 (N_34666,N_32106,N_30274);
xnor U34667 (N_34667,N_31934,N_31622);
or U34668 (N_34668,N_32017,N_31446);
and U34669 (N_34669,N_30119,N_30480);
nand U34670 (N_34670,N_31235,N_32493);
nand U34671 (N_34671,N_31611,N_32141);
nand U34672 (N_34672,N_32058,N_31655);
or U34673 (N_34673,N_30929,N_32106);
or U34674 (N_34674,N_30674,N_30837);
or U34675 (N_34675,N_31122,N_30621);
and U34676 (N_34676,N_30310,N_30864);
and U34677 (N_34677,N_32400,N_31040);
xor U34678 (N_34678,N_30227,N_30134);
and U34679 (N_34679,N_30778,N_31365);
and U34680 (N_34680,N_31010,N_31263);
or U34681 (N_34681,N_30702,N_30415);
or U34682 (N_34682,N_31455,N_30475);
or U34683 (N_34683,N_31887,N_31395);
xor U34684 (N_34684,N_32040,N_30327);
xor U34685 (N_34685,N_30901,N_32330);
or U34686 (N_34686,N_30341,N_32242);
or U34687 (N_34687,N_32205,N_32444);
xor U34688 (N_34688,N_31599,N_31460);
nor U34689 (N_34689,N_32255,N_30938);
xor U34690 (N_34690,N_30514,N_32250);
nand U34691 (N_34691,N_30219,N_32341);
nand U34692 (N_34692,N_32170,N_30954);
and U34693 (N_34693,N_32410,N_30102);
and U34694 (N_34694,N_30484,N_31250);
or U34695 (N_34695,N_32417,N_31074);
xnor U34696 (N_34696,N_30057,N_32003);
and U34697 (N_34697,N_31922,N_31834);
nor U34698 (N_34698,N_31896,N_31620);
xor U34699 (N_34699,N_32387,N_31663);
or U34700 (N_34700,N_30053,N_32140);
xnor U34701 (N_34701,N_31308,N_30600);
and U34702 (N_34702,N_31340,N_30808);
nand U34703 (N_34703,N_32394,N_30353);
or U34704 (N_34704,N_30571,N_30351);
or U34705 (N_34705,N_31029,N_31902);
nor U34706 (N_34706,N_30211,N_31542);
and U34707 (N_34707,N_30940,N_32187);
nand U34708 (N_34708,N_30338,N_31742);
or U34709 (N_34709,N_32313,N_31882);
or U34710 (N_34710,N_30597,N_32170);
or U34711 (N_34711,N_31298,N_30908);
nor U34712 (N_34712,N_31843,N_31859);
or U34713 (N_34713,N_31705,N_32486);
nand U34714 (N_34714,N_32144,N_30101);
and U34715 (N_34715,N_32091,N_30786);
nor U34716 (N_34716,N_30901,N_31909);
or U34717 (N_34717,N_30910,N_30176);
or U34718 (N_34718,N_30667,N_32079);
or U34719 (N_34719,N_30694,N_30023);
nand U34720 (N_34720,N_31667,N_30281);
and U34721 (N_34721,N_30220,N_30460);
and U34722 (N_34722,N_30800,N_32284);
xor U34723 (N_34723,N_32359,N_32280);
nand U34724 (N_34724,N_31390,N_31280);
and U34725 (N_34725,N_30182,N_30336);
and U34726 (N_34726,N_30867,N_30834);
xnor U34727 (N_34727,N_31340,N_31062);
and U34728 (N_34728,N_31570,N_31390);
xor U34729 (N_34729,N_30415,N_30729);
nand U34730 (N_34730,N_32219,N_30821);
xor U34731 (N_34731,N_32332,N_31727);
or U34732 (N_34732,N_32420,N_32319);
or U34733 (N_34733,N_32001,N_32146);
nor U34734 (N_34734,N_30542,N_32440);
or U34735 (N_34735,N_30681,N_32043);
and U34736 (N_34736,N_30839,N_31042);
and U34737 (N_34737,N_31559,N_30736);
nor U34738 (N_34738,N_30441,N_30958);
or U34739 (N_34739,N_30069,N_31247);
nand U34740 (N_34740,N_31505,N_31882);
nand U34741 (N_34741,N_31880,N_30408);
xnor U34742 (N_34742,N_30663,N_31582);
nand U34743 (N_34743,N_31940,N_32229);
and U34744 (N_34744,N_30516,N_30848);
xnor U34745 (N_34745,N_30867,N_31287);
nand U34746 (N_34746,N_31966,N_30176);
and U34747 (N_34747,N_32480,N_32189);
or U34748 (N_34748,N_31963,N_30088);
or U34749 (N_34749,N_30274,N_31144);
nand U34750 (N_34750,N_30779,N_30545);
or U34751 (N_34751,N_30842,N_32198);
and U34752 (N_34752,N_31963,N_30223);
and U34753 (N_34753,N_31060,N_30523);
nor U34754 (N_34754,N_32476,N_31377);
and U34755 (N_34755,N_31711,N_30368);
and U34756 (N_34756,N_32479,N_30937);
xor U34757 (N_34757,N_31090,N_30085);
and U34758 (N_34758,N_30937,N_32430);
or U34759 (N_34759,N_31813,N_31482);
or U34760 (N_34760,N_31066,N_32203);
and U34761 (N_34761,N_32367,N_31866);
xor U34762 (N_34762,N_30054,N_32357);
nand U34763 (N_34763,N_31378,N_30692);
nor U34764 (N_34764,N_30238,N_30821);
xnor U34765 (N_34765,N_31592,N_30308);
xnor U34766 (N_34766,N_32127,N_32425);
or U34767 (N_34767,N_30598,N_30317);
nand U34768 (N_34768,N_30260,N_31766);
and U34769 (N_34769,N_32014,N_30676);
nor U34770 (N_34770,N_30676,N_31011);
and U34771 (N_34771,N_32060,N_30470);
nor U34772 (N_34772,N_31467,N_31641);
and U34773 (N_34773,N_31509,N_32405);
nand U34774 (N_34774,N_32366,N_30806);
or U34775 (N_34775,N_31271,N_30658);
and U34776 (N_34776,N_31841,N_32330);
xnor U34777 (N_34777,N_31829,N_31315);
xor U34778 (N_34778,N_31983,N_32241);
xor U34779 (N_34779,N_31453,N_32085);
and U34780 (N_34780,N_32401,N_30650);
xnor U34781 (N_34781,N_32164,N_30427);
nand U34782 (N_34782,N_31517,N_32173);
or U34783 (N_34783,N_31322,N_30522);
nor U34784 (N_34784,N_31295,N_32093);
nand U34785 (N_34785,N_31873,N_31089);
nand U34786 (N_34786,N_30975,N_31572);
or U34787 (N_34787,N_32396,N_30947);
nand U34788 (N_34788,N_30044,N_30441);
nand U34789 (N_34789,N_32455,N_30155);
nor U34790 (N_34790,N_31935,N_30012);
or U34791 (N_34791,N_30838,N_30007);
or U34792 (N_34792,N_31437,N_31579);
xor U34793 (N_34793,N_30151,N_31614);
and U34794 (N_34794,N_31616,N_30469);
nor U34795 (N_34795,N_30862,N_30986);
nand U34796 (N_34796,N_30369,N_31742);
xnor U34797 (N_34797,N_30664,N_31181);
or U34798 (N_34798,N_30208,N_31765);
or U34799 (N_34799,N_30140,N_31493);
and U34800 (N_34800,N_31638,N_30388);
nor U34801 (N_34801,N_30894,N_30022);
nor U34802 (N_34802,N_30044,N_31849);
nand U34803 (N_34803,N_32270,N_30418);
xor U34804 (N_34804,N_30788,N_30726);
or U34805 (N_34805,N_31490,N_31954);
nand U34806 (N_34806,N_30088,N_31998);
xnor U34807 (N_34807,N_30544,N_31270);
xor U34808 (N_34808,N_30741,N_30244);
or U34809 (N_34809,N_31137,N_31388);
xnor U34810 (N_34810,N_30704,N_30971);
xor U34811 (N_34811,N_30798,N_30533);
xnor U34812 (N_34812,N_31981,N_30039);
nand U34813 (N_34813,N_31854,N_30343);
and U34814 (N_34814,N_31329,N_30557);
nand U34815 (N_34815,N_31265,N_32177);
nor U34816 (N_34816,N_32091,N_30863);
xnor U34817 (N_34817,N_30213,N_31089);
xnor U34818 (N_34818,N_32179,N_32047);
and U34819 (N_34819,N_32211,N_31733);
and U34820 (N_34820,N_31617,N_30654);
and U34821 (N_34821,N_30977,N_30974);
nand U34822 (N_34822,N_31555,N_31926);
and U34823 (N_34823,N_30874,N_32453);
or U34824 (N_34824,N_30820,N_31699);
xnor U34825 (N_34825,N_30251,N_30279);
nor U34826 (N_34826,N_31258,N_30469);
or U34827 (N_34827,N_32398,N_30682);
or U34828 (N_34828,N_30871,N_31602);
or U34829 (N_34829,N_32039,N_30931);
or U34830 (N_34830,N_31235,N_31559);
xnor U34831 (N_34831,N_32412,N_30524);
xor U34832 (N_34832,N_31031,N_31738);
xor U34833 (N_34833,N_31301,N_32107);
nor U34834 (N_34834,N_31466,N_32356);
nand U34835 (N_34835,N_30309,N_32421);
and U34836 (N_34836,N_32019,N_31072);
or U34837 (N_34837,N_32252,N_32352);
nor U34838 (N_34838,N_31742,N_31437);
nor U34839 (N_34839,N_30398,N_30943);
or U34840 (N_34840,N_32135,N_30713);
and U34841 (N_34841,N_30646,N_31289);
or U34842 (N_34842,N_32109,N_31621);
xnor U34843 (N_34843,N_31164,N_30714);
nor U34844 (N_34844,N_30446,N_30893);
nor U34845 (N_34845,N_30683,N_30996);
nor U34846 (N_34846,N_31073,N_30687);
or U34847 (N_34847,N_30003,N_32270);
nand U34848 (N_34848,N_30876,N_30692);
or U34849 (N_34849,N_31304,N_30172);
nor U34850 (N_34850,N_32498,N_30686);
nor U34851 (N_34851,N_32230,N_30462);
xnor U34852 (N_34852,N_30484,N_31785);
xnor U34853 (N_34853,N_31482,N_32210);
nand U34854 (N_34854,N_31691,N_31760);
nand U34855 (N_34855,N_31271,N_30838);
xnor U34856 (N_34856,N_32250,N_30555);
and U34857 (N_34857,N_30293,N_31328);
nand U34858 (N_34858,N_31763,N_31202);
and U34859 (N_34859,N_30111,N_32082);
nand U34860 (N_34860,N_30643,N_32386);
or U34861 (N_34861,N_31557,N_31080);
nor U34862 (N_34862,N_30326,N_32331);
or U34863 (N_34863,N_30926,N_30467);
nand U34864 (N_34864,N_30259,N_30169);
or U34865 (N_34865,N_32268,N_31059);
nor U34866 (N_34866,N_32393,N_30377);
nand U34867 (N_34867,N_31949,N_31902);
nor U34868 (N_34868,N_32451,N_30382);
and U34869 (N_34869,N_32064,N_32353);
or U34870 (N_34870,N_31745,N_30433);
nor U34871 (N_34871,N_31958,N_31385);
nand U34872 (N_34872,N_30208,N_32400);
xnor U34873 (N_34873,N_31137,N_30064);
and U34874 (N_34874,N_31484,N_31358);
nor U34875 (N_34875,N_31749,N_30060);
nor U34876 (N_34876,N_31696,N_31485);
nand U34877 (N_34877,N_30795,N_32120);
or U34878 (N_34878,N_30184,N_30469);
nand U34879 (N_34879,N_31340,N_31408);
nand U34880 (N_34880,N_31739,N_31282);
xor U34881 (N_34881,N_32097,N_30722);
nor U34882 (N_34882,N_30238,N_31233);
nand U34883 (N_34883,N_31971,N_32496);
or U34884 (N_34884,N_30630,N_31211);
nor U34885 (N_34885,N_30876,N_31314);
nand U34886 (N_34886,N_31347,N_30835);
xor U34887 (N_34887,N_30801,N_30085);
xnor U34888 (N_34888,N_32342,N_30575);
nand U34889 (N_34889,N_31543,N_30431);
nor U34890 (N_34890,N_31656,N_32182);
and U34891 (N_34891,N_31137,N_31958);
xor U34892 (N_34892,N_31810,N_30528);
nor U34893 (N_34893,N_30209,N_30738);
xor U34894 (N_34894,N_30062,N_31026);
and U34895 (N_34895,N_30137,N_30054);
and U34896 (N_34896,N_30360,N_31091);
or U34897 (N_34897,N_30798,N_32356);
nor U34898 (N_34898,N_30920,N_31237);
or U34899 (N_34899,N_30926,N_31238);
nand U34900 (N_34900,N_30709,N_31144);
or U34901 (N_34901,N_31816,N_31928);
xnor U34902 (N_34902,N_30839,N_31417);
xor U34903 (N_34903,N_30320,N_31605);
or U34904 (N_34904,N_31970,N_30134);
nor U34905 (N_34905,N_32270,N_31601);
xor U34906 (N_34906,N_30532,N_30689);
nor U34907 (N_34907,N_30090,N_30880);
and U34908 (N_34908,N_32368,N_31552);
xor U34909 (N_34909,N_31646,N_31761);
xnor U34910 (N_34910,N_32177,N_31284);
or U34911 (N_34911,N_32090,N_30889);
nor U34912 (N_34912,N_31064,N_30155);
xor U34913 (N_34913,N_31654,N_32450);
xor U34914 (N_34914,N_30085,N_32376);
or U34915 (N_34915,N_31268,N_30199);
xor U34916 (N_34916,N_30341,N_32080);
or U34917 (N_34917,N_31131,N_30097);
or U34918 (N_34918,N_31603,N_32488);
nand U34919 (N_34919,N_30542,N_30363);
nand U34920 (N_34920,N_31643,N_32385);
nor U34921 (N_34921,N_31460,N_31639);
nor U34922 (N_34922,N_30143,N_32183);
or U34923 (N_34923,N_32303,N_30566);
or U34924 (N_34924,N_32384,N_30459);
nor U34925 (N_34925,N_31684,N_32087);
xnor U34926 (N_34926,N_31969,N_31934);
xor U34927 (N_34927,N_32167,N_30545);
xor U34928 (N_34928,N_30106,N_31562);
nor U34929 (N_34929,N_32388,N_31927);
or U34930 (N_34930,N_31325,N_32054);
nand U34931 (N_34931,N_30244,N_30730);
nand U34932 (N_34932,N_31210,N_30831);
xor U34933 (N_34933,N_30849,N_30455);
nor U34934 (N_34934,N_31530,N_32101);
and U34935 (N_34935,N_31991,N_31956);
or U34936 (N_34936,N_32209,N_31315);
and U34937 (N_34937,N_31822,N_31164);
and U34938 (N_34938,N_30282,N_30280);
and U34939 (N_34939,N_30181,N_31389);
xor U34940 (N_34940,N_30887,N_30145);
nor U34941 (N_34941,N_30854,N_31419);
xor U34942 (N_34942,N_30532,N_30731);
nand U34943 (N_34943,N_30765,N_30829);
nand U34944 (N_34944,N_30746,N_31607);
and U34945 (N_34945,N_31002,N_31282);
nand U34946 (N_34946,N_31470,N_31059);
or U34947 (N_34947,N_31401,N_31298);
nor U34948 (N_34948,N_31455,N_31092);
or U34949 (N_34949,N_32128,N_31306);
or U34950 (N_34950,N_31859,N_32261);
xor U34951 (N_34951,N_31963,N_31475);
nor U34952 (N_34952,N_31225,N_32343);
and U34953 (N_34953,N_30732,N_30573);
xor U34954 (N_34954,N_30240,N_31289);
or U34955 (N_34955,N_31151,N_32100);
xor U34956 (N_34956,N_31975,N_31364);
and U34957 (N_34957,N_30758,N_30262);
nand U34958 (N_34958,N_31085,N_30176);
nand U34959 (N_34959,N_30427,N_30341);
xnor U34960 (N_34960,N_30694,N_31306);
nand U34961 (N_34961,N_31388,N_32258);
nand U34962 (N_34962,N_31090,N_31055);
nor U34963 (N_34963,N_32432,N_31000);
nand U34964 (N_34964,N_30816,N_30826);
or U34965 (N_34965,N_32100,N_31872);
nor U34966 (N_34966,N_32007,N_31724);
and U34967 (N_34967,N_31961,N_32174);
xnor U34968 (N_34968,N_31516,N_32135);
or U34969 (N_34969,N_31897,N_31747);
or U34970 (N_34970,N_31952,N_31245);
nand U34971 (N_34971,N_30711,N_30318);
xor U34972 (N_34972,N_32386,N_30207);
or U34973 (N_34973,N_30019,N_32448);
nor U34974 (N_34974,N_31204,N_30953);
nor U34975 (N_34975,N_30894,N_32292);
nand U34976 (N_34976,N_30608,N_30836);
and U34977 (N_34977,N_31743,N_31337);
xor U34978 (N_34978,N_30467,N_32392);
and U34979 (N_34979,N_32094,N_30884);
or U34980 (N_34980,N_31238,N_31077);
or U34981 (N_34981,N_31812,N_31481);
nor U34982 (N_34982,N_30450,N_31186);
nor U34983 (N_34983,N_30663,N_30591);
or U34984 (N_34984,N_31641,N_31323);
xor U34985 (N_34985,N_32154,N_31825);
nor U34986 (N_34986,N_32081,N_31221);
and U34987 (N_34987,N_32389,N_30922);
or U34988 (N_34988,N_30802,N_30548);
and U34989 (N_34989,N_30570,N_32218);
or U34990 (N_34990,N_30388,N_31302);
nor U34991 (N_34991,N_32435,N_30677);
and U34992 (N_34992,N_31646,N_30732);
xnor U34993 (N_34993,N_31326,N_32272);
nand U34994 (N_34994,N_30902,N_31935);
nor U34995 (N_34995,N_31815,N_31668);
or U34996 (N_34996,N_31693,N_31428);
and U34997 (N_34997,N_30504,N_30023);
and U34998 (N_34998,N_32249,N_30597);
nand U34999 (N_34999,N_31190,N_32015);
nor U35000 (N_35000,N_34413,N_34015);
xnor U35001 (N_35001,N_33192,N_33287);
nand U35002 (N_35002,N_33428,N_32573);
xor U35003 (N_35003,N_32843,N_32702);
and U35004 (N_35004,N_32744,N_33383);
nor U35005 (N_35005,N_34180,N_33703);
nor U35006 (N_35006,N_33567,N_34840);
xor U35007 (N_35007,N_33381,N_32775);
or U35008 (N_35008,N_34438,N_34738);
nand U35009 (N_35009,N_33384,N_34035);
xor U35010 (N_35010,N_34251,N_34950);
nand U35011 (N_35011,N_33686,N_34873);
xor U35012 (N_35012,N_34502,N_33774);
xnor U35013 (N_35013,N_34646,N_33746);
nor U35014 (N_35014,N_33433,N_32788);
or U35015 (N_35015,N_34771,N_34929);
nor U35016 (N_35016,N_33575,N_33028);
or U35017 (N_35017,N_32664,N_34360);
or U35018 (N_35018,N_34190,N_34369);
and U35019 (N_35019,N_32567,N_34570);
or U35020 (N_35020,N_33256,N_33334);
nand U35021 (N_35021,N_34158,N_33582);
or U35022 (N_35022,N_32706,N_34162);
xor U35023 (N_35023,N_32692,N_32733);
xor U35024 (N_35024,N_32509,N_33505);
nand U35025 (N_35025,N_34666,N_33648);
xnor U35026 (N_35026,N_34444,N_33612);
xor U35027 (N_35027,N_34457,N_34240);
nand U35028 (N_35028,N_32891,N_34186);
xnor U35029 (N_35029,N_34089,N_32771);
and U35030 (N_35030,N_33682,N_33123);
or U35031 (N_35031,N_33613,N_34572);
or U35032 (N_35032,N_34878,N_32711);
or U35033 (N_35033,N_32847,N_34092);
xor U35034 (N_35034,N_32660,N_32605);
xor U35035 (N_35035,N_34478,N_34963);
nand U35036 (N_35036,N_34167,N_33517);
xor U35037 (N_35037,N_32751,N_34674);
and U35038 (N_35038,N_33219,N_34611);
nor U35039 (N_35039,N_32877,N_33659);
nor U35040 (N_35040,N_33463,N_34688);
nor U35041 (N_35041,N_34494,N_32624);
xnor U35042 (N_35042,N_34227,N_33741);
or U35043 (N_35043,N_33330,N_34285);
nor U35044 (N_35044,N_34200,N_34689);
nor U35045 (N_35045,N_33088,N_33536);
and U35046 (N_35046,N_32999,N_34782);
or U35047 (N_35047,N_33504,N_32661);
or U35048 (N_35048,N_34786,N_34397);
nand U35049 (N_35049,N_33489,N_34411);
nand U35050 (N_35050,N_32838,N_33526);
or U35051 (N_35051,N_34741,N_34034);
and U35052 (N_35052,N_34521,N_34318);
or U35053 (N_35053,N_34442,N_33943);
xnor U35054 (N_35054,N_32683,N_33206);
nand U35055 (N_35055,N_34728,N_33832);
nand U35056 (N_35056,N_34255,N_34192);
nand U35057 (N_35057,N_34850,N_34648);
nor U35058 (N_35058,N_32897,N_33209);
and U35059 (N_35059,N_33542,N_34422);
nor U35060 (N_35060,N_34077,N_32929);
nand U35061 (N_35061,N_33070,N_33953);
nor U35062 (N_35062,N_33581,N_32549);
xnor U35063 (N_35063,N_32742,N_32672);
or U35064 (N_35064,N_33040,N_33823);
xor U35065 (N_35065,N_33163,N_33728);
xnor U35066 (N_35066,N_34317,N_33451);
xnor U35067 (N_35067,N_34593,N_32625);
nand U35068 (N_35068,N_33814,N_33792);
nand U35069 (N_35069,N_33726,N_34351);
and U35070 (N_35070,N_34406,N_33286);
or U35071 (N_35071,N_34199,N_33835);
nand U35072 (N_35072,N_34960,N_32765);
nand U35073 (N_35073,N_34606,N_34374);
xnor U35074 (N_35074,N_34864,N_32682);
xnor U35075 (N_35075,N_33750,N_33912);
and U35076 (N_35076,N_34335,N_34994);
nand U35077 (N_35077,N_34636,N_34177);
xor U35078 (N_35078,N_32651,N_33377);
nand U35079 (N_35079,N_33159,N_34859);
or U35080 (N_35080,N_34942,N_33514);
and U35081 (N_35081,N_34826,N_32927);
and U35082 (N_35082,N_33509,N_33050);
nor U35083 (N_35083,N_34887,N_33365);
and U35084 (N_35084,N_34590,N_32812);
nor U35085 (N_35085,N_34133,N_34690);
nor U35086 (N_35086,N_34568,N_32968);
nor U35087 (N_35087,N_34815,N_32915);
xnor U35088 (N_35088,N_34145,N_33139);
xor U35089 (N_35089,N_33197,N_34254);
and U35090 (N_35090,N_34205,N_32959);
xor U35091 (N_35091,N_33699,N_33934);
and U35092 (N_35092,N_33162,N_34224);
nand U35093 (N_35093,N_32822,N_33815);
and U35094 (N_35094,N_33578,N_33017);
and U35095 (N_35095,N_34475,N_34604);
or U35096 (N_35096,N_34029,N_32878);
or U35097 (N_35097,N_34802,N_33600);
xnor U35098 (N_35098,N_33412,N_34160);
and U35099 (N_35099,N_34157,N_34597);
nand U35100 (N_35100,N_33191,N_33390);
nand U35101 (N_35101,N_33572,N_34903);
or U35102 (N_35102,N_33900,N_33472);
xnor U35103 (N_35103,N_32791,N_34843);
xnor U35104 (N_35104,N_34816,N_34839);
and U35105 (N_35105,N_32607,N_33506);
nor U35106 (N_35106,N_33965,N_34165);
nor U35107 (N_35107,N_33131,N_34373);
or U35108 (N_35108,N_34819,N_34538);
or U35109 (N_35109,N_33760,N_32678);
nor U35110 (N_35110,N_34852,N_32740);
nand U35111 (N_35111,N_34750,N_33976);
nand U35112 (N_35112,N_34524,N_32925);
and U35113 (N_35113,N_32533,N_33193);
xnor U35114 (N_35114,N_34833,N_32813);
and U35115 (N_35115,N_34600,N_34345);
and U35116 (N_35116,N_33982,N_33491);
and U35117 (N_35117,N_33094,N_33802);
or U35118 (N_35118,N_34584,N_32787);
and U35119 (N_35119,N_34389,N_32868);
and U35120 (N_35120,N_34947,N_34208);
nor U35121 (N_35121,N_34552,N_33336);
nor U35122 (N_35122,N_34172,N_33370);
or U35123 (N_35123,N_33173,N_33441);
nand U35124 (N_35124,N_32770,N_34731);
nor U35125 (N_35125,N_34599,N_34895);
nand U35126 (N_35126,N_32537,N_34032);
nand U35127 (N_35127,N_33752,N_33853);
nand U35128 (N_35128,N_33062,N_33317);
and U35129 (N_35129,N_33171,N_33335);
or U35130 (N_35130,N_34805,N_32979);
xnor U35131 (N_35131,N_33068,N_32919);
or U35132 (N_35132,N_32650,N_34737);
or U35133 (N_35133,N_34159,N_32809);
or U35134 (N_35134,N_33115,N_33252);
and U35135 (N_35135,N_33990,N_34187);
xnor U35136 (N_35136,N_33722,N_34112);
nand U35137 (N_35137,N_32715,N_34281);
xor U35138 (N_35138,N_32559,N_32568);
nor U35139 (N_35139,N_32907,N_34797);
xnor U35140 (N_35140,N_32534,N_34679);
nand U35141 (N_35141,N_34898,N_32645);
nand U35142 (N_35142,N_33886,N_33820);
xnor U35143 (N_35143,N_32947,N_33315);
nor U35144 (N_35144,N_34639,N_32539);
nand U35145 (N_35145,N_33438,N_34354);
and U35146 (N_35146,N_34264,N_34232);
xor U35147 (N_35147,N_33615,N_34848);
nor U35148 (N_35148,N_33693,N_34783);
nor U35149 (N_35149,N_34484,N_33431);
and U35150 (N_35150,N_34935,N_33907);
or U35151 (N_35151,N_33076,N_34104);
xor U35152 (N_35152,N_33011,N_32869);
or U35153 (N_35153,N_34103,N_34900);
xor U35154 (N_35154,N_34892,N_34508);
xnor U35155 (N_35155,N_33737,N_34291);
nor U35156 (N_35156,N_33803,N_34204);
and U35157 (N_35157,N_33380,N_34314);
xnor U35158 (N_35158,N_34651,N_33666);
nand U35159 (N_35159,N_34927,N_33409);
and U35160 (N_35160,N_33913,N_34641);
xor U35161 (N_35161,N_34206,N_33013);
xnor U35162 (N_35162,N_32728,N_33200);
or U35163 (N_35163,N_32934,N_34628);
nor U35164 (N_35164,N_34353,N_33168);
nand U35165 (N_35165,N_33065,N_33174);
nor U35166 (N_35166,N_34025,N_34820);
and U35167 (N_35167,N_33633,N_34121);
xnor U35168 (N_35168,N_34723,N_34732);
nor U35169 (N_35169,N_34916,N_33022);
xor U35170 (N_35170,N_32724,N_34429);
xor U35171 (N_35171,N_34634,N_34503);
and U35172 (N_35172,N_34409,N_34488);
nor U35173 (N_35173,N_33518,N_32604);
nand U35174 (N_35174,N_33884,N_34768);
nand U35175 (N_35175,N_34548,N_34976);
and U35176 (N_35176,N_34851,N_34398);
and U35177 (N_35177,N_34617,N_32701);
nand U35178 (N_35178,N_32950,N_33083);
or U35179 (N_35179,N_32611,N_33473);
nand U35180 (N_35180,N_34505,N_33754);
nand U35181 (N_35181,N_34876,N_33766);
and U35182 (N_35182,N_34226,N_33464);
nor U35183 (N_35183,N_33704,N_33753);
xnor U35184 (N_35184,N_33324,N_33730);
and U35185 (N_35185,N_34368,N_32961);
or U35186 (N_35186,N_33051,N_32511);
nand U35187 (N_35187,N_33403,N_34303);
or U35188 (N_35188,N_32970,N_33558);
nand U35189 (N_35189,N_32516,N_34622);
nand U35190 (N_35190,N_32512,N_32839);
xnor U35191 (N_35191,N_34523,N_34662);
xnor U35192 (N_35192,N_34827,N_33087);
and U35193 (N_35193,N_34594,N_33149);
xor U35194 (N_35194,N_34344,N_33471);
xnor U35195 (N_35195,N_32563,N_33425);
xnor U35196 (N_35196,N_34233,N_33397);
and U35197 (N_35197,N_33478,N_34930);
nor U35198 (N_35198,N_32905,N_32506);
nor U35199 (N_35199,N_33119,N_34069);
nor U35200 (N_35200,N_34392,N_33074);
and U35201 (N_35201,N_32797,N_32668);
and U35202 (N_35202,N_33822,N_33981);
xnor U35203 (N_35203,N_34941,N_34076);
or U35204 (N_35204,N_32597,N_33475);
nand U35205 (N_35205,N_34117,N_32881);
or U35206 (N_35206,N_33672,N_33875);
or U35207 (N_35207,N_34765,N_33890);
xnor U35208 (N_35208,N_32756,N_33885);
or U35209 (N_35209,N_32858,N_34294);
nand U35210 (N_35210,N_34323,N_33207);
xor U35211 (N_35211,N_32519,N_34440);
xor U35212 (N_35212,N_33711,N_33418);
nor U35213 (N_35213,N_34030,N_32807);
or U35214 (N_35214,N_33539,N_32767);
nor U35215 (N_35215,N_33522,N_33279);
nand U35216 (N_35216,N_33235,N_34865);
nor U35217 (N_35217,N_33282,N_34914);
or U35218 (N_35218,N_34838,N_32599);
xnor U35219 (N_35219,N_34435,N_32933);
nand U35220 (N_35220,N_34962,N_33781);
xnor U35221 (N_35221,N_34907,N_33707);
nand U35222 (N_35222,N_33511,N_33114);
or U35223 (N_35223,N_34616,N_32614);
nor U35224 (N_35224,N_33257,N_32619);
nor U35225 (N_35225,N_33854,N_32758);
nor U35226 (N_35226,N_34319,N_33574);
nand U35227 (N_35227,N_33097,N_33332);
nor U35228 (N_35228,N_34722,N_33300);
or U35229 (N_35229,N_32956,N_33643);
xnor U35230 (N_35230,N_34210,N_34658);
nand U35231 (N_35231,N_34870,N_33841);
nand U35232 (N_35232,N_33614,N_34042);
xor U35233 (N_35233,N_34271,N_34410);
and U35234 (N_35234,N_33399,N_34202);
and U35235 (N_35235,N_34924,N_34216);
and U35236 (N_35236,N_33762,N_32875);
xnor U35237 (N_35237,N_34633,N_32923);
and U35238 (N_35238,N_33455,N_34266);
xnor U35239 (N_35239,N_34586,N_34498);
or U35240 (N_35240,N_32971,N_32783);
nand U35241 (N_35241,N_34074,N_33535);
nor U35242 (N_35242,N_33789,N_34591);
and U35243 (N_35243,N_32593,N_32883);
or U35244 (N_35244,N_33341,N_33601);
nor U35245 (N_35245,N_32964,N_34010);
xnor U35246 (N_35246,N_33165,N_34296);
and U35247 (N_35247,N_32940,N_34746);
nor U35248 (N_35248,N_34241,N_33422);
xor U35249 (N_35249,N_33790,N_33673);
nor U35250 (N_35250,N_33230,N_32543);
or U35251 (N_35251,N_34657,N_34124);
and U35252 (N_35252,N_34279,N_34808);
nand U35253 (N_35253,N_32538,N_34632);
xnor U35254 (N_35254,N_32569,N_32653);
or U35255 (N_35255,N_33047,N_33795);
and U35256 (N_35256,N_34247,N_33113);
xnor U35257 (N_35257,N_34532,N_34028);
xor U35258 (N_35258,N_33107,N_32816);
or U35259 (N_35259,N_33253,N_34024);
or U35260 (N_35260,N_33079,N_32978);
nor U35261 (N_35261,N_33530,N_32551);
nand U35262 (N_35262,N_32768,N_32866);
nor U35263 (N_35263,N_32743,N_34683);
or U35264 (N_35264,N_33836,N_34515);
xor U35265 (N_35265,N_33343,N_33089);
nor U35266 (N_35266,N_33329,N_34088);
and U35267 (N_35267,N_34618,N_34706);
or U35268 (N_35268,N_32552,N_33634);
and U35269 (N_35269,N_34763,N_32703);
or U35270 (N_35270,N_32530,N_33347);
and U35271 (N_35271,N_34402,N_33597);
nand U35272 (N_35272,N_33880,N_34635);
or U35273 (N_35273,N_33043,N_34361);
nand U35274 (N_35274,N_33321,N_34978);
xnor U35275 (N_35275,N_34672,N_33735);
nand U35276 (N_35276,N_34522,N_33671);
or U35277 (N_35277,N_33571,N_34828);
nand U35278 (N_35278,N_33521,N_34896);
xor U35279 (N_35279,N_33291,N_32795);
and U35280 (N_35280,N_34416,N_33891);
and U35281 (N_35281,N_33210,N_34625);
or U35282 (N_35282,N_34357,N_34301);
nand U35283 (N_35283,N_34268,N_32566);
nor U35284 (N_35284,N_32828,N_32615);
xnor U35285 (N_35285,N_34671,N_33631);
or U35286 (N_35286,N_33767,N_32747);
and U35287 (N_35287,N_34339,N_32688);
nand U35288 (N_35288,N_34989,N_34809);
or U35289 (N_35289,N_33967,N_34749);
or U35290 (N_35290,N_32911,N_34968);
and U35291 (N_35291,N_33893,N_33363);
nor U35292 (N_35292,N_33450,N_34821);
or U35293 (N_35293,N_33541,N_34631);
and U35294 (N_35294,N_33482,N_33679);
xor U35295 (N_35295,N_34031,N_34100);
xor U35296 (N_35296,N_33411,N_32671);
nor U35297 (N_35297,N_33142,N_33918);
xnor U35298 (N_35298,N_33716,N_32790);
or U35299 (N_35299,N_33010,N_34445);
xor U35300 (N_35300,N_34744,N_33125);
xnor U35301 (N_35301,N_33779,N_33894);
nand U35302 (N_35302,N_34707,N_33724);
nor U35303 (N_35303,N_32799,N_33467);
and U35304 (N_35304,N_33816,N_33801);
nor U35305 (N_35305,N_34918,N_34175);
xnor U35306 (N_35306,N_34877,N_33167);
nor U35307 (N_35307,N_34324,N_34882);
and U35308 (N_35308,N_34879,N_33798);
nand U35309 (N_35309,N_32677,N_34904);
xnor U35310 (N_35310,N_33231,N_34955);
and U35311 (N_35311,N_34243,N_33607);
nor U35312 (N_35312,N_33494,N_32762);
xnor U35313 (N_35313,N_33030,N_34770);
or U35314 (N_35314,N_33793,N_32718);
or U35315 (N_35315,N_33280,N_33935);
nand U35316 (N_35316,N_33447,N_34626);
and U35317 (N_35317,N_34428,N_33346);
nand U35318 (N_35318,N_33307,N_33661);
and U35319 (N_35319,N_34193,N_34005);
nor U35320 (N_35320,N_32515,N_32752);
nand U35321 (N_35321,N_32704,N_33362);
or U35322 (N_35322,N_33999,N_33106);
xnor U35323 (N_35323,N_34242,N_33553);
nor U35324 (N_35324,N_33326,N_33049);
nor U35325 (N_35325,N_33860,N_34529);
or U35326 (N_35326,N_33547,N_33453);
or U35327 (N_35327,N_33850,N_33638);
nand U35328 (N_35328,N_34979,N_34881);
xnor U35329 (N_35329,N_32895,N_34725);
xor U35330 (N_35330,N_34761,N_33290);
or U35331 (N_35331,N_34367,N_34188);
xnor U35332 (N_35332,N_33462,N_33963);
or U35333 (N_35333,N_32909,N_33695);
and U35334 (N_35334,N_34995,N_32836);
and U35335 (N_35335,N_34181,N_32990);
xor U35336 (N_35336,N_33402,N_34712);
nor U35337 (N_35337,N_33085,N_33419);
nand U35338 (N_35338,N_32835,N_34695);
nor U35339 (N_35339,N_34585,N_34541);
xnor U35340 (N_35340,N_34099,N_32522);
or U35341 (N_35341,N_33421,N_34098);
and U35342 (N_35342,N_33285,N_33947);
nor U35343 (N_35343,N_34772,N_33617);
or U35344 (N_35344,N_32556,N_34485);
nand U35345 (N_35345,N_34670,N_32606);
xnor U35346 (N_35346,N_32801,N_33372);
xor U35347 (N_35347,N_33406,N_34817);
nor U35348 (N_35348,N_34939,N_34982);
nand U35349 (N_35349,N_33873,N_34474);
xnor U35350 (N_35350,N_33899,N_34311);
nor U35351 (N_35351,N_34510,N_34215);
or U35352 (N_35352,N_34476,N_33364);
nand U35353 (N_35353,N_33158,N_33871);
and U35354 (N_35354,N_34461,N_33887);
xor U35355 (N_35355,N_34156,N_33620);
or U35356 (N_35356,N_33348,N_32738);
xor U35357 (N_35357,N_33528,N_32746);
nand U35358 (N_35358,N_33925,N_34249);
xor U35359 (N_35359,N_33996,N_34171);
and U35360 (N_35360,N_33869,N_34053);
xor U35361 (N_35361,N_33588,N_34387);
nand U35362 (N_35362,N_33249,N_34039);
or U35363 (N_35363,N_32943,N_33124);
xnor U35364 (N_35364,N_33797,N_32705);
or U35365 (N_35365,N_33901,N_34987);
xor U35366 (N_35366,N_32641,N_34528);
nor U35367 (N_35367,N_34872,N_32827);
nand U35368 (N_35368,N_34447,N_32582);
xor U35369 (N_35369,N_34275,N_33296);
xnor U35370 (N_35370,N_34282,N_33442);
xor U35371 (N_35371,N_33828,N_33497);
nand U35372 (N_35372,N_34298,N_34184);
and U35373 (N_35373,N_33217,N_33974);
xnor U35374 (N_35374,N_33810,N_34909);
xor U35375 (N_35375,N_33141,N_34095);
and U35376 (N_35376,N_32644,N_34248);
or U35377 (N_35377,N_32532,N_33989);
and U35378 (N_35378,N_32680,N_33992);
nand U35379 (N_35379,N_34997,N_34891);
nand U35380 (N_35380,N_33112,N_33202);
and U35381 (N_35381,N_32572,N_34302);
or U35382 (N_35382,N_34483,N_33400);
nor U35383 (N_35383,N_33432,N_32504);
or U35384 (N_35384,N_33586,N_34363);
nand U35385 (N_35385,N_32983,N_32842);
or U35386 (N_35386,N_32576,N_34013);
and U35387 (N_35387,N_32864,N_34463);
or U35388 (N_35388,N_34954,N_33960);
and U35389 (N_35389,N_33519,N_34705);
or U35390 (N_35390,N_32779,N_33705);
nor U35391 (N_35391,N_34992,N_34455);
and U35392 (N_35392,N_32565,N_34320);
nor U35393 (N_35393,N_34814,N_34862);
nor U35394 (N_35394,N_32712,N_32854);
and U35395 (N_35395,N_33394,N_34587);
and U35396 (N_35396,N_34333,N_33486);
nand U35397 (N_35397,N_33345,N_34304);
nor U35398 (N_35398,N_33069,N_34277);
or U35399 (N_35399,N_34493,N_33375);
and U35400 (N_35400,N_34033,N_33513);
xnor U35401 (N_35401,N_33240,N_34056);
and U35402 (N_35402,N_34734,N_34576);
or U35403 (N_35403,N_33983,N_33410);
nand U35404 (N_35404,N_33557,N_32517);
or U35405 (N_35405,N_32963,N_33032);
xnor U35406 (N_35406,N_33635,N_34348);
and U35407 (N_35407,N_32698,N_33739);
xor U35408 (N_35408,N_33005,N_34085);
and U35409 (N_35409,N_32991,N_34431);
or U35410 (N_35410,N_34423,N_33978);
xor U35411 (N_35411,N_32789,N_33580);
and U35412 (N_35412,N_34691,N_34589);
nand U35413 (N_35413,N_32764,N_33759);
xor U35414 (N_35414,N_33713,N_34880);
nand U35415 (N_35415,N_34757,N_33292);
nor U35416 (N_35416,N_33204,N_34161);
xnor U35417 (N_35417,N_32695,N_33930);
xor U35418 (N_35418,N_34472,N_32817);
xor U35419 (N_35419,N_34141,N_33026);
xor U35420 (N_35420,N_34462,N_32785);
nor U35421 (N_35421,N_32908,N_34933);
nor U35422 (N_35422,N_33593,N_34906);
and U35423 (N_35423,N_33527,N_33243);
xor U35424 (N_35424,N_34886,N_32753);
xor U35425 (N_35425,N_34059,N_33474);
nor U35426 (N_35426,N_33104,N_32887);
nand U35427 (N_35427,N_33009,N_32670);
or U35428 (N_35428,N_33311,N_34113);
and U35429 (N_35429,N_34944,N_33826);
and U35430 (N_35430,N_33904,N_34974);
and U35431 (N_35431,N_34412,N_33689);
nor U35432 (N_35432,N_32687,N_33830);
and U35433 (N_35433,N_34120,N_32571);
and U35434 (N_35434,N_34810,N_32500);
and U35435 (N_35435,N_33995,N_33772);
nand U35436 (N_35436,N_32561,N_34926);
nor U35437 (N_35437,N_32721,N_32811);
and U35438 (N_35438,N_32541,N_32823);
nor U35439 (N_35439,N_33426,N_34458);
or U35440 (N_35440,N_33595,N_33962);
nor U35441 (N_35441,N_33512,N_34060);
xor U35442 (N_35442,N_32898,N_34676);
xor U35443 (N_35443,N_32837,N_33376);
nand U35444 (N_35444,N_34747,N_34684);
nor U35445 (N_35445,N_33281,N_32725);
nand U35446 (N_35446,N_33652,N_32629);
nor U35447 (N_35447,N_33997,N_34364);
xor U35448 (N_35448,N_34779,N_32806);
and U35449 (N_35449,N_33696,N_34479);
and U35450 (N_35450,N_34014,N_34456);
or U35451 (N_35451,N_33415,N_33570);
nand U35452 (N_35452,N_33986,N_33610);
nor U35453 (N_35453,N_34306,N_33653);
nand U35454 (N_35454,N_34996,N_32932);
or U35455 (N_35455,N_32726,N_34603);
nand U35456 (N_35456,N_33550,N_34525);
xor U35457 (N_35457,N_34182,N_34842);
nand U35458 (N_35458,N_34911,N_33117);
nand U35459 (N_35459,N_34650,N_34340);
and U35460 (N_35460,N_32739,N_34535);
nor U35461 (N_35461,N_34118,N_33812);
nor U35462 (N_35462,N_34550,N_33259);
or U35463 (N_35463,N_34739,N_33312);
or U35464 (N_35464,N_32655,N_34931);
nand U35465 (N_35465,N_33319,N_34564);
nor U35466 (N_35466,N_34129,N_33023);
or U35467 (N_35467,N_33868,N_32904);
or U35468 (N_35468,N_33338,N_32942);
xnor U35469 (N_35469,N_32863,N_34228);
nor U35470 (N_35470,N_34756,N_32639);
and U35471 (N_35471,N_33765,N_33761);
xor U35472 (N_35472,N_32860,N_33045);
nand U35473 (N_35473,N_32656,N_34096);
nand U35474 (N_35474,N_33014,N_33544);
and U35475 (N_35475,N_32562,N_33157);
xnor U35476 (N_35476,N_33968,N_34107);
or U35477 (N_35477,N_34875,N_34901);
xor U35478 (N_35478,N_33680,N_33337);
xnor U35479 (N_35479,N_32781,N_33297);
nor U35480 (N_35480,N_33318,N_33706);
xor U35481 (N_35481,N_32935,N_33264);
or U35482 (N_35482,N_32918,N_33121);
and U35483 (N_35483,N_33743,N_32696);
xnor U35484 (N_35484,N_33237,N_33000);
nor U35485 (N_35485,N_33299,N_34414);
nand U35486 (N_35486,N_33920,N_33002);
xnor U35487 (N_35487,N_34534,N_34231);
and U35488 (N_35488,N_33092,N_34822);
nor U35489 (N_35489,N_32575,N_33529);
nand U35490 (N_35490,N_32989,N_33261);
or U35491 (N_35491,N_34693,N_32689);
and U35492 (N_35492,N_33099,N_34908);
nor U35493 (N_35493,N_33749,N_33993);
nor U35494 (N_35494,N_34915,N_33222);
and U35495 (N_35495,N_32826,N_33940);
nand U35496 (N_35496,N_33800,N_33538);
and U35497 (N_35497,N_34799,N_34115);
nor U35498 (N_35498,N_33923,N_33740);
nand U35499 (N_35499,N_33223,N_32857);
and U35500 (N_35500,N_32774,N_32745);
xnor U35501 (N_35501,N_33405,N_34384);
or U35502 (N_35502,N_34583,N_34936);
nand U35503 (N_35503,N_33681,N_34713);
xor U35504 (N_35504,N_32901,N_33301);
and U35505 (N_35505,N_32507,N_34379);
or U35506 (N_35506,N_33188,N_34561);
xor U35507 (N_35507,N_32798,N_33452);
xnor U35508 (N_35508,N_34919,N_34209);
and U35509 (N_35509,N_33609,N_32634);
xor U35510 (N_35510,N_34619,N_33146);
xnor U35511 (N_35511,N_32525,N_32518);
or U35512 (N_35512,N_34446,N_34263);
nor U35513 (N_35513,N_34714,N_33359);
nor U35514 (N_35514,N_33817,N_32546);
xor U35515 (N_35515,N_34064,N_33339);
or U35516 (N_35516,N_32585,N_34147);
or U35517 (N_35517,N_34405,N_33393);
and U35518 (N_35518,N_32930,N_34970);
and U35519 (N_35519,N_33477,N_34582);
or U35520 (N_35520,N_33936,N_34511);
or U35521 (N_35521,N_32876,N_32600);
xnor U35522 (N_35522,N_33247,N_32647);
and U35523 (N_35523,N_33360,N_33031);
and U35524 (N_35524,N_32808,N_34201);
nand U35525 (N_35525,N_33952,N_32865);
nand U35526 (N_35526,N_33388,N_34555);
or U35527 (N_35527,N_33769,N_33971);
and U35528 (N_35528,N_32859,N_32954);
or U35529 (N_35529,N_33733,N_34623);
xor U35530 (N_35530,N_34090,N_32952);
nand U35531 (N_35531,N_32755,N_34054);
nand U35532 (N_35532,N_32595,N_33226);
or U35533 (N_35533,N_32955,N_32621);
and U35534 (N_35534,N_33443,N_33314);
nand U35535 (N_35535,N_33594,N_32840);
nor U35536 (N_35536,N_33694,N_32759);
and U35537 (N_35537,N_33932,N_33824);
xnor U35538 (N_35538,N_34126,N_32662);
nand U35539 (N_35539,N_33794,N_32853);
nor U35540 (N_35540,N_33623,N_34718);
nor U35541 (N_35541,N_32862,N_33020);
and U35542 (N_35542,N_32659,N_34017);
xnor U35543 (N_35543,N_33732,N_34894);
and U35544 (N_35544,N_32945,N_33502);
xnor U35545 (N_35545,N_34250,N_34058);
nor U35546 (N_35546,N_34454,N_34751);
nand U35547 (N_35547,N_34038,N_33136);
nor U35548 (N_35548,N_34940,N_33184);
xor U35549 (N_35549,N_32949,N_33498);
nor U35550 (N_35550,N_34467,N_34365);
xnor U35551 (N_35551,N_32986,N_34801);
nor U35552 (N_35552,N_33130,N_34261);
or U35553 (N_35553,N_33183,N_34366);
nor U35554 (N_35554,N_32777,N_34910);
and U35555 (N_35555,N_33632,N_33355);
xnor U35556 (N_35556,N_34448,N_34834);
xnor U35557 (N_35557,N_33840,N_32592);
xor U35558 (N_35558,N_33549,N_33533);
nor U35559 (N_35559,N_33254,N_33621);
nor U35560 (N_35560,N_33651,N_33039);
or U35561 (N_35561,N_34154,N_34602);
xor U35562 (N_35562,N_33246,N_34536);
or U35563 (N_35563,N_34581,N_33306);
xnor U35564 (N_35564,N_32966,N_33273);
or U35565 (N_35565,N_33407,N_34660);
and U35566 (N_35566,N_34343,N_33236);
and U35567 (N_35567,N_32699,N_33954);
or U35568 (N_35568,N_33562,N_33021);
nand U35569 (N_35569,N_34197,N_33379);
xor U35570 (N_35570,N_34355,N_32845);
and U35571 (N_35571,N_33717,N_34152);
nand U35572 (N_35572,N_34500,N_32727);
nand U35573 (N_35573,N_32617,N_33991);
or U35574 (N_35574,N_34854,N_33082);
nand U35575 (N_35575,N_34824,N_34871);
nor U35576 (N_35576,N_33848,N_34596);
nor U35577 (N_35577,N_33701,N_34238);
or U35578 (N_35578,N_33662,N_33232);
nand U35579 (N_35579,N_33676,N_34762);
xnor U35580 (N_35580,N_33250,N_34899);
nor U35581 (N_35581,N_34800,N_33133);
nand U35582 (N_35582,N_33166,N_34776);
and U35583 (N_35583,N_34811,N_33148);
nor U35584 (N_35584,N_33373,N_34421);
nand U35585 (N_35585,N_33628,N_34399);
nand U35586 (N_35586,N_33955,N_34173);
and U35587 (N_35587,N_32818,N_32608);
and U35588 (N_35588,N_34452,N_34027);
xor U35589 (N_35589,N_33589,N_34745);
and U35590 (N_35590,N_34544,N_34174);
and U35591 (N_35591,N_33602,N_33215);
or U35592 (N_35592,N_34191,N_33646);
nor U35593 (N_35593,N_32649,N_32975);
nand U35594 (N_35594,N_32834,N_34084);
xor U35595 (N_35595,N_34066,N_33413);
xor U35596 (N_35596,N_33857,N_32673);
or U35597 (N_35597,N_34804,N_34164);
or U35598 (N_35598,N_32548,N_33941);
nand U35599 (N_35599,N_34217,N_34313);
nor U35600 (N_35600,N_34307,N_33867);
xor U35601 (N_35601,N_34563,N_33169);
nor U35602 (N_35602,N_32748,N_33046);
nor U35603 (N_35603,N_32628,N_32633);
or U35604 (N_35604,N_33378,N_34425);
and U35605 (N_35605,N_34818,N_33460);
xnor U35606 (N_35606,N_33127,N_32957);
nand U35607 (N_35607,N_32814,N_34499);
nor U35608 (N_35608,N_33189,N_33642);
or U35609 (N_35609,N_33599,N_33175);
nand U35610 (N_35610,N_34956,N_33270);
xnor U35611 (N_35611,N_34439,N_33034);
or U35612 (N_35612,N_32937,N_34308);
nand U35613 (N_35613,N_32717,N_33924);
nor U35614 (N_35614,N_32846,N_33973);
and U35615 (N_35615,N_32754,N_32855);
nor U35616 (N_35616,N_33787,N_33103);
and U35617 (N_35617,N_33523,N_32830);
or U35618 (N_35618,N_34567,N_34105);
nor U35619 (N_35619,N_34885,N_33029);
or U35620 (N_35620,N_33071,N_33342);
nand U35621 (N_35621,N_33956,N_34137);
xor U35622 (N_35622,N_34132,N_34130);
or U35623 (N_35623,N_33844,N_34959);
nor U35624 (N_35624,N_34272,N_32529);
nor U35625 (N_35625,N_34777,N_33327);
nand U35626 (N_35626,N_34984,N_33266);
xnor U35627 (N_35627,N_33663,N_32654);
nor U35628 (N_35628,N_33683,N_34265);
and U35629 (N_35629,N_34067,N_33155);
xor U35630 (N_35630,N_34858,N_33495);
or U35631 (N_35631,N_33537,N_34957);
or U35632 (N_35632,N_33898,N_33485);
or U35633 (N_35633,N_34322,N_34637);
and U35634 (N_35634,N_33786,N_34653);
nand U35635 (N_35635,N_32773,N_33416);
nor U35636 (N_35636,N_34223,N_32555);
nor U35637 (N_35637,N_34464,N_33849);
xor U35638 (N_35638,N_34775,N_34965);
nor U35639 (N_35639,N_32708,N_33058);
and U35640 (N_35640,N_34860,N_33878);
or U35641 (N_35641,N_33843,N_33889);
or U35642 (N_35642,N_33771,N_33751);
xnor U35643 (N_35643,N_34539,N_32610);
nor U35644 (N_35644,N_34480,N_32741);
and U35645 (N_35645,N_34449,N_33056);
xnor U35646 (N_35646,N_33272,N_33882);
or U35647 (N_35647,N_32697,N_33468);
nand U35648 (N_35648,N_32900,N_32716);
nor U35649 (N_35649,N_32803,N_33172);
and U35650 (N_35650,N_33922,N_33906);
or U35651 (N_35651,N_34287,N_33063);
xnor U35652 (N_35652,N_32831,N_33933);
or U35653 (N_35653,N_32872,N_34041);
xnor U35654 (N_35654,N_34486,N_34050);
or U35655 (N_35655,N_33488,N_34792);
nor U35656 (N_35656,N_33208,N_33715);
xnor U35657 (N_35657,N_34108,N_34116);
nand U35658 (N_35658,N_34884,N_33105);
and U35659 (N_35659,N_33870,N_34830);
or U35660 (N_35660,N_32734,N_33540);
or U35661 (N_35661,N_34286,N_33592);
nor U35662 (N_35662,N_33964,N_32665);
and U35663 (N_35663,N_34640,N_33697);
and U35664 (N_35664,N_32760,N_34327);
or U35665 (N_35665,N_34897,N_33080);
xor U35666 (N_35666,N_33012,N_32579);
or U35667 (N_35667,N_34315,N_34235);
nand U35668 (N_35668,N_33729,N_33685);
nor U35669 (N_35669,N_34481,N_33805);
xor U35670 (N_35670,N_34218,N_34767);
or U35671 (N_35671,N_34780,N_32545);
nand U35672 (N_35672,N_32987,N_32523);
and U35673 (N_35673,N_33234,N_32992);
or U35674 (N_35674,N_34393,N_33645);
or U35675 (N_35675,N_33825,N_33367);
nor U35676 (N_35676,N_32993,N_34813);
nand U35677 (N_35677,N_32676,N_33077);
or U35678 (N_35678,N_32769,N_34459);
nand U35679 (N_35679,N_34540,N_34874);
nand U35680 (N_35680,N_34134,N_33692);
nor U35681 (N_35681,N_32685,N_34404);
nand U35682 (N_35682,N_32632,N_32736);
xnor U35683 (N_35683,N_33624,N_34546);
nand U35684 (N_35684,N_32542,N_34111);
nor U35685 (N_35685,N_34349,N_34299);
nor U35686 (N_35686,N_33454,N_33349);
and U35687 (N_35687,N_33470,N_33093);
nand U35688 (N_35688,N_34716,N_33420);
or U35689 (N_35689,N_33356,N_33756);
nand U35690 (N_35690,N_34677,N_34473);
xnor U35691 (N_35691,N_32849,N_33161);
or U35692 (N_35692,N_32888,N_34434);
nor U35693 (N_35693,N_33298,N_32974);
nand U35694 (N_35694,N_33323,N_33690);
nand U35695 (N_35695,N_33994,N_32591);
nor U35696 (N_35696,N_33160,N_34065);
and U35697 (N_35697,N_32707,N_32889);
nor U35698 (N_35698,N_32861,N_33078);
nand U35699 (N_35699,N_33361,N_33640);
nand U35700 (N_35700,N_32792,N_33879);
nand U35701 (N_35701,N_33584,N_32782);
xor U35702 (N_35702,N_32946,N_33783);
and U35703 (N_35703,N_32879,N_34040);
nor U35704 (N_35704,N_34520,N_34295);
or U35705 (N_35705,N_34003,N_34560);
nor U35706 (N_35706,N_33914,N_33320);
and U35707 (N_35707,N_34964,N_34694);
or U35708 (N_35708,N_32960,N_32630);
xnor U35709 (N_35709,N_34889,N_33604);
or U35710 (N_35710,N_33218,N_33401);
xnor U35711 (N_35711,N_33702,N_33354);
nand U35712 (N_35712,N_34234,N_34743);
and U35713 (N_35713,N_33806,N_33132);
and U35714 (N_35714,N_33305,N_34844);
nand U35715 (N_35715,N_33603,N_34966);
nand U35716 (N_35716,N_34110,N_33972);
xnor U35717 (N_35717,N_34213,N_34849);
xor U35718 (N_35718,N_33185,N_33688);
nor U35719 (N_35719,N_34985,N_34071);
xor U35720 (N_35720,N_34341,N_34006);
nor U35721 (N_35721,N_32570,N_32962);
nand U35722 (N_35722,N_32588,N_32681);
nand U35723 (N_35723,N_32557,N_34280);
xor U35724 (N_35724,N_33241,N_34530);
and U35725 (N_35725,N_34607,N_32635);
and U35726 (N_35726,N_34605,N_33302);
nor U35727 (N_35727,N_34812,N_32719);
nand U35728 (N_35728,N_33808,N_33548);
nand U35729 (N_35729,N_33874,N_33821);
and U35730 (N_35730,N_34644,N_33700);
nand U35731 (N_35731,N_34740,N_33778);
and U35732 (N_35732,N_34183,N_33182);
or U35733 (N_35733,N_34832,N_33501);
or U35734 (N_35734,N_34578,N_32574);
nor U35735 (N_35735,N_32980,N_34922);
and U35736 (N_35736,N_34609,N_33579);
or U35737 (N_35737,N_32731,N_34736);
nand U35738 (N_35738,N_34932,N_32514);
nand U35739 (N_35739,N_34668,N_34754);
xnor U35740 (N_35740,N_33268,N_33201);
xor U35741 (N_35741,N_32602,N_34328);
or U35742 (N_35742,N_33516,N_32936);
and U35743 (N_35743,N_32772,N_32581);
nor U35744 (N_35744,N_34624,N_34052);
and U35745 (N_35745,N_33834,N_33408);
nor U35746 (N_35746,N_34386,N_33654);
xnor U35747 (N_35747,N_34545,N_32941);
or U35748 (N_35748,N_32713,N_33500);
nand U35749 (N_35749,N_32603,N_33608);
and U35750 (N_35750,N_34492,N_32833);
xnor U35751 (N_35751,N_33015,N_33274);
and U35752 (N_35752,N_33545,N_33229);
xnor U35753 (N_35753,N_33892,N_34509);
nand U35754 (N_35754,N_33476,N_32917);
or U35755 (N_35755,N_32691,N_34973);
xnor U35756 (N_35756,N_34021,N_34575);
or U35757 (N_35757,N_34504,N_32526);
nand U35758 (N_35758,N_34149,N_33525);
xnor U35759 (N_35759,N_33664,N_34420);
xnor U35760 (N_35760,N_33929,N_32666);
nand U35761 (N_35761,N_33902,N_33531);
nand U35762 (N_35762,N_33984,N_33773);
and U35763 (N_35763,N_33469,N_33507);
nor U35764 (N_35764,N_33669,N_33980);
xor U35765 (N_35765,N_34140,N_34890);
nor U35766 (N_35766,N_34061,N_33444);
nand U35767 (N_35767,N_34011,N_33086);
nand U35768 (N_35768,N_34288,N_34912);
or U35769 (N_35769,N_33658,N_34697);
and U35770 (N_35770,N_32931,N_34856);
xor U35771 (N_35771,N_34592,N_34758);
or U35772 (N_35772,N_34793,N_34857);
nand U35773 (N_35773,N_34195,N_34443);
nor U35774 (N_35774,N_32969,N_34647);
nand U35775 (N_35775,N_34554,N_33090);
and U35776 (N_35776,N_33807,N_32657);
nand U35777 (N_35777,N_33944,N_33775);
nand U35778 (N_35778,N_32669,N_32903);
nor U35779 (N_35779,N_34562,N_34376);
xor U35780 (N_35780,N_33275,N_33975);
and U35781 (N_35781,N_32675,N_33650);
or U35782 (N_35782,N_33691,N_33839);
and U35783 (N_35783,N_34664,N_33255);
nand U35784 (N_35784,N_34861,N_33573);
nor U35785 (N_35785,N_32819,N_34836);
nand U35786 (N_35786,N_32684,N_34101);
xor U35787 (N_35787,N_34390,N_34283);
xor U35788 (N_35788,N_32609,N_33979);
nor U35789 (N_35789,N_33190,N_33289);
or U35790 (N_35790,N_34533,N_34823);
nor U35791 (N_35791,N_33687,N_34598);
nand U35792 (N_35792,N_33727,N_34222);
nand U35793 (N_35793,N_32750,N_34846);
or U35794 (N_35794,N_33449,N_34612);
nand U35795 (N_35795,N_34331,N_34685);
nor U35796 (N_35796,N_34359,N_33881);
nand U35797 (N_35797,N_32892,N_33636);
and U35798 (N_35798,N_33785,N_34490);
or U35799 (N_35799,N_34142,N_32587);
or U35800 (N_35800,N_33561,N_34669);
xnor U35801 (N_35801,N_33440,N_33138);
nor U35802 (N_35802,N_34652,N_34869);
nor U35803 (N_35803,N_33177,N_34178);
nor U35804 (N_35804,N_33288,N_32914);
nor U35805 (N_35805,N_33862,N_32553);
or U35806 (N_35806,N_34293,N_33156);
xor U35807 (N_35807,N_34007,N_32578);
or U35808 (N_35808,N_33404,N_33606);
or U35809 (N_35809,N_34981,N_33265);
nor U35810 (N_35810,N_32679,N_34951);
xnor U35811 (N_35811,N_32874,N_34385);
xnor U35812 (N_35812,N_33044,N_34358);
xnor U35813 (N_35813,N_33747,N_34841);
nand U35814 (N_35814,N_33829,N_32910);
nand U35815 (N_35815,N_34225,N_33458);
nand U35816 (N_35816,N_34773,N_34913);
nor U35817 (N_35817,N_34465,N_33035);
or U35818 (N_35818,N_33027,N_32916);
nor U35819 (N_35819,N_33919,N_34253);
and U35820 (N_35820,N_32531,N_32722);
and U35821 (N_35821,N_34046,N_34292);
or U35822 (N_35822,N_33263,N_33322);
nand U35823 (N_35823,N_34553,N_32524);
nand U35824 (N_35824,N_34125,N_32805);
xor U35825 (N_35825,N_34752,N_33777);
or U35826 (N_35826,N_32658,N_33721);
or U35827 (N_35827,N_34043,N_34729);
nand U35828 (N_35828,N_34934,N_33417);
xor U35829 (N_35829,N_34023,N_32510);
nor U35830 (N_35830,N_33811,N_34441);
or U35831 (N_35831,N_33392,N_33271);
xor U35832 (N_35832,N_33796,N_33134);
xnor U35833 (N_35833,N_34866,N_34321);
or U35834 (N_35834,N_33629,N_34630);
or U35835 (N_35835,N_34256,N_33396);
nor U35836 (N_35836,N_34902,N_33718);
or U35837 (N_35837,N_33493,N_34656);
and U35838 (N_35838,N_32997,N_33024);
nand U35839 (N_35839,N_34556,N_34642);
or U35840 (N_35840,N_34131,N_32926);
nor U35841 (N_35841,N_34008,N_33780);
nand U35842 (N_35842,N_33916,N_34537);
or U35843 (N_35843,N_32844,N_33655);
and U35844 (N_35844,N_34727,N_34391);
nor U35845 (N_35845,N_34297,N_34923);
and U35846 (N_35846,N_34407,N_34274);
or U35847 (N_35847,N_32778,N_33436);
or U35848 (N_35848,N_33556,N_33846);
and U35849 (N_35849,N_34724,N_32564);
xnor U35850 (N_35850,N_34094,N_34655);
and U35851 (N_35851,N_34329,N_33496);
nand U35852 (N_35852,N_33120,N_34127);
nor U35853 (N_35853,N_33888,N_33284);
or U35854 (N_35854,N_33391,N_33374);
nor U35855 (N_35855,N_33310,N_34595);
or U35856 (N_35856,N_32505,N_34748);
or U35857 (N_35857,N_34284,N_33926);
and U35858 (N_35858,N_33126,N_33251);
xnor U35859 (N_35859,N_32508,N_33709);
nand U35860 (N_35860,N_33667,N_33845);
nor U35861 (N_35861,N_33483,N_33554);
nor U35862 (N_35862,N_34087,N_34417);
xor U35863 (N_35863,N_33742,N_32601);
nor U35864 (N_35864,N_34300,N_33019);
nand U35865 (N_35865,N_34070,N_32924);
nand U35866 (N_35866,N_33059,N_32794);
and U35867 (N_35867,N_33861,N_34527);
or U35868 (N_35868,N_33187,N_34495);
nor U35869 (N_35869,N_33038,N_33770);
and U35870 (N_35870,N_34980,N_32667);
and U35871 (N_35871,N_34721,N_32996);
nor U35872 (N_35872,N_33684,N_33057);
xnor U35873 (N_35873,N_33109,N_34109);
xor U35874 (N_35874,N_33948,N_33938);
nor U35875 (N_35875,N_32535,N_34948);
nor U35876 (N_35876,N_33366,N_33351);
nor U35877 (N_35877,N_34114,N_32620);
nor U35878 (N_35878,N_33961,N_32583);
xor U35879 (N_35879,N_34432,N_33855);
nand U35880 (N_35880,N_33164,N_32815);
and U35881 (N_35881,N_32824,N_34863);
xnor U35882 (N_35882,N_32953,N_33583);
and U35883 (N_35883,N_34571,N_34615);
xnor U35884 (N_35884,N_34289,N_33576);
xor U35885 (N_35885,N_33937,N_33480);
nor U35886 (N_35886,N_34189,N_33283);
or U35887 (N_35887,N_34993,N_34513);
and U35888 (N_35888,N_32648,N_33102);
nand U35889 (N_35889,N_34806,N_34667);
xor U35890 (N_35890,N_34557,N_34733);
nand U35891 (N_35891,N_32735,N_34062);
and U35892 (N_35892,N_34988,N_32577);
and U35893 (N_35893,N_34853,N_33001);
or U35894 (N_35894,N_33145,N_34151);
xor U35895 (N_35895,N_33837,N_34336);
xnor U35896 (N_35896,N_34424,N_33791);
nand U35897 (N_35897,N_33052,N_32749);
xor U35898 (N_35898,N_33205,N_33856);
nor U35899 (N_35899,N_34419,N_34091);
xor U35900 (N_35900,N_34991,N_33096);
nand U35901 (N_35901,N_32544,N_32985);
nand U35902 (N_35902,N_33446,N_32821);
nand U35903 (N_35903,N_34794,N_32594);
and U35904 (N_35904,N_33768,N_34259);
nand U35905 (N_35905,N_33212,N_33764);
nand U35906 (N_35906,N_32800,N_32694);
and U35907 (N_35907,N_32693,N_32804);
or U35908 (N_35908,N_33897,N_34649);
xor U35909 (N_35909,N_33585,N_32967);
nor U35910 (N_35910,N_34661,N_33515);
or U35911 (N_35911,N_34798,N_33448);
nor U35912 (N_35912,N_34645,N_33144);
or U35913 (N_35913,N_34717,N_33042);
and U35914 (N_35914,N_34588,N_34700);
nor U35915 (N_35915,N_33859,N_33872);
nor U35916 (N_35916,N_34057,N_33435);
nor U35917 (N_35917,N_32912,N_34781);
xnor U35918 (N_35918,N_33921,N_33262);
and U35919 (N_35919,N_33194,N_33465);
xor U35920 (N_35920,N_32802,N_34487);
xnor U35921 (N_35921,N_33176,N_32981);
or U35922 (N_35922,N_32732,N_33799);
nand U35923 (N_35923,N_34049,N_32984);
nand U35924 (N_35924,N_34829,N_32793);
nand U35925 (N_35925,N_32638,N_33945);
nor U35926 (N_35926,N_34305,N_32554);
and U35927 (N_35927,N_32627,N_34969);
nand U35928 (N_35928,N_34803,N_32973);
or U35929 (N_35929,N_33075,N_32870);
and U35930 (N_35930,N_33876,N_33260);
xor U35931 (N_35931,N_33784,N_34497);
and U35932 (N_35932,N_32939,N_34044);
nand U35933 (N_35933,N_33387,N_33931);
nor U35934 (N_35934,N_34791,N_32766);
nand U35935 (N_35935,N_34083,N_34045);
xnor U35936 (N_35936,N_33487,N_34477);
xor U35937 (N_35937,N_34000,N_33137);
xor U35938 (N_35938,N_33213,N_33637);
and U35939 (N_35939,N_32720,N_33758);
xor U35940 (N_35940,N_33095,N_32623);
xor U35941 (N_35941,N_33211,N_34496);
nor U35942 (N_35942,N_32893,N_34453);
xor U35943 (N_35943,N_32580,N_32832);
nand U35944 (N_35944,N_33357,N_33081);
nand U35945 (N_35945,N_33293,N_32714);
nand U35946 (N_35946,N_33178,N_33877);
nor U35947 (N_35947,N_34290,N_34971);
nor U35948 (N_35948,N_33866,N_34551);
and U35949 (N_35949,N_33564,N_32730);
nand U35950 (N_35950,N_34138,N_33675);
xor U35951 (N_35951,N_32965,N_34395);
nor U35952 (N_35952,N_34018,N_32613);
or U35953 (N_35953,N_33018,N_34144);
or U35954 (N_35954,N_33647,N_34380);
nand U35955 (N_35955,N_33227,N_34945);
and U35956 (N_35956,N_34312,N_32502);
and U35957 (N_35957,N_34450,N_34569);
nand U35958 (N_35958,N_34468,N_33143);
xor U35959 (N_35959,N_33532,N_32848);
and U35960 (N_35960,N_34401,N_34920);
nand U35961 (N_35961,N_34316,N_33569);
or U35962 (N_35962,N_33195,N_32622);
or U35963 (N_35963,N_34698,N_33568);
nor U35964 (N_35964,N_33847,N_34047);
and U35965 (N_35965,N_32616,N_34375);
and U35966 (N_35966,N_34451,N_34784);
or U35967 (N_35967,N_33755,N_32536);
nand U35968 (N_35968,N_34681,N_34847);
or U35969 (N_35969,N_33382,N_33559);
nand U35970 (N_35970,N_33959,N_33563);
nand U35971 (N_35971,N_32906,N_34489);
or U35972 (N_35972,N_32873,N_34760);
xnor U35973 (N_35973,N_32642,N_32896);
or U35974 (N_35974,N_33170,N_32618);
xnor U35975 (N_35975,N_32710,N_34139);
nor U35976 (N_35976,N_33278,N_34078);
nor U35977 (N_35977,N_34252,N_32958);
xor U35978 (N_35978,N_34938,N_34245);
nor U35979 (N_35979,N_34097,N_34119);
xnor U35980 (N_35980,N_33988,N_34659);
xnor U35981 (N_35981,N_33644,N_34501);
or U35982 (N_35982,N_33016,N_34135);
xor U35983 (N_35983,N_34418,N_34378);
nand U35984 (N_35984,N_34565,N_34888);
nand U35985 (N_35985,N_34470,N_32643);
and U35986 (N_35986,N_33551,N_34123);
or U35987 (N_35987,N_34682,N_33116);
xor U35988 (N_35988,N_33055,N_34143);
xnor U35989 (N_35989,N_34460,N_33248);
nand U35990 (N_35990,N_33061,N_33831);
and U35991 (N_35991,N_33098,N_34169);
xnor U35992 (N_35992,N_34350,N_33084);
and U35993 (N_35993,N_33757,N_32729);
nand U35994 (N_35994,N_34531,N_34807);
or U35995 (N_35995,N_34709,N_34789);
nor U35996 (N_35996,N_33484,N_33358);
and U35997 (N_35997,N_33591,N_32784);
xnor U35998 (N_35998,N_34371,N_33951);
nand U35999 (N_35999,N_34638,N_33949);
xnor U36000 (N_36000,N_34026,N_33998);
nor U36001 (N_36001,N_32652,N_34766);
or U36002 (N_36002,N_34211,N_33674);
and U36003 (N_36003,N_32674,N_33276);
nor U36004 (N_36004,N_32646,N_34517);
xor U36005 (N_36005,N_34102,N_34063);
nor U36006 (N_36006,N_33368,N_33605);
nor U36007 (N_36007,N_33838,N_34426);
and U36008 (N_36008,N_33025,N_33386);
nor U36009 (N_36009,N_33776,N_34958);
xnor U36010 (N_36010,N_33782,N_34774);
and U36011 (N_36011,N_33657,N_34610);
or U36012 (N_36012,N_33064,N_33427);
or U36013 (N_36013,N_33128,N_34437);
or U36014 (N_36014,N_33966,N_33369);
nor U36015 (N_36015,N_34837,N_34383);
xnor U36016 (N_36016,N_32709,N_34905);
and U36017 (N_36017,N_34687,N_33153);
nor U36018 (N_36018,N_33313,N_34702);
xor U36019 (N_36019,N_32558,N_34704);
or U36020 (N_36020,N_32938,N_34020);
nand U36021 (N_36021,N_32513,N_32856);
nand U36022 (N_36022,N_33985,N_33911);
and U36023 (N_36023,N_34967,N_34710);
or U36024 (N_36024,N_34608,N_34022);
nor U36025 (N_36025,N_33224,N_33225);
and U36026 (N_36026,N_32686,N_33915);
nor U36027 (N_36027,N_33596,N_33895);
xor U36028 (N_36028,N_33625,N_34278);
nand U36029 (N_36029,N_33445,N_33238);
xnor U36030 (N_36030,N_32598,N_34382);
nor U36031 (N_36031,N_33316,N_33503);
nor U36032 (N_36032,N_34867,N_34148);
xnor U36033 (N_36033,N_32810,N_33073);
nand U36034 (N_36034,N_34983,N_33245);
or U36035 (N_36035,N_34080,N_34198);
nand U36036 (N_36036,N_32637,N_33091);
and U36037 (N_36037,N_33723,N_33350);
nand U36038 (N_36038,N_34491,N_34986);
or U36039 (N_36039,N_33389,N_34999);
and U36040 (N_36040,N_33340,N_33294);
xor U36041 (N_36041,N_34427,N_33883);
and U36042 (N_36042,N_32982,N_32851);
and U36043 (N_36043,N_34961,N_33543);
nor U36044 (N_36044,N_32995,N_34019);
and U36045 (N_36045,N_32944,N_34436);
nor U36046 (N_36046,N_34893,N_34037);
xor U36047 (N_36047,N_32547,N_32763);
or U36048 (N_36048,N_34128,N_34176);
nor U36049 (N_36049,N_33946,N_34953);
xnor U36050 (N_36050,N_34566,N_34673);
and U36051 (N_36051,N_34309,N_34790);
nand U36052 (N_36052,N_34072,N_33668);
nor U36053 (N_36053,N_33457,N_33140);
and U36054 (N_36054,N_32972,N_34258);
nor U36055 (N_36055,N_34237,N_32776);
and U36056 (N_36056,N_33395,N_32612);
or U36057 (N_36057,N_34925,N_34170);
xnor U36058 (N_36058,N_34230,N_34482);
xor U36059 (N_36059,N_33748,N_33216);
xor U36060 (N_36060,N_34787,N_33977);
xor U36061 (N_36061,N_33714,N_32882);
or U36062 (N_36062,N_33371,N_33744);
nor U36063 (N_36063,N_34514,N_32560);
xnor U36064 (N_36064,N_32884,N_33698);
and U36065 (N_36065,N_34835,N_34764);
or U36066 (N_36066,N_33048,N_33180);
nand U36067 (N_36067,N_33053,N_34506);
xnor U36068 (N_36068,N_34408,N_33398);
and U36069 (N_36069,N_33186,N_33004);
or U36070 (N_36070,N_34512,N_33566);
xor U36071 (N_36071,N_32899,N_34627);
and U36072 (N_36072,N_33414,N_33560);
nor U36073 (N_36073,N_33199,N_33423);
nand U36074 (N_36074,N_34726,N_33852);
xnor U36075 (N_36075,N_34620,N_32586);
nor U36076 (N_36076,N_33524,N_33950);
xor U36077 (N_36077,N_34356,N_34778);
nor U36078 (N_36078,N_34785,N_34269);
and U36079 (N_36079,N_34203,N_34207);
nor U36080 (N_36080,N_34943,N_34883);
and U36081 (N_36081,N_34370,N_33198);
nand U36082 (N_36082,N_33490,N_34212);
or U36083 (N_36083,N_34507,N_33851);
and U36084 (N_36084,N_33033,N_34769);
xor U36085 (N_36085,N_33827,N_33534);
or U36086 (N_36086,N_34753,N_33510);
nor U36087 (N_36087,N_32921,N_33864);
nor U36088 (N_36088,N_34262,N_32786);
or U36089 (N_36089,N_34543,N_34260);
nor U36090 (N_36090,N_33430,N_32521);
nor U36091 (N_36091,N_32780,N_33269);
and U36092 (N_36092,N_32871,N_34081);
nand U36093 (N_36093,N_34155,N_32590);
nand U36094 (N_36094,N_32596,N_33110);
nor U36095 (N_36095,N_34244,N_33616);
or U36096 (N_36096,N_32920,N_33066);
nor U36097 (N_36097,N_34276,N_32852);
xnor U36098 (N_36098,N_34573,N_33958);
and U36099 (N_36099,N_34221,N_32948);
or U36100 (N_36100,N_34730,N_33712);
nor U36101 (N_36101,N_33969,N_33908);
or U36102 (N_36102,N_34004,N_34665);
nand U36103 (N_36103,N_33036,N_34310);
nor U36104 (N_36104,N_34400,N_33060);
or U36105 (N_36105,N_34788,N_33720);
or U36106 (N_36106,N_33719,N_34246);
and U36107 (N_36107,N_34715,N_32994);
nand U36108 (N_36108,N_33303,N_32829);
xnor U36109 (N_36109,N_32503,N_33809);
nor U36110 (N_36110,N_34239,N_33150);
nand U36111 (N_36111,N_34675,N_34179);
nor U36112 (N_36112,N_34559,N_33818);
nor U36113 (N_36113,N_34577,N_32902);
nor U36114 (N_36114,N_33008,N_34580);
xor U36115 (N_36115,N_33865,N_32589);
and U36116 (N_36116,N_33546,N_34621);
or U36117 (N_36117,N_34082,N_34921);
or U36118 (N_36118,N_33037,N_34601);
nand U36119 (N_36119,N_34036,N_33508);
nor U36120 (N_36120,N_33333,N_34701);
nor U36121 (N_36121,N_33957,N_33736);
nand U36122 (N_36122,N_33308,N_33677);
and U36123 (N_36123,N_34720,N_33154);
or U36124 (N_36124,N_34009,N_33481);
nor U36125 (N_36125,N_34377,N_33003);
nor U36126 (N_36126,N_33928,N_34796);
xor U36127 (N_36127,N_33221,N_32663);
xnor U36128 (N_36128,N_32977,N_33492);
nand U36129 (N_36129,N_33429,N_32850);
nor U36130 (N_36130,N_33804,N_34696);
or U36131 (N_36131,N_34719,N_34093);
nand U36132 (N_36132,N_34150,N_34519);
and U36133 (N_36133,N_34270,N_34236);
or U36134 (N_36134,N_34680,N_34654);
or U36135 (N_36135,N_33041,N_34347);
nor U36136 (N_36136,N_34998,N_34326);
nand U36137 (N_36137,N_34547,N_34825);
and U36138 (N_36138,N_34708,N_33896);
or U36139 (N_36139,N_32631,N_34220);
nand U36140 (N_36140,N_34337,N_33656);
nor U36141 (N_36141,N_33466,N_33731);
xor U36142 (N_36142,N_32928,N_34430);
nor U36143 (N_36143,N_34558,N_34342);
and U36144 (N_36144,N_34122,N_34433);
xnor U36145 (N_36145,N_34526,N_34928);
nand U36146 (N_36146,N_33054,N_34831);
or U36147 (N_36147,N_33220,N_34711);
nand U36148 (N_36148,N_34346,N_34975);
nand U36149 (N_36149,N_33678,N_32867);
nor U36150 (N_36150,N_34012,N_32998);
and U36151 (N_36151,N_34855,N_32640);
xnor U36152 (N_36152,N_33917,N_33842);
or U36153 (N_36153,N_32886,N_34002);
xnor U36154 (N_36154,N_34613,N_33072);
xnor U36155 (N_36155,N_33277,N_34471);
xnor U36156 (N_36156,N_34229,N_33111);
xor U36157 (N_36157,N_34977,N_34372);
and U36158 (N_36158,N_33179,N_33331);
and U36159 (N_36159,N_33665,N_33734);
nand U36160 (N_36160,N_33788,N_33618);
nor U36161 (N_36161,N_34153,N_34629);
and U36162 (N_36162,N_34466,N_32501);
and U36163 (N_36163,N_34579,N_32796);
xnor U36164 (N_36164,N_33987,N_33708);
nand U36165 (N_36165,N_33763,N_32757);
or U36166 (N_36166,N_34868,N_34196);
or U36167 (N_36167,N_33108,N_33590);
xnor U36168 (N_36168,N_32540,N_34267);
nand U36169 (N_36169,N_33927,N_33813);
nand U36170 (N_36170,N_34086,N_33577);
nand U36171 (N_36171,N_34168,N_34330);
or U36172 (N_36172,N_33233,N_34735);
nor U36173 (N_36173,N_34338,N_34663);
xnor U36174 (N_36174,N_33152,N_34946);
and U36175 (N_36175,N_33456,N_34396);
and U36176 (N_36176,N_33833,N_34678);
nand U36177 (N_36177,N_34549,N_32520);
nor U36178 (N_36178,N_34972,N_33598);
or U36179 (N_36179,N_33639,N_34759);
nand U36180 (N_36180,N_33738,N_33181);
nor U36181 (N_36181,N_34388,N_33006);
nand U36182 (N_36182,N_33479,N_33304);
xnor U36183 (N_36183,N_33649,N_33641);
nor U36184 (N_36184,N_33499,N_33101);
nand U36185 (N_36185,N_34643,N_34106);
xor U36186 (N_36186,N_33863,N_34469);
and U36187 (N_36187,N_32988,N_32723);
nor U36188 (N_36188,N_33325,N_33611);
nor U36189 (N_36189,N_32880,N_32737);
nand U36190 (N_36190,N_34394,N_34742);
xor U36191 (N_36191,N_32527,N_32690);
nor U36192 (N_36192,N_33203,N_33122);
and U36193 (N_36193,N_34990,N_34686);
and U36194 (N_36194,N_32761,N_33565);
nand U36195 (N_36195,N_33352,N_34185);
or U36196 (N_36196,N_32700,N_33745);
xor U36197 (N_36197,N_34001,N_33129);
nand U36198 (N_36198,N_33344,N_32841);
xnor U36199 (N_36199,N_32976,N_33424);
or U36200 (N_36200,N_33520,N_33007);
nor U36201 (N_36201,N_33151,N_33295);
and U36202 (N_36202,N_33309,N_34703);
nand U36203 (N_36203,N_34219,N_34937);
nor U36204 (N_36204,N_33939,N_33905);
nor U36205 (N_36205,N_33970,N_34845);
or U36206 (N_36206,N_33619,N_34614);
or U36207 (N_36207,N_32890,N_34917);
nand U36208 (N_36208,N_33710,N_34257);
nand U36209 (N_36209,N_32825,N_33725);
nor U36210 (N_36210,N_34163,N_33118);
nor U36211 (N_36211,N_34381,N_34051);
or U36212 (N_36212,N_34079,N_33239);
nand U36213 (N_36213,N_33555,N_33858);
or U36214 (N_36214,N_34699,N_32922);
nor U36215 (N_36215,N_33196,N_33587);
or U36216 (N_36216,N_33630,N_33100);
nand U36217 (N_36217,N_34068,N_33258);
or U36218 (N_36218,N_33903,N_33622);
xor U36219 (N_36219,N_33819,N_32951);
and U36220 (N_36220,N_34949,N_33385);
nor U36221 (N_36221,N_34542,N_34362);
and U36222 (N_36222,N_34334,N_34692);
and U36223 (N_36223,N_33910,N_33660);
nand U36224 (N_36224,N_34415,N_34075);
or U36225 (N_36225,N_34048,N_34166);
or U36226 (N_36226,N_33627,N_33242);
nor U36227 (N_36227,N_32894,N_33434);
nor U36228 (N_36228,N_34055,N_34073);
or U36229 (N_36229,N_32885,N_33067);
or U36230 (N_36230,N_32584,N_33909);
nand U36231 (N_36231,N_32636,N_34214);
and U36232 (N_36232,N_34518,N_33461);
nand U36233 (N_36233,N_33135,N_34352);
or U36234 (N_36234,N_33670,N_34574);
xor U36235 (N_36235,N_34016,N_33147);
or U36236 (N_36236,N_33244,N_34146);
nand U36237 (N_36237,N_34273,N_33439);
xnor U36238 (N_36238,N_32820,N_33228);
or U36239 (N_36239,N_32626,N_32913);
or U36240 (N_36240,N_34795,N_34332);
xnor U36241 (N_36241,N_33552,N_33437);
nor U36242 (N_36242,N_33626,N_34194);
nor U36243 (N_36243,N_34136,N_33353);
and U36244 (N_36244,N_32550,N_34755);
xor U36245 (N_36245,N_33328,N_34952);
and U36246 (N_36246,N_33267,N_34403);
and U36247 (N_36247,N_33942,N_32528);
nand U36248 (N_36248,N_34325,N_33459);
nand U36249 (N_36249,N_33214,N_34516);
or U36250 (N_36250,N_33795,N_34086);
and U36251 (N_36251,N_32627,N_34048);
or U36252 (N_36252,N_33483,N_33425);
xor U36253 (N_36253,N_32555,N_33924);
xnor U36254 (N_36254,N_34702,N_34668);
xor U36255 (N_36255,N_34098,N_33132);
and U36256 (N_36256,N_32506,N_33228);
nand U36257 (N_36257,N_32513,N_32768);
nor U36258 (N_36258,N_34755,N_34974);
or U36259 (N_36259,N_34404,N_32525);
or U36260 (N_36260,N_33819,N_32910);
nor U36261 (N_36261,N_33993,N_33664);
or U36262 (N_36262,N_32592,N_34357);
and U36263 (N_36263,N_33003,N_34080);
or U36264 (N_36264,N_33638,N_33790);
xor U36265 (N_36265,N_34528,N_33136);
or U36266 (N_36266,N_34067,N_33954);
nor U36267 (N_36267,N_34705,N_32888);
nand U36268 (N_36268,N_34128,N_33994);
or U36269 (N_36269,N_34925,N_33751);
xnor U36270 (N_36270,N_33955,N_32571);
and U36271 (N_36271,N_34105,N_34779);
nand U36272 (N_36272,N_33292,N_34410);
and U36273 (N_36273,N_34959,N_34199);
xnor U36274 (N_36274,N_34736,N_34693);
or U36275 (N_36275,N_32660,N_32983);
or U36276 (N_36276,N_33183,N_34290);
and U36277 (N_36277,N_32581,N_33984);
nor U36278 (N_36278,N_32586,N_32615);
nand U36279 (N_36279,N_33672,N_34419);
or U36280 (N_36280,N_33768,N_34526);
nand U36281 (N_36281,N_32732,N_33971);
nand U36282 (N_36282,N_33301,N_33789);
nand U36283 (N_36283,N_32818,N_34300);
and U36284 (N_36284,N_33471,N_34716);
nor U36285 (N_36285,N_32593,N_33068);
xor U36286 (N_36286,N_34547,N_32793);
nor U36287 (N_36287,N_33861,N_34544);
nand U36288 (N_36288,N_34629,N_33322);
and U36289 (N_36289,N_34045,N_34490);
or U36290 (N_36290,N_32738,N_34888);
or U36291 (N_36291,N_32886,N_33004);
xnor U36292 (N_36292,N_33913,N_32827);
nor U36293 (N_36293,N_32623,N_33840);
nor U36294 (N_36294,N_32856,N_33351);
nand U36295 (N_36295,N_32647,N_32747);
and U36296 (N_36296,N_34190,N_33752);
xor U36297 (N_36297,N_34429,N_32779);
nor U36298 (N_36298,N_34686,N_33942);
and U36299 (N_36299,N_34694,N_34223);
and U36300 (N_36300,N_33830,N_32743);
and U36301 (N_36301,N_33356,N_34665);
xnor U36302 (N_36302,N_34304,N_34699);
and U36303 (N_36303,N_33467,N_32740);
and U36304 (N_36304,N_33986,N_33056);
nor U36305 (N_36305,N_34764,N_33018);
and U36306 (N_36306,N_34510,N_32759);
and U36307 (N_36307,N_34636,N_33414);
nor U36308 (N_36308,N_33857,N_34991);
nand U36309 (N_36309,N_34225,N_33442);
or U36310 (N_36310,N_34070,N_34486);
nand U36311 (N_36311,N_33097,N_33762);
or U36312 (N_36312,N_34994,N_32636);
or U36313 (N_36313,N_33247,N_34282);
nand U36314 (N_36314,N_32706,N_32578);
or U36315 (N_36315,N_34616,N_33265);
nand U36316 (N_36316,N_34704,N_34709);
xnor U36317 (N_36317,N_34777,N_33113);
or U36318 (N_36318,N_34542,N_32505);
xnor U36319 (N_36319,N_32832,N_33249);
xor U36320 (N_36320,N_34892,N_33054);
nand U36321 (N_36321,N_33704,N_33661);
and U36322 (N_36322,N_34756,N_34665);
xnor U36323 (N_36323,N_33436,N_34455);
or U36324 (N_36324,N_34696,N_32548);
or U36325 (N_36325,N_33708,N_32688);
xor U36326 (N_36326,N_33102,N_34109);
and U36327 (N_36327,N_32710,N_34006);
and U36328 (N_36328,N_33232,N_33603);
xnor U36329 (N_36329,N_34073,N_33664);
nor U36330 (N_36330,N_32788,N_34807);
or U36331 (N_36331,N_34483,N_33372);
nor U36332 (N_36332,N_33566,N_34055);
or U36333 (N_36333,N_34849,N_34325);
nor U36334 (N_36334,N_34338,N_34135);
nor U36335 (N_36335,N_34245,N_33511);
or U36336 (N_36336,N_33905,N_33592);
nand U36337 (N_36337,N_32781,N_33123);
xnor U36338 (N_36338,N_33384,N_34695);
nand U36339 (N_36339,N_33380,N_34952);
xor U36340 (N_36340,N_32713,N_32778);
nand U36341 (N_36341,N_32692,N_32866);
xor U36342 (N_36342,N_34414,N_34950);
and U36343 (N_36343,N_33995,N_34175);
nor U36344 (N_36344,N_34813,N_33285);
nand U36345 (N_36345,N_32650,N_34449);
nor U36346 (N_36346,N_33136,N_34997);
or U36347 (N_36347,N_33892,N_34820);
and U36348 (N_36348,N_33862,N_33170);
nand U36349 (N_36349,N_32501,N_34369);
nand U36350 (N_36350,N_33230,N_34021);
xor U36351 (N_36351,N_32609,N_34876);
or U36352 (N_36352,N_32670,N_34056);
or U36353 (N_36353,N_34786,N_34161);
or U36354 (N_36354,N_33222,N_33264);
and U36355 (N_36355,N_33487,N_34960);
xnor U36356 (N_36356,N_32584,N_34132);
and U36357 (N_36357,N_33204,N_34360);
or U36358 (N_36358,N_34880,N_34944);
and U36359 (N_36359,N_34658,N_33908);
xor U36360 (N_36360,N_34656,N_33506);
nor U36361 (N_36361,N_33520,N_34941);
or U36362 (N_36362,N_32971,N_33167);
nor U36363 (N_36363,N_34949,N_32728);
xor U36364 (N_36364,N_33491,N_32683);
and U36365 (N_36365,N_34048,N_34669);
nor U36366 (N_36366,N_32749,N_32724);
or U36367 (N_36367,N_33064,N_32967);
or U36368 (N_36368,N_34791,N_33453);
or U36369 (N_36369,N_33203,N_32987);
or U36370 (N_36370,N_34638,N_33460);
and U36371 (N_36371,N_32565,N_33723);
nor U36372 (N_36372,N_32894,N_34051);
nor U36373 (N_36373,N_34821,N_34818);
nand U36374 (N_36374,N_34057,N_34668);
nand U36375 (N_36375,N_33066,N_33125);
xnor U36376 (N_36376,N_33094,N_33668);
and U36377 (N_36377,N_32874,N_33575);
xnor U36378 (N_36378,N_34674,N_34673);
or U36379 (N_36379,N_33052,N_32719);
or U36380 (N_36380,N_33270,N_34705);
xor U36381 (N_36381,N_34388,N_32623);
nand U36382 (N_36382,N_34690,N_33262);
nor U36383 (N_36383,N_34502,N_34926);
xor U36384 (N_36384,N_34209,N_34401);
or U36385 (N_36385,N_33652,N_33529);
or U36386 (N_36386,N_32568,N_32640);
or U36387 (N_36387,N_34568,N_33140);
and U36388 (N_36388,N_32749,N_34386);
nor U36389 (N_36389,N_33631,N_34582);
or U36390 (N_36390,N_34858,N_32736);
or U36391 (N_36391,N_34962,N_34441);
nor U36392 (N_36392,N_32735,N_34679);
or U36393 (N_36393,N_33277,N_33223);
nand U36394 (N_36394,N_34586,N_32748);
nor U36395 (N_36395,N_32674,N_34405);
and U36396 (N_36396,N_33146,N_33183);
nor U36397 (N_36397,N_33946,N_32958);
or U36398 (N_36398,N_32995,N_34206);
and U36399 (N_36399,N_33687,N_34989);
or U36400 (N_36400,N_33292,N_33838);
and U36401 (N_36401,N_33150,N_32554);
nand U36402 (N_36402,N_33315,N_34581);
xnor U36403 (N_36403,N_34493,N_33043);
xnor U36404 (N_36404,N_32710,N_33460);
and U36405 (N_36405,N_33488,N_32926);
nand U36406 (N_36406,N_32838,N_33351);
and U36407 (N_36407,N_34110,N_33886);
xnor U36408 (N_36408,N_32841,N_33544);
or U36409 (N_36409,N_33762,N_34591);
and U36410 (N_36410,N_32619,N_32578);
nor U36411 (N_36411,N_33435,N_32776);
nor U36412 (N_36412,N_33277,N_33759);
nor U36413 (N_36413,N_32984,N_34736);
or U36414 (N_36414,N_34860,N_33302);
nor U36415 (N_36415,N_34708,N_33681);
xor U36416 (N_36416,N_34389,N_33211);
or U36417 (N_36417,N_32896,N_34245);
and U36418 (N_36418,N_33112,N_34175);
xnor U36419 (N_36419,N_33928,N_32567);
nor U36420 (N_36420,N_33130,N_34394);
nand U36421 (N_36421,N_33910,N_33696);
and U36422 (N_36422,N_33097,N_33325);
and U36423 (N_36423,N_33197,N_33524);
xnor U36424 (N_36424,N_32857,N_33747);
xnor U36425 (N_36425,N_32645,N_33656);
and U36426 (N_36426,N_33760,N_34586);
nand U36427 (N_36427,N_33199,N_34369);
nor U36428 (N_36428,N_34858,N_33958);
or U36429 (N_36429,N_34966,N_34637);
nand U36430 (N_36430,N_34266,N_34841);
or U36431 (N_36431,N_32663,N_34356);
or U36432 (N_36432,N_34154,N_32639);
or U36433 (N_36433,N_33402,N_32541);
xnor U36434 (N_36434,N_34725,N_34076);
xnor U36435 (N_36435,N_34433,N_33992);
and U36436 (N_36436,N_33738,N_32979);
xor U36437 (N_36437,N_33495,N_34621);
and U36438 (N_36438,N_33288,N_33954);
xnor U36439 (N_36439,N_34129,N_33807);
xnor U36440 (N_36440,N_33980,N_34478);
or U36441 (N_36441,N_34648,N_32810);
and U36442 (N_36442,N_32808,N_33052);
or U36443 (N_36443,N_34984,N_32989);
nor U36444 (N_36444,N_33255,N_33225);
nor U36445 (N_36445,N_33566,N_32899);
nor U36446 (N_36446,N_34022,N_34480);
nand U36447 (N_36447,N_33495,N_34660);
and U36448 (N_36448,N_32595,N_34216);
nor U36449 (N_36449,N_33112,N_33538);
xor U36450 (N_36450,N_34415,N_34634);
or U36451 (N_36451,N_34538,N_34704);
nor U36452 (N_36452,N_33004,N_32823);
nand U36453 (N_36453,N_32988,N_33722);
and U36454 (N_36454,N_32733,N_33268);
and U36455 (N_36455,N_32969,N_32593);
nor U36456 (N_36456,N_34931,N_32657);
nand U36457 (N_36457,N_33281,N_32999);
xnor U36458 (N_36458,N_34933,N_33952);
and U36459 (N_36459,N_33500,N_33950);
nor U36460 (N_36460,N_32811,N_33583);
xnor U36461 (N_36461,N_34094,N_33409);
nor U36462 (N_36462,N_32577,N_34715);
and U36463 (N_36463,N_32658,N_34312);
nand U36464 (N_36464,N_33613,N_34732);
xnor U36465 (N_36465,N_34897,N_33100);
and U36466 (N_36466,N_34078,N_33889);
nor U36467 (N_36467,N_32870,N_33358);
nor U36468 (N_36468,N_34657,N_34786);
nor U36469 (N_36469,N_34427,N_34433);
xor U36470 (N_36470,N_33784,N_34045);
nand U36471 (N_36471,N_33833,N_32640);
nor U36472 (N_36472,N_33674,N_34786);
xor U36473 (N_36473,N_32823,N_34017);
nor U36474 (N_36474,N_34458,N_34565);
and U36475 (N_36475,N_34515,N_34912);
xnor U36476 (N_36476,N_34454,N_34982);
xnor U36477 (N_36477,N_34406,N_32832);
nor U36478 (N_36478,N_32864,N_32634);
xor U36479 (N_36479,N_32512,N_34482);
and U36480 (N_36480,N_34605,N_33933);
xor U36481 (N_36481,N_32838,N_33497);
and U36482 (N_36482,N_34011,N_33362);
nand U36483 (N_36483,N_34283,N_34466);
nand U36484 (N_36484,N_34614,N_33149);
and U36485 (N_36485,N_32759,N_32611);
and U36486 (N_36486,N_33361,N_34888);
nand U36487 (N_36487,N_33295,N_34411);
nand U36488 (N_36488,N_32991,N_34961);
nand U36489 (N_36489,N_34821,N_33237);
xnor U36490 (N_36490,N_33785,N_33258);
or U36491 (N_36491,N_33519,N_33212);
nand U36492 (N_36492,N_33194,N_34034);
xor U36493 (N_36493,N_33783,N_32603);
xnor U36494 (N_36494,N_33482,N_33662);
xor U36495 (N_36495,N_34500,N_32845);
xor U36496 (N_36496,N_34408,N_34650);
nor U36497 (N_36497,N_33136,N_34866);
or U36498 (N_36498,N_34704,N_34710);
nor U36499 (N_36499,N_33941,N_34411);
or U36500 (N_36500,N_32664,N_33222);
or U36501 (N_36501,N_34405,N_33757);
nand U36502 (N_36502,N_34940,N_33357);
and U36503 (N_36503,N_34283,N_33076);
nand U36504 (N_36504,N_34395,N_34941);
nor U36505 (N_36505,N_34817,N_32514);
nor U36506 (N_36506,N_34163,N_33435);
xnor U36507 (N_36507,N_34684,N_34060);
nand U36508 (N_36508,N_32767,N_33397);
nand U36509 (N_36509,N_33678,N_33032);
nand U36510 (N_36510,N_34046,N_34827);
or U36511 (N_36511,N_33474,N_32896);
nand U36512 (N_36512,N_33424,N_34503);
nor U36513 (N_36513,N_34252,N_34925);
or U36514 (N_36514,N_34828,N_33861);
xnor U36515 (N_36515,N_34483,N_32982);
nor U36516 (N_36516,N_34522,N_34619);
xor U36517 (N_36517,N_32985,N_32512);
or U36518 (N_36518,N_33644,N_34598);
nor U36519 (N_36519,N_34069,N_34479);
or U36520 (N_36520,N_34889,N_33108);
and U36521 (N_36521,N_33248,N_34670);
nand U36522 (N_36522,N_33593,N_32986);
xnor U36523 (N_36523,N_34414,N_34305);
nor U36524 (N_36524,N_34319,N_34724);
or U36525 (N_36525,N_33957,N_33776);
nor U36526 (N_36526,N_34100,N_34572);
nand U36527 (N_36527,N_33870,N_33218);
nand U36528 (N_36528,N_33364,N_34091);
or U36529 (N_36529,N_33493,N_33649);
nor U36530 (N_36530,N_32946,N_32695);
xnor U36531 (N_36531,N_32612,N_34211);
nor U36532 (N_36532,N_34787,N_34727);
or U36533 (N_36533,N_33159,N_33118);
xor U36534 (N_36534,N_34693,N_32639);
nor U36535 (N_36535,N_33395,N_34433);
nand U36536 (N_36536,N_33205,N_34519);
xor U36537 (N_36537,N_33517,N_33611);
nand U36538 (N_36538,N_34960,N_32597);
xor U36539 (N_36539,N_34647,N_34499);
nand U36540 (N_36540,N_33742,N_34917);
xnor U36541 (N_36541,N_34450,N_32518);
xnor U36542 (N_36542,N_33247,N_33731);
nand U36543 (N_36543,N_34880,N_33076);
or U36544 (N_36544,N_32942,N_34073);
nor U36545 (N_36545,N_34940,N_32941);
and U36546 (N_36546,N_32673,N_34369);
xnor U36547 (N_36547,N_34977,N_33990);
xnor U36548 (N_36548,N_33862,N_33453);
nand U36549 (N_36549,N_33793,N_33133);
and U36550 (N_36550,N_32634,N_32756);
nor U36551 (N_36551,N_34054,N_33446);
nand U36552 (N_36552,N_32696,N_33294);
nor U36553 (N_36553,N_34355,N_32862);
nand U36554 (N_36554,N_34294,N_34660);
nor U36555 (N_36555,N_34416,N_33906);
nand U36556 (N_36556,N_34411,N_33924);
or U36557 (N_36557,N_34755,N_33038);
and U36558 (N_36558,N_33451,N_34413);
or U36559 (N_36559,N_33845,N_32677);
nand U36560 (N_36560,N_33657,N_33196);
or U36561 (N_36561,N_34952,N_33895);
and U36562 (N_36562,N_33136,N_32607);
xor U36563 (N_36563,N_32603,N_32543);
nand U36564 (N_36564,N_34939,N_34465);
nand U36565 (N_36565,N_32516,N_33661);
nor U36566 (N_36566,N_33830,N_33103);
nand U36567 (N_36567,N_34094,N_32561);
or U36568 (N_36568,N_32711,N_32988);
or U36569 (N_36569,N_33223,N_33255);
or U36570 (N_36570,N_33987,N_33639);
and U36571 (N_36571,N_32709,N_34893);
xnor U36572 (N_36572,N_34903,N_32761);
nand U36573 (N_36573,N_34015,N_32586);
or U36574 (N_36574,N_34876,N_34990);
nand U36575 (N_36575,N_34254,N_33654);
nor U36576 (N_36576,N_32507,N_34254);
and U36577 (N_36577,N_34524,N_33702);
and U36578 (N_36578,N_34968,N_34929);
xor U36579 (N_36579,N_33907,N_33382);
or U36580 (N_36580,N_34518,N_32840);
nor U36581 (N_36581,N_33583,N_33252);
or U36582 (N_36582,N_34194,N_33798);
xor U36583 (N_36583,N_34791,N_33382);
or U36584 (N_36584,N_34287,N_33880);
and U36585 (N_36585,N_33559,N_34643);
xnor U36586 (N_36586,N_32577,N_34636);
or U36587 (N_36587,N_34249,N_34334);
nand U36588 (N_36588,N_32818,N_34194);
and U36589 (N_36589,N_32909,N_32707);
nor U36590 (N_36590,N_32966,N_34822);
xnor U36591 (N_36591,N_33790,N_34414);
and U36592 (N_36592,N_33824,N_32569);
nand U36593 (N_36593,N_33963,N_33486);
and U36594 (N_36594,N_33229,N_32810);
xnor U36595 (N_36595,N_34081,N_33469);
xor U36596 (N_36596,N_34669,N_34047);
nand U36597 (N_36597,N_33883,N_34690);
nand U36598 (N_36598,N_33898,N_33717);
and U36599 (N_36599,N_33368,N_33889);
xor U36600 (N_36600,N_32509,N_33335);
and U36601 (N_36601,N_33949,N_34791);
xnor U36602 (N_36602,N_33625,N_33064);
or U36603 (N_36603,N_32597,N_32620);
and U36604 (N_36604,N_33856,N_33373);
nand U36605 (N_36605,N_33909,N_32678);
and U36606 (N_36606,N_33698,N_33643);
nor U36607 (N_36607,N_34047,N_32907);
and U36608 (N_36608,N_32506,N_32508);
nand U36609 (N_36609,N_34480,N_33198);
and U36610 (N_36610,N_32573,N_33896);
nand U36611 (N_36611,N_32659,N_34461);
xnor U36612 (N_36612,N_33150,N_33233);
or U36613 (N_36613,N_32900,N_33590);
nand U36614 (N_36614,N_34357,N_33153);
xor U36615 (N_36615,N_33735,N_33591);
and U36616 (N_36616,N_34493,N_32959);
or U36617 (N_36617,N_34086,N_34333);
nor U36618 (N_36618,N_34275,N_33808);
and U36619 (N_36619,N_32912,N_33223);
or U36620 (N_36620,N_34784,N_33137);
nand U36621 (N_36621,N_33810,N_34159);
xor U36622 (N_36622,N_33354,N_33218);
xor U36623 (N_36623,N_32940,N_33211);
nand U36624 (N_36624,N_33413,N_34041);
nor U36625 (N_36625,N_34094,N_34818);
nand U36626 (N_36626,N_32525,N_32630);
xnor U36627 (N_36627,N_33168,N_32787);
nor U36628 (N_36628,N_34690,N_32696);
xor U36629 (N_36629,N_33942,N_32951);
nor U36630 (N_36630,N_34188,N_34168);
nor U36631 (N_36631,N_34554,N_34065);
and U36632 (N_36632,N_34262,N_34418);
nor U36633 (N_36633,N_33065,N_32831);
or U36634 (N_36634,N_34244,N_33234);
or U36635 (N_36635,N_32995,N_33093);
xor U36636 (N_36636,N_33468,N_33616);
xnor U36637 (N_36637,N_34371,N_33511);
xnor U36638 (N_36638,N_34378,N_33246);
nand U36639 (N_36639,N_34783,N_34488);
xor U36640 (N_36640,N_32875,N_34742);
or U36641 (N_36641,N_34890,N_33172);
or U36642 (N_36642,N_33127,N_33099);
xnor U36643 (N_36643,N_32736,N_34640);
xor U36644 (N_36644,N_34616,N_32939);
and U36645 (N_36645,N_34502,N_34062);
or U36646 (N_36646,N_34305,N_33190);
xnor U36647 (N_36647,N_33700,N_33405);
or U36648 (N_36648,N_33310,N_33863);
or U36649 (N_36649,N_34228,N_34135);
nor U36650 (N_36650,N_33664,N_33353);
xnor U36651 (N_36651,N_34116,N_33938);
xor U36652 (N_36652,N_34659,N_33335);
or U36653 (N_36653,N_32892,N_32731);
or U36654 (N_36654,N_34580,N_34529);
nor U36655 (N_36655,N_33091,N_34724);
nand U36656 (N_36656,N_34850,N_34804);
and U36657 (N_36657,N_33431,N_32769);
nor U36658 (N_36658,N_34715,N_34877);
and U36659 (N_36659,N_33559,N_33048);
nor U36660 (N_36660,N_32625,N_34166);
and U36661 (N_36661,N_33004,N_33356);
and U36662 (N_36662,N_33228,N_33499);
nand U36663 (N_36663,N_34189,N_34589);
nand U36664 (N_36664,N_33530,N_34062);
or U36665 (N_36665,N_33258,N_34355);
nand U36666 (N_36666,N_33970,N_33229);
xnor U36667 (N_36667,N_33054,N_33145);
or U36668 (N_36668,N_33082,N_34947);
nor U36669 (N_36669,N_34625,N_33726);
and U36670 (N_36670,N_33825,N_34720);
xor U36671 (N_36671,N_34538,N_33584);
xor U36672 (N_36672,N_34252,N_34519);
nor U36673 (N_36673,N_33403,N_32729);
nor U36674 (N_36674,N_32939,N_33576);
xor U36675 (N_36675,N_32635,N_34895);
xnor U36676 (N_36676,N_33160,N_32926);
nor U36677 (N_36677,N_33938,N_33865);
xnor U36678 (N_36678,N_32944,N_33335);
and U36679 (N_36679,N_33079,N_33571);
nor U36680 (N_36680,N_34950,N_33056);
and U36681 (N_36681,N_34294,N_34828);
nor U36682 (N_36682,N_34908,N_33926);
nor U36683 (N_36683,N_33501,N_34873);
nor U36684 (N_36684,N_33353,N_34415);
or U36685 (N_36685,N_33376,N_33870);
and U36686 (N_36686,N_33382,N_34780);
nor U36687 (N_36687,N_33613,N_34010);
nand U36688 (N_36688,N_33129,N_33866);
xor U36689 (N_36689,N_34651,N_33919);
or U36690 (N_36690,N_32838,N_33288);
xor U36691 (N_36691,N_33528,N_33592);
nand U36692 (N_36692,N_33600,N_34484);
nand U36693 (N_36693,N_33239,N_34749);
nand U36694 (N_36694,N_34283,N_32703);
nor U36695 (N_36695,N_33366,N_33696);
nand U36696 (N_36696,N_33512,N_33083);
nand U36697 (N_36697,N_34028,N_33964);
and U36698 (N_36698,N_34187,N_34995);
and U36699 (N_36699,N_33832,N_33724);
nand U36700 (N_36700,N_34772,N_34145);
and U36701 (N_36701,N_33554,N_33214);
nor U36702 (N_36702,N_34203,N_33615);
nand U36703 (N_36703,N_32863,N_33483);
nor U36704 (N_36704,N_32835,N_32704);
and U36705 (N_36705,N_33545,N_32645);
nor U36706 (N_36706,N_34199,N_34142);
or U36707 (N_36707,N_32968,N_34292);
nor U36708 (N_36708,N_32970,N_32585);
nor U36709 (N_36709,N_32635,N_34415);
nor U36710 (N_36710,N_34626,N_34233);
or U36711 (N_36711,N_33908,N_34342);
or U36712 (N_36712,N_33561,N_34838);
or U36713 (N_36713,N_34566,N_33303);
or U36714 (N_36714,N_32797,N_34115);
and U36715 (N_36715,N_33477,N_34658);
nor U36716 (N_36716,N_34553,N_34454);
and U36717 (N_36717,N_32913,N_33443);
or U36718 (N_36718,N_33799,N_34823);
or U36719 (N_36719,N_32872,N_34192);
or U36720 (N_36720,N_33711,N_33220);
xnor U36721 (N_36721,N_34369,N_32741);
and U36722 (N_36722,N_32793,N_33550);
and U36723 (N_36723,N_33295,N_32926);
nor U36724 (N_36724,N_33896,N_34913);
xor U36725 (N_36725,N_34037,N_33033);
xnor U36726 (N_36726,N_34906,N_33079);
xnor U36727 (N_36727,N_34821,N_34028);
and U36728 (N_36728,N_32815,N_32539);
or U36729 (N_36729,N_32521,N_34679);
xnor U36730 (N_36730,N_33096,N_32802);
nor U36731 (N_36731,N_33165,N_33603);
nand U36732 (N_36732,N_34633,N_33881);
and U36733 (N_36733,N_32972,N_33849);
xnor U36734 (N_36734,N_34792,N_32945);
nand U36735 (N_36735,N_34410,N_34644);
xor U36736 (N_36736,N_34913,N_34119);
xnor U36737 (N_36737,N_32780,N_33511);
nand U36738 (N_36738,N_32858,N_32957);
nor U36739 (N_36739,N_33623,N_32980);
nand U36740 (N_36740,N_34687,N_33228);
xnor U36741 (N_36741,N_33807,N_32540);
nand U36742 (N_36742,N_33663,N_33954);
nor U36743 (N_36743,N_33839,N_34884);
and U36744 (N_36744,N_34895,N_32800);
or U36745 (N_36745,N_34985,N_33689);
xnor U36746 (N_36746,N_33369,N_34900);
nand U36747 (N_36747,N_32844,N_34595);
xnor U36748 (N_36748,N_33139,N_32814);
nor U36749 (N_36749,N_34043,N_34211);
nand U36750 (N_36750,N_34757,N_34059);
and U36751 (N_36751,N_33697,N_34668);
nor U36752 (N_36752,N_34776,N_34488);
nor U36753 (N_36753,N_32734,N_33166);
xnor U36754 (N_36754,N_33087,N_34959);
xnor U36755 (N_36755,N_33344,N_34467);
and U36756 (N_36756,N_34204,N_33775);
xor U36757 (N_36757,N_33651,N_33823);
or U36758 (N_36758,N_34661,N_33493);
nand U36759 (N_36759,N_34738,N_34125);
xor U36760 (N_36760,N_34732,N_32554);
nand U36761 (N_36761,N_34866,N_33392);
xor U36762 (N_36762,N_34299,N_33887);
nor U36763 (N_36763,N_32977,N_34091);
nor U36764 (N_36764,N_32935,N_32516);
nand U36765 (N_36765,N_34782,N_34310);
xnor U36766 (N_36766,N_33428,N_32560);
nand U36767 (N_36767,N_34978,N_33525);
nor U36768 (N_36768,N_33047,N_33191);
nor U36769 (N_36769,N_34735,N_32800);
or U36770 (N_36770,N_34915,N_32539);
nor U36771 (N_36771,N_33274,N_34826);
xnor U36772 (N_36772,N_33077,N_32839);
nand U36773 (N_36773,N_33118,N_33489);
nand U36774 (N_36774,N_34265,N_34763);
xnor U36775 (N_36775,N_34535,N_34551);
nand U36776 (N_36776,N_33141,N_32817);
xnor U36777 (N_36777,N_33010,N_34393);
xor U36778 (N_36778,N_34736,N_32510);
nor U36779 (N_36779,N_34231,N_34199);
nand U36780 (N_36780,N_34350,N_33738);
xnor U36781 (N_36781,N_33426,N_32672);
or U36782 (N_36782,N_33052,N_34863);
nor U36783 (N_36783,N_32784,N_33539);
xnor U36784 (N_36784,N_34495,N_32591);
nor U36785 (N_36785,N_34636,N_33770);
and U36786 (N_36786,N_34281,N_34644);
and U36787 (N_36787,N_34053,N_33700);
xnor U36788 (N_36788,N_34246,N_34313);
and U36789 (N_36789,N_32894,N_32676);
nand U36790 (N_36790,N_34117,N_33827);
xnor U36791 (N_36791,N_33834,N_33303);
or U36792 (N_36792,N_34893,N_32847);
or U36793 (N_36793,N_33155,N_34317);
nand U36794 (N_36794,N_32967,N_33150);
xnor U36795 (N_36795,N_33412,N_33673);
and U36796 (N_36796,N_34503,N_32555);
nor U36797 (N_36797,N_33775,N_32690);
nand U36798 (N_36798,N_32939,N_33622);
and U36799 (N_36799,N_32701,N_33274);
or U36800 (N_36800,N_33636,N_34675);
xnor U36801 (N_36801,N_33202,N_32902);
xor U36802 (N_36802,N_33974,N_33264);
nand U36803 (N_36803,N_34564,N_33521);
and U36804 (N_36804,N_34227,N_32753);
and U36805 (N_36805,N_33773,N_33878);
nor U36806 (N_36806,N_32863,N_34915);
xor U36807 (N_36807,N_32628,N_32657);
and U36808 (N_36808,N_34709,N_32768);
nand U36809 (N_36809,N_33441,N_33197);
nand U36810 (N_36810,N_34318,N_33541);
or U36811 (N_36811,N_34917,N_33182);
or U36812 (N_36812,N_32659,N_34253);
or U36813 (N_36813,N_33975,N_34286);
nor U36814 (N_36814,N_32697,N_34684);
nand U36815 (N_36815,N_34129,N_33262);
xor U36816 (N_36816,N_32791,N_34753);
xor U36817 (N_36817,N_32977,N_34604);
nand U36818 (N_36818,N_34970,N_33481);
and U36819 (N_36819,N_33730,N_32760);
nor U36820 (N_36820,N_33324,N_32521);
and U36821 (N_36821,N_32670,N_32539);
or U36822 (N_36822,N_33955,N_34434);
nand U36823 (N_36823,N_34753,N_32579);
xor U36824 (N_36824,N_33597,N_34833);
xor U36825 (N_36825,N_33609,N_33329);
or U36826 (N_36826,N_33536,N_33188);
xnor U36827 (N_36827,N_32730,N_34280);
nand U36828 (N_36828,N_33702,N_34558);
xor U36829 (N_36829,N_33802,N_33293);
and U36830 (N_36830,N_32863,N_32940);
or U36831 (N_36831,N_32820,N_33769);
xor U36832 (N_36832,N_33673,N_33341);
or U36833 (N_36833,N_34042,N_33160);
or U36834 (N_36834,N_33311,N_34157);
xor U36835 (N_36835,N_34984,N_32665);
nor U36836 (N_36836,N_33247,N_33514);
and U36837 (N_36837,N_34623,N_34148);
or U36838 (N_36838,N_32560,N_33502);
and U36839 (N_36839,N_34162,N_32902);
nand U36840 (N_36840,N_34142,N_34034);
and U36841 (N_36841,N_33007,N_33154);
and U36842 (N_36842,N_33944,N_33709);
nand U36843 (N_36843,N_33575,N_33057);
xnor U36844 (N_36844,N_33801,N_33815);
or U36845 (N_36845,N_33687,N_32936);
or U36846 (N_36846,N_32577,N_32739);
xnor U36847 (N_36847,N_34872,N_32746);
xor U36848 (N_36848,N_32572,N_33785);
nor U36849 (N_36849,N_34272,N_33006);
nor U36850 (N_36850,N_32772,N_34584);
xor U36851 (N_36851,N_34426,N_34280);
xor U36852 (N_36852,N_33808,N_34850);
xor U36853 (N_36853,N_34472,N_33051);
nor U36854 (N_36854,N_33937,N_34918);
or U36855 (N_36855,N_33468,N_34994);
or U36856 (N_36856,N_34067,N_33846);
nand U36857 (N_36857,N_33556,N_33887);
and U36858 (N_36858,N_34443,N_34237);
or U36859 (N_36859,N_32765,N_32712);
xnor U36860 (N_36860,N_34010,N_34084);
or U36861 (N_36861,N_32636,N_32777);
and U36862 (N_36862,N_33597,N_34513);
and U36863 (N_36863,N_33358,N_33233);
nor U36864 (N_36864,N_34151,N_32688);
nor U36865 (N_36865,N_33547,N_34224);
or U36866 (N_36866,N_33605,N_33310);
or U36867 (N_36867,N_32566,N_34314);
nand U36868 (N_36868,N_34825,N_34086);
and U36869 (N_36869,N_34293,N_32934);
nand U36870 (N_36870,N_34864,N_33762);
xnor U36871 (N_36871,N_33796,N_33072);
or U36872 (N_36872,N_33878,N_34580);
or U36873 (N_36873,N_33016,N_32854);
nand U36874 (N_36874,N_33106,N_33456);
and U36875 (N_36875,N_34834,N_34017);
or U36876 (N_36876,N_32966,N_33229);
and U36877 (N_36877,N_34754,N_32771);
nor U36878 (N_36878,N_34560,N_33392);
xor U36879 (N_36879,N_33783,N_34326);
xnor U36880 (N_36880,N_33891,N_33025);
and U36881 (N_36881,N_33461,N_34636);
xor U36882 (N_36882,N_33564,N_32533);
xnor U36883 (N_36883,N_33264,N_34674);
nand U36884 (N_36884,N_34978,N_32559);
and U36885 (N_36885,N_34925,N_34269);
and U36886 (N_36886,N_34539,N_32848);
or U36887 (N_36887,N_32996,N_33750);
nand U36888 (N_36888,N_33443,N_32728);
nand U36889 (N_36889,N_34865,N_33618);
nor U36890 (N_36890,N_33331,N_33578);
nand U36891 (N_36891,N_33797,N_34889);
xor U36892 (N_36892,N_32678,N_33567);
and U36893 (N_36893,N_34145,N_34864);
and U36894 (N_36894,N_32827,N_33356);
and U36895 (N_36895,N_34662,N_33359);
xor U36896 (N_36896,N_34104,N_34650);
nor U36897 (N_36897,N_33233,N_33491);
xnor U36898 (N_36898,N_34729,N_33224);
nor U36899 (N_36899,N_33810,N_32803);
xnor U36900 (N_36900,N_32644,N_33105);
nor U36901 (N_36901,N_34670,N_33397);
and U36902 (N_36902,N_33343,N_33147);
or U36903 (N_36903,N_34623,N_34548);
or U36904 (N_36904,N_33597,N_34125);
nand U36905 (N_36905,N_34769,N_32545);
nand U36906 (N_36906,N_33707,N_32558);
nand U36907 (N_36907,N_34018,N_33468);
or U36908 (N_36908,N_33446,N_32541);
and U36909 (N_36909,N_33565,N_34662);
and U36910 (N_36910,N_34793,N_33102);
xnor U36911 (N_36911,N_34608,N_34667);
nand U36912 (N_36912,N_33624,N_34901);
or U36913 (N_36913,N_34896,N_34995);
nand U36914 (N_36914,N_33806,N_34032);
nor U36915 (N_36915,N_34582,N_32953);
xor U36916 (N_36916,N_32961,N_34378);
xnor U36917 (N_36917,N_33016,N_33578);
and U36918 (N_36918,N_33128,N_33054);
or U36919 (N_36919,N_32621,N_34277);
or U36920 (N_36920,N_33986,N_33635);
xnor U36921 (N_36921,N_33222,N_33337);
or U36922 (N_36922,N_34051,N_33251);
or U36923 (N_36923,N_32643,N_34531);
xor U36924 (N_36924,N_34559,N_33722);
or U36925 (N_36925,N_32909,N_33864);
nand U36926 (N_36926,N_34533,N_34695);
xor U36927 (N_36927,N_33866,N_32877);
or U36928 (N_36928,N_33242,N_34121);
nand U36929 (N_36929,N_33739,N_33104);
nand U36930 (N_36930,N_34965,N_33176);
nor U36931 (N_36931,N_34272,N_34176);
or U36932 (N_36932,N_33456,N_33745);
nand U36933 (N_36933,N_34581,N_34652);
xnor U36934 (N_36934,N_34855,N_33500);
and U36935 (N_36935,N_34075,N_32543);
nand U36936 (N_36936,N_32735,N_33594);
nor U36937 (N_36937,N_33985,N_33538);
xor U36938 (N_36938,N_33467,N_34967);
nor U36939 (N_36939,N_34512,N_34789);
xor U36940 (N_36940,N_34424,N_33693);
or U36941 (N_36941,N_34245,N_33379);
or U36942 (N_36942,N_34782,N_32814);
and U36943 (N_36943,N_34678,N_34547);
and U36944 (N_36944,N_32577,N_34594);
xor U36945 (N_36945,N_33343,N_33974);
xnor U36946 (N_36946,N_33984,N_32893);
nand U36947 (N_36947,N_34469,N_33846);
xor U36948 (N_36948,N_33899,N_34835);
xor U36949 (N_36949,N_33200,N_33803);
nor U36950 (N_36950,N_34077,N_33177);
or U36951 (N_36951,N_33713,N_33899);
and U36952 (N_36952,N_34469,N_34669);
nor U36953 (N_36953,N_33405,N_33339);
nand U36954 (N_36954,N_34802,N_34334);
nor U36955 (N_36955,N_34269,N_34754);
and U36956 (N_36956,N_33370,N_32947);
nor U36957 (N_36957,N_32858,N_32646);
nand U36958 (N_36958,N_33521,N_32852);
or U36959 (N_36959,N_33106,N_34632);
xor U36960 (N_36960,N_33761,N_32594);
xnor U36961 (N_36961,N_32865,N_34984);
xor U36962 (N_36962,N_34352,N_32966);
nand U36963 (N_36963,N_33349,N_33563);
nor U36964 (N_36964,N_32894,N_33146);
or U36965 (N_36965,N_34279,N_34337);
nor U36966 (N_36966,N_32684,N_33867);
or U36967 (N_36967,N_34650,N_33573);
nand U36968 (N_36968,N_32844,N_34293);
and U36969 (N_36969,N_34296,N_33846);
or U36970 (N_36970,N_32695,N_34695);
nor U36971 (N_36971,N_34704,N_34129);
and U36972 (N_36972,N_32672,N_34047);
nand U36973 (N_36973,N_32926,N_33258);
and U36974 (N_36974,N_34405,N_32549);
xnor U36975 (N_36975,N_32829,N_34777);
xor U36976 (N_36976,N_32690,N_34760);
or U36977 (N_36977,N_33584,N_33630);
or U36978 (N_36978,N_33098,N_33958);
nand U36979 (N_36979,N_34637,N_34002);
or U36980 (N_36980,N_34061,N_32904);
nand U36981 (N_36981,N_33468,N_33406);
and U36982 (N_36982,N_34374,N_34237);
or U36983 (N_36983,N_33227,N_34757);
nand U36984 (N_36984,N_32581,N_33738);
or U36985 (N_36985,N_33076,N_34671);
xor U36986 (N_36986,N_32731,N_32871);
and U36987 (N_36987,N_34503,N_32640);
nor U36988 (N_36988,N_34611,N_33964);
nor U36989 (N_36989,N_33620,N_32865);
nor U36990 (N_36990,N_33302,N_34342);
nor U36991 (N_36991,N_33768,N_33604);
nand U36992 (N_36992,N_34975,N_34588);
xor U36993 (N_36993,N_34357,N_34417);
and U36994 (N_36994,N_33287,N_32667);
xor U36995 (N_36995,N_32539,N_34473);
nand U36996 (N_36996,N_34826,N_33532);
or U36997 (N_36997,N_34268,N_34250);
nor U36998 (N_36998,N_33967,N_33353);
and U36999 (N_36999,N_33121,N_33047);
nand U37000 (N_37000,N_34749,N_34379);
xor U37001 (N_37001,N_33288,N_32908);
or U37002 (N_37002,N_34311,N_33310);
and U37003 (N_37003,N_32549,N_33953);
nor U37004 (N_37004,N_32737,N_33528);
or U37005 (N_37005,N_32735,N_33192);
nor U37006 (N_37006,N_33229,N_34489);
nor U37007 (N_37007,N_33208,N_33890);
nor U37008 (N_37008,N_32579,N_32789);
nand U37009 (N_37009,N_33165,N_33447);
nand U37010 (N_37010,N_33064,N_33971);
nand U37011 (N_37011,N_34182,N_32504);
nand U37012 (N_37012,N_32692,N_32873);
xnor U37013 (N_37013,N_34236,N_32698);
nor U37014 (N_37014,N_33467,N_34667);
or U37015 (N_37015,N_33649,N_33293);
nor U37016 (N_37016,N_33908,N_33618);
nand U37017 (N_37017,N_33142,N_33323);
or U37018 (N_37018,N_33398,N_34829);
xor U37019 (N_37019,N_33698,N_34541);
or U37020 (N_37020,N_34690,N_33840);
and U37021 (N_37021,N_33843,N_33026);
nor U37022 (N_37022,N_32500,N_34478);
or U37023 (N_37023,N_34924,N_34288);
or U37024 (N_37024,N_33091,N_32643);
and U37025 (N_37025,N_32624,N_34527);
nor U37026 (N_37026,N_33010,N_34259);
nand U37027 (N_37027,N_33620,N_34559);
or U37028 (N_37028,N_33032,N_33344);
or U37029 (N_37029,N_33736,N_34251);
nor U37030 (N_37030,N_32894,N_32867);
or U37031 (N_37031,N_34585,N_34879);
nand U37032 (N_37032,N_34864,N_34098);
nor U37033 (N_37033,N_34206,N_33893);
and U37034 (N_37034,N_34417,N_33694);
nand U37035 (N_37035,N_33483,N_34185);
and U37036 (N_37036,N_34835,N_34938);
and U37037 (N_37037,N_33296,N_34086);
nor U37038 (N_37038,N_33127,N_34207);
nand U37039 (N_37039,N_34064,N_32881);
or U37040 (N_37040,N_33517,N_33287);
and U37041 (N_37041,N_33282,N_33151);
or U37042 (N_37042,N_32970,N_34873);
nor U37043 (N_37043,N_34614,N_32756);
nand U37044 (N_37044,N_33427,N_33328);
or U37045 (N_37045,N_33744,N_32969);
xnor U37046 (N_37046,N_32823,N_33114);
nand U37047 (N_37047,N_32859,N_34218);
nor U37048 (N_37048,N_33440,N_33541);
xor U37049 (N_37049,N_32727,N_32651);
nor U37050 (N_37050,N_34094,N_32682);
nor U37051 (N_37051,N_34632,N_32662);
and U37052 (N_37052,N_32575,N_34351);
nor U37053 (N_37053,N_34908,N_33707);
and U37054 (N_37054,N_33896,N_32967);
and U37055 (N_37055,N_32694,N_33911);
nand U37056 (N_37056,N_34424,N_33509);
and U37057 (N_37057,N_32754,N_32842);
or U37058 (N_37058,N_34549,N_32766);
nand U37059 (N_37059,N_33056,N_34206);
nand U37060 (N_37060,N_32628,N_34071);
nor U37061 (N_37061,N_33964,N_34166);
nor U37062 (N_37062,N_33334,N_34185);
and U37063 (N_37063,N_33885,N_33392);
nand U37064 (N_37064,N_33722,N_33846);
nor U37065 (N_37065,N_33846,N_34784);
and U37066 (N_37066,N_33710,N_34290);
nor U37067 (N_37067,N_33428,N_34180);
and U37068 (N_37068,N_33950,N_33593);
nor U37069 (N_37069,N_34718,N_33347);
or U37070 (N_37070,N_32700,N_33926);
or U37071 (N_37071,N_33913,N_33030);
nand U37072 (N_37072,N_32760,N_34078);
nand U37073 (N_37073,N_34150,N_34078);
nor U37074 (N_37074,N_34574,N_33471);
nor U37075 (N_37075,N_33479,N_33818);
nor U37076 (N_37076,N_34932,N_33329);
and U37077 (N_37077,N_33078,N_34382);
nand U37078 (N_37078,N_32734,N_33956);
and U37079 (N_37079,N_33285,N_33673);
and U37080 (N_37080,N_33115,N_33366);
nor U37081 (N_37081,N_34416,N_33425);
nand U37082 (N_37082,N_34977,N_33103);
and U37083 (N_37083,N_34269,N_33147);
nand U37084 (N_37084,N_33106,N_34033);
nor U37085 (N_37085,N_32703,N_33042);
nand U37086 (N_37086,N_33975,N_34844);
xor U37087 (N_37087,N_33803,N_33541);
nand U37088 (N_37088,N_33813,N_32838);
or U37089 (N_37089,N_34974,N_34611);
or U37090 (N_37090,N_34028,N_32523);
and U37091 (N_37091,N_33564,N_33346);
nand U37092 (N_37092,N_32632,N_34500);
and U37093 (N_37093,N_34231,N_33087);
nor U37094 (N_37094,N_32671,N_32573);
nor U37095 (N_37095,N_34054,N_34130);
nor U37096 (N_37096,N_33786,N_34061);
or U37097 (N_37097,N_34241,N_33665);
or U37098 (N_37098,N_34138,N_33141);
or U37099 (N_37099,N_33407,N_34381);
and U37100 (N_37100,N_34705,N_34460);
nor U37101 (N_37101,N_34972,N_33813);
xor U37102 (N_37102,N_34192,N_32857);
xnor U37103 (N_37103,N_33436,N_32563);
nand U37104 (N_37104,N_34304,N_34152);
nand U37105 (N_37105,N_33957,N_34242);
nand U37106 (N_37106,N_34361,N_34682);
nor U37107 (N_37107,N_34236,N_34521);
xor U37108 (N_37108,N_33957,N_34255);
or U37109 (N_37109,N_34365,N_34176);
nor U37110 (N_37110,N_34060,N_33949);
and U37111 (N_37111,N_33266,N_33524);
nand U37112 (N_37112,N_33231,N_32613);
or U37113 (N_37113,N_32989,N_34242);
and U37114 (N_37114,N_34304,N_33476);
nand U37115 (N_37115,N_32964,N_33995);
nand U37116 (N_37116,N_33510,N_33768);
and U37117 (N_37117,N_34691,N_33855);
xor U37118 (N_37118,N_33502,N_33677);
nor U37119 (N_37119,N_32976,N_34292);
or U37120 (N_37120,N_33170,N_34779);
or U37121 (N_37121,N_32687,N_34614);
or U37122 (N_37122,N_34893,N_33340);
or U37123 (N_37123,N_32808,N_33628);
nor U37124 (N_37124,N_33999,N_32714);
nand U37125 (N_37125,N_34232,N_34652);
or U37126 (N_37126,N_33255,N_33440);
nor U37127 (N_37127,N_34244,N_34266);
xor U37128 (N_37128,N_34757,N_33569);
or U37129 (N_37129,N_34899,N_34660);
and U37130 (N_37130,N_34239,N_33082);
or U37131 (N_37131,N_33494,N_34854);
or U37132 (N_37132,N_33829,N_32810);
and U37133 (N_37133,N_32842,N_33301);
and U37134 (N_37134,N_34006,N_34860);
xor U37135 (N_37135,N_34022,N_33131);
nor U37136 (N_37136,N_33850,N_33413);
nor U37137 (N_37137,N_33457,N_33918);
and U37138 (N_37138,N_34932,N_33081);
or U37139 (N_37139,N_34785,N_33324);
nand U37140 (N_37140,N_33237,N_34227);
nand U37141 (N_37141,N_34502,N_33499);
nand U37142 (N_37142,N_34260,N_33211);
or U37143 (N_37143,N_34145,N_33317);
and U37144 (N_37144,N_32747,N_32666);
nor U37145 (N_37145,N_33961,N_34756);
or U37146 (N_37146,N_32595,N_34562);
and U37147 (N_37147,N_34815,N_33889);
and U37148 (N_37148,N_33755,N_32531);
nor U37149 (N_37149,N_33229,N_32529);
nand U37150 (N_37150,N_34657,N_33714);
nor U37151 (N_37151,N_33949,N_32662);
nor U37152 (N_37152,N_34133,N_34428);
nand U37153 (N_37153,N_33287,N_32932);
xor U37154 (N_37154,N_32509,N_32767);
nor U37155 (N_37155,N_32996,N_33591);
and U37156 (N_37156,N_32506,N_33547);
and U37157 (N_37157,N_34401,N_34826);
nor U37158 (N_37158,N_32767,N_34871);
xnor U37159 (N_37159,N_34748,N_33753);
nand U37160 (N_37160,N_34347,N_33996);
nor U37161 (N_37161,N_32973,N_34718);
or U37162 (N_37162,N_34428,N_32754);
xnor U37163 (N_37163,N_33140,N_32978);
xor U37164 (N_37164,N_34983,N_34780);
xor U37165 (N_37165,N_33197,N_33271);
and U37166 (N_37166,N_34016,N_34048);
and U37167 (N_37167,N_34015,N_34913);
nor U37168 (N_37168,N_34128,N_32842);
xnor U37169 (N_37169,N_34251,N_34918);
or U37170 (N_37170,N_33910,N_34784);
and U37171 (N_37171,N_33966,N_33382);
nand U37172 (N_37172,N_33902,N_33578);
and U37173 (N_37173,N_34255,N_33896);
nand U37174 (N_37174,N_34341,N_34138);
nor U37175 (N_37175,N_32791,N_33846);
and U37176 (N_37176,N_34049,N_34327);
nand U37177 (N_37177,N_34280,N_33434);
nand U37178 (N_37178,N_34593,N_32942);
or U37179 (N_37179,N_34174,N_34841);
nor U37180 (N_37180,N_33128,N_33426);
and U37181 (N_37181,N_34725,N_33005);
or U37182 (N_37182,N_33468,N_32972);
and U37183 (N_37183,N_34402,N_34200);
and U37184 (N_37184,N_34401,N_32764);
nand U37185 (N_37185,N_33913,N_33417);
nand U37186 (N_37186,N_33927,N_32804);
nor U37187 (N_37187,N_34241,N_33307);
nor U37188 (N_37188,N_34894,N_34846);
xor U37189 (N_37189,N_33400,N_33690);
or U37190 (N_37190,N_33058,N_34418);
and U37191 (N_37191,N_33118,N_34813);
xnor U37192 (N_37192,N_33013,N_33693);
or U37193 (N_37193,N_33292,N_33925);
nand U37194 (N_37194,N_34002,N_34263);
or U37195 (N_37195,N_34705,N_33025);
nor U37196 (N_37196,N_34214,N_34055);
nand U37197 (N_37197,N_32731,N_33366);
and U37198 (N_37198,N_34257,N_33957);
nand U37199 (N_37199,N_34033,N_33666);
and U37200 (N_37200,N_34359,N_32774);
or U37201 (N_37201,N_33921,N_33159);
nand U37202 (N_37202,N_32506,N_34722);
and U37203 (N_37203,N_33229,N_33376);
nand U37204 (N_37204,N_32735,N_34248);
or U37205 (N_37205,N_33274,N_34236);
nand U37206 (N_37206,N_33074,N_33292);
nor U37207 (N_37207,N_34824,N_34313);
xnor U37208 (N_37208,N_33912,N_34821);
or U37209 (N_37209,N_34880,N_32609);
and U37210 (N_37210,N_32622,N_34587);
nand U37211 (N_37211,N_34751,N_34102);
or U37212 (N_37212,N_33208,N_34301);
nand U37213 (N_37213,N_32905,N_32881);
and U37214 (N_37214,N_33046,N_33765);
and U37215 (N_37215,N_33943,N_34036);
xor U37216 (N_37216,N_34190,N_34159);
or U37217 (N_37217,N_32812,N_33918);
xor U37218 (N_37218,N_33238,N_33280);
nand U37219 (N_37219,N_34188,N_32693);
xnor U37220 (N_37220,N_33209,N_33365);
and U37221 (N_37221,N_33189,N_33558);
nand U37222 (N_37222,N_32893,N_32730);
xnor U37223 (N_37223,N_33007,N_32651);
xor U37224 (N_37224,N_34487,N_33552);
xnor U37225 (N_37225,N_33651,N_34751);
xor U37226 (N_37226,N_34015,N_34387);
nand U37227 (N_37227,N_33641,N_33877);
nor U37228 (N_37228,N_32848,N_33653);
and U37229 (N_37229,N_32592,N_33690);
or U37230 (N_37230,N_32707,N_33289);
and U37231 (N_37231,N_32927,N_34029);
xor U37232 (N_37232,N_33085,N_32739);
and U37233 (N_37233,N_34231,N_34211);
or U37234 (N_37234,N_33034,N_32942);
nor U37235 (N_37235,N_33170,N_34786);
nand U37236 (N_37236,N_33314,N_32803);
nor U37237 (N_37237,N_33244,N_34193);
nor U37238 (N_37238,N_32569,N_33091);
nand U37239 (N_37239,N_34461,N_33874);
xor U37240 (N_37240,N_34399,N_32862);
nand U37241 (N_37241,N_34793,N_34969);
xnor U37242 (N_37242,N_33506,N_34758);
xnor U37243 (N_37243,N_32863,N_33724);
nor U37244 (N_37244,N_34683,N_34005);
and U37245 (N_37245,N_33465,N_33751);
nor U37246 (N_37246,N_32541,N_33917);
nand U37247 (N_37247,N_34906,N_34119);
xor U37248 (N_37248,N_33338,N_32561);
nor U37249 (N_37249,N_34330,N_32806);
nor U37250 (N_37250,N_33159,N_32972);
and U37251 (N_37251,N_33865,N_33399);
or U37252 (N_37252,N_32764,N_32699);
or U37253 (N_37253,N_33920,N_34029);
or U37254 (N_37254,N_33631,N_34738);
nand U37255 (N_37255,N_32997,N_33021);
nor U37256 (N_37256,N_34034,N_33392);
xor U37257 (N_37257,N_34194,N_34700);
nand U37258 (N_37258,N_33079,N_33430);
nand U37259 (N_37259,N_34367,N_32614);
nor U37260 (N_37260,N_34236,N_32608);
nor U37261 (N_37261,N_33999,N_34357);
and U37262 (N_37262,N_33171,N_33351);
nor U37263 (N_37263,N_34528,N_34962);
and U37264 (N_37264,N_33970,N_33252);
xnor U37265 (N_37265,N_33198,N_33805);
xor U37266 (N_37266,N_34081,N_33050);
nor U37267 (N_37267,N_34230,N_32588);
nand U37268 (N_37268,N_34319,N_32874);
xnor U37269 (N_37269,N_34092,N_34679);
nand U37270 (N_37270,N_34450,N_33987);
nor U37271 (N_37271,N_33045,N_32910);
or U37272 (N_37272,N_32775,N_32989);
nor U37273 (N_37273,N_33217,N_34932);
or U37274 (N_37274,N_33352,N_33016);
or U37275 (N_37275,N_34114,N_32616);
xnor U37276 (N_37276,N_33545,N_34959);
nand U37277 (N_37277,N_34433,N_33964);
and U37278 (N_37278,N_32522,N_32932);
xnor U37279 (N_37279,N_33337,N_32903);
xor U37280 (N_37280,N_34416,N_33044);
nor U37281 (N_37281,N_33685,N_34793);
or U37282 (N_37282,N_34622,N_32737);
nand U37283 (N_37283,N_34065,N_34969);
and U37284 (N_37284,N_32705,N_34735);
nand U37285 (N_37285,N_32923,N_34398);
nand U37286 (N_37286,N_32631,N_33844);
nor U37287 (N_37287,N_33051,N_34251);
xnor U37288 (N_37288,N_33653,N_33941);
xnor U37289 (N_37289,N_32738,N_34723);
nor U37290 (N_37290,N_33787,N_33449);
or U37291 (N_37291,N_34813,N_32662);
nor U37292 (N_37292,N_34071,N_34658);
xnor U37293 (N_37293,N_34703,N_33497);
nand U37294 (N_37294,N_33732,N_33811);
nand U37295 (N_37295,N_34852,N_33314);
xnor U37296 (N_37296,N_33312,N_33548);
nand U37297 (N_37297,N_33202,N_33920);
xnor U37298 (N_37298,N_34715,N_33760);
and U37299 (N_37299,N_33376,N_34443);
xnor U37300 (N_37300,N_33205,N_33178);
nor U37301 (N_37301,N_32758,N_33460);
nor U37302 (N_37302,N_34858,N_33568);
and U37303 (N_37303,N_33336,N_33461);
and U37304 (N_37304,N_34527,N_33007);
nand U37305 (N_37305,N_34577,N_33232);
and U37306 (N_37306,N_34381,N_33883);
or U37307 (N_37307,N_33854,N_33053);
and U37308 (N_37308,N_32571,N_32907);
xnor U37309 (N_37309,N_34242,N_34760);
xnor U37310 (N_37310,N_34231,N_34841);
and U37311 (N_37311,N_34495,N_34420);
and U37312 (N_37312,N_33959,N_33335);
nor U37313 (N_37313,N_33929,N_34757);
xor U37314 (N_37314,N_34762,N_33438);
nor U37315 (N_37315,N_33746,N_33417);
and U37316 (N_37316,N_33276,N_34508);
nor U37317 (N_37317,N_34560,N_33549);
or U37318 (N_37318,N_33802,N_33614);
and U37319 (N_37319,N_32920,N_32698);
nand U37320 (N_37320,N_33419,N_32734);
or U37321 (N_37321,N_34819,N_34934);
nor U37322 (N_37322,N_34039,N_33744);
nand U37323 (N_37323,N_33153,N_34757);
xor U37324 (N_37324,N_33581,N_32748);
xor U37325 (N_37325,N_34441,N_34423);
xor U37326 (N_37326,N_32699,N_33697);
nand U37327 (N_37327,N_34841,N_34738);
nor U37328 (N_37328,N_33460,N_33950);
and U37329 (N_37329,N_34124,N_32884);
xnor U37330 (N_37330,N_34068,N_32879);
and U37331 (N_37331,N_32770,N_34329);
nand U37332 (N_37332,N_32531,N_32561);
nor U37333 (N_37333,N_32567,N_34001);
nand U37334 (N_37334,N_32747,N_34474);
nor U37335 (N_37335,N_33945,N_34666);
or U37336 (N_37336,N_33949,N_33937);
or U37337 (N_37337,N_34277,N_33492);
xor U37338 (N_37338,N_34259,N_34971);
nor U37339 (N_37339,N_32524,N_34019);
xor U37340 (N_37340,N_33320,N_33156);
xor U37341 (N_37341,N_33960,N_34138);
or U37342 (N_37342,N_33314,N_33634);
xor U37343 (N_37343,N_34764,N_34655);
or U37344 (N_37344,N_32534,N_34349);
nor U37345 (N_37345,N_33609,N_34503);
nor U37346 (N_37346,N_34537,N_32677);
and U37347 (N_37347,N_33392,N_34588);
and U37348 (N_37348,N_34658,N_32928);
nand U37349 (N_37349,N_34411,N_34423);
and U37350 (N_37350,N_33583,N_32911);
or U37351 (N_37351,N_33716,N_34285);
nor U37352 (N_37352,N_34921,N_32960);
and U37353 (N_37353,N_32575,N_32825);
xnor U37354 (N_37354,N_34493,N_32885);
or U37355 (N_37355,N_33867,N_34179);
nand U37356 (N_37356,N_33629,N_34839);
and U37357 (N_37357,N_32721,N_33651);
nand U37358 (N_37358,N_34103,N_34870);
and U37359 (N_37359,N_33524,N_32517);
or U37360 (N_37360,N_33999,N_34183);
xnor U37361 (N_37361,N_34957,N_32525);
and U37362 (N_37362,N_34256,N_33690);
or U37363 (N_37363,N_34568,N_34070);
nand U37364 (N_37364,N_34887,N_32871);
and U37365 (N_37365,N_32996,N_33830);
nor U37366 (N_37366,N_34439,N_34066);
or U37367 (N_37367,N_32979,N_34279);
xnor U37368 (N_37368,N_33838,N_34741);
xnor U37369 (N_37369,N_32788,N_32731);
nand U37370 (N_37370,N_33061,N_33343);
nor U37371 (N_37371,N_34081,N_34634);
nand U37372 (N_37372,N_33748,N_34007);
nand U37373 (N_37373,N_33336,N_33735);
xor U37374 (N_37374,N_33794,N_33038);
or U37375 (N_37375,N_32956,N_32550);
and U37376 (N_37376,N_33282,N_34187);
nor U37377 (N_37377,N_32532,N_34759);
nor U37378 (N_37378,N_34670,N_34364);
or U37379 (N_37379,N_33605,N_33160);
xnor U37380 (N_37380,N_33525,N_33520);
xor U37381 (N_37381,N_33038,N_32828);
xor U37382 (N_37382,N_33224,N_34759);
xnor U37383 (N_37383,N_32565,N_34884);
and U37384 (N_37384,N_33479,N_33809);
and U37385 (N_37385,N_33399,N_33342);
nand U37386 (N_37386,N_33709,N_32592);
and U37387 (N_37387,N_32844,N_34093);
or U37388 (N_37388,N_33983,N_32870);
nand U37389 (N_37389,N_33228,N_32700);
and U37390 (N_37390,N_33786,N_33300);
xor U37391 (N_37391,N_33848,N_34309);
xnor U37392 (N_37392,N_34273,N_33622);
nand U37393 (N_37393,N_33812,N_32874);
or U37394 (N_37394,N_32789,N_33741);
xnor U37395 (N_37395,N_33005,N_32820);
xor U37396 (N_37396,N_33914,N_33260);
and U37397 (N_37397,N_34701,N_33469);
xnor U37398 (N_37398,N_34225,N_34480);
nand U37399 (N_37399,N_32830,N_34278);
nand U37400 (N_37400,N_32555,N_34245);
nand U37401 (N_37401,N_33245,N_34825);
nor U37402 (N_37402,N_34082,N_33876);
nor U37403 (N_37403,N_34689,N_34729);
and U37404 (N_37404,N_33931,N_33731);
or U37405 (N_37405,N_32773,N_34209);
and U37406 (N_37406,N_32524,N_32730);
and U37407 (N_37407,N_34190,N_33630);
or U37408 (N_37408,N_33960,N_32510);
and U37409 (N_37409,N_33241,N_34055);
nor U37410 (N_37410,N_33049,N_34756);
and U37411 (N_37411,N_32828,N_34578);
xnor U37412 (N_37412,N_33196,N_34102);
xor U37413 (N_37413,N_34651,N_33929);
and U37414 (N_37414,N_34147,N_33216);
nand U37415 (N_37415,N_34504,N_34945);
xnor U37416 (N_37416,N_33644,N_33673);
or U37417 (N_37417,N_33191,N_33517);
xor U37418 (N_37418,N_34546,N_34324);
xor U37419 (N_37419,N_34016,N_34297);
nand U37420 (N_37420,N_34499,N_34428);
nand U37421 (N_37421,N_33447,N_34711);
xor U37422 (N_37422,N_33015,N_32731);
xor U37423 (N_37423,N_34126,N_32550);
nor U37424 (N_37424,N_34157,N_33974);
nand U37425 (N_37425,N_33634,N_32502);
nor U37426 (N_37426,N_33595,N_33022);
xnor U37427 (N_37427,N_34285,N_34730);
xnor U37428 (N_37428,N_34822,N_33314);
and U37429 (N_37429,N_33216,N_34780);
and U37430 (N_37430,N_32895,N_33216);
and U37431 (N_37431,N_33667,N_34891);
nor U37432 (N_37432,N_32816,N_33480);
nand U37433 (N_37433,N_33701,N_32858);
nor U37434 (N_37434,N_33725,N_32972);
xnor U37435 (N_37435,N_34040,N_34497);
nand U37436 (N_37436,N_34704,N_34574);
or U37437 (N_37437,N_32993,N_33538);
nor U37438 (N_37438,N_33115,N_32981);
nor U37439 (N_37439,N_33357,N_34330);
nor U37440 (N_37440,N_34093,N_34257);
nand U37441 (N_37441,N_32825,N_32913);
and U37442 (N_37442,N_33480,N_33880);
nand U37443 (N_37443,N_34059,N_34277);
or U37444 (N_37444,N_32823,N_33390);
or U37445 (N_37445,N_34104,N_34328);
and U37446 (N_37446,N_32709,N_33632);
and U37447 (N_37447,N_34478,N_34218);
and U37448 (N_37448,N_32915,N_33898);
and U37449 (N_37449,N_34498,N_32624);
nand U37450 (N_37450,N_32794,N_32757);
or U37451 (N_37451,N_32819,N_32640);
and U37452 (N_37452,N_34790,N_33507);
and U37453 (N_37453,N_33552,N_32707);
nand U37454 (N_37454,N_34413,N_33609);
nand U37455 (N_37455,N_34995,N_33183);
or U37456 (N_37456,N_34216,N_34173);
and U37457 (N_37457,N_33961,N_33526);
xor U37458 (N_37458,N_34156,N_32838);
nand U37459 (N_37459,N_34617,N_33890);
nand U37460 (N_37460,N_34201,N_33352);
and U37461 (N_37461,N_34643,N_32715);
nor U37462 (N_37462,N_33080,N_34775);
nor U37463 (N_37463,N_34649,N_34286);
or U37464 (N_37464,N_33544,N_34501);
nand U37465 (N_37465,N_34380,N_32915);
nor U37466 (N_37466,N_32559,N_33882);
nand U37467 (N_37467,N_32880,N_33986);
nand U37468 (N_37468,N_34842,N_34098);
or U37469 (N_37469,N_33869,N_33008);
xor U37470 (N_37470,N_33836,N_33362);
and U37471 (N_37471,N_33914,N_34708);
and U37472 (N_37472,N_33423,N_34784);
or U37473 (N_37473,N_34490,N_32831);
nand U37474 (N_37474,N_33860,N_34104);
nand U37475 (N_37475,N_33132,N_32963);
nor U37476 (N_37476,N_33590,N_34087);
and U37477 (N_37477,N_32756,N_34365);
nand U37478 (N_37478,N_34171,N_33422);
xor U37479 (N_37479,N_33687,N_34522);
xnor U37480 (N_37480,N_34988,N_33966);
or U37481 (N_37481,N_34822,N_34343);
nand U37482 (N_37482,N_34427,N_33099);
and U37483 (N_37483,N_33134,N_34328);
or U37484 (N_37484,N_34587,N_34035);
xnor U37485 (N_37485,N_32837,N_33514);
nand U37486 (N_37486,N_34170,N_32651);
nand U37487 (N_37487,N_34846,N_34513);
or U37488 (N_37488,N_34006,N_32806);
and U37489 (N_37489,N_33665,N_34423);
or U37490 (N_37490,N_34599,N_32878);
nor U37491 (N_37491,N_32628,N_34916);
xnor U37492 (N_37492,N_32926,N_34409);
nand U37493 (N_37493,N_34005,N_33968);
or U37494 (N_37494,N_34078,N_34720);
nand U37495 (N_37495,N_34085,N_34044);
nand U37496 (N_37496,N_33051,N_34037);
or U37497 (N_37497,N_33427,N_33672);
nand U37498 (N_37498,N_33313,N_34985);
or U37499 (N_37499,N_32723,N_32809);
and U37500 (N_37500,N_35501,N_35878);
or U37501 (N_37501,N_35049,N_36805);
nand U37502 (N_37502,N_35992,N_35456);
nor U37503 (N_37503,N_37254,N_35660);
xor U37504 (N_37504,N_35875,N_36452);
and U37505 (N_37505,N_37287,N_36754);
nand U37506 (N_37506,N_35328,N_37360);
xnor U37507 (N_37507,N_35154,N_35936);
or U37508 (N_37508,N_35063,N_37456);
and U37509 (N_37509,N_36009,N_36467);
or U37510 (N_37510,N_36546,N_37402);
nand U37511 (N_37511,N_37374,N_36572);
xor U37512 (N_37512,N_36534,N_37261);
nand U37513 (N_37513,N_35655,N_35443);
nor U37514 (N_37514,N_36547,N_36428);
nor U37515 (N_37515,N_36336,N_35712);
or U37516 (N_37516,N_36440,N_36111);
xnor U37517 (N_37517,N_35953,N_35293);
xor U37518 (N_37518,N_35637,N_35190);
and U37519 (N_37519,N_37293,N_36846);
xnor U37520 (N_37520,N_35414,N_36792);
xnor U37521 (N_37521,N_36594,N_35177);
nand U37522 (N_37522,N_36222,N_37325);
nand U37523 (N_37523,N_36512,N_35740);
xor U37524 (N_37524,N_35096,N_36983);
and U37525 (N_37525,N_36378,N_35641);
xor U37526 (N_37526,N_36849,N_35382);
and U37527 (N_37527,N_37055,N_37314);
or U37528 (N_37528,N_37337,N_35839);
nor U37529 (N_37529,N_35672,N_37089);
nand U37530 (N_37530,N_36901,N_35753);
or U37531 (N_37531,N_35691,N_35990);
xor U37532 (N_37532,N_37058,N_36684);
nand U37533 (N_37533,N_35576,N_36844);
nor U37534 (N_37534,N_35174,N_36479);
or U37535 (N_37535,N_37297,N_36880);
nand U37536 (N_37536,N_35368,N_36298);
nor U37537 (N_37537,N_36242,N_35998);
and U37538 (N_37538,N_35013,N_36410);
xor U37539 (N_37539,N_37029,N_36851);
and U37540 (N_37540,N_37198,N_37018);
nand U37541 (N_37541,N_35694,N_36885);
xor U37542 (N_37542,N_36682,N_36184);
and U37543 (N_37543,N_36550,N_36231);
xnor U37544 (N_37544,N_37171,N_35789);
nor U37545 (N_37545,N_37070,N_36155);
or U37546 (N_37546,N_35234,N_35794);
nor U37547 (N_37547,N_35250,N_37117);
xnor U37548 (N_37548,N_35405,N_37017);
or U37549 (N_37549,N_36059,N_36913);
xnor U37550 (N_37550,N_37066,N_37243);
nor U37551 (N_37551,N_35764,N_37026);
xnor U37552 (N_37552,N_36283,N_35937);
nor U37553 (N_37553,N_36940,N_36210);
xnor U37554 (N_37554,N_35522,N_35976);
nor U37555 (N_37555,N_37447,N_37344);
and U37556 (N_37556,N_36032,N_36074);
or U37557 (N_37557,N_36172,N_36267);
nor U37558 (N_37558,N_35084,N_36904);
nand U37559 (N_37559,N_37274,N_35244);
nand U37560 (N_37560,N_37087,N_35273);
nor U37561 (N_37561,N_36284,N_37386);
nor U37562 (N_37562,N_35553,N_36365);
xnor U37563 (N_37563,N_35578,N_37049);
nand U37564 (N_37564,N_37399,N_36102);
xnor U37565 (N_37565,N_36384,N_35823);
nand U37566 (N_37566,N_36946,N_36789);
nand U37567 (N_37567,N_37455,N_35934);
and U37568 (N_37568,N_37033,N_35149);
xnor U37569 (N_37569,N_35054,N_36943);
nor U37570 (N_37570,N_37236,N_35082);
nand U37571 (N_37571,N_36625,N_35667);
nor U37572 (N_37572,N_35502,N_37179);
nor U37573 (N_37573,N_35097,N_35530);
xnor U37574 (N_37574,N_36918,N_35706);
nor U37575 (N_37575,N_35949,N_36910);
or U37576 (N_37576,N_35886,N_36592);
nor U37577 (N_37577,N_37301,N_36709);
nor U37578 (N_37578,N_36543,N_36109);
nand U37579 (N_37579,N_35125,N_35735);
nand U37580 (N_37580,N_36502,N_35561);
xnor U37581 (N_37581,N_36574,N_37030);
and U37582 (N_37582,N_35591,N_35338);
or U37583 (N_37583,N_37095,N_36873);
nand U37584 (N_37584,N_37013,N_37356);
nand U37585 (N_37585,N_36416,N_36016);
and U37586 (N_37586,N_37183,N_36066);
or U37587 (N_37587,N_36388,N_35803);
nand U37588 (N_37588,N_35301,N_36786);
and U37589 (N_37589,N_35046,N_36215);
and U37590 (N_37590,N_36887,N_36347);
or U37591 (N_37591,N_36319,N_35281);
xor U37592 (N_37592,N_37253,N_35772);
xor U37593 (N_37593,N_37315,N_35164);
nor U37594 (N_37594,N_36176,N_35972);
xnor U37595 (N_37595,N_36957,N_36049);
nor U37596 (N_37596,N_36180,N_35123);
xor U37597 (N_37597,N_35081,N_37387);
and U37598 (N_37598,N_36586,N_35243);
and U37599 (N_37599,N_37383,N_36896);
nand U37600 (N_37600,N_35488,N_37372);
nor U37601 (N_37601,N_35138,N_35478);
or U37602 (N_37602,N_35342,N_37234);
nand U37603 (N_37603,N_35151,N_36361);
nand U37604 (N_37604,N_35284,N_36251);
or U37605 (N_37605,N_35588,N_35736);
and U37606 (N_37606,N_37318,N_37457);
and U37607 (N_37607,N_36099,N_35481);
nand U37608 (N_37608,N_35091,N_37047);
or U37609 (N_37609,N_36316,N_35978);
or U37610 (N_37610,N_36984,N_36480);
and U37611 (N_37611,N_36633,N_36986);
or U37612 (N_37612,N_37131,N_36152);
or U37613 (N_37613,N_35716,N_36532);
or U37614 (N_37614,N_36490,N_36756);
xnor U37615 (N_37615,N_35459,N_36446);
and U37616 (N_37616,N_36076,N_36667);
and U37617 (N_37617,N_35272,N_35916);
or U37618 (N_37618,N_36856,N_35348);
or U37619 (N_37619,N_35639,N_37227);
and U37620 (N_37620,N_37078,N_36127);
nor U37621 (N_37621,N_36160,N_36411);
nand U37622 (N_37622,N_35506,N_35683);
xnor U37623 (N_37623,N_36517,N_36657);
and U37624 (N_37624,N_37275,N_37186);
and U37625 (N_37625,N_36954,N_35027);
and U37626 (N_37626,N_35634,N_36005);
or U37627 (N_37627,N_35836,N_35408);
xnor U37628 (N_37628,N_37453,N_36393);
and U37629 (N_37629,N_37040,N_35323);
nor U37630 (N_37630,N_36370,N_35883);
and U37631 (N_37631,N_36023,N_36084);
and U37632 (N_37632,N_35783,N_36335);
nor U37633 (N_37633,N_35782,N_35833);
nor U37634 (N_37634,N_35673,N_35665);
xor U37635 (N_37635,N_35028,N_36027);
and U37636 (N_37636,N_35067,N_36513);
and U37637 (N_37637,N_35142,N_37022);
or U37638 (N_37638,N_37020,N_35445);
nand U37639 (N_37639,N_36566,N_36068);
and U37640 (N_37640,N_35322,N_36130);
xor U37641 (N_37641,N_35264,N_35024);
and U37642 (N_37642,N_36445,N_36292);
nand U37643 (N_37643,N_35423,N_35601);
or U37644 (N_37644,N_36585,N_36028);
nand U37645 (N_37645,N_35629,N_37438);
and U37646 (N_37646,N_37223,N_35043);
or U37647 (N_37647,N_36404,N_36529);
xor U37648 (N_37648,N_36829,N_36795);
and U37649 (N_37649,N_36002,N_36510);
and U37650 (N_37650,N_37061,N_36826);
or U37651 (N_37651,N_37146,N_35044);
or U37652 (N_37652,N_35473,N_36746);
nor U37653 (N_37653,N_35714,N_36649);
nand U37654 (N_37654,N_35065,N_35625);
or U37655 (N_37655,N_35393,N_35179);
or U37656 (N_37656,N_36342,N_35677);
nand U37657 (N_37657,N_35367,N_36471);
or U37658 (N_37658,N_36775,N_36807);
or U37659 (N_37659,N_35358,N_35023);
or U37660 (N_37660,N_37357,N_36836);
nand U37661 (N_37661,N_36634,N_36401);
or U37662 (N_37662,N_35713,N_35186);
and U37663 (N_37663,N_36724,N_36992);
nor U37664 (N_37664,N_36080,N_36942);
and U37665 (N_37665,N_37039,N_37370);
or U37666 (N_37666,N_37333,N_35104);
nand U37667 (N_37667,N_35214,N_35416);
and U37668 (N_37668,N_36168,N_35858);
and U37669 (N_37669,N_35490,N_35732);
nor U37670 (N_37670,N_36647,N_36728);
nor U37671 (N_37671,N_35961,N_35757);
nor U37672 (N_37672,N_36493,N_36835);
and U37673 (N_37673,N_35194,N_37232);
nor U37674 (N_37674,N_36619,N_37156);
or U37675 (N_37675,N_35633,N_36762);
or U37676 (N_37676,N_35837,N_37401);
and U37677 (N_37677,N_35927,N_36922);
or U37678 (N_37678,N_36266,N_35958);
nor U37679 (N_37679,N_36320,N_36958);
xor U37680 (N_37680,N_36978,N_37273);
nor U37681 (N_37681,N_35627,N_35769);
or U37682 (N_37682,N_37104,N_36987);
or U37683 (N_37683,N_37365,N_36257);
nor U37684 (N_37684,N_37221,N_35771);
and U37685 (N_37685,N_36816,N_36469);
or U37686 (N_37686,N_37220,N_37099);
and U37687 (N_37687,N_35465,N_36607);
xnor U37688 (N_37688,N_37413,N_35640);
and U37689 (N_37689,N_36663,N_35040);
xor U37690 (N_37690,N_36389,N_37176);
xor U37691 (N_37691,N_37385,N_37340);
nand U37692 (N_37692,N_36899,N_37391);
xor U37693 (N_37693,N_35954,N_37027);
nor U37694 (N_37694,N_35289,N_35513);
nand U37695 (N_37695,N_36761,N_35538);
nand U37696 (N_37696,N_36845,N_36536);
and U37697 (N_37697,N_36259,N_36610);
xnor U37698 (N_37698,N_35910,N_36577);
and U37699 (N_37699,N_35652,N_35185);
and U37700 (N_37700,N_35122,N_37244);
and U37701 (N_37701,N_36293,N_35434);
or U37702 (N_37702,N_36595,N_36148);
and U37703 (N_37703,N_35071,N_36772);
nand U37704 (N_37704,N_35425,N_35666);
xor U37705 (N_37705,N_36631,N_36158);
nand U37706 (N_37706,N_36092,N_35241);
xnor U37707 (N_37707,N_36057,N_37353);
nor U37708 (N_37708,N_35001,N_35285);
xnor U37709 (N_37709,N_36246,N_36900);
nor U37710 (N_37710,N_36011,N_36313);
nand U37711 (N_37711,N_35215,N_37369);
nand U37712 (N_37712,N_36993,N_35535);
nor U37713 (N_37713,N_35815,N_35008);
and U37714 (N_37714,N_36179,N_36110);
xor U37715 (N_37715,N_35150,N_35620);
or U37716 (N_37716,N_35623,N_37126);
or U37717 (N_37717,N_37120,N_35577);
nor U37718 (N_37718,N_35055,N_35507);
nand U37719 (N_37719,N_36650,N_35860);
nor U37720 (N_37720,N_36159,N_37488);
or U37721 (N_37721,N_36237,N_35569);
nor U37722 (N_37722,N_37125,N_37056);
or U37723 (N_37723,N_36914,N_35482);
nor U37724 (N_37724,N_35339,N_35240);
or U37725 (N_37725,N_36124,N_35221);
nor U37726 (N_37726,N_36424,N_35454);
xnor U37727 (N_37727,N_36858,N_37487);
or U37728 (N_37728,N_37317,N_35356);
nand U37729 (N_37729,N_36869,N_36980);
or U37730 (N_37730,N_36484,N_35907);
nand U37731 (N_37731,N_36483,N_36804);
or U37732 (N_37732,N_35995,N_36919);
xor U37733 (N_37733,N_35919,N_35187);
xnor U37734 (N_37734,N_35183,N_35156);
nor U37735 (N_37735,N_37113,N_36321);
nor U37736 (N_37736,N_35099,N_36421);
nand U37737 (N_37737,N_37000,N_35671);
nor U37738 (N_37738,N_36809,N_36225);
xnor U37739 (N_37739,N_35840,N_36056);
nand U37740 (N_37740,N_35231,N_36680);
nor U37741 (N_37741,N_37256,N_36010);
or U37742 (N_37742,N_35057,N_36422);
nor U37743 (N_37743,N_35543,N_35135);
nor U37744 (N_37744,N_36455,N_35257);
nor U37745 (N_37745,N_35074,N_37281);
nor U37746 (N_37746,N_36138,N_36275);
or U37747 (N_37747,N_37334,N_35778);
xor U37748 (N_37748,N_36596,N_35517);
xor U37749 (N_37749,N_37375,N_35102);
and U37750 (N_37750,N_36977,N_36258);
or U37751 (N_37751,N_37467,N_35238);
nor U37752 (N_37752,N_36812,N_35015);
or U37753 (N_37753,N_35011,N_35765);
nand U37754 (N_37754,N_37276,N_36306);
nor U37755 (N_37755,N_37139,N_35668);
nand U37756 (N_37756,N_35369,N_37187);
or U37757 (N_37757,N_35977,N_35030);
nand U37758 (N_37758,N_36202,N_35451);
and U37759 (N_37759,N_35426,N_37133);
nor U37760 (N_37760,N_36163,N_36438);
xor U37761 (N_37761,N_36831,N_36850);
xnor U37762 (N_37762,N_36832,N_37486);
or U37763 (N_37763,N_36398,N_36117);
or U37764 (N_37764,N_36509,N_36748);
nor U37765 (N_37765,N_37392,N_36432);
and U37766 (N_37766,N_36938,N_35471);
nand U37767 (N_37767,N_35754,N_37433);
nor U37768 (N_37768,N_37436,N_35440);
or U37769 (N_37769,N_37425,N_36119);
xor U37770 (N_37770,N_36195,N_37192);
and U37771 (N_37771,N_35755,N_37248);
nor U37772 (N_37772,N_35832,N_35497);
nor U37773 (N_37773,N_37212,N_36482);
or U37774 (N_37774,N_37440,N_37348);
and U37775 (N_37775,N_35865,N_36898);
nor U37776 (N_37776,N_36248,N_37366);
and U37777 (N_37777,N_35986,N_37045);
and U37778 (N_37778,N_36808,N_35882);
xnor U37779 (N_37779,N_35470,N_36055);
xnor U37780 (N_37780,N_35575,N_35290);
xnor U37781 (N_37781,N_35038,N_37382);
nand U37782 (N_37782,N_35618,N_35642);
nor U37783 (N_37783,N_36605,N_36396);
xnor U37784 (N_37784,N_35511,N_36722);
or U37785 (N_37785,N_36953,N_36192);
nand U37786 (N_37786,N_35029,N_36371);
or U37787 (N_37787,N_36095,N_36841);
nor U37788 (N_37788,N_37312,N_35255);
nor U37789 (N_37789,N_36311,N_37483);
and U37790 (N_37790,N_35495,N_35628);
xnor U37791 (N_37791,N_35559,N_37259);
nor U37792 (N_37792,N_36417,N_35321);
and U37793 (N_37793,N_35926,N_35377);
nand U37794 (N_37794,N_37480,N_35894);
nand U37795 (N_37795,N_35217,N_36329);
or U37796 (N_37796,N_35862,N_35945);
nand U37797 (N_37797,N_35076,N_35205);
nand U37798 (N_37798,N_36583,N_35831);
nor U37799 (N_37799,N_36046,N_36048);
xor U37800 (N_37800,N_36414,N_35996);
nand U37801 (N_37801,N_35311,N_36867);
nor U37802 (N_37802,N_36140,N_35020);
xnor U37803 (N_37803,N_35643,N_35848);
nor U37804 (N_37804,N_36305,N_36139);
nor U37805 (N_37805,N_36810,N_36956);
xnor U37806 (N_37806,N_35825,N_35093);
nor U37807 (N_37807,N_35401,N_36462);
or U37808 (N_37808,N_35702,N_36769);
nor U37809 (N_37809,N_36333,N_35903);
nand U37810 (N_37810,N_36862,N_35776);
nor U37811 (N_37811,N_35604,N_36357);
and U37812 (N_37812,N_35924,N_36656);
and U37813 (N_37813,N_37052,N_37485);
and U37814 (N_37814,N_36077,N_35647);
or U37815 (N_37815,N_37422,N_35347);
and U37816 (N_37816,N_35879,N_37410);
or U37817 (N_37817,N_37412,N_35376);
xor U37818 (N_37818,N_37294,N_37137);
nor U37819 (N_37819,N_35827,N_35133);
and U37820 (N_37820,N_36505,N_35058);
and U37821 (N_37821,N_35844,N_36271);
or U37822 (N_37822,N_37172,N_36475);
or U37823 (N_37823,N_36552,N_36064);
and U37824 (N_37824,N_36343,N_35457);
or U37825 (N_37825,N_36963,N_35876);
or U37826 (N_37826,N_37368,N_37199);
xor U37827 (N_37827,N_36129,N_36955);
and U37828 (N_37828,N_37124,N_35357);
xor U37829 (N_37829,N_37106,N_35994);
or U37830 (N_37830,N_36527,N_36995);
or U37831 (N_37831,N_36670,N_36638);
xnor U37832 (N_37832,N_36753,N_36137);
nand U37833 (N_37833,N_37466,N_37462);
nor U37834 (N_37834,N_37228,N_37147);
and U37835 (N_37835,N_35563,N_37381);
or U37836 (N_37836,N_35545,N_37477);
and U37837 (N_37837,N_35942,N_35514);
xnor U37838 (N_37838,N_37464,N_35370);
and U37839 (N_37839,N_36923,N_35959);
or U37840 (N_37840,N_35654,N_35867);
xnor U37841 (N_37841,N_35399,N_37128);
nand U37842 (N_37842,N_35315,N_35430);
and U37843 (N_37843,N_36972,N_36042);
nand U37844 (N_37844,N_35254,N_35365);
and U37845 (N_37845,N_36537,N_37307);
and U37846 (N_37846,N_37157,N_35303);
nor U37847 (N_37847,N_37028,N_37012);
and U37848 (N_37848,N_35944,N_37148);
nor U37849 (N_37849,N_35474,N_36823);
nand U37850 (N_37850,N_36228,N_37389);
nor U37851 (N_37851,N_36456,N_36058);
or U37852 (N_37852,N_35325,N_36830);
and U37853 (N_37853,N_37491,N_36413);
xnor U37854 (N_37854,N_36661,N_35230);
xor U37855 (N_37855,N_36576,N_37005);
nor U37856 (N_37856,N_36526,N_36133);
and U37857 (N_37857,N_36929,N_36701);
and U37858 (N_37858,N_37072,N_36582);
xnor U37859 (N_37859,N_35048,N_36544);
and U37860 (N_37860,N_35503,N_37063);
xor U37861 (N_37861,N_35178,N_35816);
or U37862 (N_37862,N_36403,N_35120);
nor U37863 (N_37863,N_36406,N_37398);
xor U37864 (N_37864,N_35790,N_36377);
nand U37865 (N_37865,N_37037,N_36698);
or U37866 (N_37866,N_35658,N_37135);
and U37867 (N_37867,N_37068,N_37100);
xnor U37868 (N_37868,N_35180,N_35010);
and U37869 (N_37869,N_37423,N_35873);
or U37870 (N_37870,N_36031,N_35251);
xnor U37871 (N_37871,N_36491,N_35220);
nor U37872 (N_37872,N_37308,N_36936);
xnor U37873 (N_37873,N_35870,N_35492);
nand U37874 (N_37874,N_36103,N_36535);
nand U37875 (N_37875,N_36557,N_36962);
or U37876 (N_37876,N_35664,N_37379);
or U37877 (N_37877,N_36330,N_35928);
xor U37878 (N_37878,N_35042,N_35302);
and U37879 (N_37879,N_36514,N_36603);
or U37880 (N_37880,N_35341,N_35610);
xnor U37881 (N_37881,N_35450,N_37160);
nand U37882 (N_37882,N_36508,N_36920);
and U37883 (N_37883,N_35419,N_35644);
xnor U37884 (N_37884,N_36883,N_35391);
and U37885 (N_37885,N_37323,N_35531);
xor U37886 (N_37886,N_35609,N_37154);
and U37887 (N_37887,N_36207,N_35512);
and U37888 (N_37888,N_36079,N_35971);
and U37889 (N_37889,N_35745,N_36038);
or U37890 (N_37890,N_36981,N_35314);
nand U37891 (N_37891,N_36397,N_37180);
and U37892 (N_37892,N_37222,N_36533);
and U37893 (N_37893,N_35760,N_36803);
and U37894 (N_37894,N_35016,N_36648);
nand U37895 (N_37895,N_37170,N_35005);
and U37896 (N_37896,N_35534,N_35022);
xnor U37897 (N_37897,N_35843,N_35869);
xor U37898 (N_37898,N_36782,N_35593);
xnor U37899 (N_37899,N_35116,N_36354);
and U37900 (N_37900,N_37065,N_35900);
xor U37901 (N_37901,N_36645,N_35520);
nor U37902 (N_37902,N_36615,N_35246);
and U37903 (N_37903,N_37409,N_35300);
nor U37904 (N_37904,N_35617,N_37107);
or U37905 (N_37905,N_37494,N_36538);
nor U37906 (N_37906,N_36857,N_36617);
xnor U37907 (N_37907,N_36798,N_35306);
nor U37908 (N_37908,N_35785,N_36249);
nand U37909 (N_37909,N_35568,N_37364);
xor U37910 (N_37910,N_35447,N_36771);
or U37911 (N_37911,N_35162,N_35761);
nand U37912 (N_37912,N_36628,N_36852);
nor U37913 (N_37913,N_36255,N_36262);
nor U37914 (N_37914,N_36945,N_35747);
nand U37915 (N_37915,N_37151,N_35859);
or U37916 (N_37916,N_35309,N_36345);
or U37917 (N_37917,N_35899,N_37255);
nor U37918 (N_37918,N_36036,N_35332);
and U37919 (N_37919,N_35547,N_35045);
and U37920 (N_37920,N_36496,N_37197);
or U37921 (N_37921,N_36646,N_36640);
nand U37922 (N_37922,N_35788,N_35235);
nor U37923 (N_37923,N_35441,N_35458);
nor U37924 (N_37924,N_35897,N_36518);
nand U37925 (N_37925,N_37109,N_35468);
and U37926 (N_37926,N_35117,N_35033);
and U37927 (N_37927,N_35312,N_36905);
xor U37928 (N_37928,N_36000,N_36004);
or U37929 (N_37929,N_36916,N_35948);
and U37930 (N_37930,N_36620,N_36608);
and U37931 (N_37931,N_35731,N_36530);
nand U37932 (N_37932,N_36463,N_36924);
or U37933 (N_37933,N_36501,N_37388);
or U37934 (N_37934,N_35494,N_36815);
or U37935 (N_37935,N_35619,N_35527);
or U37936 (N_37936,N_36276,N_36908);
and U37937 (N_37937,N_36244,N_35041);
xnor U37938 (N_37938,N_36928,N_35239);
xnor U37939 (N_37939,N_35508,N_35103);
nor U37940 (N_37940,N_35261,N_36691);
and U37941 (N_37941,N_35855,N_35227);
xnor U37942 (N_37942,N_36794,N_35153);
and U37943 (N_37943,N_36256,N_36156);
nand U37944 (N_37944,N_35612,N_35930);
or U37945 (N_37945,N_36128,N_35108);
and U37946 (N_37946,N_36553,N_37446);
or U37947 (N_37947,N_36551,N_36597);
or U37948 (N_37948,N_37418,N_36081);
and U37949 (N_37949,N_35518,N_36717);
nand U37950 (N_37950,N_37341,N_35931);
or U37951 (N_37951,N_35307,N_36265);
or U37952 (N_37952,N_36328,N_35337);
nand U37953 (N_37953,N_35955,N_35113);
nand U37954 (N_37954,N_36740,N_36211);
nand U37955 (N_37955,N_36374,N_36668);
and U37956 (N_37956,N_35586,N_35087);
or U37957 (N_37957,N_36126,N_36239);
and U37958 (N_37958,N_35722,N_35528);
or U37959 (N_37959,N_35463,N_37302);
or U37960 (N_37960,N_36190,N_35274);
nand U37961 (N_37961,N_36203,N_35266);
xor U37962 (N_37962,N_37240,N_36040);
nor U37963 (N_37963,N_36948,N_36886);
nand U37964 (N_37964,N_35824,N_35596);
or U37965 (N_37965,N_36870,N_36976);
and U37966 (N_37966,N_35509,N_35236);
or U37967 (N_37967,N_35319,N_36690);
xnor U37968 (N_37968,N_36712,N_37292);
nor U37969 (N_37969,N_36708,N_36863);
or U37970 (N_37970,N_35160,N_36768);
and U37971 (N_37971,N_35064,N_37326);
xor U37972 (N_37972,N_35709,N_36145);
nor U37973 (N_37973,N_36008,N_37075);
and U37974 (N_37974,N_35019,N_35678);
or U37975 (N_37975,N_36934,N_37437);
xor U37976 (N_37976,N_36704,N_37168);
or U37977 (N_37977,N_35085,N_36659);
and U37978 (N_37978,N_35820,N_35263);
nor U37979 (N_37979,N_36689,N_35397);
nor U37980 (N_37980,N_36442,N_36308);
xnor U37981 (N_37981,N_35805,N_35964);
nand U37982 (N_37982,N_37111,N_36162);
xnor U37983 (N_37983,N_35432,N_35810);
nor U37984 (N_37984,N_36776,N_35453);
or U37985 (N_37985,N_36729,N_35409);
nor U37986 (N_37986,N_35693,N_35940);
or U37987 (N_37987,N_37233,N_37114);
nor U37988 (N_37988,N_36895,N_35101);
and U37989 (N_37989,N_36499,N_35168);
and U37990 (N_37990,N_35602,N_35991);
or U37991 (N_37991,N_37134,N_36965);
nand U37992 (N_37992,N_36889,N_36664);
or U37993 (N_37993,N_35988,N_35562);
and U37994 (N_37994,N_36531,N_36083);
xor U37995 (N_37995,N_36627,N_36075);
xor U37996 (N_37996,N_35193,N_37451);
and U37997 (N_37997,N_37450,N_35202);
xor U37998 (N_37998,N_36189,N_36568);
xnor U37999 (N_37999,N_35830,N_35599);
nor U38000 (N_38000,N_35580,N_36121);
and U38001 (N_38001,N_36315,N_37144);
xor U38002 (N_38002,N_36476,N_37478);
or U38003 (N_38003,N_36318,N_37469);
or U38004 (N_38004,N_35885,N_37110);
nand U38005 (N_38005,N_35615,N_36487);
or U38006 (N_38006,N_35105,N_35390);
and U38007 (N_38007,N_36730,N_37059);
or U38008 (N_38008,N_36504,N_36695);
and U38009 (N_38009,N_36287,N_35184);
xor U38010 (N_38010,N_36497,N_36299);
xnor U38011 (N_38011,N_36274,N_35283);
nand U38012 (N_38012,N_36104,N_35963);
and U38013 (N_38013,N_35075,N_37130);
or U38014 (N_38014,N_35126,N_37143);
nor U38015 (N_38015,N_37214,N_36599);
nor U38016 (N_38016,N_36665,N_35410);
nor U38017 (N_38017,N_36261,N_35965);
xor U38018 (N_38018,N_35932,N_36584);
or U38019 (N_38019,N_36834,N_37286);
and U38020 (N_38020,N_36797,N_36216);
or U38021 (N_38021,N_36353,N_35427);
nand U38022 (N_38022,N_35587,N_35143);
or U38023 (N_38023,N_35649,N_36975);
or U38024 (N_38024,N_35326,N_36653);
nor U38025 (N_38025,N_37034,N_35389);
and U38026 (N_38026,N_36985,N_36383);
and U38027 (N_38027,N_37299,N_36521);
and U38028 (N_38028,N_35925,N_36473);
and U38029 (N_38029,N_36894,N_36279);
nor U38030 (N_38030,N_35717,N_37041);
nand U38031 (N_38031,N_36108,N_35051);
and U38032 (N_38032,N_36498,N_36988);
or U38033 (N_38033,N_36094,N_35475);
nor U38034 (N_38034,N_35224,N_35025);
xnor U38035 (N_38035,N_36777,N_37354);
xor U38036 (N_38036,N_36485,N_36604);
or U38037 (N_38037,N_36391,N_35871);
nor U38038 (N_38038,N_35216,N_37495);
xor U38039 (N_38039,N_36824,N_37430);
xnor U38040 (N_38040,N_36142,N_37088);
xor U38041 (N_38041,N_35504,N_37121);
nand U38042 (N_38042,N_35203,N_36593);
nor U38043 (N_38043,N_35404,N_36629);
nor U38044 (N_38044,N_36454,N_37439);
xor U38045 (N_38045,N_36486,N_35851);
or U38046 (N_38046,N_36655,N_37246);
nor U38047 (N_38047,N_37355,N_36500);
or U38048 (N_38048,N_36932,N_36478);
xor U38049 (N_38049,N_36018,N_37190);
and U38050 (N_38050,N_36718,N_36524);
xnor U38051 (N_38051,N_35139,N_35645);
and U38052 (N_38052,N_36441,N_36070);
nor U38053 (N_38053,N_37153,N_36314);
xnor U38054 (N_38054,N_35298,N_35519);
or U38055 (N_38055,N_35768,N_36495);
nor U38056 (N_38056,N_37400,N_35489);
or U38057 (N_38057,N_35464,N_35699);
nor U38058 (N_38058,N_36020,N_36738);
and U38059 (N_38059,N_36970,N_35191);
nand U38060 (N_38060,N_36296,N_35249);
or U38061 (N_38061,N_36833,N_37024);
or U38062 (N_38062,N_35491,N_36840);
and U38063 (N_38063,N_35477,N_36893);
nand U38064 (N_38064,N_37225,N_35774);
or U38065 (N_38065,N_37174,N_36426);
and U38066 (N_38066,N_35938,N_35291);
nand U38067 (N_38067,N_35962,N_36186);
xnor U38068 (N_38068,N_36523,N_35002);
nor U38069 (N_38069,N_35137,N_37102);
nor U38070 (N_38070,N_35841,N_35260);
and U38071 (N_38071,N_37295,N_35555);
xnor U38072 (N_38072,N_35539,N_36150);
or U38073 (N_38073,N_36519,N_36892);
xor U38074 (N_38074,N_36326,N_35812);
nor U38075 (N_38075,N_35868,N_36540);
or U38076 (N_38076,N_36096,N_37482);
nor U38077 (N_38077,N_36707,N_37169);
xor U38078 (N_38078,N_36906,N_37090);
xor U38079 (N_38079,N_36147,N_35554);
and U38080 (N_38080,N_35797,N_37008);
nor U38081 (N_38081,N_35983,N_36939);
or U38082 (N_38082,N_35159,N_35698);
or U38083 (N_38083,N_36811,N_36800);
or U38084 (N_38084,N_35838,N_35711);
or U38085 (N_38085,N_35305,N_35737);
nand U38086 (N_38086,N_36060,N_35756);
xor U38087 (N_38087,N_35429,N_35346);
and U38088 (N_38088,N_35182,N_37205);
and U38089 (N_38089,N_35455,N_37347);
xor U38090 (N_38090,N_35638,N_35741);
or U38091 (N_38091,N_35480,N_36624);
and U38092 (N_38092,N_36721,N_35072);
nor U38093 (N_38093,N_36613,N_37263);
xnor U38094 (N_38094,N_36412,N_37003);
and U38095 (N_38095,N_36364,N_35687);
nor U38096 (N_38096,N_35802,N_35222);
and U38097 (N_38097,N_35355,N_35526);
or U38098 (N_38098,N_36359,N_35877);
xor U38099 (N_38099,N_35158,N_36218);
nand U38100 (N_38100,N_36959,N_36884);
nor U38101 (N_38101,N_36012,N_35728);
nor U38102 (N_38102,N_35536,N_36658);
or U38103 (N_38103,N_35237,N_37460);
or U38104 (N_38104,N_37097,N_36881);
xor U38105 (N_38105,N_36644,N_35310);
nor U38106 (N_38106,N_37091,N_36488);
xnor U38107 (N_38107,N_36304,N_36285);
nand U38108 (N_38108,N_36755,N_37159);
nor U38109 (N_38109,N_35856,N_36091);
or U38110 (N_38110,N_35189,N_35493);
xnor U38111 (N_38111,N_35595,N_37152);
or U38112 (N_38112,N_35787,N_37285);
nand U38113 (N_38113,N_36144,N_35299);
xnor U38114 (N_38114,N_35516,N_35204);
and U38115 (N_38115,N_36164,N_36790);
xor U38116 (N_38116,N_35098,N_37417);
nor U38117 (N_38117,N_35228,N_37250);
nand U38118 (N_38118,N_36420,N_37441);
xor U38119 (N_38119,N_36146,N_37435);
nor U38120 (N_38120,N_35887,N_36107);
nor U38121 (N_38121,N_37284,N_36861);
or U38122 (N_38122,N_36199,N_37081);
nand U38123 (N_38123,N_35280,N_35373);
nand U38124 (N_38124,N_35594,N_36522);
or U38125 (N_38125,N_36072,N_36611);
or U38126 (N_38126,N_36209,N_35361);
or U38127 (N_38127,N_35669,N_35288);
nor U38128 (N_38128,N_36766,N_36864);
nor U38129 (N_38129,N_36859,N_35570);
or U38130 (N_38130,N_35380,N_35115);
nor U38131 (N_38131,N_36214,N_37394);
xnor U38132 (N_38132,N_36503,N_35791);
nand U38133 (N_38133,N_35026,N_35720);
and U38134 (N_38134,N_36726,N_36078);
nor U38135 (N_38135,N_37165,N_35210);
nor U38136 (N_38136,N_37378,N_37459);
and U38137 (N_38137,N_36101,N_36838);
nand U38138 (N_38138,N_36300,N_35050);
and U38139 (N_38139,N_36088,N_35060);
nand U38140 (N_38140,N_35066,N_35172);
xnor U38141 (N_38141,N_35857,N_36589);
nand U38142 (N_38142,N_35371,N_37231);
or U38143 (N_38143,N_37092,N_37031);
nor U38144 (N_38144,N_35541,N_36868);
and U38145 (N_38145,N_35917,N_36071);
and U38146 (N_38146,N_36431,N_35386);
or U38147 (N_38147,N_35375,N_37452);
xnor U38148 (N_38148,N_35866,N_37497);
xor U38149 (N_38149,N_37468,N_35487);
nor U38150 (N_38150,N_37342,N_36037);
or U38151 (N_38151,N_35792,N_36773);
nand U38152 (N_38152,N_35829,N_37443);
and U38153 (N_38153,N_36506,N_36710);
or U38154 (N_38154,N_35335,N_35021);
and U38155 (N_38155,N_35630,N_37331);
and U38156 (N_38156,N_35814,N_35056);
nor U38157 (N_38157,N_35786,N_35579);
xnor U38158 (N_38158,N_35676,N_36787);
or U38159 (N_38159,N_36024,N_36015);
xor U38160 (N_38160,N_37496,N_37046);
nand U38161 (N_38161,N_35324,N_36052);
nor U38162 (N_38162,N_36778,N_36964);
nand U38163 (N_38163,N_37310,N_35004);
nand U38164 (N_38164,N_35031,N_35659);
xor U38165 (N_38165,N_37463,N_37290);
or U38166 (N_38166,N_36181,N_35564);
xor U38167 (N_38167,N_35388,N_35061);
and U38168 (N_38168,N_37258,N_35544);
or U38169 (N_38169,N_35006,N_37162);
nor U38170 (N_38170,N_37112,N_36783);
nand U38171 (N_38171,N_36720,N_36050);
nor U38172 (N_38172,N_36301,N_36796);
and U38173 (N_38173,N_35707,N_35350);
and U38174 (N_38174,N_37119,N_36234);
xor U38175 (N_38175,N_35981,N_36044);
and U38176 (N_38176,N_36219,N_36436);
and U38177 (N_38177,N_35929,N_37434);
nand U38178 (N_38178,N_35718,N_35229);
and U38179 (N_38179,N_37311,N_35605);
nor U38180 (N_38180,N_36666,N_36930);
nor U38181 (N_38181,N_36950,N_35403);
xnor U38182 (N_38182,N_36322,N_37206);
nor U38183 (N_38183,N_37136,N_37141);
xor U38184 (N_38184,N_37229,N_36460);
nand U38185 (N_38185,N_35384,N_36171);
nand U38186 (N_38186,N_35846,N_36575);
and U38187 (N_38187,N_35796,N_36632);
nand U38188 (N_38188,N_36685,N_35018);
or U38189 (N_38189,N_36451,N_35253);
xor U38190 (N_38190,N_35550,N_35906);
nor U38191 (N_38191,N_35320,N_36732);
or U38192 (N_38192,N_35157,N_37373);
nor U38193 (N_38193,N_36423,N_37484);
nand U38194 (N_38194,N_35278,N_36866);
xor U38195 (N_38195,N_36865,N_35279);
or U38196 (N_38196,N_35912,N_35675);
or U38197 (N_38197,N_37086,N_36385);
nor U38198 (N_38198,N_35585,N_36872);
nand U38199 (N_38199,N_37411,N_37329);
nor U38200 (N_38200,N_36814,N_35679);
and U38201 (N_38201,N_35681,N_36114);
nor U38202 (N_38202,N_37336,N_37473);
and U38203 (N_38203,N_37208,N_36453);
or U38204 (N_38204,N_35874,N_35413);
or U38205 (N_38205,N_36779,N_35400);
nand U38206 (N_38206,N_37011,N_37094);
and U38207 (N_38207,N_35556,N_36232);
nand U38208 (N_38208,N_35366,N_37257);
xnor U38209 (N_38209,N_36363,N_35420);
nor U38210 (N_38210,N_36220,N_37235);
nand U38211 (N_38211,N_35546,N_36917);
or U38212 (N_38212,N_35444,N_37115);
and U38213 (N_38213,N_36528,N_35584);
xnor U38214 (N_38214,N_35127,N_36686);
and U38215 (N_38215,N_36399,N_36562);
or U38216 (N_38216,N_37406,N_37461);
nand U38217 (N_38217,N_36548,N_36817);
or U38218 (N_38218,N_36912,N_36332);
nand U38219 (N_38219,N_37277,N_35363);
xor U38220 (N_38220,N_37238,N_36618);
or U38221 (N_38221,N_36801,N_35670);
and U38222 (N_38222,N_37010,N_36039);
or U38223 (N_38223,N_37249,N_36947);
nand U38224 (N_38224,N_36358,N_37188);
and U38225 (N_38225,N_36780,N_36021);
and U38226 (N_38226,N_36245,N_37303);
nand U38227 (N_38227,N_36520,N_35686);
xnor U38228 (N_38228,N_37271,N_37071);
xor U38229 (N_38229,N_37194,N_35734);
xnor U38230 (N_38230,N_36444,N_35148);
or U38231 (N_38231,N_35766,N_35549);
xor U38232 (N_38232,N_37239,N_36310);
and U38233 (N_38233,N_36806,N_35385);
or U38234 (N_38234,N_36187,N_37479);
or U38235 (N_38235,N_37201,N_36570);
xnor U38236 (N_38236,N_35068,N_35262);
nor U38237 (N_38237,N_35308,N_37132);
nand U38238 (N_38238,N_37445,N_36591);
and U38239 (N_38239,N_37116,N_35793);
or U38240 (N_38240,N_36903,N_36821);
nand U38241 (N_38241,N_37062,N_36001);
nor U38242 (N_38242,N_36693,N_35529);
xnor U38243 (N_38243,N_35721,N_35079);
xnor U38244 (N_38244,N_37077,N_36415);
nor U38245 (N_38245,N_37309,N_37359);
xor U38246 (N_38246,N_36937,N_37006);
and U38247 (N_38247,N_37270,N_35083);
nand U38248 (N_38248,N_36349,N_35613);
nand U38249 (N_38249,N_36229,N_37390);
xnor U38250 (N_38250,N_35132,N_36989);
nor U38251 (N_38251,N_36758,N_36590);
nor U38252 (N_38252,N_35206,N_36323);
and U38253 (N_38253,N_37377,N_36307);
nor U38254 (N_38254,N_36825,N_36067);
nor U38255 (N_38255,N_37332,N_36681);
or U38256 (N_38256,N_35565,N_37304);
xor U38257 (N_38257,N_36191,N_36418);
nand U38258 (N_38258,N_36073,N_35566);
xnor U38259 (N_38259,N_36601,N_35292);
nor U38260 (N_38260,N_35852,N_37428);
xnor U38261 (N_38261,N_35073,N_37324);
nand U38262 (N_38262,N_37185,N_35232);
nand U38263 (N_38263,N_35110,N_36344);
nor U38264 (N_38264,N_36429,N_35438);
xor U38265 (N_38265,N_35484,N_36630);
or U38266 (N_38266,N_35653,N_36230);
or U38267 (N_38267,N_36991,N_37079);
and U38268 (N_38268,N_36448,N_37358);
xor U38269 (N_38269,N_35684,N_35152);
and U38270 (N_38270,N_36637,N_36141);
and U38271 (N_38271,N_36062,N_37426);
nor U38272 (N_38272,N_36752,N_37166);
nor U38273 (N_38273,N_35724,N_35297);
xnor U38274 (N_38274,N_36888,N_37371);
and U38275 (N_38275,N_35197,N_35726);
nor U38276 (N_38276,N_35362,N_35131);
and U38277 (N_38277,N_37101,N_35089);
nor U38278 (N_38278,N_36639,N_36029);
nand U38279 (N_38279,N_36606,N_35943);
and U38280 (N_38280,N_35607,N_35742);
xnor U38281 (N_38281,N_35656,N_35012);
xor U38282 (N_38282,N_35880,N_35746);
nand U38283 (N_38283,N_36820,N_35287);
and U38284 (N_38284,N_35819,N_37224);
or U38285 (N_38285,N_35198,N_36132);
and U38286 (N_38286,N_36193,N_35052);
nor U38287 (N_38287,N_35704,N_36376);
and U38288 (N_38288,N_36026,N_37471);
and U38289 (N_38289,N_35795,N_36100);
nor U38290 (N_38290,N_35462,N_35446);
nand U38291 (N_38291,N_35379,N_35394);
or U38292 (N_38292,N_36053,N_37064);
and U38293 (N_38293,N_36182,N_36459);
or U38294 (N_38294,N_37367,N_37362);
or U38295 (N_38295,N_37050,N_35500);
or U38296 (N_38296,N_35329,N_36470);
xor U38297 (N_38297,N_37096,N_35140);
xnor U38298 (N_38298,N_37395,N_37004);
or U38299 (N_38299,N_35398,N_36472);
xnor U38300 (N_38300,N_37127,N_35956);
nand U38301 (N_38301,N_37213,N_36902);
and U38302 (N_38302,N_36974,N_37403);
or U38303 (N_38303,N_35469,N_37320);
xor U38304 (N_38304,N_35674,N_36263);
and U38305 (N_38305,N_35733,N_35062);
xor U38306 (N_38306,N_37175,N_36188);
nor U38307 (N_38307,N_36545,N_37189);
xnor U38308 (N_38308,N_36791,N_35881);
nand U38309 (N_38309,N_37330,N_35351);
xor U38310 (N_38310,N_37416,N_35902);
and U38311 (N_38311,N_36558,N_35165);
nor U38312 (N_38312,N_37442,N_35395);
and U38313 (N_38313,N_36045,N_35861);
or U38314 (N_38314,N_36233,N_36477);
and U38315 (N_38315,N_35176,N_35960);
nand U38316 (N_38316,N_35540,N_35571);
or U38317 (N_38317,N_36106,N_35891);
nor U38318 (N_38318,N_36642,N_37016);
and U38319 (N_38319,N_36047,N_35100);
nand U38320 (N_38320,N_36273,N_35779);
nand U38321 (N_38321,N_36034,N_35247);
or U38322 (N_38322,N_37080,N_37498);
nor U38323 (N_38323,N_35775,N_35295);
and U38324 (N_38324,N_36270,N_37282);
or U38325 (N_38325,N_36289,N_36390);
nand U38326 (N_38326,N_37499,N_36723);
or U38327 (N_38327,N_36173,N_35424);
nor U38328 (N_38328,N_35449,N_37138);
and U38329 (N_38329,N_37002,N_35161);
nand U38330 (N_38330,N_35853,N_36356);
nand U38331 (N_38331,N_37177,N_36204);
nor U38332 (N_38332,N_35047,N_36433);
nand U38333 (N_38333,N_37038,N_35134);
nor U38334 (N_38334,N_35258,N_35781);
nor U38335 (N_38335,N_35624,N_35485);
xnor U38336 (N_38336,N_35442,N_36386);
nor U38337 (N_38337,N_35818,N_36871);
nor U38338 (N_38338,N_35979,N_35533);
xor U38339 (N_38339,N_35648,N_36507);
nor U38340 (N_38340,N_35767,N_36781);
nor U38341 (N_38341,N_36669,N_37001);
or U38342 (N_38342,N_35188,N_35558);
nor U38343 (N_38343,N_35422,N_35583);
or U38344 (N_38344,N_36346,N_36994);
and U38345 (N_38345,N_35207,N_36253);
xnor U38346 (N_38346,N_37237,N_35146);
and U38347 (N_38347,N_36588,N_36759);
nand U38348 (N_38348,N_36793,N_35496);
nor U38349 (N_38349,N_35036,N_36967);
nand U38350 (N_38350,N_35169,N_35141);
and U38351 (N_38351,N_36678,N_37431);
and U38352 (N_38352,N_36671,N_36750);
xnor U38353 (N_38353,N_37182,N_37300);
and U38354 (N_38354,N_35770,N_37021);
nor U38355 (N_38355,N_37465,N_37279);
and U38356 (N_38356,N_35589,N_35039);
or U38357 (N_38357,N_37036,N_35317);
nor U38358 (N_38358,N_36268,N_35708);
and U38359 (N_38359,N_36683,N_35213);
nor U38360 (N_38360,N_36555,N_37476);
xor U38361 (N_38361,N_35195,N_35923);
or U38362 (N_38362,N_36025,N_35353);
nor U38363 (N_38363,N_35035,N_35479);
nor U38364 (N_38364,N_35700,N_37123);
and U38365 (N_38365,N_35354,N_36465);
or U38366 (N_38366,N_36692,N_36286);
and U38367 (N_38367,N_35275,N_35175);
nand U38368 (N_38368,N_35037,N_36362);
xor U38369 (N_38369,N_35974,N_35758);
xnor U38370 (N_38370,N_35572,N_37493);
and U38371 (N_38371,N_36481,N_37351);
nand U38372 (N_38372,N_36719,N_37073);
and U38373 (N_38373,N_36969,N_36641);
nor U38374 (N_38374,N_35826,N_36427);
or U38375 (N_38375,N_35270,N_35466);
nor U38376 (N_38376,N_35017,N_35759);
and U38377 (N_38377,N_37053,N_35997);
or U38378 (N_38378,N_35581,N_36120);
or U38379 (N_38379,N_36457,N_36167);
xor U38380 (N_38380,N_36979,N_36677);
nand U38381 (N_38381,N_36643,N_35892);
nand U38382 (N_38382,N_37191,N_36051);
and U38383 (N_38383,N_37339,N_37245);
and U38384 (N_38384,N_36602,N_37252);
nand U38385 (N_38385,N_36105,N_36334);
xnor U38386 (N_38386,N_35523,N_36662);
and U38387 (N_38387,N_37015,N_36725);
nand U38388 (N_38388,N_35106,N_37155);
nor U38389 (N_38389,N_36563,N_36085);
xor U38390 (N_38390,N_36118,N_36854);
and U38391 (N_38391,N_37242,N_35603);
or U38392 (N_38392,N_35600,N_36636);
and U38393 (N_38393,N_35223,N_35381);
or U38394 (N_38394,N_35989,N_37149);
xor U38395 (N_38395,N_35933,N_35428);
xnor U38396 (N_38396,N_35472,N_36579);
and U38397 (N_38397,N_36822,N_37076);
and U38398 (N_38398,N_36578,N_36911);
or U38399 (N_38399,N_37200,N_35597);
and U38400 (N_38400,N_37105,N_36688);
nand U38401 (N_38401,N_35211,N_35967);
or U38402 (N_38402,N_36408,N_36198);
nand U38403 (N_38403,N_36288,N_36425);
and U38404 (N_38404,N_36944,N_35715);
or U38405 (N_38405,N_37490,N_35407);
xnor U38406 (N_38406,N_36694,N_36157);
and U38407 (N_38407,N_36395,N_35590);
nand U38408 (N_38408,N_35636,N_35573);
nor U38409 (N_38409,N_37195,N_36317);
and U38410 (N_38410,N_36554,N_36968);
or U38411 (N_38411,N_36097,N_35809);
xnor U38412 (N_38412,N_36458,N_35080);
xor U38413 (N_38413,N_36587,N_36447);
or U38414 (N_38414,N_36654,N_35269);
and U38415 (N_38415,N_35898,N_35499);
nand U38416 (N_38416,N_36030,N_35417);
xor U38417 (N_38417,N_37404,N_36115);
xnor U38418 (N_38418,N_35032,N_37241);
and U38419 (N_38419,N_35107,N_36197);
nand U38420 (N_38420,N_36351,N_35893);
and U38421 (N_38421,N_36407,N_35727);
nor U38422 (N_38422,N_35896,N_36567);
xor U38423 (N_38423,N_37345,N_35483);
xor U38424 (N_38424,N_37145,N_36294);
nor U38425 (N_38425,N_35256,N_35345);
and U38426 (N_38426,N_36221,N_35316);
nor U38427 (N_38427,N_35111,N_35985);
xnor U38428 (N_38428,N_36734,N_35730);
and U38429 (N_38429,N_36843,N_35697);
nor U38430 (N_38430,N_35947,N_37048);
xor U38431 (N_38431,N_35070,N_35537);
or U38432 (N_38432,N_35336,N_37419);
and U38433 (N_38433,N_36043,N_37202);
and U38434 (N_38434,N_35510,N_35662);
nor U38435 (N_38435,N_36063,N_36837);
nor U38436 (N_38436,N_37218,N_36098);
nor U38437 (N_38437,N_36933,N_37432);
xor U38438 (N_38438,N_37350,N_35946);
or U38439 (N_38439,N_35411,N_37226);
xnor U38440 (N_38440,N_36461,N_36561);
and U38441 (N_38441,N_36254,N_35248);
xnor U38442 (N_38442,N_36788,N_35606);
and U38443 (N_38443,N_35128,N_36973);
and U38444 (N_38444,N_36941,N_36166);
xor U38445 (N_38445,N_35208,N_36013);
xnor U38446 (N_38446,N_35828,N_36569);
nor U38447 (N_38447,N_36238,N_36183);
nand U38448 (N_38448,N_37444,N_36614);
and U38449 (N_38449,N_36054,N_36019);
nand U38450 (N_38450,N_36269,N_36971);
nand U38451 (N_38451,N_36200,N_35970);
nor U38452 (N_38452,N_36303,N_35034);
nand U38453 (N_38453,N_35913,N_37283);
nand U38454 (N_38454,N_37023,N_37207);
nand U38455 (N_38455,N_36069,N_36082);
nor U38456 (N_38456,N_35252,N_35092);
nand U38457 (N_38457,N_36260,N_36571);
nor U38458 (N_38458,N_35650,N_36089);
xor U38459 (N_38459,N_37380,N_36201);
nor U38460 (N_38460,N_35952,N_37203);
xnor U38461 (N_38461,N_36706,N_36679);
nand U38462 (N_38462,N_35657,N_35276);
nand U38463 (N_38463,N_37129,N_36131);
or U38464 (N_38464,N_36090,N_35705);
nor U38465 (N_38465,N_37421,N_37167);
nor U38466 (N_38466,N_35918,N_35941);
and U38467 (N_38467,N_35811,N_36302);
nand U38468 (N_38468,N_35359,N_35849);
and U38469 (N_38469,N_36093,N_35452);
xnor U38470 (N_38470,N_37481,N_36672);
and U38471 (N_38471,N_35267,N_35751);
xor U38472 (N_38472,N_35435,N_35850);
nand U38473 (N_38473,N_36022,N_35574);
and U38474 (N_38474,N_36999,N_35218);
xor U38475 (N_38475,N_35349,N_36017);
nand U38476 (N_38476,N_35725,N_36405);
xor U38477 (N_38477,N_36581,N_36623);
xnor U38478 (N_38478,N_37288,N_35632);
or U38479 (N_38479,N_36699,N_37074);
and U38480 (N_38480,N_35626,N_35762);
and U38481 (N_38481,N_36765,N_35521);
and U38482 (N_38482,N_37338,N_35069);
and U38483 (N_38483,N_36331,N_36372);
and U38484 (N_38484,N_35212,N_37475);
nand U38485 (N_38485,N_37420,N_37489);
xor U38486 (N_38486,N_36135,N_36290);
nor U38487 (N_38487,N_36549,N_37458);
nand U38488 (N_38488,N_35980,N_36250);
nor U38489 (N_38489,N_36402,N_36175);
or U38490 (N_38490,N_36380,N_36205);
and U38491 (N_38491,N_36369,N_36061);
nor U38492 (N_38492,N_36897,N_35822);
or U38493 (N_38493,N_36996,N_35167);
or U38494 (N_38494,N_35889,N_35436);
nand U38495 (N_38495,N_35922,N_35743);
or U38496 (N_38496,N_36151,N_36224);
xnor U38497 (N_38497,N_35119,N_36700);
or U38498 (N_38498,N_35334,N_36813);
nor U38499 (N_38499,N_36714,N_36839);
or U38500 (N_38500,N_36716,N_37280);
nor U38501 (N_38501,N_37393,N_35987);
nor U38502 (N_38502,N_36622,N_36337);
xnor U38503 (N_38503,N_36282,N_36241);
and U38504 (N_38504,N_36515,N_35800);
and U38505 (N_38505,N_35327,N_35611);
nor U38506 (N_38506,N_36400,N_35614);
or U38507 (N_38507,N_37429,N_36373);
or U38508 (N_38508,N_35845,N_36212);
and U38509 (N_38509,N_37448,N_35130);
and U38510 (N_38510,N_37415,N_36676);
or U38511 (N_38511,N_36760,N_36264);
and U38512 (N_38512,N_36616,N_36674);
nand U38513 (N_38513,N_37266,N_36878);
or U38514 (N_38514,N_36848,N_35548);
nand U38515 (N_38515,N_36277,N_36240);
xor U38516 (N_38516,N_35294,N_37474);
xnor U38517 (N_38517,N_36489,N_36170);
or U38518 (N_38518,N_36785,N_35014);
nand U38519 (N_38519,N_37204,N_37142);
or U38520 (N_38520,N_36565,N_35259);
and U38521 (N_38521,N_35155,N_36731);
and U38522 (N_38522,N_36711,N_37264);
and U38523 (N_38523,N_35915,N_37472);
nor U38524 (N_38524,N_35170,N_36635);
xnor U38525 (N_38525,N_36556,N_35431);
or U38526 (N_38526,N_37103,N_36466);
or U38527 (N_38527,N_35739,N_36443);
nor U38528 (N_38528,N_36136,N_35461);
or U38529 (N_38529,N_37163,N_35557);
or U38530 (N_38530,N_37327,N_37316);
and U38531 (N_38531,N_36086,N_37298);
xnor U38532 (N_38532,N_36394,N_36409);
nor U38533 (N_38533,N_35842,N_35560);
or U38534 (N_38534,N_35486,N_36367);
nand U38535 (N_38535,N_36915,N_37150);
xor U38536 (N_38536,N_36312,N_35525);
nand U38537 (N_38537,N_35680,N_36185);
xnor U38538 (N_38538,N_35968,N_36651);
nand U38539 (N_38539,N_35124,N_36802);
xnor U38540 (N_38540,N_35616,N_35863);
nor U38541 (N_38541,N_36763,N_35009);
and U38542 (N_38542,N_35201,N_35723);
and U38543 (N_38543,N_35817,N_36474);
nand U38544 (N_38544,N_35225,N_37278);
and U38545 (N_38545,N_35748,N_37251);
xnor U38546 (N_38546,N_37085,N_36855);
or U38547 (N_38547,N_35982,N_35777);
or U38548 (N_38548,N_37043,N_36169);
and U38549 (N_38549,N_36961,N_35059);
xnor U38550 (N_38550,N_36727,N_36739);
nand U38551 (N_38551,N_36774,N_36687);
nor U38552 (N_38552,N_35984,N_36194);
or U38553 (N_38553,N_36742,N_36935);
nor U38554 (N_38554,N_36951,N_37051);
nand U38555 (N_38555,N_35421,N_35864);
xnor U38556 (N_38556,N_36673,N_36874);
xor U38557 (N_38557,N_36324,N_36621);
nand U38558 (N_38558,N_36612,N_36702);
xnor U38559 (N_38559,N_36113,N_35114);
or U38560 (N_38560,N_35392,N_36882);
nor U38561 (N_38561,N_36153,N_35088);
xor U38562 (N_38562,N_37042,N_37007);
nand U38563 (N_38563,N_36741,N_35181);
or U38564 (N_38564,N_36675,N_36041);
nand U38565 (N_38565,N_35999,N_37343);
or U38566 (N_38566,N_35801,N_35166);
or U38567 (N_38567,N_36434,N_36997);
and U38568 (N_38568,N_36006,N_36697);
nor U38569 (N_38569,N_36278,N_36860);
nor U38570 (N_38570,N_35710,N_37014);
nor U38571 (N_38571,N_36875,N_35467);
nor U38572 (N_38572,N_36123,N_35402);
and U38573 (N_38573,N_35415,N_35551);
xnor U38574 (N_38574,N_35834,N_36355);
nor U38575 (N_38575,N_35147,N_35935);
xor U38576 (N_38576,N_36652,N_36736);
nor U38577 (N_38577,N_36767,N_37272);
or U38578 (N_38578,N_36379,N_37161);
or U38579 (N_38579,N_35622,N_35872);
xnor U38580 (N_38580,N_35854,N_36770);
nor U38581 (N_38581,N_37184,N_37407);
or U38582 (N_38582,N_36177,N_35476);
nand U38583 (N_38583,N_37269,N_35806);
xor U38584 (N_38584,N_35226,N_36352);
and U38585 (N_38585,N_37158,N_36003);
nand U38586 (N_38586,N_35592,N_35387);
nor U38587 (N_38587,N_36696,N_36435);
nor U38588 (N_38588,N_35692,N_36430);
or U38589 (N_38589,N_35219,N_36879);
nor U38590 (N_38590,N_37427,N_35372);
or U38591 (N_38591,N_36134,N_36982);
nand U38592 (N_38592,N_35448,N_37313);
nor U38593 (N_38593,N_35719,N_36252);
nand U38594 (N_38594,N_35905,N_36926);
xor U38595 (N_38595,N_36309,N_36213);
nand U38596 (N_38596,N_35343,N_36007);
or U38597 (N_38597,N_35163,N_36609);
or U38598 (N_38598,N_37069,N_37384);
nand U38599 (N_38599,N_36226,N_37025);
and U38600 (N_38600,N_36847,N_36764);
nor U38601 (N_38601,N_37210,N_37217);
nand U38602 (N_38602,N_36382,N_35750);
and U38603 (N_38603,N_35689,N_35909);
and U38604 (N_38604,N_35209,N_37019);
or U38605 (N_38605,N_37267,N_35621);
nand U38606 (N_38606,N_36295,N_35780);
xor U38607 (N_38607,N_35505,N_35582);
nand U38608 (N_38608,N_35333,N_35631);
xnor U38609 (N_38609,N_37044,N_37230);
and U38610 (N_38610,N_35608,N_35118);
and U38611 (N_38611,N_37260,N_35112);
or U38612 (N_38612,N_36392,N_35682);
and U38613 (N_38613,N_35663,N_37352);
nor U38614 (N_38614,N_37454,N_37215);
nor U38615 (N_38615,N_36511,N_36818);
xnor U38616 (N_38616,N_35950,N_36737);
and U38617 (N_38617,N_35695,N_36966);
nor U38618 (N_38618,N_37193,N_36542);
nor U38619 (N_38619,N_37181,N_37093);
and U38620 (N_38620,N_37405,N_36338);
nor U38621 (N_38621,N_36799,N_35966);
xor U38622 (N_38622,N_37396,N_36174);
nand U38623 (N_38623,N_36217,N_37219);
or U38624 (N_38624,N_36227,N_35973);
nor U38625 (N_38625,N_35498,N_35245);
nand U38626 (N_38626,N_35939,N_37328);
nor U38627 (N_38627,N_36819,N_35412);
xnor U38628 (N_38628,N_35799,N_36112);
xor U38629 (N_38629,N_35532,N_35077);
xnor U38630 (N_38630,N_35265,N_35661);
nand U38631 (N_38631,N_36247,N_35313);
nand U38632 (N_38632,N_35383,N_36143);
and U38633 (N_38633,N_35271,N_37319);
xor U38634 (N_38634,N_35086,N_37083);
or U38635 (N_38635,N_36339,N_36998);
or U38636 (N_38636,N_37321,N_36907);
and U38637 (N_38637,N_37140,N_36366);
and U38638 (N_38638,N_36165,N_35975);
or U38639 (N_38639,N_35744,N_36196);
and U38640 (N_38640,N_36125,N_37305);
nand U38641 (N_38641,N_36340,N_36065);
nand U38642 (N_38642,N_35835,N_36559);
nand U38643 (N_38643,N_35090,N_36952);
and U38644 (N_38644,N_36516,N_36281);
or U38645 (N_38645,N_35784,N_35911);
and U38646 (N_38646,N_36745,N_37414);
and U38647 (N_38647,N_36743,N_36464);
nor U38648 (N_38648,N_36014,N_37209);
and U38649 (N_38649,N_37098,N_37449);
nand U38650 (N_38650,N_35690,N_36598);
nor U38651 (N_38651,N_35515,N_36626);
nor U38652 (N_38652,N_35908,N_36468);
and U38653 (N_38653,N_35808,N_36291);
xnor U38654 (N_38654,N_35890,N_35703);
and U38655 (N_38655,N_35920,N_35460);
xor U38656 (N_38656,N_36747,N_37211);
or U38657 (N_38657,N_35145,N_35439);
or U38658 (N_38658,N_37289,N_35685);
and U38659 (N_38659,N_36236,N_35993);
nor U38660 (N_38660,N_36360,N_35542);
and U38661 (N_38661,N_35374,N_36949);
nand U38662 (N_38662,N_35000,N_36990);
nand U38663 (N_38663,N_37164,N_37363);
or U38664 (N_38664,N_35242,N_36921);
nand U38665 (N_38665,N_36827,N_36757);
nor U38666 (N_38666,N_35109,N_36580);
nand U38667 (N_38667,N_37346,N_36035);
xor U38668 (N_38668,N_37054,N_35136);
nand U38669 (N_38669,N_35352,N_36744);
and U38670 (N_38670,N_37361,N_36492);
nor U38671 (N_38671,N_35895,N_36733);
xor U38672 (N_38672,N_35331,N_36715);
and U38673 (N_38673,N_36573,N_35196);
and U38674 (N_38674,N_35701,N_37349);
xor U38675 (N_38675,N_36842,N_35360);
xor U38676 (N_38676,N_35729,N_37424);
nand U38677 (N_38677,N_35406,N_35053);
or U38678 (N_38678,N_37060,N_35173);
or U38679 (N_38679,N_35951,N_35433);
nand U38680 (N_38680,N_35144,N_37216);
nor U38681 (N_38681,N_35129,N_35598);
nor U38682 (N_38682,N_35418,N_35233);
nor U38683 (N_38683,N_35798,N_36243);
nand U38684 (N_38684,N_35121,N_36564);
or U38685 (N_38685,N_35524,N_35821);
or U38686 (N_38686,N_35804,N_35901);
and U38687 (N_38687,N_35651,N_36327);
nor U38688 (N_38688,N_36439,N_36703);
nand U38689 (N_38689,N_36223,N_36235);
nand U38690 (N_38690,N_36348,N_37118);
and U38691 (N_38691,N_37009,N_36494);
and U38692 (N_38692,N_35095,N_35003);
nand U38693 (N_38693,N_37291,N_37035);
and U38694 (N_38694,N_36853,N_35296);
nand U38695 (N_38695,N_35763,N_35957);
nand U38696 (N_38696,N_36116,N_35635);
xor U38697 (N_38697,N_37268,N_36437);
xor U38698 (N_38698,N_35268,N_36272);
nand U38699 (N_38699,N_37470,N_36600);
xnor U38700 (N_38700,N_37376,N_35738);
nor U38701 (N_38701,N_36705,N_37067);
xor U38702 (N_38702,N_36960,N_36297);
or U38703 (N_38703,N_35304,N_37492);
or U38704 (N_38704,N_35437,N_36909);
xnor U38705 (N_38705,N_36450,N_35277);
or U38706 (N_38706,N_37247,N_36368);
and U38707 (N_38707,N_36161,N_37265);
nor U38708 (N_38708,N_36660,N_37408);
or U38709 (N_38709,N_36784,N_37032);
xnor U38710 (N_38710,N_36751,N_36280);
or U38711 (N_38711,N_35847,N_35282);
xor U38712 (N_38712,N_35192,N_36749);
and U38713 (N_38713,N_35884,N_36828);
or U38714 (N_38714,N_36178,N_35969);
nand U38715 (N_38715,N_35552,N_37322);
nor U38716 (N_38716,N_35007,N_35921);
nand U38717 (N_38717,N_37296,N_36375);
xnor U38718 (N_38718,N_37173,N_36087);
xnor U38719 (N_38719,N_36154,N_37122);
and U38720 (N_38720,N_37196,N_35914);
nand U38721 (N_38721,N_36890,N_36539);
nand U38722 (N_38722,N_36876,N_36387);
or U38723 (N_38723,N_36925,N_35396);
xnor U38724 (N_38724,N_36891,N_35094);
nand U38725 (N_38725,N_35286,N_37397);
or U38726 (N_38726,N_36419,N_37306);
nand U38727 (N_38727,N_35888,N_36341);
nor U38728 (N_38728,N_35807,N_35078);
nor U38729 (N_38729,N_37108,N_35344);
nand U38730 (N_38730,N_36927,N_36713);
nor U38731 (N_38731,N_35696,N_35199);
nand U38732 (N_38732,N_36350,N_36541);
and U38733 (N_38733,N_37335,N_35200);
nand U38734 (N_38734,N_35688,N_35646);
nor U38735 (N_38735,N_37057,N_35904);
and U38736 (N_38736,N_36208,N_36560);
nand U38737 (N_38737,N_35813,N_35171);
and U38738 (N_38738,N_37084,N_36877);
and U38739 (N_38739,N_36525,N_35749);
and U38740 (N_38740,N_36206,N_36449);
nand U38741 (N_38741,N_35773,N_35378);
and U38742 (N_38742,N_35567,N_37082);
or U38743 (N_38743,N_37262,N_35364);
and U38744 (N_38744,N_35318,N_35330);
nor U38745 (N_38745,N_36931,N_36735);
or U38746 (N_38746,N_36149,N_36033);
nor U38747 (N_38747,N_36381,N_36325);
nand U38748 (N_38748,N_36122,N_35340);
or U38749 (N_38749,N_35752,N_37178);
and U38750 (N_38750,N_35608,N_37205);
or U38751 (N_38751,N_35643,N_35788);
or U38752 (N_38752,N_35198,N_35071);
xor U38753 (N_38753,N_35865,N_35367);
or U38754 (N_38754,N_36133,N_35706);
xor U38755 (N_38755,N_36376,N_35470);
and U38756 (N_38756,N_37313,N_37173);
and U38757 (N_38757,N_35287,N_36358);
nand U38758 (N_38758,N_35372,N_35862);
or U38759 (N_38759,N_35972,N_35786);
or U38760 (N_38760,N_35844,N_35736);
or U38761 (N_38761,N_35747,N_35585);
nand U38762 (N_38762,N_37461,N_37140);
nand U38763 (N_38763,N_36039,N_35060);
xnor U38764 (N_38764,N_35943,N_37399);
xnor U38765 (N_38765,N_37185,N_36931);
nor U38766 (N_38766,N_35452,N_37156);
or U38767 (N_38767,N_35449,N_37316);
xnor U38768 (N_38768,N_35725,N_36997);
nor U38769 (N_38769,N_36616,N_35894);
or U38770 (N_38770,N_36298,N_35212);
or U38771 (N_38771,N_35233,N_36922);
nand U38772 (N_38772,N_35777,N_37133);
and U38773 (N_38773,N_35128,N_36963);
or U38774 (N_38774,N_37231,N_37237);
xnor U38775 (N_38775,N_35874,N_36030);
and U38776 (N_38776,N_35613,N_36704);
and U38777 (N_38777,N_36770,N_35195);
xor U38778 (N_38778,N_36426,N_35318);
nor U38779 (N_38779,N_35588,N_37403);
nor U38780 (N_38780,N_36268,N_35865);
and U38781 (N_38781,N_35819,N_36108);
nand U38782 (N_38782,N_36287,N_36985);
or U38783 (N_38783,N_37427,N_37284);
nand U38784 (N_38784,N_36589,N_36431);
nand U38785 (N_38785,N_35668,N_35815);
and U38786 (N_38786,N_35066,N_36222);
xor U38787 (N_38787,N_36574,N_35627);
and U38788 (N_38788,N_36860,N_36000);
nor U38789 (N_38789,N_35581,N_37415);
and U38790 (N_38790,N_36430,N_35229);
xor U38791 (N_38791,N_35219,N_36529);
nand U38792 (N_38792,N_36207,N_35264);
xnor U38793 (N_38793,N_36223,N_37278);
nand U38794 (N_38794,N_37360,N_36055);
nand U38795 (N_38795,N_36301,N_37232);
xnor U38796 (N_38796,N_36295,N_35005);
and U38797 (N_38797,N_37067,N_36262);
nor U38798 (N_38798,N_36364,N_35016);
xnor U38799 (N_38799,N_35239,N_35071);
nor U38800 (N_38800,N_37240,N_35759);
xor U38801 (N_38801,N_37453,N_35494);
or U38802 (N_38802,N_36707,N_36862);
or U38803 (N_38803,N_35811,N_35159);
nand U38804 (N_38804,N_37420,N_35028);
and U38805 (N_38805,N_36081,N_35656);
or U38806 (N_38806,N_37364,N_37260);
nor U38807 (N_38807,N_37361,N_35958);
xnor U38808 (N_38808,N_37124,N_35477);
nand U38809 (N_38809,N_35178,N_36205);
or U38810 (N_38810,N_35194,N_37141);
nand U38811 (N_38811,N_37036,N_35446);
or U38812 (N_38812,N_35214,N_36265);
or U38813 (N_38813,N_36030,N_35770);
or U38814 (N_38814,N_35018,N_37102);
or U38815 (N_38815,N_37356,N_36698);
xnor U38816 (N_38816,N_36532,N_37111);
and U38817 (N_38817,N_37181,N_35092);
xnor U38818 (N_38818,N_35777,N_36675);
and U38819 (N_38819,N_35040,N_35089);
nor U38820 (N_38820,N_35511,N_37262);
nand U38821 (N_38821,N_36464,N_37407);
nand U38822 (N_38822,N_35107,N_35089);
and U38823 (N_38823,N_36294,N_36659);
xor U38824 (N_38824,N_36063,N_35227);
xor U38825 (N_38825,N_37216,N_35286);
nand U38826 (N_38826,N_36034,N_36686);
nor U38827 (N_38827,N_36842,N_37397);
nand U38828 (N_38828,N_36849,N_36304);
and U38829 (N_38829,N_35719,N_36009);
nor U38830 (N_38830,N_35262,N_37398);
and U38831 (N_38831,N_36250,N_36540);
and U38832 (N_38832,N_35138,N_36121);
or U38833 (N_38833,N_35073,N_35133);
and U38834 (N_38834,N_36249,N_35798);
xnor U38835 (N_38835,N_35743,N_35456);
xnor U38836 (N_38836,N_36999,N_35086);
xor U38837 (N_38837,N_35747,N_35860);
and U38838 (N_38838,N_35122,N_36815);
xnor U38839 (N_38839,N_35086,N_37054);
nand U38840 (N_38840,N_37156,N_35287);
xor U38841 (N_38841,N_35883,N_35546);
xor U38842 (N_38842,N_36514,N_36554);
nand U38843 (N_38843,N_36056,N_37041);
nand U38844 (N_38844,N_35126,N_35242);
xnor U38845 (N_38845,N_36549,N_36673);
or U38846 (N_38846,N_36498,N_36222);
and U38847 (N_38847,N_36614,N_35801);
nor U38848 (N_38848,N_37188,N_35034);
nor U38849 (N_38849,N_35246,N_35614);
xnor U38850 (N_38850,N_35331,N_35163);
or U38851 (N_38851,N_36627,N_36172);
and U38852 (N_38852,N_35325,N_35141);
nor U38853 (N_38853,N_36901,N_36812);
or U38854 (N_38854,N_35367,N_37066);
nand U38855 (N_38855,N_36472,N_36429);
or U38856 (N_38856,N_36303,N_36826);
xor U38857 (N_38857,N_35011,N_35802);
and U38858 (N_38858,N_35464,N_36790);
xnor U38859 (N_38859,N_36464,N_36673);
nand U38860 (N_38860,N_36604,N_37363);
or U38861 (N_38861,N_36261,N_36204);
nor U38862 (N_38862,N_36714,N_35667);
or U38863 (N_38863,N_35189,N_35385);
nand U38864 (N_38864,N_36287,N_36492);
nand U38865 (N_38865,N_36203,N_35818);
or U38866 (N_38866,N_36034,N_36596);
and U38867 (N_38867,N_35471,N_37479);
nor U38868 (N_38868,N_36745,N_36813);
xnor U38869 (N_38869,N_35939,N_36962);
or U38870 (N_38870,N_37229,N_36795);
nand U38871 (N_38871,N_36829,N_37426);
and U38872 (N_38872,N_37202,N_35305);
and U38873 (N_38873,N_35160,N_35296);
xor U38874 (N_38874,N_35959,N_36722);
xnor U38875 (N_38875,N_35854,N_35432);
or U38876 (N_38876,N_36828,N_36703);
nand U38877 (N_38877,N_35014,N_35290);
nor U38878 (N_38878,N_35269,N_36331);
nor U38879 (N_38879,N_35131,N_37338);
or U38880 (N_38880,N_35583,N_36775);
xor U38881 (N_38881,N_37082,N_37151);
xnor U38882 (N_38882,N_35099,N_36793);
nor U38883 (N_38883,N_35222,N_37043);
or U38884 (N_38884,N_36006,N_37390);
and U38885 (N_38885,N_35380,N_36235);
or U38886 (N_38886,N_35116,N_36428);
or U38887 (N_38887,N_35727,N_37476);
or U38888 (N_38888,N_36442,N_36222);
and U38889 (N_38889,N_36771,N_35431);
nand U38890 (N_38890,N_35794,N_37214);
nand U38891 (N_38891,N_35557,N_36393);
nand U38892 (N_38892,N_35591,N_36949);
and U38893 (N_38893,N_36310,N_36228);
xnor U38894 (N_38894,N_36854,N_36551);
nand U38895 (N_38895,N_35751,N_36250);
nand U38896 (N_38896,N_36530,N_37158);
nor U38897 (N_38897,N_36410,N_36803);
nor U38898 (N_38898,N_36732,N_36894);
nor U38899 (N_38899,N_37494,N_37169);
nand U38900 (N_38900,N_36952,N_36367);
and U38901 (N_38901,N_35238,N_35248);
nand U38902 (N_38902,N_35450,N_35643);
nor U38903 (N_38903,N_37095,N_35912);
nand U38904 (N_38904,N_36299,N_35789);
nor U38905 (N_38905,N_37022,N_36819);
nor U38906 (N_38906,N_37263,N_36647);
nor U38907 (N_38907,N_37082,N_37023);
and U38908 (N_38908,N_36982,N_35445);
nor U38909 (N_38909,N_36843,N_36633);
and U38910 (N_38910,N_36893,N_35812);
and U38911 (N_38911,N_35969,N_35864);
or U38912 (N_38912,N_37176,N_35234);
or U38913 (N_38913,N_37159,N_36739);
nand U38914 (N_38914,N_36049,N_35514);
xor U38915 (N_38915,N_36715,N_36716);
nand U38916 (N_38916,N_36342,N_35062);
or U38917 (N_38917,N_37384,N_36650);
and U38918 (N_38918,N_36957,N_36799);
or U38919 (N_38919,N_37497,N_35772);
and U38920 (N_38920,N_36385,N_37499);
xnor U38921 (N_38921,N_35735,N_36261);
or U38922 (N_38922,N_36275,N_35457);
nand U38923 (N_38923,N_36219,N_36741);
xor U38924 (N_38924,N_36681,N_36595);
or U38925 (N_38925,N_37352,N_35706);
or U38926 (N_38926,N_35216,N_37085);
nand U38927 (N_38927,N_36488,N_35441);
or U38928 (N_38928,N_37312,N_36387);
xor U38929 (N_38929,N_37233,N_35619);
nor U38930 (N_38930,N_37190,N_36698);
xnor U38931 (N_38931,N_35110,N_36577);
xor U38932 (N_38932,N_35519,N_36442);
nor U38933 (N_38933,N_36443,N_36298);
nand U38934 (N_38934,N_36956,N_36391);
nand U38935 (N_38935,N_35842,N_35788);
and U38936 (N_38936,N_36857,N_37492);
nand U38937 (N_38937,N_37327,N_37177);
xor U38938 (N_38938,N_36784,N_36587);
or U38939 (N_38939,N_35635,N_35471);
or U38940 (N_38940,N_37180,N_36068);
or U38941 (N_38941,N_35304,N_35135);
nor U38942 (N_38942,N_36494,N_37086);
nand U38943 (N_38943,N_36446,N_36238);
and U38944 (N_38944,N_37314,N_35289);
nor U38945 (N_38945,N_35879,N_37049);
nand U38946 (N_38946,N_35513,N_36307);
xnor U38947 (N_38947,N_35480,N_36359);
nand U38948 (N_38948,N_36263,N_36406);
nor U38949 (N_38949,N_36553,N_36394);
or U38950 (N_38950,N_36312,N_35075);
or U38951 (N_38951,N_37129,N_36806);
nand U38952 (N_38952,N_36568,N_35167);
nor U38953 (N_38953,N_35122,N_35528);
or U38954 (N_38954,N_36241,N_37288);
nand U38955 (N_38955,N_36998,N_37041);
xor U38956 (N_38956,N_36167,N_36271);
and U38957 (N_38957,N_35440,N_36378);
nor U38958 (N_38958,N_36403,N_37480);
nor U38959 (N_38959,N_37031,N_35574);
or U38960 (N_38960,N_35387,N_35532);
nand U38961 (N_38961,N_35881,N_35065);
nand U38962 (N_38962,N_37458,N_36006);
and U38963 (N_38963,N_36465,N_37060);
xor U38964 (N_38964,N_37495,N_37470);
or U38965 (N_38965,N_35473,N_35521);
and U38966 (N_38966,N_36082,N_35260);
nor U38967 (N_38967,N_37197,N_35983);
nand U38968 (N_38968,N_35648,N_36404);
and U38969 (N_38969,N_36079,N_36132);
or U38970 (N_38970,N_35447,N_37021);
nand U38971 (N_38971,N_35779,N_35406);
nand U38972 (N_38972,N_36377,N_37003);
nand U38973 (N_38973,N_37079,N_36047);
nor U38974 (N_38974,N_37304,N_35705);
or U38975 (N_38975,N_37391,N_36972);
and U38976 (N_38976,N_35147,N_37047);
xnor U38977 (N_38977,N_37216,N_37128);
nand U38978 (N_38978,N_35635,N_35146);
or U38979 (N_38979,N_36777,N_35561);
xnor U38980 (N_38980,N_35239,N_37340);
or U38981 (N_38981,N_36176,N_35150);
xor U38982 (N_38982,N_36115,N_35455);
xor U38983 (N_38983,N_36474,N_36250);
xnor U38984 (N_38984,N_35324,N_35592);
or U38985 (N_38985,N_35366,N_36966);
nor U38986 (N_38986,N_36583,N_37019);
or U38987 (N_38987,N_36410,N_35201);
xor U38988 (N_38988,N_37296,N_35200);
nand U38989 (N_38989,N_36592,N_37221);
xor U38990 (N_38990,N_36865,N_36626);
nand U38991 (N_38991,N_36753,N_36873);
nor U38992 (N_38992,N_36533,N_37118);
nor U38993 (N_38993,N_36188,N_35358);
nor U38994 (N_38994,N_36161,N_36073);
nand U38995 (N_38995,N_35073,N_36200);
and U38996 (N_38996,N_36496,N_35672);
or U38997 (N_38997,N_36043,N_35355);
nand U38998 (N_38998,N_35979,N_35609);
and U38999 (N_38999,N_36356,N_36960);
and U39000 (N_39000,N_35030,N_35846);
xor U39001 (N_39001,N_36944,N_35178);
nand U39002 (N_39002,N_36359,N_36380);
nand U39003 (N_39003,N_35372,N_36210);
or U39004 (N_39004,N_35526,N_35315);
nand U39005 (N_39005,N_35230,N_35069);
or U39006 (N_39006,N_36648,N_36306);
nand U39007 (N_39007,N_36745,N_37267);
xor U39008 (N_39008,N_36997,N_36714);
and U39009 (N_39009,N_37283,N_35883);
or U39010 (N_39010,N_36682,N_36227);
or U39011 (N_39011,N_36762,N_36389);
xor U39012 (N_39012,N_36557,N_37390);
nor U39013 (N_39013,N_35174,N_36123);
and U39014 (N_39014,N_36775,N_36606);
nor U39015 (N_39015,N_35557,N_37346);
nor U39016 (N_39016,N_36814,N_35965);
xnor U39017 (N_39017,N_35345,N_36422);
nand U39018 (N_39018,N_36852,N_35830);
xnor U39019 (N_39019,N_37129,N_35305);
nor U39020 (N_39020,N_36903,N_35131);
or U39021 (N_39021,N_37181,N_37420);
nand U39022 (N_39022,N_36698,N_36076);
or U39023 (N_39023,N_36451,N_36627);
and U39024 (N_39024,N_36713,N_35736);
nor U39025 (N_39025,N_35773,N_37138);
nor U39026 (N_39026,N_37285,N_37167);
xnor U39027 (N_39027,N_35375,N_36228);
and U39028 (N_39028,N_35982,N_37265);
nand U39029 (N_39029,N_35451,N_37491);
and U39030 (N_39030,N_37449,N_35266);
nor U39031 (N_39031,N_35140,N_35586);
nor U39032 (N_39032,N_35667,N_37104);
and U39033 (N_39033,N_37049,N_36274);
nor U39034 (N_39034,N_35978,N_37080);
or U39035 (N_39035,N_35972,N_36097);
nand U39036 (N_39036,N_35616,N_36474);
or U39037 (N_39037,N_35386,N_35351);
and U39038 (N_39038,N_37024,N_35937);
and U39039 (N_39039,N_35582,N_35296);
nor U39040 (N_39040,N_36542,N_37051);
xnor U39041 (N_39041,N_35884,N_36259);
xnor U39042 (N_39042,N_36045,N_35067);
or U39043 (N_39043,N_36371,N_36695);
nor U39044 (N_39044,N_36603,N_35659);
and U39045 (N_39045,N_35370,N_36757);
and U39046 (N_39046,N_36108,N_35766);
nand U39047 (N_39047,N_35894,N_35163);
or U39048 (N_39048,N_37008,N_36459);
and U39049 (N_39049,N_35153,N_36630);
xor U39050 (N_39050,N_36990,N_37016);
nand U39051 (N_39051,N_36491,N_35248);
xor U39052 (N_39052,N_35864,N_35740);
nand U39053 (N_39053,N_36823,N_36690);
nand U39054 (N_39054,N_35583,N_36389);
or U39055 (N_39055,N_36265,N_36456);
nor U39056 (N_39056,N_36868,N_36398);
nand U39057 (N_39057,N_35150,N_36397);
and U39058 (N_39058,N_36020,N_35483);
nor U39059 (N_39059,N_35982,N_37466);
or U39060 (N_39060,N_36743,N_36171);
nor U39061 (N_39061,N_35774,N_35646);
xnor U39062 (N_39062,N_36560,N_35091);
nor U39063 (N_39063,N_35897,N_35071);
nand U39064 (N_39064,N_35529,N_35111);
xor U39065 (N_39065,N_35843,N_36890);
nand U39066 (N_39066,N_35592,N_35015);
nor U39067 (N_39067,N_35539,N_37151);
or U39068 (N_39068,N_35786,N_36510);
xor U39069 (N_39069,N_36339,N_35930);
xnor U39070 (N_39070,N_36137,N_36857);
nor U39071 (N_39071,N_35610,N_36966);
or U39072 (N_39072,N_35036,N_37309);
nor U39073 (N_39073,N_35100,N_35692);
nor U39074 (N_39074,N_36997,N_36844);
xnor U39075 (N_39075,N_36057,N_37410);
or U39076 (N_39076,N_36293,N_35643);
nand U39077 (N_39077,N_36500,N_37087);
or U39078 (N_39078,N_35920,N_35675);
or U39079 (N_39079,N_35946,N_36141);
xor U39080 (N_39080,N_36043,N_36246);
xnor U39081 (N_39081,N_37315,N_37380);
nor U39082 (N_39082,N_35079,N_36604);
nor U39083 (N_39083,N_36006,N_35271);
xor U39084 (N_39084,N_37394,N_35007);
xnor U39085 (N_39085,N_35897,N_35628);
and U39086 (N_39086,N_35420,N_37075);
and U39087 (N_39087,N_35074,N_36825);
nand U39088 (N_39088,N_35135,N_35254);
and U39089 (N_39089,N_36564,N_37062);
nand U39090 (N_39090,N_35019,N_36642);
xor U39091 (N_39091,N_36717,N_37164);
and U39092 (N_39092,N_35261,N_36640);
nor U39093 (N_39093,N_35381,N_36254);
xor U39094 (N_39094,N_37160,N_36956);
nor U39095 (N_39095,N_35107,N_35176);
xnor U39096 (N_39096,N_36234,N_37472);
and U39097 (N_39097,N_36642,N_35088);
nand U39098 (N_39098,N_35935,N_36929);
or U39099 (N_39099,N_35782,N_37106);
or U39100 (N_39100,N_35431,N_36479);
or U39101 (N_39101,N_35666,N_37257);
or U39102 (N_39102,N_35572,N_35358);
xnor U39103 (N_39103,N_36052,N_37231);
nor U39104 (N_39104,N_35724,N_35126);
nand U39105 (N_39105,N_37085,N_35002);
xor U39106 (N_39106,N_36126,N_35556);
xnor U39107 (N_39107,N_35353,N_35845);
nand U39108 (N_39108,N_37310,N_36649);
and U39109 (N_39109,N_35331,N_36825);
and U39110 (N_39110,N_35350,N_36129);
nor U39111 (N_39111,N_36638,N_36506);
nor U39112 (N_39112,N_35286,N_35019);
nor U39113 (N_39113,N_36682,N_35011);
or U39114 (N_39114,N_35859,N_37078);
and U39115 (N_39115,N_36376,N_35307);
or U39116 (N_39116,N_37073,N_36950);
nor U39117 (N_39117,N_37146,N_37302);
and U39118 (N_39118,N_35148,N_36505);
xnor U39119 (N_39119,N_36938,N_35413);
nor U39120 (N_39120,N_37212,N_36551);
or U39121 (N_39121,N_35358,N_35177);
xor U39122 (N_39122,N_35922,N_36089);
nor U39123 (N_39123,N_36544,N_35039);
nor U39124 (N_39124,N_35219,N_35910);
xor U39125 (N_39125,N_35901,N_37326);
and U39126 (N_39126,N_36680,N_35337);
nor U39127 (N_39127,N_36325,N_36490);
and U39128 (N_39128,N_35179,N_36209);
or U39129 (N_39129,N_37242,N_36082);
nor U39130 (N_39130,N_35627,N_36793);
and U39131 (N_39131,N_36817,N_35216);
nand U39132 (N_39132,N_35148,N_35845);
xnor U39133 (N_39133,N_35230,N_37109);
nand U39134 (N_39134,N_35581,N_36327);
nand U39135 (N_39135,N_37358,N_35889);
nor U39136 (N_39136,N_35141,N_37440);
or U39137 (N_39137,N_35210,N_35786);
or U39138 (N_39138,N_35046,N_35220);
nor U39139 (N_39139,N_35888,N_36707);
and U39140 (N_39140,N_35595,N_35958);
xor U39141 (N_39141,N_35370,N_35063);
xor U39142 (N_39142,N_36256,N_35040);
or U39143 (N_39143,N_35741,N_35943);
or U39144 (N_39144,N_36972,N_37411);
or U39145 (N_39145,N_36765,N_35587);
xor U39146 (N_39146,N_35449,N_35619);
xnor U39147 (N_39147,N_36941,N_36219);
nor U39148 (N_39148,N_37247,N_35248);
nor U39149 (N_39149,N_36118,N_37172);
nor U39150 (N_39150,N_36490,N_36182);
nand U39151 (N_39151,N_37467,N_37098);
nand U39152 (N_39152,N_36937,N_37354);
or U39153 (N_39153,N_36616,N_35668);
or U39154 (N_39154,N_36138,N_35393);
and U39155 (N_39155,N_36817,N_37097);
or U39156 (N_39156,N_36607,N_35753);
and U39157 (N_39157,N_36166,N_35452);
or U39158 (N_39158,N_36495,N_35800);
nand U39159 (N_39159,N_35858,N_36303);
and U39160 (N_39160,N_36922,N_36665);
xnor U39161 (N_39161,N_35508,N_35837);
nor U39162 (N_39162,N_36114,N_35209);
or U39163 (N_39163,N_35149,N_36893);
xnor U39164 (N_39164,N_35467,N_36732);
and U39165 (N_39165,N_35282,N_36196);
nor U39166 (N_39166,N_36339,N_35626);
or U39167 (N_39167,N_35956,N_35875);
or U39168 (N_39168,N_36649,N_35464);
and U39169 (N_39169,N_35583,N_35987);
xor U39170 (N_39170,N_36473,N_36453);
and U39171 (N_39171,N_36277,N_35788);
or U39172 (N_39172,N_35625,N_35344);
and U39173 (N_39173,N_36805,N_35783);
and U39174 (N_39174,N_35768,N_35619);
nor U39175 (N_39175,N_35563,N_36608);
nor U39176 (N_39176,N_35556,N_35741);
nand U39177 (N_39177,N_36079,N_36516);
xnor U39178 (N_39178,N_35335,N_36494);
or U39179 (N_39179,N_37325,N_37346);
xor U39180 (N_39180,N_36361,N_36121);
xor U39181 (N_39181,N_35686,N_37192);
nand U39182 (N_39182,N_36358,N_36355);
nand U39183 (N_39183,N_35935,N_35201);
xor U39184 (N_39184,N_36305,N_36196);
nor U39185 (N_39185,N_35615,N_35774);
xnor U39186 (N_39186,N_35209,N_36632);
nand U39187 (N_39187,N_35676,N_36902);
nand U39188 (N_39188,N_35300,N_35342);
xor U39189 (N_39189,N_37205,N_35867);
nor U39190 (N_39190,N_37482,N_36206);
xnor U39191 (N_39191,N_36054,N_36282);
xor U39192 (N_39192,N_36408,N_36152);
xnor U39193 (N_39193,N_35928,N_35678);
and U39194 (N_39194,N_36818,N_37020);
or U39195 (N_39195,N_36651,N_36693);
and U39196 (N_39196,N_35638,N_35000);
nand U39197 (N_39197,N_36908,N_35984);
and U39198 (N_39198,N_36441,N_37181);
xor U39199 (N_39199,N_35470,N_37248);
and U39200 (N_39200,N_35922,N_37077);
or U39201 (N_39201,N_36987,N_36067);
xor U39202 (N_39202,N_35398,N_36547);
xnor U39203 (N_39203,N_36159,N_37450);
xor U39204 (N_39204,N_36641,N_35844);
and U39205 (N_39205,N_36312,N_35553);
and U39206 (N_39206,N_35332,N_35576);
nor U39207 (N_39207,N_36449,N_37171);
and U39208 (N_39208,N_35200,N_35880);
xor U39209 (N_39209,N_35686,N_36261);
or U39210 (N_39210,N_36777,N_35374);
nor U39211 (N_39211,N_37332,N_35682);
xor U39212 (N_39212,N_36136,N_37412);
and U39213 (N_39213,N_35187,N_35687);
nand U39214 (N_39214,N_35224,N_35059);
nor U39215 (N_39215,N_35718,N_35100);
or U39216 (N_39216,N_37339,N_36210);
xor U39217 (N_39217,N_36239,N_37164);
or U39218 (N_39218,N_35004,N_35922);
or U39219 (N_39219,N_36910,N_36068);
or U39220 (N_39220,N_35961,N_37251);
nor U39221 (N_39221,N_36698,N_35348);
nor U39222 (N_39222,N_36885,N_35129);
or U39223 (N_39223,N_35302,N_35884);
nor U39224 (N_39224,N_36151,N_36271);
and U39225 (N_39225,N_37189,N_35141);
xnor U39226 (N_39226,N_36567,N_36980);
xnor U39227 (N_39227,N_36337,N_36383);
nor U39228 (N_39228,N_35491,N_37028);
or U39229 (N_39229,N_37395,N_35492);
nor U39230 (N_39230,N_35786,N_35911);
nor U39231 (N_39231,N_35724,N_35015);
nand U39232 (N_39232,N_36220,N_37116);
and U39233 (N_39233,N_37286,N_35637);
and U39234 (N_39234,N_35152,N_36686);
xor U39235 (N_39235,N_37136,N_35525);
nor U39236 (N_39236,N_35882,N_37391);
nor U39237 (N_39237,N_36616,N_37253);
nor U39238 (N_39238,N_37261,N_35580);
nor U39239 (N_39239,N_37415,N_36219);
or U39240 (N_39240,N_37372,N_35725);
nand U39241 (N_39241,N_36462,N_36800);
or U39242 (N_39242,N_35983,N_37415);
nor U39243 (N_39243,N_35645,N_35305);
or U39244 (N_39244,N_36200,N_37201);
and U39245 (N_39245,N_37185,N_36246);
and U39246 (N_39246,N_37073,N_35654);
nor U39247 (N_39247,N_36153,N_36224);
nor U39248 (N_39248,N_35240,N_36732);
and U39249 (N_39249,N_36785,N_36822);
or U39250 (N_39250,N_36333,N_36341);
xnor U39251 (N_39251,N_35568,N_35904);
xnor U39252 (N_39252,N_36031,N_35589);
and U39253 (N_39253,N_36641,N_36111);
nor U39254 (N_39254,N_37406,N_35757);
and U39255 (N_39255,N_36379,N_35826);
nor U39256 (N_39256,N_35349,N_37441);
or U39257 (N_39257,N_35669,N_35079);
nor U39258 (N_39258,N_37359,N_36251);
and U39259 (N_39259,N_35344,N_36527);
nand U39260 (N_39260,N_36267,N_35801);
nor U39261 (N_39261,N_37311,N_35879);
nor U39262 (N_39262,N_35282,N_35108);
xor U39263 (N_39263,N_36500,N_35584);
or U39264 (N_39264,N_36655,N_36602);
nor U39265 (N_39265,N_35651,N_35376);
nand U39266 (N_39266,N_37406,N_35990);
xnor U39267 (N_39267,N_36778,N_35229);
or U39268 (N_39268,N_37101,N_36493);
and U39269 (N_39269,N_35971,N_35283);
nor U39270 (N_39270,N_37221,N_35465);
and U39271 (N_39271,N_37134,N_35327);
or U39272 (N_39272,N_36598,N_36399);
or U39273 (N_39273,N_37462,N_36015);
or U39274 (N_39274,N_36475,N_35058);
nand U39275 (N_39275,N_36312,N_36264);
or U39276 (N_39276,N_35102,N_36171);
and U39277 (N_39277,N_36059,N_36463);
xor U39278 (N_39278,N_36019,N_37378);
and U39279 (N_39279,N_36395,N_37098);
nand U39280 (N_39280,N_36554,N_37379);
xnor U39281 (N_39281,N_36658,N_36064);
and U39282 (N_39282,N_36370,N_35121);
nand U39283 (N_39283,N_36276,N_37159);
xor U39284 (N_39284,N_35523,N_35290);
xor U39285 (N_39285,N_35370,N_37204);
nand U39286 (N_39286,N_35341,N_35448);
or U39287 (N_39287,N_35363,N_36046);
or U39288 (N_39288,N_36669,N_36580);
nor U39289 (N_39289,N_36636,N_36520);
and U39290 (N_39290,N_36048,N_36868);
nor U39291 (N_39291,N_35213,N_35361);
and U39292 (N_39292,N_37190,N_35193);
nor U39293 (N_39293,N_35959,N_36577);
nor U39294 (N_39294,N_35982,N_37187);
nand U39295 (N_39295,N_36495,N_35854);
and U39296 (N_39296,N_36540,N_37498);
nand U39297 (N_39297,N_36921,N_35281);
nand U39298 (N_39298,N_36740,N_35364);
and U39299 (N_39299,N_35382,N_36524);
or U39300 (N_39300,N_37285,N_35480);
nand U39301 (N_39301,N_36803,N_36559);
xnor U39302 (N_39302,N_36214,N_37306);
nor U39303 (N_39303,N_35761,N_35613);
and U39304 (N_39304,N_37135,N_36309);
and U39305 (N_39305,N_37444,N_36177);
or U39306 (N_39306,N_36279,N_35108);
xnor U39307 (N_39307,N_37097,N_36833);
and U39308 (N_39308,N_36804,N_36947);
nor U39309 (N_39309,N_36031,N_35891);
xnor U39310 (N_39310,N_35122,N_37493);
and U39311 (N_39311,N_37439,N_35611);
or U39312 (N_39312,N_35418,N_35664);
nand U39313 (N_39313,N_37043,N_35479);
xor U39314 (N_39314,N_36019,N_35152);
and U39315 (N_39315,N_37171,N_36350);
nand U39316 (N_39316,N_37247,N_37460);
or U39317 (N_39317,N_36071,N_37309);
and U39318 (N_39318,N_36413,N_36878);
nor U39319 (N_39319,N_36418,N_36090);
or U39320 (N_39320,N_36352,N_35530);
nand U39321 (N_39321,N_36080,N_37039);
and U39322 (N_39322,N_35949,N_35132);
or U39323 (N_39323,N_35647,N_35337);
nand U39324 (N_39324,N_36551,N_36898);
nand U39325 (N_39325,N_35872,N_36703);
or U39326 (N_39326,N_35975,N_36728);
or U39327 (N_39327,N_37064,N_36826);
and U39328 (N_39328,N_36517,N_35219);
xnor U39329 (N_39329,N_35614,N_37103);
nor U39330 (N_39330,N_36437,N_36645);
xnor U39331 (N_39331,N_36030,N_36715);
nand U39332 (N_39332,N_36933,N_35087);
nor U39333 (N_39333,N_36567,N_37495);
nand U39334 (N_39334,N_35169,N_36237);
xor U39335 (N_39335,N_37025,N_35498);
nand U39336 (N_39336,N_35026,N_35666);
nor U39337 (N_39337,N_35833,N_36236);
and U39338 (N_39338,N_35576,N_36826);
and U39339 (N_39339,N_36168,N_36761);
nand U39340 (N_39340,N_35856,N_35615);
nand U39341 (N_39341,N_36893,N_35830);
and U39342 (N_39342,N_35436,N_35917);
nand U39343 (N_39343,N_36844,N_35462);
or U39344 (N_39344,N_36711,N_35905);
nor U39345 (N_39345,N_36457,N_37228);
nand U39346 (N_39346,N_36236,N_36945);
or U39347 (N_39347,N_36532,N_36947);
nand U39348 (N_39348,N_36035,N_37121);
and U39349 (N_39349,N_36521,N_37142);
xor U39350 (N_39350,N_35100,N_37253);
or U39351 (N_39351,N_37161,N_36210);
nand U39352 (N_39352,N_37355,N_35414);
xor U39353 (N_39353,N_37434,N_36122);
nor U39354 (N_39354,N_37296,N_35282);
nor U39355 (N_39355,N_35387,N_36457);
nor U39356 (N_39356,N_36169,N_35549);
nand U39357 (N_39357,N_35918,N_35995);
or U39358 (N_39358,N_36685,N_35026);
or U39359 (N_39359,N_36949,N_36426);
nor U39360 (N_39360,N_35078,N_36442);
and U39361 (N_39361,N_36212,N_36123);
and U39362 (N_39362,N_36297,N_37080);
nor U39363 (N_39363,N_36829,N_36015);
nor U39364 (N_39364,N_35945,N_37280);
nand U39365 (N_39365,N_36277,N_35443);
nor U39366 (N_39366,N_36410,N_37141);
or U39367 (N_39367,N_37257,N_37370);
and U39368 (N_39368,N_36757,N_36606);
and U39369 (N_39369,N_35369,N_36516);
nand U39370 (N_39370,N_35820,N_36336);
nor U39371 (N_39371,N_35128,N_35467);
nor U39372 (N_39372,N_37486,N_35494);
nor U39373 (N_39373,N_36233,N_37049);
or U39374 (N_39374,N_36738,N_37457);
xor U39375 (N_39375,N_35375,N_36844);
and U39376 (N_39376,N_35013,N_36275);
nor U39377 (N_39377,N_36457,N_36012);
nand U39378 (N_39378,N_36736,N_37349);
and U39379 (N_39379,N_37059,N_35230);
xor U39380 (N_39380,N_37441,N_37022);
nor U39381 (N_39381,N_37150,N_36730);
or U39382 (N_39382,N_36267,N_35970);
nor U39383 (N_39383,N_35918,N_37190);
nand U39384 (N_39384,N_35293,N_37471);
nand U39385 (N_39385,N_36222,N_36744);
nor U39386 (N_39386,N_36784,N_37330);
nor U39387 (N_39387,N_37146,N_36873);
xor U39388 (N_39388,N_36074,N_37241);
nor U39389 (N_39389,N_36696,N_37406);
and U39390 (N_39390,N_37017,N_36793);
or U39391 (N_39391,N_35744,N_35357);
nor U39392 (N_39392,N_35203,N_35250);
or U39393 (N_39393,N_37151,N_37471);
xor U39394 (N_39394,N_36932,N_36261);
or U39395 (N_39395,N_37383,N_37387);
nand U39396 (N_39396,N_35079,N_36955);
and U39397 (N_39397,N_36597,N_35749);
xnor U39398 (N_39398,N_37192,N_35787);
or U39399 (N_39399,N_35489,N_35642);
xor U39400 (N_39400,N_35802,N_35428);
and U39401 (N_39401,N_35081,N_35296);
and U39402 (N_39402,N_37047,N_35835);
and U39403 (N_39403,N_35208,N_37015);
nor U39404 (N_39404,N_36930,N_36751);
and U39405 (N_39405,N_35886,N_37121);
and U39406 (N_39406,N_36351,N_36765);
and U39407 (N_39407,N_36021,N_35482);
nor U39408 (N_39408,N_37056,N_36978);
xor U39409 (N_39409,N_35112,N_35263);
and U39410 (N_39410,N_36507,N_36350);
nand U39411 (N_39411,N_36126,N_35104);
nand U39412 (N_39412,N_35673,N_36624);
and U39413 (N_39413,N_35729,N_36197);
nor U39414 (N_39414,N_36079,N_36993);
and U39415 (N_39415,N_37213,N_35513);
or U39416 (N_39416,N_35414,N_35374);
nor U39417 (N_39417,N_35963,N_36692);
nand U39418 (N_39418,N_35359,N_35832);
xnor U39419 (N_39419,N_35317,N_35689);
nand U39420 (N_39420,N_35839,N_36429);
nand U39421 (N_39421,N_36858,N_37228);
nor U39422 (N_39422,N_37422,N_36523);
xor U39423 (N_39423,N_36085,N_37415);
xnor U39424 (N_39424,N_35218,N_37435);
or U39425 (N_39425,N_35704,N_36614);
nand U39426 (N_39426,N_36125,N_35077);
xor U39427 (N_39427,N_36849,N_36430);
or U39428 (N_39428,N_35962,N_36040);
and U39429 (N_39429,N_36173,N_36981);
and U39430 (N_39430,N_35876,N_36070);
nand U39431 (N_39431,N_35064,N_35617);
or U39432 (N_39432,N_36720,N_35104);
nor U39433 (N_39433,N_37469,N_35700);
or U39434 (N_39434,N_35486,N_35159);
xor U39435 (N_39435,N_36792,N_35367);
xnor U39436 (N_39436,N_35658,N_35522);
xnor U39437 (N_39437,N_35279,N_35042);
and U39438 (N_39438,N_37292,N_35540);
and U39439 (N_39439,N_35919,N_35331);
nand U39440 (N_39440,N_36848,N_36931);
xor U39441 (N_39441,N_36867,N_37269);
xor U39442 (N_39442,N_36558,N_36696);
or U39443 (N_39443,N_37034,N_36133);
and U39444 (N_39444,N_36778,N_36414);
xnor U39445 (N_39445,N_35097,N_36128);
and U39446 (N_39446,N_37088,N_36572);
and U39447 (N_39447,N_35676,N_37028);
xor U39448 (N_39448,N_35231,N_35699);
nor U39449 (N_39449,N_36706,N_35685);
xor U39450 (N_39450,N_35069,N_37346);
nand U39451 (N_39451,N_36938,N_36309);
xor U39452 (N_39452,N_35446,N_35326);
nand U39453 (N_39453,N_36640,N_35797);
nor U39454 (N_39454,N_36895,N_35012);
nand U39455 (N_39455,N_35678,N_35870);
or U39456 (N_39456,N_35423,N_37034);
nor U39457 (N_39457,N_36221,N_36824);
nand U39458 (N_39458,N_35999,N_36119);
nand U39459 (N_39459,N_35071,N_35597);
xor U39460 (N_39460,N_37333,N_37240);
xnor U39461 (N_39461,N_36134,N_35485);
or U39462 (N_39462,N_35076,N_37008);
and U39463 (N_39463,N_35025,N_35558);
nor U39464 (N_39464,N_35585,N_36251);
or U39465 (N_39465,N_35053,N_37311);
nand U39466 (N_39466,N_36494,N_35830);
and U39467 (N_39467,N_35612,N_37082);
nor U39468 (N_39468,N_36902,N_35173);
nand U39469 (N_39469,N_35189,N_35289);
and U39470 (N_39470,N_36346,N_36116);
and U39471 (N_39471,N_35128,N_36427);
nor U39472 (N_39472,N_35397,N_37248);
xnor U39473 (N_39473,N_36658,N_37385);
or U39474 (N_39474,N_37442,N_35142);
and U39475 (N_39475,N_35579,N_37394);
and U39476 (N_39476,N_36708,N_36529);
xor U39477 (N_39477,N_36485,N_37372);
nor U39478 (N_39478,N_37313,N_35324);
nand U39479 (N_39479,N_35070,N_35988);
xor U39480 (N_39480,N_36140,N_36727);
or U39481 (N_39481,N_35689,N_35740);
xnor U39482 (N_39482,N_36170,N_35996);
and U39483 (N_39483,N_35749,N_35632);
or U39484 (N_39484,N_36767,N_36293);
and U39485 (N_39485,N_37078,N_35328);
nor U39486 (N_39486,N_36297,N_36003);
and U39487 (N_39487,N_35445,N_36519);
and U39488 (N_39488,N_36281,N_35013);
or U39489 (N_39489,N_36527,N_36132);
nor U39490 (N_39490,N_37408,N_35193);
or U39491 (N_39491,N_36959,N_37178);
nand U39492 (N_39492,N_35385,N_37080);
nand U39493 (N_39493,N_37132,N_37447);
and U39494 (N_39494,N_36045,N_35130);
xnor U39495 (N_39495,N_36190,N_35985);
xnor U39496 (N_39496,N_35028,N_35383);
xnor U39497 (N_39497,N_37176,N_37075);
or U39498 (N_39498,N_37202,N_36589);
nor U39499 (N_39499,N_36677,N_36697);
xor U39500 (N_39500,N_36474,N_35037);
or U39501 (N_39501,N_36695,N_36726);
and U39502 (N_39502,N_37404,N_36875);
xor U39503 (N_39503,N_37425,N_35130);
nor U39504 (N_39504,N_36044,N_36355);
nor U39505 (N_39505,N_35150,N_37111);
xor U39506 (N_39506,N_36121,N_35647);
or U39507 (N_39507,N_35865,N_36025);
and U39508 (N_39508,N_35959,N_35728);
or U39509 (N_39509,N_35248,N_35233);
or U39510 (N_39510,N_35745,N_36383);
xnor U39511 (N_39511,N_36096,N_36539);
and U39512 (N_39512,N_36687,N_35549);
and U39513 (N_39513,N_36230,N_36049);
xnor U39514 (N_39514,N_35675,N_36659);
nand U39515 (N_39515,N_35476,N_36384);
and U39516 (N_39516,N_35043,N_36538);
nor U39517 (N_39517,N_36224,N_37356);
xnor U39518 (N_39518,N_35665,N_35269);
nor U39519 (N_39519,N_35626,N_36419);
nand U39520 (N_39520,N_37133,N_35583);
and U39521 (N_39521,N_35616,N_35930);
or U39522 (N_39522,N_36100,N_36735);
or U39523 (N_39523,N_37489,N_35748);
and U39524 (N_39524,N_37025,N_35805);
nand U39525 (N_39525,N_35843,N_36097);
or U39526 (N_39526,N_37311,N_35845);
nand U39527 (N_39527,N_35354,N_35104);
nor U39528 (N_39528,N_36415,N_35863);
and U39529 (N_39529,N_36297,N_37279);
and U39530 (N_39530,N_35469,N_37370);
nor U39531 (N_39531,N_36445,N_37179);
and U39532 (N_39532,N_36684,N_35587);
and U39533 (N_39533,N_36787,N_36545);
or U39534 (N_39534,N_35472,N_36787);
nand U39535 (N_39535,N_35153,N_36684);
xnor U39536 (N_39536,N_37307,N_35507);
nor U39537 (N_39537,N_35885,N_36990);
xnor U39538 (N_39538,N_35015,N_35333);
nor U39539 (N_39539,N_36398,N_37063);
nand U39540 (N_39540,N_36390,N_36172);
xnor U39541 (N_39541,N_36003,N_35857);
xor U39542 (N_39542,N_36771,N_36977);
xnor U39543 (N_39543,N_37237,N_36186);
nand U39544 (N_39544,N_35057,N_35665);
or U39545 (N_39545,N_35805,N_37490);
or U39546 (N_39546,N_35449,N_36625);
xnor U39547 (N_39547,N_35891,N_37451);
or U39548 (N_39548,N_35440,N_37439);
and U39549 (N_39549,N_35812,N_36239);
nor U39550 (N_39550,N_36928,N_36118);
nor U39551 (N_39551,N_36745,N_36363);
and U39552 (N_39552,N_36334,N_37257);
and U39553 (N_39553,N_36293,N_37016);
and U39554 (N_39554,N_35614,N_35471);
and U39555 (N_39555,N_35164,N_36250);
or U39556 (N_39556,N_37102,N_36186);
nor U39557 (N_39557,N_37465,N_36434);
nand U39558 (N_39558,N_35232,N_36739);
nand U39559 (N_39559,N_35239,N_36538);
and U39560 (N_39560,N_37076,N_37354);
nand U39561 (N_39561,N_35334,N_36344);
xor U39562 (N_39562,N_36125,N_35315);
or U39563 (N_39563,N_35307,N_36711);
nor U39564 (N_39564,N_36628,N_35973);
nand U39565 (N_39565,N_35923,N_35409);
nor U39566 (N_39566,N_35418,N_35279);
nor U39567 (N_39567,N_35767,N_35613);
nor U39568 (N_39568,N_36436,N_36776);
nor U39569 (N_39569,N_36613,N_35296);
or U39570 (N_39570,N_35728,N_35518);
nand U39571 (N_39571,N_35779,N_35951);
nor U39572 (N_39572,N_35663,N_36015);
nand U39573 (N_39573,N_37109,N_35430);
and U39574 (N_39574,N_36321,N_35644);
or U39575 (N_39575,N_35404,N_37495);
nand U39576 (N_39576,N_37353,N_35139);
and U39577 (N_39577,N_36923,N_36011);
or U39578 (N_39578,N_36388,N_37093);
nand U39579 (N_39579,N_35093,N_35294);
nand U39580 (N_39580,N_37120,N_36039);
nor U39581 (N_39581,N_35759,N_35238);
or U39582 (N_39582,N_36904,N_36528);
nor U39583 (N_39583,N_36923,N_35352);
xnor U39584 (N_39584,N_36066,N_36318);
nand U39585 (N_39585,N_35539,N_36422);
xnor U39586 (N_39586,N_35734,N_35889);
nand U39587 (N_39587,N_36614,N_37170);
or U39588 (N_39588,N_35198,N_36371);
or U39589 (N_39589,N_36903,N_37298);
nand U39590 (N_39590,N_35252,N_36460);
or U39591 (N_39591,N_35669,N_37068);
and U39592 (N_39592,N_36736,N_36067);
xnor U39593 (N_39593,N_37464,N_37121);
nand U39594 (N_39594,N_35523,N_37133);
or U39595 (N_39595,N_36727,N_36882);
nand U39596 (N_39596,N_35358,N_35401);
xor U39597 (N_39597,N_36174,N_36559);
or U39598 (N_39598,N_36766,N_37088);
or U39599 (N_39599,N_36982,N_36612);
nand U39600 (N_39600,N_37253,N_37344);
and U39601 (N_39601,N_35717,N_35830);
and U39602 (N_39602,N_35307,N_35386);
or U39603 (N_39603,N_35907,N_35067);
nand U39604 (N_39604,N_35126,N_35324);
nor U39605 (N_39605,N_36229,N_35128);
and U39606 (N_39606,N_36484,N_35640);
nor U39607 (N_39607,N_35385,N_36544);
xor U39608 (N_39608,N_36298,N_36001);
nor U39609 (N_39609,N_35379,N_36261);
nand U39610 (N_39610,N_37467,N_36558);
nor U39611 (N_39611,N_35994,N_36173);
nand U39612 (N_39612,N_35142,N_35875);
or U39613 (N_39613,N_35078,N_35039);
or U39614 (N_39614,N_37364,N_37080);
nor U39615 (N_39615,N_37346,N_36104);
and U39616 (N_39616,N_35874,N_35338);
or U39617 (N_39617,N_36601,N_36623);
or U39618 (N_39618,N_37352,N_36706);
nand U39619 (N_39619,N_36213,N_36434);
nand U39620 (N_39620,N_35744,N_35573);
nor U39621 (N_39621,N_37468,N_35624);
nand U39622 (N_39622,N_35418,N_37041);
or U39623 (N_39623,N_37497,N_36093);
nand U39624 (N_39624,N_36658,N_37375);
nor U39625 (N_39625,N_35761,N_37054);
nor U39626 (N_39626,N_35832,N_37107);
nand U39627 (N_39627,N_35369,N_35703);
nand U39628 (N_39628,N_36456,N_35385);
or U39629 (N_39629,N_35197,N_35480);
or U39630 (N_39630,N_35151,N_37419);
xor U39631 (N_39631,N_35579,N_36692);
nand U39632 (N_39632,N_37211,N_37075);
and U39633 (N_39633,N_36052,N_36112);
and U39634 (N_39634,N_36911,N_35896);
and U39635 (N_39635,N_36186,N_36383);
nand U39636 (N_39636,N_35734,N_36633);
or U39637 (N_39637,N_37235,N_35591);
xnor U39638 (N_39638,N_36102,N_35314);
and U39639 (N_39639,N_36084,N_37371);
nor U39640 (N_39640,N_36811,N_36305);
and U39641 (N_39641,N_36404,N_35871);
or U39642 (N_39642,N_36789,N_35404);
xnor U39643 (N_39643,N_36757,N_36842);
nor U39644 (N_39644,N_36514,N_35967);
nand U39645 (N_39645,N_37427,N_35782);
nand U39646 (N_39646,N_35116,N_35674);
or U39647 (N_39647,N_35985,N_35581);
nor U39648 (N_39648,N_35776,N_35534);
nor U39649 (N_39649,N_35480,N_36955);
or U39650 (N_39650,N_35854,N_35248);
nor U39651 (N_39651,N_35851,N_35650);
nor U39652 (N_39652,N_35667,N_37380);
or U39653 (N_39653,N_35023,N_35924);
xor U39654 (N_39654,N_36972,N_35557);
nand U39655 (N_39655,N_35385,N_36126);
nor U39656 (N_39656,N_35177,N_37422);
or U39657 (N_39657,N_37218,N_36277);
nand U39658 (N_39658,N_36000,N_37439);
or U39659 (N_39659,N_36841,N_37438);
and U39660 (N_39660,N_35436,N_36343);
and U39661 (N_39661,N_35087,N_36596);
nor U39662 (N_39662,N_36037,N_36499);
or U39663 (N_39663,N_37490,N_35647);
nand U39664 (N_39664,N_35391,N_35538);
and U39665 (N_39665,N_35873,N_36296);
xnor U39666 (N_39666,N_36929,N_37120);
and U39667 (N_39667,N_37459,N_35743);
or U39668 (N_39668,N_35485,N_37260);
or U39669 (N_39669,N_36901,N_36487);
or U39670 (N_39670,N_36547,N_37284);
nand U39671 (N_39671,N_35747,N_36005);
nand U39672 (N_39672,N_35244,N_36341);
or U39673 (N_39673,N_36722,N_36320);
nand U39674 (N_39674,N_35333,N_35517);
and U39675 (N_39675,N_36343,N_35994);
or U39676 (N_39676,N_37056,N_37160);
or U39677 (N_39677,N_35937,N_36442);
nand U39678 (N_39678,N_35543,N_36636);
and U39679 (N_39679,N_35385,N_36931);
xnor U39680 (N_39680,N_37425,N_36496);
and U39681 (N_39681,N_37048,N_36508);
nor U39682 (N_39682,N_37105,N_35934);
and U39683 (N_39683,N_36915,N_36585);
nor U39684 (N_39684,N_36303,N_35227);
and U39685 (N_39685,N_35943,N_37181);
and U39686 (N_39686,N_36891,N_37194);
xor U39687 (N_39687,N_35014,N_35591);
nand U39688 (N_39688,N_36917,N_37069);
nand U39689 (N_39689,N_36928,N_37488);
or U39690 (N_39690,N_37029,N_35622);
or U39691 (N_39691,N_37386,N_37373);
xor U39692 (N_39692,N_36076,N_37008);
nor U39693 (N_39693,N_35550,N_37148);
and U39694 (N_39694,N_36478,N_36937);
xnor U39695 (N_39695,N_36624,N_37431);
nor U39696 (N_39696,N_35022,N_35395);
xor U39697 (N_39697,N_36872,N_35238);
nor U39698 (N_39698,N_36847,N_36897);
nor U39699 (N_39699,N_36589,N_35818);
nand U39700 (N_39700,N_36757,N_36060);
nor U39701 (N_39701,N_35455,N_37021);
nand U39702 (N_39702,N_37333,N_35174);
and U39703 (N_39703,N_36318,N_35406);
and U39704 (N_39704,N_37173,N_35255);
nor U39705 (N_39705,N_36834,N_37454);
nand U39706 (N_39706,N_36286,N_35672);
nand U39707 (N_39707,N_35016,N_36327);
and U39708 (N_39708,N_37089,N_36427);
nor U39709 (N_39709,N_37155,N_35241);
nor U39710 (N_39710,N_37318,N_37166);
and U39711 (N_39711,N_36895,N_36938);
xnor U39712 (N_39712,N_35723,N_35196);
nor U39713 (N_39713,N_37296,N_36988);
nand U39714 (N_39714,N_35065,N_36332);
and U39715 (N_39715,N_36338,N_35020);
xnor U39716 (N_39716,N_36706,N_36897);
nand U39717 (N_39717,N_35489,N_36611);
xor U39718 (N_39718,N_35522,N_36138);
nand U39719 (N_39719,N_37179,N_35590);
nand U39720 (N_39720,N_36866,N_37457);
nand U39721 (N_39721,N_37169,N_35255);
nand U39722 (N_39722,N_35609,N_36844);
nor U39723 (N_39723,N_36416,N_35205);
or U39724 (N_39724,N_35058,N_37100);
xor U39725 (N_39725,N_37121,N_35119);
nand U39726 (N_39726,N_35060,N_37057);
or U39727 (N_39727,N_37270,N_36772);
nor U39728 (N_39728,N_37121,N_35140);
nand U39729 (N_39729,N_36001,N_35099);
or U39730 (N_39730,N_36445,N_37249);
xor U39731 (N_39731,N_37332,N_36456);
or U39732 (N_39732,N_37049,N_35134);
nand U39733 (N_39733,N_37366,N_35552);
xor U39734 (N_39734,N_35489,N_35233);
xor U39735 (N_39735,N_35453,N_35374);
or U39736 (N_39736,N_35344,N_36330);
or U39737 (N_39737,N_35881,N_36653);
nand U39738 (N_39738,N_36755,N_35034);
and U39739 (N_39739,N_36760,N_36938);
or U39740 (N_39740,N_35244,N_36844);
or U39741 (N_39741,N_36736,N_35271);
nor U39742 (N_39742,N_35769,N_37319);
or U39743 (N_39743,N_35864,N_35034);
nor U39744 (N_39744,N_36130,N_36650);
nand U39745 (N_39745,N_37233,N_37254);
nand U39746 (N_39746,N_35174,N_35469);
nand U39747 (N_39747,N_35478,N_36698);
nor U39748 (N_39748,N_36751,N_37316);
nand U39749 (N_39749,N_35157,N_37341);
and U39750 (N_39750,N_37133,N_37422);
or U39751 (N_39751,N_35072,N_35565);
and U39752 (N_39752,N_36398,N_37378);
and U39753 (N_39753,N_35054,N_36492);
and U39754 (N_39754,N_37000,N_35546);
xnor U39755 (N_39755,N_36569,N_36253);
and U39756 (N_39756,N_36608,N_37158);
nand U39757 (N_39757,N_36395,N_37116);
nor U39758 (N_39758,N_36036,N_36504);
nor U39759 (N_39759,N_35524,N_36021);
and U39760 (N_39760,N_36330,N_35981);
xnor U39761 (N_39761,N_35469,N_37345);
xor U39762 (N_39762,N_35456,N_36851);
nor U39763 (N_39763,N_35603,N_35218);
xor U39764 (N_39764,N_37423,N_35669);
and U39765 (N_39765,N_36889,N_36723);
nand U39766 (N_39766,N_36344,N_35703);
nand U39767 (N_39767,N_35706,N_36617);
xor U39768 (N_39768,N_36353,N_35990);
and U39769 (N_39769,N_35305,N_36673);
or U39770 (N_39770,N_37344,N_35092);
and U39771 (N_39771,N_35226,N_35845);
and U39772 (N_39772,N_35847,N_37159);
xnor U39773 (N_39773,N_35030,N_37490);
xnor U39774 (N_39774,N_36071,N_35752);
and U39775 (N_39775,N_37180,N_36417);
xor U39776 (N_39776,N_36754,N_36424);
and U39777 (N_39777,N_35498,N_37304);
or U39778 (N_39778,N_37115,N_35192);
xor U39779 (N_39779,N_36581,N_35302);
and U39780 (N_39780,N_35976,N_37180);
xnor U39781 (N_39781,N_36533,N_37421);
nand U39782 (N_39782,N_35028,N_36502);
xnor U39783 (N_39783,N_35261,N_37074);
nand U39784 (N_39784,N_36392,N_36054);
nand U39785 (N_39785,N_36056,N_35931);
nand U39786 (N_39786,N_35555,N_36311);
nand U39787 (N_39787,N_36922,N_35146);
or U39788 (N_39788,N_36715,N_37216);
nor U39789 (N_39789,N_35195,N_36372);
xnor U39790 (N_39790,N_36757,N_37303);
and U39791 (N_39791,N_35768,N_36426);
nand U39792 (N_39792,N_35585,N_36665);
and U39793 (N_39793,N_35316,N_35220);
or U39794 (N_39794,N_36971,N_36713);
nor U39795 (N_39795,N_36100,N_36026);
or U39796 (N_39796,N_36375,N_37126);
or U39797 (N_39797,N_36761,N_36252);
xnor U39798 (N_39798,N_35961,N_35462);
or U39799 (N_39799,N_36379,N_35908);
xnor U39800 (N_39800,N_35545,N_35199);
nand U39801 (N_39801,N_36369,N_35988);
or U39802 (N_39802,N_37002,N_36749);
or U39803 (N_39803,N_35309,N_36245);
nand U39804 (N_39804,N_37226,N_36980);
xnor U39805 (N_39805,N_36128,N_36627);
or U39806 (N_39806,N_37193,N_35364);
xnor U39807 (N_39807,N_35258,N_35739);
nor U39808 (N_39808,N_37031,N_37304);
nor U39809 (N_39809,N_37085,N_37252);
nand U39810 (N_39810,N_35979,N_36331);
nor U39811 (N_39811,N_35219,N_36568);
xor U39812 (N_39812,N_35974,N_36027);
and U39813 (N_39813,N_37039,N_35819);
or U39814 (N_39814,N_35807,N_36523);
xnor U39815 (N_39815,N_37488,N_36760);
or U39816 (N_39816,N_35056,N_36913);
nor U39817 (N_39817,N_36347,N_36305);
nand U39818 (N_39818,N_36901,N_35410);
xor U39819 (N_39819,N_36618,N_36251);
or U39820 (N_39820,N_36529,N_36043);
or U39821 (N_39821,N_36062,N_35801);
nor U39822 (N_39822,N_37034,N_36915);
or U39823 (N_39823,N_36483,N_35525);
nor U39824 (N_39824,N_36471,N_35772);
or U39825 (N_39825,N_36625,N_36063);
xor U39826 (N_39826,N_36830,N_35023);
nor U39827 (N_39827,N_35286,N_36678);
or U39828 (N_39828,N_36572,N_35353);
nor U39829 (N_39829,N_35268,N_37296);
xor U39830 (N_39830,N_35695,N_37069);
nor U39831 (N_39831,N_35093,N_36747);
or U39832 (N_39832,N_37244,N_36596);
or U39833 (N_39833,N_36766,N_35343);
nor U39834 (N_39834,N_35757,N_35646);
nand U39835 (N_39835,N_36281,N_36655);
nor U39836 (N_39836,N_37100,N_35350);
nand U39837 (N_39837,N_37470,N_36113);
xor U39838 (N_39838,N_36485,N_36082);
xnor U39839 (N_39839,N_35429,N_35138);
nand U39840 (N_39840,N_35914,N_36088);
nand U39841 (N_39841,N_35626,N_35023);
xor U39842 (N_39842,N_37059,N_35519);
nand U39843 (N_39843,N_36116,N_35795);
xor U39844 (N_39844,N_35356,N_35073);
nor U39845 (N_39845,N_36552,N_35378);
nand U39846 (N_39846,N_35068,N_35945);
nand U39847 (N_39847,N_36243,N_35706);
nor U39848 (N_39848,N_37012,N_36186);
xor U39849 (N_39849,N_35232,N_36727);
and U39850 (N_39850,N_36784,N_35844);
and U39851 (N_39851,N_37450,N_35345);
nand U39852 (N_39852,N_36755,N_35846);
nand U39853 (N_39853,N_37188,N_35128);
nand U39854 (N_39854,N_36073,N_36128);
xnor U39855 (N_39855,N_37271,N_35227);
nor U39856 (N_39856,N_36376,N_35637);
nand U39857 (N_39857,N_36750,N_36374);
nand U39858 (N_39858,N_37095,N_37079);
nand U39859 (N_39859,N_35847,N_36132);
nand U39860 (N_39860,N_35740,N_35019);
nor U39861 (N_39861,N_36033,N_35020);
xor U39862 (N_39862,N_37473,N_36962);
xnor U39863 (N_39863,N_35967,N_35748);
xor U39864 (N_39864,N_37361,N_35452);
nand U39865 (N_39865,N_37027,N_37271);
xor U39866 (N_39866,N_36188,N_36576);
nor U39867 (N_39867,N_35991,N_35477);
nand U39868 (N_39868,N_35086,N_36803);
nand U39869 (N_39869,N_36224,N_35942);
xnor U39870 (N_39870,N_37463,N_37166);
and U39871 (N_39871,N_36488,N_36445);
xnor U39872 (N_39872,N_35524,N_36524);
and U39873 (N_39873,N_37386,N_36564);
or U39874 (N_39874,N_36212,N_36452);
nand U39875 (N_39875,N_36702,N_36560);
and U39876 (N_39876,N_36663,N_35793);
and U39877 (N_39877,N_36261,N_36861);
and U39878 (N_39878,N_36795,N_35824);
nand U39879 (N_39879,N_37476,N_36153);
and U39880 (N_39880,N_36593,N_35863);
or U39881 (N_39881,N_36731,N_35641);
nor U39882 (N_39882,N_37070,N_36332);
nor U39883 (N_39883,N_36783,N_35649);
and U39884 (N_39884,N_35481,N_37066);
nor U39885 (N_39885,N_35432,N_36145);
nor U39886 (N_39886,N_36418,N_35048);
or U39887 (N_39887,N_37241,N_37329);
nor U39888 (N_39888,N_35508,N_37422);
or U39889 (N_39889,N_36224,N_35999);
xor U39890 (N_39890,N_35687,N_35041);
nor U39891 (N_39891,N_35066,N_37303);
or U39892 (N_39892,N_35850,N_35691);
and U39893 (N_39893,N_35265,N_36519);
xor U39894 (N_39894,N_37445,N_36340);
and U39895 (N_39895,N_36862,N_36520);
xnor U39896 (N_39896,N_35696,N_36991);
nand U39897 (N_39897,N_35792,N_36911);
nand U39898 (N_39898,N_35216,N_35915);
nor U39899 (N_39899,N_36643,N_37085);
xor U39900 (N_39900,N_35095,N_36696);
xnor U39901 (N_39901,N_36087,N_35885);
or U39902 (N_39902,N_37177,N_37415);
and U39903 (N_39903,N_36984,N_36256);
nand U39904 (N_39904,N_35407,N_36565);
xor U39905 (N_39905,N_36866,N_35607);
or U39906 (N_39906,N_35637,N_36852);
xor U39907 (N_39907,N_36606,N_35813);
and U39908 (N_39908,N_35679,N_35859);
xnor U39909 (N_39909,N_36829,N_36251);
nand U39910 (N_39910,N_35986,N_35400);
nand U39911 (N_39911,N_37292,N_36027);
or U39912 (N_39912,N_36530,N_36409);
xor U39913 (N_39913,N_36717,N_36578);
and U39914 (N_39914,N_36875,N_37020);
nand U39915 (N_39915,N_37423,N_37204);
and U39916 (N_39916,N_35742,N_35612);
or U39917 (N_39917,N_35061,N_36908);
nand U39918 (N_39918,N_35845,N_36387);
or U39919 (N_39919,N_36502,N_35161);
or U39920 (N_39920,N_37061,N_35406);
xnor U39921 (N_39921,N_36718,N_36766);
nor U39922 (N_39922,N_37141,N_36011);
or U39923 (N_39923,N_35582,N_37148);
xor U39924 (N_39924,N_35345,N_37499);
nor U39925 (N_39925,N_36878,N_36514);
xor U39926 (N_39926,N_36972,N_35351);
nand U39927 (N_39927,N_35233,N_36778);
or U39928 (N_39928,N_36286,N_35576);
xnor U39929 (N_39929,N_35870,N_36111);
and U39930 (N_39930,N_37049,N_36893);
xor U39931 (N_39931,N_36371,N_35321);
nor U39932 (N_39932,N_36506,N_37038);
and U39933 (N_39933,N_37118,N_35892);
and U39934 (N_39934,N_36711,N_36020);
xnor U39935 (N_39935,N_36068,N_35489);
nor U39936 (N_39936,N_36927,N_35520);
and U39937 (N_39937,N_35745,N_35599);
or U39938 (N_39938,N_35044,N_37090);
nand U39939 (N_39939,N_35398,N_36856);
nor U39940 (N_39940,N_37012,N_36628);
xor U39941 (N_39941,N_36152,N_37411);
nand U39942 (N_39942,N_37025,N_36211);
nand U39943 (N_39943,N_35067,N_35333);
xnor U39944 (N_39944,N_36766,N_36324);
and U39945 (N_39945,N_35769,N_35492);
or U39946 (N_39946,N_35284,N_35267);
nor U39947 (N_39947,N_36195,N_35338);
nor U39948 (N_39948,N_36705,N_36531);
xor U39949 (N_39949,N_37143,N_35436);
or U39950 (N_39950,N_37321,N_37445);
nor U39951 (N_39951,N_35436,N_35722);
and U39952 (N_39952,N_35269,N_36132);
xor U39953 (N_39953,N_35646,N_35259);
and U39954 (N_39954,N_35435,N_35715);
and U39955 (N_39955,N_35003,N_35934);
xnor U39956 (N_39956,N_35040,N_35890);
nor U39957 (N_39957,N_36973,N_36437);
nor U39958 (N_39958,N_35577,N_35299);
xor U39959 (N_39959,N_36716,N_37202);
xnor U39960 (N_39960,N_35932,N_36479);
or U39961 (N_39961,N_35379,N_37089);
xnor U39962 (N_39962,N_36104,N_37074);
and U39963 (N_39963,N_35209,N_36400);
nand U39964 (N_39964,N_35300,N_35663);
nand U39965 (N_39965,N_35030,N_37123);
or U39966 (N_39966,N_35610,N_35045);
nor U39967 (N_39967,N_35157,N_36899);
nand U39968 (N_39968,N_36911,N_35229);
and U39969 (N_39969,N_36892,N_36579);
xnor U39970 (N_39970,N_37236,N_35412);
nand U39971 (N_39971,N_36972,N_37112);
nor U39972 (N_39972,N_35815,N_36334);
nand U39973 (N_39973,N_37083,N_36983);
nor U39974 (N_39974,N_36084,N_35633);
xnor U39975 (N_39975,N_35764,N_37328);
nor U39976 (N_39976,N_35851,N_35117);
nand U39977 (N_39977,N_37040,N_36309);
and U39978 (N_39978,N_35710,N_36279);
nor U39979 (N_39979,N_36462,N_36153);
nand U39980 (N_39980,N_36603,N_36112);
nand U39981 (N_39981,N_36962,N_36417);
xnor U39982 (N_39982,N_36728,N_36020);
nand U39983 (N_39983,N_37052,N_36811);
or U39984 (N_39984,N_36690,N_37185);
or U39985 (N_39985,N_36209,N_37467);
nand U39986 (N_39986,N_36869,N_36227);
nor U39987 (N_39987,N_37333,N_36727);
or U39988 (N_39988,N_35255,N_37013);
or U39989 (N_39989,N_35795,N_35550);
or U39990 (N_39990,N_35863,N_36276);
nor U39991 (N_39991,N_36077,N_35977);
nand U39992 (N_39992,N_35533,N_35961);
nand U39993 (N_39993,N_35082,N_36743);
nand U39994 (N_39994,N_36171,N_35581);
nand U39995 (N_39995,N_36397,N_35718);
and U39996 (N_39996,N_36815,N_37152);
nand U39997 (N_39997,N_35432,N_35212);
nor U39998 (N_39998,N_35496,N_36397);
nand U39999 (N_39999,N_37087,N_36763);
xnor U40000 (N_40000,N_37625,N_39083);
and U40001 (N_40001,N_38367,N_38083);
and U40002 (N_40002,N_39466,N_38978);
xnor U40003 (N_40003,N_39512,N_37721);
xnor U40004 (N_40004,N_38744,N_39582);
nand U40005 (N_40005,N_38248,N_37783);
or U40006 (N_40006,N_39013,N_39643);
nor U40007 (N_40007,N_37997,N_37774);
or U40008 (N_40008,N_39758,N_39366);
and U40009 (N_40009,N_38280,N_39952);
and U40010 (N_40010,N_39750,N_39834);
nand U40011 (N_40011,N_38608,N_37862);
nand U40012 (N_40012,N_39222,N_39398);
nand U40013 (N_40013,N_37856,N_39339);
nand U40014 (N_40014,N_38737,N_37697);
xor U40015 (N_40015,N_37883,N_38579);
nor U40016 (N_40016,N_38309,N_38164);
nand U40017 (N_40017,N_39575,N_38637);
nor U40018 (N_40018,N_38038,N_37849);
nor U40019 (N_40019,N_37521,N_39263);
and U40020 (N_40020,N_38117,N_39132);
nand U40021 (N_40021,N_37688,N_38994);
and U40022 (N_40022,N_39184,N_37946);
and U40023 (N_40023,N_39298,N_39346);
nand U40024 (N_40024,N_39563,N_39247);
nand U40025 (N_40025,N_39252,N_37800);
or U40026 (N_40026,N_37757,N_39026);
nor U40027 (N_40027,N_39332,N_39790);
or U40028 (N_40028,N_37571,N_38125);
xor U40029 (N_40029,N_39255,N_38364);
nor U40030 (N_40030,N_39015,N_37704);
xor U40031 (N_40031,N_38497,N_39814);
nand U40032 (N_40032,N_38318,N_37799);
and U40033 (N_40033,N_39186,N_38936);
nor U40034 (N_40034,N_38422,N_38738);
nor U40035 (N_40035,N_38640,N_38271);
nor U40036 (N_40036,N_37941,N_39437);
xor U40037 (N_40037,N_39793,N_39772);
nand U40038 (N_40038,N_39344,N_38003);
or U40039 (N_40039,N_38325,N_37661);
or U40040 (N_40040,N_39097,N_37846);
nand U40041 (N_40041,N_39125,N_39014);
nand U40042 (N_40042,N_37879,N_39858);
nor U40043 (N_40043,N_39562,N_37620);
nor U40044 (N_40044,N_37703,N_38577);
and U40045 (N_40045,N_39345,N_38075);
xnor U40046 (N_40046,N_39866,N_39987);
and U40047 (N_40047,N_37589,N_37985);
xnor U40048 (N_40048,N_38594,N_38473);
or U40049 (N_40049,N_37554,N_37833);
nor U40050 (N_40050,N_38867,N_38948);
or U40051 (N_40051,N_39274,N_39962);
xnor U40052 (N_40052,N_38079,N_39146);
nor U40053 (N_40053,N_37788,N_38427);
and U40054 (N_40054,N_39386,N_39107);
xor U40055 (N_40055,N_39913,N_38006);
xor U40056 (N_40056,N_39804,N_39170);
or U40057 (N_40057,N_39285,N_38277);
or U40058 (N_40058,N_38301,N_39825);
nand U40059 (N_40059,N_38055,N_38910);
or U40060 (N_40060,N_37926,N_37951);
nand U40061 (N_40061,N_39100,N_38952);
nand U40062 (N_40062,N_38760,N_38890);
xnor U40063 (N_40063,N_39579,N_38505);
and U40064 (N_40064,N_38287,N_39592);
xor U40065 (N_40065,N_38415,N_39304);
or U40066 (N_40066,N_39647,N_39686);
nor U40067 (N_40067,N_38487,N_38391);
or U40068 (N_40068,N_37715,N_39526);
nor U40069 (N_40069,N_37840,N_39728);
nand U40070 (N_40070,N_38866,N_37780);
xnor U40071 (N_40071,N_38990,N_38908);
xor U40072 (N_40072,N_39847,N_37513);
xnor U40073 (N_40073,N_39240,N_39150);
nor U40074 (N_40074,N_39494,N_38369);
nor U40075 (N_40075,N_39432,N_38719);
xnor U40076 (N_40076,N_37515,N_38360);
or U40077 (N_40077,N_39017,N_38884);
nor U40078 (N_40078,N_38353,N_38781);
or U40079 (N_40079,N_39042,N_37938);
xor U40080 (N_40080,N_37547,N_38530);
nand U40081 (N_40081,N_38545,N_38976);
nor U40082 (N_40082,N_39970,N_37669);
nor U40083 (N_40083,N_38447,N_39397);
nand U40084 (N_40084,N_38950,N_39675);
or U40085 (N_40085,N_38587,N_39223);
and U40086 (N_40086,N_38971,N_38151);
xor U40087 (N_40087,N_38389,N_39444);
nor U40088 (N_40088,N_39238,N_39160);
xnor U40089 (N_40089,N_38892,N_39764);
and U40090 (N_40090,N_39785,N_38157);
and U40091 (N_40091,N_37742,N_39174);
or U40092 (N_40092,N_37972,N_38399);
and U40093 (N_40093,N_38897,N_37709);
nand U40094 (N_40094,N_39771,N_38928);
or U40095 (N_40095,N_38463,N_37749);
nor U40096 (N_40096,N_38670,N_38090);
nand U40097 (N_40097,N_38762,N_38663);
or U40098 (N_40098,N_38102,N_38105);
nand U40099 (N_40099,N_37698,N_38642);
nand U40100 (N_40100,N_38929,N_39354);
and U40101 (N_40101,N_39951,N_38787);
or U40102 (N_40102,N_39896,N_38080);
nor U40103 (N_40103,N_39551,N_39571);
nand U40104 (N_40104,N_38288,N_39634);
and U40105 (N_40105,N_37700,N_37878);
and U40106 (N_40106,N_38882,N_38334);
or U40107 (N_40107,N_37930,N_37854);
nor U40108 (N_40108,N_38158,N_37586);
nand U40109 (N_40109,N_39070,N_39038);
nand U40110 (N_40110,N_37762,N_38124);
or U40111 (N_40111,N_39064,N_38071);
or U40112 (N_40112,N_39450,N_39802);
or U40113 (N_40113,N_38667,N_39996);
xnor U40114 (N_40114,N_38534,N_37570);
or U40115 (N_40115,N_37936,N_39650);
xor U40116 (N_40116,N_38464,N_37577);
and U40117 (N_40117,N_38911,N_37811);
and U40118 (N_40118,N_39018,N_38688);
and U40119 (N_40119,N_37518,N_39917);
nor U40120 (N_40120,N_39608,N_37770);
and U40121 (N_40121,N_39370,N_38173);
xor U40122 (N_40122,N_37502,N_39912);
xnor U40123 (N_40123,N_37771,N_39388);
or U40124 (N_40124,N_38586,N_39248);
xnor U40125 (N_40125,N_38380,N_37587);
nand U40126 (N_40126,N_38596,N_39969);
nand U40127 (N_40127,N_39200,N_39074);
or U40128 (N_40128,N_39715,N_39947);
and U40129 (N_40129,N_37575,N_39697);
nor U40130 (N_40130,N_38436,N_39309);
and U40131 (N_40131,N_38032,N_38664);
nor U40132 (N_40132,N_39929,N_39975);
and U40133 (N_40133,N_39135,N_38120);
or U40134 (N_40134,N_37973,N_39747);
xor U40135 (N_40135,N_38654,N_39797);
and U40136 (N_40136,N_38605,N_37735);
or U40137 (N_40137,N_37777,N_38222);
or U40138 (N_40138,N_39843,N_37986);
or U40139 (N_40139,N_37543,N_37702);
nor U40140 (N_40140,N_38557,N_39221);
or U40141 (N_40141,N_38330,N_38400);
and U40142 (N_40142,N_38802,N_38740);
nand U40143 (N_40143,N_39932,N_38969);
xor U40144 (N_40144,N_37616,N_38792);
xnor U40145 (N_40145,N_39203,N_38509);
or U40146 (N_40146,N_38123,N_38894);
xnor U40147 (N_40147,N_38304,N_39211);
nand U40148 (N_40148,N_37939,N_37648);
xor U40149 (N_40149,N_39404,N_39046);
xor U40150 (N_40150,N_38841,N_38235);
xnor U40151 (N_40151,N_39462,N_38915);
or U40152 (N_40152,N_38553,N_38838);
nor U40153 (N_40153,N_37809,N_39387);
and U40154 (N_40154,N_39201,N_37782);
nor U40155 (N_40155,N_39262,N_38923);
nor U40156 (N_40156,N_39841,N_38212);
nor U40157 (N_40157,N_38457,N_37815);
nand U40158 (N_40158,N_37823,N_39180);
nor U40159 (N_40159,N_38808,N_39627);
and U40160 (N_40160,N_37510,N_38960);
or U40161 (N_40161,N_39860,N_39773);
and U40162 (N_40162,N_37566,N_38517);
or U40163 (N_40163,N_38216,N_39130);
and U40164 (N_40164,N_38413,N_39905);
and U40165 (N_40165,N_39899,N_38332);
and U40166 (N_40166,N_39369,N_39737);
xnor U40167 (N_40167,N_38885,N_38603);
xnor U40168 (N_40168,N_37601,N_38804);
and U40169 (N_40169,N_38653,N_38982);
or U40170 (N_40170,N_37987,N_38562);
xnor U40171 (N_40171,N_39084,N_39002);
nand U40172 (N_40172,N_38788,N_39991);
nor U40173 (N_40173,N_37569,N_39204);
xor U40174 (N_40174,N_39090,N_39328);
nand U40175 (N_40175,N_37596,N_39883);
nand U40176 (N_40176,N_38523,N_38429);
xnor U40177 (N_40177,N_38730,N_39663);
xnor U40178 (N_40178,N_39024,N_38350);
nand U40179 (N_40179,N_37608,N_37606);
or U40180 (N_40180,N_39840,N_39464);
nand U40181 (N_40181,N_37804,N_38543);
and U40182 (N_40182,N_38725,N_38856);
and U40183 (N_40183,N_39009,N_39229);
and U40184 (N_40184,N_37567,N_39667);
xor U40185 (N_40185,N_39817,N_37597);
and U40186 (N_40186,N_38626,N_39067);
or U40187 (N_40187,N_38863,N_39903);
and U40188 (N_40188,N_39482,N_38133);
xnor U40189 (N_40189,N_38308,N_39420);
and U40190 (N_40190,N_38002,N_39406);
and U40191 (N_40191,N_39336,N_38009);
nor U40192 (N_40192,N_38270,N_39861);
nor U40193 (N_40193,N_38272,N_37656);
and U40194 (N_40194,N_37867,N_39727);
and U40195 (N_40195,N_38879,N_38257);
xor U40196 (N_40196,N_38476,N_39691);
or U40197 (N_40197,N_37536,N_38076);
nand U40198 (N_40198,N_38860,N_37713);
and U40199 (N_40199,N_39515,N_39392);
xor U40200 (N_40200,N_38130,N_37754);
or U40201 (N_40201,N_39609,N_37966);
or U40202 (N_40202,N_38366,N_38933);
or U40203 (N_40203,N_39974,N_38278);
nor U40204 (N_40204,N_38453,N_38414);
nand U40205 (N_40205,N_38115,N_38970);
nand U40206 (N_40206,N_39141,N_38592);
xor U40207 (N_40207,N_39053,N_39548);
xor U40208 (N_40208,N_39473,N_37741);
and U40209 (N_40209,N_39557,N_39657);
or U40210 (N_40210,N_39760,N_39008);
or U40211 (N_40211,N_38250,N_39955);
xor U40212 (N_40212,N_38358,N_37671);
nor U40213 (N_40213,N_37786,N_38612);
or U40214 (N_40214,N_37858,N_38137);
xor U40215 (N_40215,N_38239,N_39517);
nor U40216 (N_40216,N_38710,N_38062);
and U40217 (N_40217,N_39765,N_38700);
nor U40218 (N_40218,N_39811,N_37590);
nand U40219 (N_40219,N_39256,N_39536);
and U40220 (N_40220,N_39753,N_38515);
xor U40221 (N_40221,N_37512,N_39664);
or U40222 (N_40222,N_38508,N_38786);
nand U40223 (N_40223,N_39845,N_37537);
nand U40224 (N_40224,N_38861,N_38217);
xnor U40225 (N_40225,N_39377,N_38481);
nand U40226 (N_40226,N_38683,N_37801);
nor U40227 (N_40227,N_39671,N_39230);
nand U40228 (N_40228,N_38474,N_38997);
nand U40229 (N_40229,N_39058,N_38716);
nor U40230 (N_40230,N_39720,N_38973);
nand U40231 (N_40231,N_39079,N_39893);
or U40232 (N_40232,N_39214,N_38004);
and U40233 (N_40233,N_38251,N_37645);
nand U40234 (N_40234,N_38576,N_39799);
nand U40235 (N_40235,N_38578,N_39601);
xor U40236 (N_40236,N_38968,N_37505);
and U40237 (N_40237,N_38489,N_38636);
and U40238 (N_40238,N_38518,N_37503);
xnor U40239 (N_40239,N_39091,N_37772);
or U40240 (N_40240,N_39489,N_38706);
nand U40241 (N_40241,N_39836,N_39908);
nand U40242 (N_40242,N_39049,N_38247);
xnor U40243 (N_40243,N_37884,N_38975);
xor U40244 (N_40244,N_39436,N_38116);
nand U40245 (N_40245,N_39380,N_39164);
nand U40246 (N_40246,N_38862,N_39142);
nor U40247 (N_40247,N_39407,N_38305);
or U40248 (N_40248,N_39463,N_38434);
nand U40249 (N_40249,N_38063,N_37506);
or U40250 (N_40250,N_39080,N_37865);
or U40251 (N_40251,N_37773,N_39340);
nand U40252 (N_40252,N_38046,N_39851);
nor U40253 (N_40253,N_39796,N_37984);
nor U40254 (N_40254,N_39351,N_38896);
nand U40255 (N_40255,N_38727,N_38827);
nand U40256 (N_40256,N_39265,N_39076);
and U40257 (N_40257,N_39971,N_39568);
or U40258 (N_40258,N_38539,N_39030);
nor U40259 (N_40259,N_39740,N_38947);
nor U40260 (N_40260,N_39930,N_37903);
nor U40261 (N_40261,N_38850,N_39514);
nand U40262 (N_40262,N_39885,N_38182);
or U40263 (N_40263,N_39754,N_38091);
nor U40264 (N_40264,N_38561,N_39061);
or U40265 (N_40265,N_37841,N_39721);
xnor U40266 (N_40266,N_38547,N_38281);
nor U40267 (N_40267,N_38629,N_38972);
xnor U40268 (N_40268,N_39874,N_37790);
nor U40269 (N_40269,N_37836,N_38864);
nor U40270 (N_40270,N_38849,N_38153);
xnor U40271 (N_40271,N_38671,N_38768);
or U40272 (N_40272,N_39685,N_39358);
or U40273 (N_40273,N_39870,N_39706);
nor U40274 (N_40274,N_38757,N_39645);
nand U40275 (N_40275,N_38844,N_37759);
or U40276 (N_40276,N_37684,N_38624);
nor U40277 (N_40277,N_37827,N_38410);
xor U40278 (N_40278,N_39538,N_39939);
nor U40279 (N_40279,N_37766,N_39389);
nand U40280 (N_40280,N_38949,N_38643);
nor U40281 (N_40281,N_38584,N_37725);
or U40282 (N_40282,N_37821,N_39362);
nand U40283 (N_40283,N_37922,N_38502);
nor U40284 (N_40284,N_39424,N_38313);
xor U40285 (N_40285,N_39842,N_39698);
or U40286 (N_40286,N_37893,N_39776);
or U40287 (N_40287,N_39660,N_37612);
nor U40288 (N_40288,N_37663,N_39367);
or U40289 (N_40289,N_38229,N_39999);
or U40290 (N_40290,N_38172,N_37962);
nand U40291 (N_40291,N_39622,N_39960);
xor U40292 (N_40292,N_39949,N_39537);
nand U40293 (N_40293,N_37864,N_37542);
nor U40294 (N_40294,N_37541,N_39147);
and U40295 (N_40295,N_38296,N_39162);
nand U40296 (N_40296,N_38668,N_39126);
nand U40297 (N_40297,N_38319,N_38220);
or U40298 (N_40298,N_39990,N_38461);
nand U40299 (N_40299,N_39504,N_39054);
and U40300 (N_40300,N_39029,N_38168);
or U40301 (N_40301,N_38241,N_39266);
xnor U40302 (N_40302,N_38857,N_38101);
nor U40303 (N_40303,N_38338,N_39816);
and U40304 (N_40304,N_39086,N_38828);
or U40305 (N_40305,N_39488,N_38451);
or U40306 (N_40306,N_39003,N_39684);
and U40307 (N_40307,N_39102,N_37853);
or U40308 (N_40308,N_39486,N_39154);
nand U40309 (N_40309,N_38407,N_39277);
and U40310 (N_40310,N_38078,N_38430);
xnor U40311 (N_40311,N_38185,N_38139);
nand U40312 (N_40312,N_38805,N_39759);
or U40313 (N_40313,N_38526,N_38349);
xnor U40314 (N_40314,N_39964,N_38356);
or U40315 (N_40315,N_39206,N_39978);
xnor U40316 (N_40316,N_38814,N_38135);
and U40317 (N_40317,N_39881,N_38681);
xor U40318 (N_40318,N_37643,N_39900);
or U40319 (N_40319,N_38174,N_38020);
nand U40320 (N_40320,N_38782,N_37696);
xor U40321 (N_40321,N_37959,N_39532);
and U40322 (N_40322,N_38913,N_39510);
and U40323 (N_40323,N_37999,N_39272);
xor U40324 (N_40324,N_37523,N_39469);
xnor U40325 (N_40325,N_39348,N_38550);
and U40326 (N_40326,N_38256,N_38765);
or U40327 (N_40327,N_37927,N_39607);
and U40328 (N_40328,N_39022,N_39335);
xor U40329 (N_40329,N_38103,N_38482);
nand U40330 (N_40330,N_38218,N_39449);
or U40331 (N_40331,N_39926,N_38618);
and U40332 (N_40332,N_39722,N_39636);
nand U40333 (N_40333,N_37842,N_39421);
nor U40334 (N_40334,N_38563,N_39457);
nand U40335 (N_40335,N_38466,N_39499);
nor U40336 (N_40336,N_39423,N_37658);
or U40337 (N_40337,N_38465,N_38459);
or U40338 (N_40338,N_38086,N_38477);
or U40339 (N_40339,N_38480,N_37699);
xnor U40340 (N_40340,N_39605,N_39716);
xnor U40341 (N_40341,N_39195,N_38484);
nor U40342 (N_40342,N_38494,N_38190);
or U40343 (N_40343,N_39723,N_39835);
nand U40344 (N_40344,N_37904,N_38581);
nor U40345 (N_40345,N_37796,N_37717);
or U40346 (N_40346,N_39063,N_38832);
nor U40347 (N_40347,N_39487,N_37998);
or U40348 (N_40348,N_39808,N_39258);
or U40349 (N_40349,N_39081,N_38162);
xnor U40350 (N_40350,N_39276,N_38816);
nand U40351 (N_40351,N_39872,N_38373);
and U40352 (N_40352,N_39876,N_38385);
nor U40353 (N_40353,N_37923,N_38211);
or U40354 (N_40354,N_39873,N_38927);
or U40355 (N_40355,N_38416,N_37739);
xnor U40356 (N_40356,N_39789,N_38026);
or U40357 (N_40357,N_39139,N_38284);
nor U40358 (N_40358,N_38796,N_38417);
or U40359 (N_40359,N_38470,N_38485);
and U40360 (N_40360,N_37637,N_38945);
or U40361 (N_40361,N_38294,N_39670);
xor U40362 (N_40362,N_38395,N_37588);
xnor U40363 (N_40363,N_38843,N_39687);
xor U40364 (N_40364,N_39922,N_38265);
nand U40365 (N_40365,N_38205,N_39173);
or U40366 (N_40366,N_38452,N_39662);
or U40367 (N_40367,N_38876,N_38917);
and U40368 (N_40368,N_38344,N_37957);
or U40369 (N_40369,N_39734,N_37555);
nor U40370 (N_40370,N_39227,N_38067);
or U40371 (N_40371,N_37955,N_37574);
nor U40372 (N_40372,N_39465,N_38535);
nand U40373 (N_40373,N_38094,N_37716);
nor U40374 (N_40374,N_38300,N_38444);
nor U40375 (N_40375,N_37909,N_39738);
nor U40376 (N_40376,N_39429,N_38893);
xnor U40377 (N_40377,N_37655,N_37581);
or U40378 (N_40378,N_38479,N_39882);
and U40379 (N_40379,N_39787,N_39756);
or U40380 (N_40380,N_38337,N_38743);
xnor U40381 (N_40381,N_39178,N_39616);
and U40382 (N_40382,N_37814,N_38602);
nor U40383 (N_40383,N_38818,N_38993);
nand U40384 (N_40384,N_38819,N_39295);
and U40385 (N_40385,N_39493,N_39792);
xnor U40386 (N_40386,N_39649,N_38995);
xnor U40387 (N_40387,N_39973,N_39937);
or U40388 (N_40388,N_39190,N_39729);
and U40389 (N_40389,N_38833,N_39123);
xor U40390 (N_40390,N_39057,N_37851);
xor U40391 (N_40391,N_38161,N_38571);
and U40392 (N_40392,N_39784,N_39192);
nor U40393 (N_40393,N_38312,N_37641);
xnor U40394 (N_40394,N_39481,N_38336);
and U40395 (N_40395,N_38815,N_38230);
nor U40396 (N_40396,N_39060,N_38213);
or U40397 (N_40397,N_38696,N_38154);
nor U40398 (N_40398,N_38333,N_38449);
and U40399 (N_40399,N_39467,N_39587);
nor U40400 (N_40400,N_39919,N_39599);
nand U40401 (N_40401,N_39128,N_38495);
and U40402 (N_40402,N_38785,N_38544);
xnor U40403 (N_40403,N_39516,N_37852);
or U40404 (N_40404,N_39143,N_38348);
and U40405 (N_40405,N_39925,N_39168);
or U40406 (N_40406,N_38641,N_39950);
and U40407 (N_40407,N_38741,N_37524);
and U40408 (N_40408,N_39642,N_39391);
nand U40409 (N_40409,N_38420,N_37507);
xnor U40410 (N_40410,N_37929,N_37560);
or U40411 (N_40411,N_39144,N_38089);
or U40412 (N_40412,N_39148,N_37873);
or U40413 (N_40413,N_38315,N_38858);
or U40414 (N_40414,N_38891,N_37679);
nor U40415 (N_40415,N_38321,N_38049);
nand U40416 (N_40416,N_38274,N_39875);
nand U40417 (N_40417,N_37647,N_39373);
or U40418 (N_40418,N_38263,N_39381);
or U40419 (N_40419,N_39155,N_38027);
nand U40420 (N_40420,N_39131,N_38351);
or U40421 (N_40421,N_37806,N_39541);
nor U40422 (N_40422,N_39218,N_38191);
nand U40423 (N_40423,N_38327,N_39689);
or U40424 (N_40424,N_37914,N_38524);
nor U40425 (N_40425,N_38082,N_38469);
or U40426 (N_40426,N_37874,N_38156);
nor U40427 (N_40427,N_37611,N_37732);
nand U40428 (N_40428,N_37990,N_37731);
or U40429 (N_40429,N_38432,N_38835);
nor U40430 (N_40430,N_38058,N_39591);
and U40431 (N_40431,N_37745,N_38873);
and U40432 (N_40432,N_37660,N_38692);
or U40433 (N_40433,N_38111,N_37551);
and U40434 (N_40434,N_38215,N_39658);
nor U40435 (N_40435,N_37869,N_39428);
or U40436 (N_40436,N_37794,N_38013);
and U40437 (N_40437,N_37609,N_39246);
nor U40438 (N_40438,N_39880,N_37561);
xor U40439 (N_40439,N_39068,N_38140);
and U40440 (N_40440,N_38519,N_39307);
and U40441 (N_40441,N_38783,N_37859);
xor U40442 (N_40442,N_38219,N_39701);
or U40443 (N_40443,N_38661,N_37582);
and U40444 (N_40444,N_39242,N_39549);
nand U40445 (N_40445,N_39055,N_39826);
and U40446 (N_40446,N_38203,N_37664);
or U40447 (N_40447,N_39709,N_38023);
nor U40448 (N_40448,N_37969,N_38655);
nand U40449 (N_40449,N_37708,N_38677);
xnor U40450 (N_40450,N_38113,N_38572);
nor U40451 (N_40451,N_37714,N_39830);
nand U40452 (N_40452,N_38110,N_39172);
and U40453 (N_40453,N_37863,N_37564);
nor U40454 (N_40454,N_39496,N_39692);
nor U40455 (N_40455,N_38980,N_38488);
and U40456 (N_40456,N_38099,N_37935);
xor U40457 (N_40457,N_37548,N_39824);
or U40458 (N_40458,N_38817,N_38266);
and U40459 (N_40459,N_38492,N_39451);
nor U40460 (N_40460,N_38918,N_39837);
nor U40461 (N_40461,N_39672,N_38634);
and U40462 (N_40462,N_39495,N_39606);
nand U40463 (N_40463,N_39244,N_39213);
nand U40464 (N_40464,N_38875,N_38468);
or U40465 (N_40465,N_39048,N_39619);
and U40466 (N_40466,N_37644,N_39232);
and U40467 (N_40467,N_39602,N_38383);
xor U40468 (N_40468,N_39426,N_38254);
xor U40469 (N_40469,N_38529,N_38109);
and U40470 (N_40470,N_39507,N_37653);
nor U40471 (N_40471,N_39928,N_39547);
nand U40472 (N_40472,N_39525,N_38905);
or U40473 (N_40473,N_38921,N_39864);
nor U40474 (N_40474,N_39791,N_38043);
or U40475 (N_40475,N_39566,N_38575);
and U40476 (N_40476,N_37520,N_38379);
or U40477 (N_40477,N_37813,N_38503);
and U40478 (N_40478,N_39231,N_38999);
or U40479 (N_40479,N_39944,N_38702);
xor U40480 (N_40480,N_38121,N_37701);
nor U40481 (N_40481,N_38225,N_39795);
or U40482 (N_40482,N_39359,N_37876);
or U40483 (N_40483,N_38690,N_39207);
nor U40484 (N_40484,N_37940,N_39124);
xor U40485 (N_40485,N_39593,N_38522);
nand U40486 (N_40486,N_37820,N_38180);
and U40487 (N_40487,N_39934,N_39092);
and U40488 (N_40488,N_38958,N_38255);
or U40489 (N_40489,N_37958,N_39564);
and U40490 (N_40490,N_39777,N_38345);
and U40491 (N_40491,N_38398,N_38695);
nand U40492 (N_40492,N_38542,N_39176);
nand U40493 (N_40493,N_38651,N_38051);
nand U40494 (N_40494,N_37710,N_39803);
nor U40495 (N_40495,N_39477,N_39600);
nand U40496 (N_40496,N_38648,N_38514);
nor U40497 (N_40497,N_37952,N_39025);
xnor U40498 (N_40498,N_39646,N_37585);
nor U40499 (N_40499,N_38098,N_39577);
nor U40500 (N_40500,N_39183,N_39217);
nand U40501 (N_40501,N_39767,N_38650);
or U40502 (N_40502,N_38824,N_39977);
nand U40503 (N_40503,N_38983,N_39134);
nor U40504 (N_40504,N_39405,N_39438);
nand U40505 (N_40505,N_39783,N_39108);
or U40506 (N_40506,N_38412,N_39019);
xnor U40507 (N_40507,N_39316,N_38742);
nand U40508 (N_40508,N_39623,N_38018);
xnor U40509 (N_40509,N_38186,N_38516);
nor U40510 (N_40510,N_39942,N_37627);
nor U40511 (N_40511,N_39800,N_38194);
nand U40512 (N_40512,N_39430,N_37534);
nor U40513 (N_40513,N_39376,N_38834);
or U40514 (N_40514,N_38386,N_38246);
and U40515 (N_40515,N_38008,N_38682);
nor U40516 (N_40516,N_39078,N_39979);
and U40517 (N_40517,N_39313,N_39981);
nor U40518 (N_40518,N_39719,N_37634);
nand U40519 (N_40519,N_37584,N_37746);
or U40520 (N_40520,N_39745,N_39169);
nand U40521 (N_40521,N_39630,N_39396);
nand U40522 (N_40522,N_39574,N_39610);
and U40523 (N_40523,N_38527,N_37681);
and U40524 (N_40524,N_38633,N_38736);
or U40525 (N_40525,N_39572,N_39158);
and U40526 (N_40526,N_38604,N_39419);
or U40527 (N_40527,N_38289,N_38310);
nor U40528 (N_40528,N_38152,N_38165);
nor U40529 (N_40529,N_39781,N_38475);
xnor U40530 (N_40530,N_37765,N_37600);
nand U40531 (N_40531,N_38619,N_39197);
xnor U40532 (N_40532,N_37924,N_39933);
nor U40533 (N_40533,N_38507,N_37756);
and U40534 (N_40534,N_39699,N_39674);
or U40535 (N_40535,N_37850,N_38189);
or U40536 (N_40536,N_38314,N_37638);
nand U40537 (N_40537,N_39250,N_38902);
and U40538 (N_40538,N_37818,N_38423);
nand U40539 (N_40539,N_37798,N_37830);
xnor U40540 (N_40540,N_39374,N_38025);
and U40541 (N_40541,N_38253,N_38946);
and U40542 (N_40542,N_38877,N_38401);
xor U40543 (N_40543,N_38937,N_39554);
and U40544 (N_40544,N_37921,N_39603);
nand U40545 (N_40545,N_39205,N_38317);
xnor U40546 (N_40546,N_39484,N_39371);
nor U40547 (N_40547,N_38580,N_39655);
xnor U40548 (N_40548,N_39403,N_39614);
or U40549 (N_40549,N_39539,N_39820);
xor U40550 (N_40550,N_37916,N_39902);
nor U40551 (N_40551,N_37562,N_38570);
and U40552 (N_40552,N_38262,N_39333);
or U40553 (N_40553,N_39196,N_38033);
or U40554 (N_40554,N_38698,N_39077);
nand U40555 (N_40555,N_37605,N_37763);
nor U40556 (N_40556,N_39453,N_38678);
nor U40557 (N_40557,N_38617,N_39807);
nor U40558 (N_40558,N_39597,N_38822);
or U40559 (N_40559,N_38701,N_38405);
xor U40560 (N_40560,N_39770,N_38721);
nand U40561 (N_40561,N_38541,N_39513);
nor U40562 (N_40562,N_39032,N_39361);
nand U40563 (N_40563,N_39819,N_38703);
nand U40564 (N_40564,N_39443,N_37963);
or U40565 (N_40565,N_38599,N_38493);
xnor U40566 (N_40566,N_39356,N_37508);
or U40567 (N_40567,N_38647,N_38201);
or U40568 (N_40568,N_37769,N_38615);
and U40569 (N_40569,N_37953,N_39561);
nand U40570 (N_40570,N_38331,N_37913);
and U40571 (N_40571,N_39818,N_38059);
nor U40572 (N_40572,N_37885,N_39113);
and U40573 (N_40573,N_38799,N_38170);
nor U40574 (N_40574,N_38329,N_38127);
or U40575 (N_40575,N_37624,N_39596);
or U40576 (N_40576,N_39310,N_39637);
xnor U40577 (N_40577,N_37672,N_38748);
nand U40578 (N_40578,N_37517,N_39744);
or U40579 (N_40579,N_39290,N_39878);
nor U40580 (N_40580,N_37971,N_38689);
nor U40581 (N_40581,N_39257,N_38595);
or U40582 (N_40582,N_38558,N_37889);
and U40583 (N_40583,N_38724,N_39898);
nor U40584 (N_40584,N_39326,N_37925);
nand U40585 (N_40585,N_39312,N_39794);
nand U40586 (N_40586,N_39268,N_39530);
nor U40587 (N_40587,N_38813,N_39341);
and U40588 (N_40588,N_39209,N_37824);
xor U40589 (N_40589,N_38922,N_37797);
or U40590 (N_40590,N_39661,N_38138);
or U40591 (N_40591,N_37683,N_38644);
nand U40592 (N_40592,N_39065,N_39520);
nor U40593 (N_40593,N_37516,N_37857);
or U40594 (N_40594,N_39112,N_39501);
xnor U40595 (N_40595,N_39039,N_39895);
and U40596 (N_40596,N_37689,N_37712);
nor U40597 (N_40597,N_39518,N_39459);
nand U40598 (N_40598,N_38145,N_38623);
nand U40599 (N_40599,N_37808,N_39641);
and U40600 (N_40600,N_38209,N_37881);
xor U40601 (N_40601,N_37636,N_39439);
or U40602 (N_40602,N_39761,N_38437);
xor U40603 (N_40603,N_38895,N_39357);
xor U40604 (N_40604,N_39305,N_39527);
nand U40605 (N_40605,N_39286,N_38754);
nand U40606 (N_40606,N_38900,N_39115);
xnor U40607 (N_40607,N_38149,N_39393);
xnor U40608 (N_40608,N_39941,N_37632);
xnor U40609 (N_40609,N_38061,N_38717);
or U40610 (N_40610,N_38538,N_39251);
or U40611 (N_40611,N_37583,N_37615);
and U40612 (N_40612,N_38583,N_39301);
nor U40613 (N_40613,N_39543,N_39553);
nand U40614 (N_40614,N_38340,N_39352);
nand U40615 (N_40615,N_39047,N_38951);
nand U40616 (N_40616,N_39347,N_38954);
and U40617 (N_40617,N_37908,N_39167);
nor U40618 (N_40618,N_39702,N_38378);
xor U40619 (N_40619,N_39531,N_39275);
nor U40620 (N_40620,N_38820,N_38546);
or U40621 (N_40621,N_39349,N_38326);
xor U40622 (N_40622,N_39474,N_39631);
nand U40623 (N_40623,N_37723,N_39544);
nand U40624 (N_40624,N_38045,N_39976);
or U40625 (N_40625,N_39748,N_37890);
xor U40626 (N_40626,N_38590,N_39093);
nand U40627 (N_40627,N_38299,N_39897);
xnor U40628 (N_40628,N_38347,N_39021);
xnor U40629 (N_40629,N_38930,N_38693);
nor U40630 (N_40630,N_38372,N_39435);
xnor U40631 (N_40631,N_38088,N_38658);
nor U40632 (N_40632,N_39613,N_37928);
and U40633 (N_40633,N_37651,N_39573);
and U40634 (N_40634,N_38195,N_38674);
xnor U40635 (N_40635,N_37744,N_38448);
nand U40636 (N_40636,N_39468,N_37686);
nor U40637 (N_40637,N_39085,N_39559);
nor U40638 (N_40638,N_39712,N_39300);
nor U40639 (N_40639,N_38766,N_38840);
nand U40640 (N_40640,N_39681,N_38243);
or U40641 (N_40641,N_38167,N_39177);
and U40642 (N_40642,N_39422,N_37918);
nand U40643 (N_40643,N_39628,N_38460);
nand U40644 (N_40644,N_39099,N_39120);
or U40645 (N_40645,N_39498,N_38780);
and U40646 (N_40646,N_37610,N_38368);
or U40647 (N_40647,N_38992,N_38286);
and U40648 (N_40648,N_39534,N_38097);
nor U40649 (N_40649,N_39743,N_38837);
and U40650 (N_40650,N_38582,N_39492);
and U40651 (N_40651,N_38772,N_37981);
nand U40652 (N_40652,N_38746,N_37527);
or U40653 (N_40653,N_39589,N_38732);
xnor U40654 (N_40654,N_38851,N_39782);
xnor U40655 (N_40655,N_37896,N_38322);
or U40656 (N_40656,N_39145,N_38419);
nand U40657 (N_40657,N_39624,N_39774);
nor U40658 (N_40658,N_39062,N_38390);
nand U40659 (N_40659,N_39988,N_37572);
and U40660 (N_40660,N_37740,N_39894);
and U40661 (N_40661,N_37525,N_38342);
xnor U40662 (N_40662,N_38791,N_39253);
nor U40663 (N_40663,N_38979,N_39718);
nor U40664 (N_40664,N_39210,N_38549);
nor U40665 (N_40665,N_39045,N_38868);
and U40666 (N_40666,N_37694,N_38311);
nand U40667 (N_40667,N_38649,N_39786);
nor U40668 (N_40668,N_39746,N_37855);
nor U40669 (N_40669,N_38136,N_38260);
xnor U40670 (N_40670,N_38961,N_39005);
nor U40671 (N_40671,N_38030,N_39936);
nand U40672 (N_40672,N_38707,N_39117);
and U40673 (N_40673,N_39271,N_37670);
xor U40674 (N_40674,N_38285,N_39094);
xor U40675 (N_40675,N_38715,N_37743);
and U40676 (N_40676,N_39226,N_38709);
xor U40677 (N_40677,N_37598,N_39682);
nand U40678 (N_40678,N_38069,N_37533);
nand U40679 (N_40679,N_38723,N_38499);
xnor U40680 (N_40680,N_39331,N_39334);
and U40681 (N_40681,N_39136,N_39318);
nor U40682 (N_40682,N_38940,N_37956);
and U40683 (N_40683,N_39188,N_38609);
and U40684 (N_40684,N_39983,N_37552);
nand U40685 (N_40685,N_38962,N_39004);
and U40686 (N_40686,N_38751,N_39871);
nand U40687 (N_40687,N_37729,N_37880);
and U40688 (N_40688,N_39325,N_38984);
xnor U40689 (N_40689,N_38865,N_39779);
nor U40690 (N_40690,N_39306,N_37675);
nand U40691 (N_40691,N_38797,N_39626);
and U40692 (N_40692,N_38403,N_38888);
and U40693 (N_40693,N_39923,N_37785);
and U40694 (N_40694,N_39111,N_39909);
xor U40695 (N_40695,N_37901,N_38108);
xnor U40696 (N_40696,N_37948,N_37539);
and U40697 (N_40697,N_39409,N_38621);
or U40698 (N_40698,N_39417,N_38100);
or U40699 (N_40699,N_39965,N_38996);
xor U40700 (N_40700,N_39446,N_39653);
or U40701 (N_40701,N_37768,N_39412);
xor U40702 (N_40702,N_38394,N_37900);
and U40703 (N_40703,N_39920,N_37915);
nor U40704 (N_40704,N_38129,N_37538);
nand U40705 (N_40705,N_39831,N_39216);
and U40706 (N_40706,N_38374,N_39832);
nor U40707 (N_40707,N_38126,N_37795);
nor U40708 (N_40708,N_39683,N_37778);
and U40709 (N_40709,N_39854,N_38775);
nand U40710 (N_40710,N_38622,N_38699);
or U40711 (N_40711,N_37949,N_38790);
nand U40712 (N_40712,N_38048,N_38224);
nor U40713 (N_40713,N_38392,N_39153);
nor U40714 (N_40714,N_37767,N_39279);
nor U40715 (N_40715,N_37974,N_39043);
or U40716 (N_40716,N_39324,N_39040);
and U40717 (N_40717,N_38639,N_37898);
xnor U40718 (N_40718,N_37528,N_39219);
xor U40719 (N_40719,N_38483,N_39927);
nand U40720 (N_40720,N_38907,N_38774);
or U40721 (N_40721,N_38259,N_37707);
or U40722 (N_40722,N_37781,N_38238);
xnor U40723 (N_40723,N_37722,N_39924);
xnor U40724 (N_40724,N_38268,N_38845);
nand U40725 (N_40725,N_39337,N_39717);
and U40726 (N_40726,N_39296,N_38258);
or U40727 (N_40727,N_38144,N_37691);
xnor U40728 (N_40728,N_37737,N_38060);
or U40729 (N_40729,N_37882,N_37595);
nand U40730 (N_40730,N_38192,N_38335);
or U40731 (N_40731,N_38686,N_38520);
nand U40732 (N_40732,N_39254,N_38778);
nand U40733 (N_40733,N_38914,N_39220);
xor U40734 (N_40734,N_38231,N_37819);
nand U40735 (N_40735,N_38665,N_39273);
or U40736 (N_40736,N_39129,N_39282);
nor U40737 (N_40737,N_39654,N_37860);
nand U40738 (N_40738,N_38755,N_39580);
nor U40739 (N_40739,N_38662,N_38931);
nor U40740 (N_40740,N_38713,N_37592);
or U40741 (N_40741,N_38223,N_38635);
and U40742 (N_40742,N_39680,N_39710);
nand U40743 (N_40743,N_38953,N_38988);
xor U40744 (N_40744,N_39506,N_39567);
nand U40745 (N_40745,N_38631,N_38150);
nor U40746 (N_40746,N_38316,N_38598);
and U40747 (N_40747,N_39766,N_38745);
xor U40748 (N_40748,N_37758,N_37943);
nand U40749 (N_40749,N_39327,N_39522);
nand U40750 (N_40750,N_38183,N_38179);
and U40751 (N_40751,N_38564,N_39644);
nor U40752 (N_40752,N_39011,N_37843);
or U40753 (N_40753,N_38017,N_38532);
and U40754 (N_40754,N_38901,N_39911);
and U40755 (N_40755,N_38718,N_39311);
nand U40756 (N_40756,N_39485,N_39914);
nor U40757 (N_40757,N_38122,N_39980);
and U40758 (N_40758,N_38638,N_38759);
nand U40759 (N_40759,N_38957,N_38869);
nand U40760 (N_40760,N_38540,N_38944);
and U40761 (N_40761,N_39752,N_39259);
and U40762 (N_40762,N_38769,N_39827);
nand U40763 (N_40763,N_38705,N_37835);
or U40764 (N_40764,N_38324,N_39191);
or U40765 (N_40765,N_39958,N_38898);
xnor U40766 (N_40766,N_39110,N_39956);
xnor U40767 (N_40767,N_38903,N_38200);
or U40768 (N_40768,N_38019,N_39998);
xor U40769 (N_40769,N_38068,N_39497);
nor U40770 (N_40770,N_38292,N_39838);
xnor U40771 (N_40771,N_38513,N_37871);
nand U40772 (N_40772,N_39500,N_39617);
or U40773 (N_40773,N_39303,N_38029);
or U40774 (N_40774,N_38440,N_39901);
and U40775 (N_40775,N_39550,N_39483);
nor U40776 (N_40776,N_39088,N_39997);
and U40777 (N_40777,N_38645,N_39673);
and U40778 (N_40778,N_38853,N_39724);
or U40779 (N_40779,N_39400,N_38704);
and U40780 (N_40780,N_39966,N_38066);
and U40781 (N_40781,N_38981,N_39137);
xnor U40782 (N_40782,N_37931,N_39569);
or U40783 (N_40783,N_39732,N_39528);
nor U40784 (N_40784,N_38036,N_37895);
and U40785 (N_40785,N_39452,N_38756);
and U40786 (N_40786,N_39414,N_37888);
nand U40787 (N_40787,N_37705,N_39780);
nor U40788 (N_40788,N_39906,N_39471);
and U40789 (N_40789,N_39879,N_38007);
xor U40790 (N_40790,N_39103,N_38731);
nand U40791 (N_40791,N_37747,N_38226);
and U40792 (N_40792,N_39865,N_39052);
nor U40793 (N_40793,N_38204,N_38387);
nand U40794 (N_40794,N_37668,N_37614);
or U40795 (N_40795,N_39442,N_38767);
nor U40796 (N_40796,N_37695,N_39478);
nand U40797 (N_40797,N_38925,N_39695);
xor U40798 (N_40798,N_38166,N_39801);
nor U40799 (N_40799,N_38684,N_39199);
and U40800 (N_40800,N_39343,N_39852);
xnor U40801 (N_40801,N_38039,N_38443);
xor U40802 (N_40802,N_37665,N_38628);
nand U40803 (N_40803,N_38169,N_37776);
xor U40804 (N_40804,N_38357,N_39384);
or U40805 (N_40805,N_39161,N_39535);
or U40806 (N_40806,N_37718,N_39490);
or U40807 (N_40807,N_37894,N_39954);
nor U40808 (N_40808,N_38600,N_39089);
xnor U40809 (N_40809,N_39665,N_38376);
xnor U40810 (N_40810,N_39104,N_37965);
or U40811 (N_40811,N_39031,N_37604);
or U40812 (N_40812,N_38986,N_37531);
xor U40813 (N_40813,N_37591,N_39171);
xnor U40814 (N_40814,N_38714,N_39269);
nand U40815 (N_40815,N_38846,N_39935);
nand U40816 (N_40816,N_37832,N_38501);
nand U40817 (N_40817,N_39558,N_37557);
and U40818 (N_40818,N_37907,N_38445);
and U40819 (N_40819,N_38825,N_39292);
xor U40820 (N_40820,N_38455,N_39586);
nor U40821 (N_40821,N_38052,N_38601);
or U40822 (N_40822,N_39035,N_39302);
or U40823 (N_40823,N_39297,N_37787);
or U40824 (N_40824,N_39000,N_39291);
and U40825 (N_40825,N_38016,N_38672);
xor U40826 (N_40826,N_39458,N_39968);
nor U40827 (N_40827,N_37511,N_39368);
nand U40828 (N_40828,N_37626,N_37937);
nand U40829 (N_40829,N_37912,N_39447);
nor U40830 (N_40830,N_39208,N_39757);
or U40831 (N_40831,N_39338,N_38072);
xnor U40832 (N_40832,N_37736,N_38566);
or U40833 (N_40833,N_38276,N_37872);
nand U40834 (N_40834,N_37793,N_37594);
or U40835 (N_40835,N_38722,N_38143);
or U40836 (N_40836,N_38597,N_39007);
xor U40837 (N_40837,N_39884,N_38196);
nand U40838 (N_40838,N_39688,N_37628);
or U40839 (N_40839,N_38221,N_38454);
xnor U40840 (N_40840,N_39122,N_37810);
xor U40841 (N_40841,N_37727,N_39651);
or U40842 (N_40842,N_39239,N_39633);
and U40843 (N_40843,N_38531,N_38354);
xnor U40844 (N_40844,N_39711,N_39156);
nand U40845 (N_40845,N_38290,N_39850);
xnor U40846 (N_40846,N_39267,N_39769);
or U40847 (N_40847,N_37690,N_38498);
xnor U40848 (N_40848,N_38750,N_39853);
or U40849 (N_40849,N_39540,N_39087);
nor U40850 (N_40850,N_39730,N_38396);
nand U40851 (N_40851,N_37803,N_38559);
xnor U40852 (N_40852,N_37532,N_39027);
nor U40853 (N_40853,N_39491,N_39411);
and U40854 (N_40854,N_39119,N_39788);
xnor U40855 (N_40855,N_38159,N_39555);
nor U40856 (N_40856,N_38382,N_39815);
or U40857 (N_40857,N_37646,N_37932);
and U40858 (N_40858,N_39072,N_38966);
nor U40859 (N_40859,N_38408,N_38685);
and U40860 (N_40860,N_38967,N_38273);
or U40861 (N_40861,N_37917,N_39116);
or U40862 (N_40862,N_39082,N_39829);
nand U40863 (N_40863,N_38393,N_39166);
nor U40864 (N_40864,N_39163,N_38433);
or U40865 (N_40865,N_37829,N_38776);
or U40866 (N_40866,N_39372,N_39581);
or U40867 (N_40867,N_38491,N_39867);
xnor U40868 (N_40868,N_38021,N_39620);
xor U40869 (N_40869,N_39408,N_39460);
or U40870 (N_40870,N_39194,N_39763);
and U40871 (N_40871,N_39666,N_37685);
nor U40872 (N_40872,N_38237,N_37526);
and U40873 (N_40873,N_37509,N_39886);
nor U40874 (N_40874,N_38442,N_39441);
xnor U40875 (N_40875,N_39159,N_37791);
and U40876 (N_40876,N_37942,N_38264);
nand U40877 (N_40877,N_38184,N_38462);
nand U40878 (N_40878,N_38198,N_37822);
and U40879 (N_40879,N_39545,N_37968);
nand U40880 (N_40880,N_37639,N_38472);
or U40881 (N_40881,N_37812,N_39749);
nand U40882 (N_40882,N_39669,N_37540);
xor U40883 (N_40883,N_37784,N_37792);
or U40884 (N_40884,N_39931,N_38812);
and U40885 (N_40885,N_39529,N_39805);
nand U40886 (N_40886,N_38801,N_38512);
nor U40887 (N_40887,N_39010,N_37817);
nand U40888 (N_40888,N_39533,N_39963);
xnor U40889 (N_40889,N_38771,N_38998);
or U40890 (N_40890,N_38282,N_38676);
xor U40891 (N_40891,N_39050,N_39813);
nand U40892 (N_40892,N_38411,N_39806);
nand U40893 (N_40893,N_39678,N_38852);
or U40894 (N_40894,N_38269,N_37607);
nor U40895 (N_40895,N_38346,N_39703);
xor U40896 (N_40896,N_38343,N_37964);
or U40897 (N_40897,N_39319,N_38096);
nand U40898 (N_40898,N_38056,N_39378);
xnor U40899 (N_40899,N_39993,N_37662);
nand U40900 (N_40900,N_38839,N_39382);
xnor U40901 (N_40901,N_38131,N_38015);
or U40902 (N_40902,N_39364,N_39961);
nand U40903 (N_40903,N_38831,N_39385);
xnor U40904 (N_40904,N_39402,N_37559);
and U40905 (N_40905,N_37706,N_38652);
and U40906 (N_40906,N_37733,N_39012);
or U40907 (N_40907,N_37748,N_38252);
nor U40908 (N_40908,N_38965,N_38160);
or U40909 (N_40909,N_37535,N_39243);
or U40910 (N_40910,N_37734,N_37831);
nor U40911 (N_40911,N_38320,N_38630);
or U40912 (N_40912,N_37779,N_39224);
xor U40913 (N_40913,N_38607,N_39989);
nor U40914 (N_40914,N_37579,N_37667);
nand U40915 (N_40915,N_38613,N_37875);
nand U40916 (N_40916,N_37613,N_39140);
or U40917 (N_40917,N_38886,N_37522);
or U40918 (N_40918,N_38823,N_37652);
nor U40919 (N_40919,N_39193,N_38625);
and U40920 (N_40920,N_38926,N_38104);
xor U40921 (N_40921,N_39888,N_39461);
nand U40922 (N_40922,N_38409,N_38614);
nor U40923 (N_40923,N_38147,N_38871);
or U40924 (N_40924,N_37514,N_39006);
xor U40925 (N_40925,N_37847,N_39921);
xor U40926 (N_40926,N_37635,N_38795);
nand U40927 (N_40927,N_37845,N_38438);
xor U40928 (N_40928,N_38233,N_38803);
xnor U40929 (N_40929,N_37619,N_39314);
and U40930 (N_40930,N_38548,N_39798);
xnor U40931 (N_40931,N_39016,N_38044);
or U40932 (N_40932,N_39001,N_38085);
xor U40933 (N_40933,N_37500,N_38249);
xor U40934 (N_40934,N_38806,N_39098);
or U40935 (N_40935,N_39315,N_37550);
xnor U40936 (N_40936,N_39233,N_39383);
nor U40937 (N_40937,N_38275,N_39101);
xnor U40938 (N_40938,N_38298,N_37544);
or U40939 (N_40939,N_37868,N_39855);
nor U40940 (N_40940,N_38588,N_37659);
nor U40941 (N_40941,N_38989,N_37565);
nor U40942 (N_40942,N_37807,N_38388);
nand U40943 (N_40943,N_39648,N_38279);
nand U40944 (N_40944,N_39479,N_38283);
nand U40945 (N_40945,N_39953,N_38074);
or U40946 (N_40946,N_38424,N_39245);
or U40947 (N_40947,N_38307,N_39833);
nand U40948 (N_40948,N_37631,N_38355);
xnor U40949 (N_40949,N_39329,N_38729);
or U40950 (N_40950,N_39844,N_39552);
xnor U40951 (N_40951,N_37755,N_37719);
or U40952 (N_40952,N_38753,N_39410);
or U40953 (N_40953,N_38821,N_38536);
nand U40954 (N_40954,N_39431,N_38486);
xnor U40955 (N_40955,N_39707,N_38720);
xor U40956 (N_40956,N_38573,N_38589);
nand U40957 (N_40957,N_37834,N_37504);
or U40958 (N_40958,N_37897,N_39676);
xnor U40959 (N_40959,N_38328,N_38377);
xor U40960 (N_40960,N_39360,N_39059);
and U40961 (N_40961,N_37687,N_38859);
and U40962 (N_40962,N_38341,N_39524);
nand U40963 (N_40963,N_38034,N_39225);
xnor U40964 (N_40964,N_38471,N_38132);
nand U40965 (N_40965,N_38726,N_38496);
nor U40966 (N_40966,N_38240,N_37674);
nor U40967 (N_40967,N_38525,N_39375);
nor U40968 (N_40968,N_38001,N_37558);
xnor U40969 (N_40969,N_39809,N_38565);
nand U40970 (N_40970,N_37899,N_39594);
and U40971 (N_40971,N_39321,N_37996);
nand U40972 (N_40972,N_38093,N_38490);
or U40973 (N_40973,N_39868,N_39604);
and U40974 (N_40974,N_39353,N_37980);
and U40975 (N_40975,N_38303,N_39394);
and U40976 (N_40976,N_38585,N_38406);
xor U40977 (N_40977,N_38000,N_38593);
xor U40978 (N_40978,N_39157,N_39249);
nand U40979 (N_40979,N_39891,N_37568);
and U40980 (N_40980,N_39187,N_39621);
xnor U40981 (N_40981,N_38175,N_38381);
and U40982 (N_40982,N_38242,N_37753);
xnor U40983 (N_40983,N_39308,N_38010);
nand U40984 (N_40984,N_39959,N_39202);
or U40985 (N_40985,N_38943,N_37553);
and U40986 (N_40986,N_39615,N_38606);
xnor U40987 (N_40987,N_39679,N_38556);
xnor U40988 (N_40988,N_38974,N_39957);
xor U40989 (N_40989,N_38084,N_38809);
nand U40990 (N_40990,N_38675,N_38712);
nor U40991 (N_40991,N_38053,N_38365);
nand U40992 (N_40992,N_39938,N_39762);
nor U40993 (N_40993,N_37556,N_38095);
xor U40994 (N_40994,N_38214,N_39152);
or U40995 (N_40995,N_38426,N_38899);
nor U40996 (N_40996,N_38397,N_39521);
and U40997 (N_40997,N_39848,N_39863);
and U40998 (N_40998,N_38236,N_38881);
or U40999 (N_40999,N_39611,N_38171);
xnor U41000 (N_41000,N_38554,N_39565);
and U41001 (N_41001,N_37789,N_38187);
nand U41002 (N_41002,N_38938,N_39556);
or U41003 (N_41003,N_38510,N_39857);
nand U41004 (N_41004,N_39668,N_38087);
and U41005 (N_41005,N_38620,N_38370);
nor U41006 (N_41006,N_38037,N_39480);
xor U41007 (N_41007,N_39138,N_39342);
or U41008 (N_41008,N_39994,N_39363);
nor U41009 (N_41009,N_39322,N_39415);
nor U41010 (N_41010,N_38118,N_38679);
nor U41011 (N_41011,N_37563,N_37738);
nor U41012 (N_41012,N_37870,N_37961);
xor U41013 (N_41013,N_38777,N_39281);
nand U41014 (N_41014,N_38784,N_37720);
nand U41015 (N_41015,N_39612,N_39992);
nor U41016 (N_41016,N_38005,N_38912);
nand U41017 (N_41017,N_39892,N_38528);
xor U41018 (N_41018,N_38193,N_38874);
or U41019 (N_41019,N_39690,N_38146);
nand U41020 (N_41020,N_38789,N_39427);
nand U41021 (N_41021,N_38402,N_38361);
nor U41022 (N_41022,N_39425,N_39355);
or U41023 (N_41023,N_39751,N_38734);
or U41024 (N_41024,N_39456,N_38627);
and U41025 (N_41025,N_39033,N_39165);
nor U41026 (N_41026,N_39948,N_39179);
xnor U41027 (N_41027,N_39869,N_37657);
or U41028 (N_41028,N_39260,N_39476);
nand U41029 (N_41029,N_39028,N_38855);
or U41030 (N_41030,N_38810,N_38206);
nor U41031 (N_41031,N_37654,N_38569);
and U41032 (N_41032,N_37947,N_38826);
nor U41033 (N_41033,N_37861,N_39434);
or U41034 (N_41034,N_38181,N_39940);
or U41035 (N_41035,N_38752,N_38919);
or U41036 (N_41036,N_38064,N_38610);
xnor U41037 (N_41037,N_38904,N_38261);
nor U41038 (N_41038,N_37944,N_38939);
nor U41039 (N_41039,N_39638,N_39241);
nand U41040 (N_41040,N_39731,N_38141);
nand U41041 (N_41041,N_38728,N_39705);
nand U41042 (N_41042,N_38128,N_38511);
nor U41043 (N_41043,N_38574,N_38446);
and U41044 (N_41044,N_38761,N_39293);
or U41045 (N_41045,N_39264,N_38616);
nand U41046 (N_41046,N_37692,N_38352);
and U41047 (N_41047,N_39810,N_39470);
or U41048 (N_41048,N_39945,N_38521);
and U41049 (N_41049,N_38042,N_38012);
xnor U41050 (N_41050,N_38425,N_39625);
xnor U41051 (N_41051,N_38107,N_39972);
and U41052 (N_41052,N_38456,N_38031);
nand U41053 (N_41053,N_37977,N_37905);
nor U41054 (N_41054,N_38458,N_38050);
or U41055 (N_41055,N_39659,N_38872);
nand U41056 (N_41056,N_39284,N_38057);
xnor U41057 (N_41057,N_37848,N_38163);
nand U41058 (N_41058,N_38924,N_38847);
and U41059 (N_41059,N_38267,N_39133);
or U41060 (N_41060,N_38450,N_38985);
nand U41061 (N_41061,N_37877,N_39198);
xnor U41062 (N_41062,N_39704,N_38028);
xor U41063 (N_41063,N_37678,N_39739);
nand U41064 (N_41064,N_37649,N_39235);
nand U41065 (N_41065,N_38842,N_38297);
nor U41066 (N_41066,N_39234,N_39288);
or U41067 (N_41067,N_37623,N_39778);
nand U41068 (N_41068,N_38176,N_38418);
and U41069 (N_41069,N_38829,N_39215);
xor U41070 (N_41070,N_39365,N_38657);
and U41071 (N_41071,N_39910,N_39270);
and U41072 (N_41072,N_39228,N_38533);
nand U41073 (N_41073,N_39725,N_38591);
nor U41074 (N_41074,N_39320,N_38552);
or U41075 (N_41075,N_38632,N_39454);
nor U41076 (N_41076,N_39887,N_37995);
nand U41077 (N_41077,N_39236,N_38920);
nand U41078 (N_41078,N_39656,N_38793);
and U41079 (N_41079,N_38363,N_38807);
and U41080 (N_41080,N_39317,N_38935);
and U41081 (N_41081,N_39505,N_37650);
xnor U41082 (N_41082,N_39708,N_38035);
xor U41083 (N_41083,N_38177,N_39416);
or U41084 (N_41084,N_39755,N_38878);
nor U41085 (N_41085,N_37673,N_37910);
nand U41086 (N_41086,N_37991,N_37982);
or U41087 (N_41087,N_37802,N_37693);
or U41088 (N_41088,N_38830,N_39299);
or U41089 (N_41089,N_38747,N_37680);
and U41090 (N_41090,N_39023,N_38228);
or U41091 (N_41091,N_39812,N_39639);
and U41092 (N_41092,N_37839,N_38941);
and U41093 (N_41093,N_39694,N_39618);
nor U41094 (N_41094,N_38735,N_39775);
nor U41095 (N_41095,N_39181,N_39570);
xor U41096 (N_41096,N_39109,N_39105);
nand U41097 (N_41097,N_39503,N_39287);
nand U41098 (N_41098,N_39904,N_37886);
and U41099 (N_41099,N_38555,N_39523);
or U41100 (N_41100,N_39696,N_39823);
and U41101 (N_41101,N_38119,N_39118);
nor U41102 (N_41102,N_39066,N_37750);
nor U41103 (N_41103,N_39502,N_38773);
and U41104 (N_41104,N_38142,N_39726);
nor U41105 (N_41105,N_37954,N_39034);
nor U41106 (N_41106,N_39943,N_37501);
or U41107 (N_41107,N_38567,N_38660);
or U41108 (N_41108,N_39069,N_39822);
nand U41109 (N_41109,N_39455,N_38500);
or U41110 (N_41110,N_38880,N_37642);
nor U41111 (N_41111,N_38568,N_38848);
or U41112 (N_41112,N_38047,N_37640);
nand U41113 (N_41113,N_38977,N_38794);
xnor U41114 (N_41114,N_39598,N_38202);
xnor U41115 (N_41115,N_38551,N_37967);
or U41116 (N_41116,N_38197,N_39714);
nor U41117 (N_41117,N_37618,N_39986);
and U41118 (N_41118,N_39445,N_38022);
nor U41119 (N_41119,N_39095,N_39175);
nand U41120 (N_41120,N_39071,N_39713);
and U41121 (N_41121,N_38749,N_37950);
nor U41122 (N_41122,N_38054,N_37573);
nor U41123 (N_41123,N_37992,N_37760);
and U41124 (N_41124,N_39390,N_38560);
nand U41125 (N_41125,N_39051,N_38293);
and U41126 (N_41126,N_38439,N_37549);
and U41127 (N_41127,N_38659,N_39020);
xor U41128 (N_41128,N_39629,N_39849);
or U41129 (N_41129,N_37593,N_39096);
xnor U41130 (N_41130,N_38041,N_37919);
nand U41131 (N_41131,N_37838,N_37844);
nand U41132 (N_41132,N_38178,N_39448);
and U41133 (N_41133,N_39590,N_39546);
and U41134 (N_41134,N_37891,N_38963);
xor U41135 (N_41135,N_38339,N_38956);
or U41136 (N_41136,N_39511,N_39877);
or U41137 (N_41137,N_38763,N_38435);
and U41138 (N_41138,N_38081,N_39584);
and U41139 (N_41139,N_38733,N_37633);
nand U41140 (N_41140,N_38208,N_37629);
nand U41141 (N_41141,N_37945,N_37983);
or U41142 (N_41142,N_38964,N_37711);
or U41143 (N_41143,N_39379,N_39106);
or U41144 (N_41144,N_39350,N_37866);
xor U41145 (N_41145,N_38404,N_37519);
nand U41146 (N_41146,N_37599,N_39890);
and U41147 (N_41147,N_39475,N_38764);
nand U41148 (N_41148,N_39542,N_37576);
nor U41149 (N_41149,N_39508,N_38295);
and U41150 (N_41150,N_39635,N_37630);
or U41151 (N_41151,N_39859,N_38077);
xnor U41152 (N_41152,N_38666,N_39433);
or U41153 (N_41153,N_37546,N_39862);
nor U41154 (N_41154,N_37752,N_39323);
nand U41155 (N_41155,N_39984,N_38302);
or U41156 (N_41156,N_38323,N_38656);
xnor U41157 (N_41157,N_39330,N_39846);
nand U41158 (N_41158,N_39037,N_37970);
nor U41159 (N_41159,N_37666,N_38987);
xor U41160 (N_41160,N_39280,N_38800);
nor U41161 (N_41161,N_39294,N_39073);
nor U41162 (N_41162,N_37730,N_38854);
nor U41163 (N_41163,N_39967,N_38906);
nand U41164 (N_41164,N_37545,N_39576);
xnor U41165 (N_41165,N_38011,N_38112);
xnor U41166 (N_41166,N_39237,N_38245);
or U41167 (N_41167,N_37580,N_39509);
xnor U41168 (N_41168,N_38065,N_38467);
and U41169 (N_41169,N_38739,N_38148);
nand U41170 (N_41170,N_37530,N_39121);
and U41171 (N_41171,N_39044,N_39733);
and U41172 (N_41172,N_39640,N_39261);
and U41173 (N_41173,N_38134,N_38506);
or U41174 (N_41174,N_38362,N_38673);
nand U41175 (N_41175,N_38694,N_38227);
nand U41176 (N_41176,N_38359,N_39114);
nand U41177 (N_41177,N_38232,N_38811);
or U41178 (N_41178,N_39839,N_37728);
xor U41179 (N_41179,N_39056,N_37993);
xor U41180 (N_41180,N_39585,N_37825);
and U41181 (N_41181,N_38959,N_37677);
or U41182 (N_41182,N_39907,N_38955);
or U41183 (N_41183,N_39560,N_37816);
xor U41184 (N_41184,N_38244,N_38611);
or U41185 (N_41185,N_39828,N_38040);
xor U41186 (N_41186,N_38669,N_38199);
and U41187 (N_41187,N_37676,N_39915);
or U41188 (N_41188,N_37976,N_37887);
nor U41189 (N_41189,N_38106,N_39413);
nand U41190 (N_41190,N_39982,N_39278);
and U41191 (N_41191,N_39693,N_37529);
nor U41192 (N_41192,N_37602,N_38646);
or U41193 (N_41193,N_38210,N_39189);
xor U41194 (N_41194,N_37622,N_37892);
nand U41195 (N_41195,N_37979,N_37988);
nor U41196 (N_41196,N_39918,N_38371);
nor U41197 (N_41197,N_39889,N_38155);
or U41198 (N_41198,N_38708,N_37578);
nand U41199 (N_41199,N_37621,N_39036);
and U41200 (N_41200,N_39212,N_38537);
and U41201 (N_41201,N_39149,N_38758);
nand U41202 (N_41202,N_39283,N_39185);
xor U41203 (N_41203,N_37934,N_37682);
nand U41204 (N_41204,N_38114,N_39856);
and U41205 (N_41205,N_37837,N_39652);
xor U41206 (N_41206,N_38836,N_39401);
nand U41207 (N_41207,N_37726,N_39075);
or U41208 (N_41208,N_37617,N_37978);
nor U41209 (N_41209,N_39768,N_39578);
nor U41210 (N_41210,N_39595,N_38188);
or U41211 (N_41211,N_38014,N_38889);
and U41212 (N_41212,N_39151,N_39583);
or U41213 (N_41213,N_39742,N_38421);
nor U41214 (N_41214,N_38932,N_37751);
xnor U41215 (N_41215,N_39395,N_38798);
nand U41216 (N_41216,N_39289,N_38384);
nor U41217 (N_41217,N_39127,N_38909);
nor U41218 (N_41218,N_38375,N_37724);
nor U41219 (N_41219,N_39440,N_39995);
nand U41220 (N_41220,N_38478,N_38870);
or U41221 (N_41221,N_38711,N_38934);
and U41222 (N_41222,N_39741,N_38070);
nor U41223 (N_41223,N_39418,N_38680);
or U41224 (N_41224,N_39632,N_38779);
nand U41225 (N_41225,N_38431,N_37775);
or U41226 (N_41226,N_39399,N_37603);
and U41227 (N_41227,N_37902,N_38073);
or U41228 (N_41228,N_38887,N_38441);
and U41229 (N_41229,N_38092,N_39736);
nor U41230 (N_41230,N_38991,N_38691);
and U41231 (N_41231,N_37911,N_38024);
or U41232 (N_41232,N_39519,N_38942);
nor U41233 (N_41233,N_38428,N_37994);
or U41234 (N_41234,N_38207,N_38306);
nor U41235 (N_41235,N_39182,N_39916);
and U41236 (N_41236,N_39677,N_39588);
nand U41237 (N_41237,N_39735,N_37933);
xnor U41238 (N_41238,N_38770,N_38291);
and U41239 (N_41239,N_39700,N_37920);
xor U41240 (N_41240,N_39946,N_38883);
or U41241 (N_41241,N_38504,N_38697);
xor U41242 (N_41242,N_37764,N_37975);
xor U41243 (N_41243,N_37906,N_39472);
or U41244 (N_41244,N_39041,N_37989);
and U41245 (N_41245,N_37761,N_38687);
nor U41246 (N_41246,N_39985,N_38234);
nor U41247 (N_41247,N_39821,N_38916);
nor U41248 (N_41248,N_37805,N_37960);
or U41249 (N_41249,N_37828,N_37826);
and U41250 (N_41250,N_38114,N_38567);
nor U41251 (N_41251,N_38098,N_38948);
and U41252 (N_41252,N_38921,N_39692);
nor U41253 (N_41253,N_39304,N_39478);
xor U41254 (N_41254,N_39565,N_39592);
or U41255 (N_41255,N_39503,N_38043);
nor U41256 (N_41256,N_38824,N_38961);
and U41257 (N_41257,N_39454,N_39925);
nor U41258 (N_41258,N_38721,N_39814);
nand U41259 (N_41259,N_39576,N_37966);
or U41260 (N_41260,N_38369,N_38535);
nand U41261 (N_41261,N_39891,N_38185);
and U41262 (N_41262,N_38715,N_39355);
xnor U41263 (N_41263,N_39363,N_39213);
xor U41264 (N_41264,N_39383,N_39535);
or U41265 (N_41265,N_39167,N_38102);
and U41266 (N_41266,N_38397,N_39390);
or U41267 (N_41267,N_39545,N_38089);
nor U41268 (N_41268,N_38414,N_37661);
and U41269 (N_41269,N_38314,N_39522);
nor U41270 (N_41270,N_39306,N_39901);
or U41271 (N_41271,N_38271,N_37995);
xnor U41272 (N_41272,N_37983,N_39938);
nor U41273 (N_41273,N_39538,N_38642);
nand U41274 (N_41274,N_38526,N_39038);
and U41275 (N_41275,N_38165,N_38091);
nand U41276 (N_41276,N_39931,N_38053);
and U41277 (N_41277,N_39356,N_37748);
nand U41278 (N_41278,N_39961,N_38298);
or U41279 (N_41279,N_37849,N_38816);
xor U41280 (N_41280,N_39765,N_37984);
nor U41281 (N_41281,N_39000,N_38894);
nand U41282 (N_41282,N_37717,N_37610);
nor U41283 (N_41283,N_37518,N_39494);
nor U41284 (N_41284,N_38583,N_39619);
or U41285 (N_41285,N_38000,N_39091);
xnor U41286 (N_41286,N_38544,N_37520);
nand U41287 (N_41287,N_39501,N_38727);
or U41288 (N_41288,N_39751,N_39284);
or U41289 (N_41289,N_38048,N_39987);
nor U41290 (N_41290,N_39938,N_37581);
or U41291 (N_41291,N_38803,N_37828);
and U41292 (N_41292,N_38515,N_39271);
nor U41293 (N_41293,N_38177,N_39094);
nand U41294 (N_41294,N_39953,N_39819);
or U41295 (N_41295,N_39725,N_37796);
or U41296 (N_41296,N_38254,N_38919);
nor U41297 (N_41297,N_38392,N_38779);
xor U41298 (N_41298,N_39808,N_39498);
nor U41299 (N_41299,N_37794,N_38120);
and U41300 (N_41300,N_38249,N_38448);
nor U41301 (N_41301,N_38704,N_38649);
or U41302 (N_41302,N_39614,N_37863);
nor U41303 (N_41303,N_38883,N_38992);
or U41304 (N_41304,N_38581,N_38037);
xnor U41305 (N_41305,N_39846,N_38405);
nand U41306 (N_41306,N_38559,N_39360);
nand U41307 (N_41307,N_38710,N_37809);
xnor U41308 (N_41308,N_39788,N_37721);
nand U41309 (N_41309,N_37985,N_39155);
nand U41310 (N_41310,N_38537,N_38571);
xor U41311 (N_41311,N_37648,N_38257);
nor U41312 (N_41312,N_38321,N_38821);
nor U41313 (N_41313,N_37631,N_39250);
nand U41314 (N_41314,N_39203,N_38225);
or U41315 (N_41315,N_39885,N_38268);
nor U41316 (N_41316,N_39603,N_39771);
nor U41317 (N_41317,N_39596,N_38597);
and U41318 (N_41318,N_38135,N_39136);
nand U41319 (N_41319,N_39533,N_38282);
or U41320 (N_41320,N_38081,N_38643);
nor U41321 (N_41321,N_38991,N_39133);
xor U41322 (N_41322,N_38215,N_38346);
or U41323 (N_41323,N_38303,N_38043);
nor U41324 (N_41324,N_38577,N_39832);
or U41325 (N_41325,N_38507,N_38817);
xnor U41326 (N_41326,N_38460,N_38663);
or U41327 (N_41327,N_39330,N_37891);
nand U41328 (N_41328,N_37808,N_39929);
nor U41329 (N_41329,N_39994,N_37984);
xor U41330 (N_41330,N_38579,N_39840);
xnor U41331 (N_41331,N_38089,N_38095);
xnor U41332 (N_41332,N_37646,N_37751);
nor U41333 (N_41333,N_38228,N_37636);
xnor U41334 (N_41334,N_38638,N_39734);
nor U41335 (N_41335,N_39704,N_37632);
or U41336 (N_41336,N_39107,N_38747);
and U41337 (N_41337,N_37930,N_38818);
and U41338 (N_41338,N_37880,N_39689);
nor U41339 (N_41339,N_38331,N_38366);
nor U41340 (N_41340,N_38618,N_38709);
or U41341 (N_41341,N_39399,N_39306);
or U41342 (N_41342,N_38512,N_39564);
or U41343 (N_41343,N_39323,N_37675);
and U41344 (N_41344,N_37560,N_37648);
and U41345 (N_41345,N_38828,N_37757);
xnor U41346 (N_41346,N_39338,N_39369);
nor U41347 (N_41347,N_39274,N_38593);
nor U41348 (N_41348,N_37552,N_37616);
nand U41349 (N_41349,N_39587,N_39800);
nand U41350 (N_41350,N_39357,N_38065);
nand U41351 (N_41351,N_38766,N_39966);
nand U41352 (N_41352,N_38278,N_38938);
nand U41353 (N_41353,N_38234,N_39095);
nor U41354 (N_41354,N_39553,N_39025);
xnor U41355 (N_41355,N_38900,N_38447);
or U41356 (N_41356,N_39007,N_39259);
nand U41357 (N_41357,N_39983,N_38334);
and U41358 (N_41358,N_39354,N_37580);
xor U41359 (N_41359,N_38140,N_38373);
nand U41360 (N_41360,N_39275,N_39559);
nor U41361 (N_41361,N_37543,N_39884);
or U41362 (N_41362,N_39298,N_37897);
xnor U41363 (N_41363,N_39219,N_39630);
and U41364 (N_41364,N_39995,N_39268);
nand U41365 (N_41365,N_39824,N_38163);
nor U41366 (N_41366,N_38306,N_38242);
nand U41367 (N_41367,N_38519,N_39721);
or U41368 (N_41368,N_39020,N_39135);
nor U41369 (N_41369,N_38465,N_37889);
or U41370 (N_41370,N_39999,N_38435);
or U41371 (N_41371,N_37999,N_38032);
nand U41372 (N_41372,N_38886,N_39775);
or U41373 (N_41373,N_37506,N_38648);
and U41374 (N_41374,N_39336,N_38317);
nor U41375 (N_41375,N_37664,N_37910);
xnor U41376 (N_41376,N_39006,N_38816);
or U41377 (N_41377,N_39965,N_38857);
or U41378 (N_41378,N_38351,N_39058);
nand U41379 (N_41379,N_39174,N_38970);
or U41380 (N_41380,N_39406,N_39404);
or U41381 (N_41381,N_39368,N_38860);
and U41382 (N_41382,N_38082,N_39542);
and U41383 (N_41383,N_38258,N_37702);
and U41384 (N_41384,N_39089,N_38804);
nand U41385 (N_41385,N_38145,N_39487);
and U41386 (N_41386,N_39188,N_38831);
xor U41387 (N_41387,N_38492,N_38653);
nor U41388 (N_41388,N_39649,N_39959);
xor U41389 (N_41389,N_39767,N_37544);
or U41390 (N_41390,N_39066,N_39907);
nor U41391 (N_41391,N_39647,N_39063);
and U41392 (N_41392,N_37851,N_39674);
and U41393 (N_41393,N_37755,N_37725);
and U41394 (N_41394,N_38299,N_37678);
xor U41395 (N_41395,N_37521,N_39240);
xnor U41396 (N_41396,N_38288,N_39751);
and U41397 (N_41397,N_38856,N_39075);
and U41398 (N_41398,N_38777,N_39433);
nor U41399 (N_41399,N_39575,N_38672);
nand U41400 (N_41400,N_38442,N_39058);
nor U41401 (N_41401,N_38999,N_39074);
or U41402 (N_41402,N_38564,N_39533);
or U41403 (N_41403,N_38666,N_39891);
and U41404 (N_41404,N_39347,N_38781);
nor U41405 (N_41405,N_39799,N_37651);
xor U41406 (N_41406,N_39879,N_39920);
or U41407 (N_41407,N_39281,N_37933);
nand U41408 (N_41408,N_39576,N_39735);
nor U41409 (N_41409,N_38002,N_39804);
or U41410 (N_41410,N_37874,N_37832);
or U41411 (N_41411,N_39983,N_39897);
nor U41412 (N_41412,N_39014,N_38211);
or U41413 (N_41413,N_38887,N_39080);
and U41414 (N_41414,N_38897,N_39793);
xnor U41415 (N_41415,N_37736,N_37695);
nor U41416 (N_41416,N_38658,N_38389);
nor U41417 (N_41417,N_38444,N_38826);
xor U41418 (N_41418,N_38827,N_37850);
nand U41419 (N_41419,N_39949,N_38339);
nor U41420 (N_41420,N_38744,N_39109);
nand U41421 (N_41421,N_38458,N_38037);
xnor U41422 (N_41422,N_39710,N_38495);
or U41423 (N_41423,N_38667,N_37882);
nor U41424 (N_41424,N_37693,N_37607);
xnor U41425 (N_41425,N_38082,N_38508);
or U41426 (N_41426,N_37539,N_39664);
and U41427 (N_41427,N_37520,N_38336);
nor U41428 (N_41428,N_37925,N_39350);
or U41429 (N_41429,N_37819,N_39861);
and U41430 (N_41430,N_38865,N_38357);
and U41431 (N_41431,N_38972,N_39931);
or U41432 (N_41432,N_39048,N_39523);
nor U41433 (N_41433,N_37941,N_38966);
nor U41434 (N_41434,N_38039,N_39276);
nand U41435 (N_41435,N_39015,N_38951);
or U41436 (N_41436,N_38431,N_38556);
nand U41437 (N_41437,N_39162,N_39664);
xor U41438 (N_41438,N_38660,N_39782);
nand U41439 (N_41439,N_37916,N_37864);
or U41440 (N_41440,N_38508,N_39179);
nor U41441 (N_41441,N_39370,N_37928);
nor U41442 (N_41442,N_39793,N_39618);
nor U41443 (N_41443,N_37562,N_39225);
and U41444 (N_41444,N_38136,N_38382);
nand U41445 (N_41445,N_37704,N_39626);
and U41446 (N_41446,N_37742,N_39071);
and U41447 (N_41447,N_37786,N_38595);
nor U41448 (N_41448,N_38902,N_39602);
nand U41449 (N_41449,N_37957,N_37933);
xor U41450 (N_41450,N_39626,N_39717);
xnor U41451 (N_41451,N_38637,N_38729);
or U41452 (N_41452,N_37669,N_38734);
xor U41453 (N_41453,N_38259,N_39718);
nor U41454 (N_41454,N_39175,N_39367);
nand U41455 (N_41455,N_39887,N_39916);
nand U41456 (N_41456,N_37560,N_38794);
nor U41457 (N_41457,N_38201,N_38515);
xor U41458 (N_41458,N_38258,N_38843);
nand U41459 (N_41459,N_38970,N_38755);
nor U41460 (N_41460,N_38452,N_38450);
and U41461 (N_41461,N_37991,N_38908);
nand U41462 (N_41462,N_38774,N_39870);
nand U41463 (N_41463,N_38532,N_39275);
nor U41464 (N_41464,N_39849,N_39182);
nand U41465 (N_41465,N_39183,N_37736);
and U41466 (N_41466,N_39900,N_37592);
nand U41467 (N_41467,N_38521,N_38655);
nand U41468 (N_41468,N_39144,N_37753);
nor U41469 (N_41469,N_37638,N_39280);
and U41470 (N_41470,N_37756,N_39410);
xor U41471 (N_41471,N_37531,N_37538);
or U41472 (N_41472,N_38390,N_38048);
or U41473 (N_41473,N_39922,N_38762);
and U41474 (N_41474,N_39500,N_38424);
nand U41475 (N_41475,N_39701,N_39643);
or U41476 (N_41476,N_39546,N_38029);
or U41477 (N_41477,N_39667,N_39069);
xnor U41478 (N_41478,N_38564,N_38027);
nand U41479 (N_41479,N_39666,N_37625);
nor U41480 (N_41480,N_38781,N_38108);
nand U41481 (N_41481,N_37995,N_39314);
or U41482 (N_41482,N_38324,N_39887);
or U41483 (N_41483,N_37944,N_39839);
nand U41484 (N_41484,N_39402,N_38232);
nor U41485 (N_41485,N_39467,N_38056);
nor U41486 (N_41486,N_38475,N_39445);
xnor U41487 (N_41487,N_37924,N_38391);
nor U41488 (N_41488,N_38540,N_39135);
and U41489 (N_41489,N_38489,N_39822);
xor U41490 (N_41490,N_39351,N_37710);
or U41491 (N_41491,N_38484,N_39404);
and U41492 (N_41492,N_39134,N_38038);
xnor U41493 (N_41493,N_37643,N_38983);
or U41494 (N_41494,N_38354,N_37729);
xor U41495 (N_41495,N_38463,N_38370);
and U41496 (N_41496,N_39454,N_39054);
xnor U41497 (N_41497,N_39387,N_39399);
xor U41498 (N_41498,N_39401,N_38035);
or U41499 (N_41499,N_38311,N_39530);
nor U41500 (N_41500,N_37573,N_39879);
or U41501 (N_41501,N_39914,N_39639);
xnor U41502 (N_41502,N_39910,N_39963);
nand U41503 (N_41503,N_39455,N_39210);
or U41504 (N_41504,N_37961,N_37563);
xnor U41505 (N_41505,N_38950,N_39539);
nand U41506 (N_41506,N_38396,N_39450);
and U41507 (N_41507,N_38433,N_38191);
xnor U41508 (N_41508,N_38922,N_38018);
or U41509 (N_41509,N_37680,N_39484);
nand U41510 (N_41510,N_39024,N_38743);
and U41511 (N_41511,N_39890,N_39050);
nand U41512 (N_41512,N_39589,N_39217);
or U41513 (N_41513,N_39648,N_39828);
and U41514 (N_41514,N_39106,N_38224);
nor U41515 (N_41515,N_37925,N_39640);
nand U41516 (N_41516,N_39884,N_39407);
nand U41517 (N_41517,N_39196,N_38349);
or U41518 (N_41518,N_39403,N_37557);
and U41519 (N_41519,N_37728,N_39317);
nor U41520 (N_41520,N_38651,N_38196);
nand U41521 (N_41521,N_37629,N_39666);
and U41522 (N_41522,N_38492,N_39982);
or U41523 (N_41523,N_39741,N_39160);
or U41524 (N_41524,N_37665,N_38788);
nor U41525 (N_41525,N_38372,N_38264);
and U41526 (N_41526,N_37790,N_39781);
xnor U41527 (N_41527,N_38103,N_38390);
nand U41528 (N_41528,N_39656,N_38730);
xor U41529 (N_41529,N_38783,N_38611);
xnor U41530 (N_41530,N_39241,N_37713);
nor U41531 (N_41531,N_38464,N_38322);
and U41532 (N_41532,N_37927,N_38844);
and U41533 (N_41533,N_39830,N_39928);
nor U41534 (N_41534,N_39100,N_37846);
nor U41535 (N_41535,N_39211,N_38613);
and U41536 (N_41536,N_38043,N_37902);
or U41537 (N_41537,N_38287,N_38359);
nor U41538 (N_41538,N_39432,N_39737);
or U41539 (N_41539,N_39054,N_39774);
xnor U41540 (N_41540,N_38395,N_38405);
nor U41541 (N_41541,N_38171,N_39542);
nor U41542 (N_41542,N_39315,N_39944);
and U41543 (N_41543,N_38446,N_37797);
nor U41544 (N_41544,N_38057,N_38799);
and U41545 (N_41545,N_37829,N_38145);
xnor U41546 (N_41546,N_39861,N_38093);
nor U41547 (N_41547,N_38554,N_37692);
nand U41548 (N_41548,N_37925,N_39016);
or U41549 (N_41549,N_38012,N_39632);
nor U41550 (N_41550,N_39288,N_38871);
nand U41551 (N_41551,N_38744,N_38997);
xor U41552 (N_41552,N_38844,N_38445);
nand U41553 (N_41553,N_39179,N_38298);
nand U41554 (N_41554,N_37551,N_37804);
or U41555 (N_41555,N_39280,N_38888);
and U41556 (N_41556,N_39547,N_37696);
or U41557 (N_41557,N_38312,N_38692);
nor U41558 (N_41558,N_39748,N_38676);
nor U41559 (N_41559,N_38730,N_38370);
and U41560 (N_41560,N_38248,N_39488);
nand U41561 (N_41561,N_38834,N_39549);
nand U41562 (N_41562,N_38403,N_39672);
nor U41563 (N_41563,N_38239,N_38154);
and U41564 (N_41564,N_39095,N_37864);
nor U41565 (N_41565,N_37798,N_37800);
xor U41566 (N_41566,N_37858,N_38034);
nand U41567 (N_41567,N_37726,N_38222);
nor U41568 (N_41568,N_38727,N_39077);
and U41569 (N_41569,N_37991,N_37639);
xor U41570 (N_41570,N_37735,N_39433);
nand U41571 (N_41571,N_38331,N_37567);
nand U41572 (N_41572,N_37504,N_37646);
and U41573 (N_41573,N_38148,N_38485);
nand U41574 (N_41574,N_38031,N_38567);
nand U41575 (N_41575,N_38936,N_39085);
nor U41576 (N_41576,N_37972,N_38013);
and U41577 (N_41577,N_37910,N_38309);
xnor U41578 (N_41578,N_39369,N_38839);
nand U41579 (N_41579,N_38218,N_39162);
xor U41580 (N_41580,N_37660,N_38827);
and U41581 (N_41581,N_39166,N_38532);
or U41582 (N_41582,N_39352,N_38867);
nor U41583 (N_41583,N_37940,N_38381);
or U41584 (N_41584,N_39819,N_38243);
or U41585 (N_41585,N_39821,N_38974);
or U41586 (N_41586,N_39394,N_39603);
or U41587 (N_41587,N_37656,N_38301);
or U41588 (N_41588,N_39698,N_37908);
nor U41589 (N_41589,N_38530,N_39007);
nor U41590 (N_41590,N_39415,N_39647);
xor U41591 (N_41591,N_38934,N_39713);
or U41592 (N_41592,N_39498,N_37918);
nand U41593 (N_41593,N_38037,N_38298);
and U41594 (N_41594,N_39749,N_39921);
xnor U41595 (N_41595,N_38037,N_38717);
nand U41596 (N_41596,N_37585,N_39054);
nand U41597 (N_41597,N_38381,N_39784);
nor U41598 (N_41598,N_38634,N_39373);
nand U41599 (N_41599,N_39162,N_39623);
nor U41600 (N_41600,N_39670,N_37882);
xnor U41601 (N_41601,N_37747,N_38550);
xor U41602 (N_41602,N_39908,N_39033);
or U41603 (N_41603,N_38617,N_39668);
xnor U41604 (N_41604,N_38393,N_37580);
nor U41605 (N_41605,N_37508,N_38292);
xor U41606 (N_41606,N_38444,N_37977);
or U41607 (N_41607,N_39531,N_38906);
nand U41608 (N_41608,N_38728,N_39055);
xnor U41609 (N_41609,N_39997,N_39768);
xor U41610 (N_41610,N_38783,N_38286);
nor U41611 (N_41611,N_38709,N_39976);
nand U41612 (N_41612,N_38459,N_38858);
or U41613 (N_41613,N_39292,N_39340);
nand U41614 (N_41614,N_37867,N_39650);
and U41615 (N_41615,N_39778,N_37533);
nand U41616 (N_41616,N_38232,N_39981);
xnor U41617 (N_41617,N_37735,N_39965);
nor U41618 (N_41618,N_39921,N_38177);
or U41619 (N_41619,N_38174,N_39574);
nand U41620 (N_41620,N_38127,N_39487);
nand U41621 (N_41621,N_38909,N_39618);
and U41622 (N_41622,N_39122,N_38953);
nand U41623 (N_41623,N_37660,N_38805);
xnor U41624 (N_41624,N_39979,N_38181);
or U41625 (N_41625,N_38808,N_39048);
or U41626 (N_41626,N_38576,N_37519);
or U41627 (N_41627,N_39029,N_38750);
xnor U41628 (N_41628,N_39905,N_39145);
nor U41629 (N_41629,N_37715,N_39981);
and U41630 (N_41630,N_37590,N_39243);
nand U41631 (N_41631,N_38398,N_38145);
or U41632 (N_41632,N_37600,N_39076);
xor U41633 (N_41633,N_39057,N_39076);
nor U41634 (N_41634,N_38817,N_38191);
xor U41635 (N_41635,N_39675,N_39437);
and U41636 (N_41636,N_37663,N_39881);
nand U41637 (N_41637,N_37764,N_38843);
and U41638 (N_41638,N_39371,N_37501);
xor U41639 (N_41639,N_37695,N_39832);
nor U41640 (N_41640,N_37533,N_38570);
and U41641 (N_41641,N_37543,N_39447);
and U41642 (N_41642,N_38790,N_37746);
nor U41643 (N_41643,N_39722,N_39557);
nor U41644 (N_41644,N_39703,N_38479);
xnor U41645 (N_41645,N_38219,N_37526);
nor U41646 (N_41646,N_38980,N_37749);
and U41647 (N_41647,N_39806,N_39809);
or U41648 (N_41648,N_39409,N_39896);
nand U41649 (N_41649,N_39908,N_38164);
nor U41650 (N_41650,N_39293,N_38328);
and U41651 (N_41651,N_39108,N_37953);
xor U41652 (N_41652,N_39937,N_39444);
nand U41653 (N_41653,N_38411,N_38461);
and U41654 (N_41654,N_39997,N_38574);
xnor U41655 (N_41655,N_38351,N_37785);
xnor U41656 (N_41656,N_39003,N_39385);
nor U41657 (N_41657,N_39405,N_38418);
or U41658 (N_41658,N_38441,N_38594);
or U41659 (N_41659,N_38392,N_39529);
or U41660 (N_41660,N_39080,N_37602);
nand U41661 (N_41661,N_38509,N_38146);
or U41662 (N_41662,N_38948,N_39365);
nand U41663 (N_41663,N_38133,N_38468);
xnor U41664 (N_41664,N_37708,N_39469);
nand U41665 (N_41665,N_38964,N_38775);
xor U41666 (N_41666,N_38416,N_39232);
xnor U41667 (N_41667,N_38454,N_39457);
or U41668 (N_41668,N_39526,N_39560);
xor U41669 (N_41669,N_38914,N_39629);
or U41670 (N_41670,N_38827,N_39367);
and U41671 (N_41671,N_38450,N_37803);
nor U41672 (N_41672,N_38963,N_39735);
and U41673 (N_41673,N_39290,N_38056);
or U41674 (N_41674,N_39366,N_39401);
and U41675 (N_41675,N_37761,N_37510);
or U41676 (N_41676,N_38415,N_38502);
xnor U41677 (N_41677,N_39990,N_38304);
xor U41678 (N_41678,N_39459,N_39297);
and U41679 (N_41679,N_38798,N_37572);
xnor U41680 (N_41680,N_38084,N_39808);
nand U41681 (N_41681,N_38317,N_37710);
nor U41682 (N_41682,N_38043,N_38502);
nand U41683 (N_41683,N_38602,N_38398);
and U41684 (N_41684,N_38002,N_38577);
xor U41685 (N_41685,N_39651,N_39410);
and U41686 (N_41686,N_38456,N_39687);
nand U41687 (N_41687,N_39149,N_39068);
nor U41688 (N_41688,N_38284,N_38038);
nor U41689 (N_41689,N_39252,N_38525);
and U41690 (N_41690,N_38697,N_37756);
xor U41691 (N_41691,N_38637,N_37968);
nand U41692 (N_41692,N_38633,N_38744);
or U41693 (N_41693,N_39355,N_38329);
nand U41694 (N_41694,N_39319,N_39580);
or U41695 (N_41695,N_39278,N_39774);
xnor U41696 (N_41696,N_39637,N_37679);
nor U41697 (N_41697,N_39029,N_37669);
and U41698 (N_41698,N_37945,N_39623);
nand U41699 (N_41699,N_37888,N_37781);
or U41700 (N_41700,N_38246,N_39301);
xor U41701 (N_41701,N_39919,N_39715);
nand U41702 (N_41702,N_39890,N_37803);
and U41703 (N_41703,N_38375,N_37899);
xor U41704 (N_41704,N_37892,N_37800);
nor U41705 (N_41705,N_38304,N_38507);
xor U41706 (N_41706,N_39319,N_38202);
nand U41707 (N_41707,N_37726,N_39944);
nand U41708 (N_41708,N_39849,N_38135);
nor U41709 (N_41709,N_38475,N_39846);
nand U41710 (N_41710,N_38146,N_39426);
nand U41711 (N_41711,N_38616,N_38144);
or U41712 (N_41712,N_37973,N_39126);
nor U41713 (N_41713,N_38459,N_38933);
nand U41714 (N_41714,N_38147,N_38413);
xor U41715 (N_41715,N_38341,N_38320);
xor U41716 (N_41716,N_37851,N_39897);
and U41717 (N_41717,N_39163,N_38456);
nor U41718 (N_41718,N_38416,N_38047);
nand U41719 (N_41719,N_39781,N_39875);
nor U41720 (N_41720,N_39830,N_39083);
xnor U41721 (N_41721,N_39667,N_39171);
xnor U41722 (N_41722,N_37989,N_37914);
and U41723 (N_41723,N_38134,N_37686);
nand U41724 (N_41724,N_38699,N_39053);
nand U41725 (N_41725,N_37602,N_37795);
nand U41726 (N_41726,N_39919,N_38177);
nand U41727 (N_41727,N_37523,N_37549);
nor U41728 (N_41728,N_38534,N_39513);
or U41729 (N_41729,N_37587,N_39940);
nand U41730 (N_41730,N_37724,N_39396);
nor U41731 (N_41731,N_37824,N_37877);
nor U41732 (N_41732,N_37919,N_38721);
nand U41733 (N_41733,N_39085,N_39545);
or U41734 (N_41734,N_39961,N_37789);
nand U41735 (N_41735,N_38797,N_39382);
nand U41736 (N_41736,N_39771,N_39179);
and U41737 (N_41737,N_38009,N_38377);
and U41738 (N_41738,N_39244,N_38688);
xnor U41739 (N_41739,N_37746,N_38711);
nand U41740 (N_41740,N_37915,N_39904);
or U41741 (N_41741,N_37776,N_39451);
xnor U41742 (N_41742,N_38962,N_39682);
nor U41743 (N_41743,N_37677,N_38682);
or U41744 (N_41744,N_37925,N_37558);
nor U41745 (N_41745,N_38559,N_39050);
or U41746 (N_41746,N_38475,N_37657);
nor U41747 (N_41747,N_37966,N_38823);
or U41748 (N_41748,N_39461,N_39199);
xor U41749 (N_41749,N_38143,N_38339);
and U41750 (N_41750,N_39671,N_38963);
xnor U41751 (N_41751,N_39460,N_38705);
nor U41752 (N_41752,N_39193,N_39610);
and U41753 (N_41753,N_37656,N_39637);
nor U41754 (N_41754,N_37621,N_39350);
nand U41755 (N_41755,N_37806,N_39101);
and U41756 (N_41756,N_39020,N_38245);
nor U41757 (N_41757,N_39048,N_38977);
nor U41758 (N_41758,N_38582,N_39108);
nand U41759 (N_41759,N_37603,N_37789);
or U41760 (N_41760,N_37818,N_39898);
or U41761 (N_41761,N_37552,N_39483);
or U41762 (N_41762,N_38599,N_37815);
nand U41763 (N_41763,N_38856,N_38694);
or U41764 (N_41764,N_38625,N_38696);
nor U41765 (N_41765,N_38358,N_38545);
nor U41766 (N_41766,N_39833,N_38890);
xor U41767 (N_41767,N_39769,N_38251);
xor U41768 (N_41768,N_38522,N_39306);
nor U41769 (N_41769,N_39502,N_37767);
nor U41770 (N_41770,N_38701,N_38465);
or U41771 (N_41771,N_39794,N_39778);
nand U41772 (N_41772,N_39273,N_39233);
nand U41773 (N_41773,N_38482,N_39467);
xor U41774 (N_41774,N_39117,N_38749);
xnor U41775 (N_41775,N_38940,N_39474);
and U41776 (N_41776,N_39199,N_39585);
nor U41777 (N_41777,N_38025,N_38050);
and U41778 (N_41778,N_38265,N_37869);
nand U41779 (N_41779,N_38724,N_39715);
nor U41780 (N_41780,N_38578,N_39161);
nor U41781 (N_41781,N_37635,N_39773);
or U41782 (N_41782,N_38695,N_38683);
nand U41783 (N_41783,N_37512,N_38502);
xor U41784 (N_41784,N_38879,N_38443);
xor U41785 (N_41785,N_39025,N_38297);
and U41786 (N_41786,N_38075,N_39209);
and U41787 (N_41787,N_39387,N_37841);
nand U41788 (N_41788,N_37520,N_38903);
or U41789 (N_41789,N_37719,N_39051);
xnor U41790 (N_41790,N_39937,N_38223);
or U41791 (N_41791,N_37599,N_39930);
and U41792 (N_41792,N_37724,N_38162);
and U41793 (N_41793,N_38276,N_39998);
xnor U41794 (N_41794,N_39493,N_38609);
nor U41795 (N_41795,N_39741,N_38967);
xnor U41796 (N_41796,N_38611,N_39390);
and U41797 (N_41797,N_38868,N_38066);
nand U41798 (N_41798,N_38700,N_39663);
xor U41799 (N_41799,N_39461,N_38925);
nor U41800 (N_41800,N_38735,N_39189);
and U41801 (N_41801,N_39381,N_38646);
xnor U41802 (N_41802,N_39787,N_38718);
or U41803 (N_41803,N_38378,N_39342);
and U41804 (N_41804,N_37625,N_37552);
nor U41805 (N_41805,N_37829,N_39607);
xor U41806 (N_41806,N_37981,N_38897);
or U41807 (N_41807,N_37849,N_39957);
xor U41808 (N_41808,N_37717,N_39259);
or U41809 (N_41809,N_38621,N_38066);
and U41810 (N_41810,N_39873,N_39021);
or U41811 (N_41811,N_38409,N_38804);
and U41812 (N_41812,N_38512,N_39423);
nand U41813 (N_41813,N_39458,N_39016);
nand U41814 (N_41814,N_38127,N_39793);
nor U41815 (N_41815,N_38814,N_38061);
xnor U41816 (N_41816,N_37825,N_39363);
or U41817 (N_41817,N_39532,N_37693);
nor U41818 (N_41818,N_38653,N_38097);
and U41819 (N_41819,N_38892,N_39513);
xnor U41820 (N_41820,N_37892,N_38451);
and U41821 (N_41821,N_37980,N_37886);
nor U41822 (N_41822,N_39777,N_39559);
nand U41823 (N_41823,N_39306,N_38404);
nor U41824 (N_41824,N_37786,N_38981);
xor U41825 (N_41825,N_39701,N_38204);
or U41826 (N_41826,N_39356,N_37714);
or U41827 (N_41827,N_37948,N_37684);
and U41828 (N_41828,N_39374,N_38394);
nor U41829 (N_41829,N_39856,N_39152);
and U41830 (N_41830,N_37897,N_38343);
xor U41831 (N_41831,N_38469,N_37844);
or U41832 (N_41832,N_38665,N_38950);
nor U41833 (N_41833,N_37881,N_39839);
nor U41834 (N_41834,N_37891,N_37737);
nand U41835 (N_41835,N_39142,N_39761);
and U41836 (N_41836,N_37942,N_37704);
xor U41837 (N_41837,N_39746,N_39900);
or U41838 (N_41838,N_39742,N_38795);
nand U41839 (N_41839,N_38635,N_39008);
or U41840 (N_41840,N_37593,N_38470);
nor U41841 (N_41841,N_39650,N_38994);
nor U41842 (N_41842,N_39578,N_38283);
xnor U41843 (N_41843,N_37567,N_39055);
nor U41844 (N_41844,N_38099,N_38058);
nor U41845 (N_41845,N_37944,N_38025);
or U41846 (N_41846,N_39715,N_39826);
and U41847 (N_41847,N_38091,N_39505);
nand U41848 (N_41848,N_38266,N_38253);
xor U41849 (N_41849,N_38167,N_38617);
and U41850 (N_41850,N_39436,N_37837);
and U41851 (N_41851,N_38714,N_38617);
nor U41852 (N_41852,N_39992,N_37935);
nand U41853 (N_41853,N_39977,N_39183);
nor U41854 (N_41854,N_38172,N_37936);
nor U41855 (N_41855,N_39054,N_39390);
xnor U41856 (N_41856,N_38896,N_39500);
and U41857 (N_41857,N_39742,N_39945);
and U41858 (N_41858,N_39553,N_37812);
and U41859 (N_41859,N_38227,N_39679);
and U41860 (N_41860,N_38157,N_39334);
nand U41861 (N_41861,N_37701,N_37847);
xnor U41862 (N_41862,N_38912,N_37707);
and U41863 (N_41863,N_39041,N_38413);
nor U41864 (N_41864,N_38392,N_38802);
and U41865 (N_41865,N_37732,N_37530);
nand U41866 (N_41866,N_39392,N_38809);
and U41867 (N_41867,N_38114,N_38990);
and U41868 (N_41868,N_39602,N_38045);
nand U41869 (N_41869,N_39731,N_38636);
and U41870 (N_41870,N_39265,N_37900);
nor U41871 (N_41871,N_39248,N_38312);
nand U41872 (N_41872,N_38588,N_37657);
nand U41873 (N_41873,N_38375,N_37896);
and U41874 (N_41874,N_39709,N_37738);
and U41875 (N_41875,N_39733,N_38796);
xnor U41876 (N_41876,N_39736,N_38294);
xnor U41877 (N_41877,N_39518,N_38598);
nor U41878 (N_41878,N_38755,N_38500);
or U41879 (N_41879,N_37639,N_39643);
and U41880 (N_41880,N_39973,N_38534);
nor U41881 (N_41881,N_39910,N_39140);
or U41882 (N_41882,N_38222,N_38977);
or U41883 (N_41883,N_37669,N_39738);
or U41884 (N_41884,N_38364,N_38055);
nand U41885 (N_41885,N_37562,N_37950);
nand U41886 (N_41886,N_39756,N_39215);
and U41887 (N_41887,N_37517,N_38505);
nand U41888 (N_41888,N_39086,N_39586);
nand U41889 (N_41889,N_39376,N_38555);
nand U41890 (N_41890,N_37558,N_39108);
and U41891 (N_41891,N_38900,N_39893);
nand U41892 (N_41892,N_39303,N_39136);
xor U41893 (N_41893,N_38718,N_37910);
nor U41894 (N_41894,N_39924,N_38932);
xor U41895 (N_41895,N_37900,N_38015);
nor U41896 (N_41896,N_39630,N_38899);
nor U41897 (N_41897,N_38162,N_39123);
nor U41898 (N_41898,N_38140,N_38712);
nand U41899 (N_41899,N_39858,N_38950);
xnor U41900 (N_41900,N_39734,N_38074);
nand U41901 (N_41901,N_38697,N_37658);
xor U41902 (N_41902,N_39748,N_38683);
and U41903 (N_41903,N_37551,N_38936);
nand U41904 (N_41904,N_39086,N_37519);
xor U41905 (N_41905,N_39232,N_37642);
xnor U41906 (N_41906,N_39840,N_39195);
or U41907 (N_41907,N_38511,N_37727);
and U41908 (N_41908,N_39015,N_38667);
xnor U41909 (N_41909,N_38160,N_39517);
nor U41910 (N_41910,N_37928,N_38912);
nand U41911 (N_41911,N_37536,N_38490);
nand U41912 (N_41912,N_39222,N_38053);
or U41913 (N_41913,N_38067,N_39563);
or U41914 (N_41914,N_39437,N_39612);
nor U41915 (N_41915,N_39529,N_38283);
nand U41916 (N_41916,N_38691,N_39952);
or U41917 (N_41917,N_38673,N_38729);
or U41918 (N_41918,N_38348,N_39292);
and U41919 (N_41919,N_38954,N_38276);
or U41920 (N_41920,N_37883,N_38555);
nand U41921 (N_41921,N_38258,N_39226);
xnor U41922 (N_41922,N_37617,N_38202);
nor U41923 (N_41923,N_39121,N_38034);
xnor U41924 (N_41924,N_39514,N_39838);
nor U41925 (N_41925,N_39122,N_39361);
xor U41926 (N_41926,N_37687,N_38328);
nor U41927 (N_41927,N_38403,N_38414);
xor U41928 (N_41928,N_37632,N_37914);
nand U41929 (N_41929,N_38008,N_39125);
nand U41930 (N_41930,N_39591,N_38928);
or U41931 (N_41931,N_39349,N_38338);
or U41932 (N_41932,N_38741,N_38133);
or U41933 (N_41933,N_39098,N_39687);
or U41934 (N_41934,N_38748,N_39285);
nor U41935 (N_41935,N_39128,N_38947);
or U41936 (N_41936,N_38303,N_37812);
and U41937 (N_41937,N_38006,N_38849);
nor U41938 (N_41938,N_37650,N_38303);
and U41939 (N_41939,N_39907,N_38434);
nor U41940 (N_41940,N_39846,N_39614);
and U41941 (N_41941,N_39622,N_38262);
or U41942 (N_41942,N_39134,N_39809);
xor U41943 (N_41943,N_38268,N_38804);
nor U41944 (N_41944,N_39273,N_39948);
or U41945 (N_41945,N_39140,N_38383);
nor U41946 (N_41946,N_39887,N_39377);
and U41947 (N_41947,N_39035,N_38614);
or U41948 (N_41948,N_38893,N_38154);
and U41949 (N_41949,N_39461,N_37779);
xor U41950 (N_41950,N_37571,N_38958);
nand U41951 (N_41951,N_38259,N_37965);
or U41952 (N_41952,N_39256,N_39575);
or U41953 (N_41953,N_39120,N_37865);
or U41954 (N_41954,N_37682,N_38092);
nand U41955 (N_41955,N_38368,N_38417);
nand U41956 (N_41956,N_37582,N_38558);
and U41957 (N_41957,N_38748,N_38585);
xnor U41958 (N_41958,N_38761,N_39131);
xor U41959 (N_41959,N_38326,N_38551);
or U41960 (N_41960,N_38245,N_39011);
and U41961 (N_41961,N_39614,N_39245);
xor U41962 (N_41962,N_39594,N_38945);
nor U41963 (N_41963,N_38100,N_39097);
and U41964 (N_41964,N_39976,N_37690);
nand U41965 (N_41965,N_39090,N_38643);
or U41966 (N_41966,N_39931,N_39977);
or U41967 (N_41967,N_39902,N_39412);
nor U41968 (N_41968,N_37863,N_38822);
and U41969 (N_41969,N_37600,N_39493);
nand U41970 (N_41970,N_37781,N_39603);
nor U41971 (N_41971,N_38350,N_39809);
nand U41972 (N_41972,N_38369,N_38391);
nor U41973 (N_41973,N_37933,N_39568);
xor U41974 (N_41974,N_38950,N_39387);
xnor U41975 (N_41975,N_38481,N_37877);
nor U41976 (N_41976,N_38190,N_37504);
nand U41977 (N_41977,N_37581,N_39087);
xor U41978 (N_41978,N_38283,N_38203);
and U41979 (N_41979,N_38335,N_37666);
xnor U41980 (N_41980,N_38413,N_39568);
nand U41981 (N_41981,N_37722,N_39807);
and U41982 (N_41982,N_39805,N_38208);
or U41983 (N_41983,N_39761,N_39586);
or U41984 (N_41984,N_38853,N_38958);
xor U41985 (N_41985,N_39194,N_38943);
nand U41986 (N_41986,N_39082,N_38459);
or U41987 (N_41987,N_39930,N_38127);
or U41988 (N_41988,N_39943,N_38667);
or U41989 (N_41989,N_39623,N_38349);
nor U41990 (N_41990,N_38739,N_38484);
nand U41991 (N_41991,N_39973,N_37701);
nor U41992 (N_41992,N_38281,N_38425);
nor U41993 (N_41993,N_39380,N_39661);
and U41994 (N_41994,N_38322,N_39002);
and U41995 (N_41995,N_37703,N_38413);
nor U41996 (N_41996,N_38460,N_39585);
and U41997 (N_41997,N_38316,N_39600);
nand U41998 (N_41998,N_37973,N_38800);
nor U41999 (N_41999,N_39205,N_39279);
or U42000 (N_42000,N_38237,N_38630);
or U42001 (N_42001,N_37977,N_38092);
xnor U42002 (N_42002,N_39081,N_38171);
and U42003 (N_42003,N_38368,N_38464);
or U42004 (N_42004,N_39447,N_37894);
and U42005 (N_42005,N_37626,N_38689);
xnor U42006 (N_42006,N_37831,N_37616);
and U42007 (N_42007,N_37648,N_39754);
or U42008 (N_42008,N_39421,N_38692);
or U42009 (N_42009,N_38710,N_38084);
or U42010 (N_42010,N_39665,N_38846);
xor U42011 (N_42011,N_38135,N_38230);
xor U42012 (N_42012,N_38788,N_38879);
nand U42013 (N_42013,N_39968,N_38197);
nand U42014 (N_42014,N_39834,N_39133);
xnor U42015 (N_42015,N_37507,N_38149);
or U42016 (N_42016,N_39847,N_39520);
nor U42017 (N_42017,N_39706,N_39793);
or U42018 (N_42018,N_38010,N_39082);
xnor U42019 (N_42019,N_38317,N_39334);
nand U42020 (N_42020,N_39848,N_39934);
nor U42021 (N_42021,N_38328,N_38799);
nor U42022 (N_42022,N_38148,N_37676);
nand U42023 (N_42023,N_39972,N_38687);
and U42024 (N_42024,N_38393,N_39405);
nor U42025 (N_42025,N_38485,N_39322);
and U42026 (N_42026,N_37565,N_39855);
or U42027 (N_42027,N_37797,N_37833);
nor U42028 (N_42028,N_39771,N_38149);
nor U42029 (N_42029,N_39880,N_38214);
and U42030 (N_42030,N_39404,N_38357);
and U42031 (N_42031,N_39537,N_39752);
nor U42032 (N_42032,N_38631,N_39411);
or U42033 (N_42033,N_39602,N_37557);
xor U42034 (N_42034,N_38310,N_37593);
xor U42035 (N_42035,N_38181,N_38657);
and U42036 (N_42036,N_39735,N_38049);
and U42037 (N_42037,N_37881,N_38628);
nand U42038 (N_42038,N_39961,N_37771);
nor U42039 (N_42039,N_38142,N_37739);
nand U42040 (N_42040,N_38845,N_38402);
and U42041 (N_42041,N_37905,N_38437);
xor U42042 (N_42042,N_38450,N_38081);
and U42043 (N_42043,N_39443,N_38264);
xnor U42044 (N_42044,N_38584,N_39684);
or U42045 (N_42045,N_38685,N_37691);
or U42046 (N_42046,N_39587,N_38545);
or U42047 (N_42047,N_38951,N_37520);
or U42048 (N_42048,N_37740,N_39642);
nand U42049 (N_42049,N_39132,N_39914);
nand U42050 (N_42050,N_38540,N_37537);
nor U42051 (N_42051,N_38313,N_37839);
and U42052 (N_42052,N_39735,N_39329);
nand U42053 (N_42053,N_39320,N_37872);
xnor U42054 (N_42054,N_38573,N_39340);
and U42055 (N_42055,N_38881,N_38411);
nor U42056 (N_42056,N_37625,N_37985);
or U42057 (N_42057,N_39186,N_37637);
nand U42058 (N_42058,N_37622,N_38732);
nand U42059 (N_42059,N_38949,N_38728);
nor U42060 (N_42060,N_39575,N_39904);
xor U42061 (N_42061,N_38824,N_38466);
xnor U42062 (N_42062,N_38724,N_39775);
nand U42063 (N_42063,N_38921,N_38546);
and U42064 (N_42064,N_38603,N_38217);
and U42065 (N_42065,N_38114,N_38955);
and U42066 (N_42066,N_39657,N_37599);
and U42067 (N_42067,N_39334,N_38081);
or U42068 (N_42068,N_39364,N_37607);
or U42069 (N_42069,N_39460,N_39797);
xnor U42070 (N_42070,N_39333,N_39225);
nor U42071 (N_42071,N_37826,N_38030);
or U42072 (N_42072,N_38810,N_37664);
nor U42073 (N_42073,N_39091,N_39664);
xnor U42074 (N_42074,N_39287,N_39087);
or U42075 (N_42075,N_37948,N_39145);
or U42076 (N_42076,N_37842,N_38421);
nor U42077 (N_42077,N_39782,N_39389);
nand U42078 (N_42078,N_39132,N_37613);
nand U42079 (N_42079,N_37944,N_39096);
nor U42080 (N_42080,N_38787,N_38706);
or U42081 (N_42081,N_38644,N_38985);
nand U42082 (N_42082,N_37705,N_37953);
xor U42083 (N_42083,N_37670,N_38390);
xor U42084 (N_42084,N_37959,N_38748);
nand U42085 (N_42085,N_37524,N_38975);
xor U42086 (N_42086,N_38669,N_38334);
nor U42087 (N_42087,N_38849,N_38857);
nand U42088 (N_42088,N_38352,N_37992);
xor U42089 (N_42089,N_37781,N_37843);
and U42090 (N_42090,N_37562,N_38798);
nor U42091 (N_42091,N_38092,N_39698);
or U42092 (N_42092,N_39426,N_37631);
nand U42093 (N_42093,N_38293,N_39062);
or U42094 (N_42094,N_37982,N_38998);
and U42095 (N_42095,N_39106,N_39474);
and U42096 (N_42096,N_37784,N_38882);
nor U42097 (N_42097,N_38487,N_39165);
xnor U42098 (N_42098,N_39019,N_38232);
xnor U42099 (N_42099,N_38622,N_38914);
nor U42100 (N_42100,N_38739,N_38276);
and U42101 (N_42101,N_39434,N_37522);
and U42102 (N_42102,N_39334,N_37739);
or U42103 (N_42103,N_38373,N_38933);
nand U42104 (N_42104,N_38308,N_38122);
nor U42105 (N_42105,N_37938,N_38887);
nand U42106 (N_42106,N_39847,N_39709);
nor U42107 (N_42107,N_39279,N_38637);
nand U42108 (N_42108,N_38924,N_37841);
nand U42109 (N_42109,N_37986,N_39642);
nand U42110 (N_42110,N_38791,N_38888);
nor U42111 (N_42111,N_37979,N_39960);
or U42112 (N_42112,N_39765,N_37799);
nor U42113 (N_42113,N_39365,N_37957);
nand U42114 (N_42114,N_38610,N_37955);
and U42115 (N_42115,N_37994,N_39090);
nor U42116 (N_42116,N_38604,N_39173);
and U42117 (N_42117,N_38056,N_39426);
or U42118 (N_42118,N_39915,N_39618);
or U42119 (N_42119,N_38246,N_39793);
and U42120 (N_42120,N_39901,N_37778);
xor U42121 (N_42121,N_39782,N_39557);
nor U42122 (N_42122,N_38994,N_38662);
or U42123 (N_42123,N_37584,N_39211);
nand U42124 (N_42124,N_39774,N_39847);
xnor U42125 (N_42125,N_38930,N_38238);
or U42126 (N_42126,N_39380,N_37657);
xor U42127 (N_42127,N_38540,N_37872);
and U42128 (N_42128,N_38439,N_39985);
xnor U42129 (N_42129,N_39455,N_38468);
nor U42130 (N_42130,N_38177,N_39981);
or U42131 (N_42131,N_38642,N_37677);
nand U42132 (N_42132,N_39991,N_39217);
xnor U42133 (N_42133,N_38554,N_38121);
and U42134 (N_42134,N_37769,N_39828);
nor U42135 (N_42135,N_39817,N_38170);
nor U42136 (N_42136,N_38947,N_38980);
nand U42137 (N_42137,N_39436,N_39696);
and U42138 (N_42138,N_37963,N_38147);
nand U42139 (N_42139,N_38079,N_39892);
nor U42140 (N_42140,N_39158,N_38975);
xnor U42141 (N_42141,N_37517,N_39214);
nand U42142 (N_42142,N_38461,N_39201);
nand U42143 (N_42143,N_39325,N_39743);
xor U42144 (N_42144,N_38311,N_39278);
xnor U42145 (N_42145,N_38189,N_39558);
xor U42146 (N_42146,N_37760,N_39665);
or U42147 (N_42147,N_37688,N_37703);
nand U42148 (N_42148,N_39562,N_39288);
nor U42149 (N_42149,N_39380,N_39356);
nor U42150 (N_42150,N_39973,N_38218);
or U42151 (N_42151,N_38982,N_38385);
or U42152 (N_42152,N_38066,N_38660);
xnor U42153 (N_42153,N_39788,N_38712);
nand U42154 (N_42154,N_37928,N_39681);
and U42155 (N_42155,N_38693,N_38417);
and U42156 (N_42156,N_38729,N_38411);
nand U42157 (N_42157,N_39450,N_38452);
nor U42158 (N_42158,N_39333,N_37832);
nand U42159 (N_42159,N_38432,N_39623);
xor U42160 (N_42160,N_39726,N_37848);
or U42161 (N_42161,N_39622,N_39948);
xor U42162 (N_42162,N_39661,N_38519);
xnor U42163 (N_42163,N_38055,N_39542);
xnor U42164 (N_42164,N_39051,N_39292);
xnor U42165 (N_42165,N_38484,N_38514);
and U42166 (N_42166,N_38336,N_37693);
and U42167 (N_42167,N_39548,N_38866);
nand U42168 (N_42168,N_37767,N_38744);
or U42169 (N_42169,N_38870,N_39287);
nand U42170 (N_42170,N_38608,N_39183);
or U42171 (N_42171,N_38431,N_38930);
and U42172 (N_42172,N_39984,N_39711);
and U42173 (N_42173,N_39651,N_37557);
or U42174 (N_42174,N_38122,N_38434);
nor U42175 (N_42175,N_39856,N_38916);
nor U42176 (N_42176,N_39687,N_38836);
or U42177 (N_42177,N_38343,N_39222);
xnor U42178 (N_42178,N_39012,N_37535);
or U42179 (N_42179,N_38697,N_37885);
nand U42180 (N_42180,N_38701,N_38603);
or U42181 (N_42181,N_37722,N_38863);
or U42182 (N_42182,N_39282,N_38451);
nand U42183 (N_42183,N_39246,N_38118);
xnor U42184 (N_42184,N_38355,N_39340);
xor U42185 (N_42185,N_38201,N_38697);
nor U42186 (N_42186,N_39913,N_39008);
xor U42187 (N_42187,N_39933,N_38039);
or U42188 (N_42188,N_38955,N_38880);
nor U42189 (N_42189,N_37517,N_39402);
nor U42190 (N_42190,N_39669,N_39342);
or U42191 (N_42191,N_37883,N_37906);
or U42192 (N_42192,N_38565,N_38300);
nand U42193 (N_42193,N_37699,N_38257);
or U42194 (N_42194,N_39552,N_38497);
xnor U42195 (N_42195,N_39126,N_39727);
or U42196 (N_42196,N_39809,N_39412);
xor U42197 (N_42197,N_37997,N_38579);
and U42198 (N_42198,N_38434,N_38017);
nor U42199 (N_42199,N_38912,N_37961);
nor U42200 (N_42200,N_38767,N_37531);
nor U42201 (N_42201,N_39191,N_39820);
and U42202 (N_42202,N_39585,N_37905);
nand U42203 (N_42203,N_37782,N_38996);
nor U42204 (N_42204,N_39105,N_39789);
and U42205 (N_42205,N_39105,N_38796);
nor U42206 (N_42206,N_37602,N_39743);
xor U42207 (N_42207,N_39497,N_39154);
nor U42208 (N_42208,N_39241,N_39342);
nand U42209 (N_42209,N_39039,N_37532);
or U42210 (N_42210,N_38079,N_39317);
xor U42211 (N_42211,N_39547,N_38354);
xnor U42212 (N_42212,N_38701,N_37772);
and U42213 (N_42213,N_37775,N_39659);
nor U42214 (N_42214,N_38415,N_37748);
or U42215 (N_42215,N_38914,N_39453);
nor U42216 (N_42216,N_38822,N_37984);
and U42217 (N_42217,N_37856,N_39492);
xor U42218 (N_42218,N_38136,N_38272);
nand U42219 (N_42219,N_37987,N_37562);
nand U42220 (N_42220,N_39057,N_39224);
xor U42221 (N_42221,N_39887,N_37901);
nor U42222 (N_42222,N_39373,N_39538);
xnor U42223 (N_42223,N_38547,N_39585);
xor U42224 (N_42224,N_38830,N_38964);
and U42225 (N_42225,N_39886,N_39432);
xnor U42226 (N_42226,N_39951,N_37854);
xnor U42227 (N_42227,N_39570,N_38405);
xor U42228 (N_42228,N_37706,N_37529);
nor U42229 (N_42229,N_39232,N_37961);
nor U42230 (N_42230,N_38192,N_39346);
nor U42231 (N_42231,N_39407,N_39490);
or U42232 (N_42232,N_39985,N_38646);
nor U42233 (N_42233,N_37966,N_37897);
and U42234 (N_42234,N_38301,N_39928);
xnor U42235 (N_42235,N_37796,N_38402);
nor U42236 (N_42236,N_39704,N_38472);
and U42237 (N_42237,N_39856,N_39218);
and U42238 (N_42238,N_39660,N_38731);
and U42239 (N_42239,N_39532,N_37981);
xor U42240 (N_42240,N_39474,N_39100);
and U42241 (N_42241,N_37699,N_39491);
nand U42242 (N_42242,N_38067,N_37743);
xor U42243 (N_42243,N_38868,N_38166);
or U42244 (N_42244,N_39452,N_39765);
nand U42245 (N_42245,N_37904,N_37675);
or U42246 (N_42246,N_39265,N_38313);
and U42247 (N_42247,N_37855,N_37879);
nand U42248 (N_42248,N_39970,N_38279);
nor U42249 (N_42249,N_38229,N_38749);
and U42250 (N_42250,N_39490,N_39765);
nand U42251 (N_42251,N_39881,N_37681);
xor U42252 (N_42252,N_38609,N_38449);
nand U42253 (N_42253,N_38532,N_38379);
and U42254 (N_42254,N_37684,N_38171);
and U42255 (N_42255,N_38321,N_37649);
nand U42256 (N_42256,N_39736,N_39003);
xnor U42257 (N_42257,N_39442,N_38471);
nor U42258 (N_42258,N_39412,N_39260);
nor U42259 (N_42259,N_39119,N_38911);
and U42260 (N_42260,N_38647,N_39323);
or U42261 (N_42261,N_39389,N_39018);
xor U42262 (N_42262,N_39004,N_38860);
and U42263 (N_42263,N_37673,N_38756);
or U42264 (N_42264,N_39543,N_38738);
or U42265 (N_42265,N_39285,N_39844);
or U42266 (N_42266,N_39489,N_39831);
nand U42267 (N_42267,N_39521,N_39978);
xor U42268 (N_42268,N_38779,N_39474);
xnor U42269 (N_42269,N_38153,N_37738);
xor U42270 (N_42270,N_39494,N_37512);
nor U42271 (N_42271,N_37819,N_37728);
xnor U42272 (N_42272,N_37796,N_37574);
and U42273 (N_42273,N_39044,N_39810);
xor U42274 (N_42274,N_37781,N_38248);
nand U42275 (N_42275,N_39809,N_38560);
xor U42276 (N_42276,N_38062,N_37967);
nand U42277 (N_42277,N_38830,N_38460);
or U42278 (N_42278,N_39272,N_37602);
nor U42279 (N_42279,N_39766,N_39458);
xor U42280 (N_42280,N_38520,N_38473);
nand U42281 (N_42281,N_39801,N_38558);
xor U42282 (N_42282,N_39836,N_38002);
xnor U42283 (N_42283,N_39259,N_38735);
xor U42284 (N_42284,N_39092,N_37684);
nor U42285 (N_42285,N_38709,N_38842);
nand U42286 (N_42286,N_39042,N_39698);
nor U42287 (N_42287,N_39048,N_39420);
xnor U42288 (N_42288,N_37912,N_39927);
and U42289 (N_42289,N_37550,N_37563);
xor U42290 (N_42290,N_38409,N_38424);
or U42291 (N_42291,N_38072,N_39811);
nor U42292 (N_42292,N_38460,N_37841);
and U42293 (N_42293,N_39515,N_37882);
and U42294 (N_42294,N_38984,N_39453);
or U42295 (N_42295,N_39067,N_38700);
and U42296 (N_42296,N_39996,N_39866);
nor U42297 (N_42297,N_38912,N_39888);
or U42298 (N_42298,N_39019,N_39956);
or U42299 (N_42299,N_39198,N_37879);
or U42300 (N_42300,N_37743,N_38335);
nand U42301 (N_42301,N_38671,N_38942);
nand U42302 (N_42302,N_38380,N_39564);
and U42303 (N_42303,N_38598,N_39117);
xor U42304 (N_42304,N_39463,N_37960);
nor U42305 (N_42305,N_38403,N_39041);
and U42306 (N_42306,N_39360,N_38054);
nand U42307 (N_42307,N_38928,N_37989);
nor U42308 (N_42308,N_37922,N_38043);
or U42309 (N_42309,N_38698,N_38341);
and U42310 (N_42310,N_38532,N_39080);
xor U42311 (N_42311,N_38844,N_39189);
nor U42312 (N_42312,N_38113,N_37857);
or U42313 (N_42313,N_37893,N_39942);
xnor U42314 (N_42314,N_37831,N_38168);
nor U42315 (N_42315,N_39545,N_38913);
nand U42316 (N_42316,N_39246,N_39219);
nor U42317 (N_42317,N_39466,N_38887);
or U42318 (N_42318,N_38783,N_39476);
and U42319 (N_42319,N_39120,N_38872);
or U42320 (N_42320,N_38197,N_38657);
nand U42321 (N_42321,N_37888,N_37743);
and U42322 (N_42322,N_38665,N_38943);
and U42323 (N_42323,N_38390,N_37653);
or U42324 (N_42324,N_38040,N_38479);
and U42325 (N_42325,N_39077,N_38197);
nor U42326 (N_42326,N_39713,N_38784);
nand U42327 (N_42327,N_38359,N_39499);
and U42328 (N_42328,N_39151,N_37648);
xnor U42329 (N_42329,N_39196,N_39668);
or U42330 (N_42330,N_37638,N_37521);
nor U42331 (N_42331,N_38489,N_38704);
nand U42332 (N_42332,N_38182,N_39048);
and U42333 (N_42333,N_38116,N_39279);
and U42334 (N_42334,N_39819,N_39913);
or U42335 (N_42335,N_39648,N_38984);
nand U42336 (N_42336,N_39383,N_38089);
nand U42337 (N_42337,N_37536,N_37581);
nand U42338 (N_42338,N_39714,N_39973);
nor U42339 (N_42339,N_39516,N_39323);
or U42340 (N_42340,N_38429,N_39422);
xnor U42341 (N_42341,N_38153,N_38674);
or U42342 (N_42342,N_39728,N_38464);
and U42343 (N_42343,N_39258,N_38912);
nand U42344 (N_42344,N_38361,N_38017);
nor U42345 (N_42345,N_38888,N_38591);
or U42346 (N_42346,N_39396,N_39672);
nand U42347 (N_42347,N_38761,N_37532);
xnor U42348 (N_42348,N_38551,N_38839);
and U42349 (N_42349,N_37945,N_39729);
and U42350 (N_42350,N_38846,N_39934);
or U42351 (N_42351,N_37810,N_39960);
nor U42352 (N_42352,N_39463,N_39393);
nand U42353 (N_42353,N_37810,N_38053);
or U42354 (N_42354,N_38585,N_38517);
or U42355 (N_42355,N_38788,N_39099);
and U42356 (N_42356,N_37510,N_38585);
xnor U42357 (N_42357,N_38716,N_38004);
nor U42358 (N_42358,N_39604,N_39482);
xnor U42359 (N_42359,N_38848,N_39162);
xnor U42360 (N_42360,N_37995,N_38023);
and U42361 (N_42361,N_38056,N_39821);
or U42362 (N_42362,N_37798,N_38045);
or U42363 (N_42363,N_39724,N_38812);
nand U42364 (N_42364,N_38411,N_39047);
nor U42365 (N_42365,N_39727,N_38080);
xnor U42366 (N_42366,N_38622,N_39865);
xor U42367 (N_42367,N_39839,N_37957);
and U42368 (N_42368,N_38130,N_37974);
nor U42369 (N_42369,N_38021,N_39361);
nand U42370 (N_42370,N_38771,N_39473);
nand U42371 (N_42371,N_38057,N_39750);
and U42372 (N_42372,N_39406,N_39830);
or U42373 (N_42373,N_38840,N_38216);
nor U42374 (N_42374,N_39370,N_39953);
and U42375 (N_42375,N_38472,N_39276);
nor U42376 (N_42376,N_39035,N_39845);
and U42377 (N_42377,N_39717,N_37742);
nor U42378 (N_42378,N_39751,N_38623);
nor U42379 (N_42379,N_38121,N_38713);
or U42380 (N_42380,N_39370,N_37786);
or U42381 (N_42381,N_37944,N_38865);
xnor U42382 (N_42382,N_38417,N_38211);
xor U42383 (N_42383,N_38953,N_38110);
nand U42384 (N_42384,N_37705,N_39233);
or U42385 (N_42385,N_38447,N_37704);
nor U42386 (N_42386,N_39654,N_39020);
or U42387 (N_42387,N_39684,N_38785);
nor U42388 (N_42388,N_38446,N_39570);
and U42389 (N_42389,N_38716,N_39112);
xor U42390 (N_42390,N_38117,N_38602);
xor U42391 (N_42391,N_37525,N_38376);
and U42392 (N_42392,N_37776,N_38389);
and U42393 (N_42393,N_38565,N_38926);
nand U42394 (N_42394,N_39935,N_38821);
nand U42395 (N_42395,N_39532,N_38682);
xor U42396 (N_42396,N_37569,N_39038);
nand U42397 (N_42397,N_37513,N_38410);
xor U42398 (N_42398,N_39973,N_39309);
nor U42399 (N_42399,N_38826,N_38614);
or U42400 (N_42400,N_38447,N_38135);
and U42401 (N_42401,N_38905,N_39461);
or U42402 (N_42402,N_37890,N_38942);
nor U42403 (N_42403,N_37916,N_38597);
nor U42404 (N_42404,N_37599,N_39398);
or U42405 (N_42405,N_39202,N_38443);
xor U42406 (N_42406,N_39998,N_39900);
or U42407 (N_42407,N_39934,N_39973);
xnor U42408 (N_42408,N_39215,N_39994);
xor U42409 (N_42409,N_39557,N_39987);
nor U42410 (N_42410,N_39953,N_39367);
nand U42411 (N_42411,N_38786,N_38772);
or U42412 (N_42412,N_39401,N_39545);
and U42413 (N_42413,N_38334,N_39661);
nor U42414 (N_42414,N_38678,N_38065);
or U42415 (N_42415,N_38665,N_39473);
or U42416 (N_42416,N_39533,N_39064);
xnor U42417 (N_42417,N_38453,N_38968);
or U42418 (N_42418,N_39480,N_39891);
or U42419 (N_42419,N_39465,N_39099);
nand U42420 (N_42420,N_38396,N_38056);
and U42421 (N_42421,N_39187,N_39485);
or U42422 (N_42422,N_37531,N_37660);
nand U42423 (N_42423,N_39206,N_38861);
or U42424 (N_42424,N_39295,N_39230);
xnor U42425 (N_42425,N_39506,N_39510);
or U42426 (N_42426,N_37640,N_39177);
or U42427 (N_42427,N_38589,N_39207);
or U42428 (N_42428,N_37901,N_37510);
xor U42429 (N_42429,N_37695,N_38679);
nor U42430 (N_42430,N_38129,N_38784);
nor U42431 (N_42431,N_38070,N_39103);
xor U42432 (N_42432,N_37718,N_37681);
or U42433 (N_42433,N_39919,N_38522);
xnor U42434 (N_42434,N_38436,N_38980);
nand U42435 (N_42435,N_39959,N_37582);
nor U42436 (N_42436,N_39621,N_39785);
nor U42437 (N_42437,N_38322,N_39300);
nand U42438 (N_42438,N_39916,N_39305);
nand U42439 (N_42439,N_38476,N_38254);
or U42440 (N_42440,N_38573,N_39261);
nand U42441 (N_42441,N_39224,N_38448);
or U42442 (N_42442,N_38161,N_37880);
xor U42443 (N_42443,N_39239,N_38712);
nand U42444 (N_42444,N_39422,N_37688);
nor U42445 (N_42445,N_39168,N_39463);
or U42446 (N_42446,N_37837,N_37960);
and U42447 (N_42447,N_37531,N_38469);
xor U42448 (N_42448,N_39552,N_39930);
nand U42449 (N_42449,N_38398,N_39560);
or U42450 (N_42450,N_37507,N_38859);
or U42451 (N_42451,N_38030,N_39641);
or U42452 (N_42452,N_38475,N_37841);
xnor U42453 (N_42453,N_38524,N_37954);
and U42454 (N_42454,N_37607,N_39706);
and U42455 (N_42455,N_39215,N_39591);
nor U42456 (N_42456,N_38139,N_38511);
nor U42457 (N_42457,N_37802,N_38616);
nand U42458 (N_42458,N_39189,N_38125);
nor U42459 (N_42459,N_39288,N_39561);
xnor U42460 (N_42460,N_39955,N_38099);
or U42461 (N_42461,N_39486,N_37649);
and U42462 (N_42462,N_37868,N_37975);
or U42463 (N_42463,N_39517,N_38968);
nand U42464 (N_42464,N_38858,N_37688);
or U42465 (N_42465,N_39204,N_39012);
nor U42466 (N_42466,N_39372,N_38866);
nand U42467 (N_42467,N_38159,N_39132);
xor U42468 (N_42468,N_38309,N_38961);
nor U42469 (N_42469,N_39231,N_39257);
and U42470 (N_42470,N_38361,N_37942);
nand U42471 (N_42471,N_37935,N_39216);
nor U42472 (N_42472,N_39238,N_39771);
nor U42473 (N_42473,N_39407,N_39143);
xor U42474 (N_42474,N_39545,N_38613);
nand U42475 (N_42475,N_38382,N_38915);
nand U42476 (N_42476,N_37883,N_39632);
xnor U42477 (N_42477,N_37984,N_37664);
nand U42478 (N_42478,N_39859,N_38622);
and U42479 (N_42479,N_38334,N_37720);
or U42480 (N_42480,N_39270,N_37588);
xor U42481 (N_42481,N_39855,N_39794);
or U42482 (N_42482,N_37612,N_39324);
nor U42483 (N_42483,N_37639,N_38013);
or U42484 (N_42484,N_39789,N_38953);
nor U42485 (N_42485,N_39125,N_38559);
xor U42486 (N_42486,N_39171,N_39497);
or U42487 (N_42487,N_39628,N_39554);
and U42488 (N_42488,N_37727,N_38305);
or U42489 (N_42489,N_37692,N_38975);
nand U42490 (N_42490,N_39649,N_38129);
and U42491 (N_42491,N_39240,N_39751);
nor U42492 (N_42492,N_37869,N_39118);
and U42493 (N_42493,N_39431,N_38702);
nor U42494 (N_42494,N_39005,N_37899);
xnor U42495 (N_42495,N_39082,N_39610);
nor U42496 (N_42496,N_38456,N_39072);
nor U42497 (N_42497,N_38776,N_38164);
nor U42498 (N_42498,N_37972,N_39344);
or U42499 (N_42499,N_38858,N_38943);
and U42500 (N_42500,N_41683,N_41065);
nor U42501 (N_42501,N_41482,N_40993);
nand U42502 (N_42502,N_40854,N_40347);
or U42503 (N_42503,N_40122,N_40775);
or U42504 (N_42504,N_42191,N_41173);
nand U42505 (N_42505,N_42114,N_41381);
or U42506 (N_42506,N_40057,N_42086);
nand U42507 (N_42507,N_41473,N_42117);
or U42508 (N_42508,N_40178,N_40628);
nand U42509 (N_42509,N_41623,N_41704);
nor U42510 (N_42510,N_40911,N_41710);
nand U42511 (N_42511,N_41123,N_40019);
and U42512 (N_42512,N_42095,N_42015);
or U42513 (N_42513,N_41736,N_41273);
or U42514 (N_42514,N_41046,N_42044);
and U42515 (N_42515,N_40507,N_42097);
and U42516 (N_42516,N_40204,N_42367);
nand U42517 (N_42517,N_41648,N_40514);
xnor U42518 (N_42518,N_41245,N_41546);
and U42519 (N_42519,N_41628,N_40888);
nor U42520 (N_42520,N_40815,N_42311);
and U42521 (N_42521,N_41384,N_41706);
and U42522 (N_42522,N_42482,N_41616);
xnor U42523 (N_42523,N_42380,N_41576);
xor U42524 (N_42524,N_41768,N_40327);
nand U42525 (N_42525,N_41760,N_41329);
nor U42526 (N_42526,N_41400,N_40060);
xor U42527 (N_42527,N_41861,N_40937);
nand U42528 (N_42528,N_40211,N_40494);
and U42529 (N_42529,N_41205,N_42271);
xor U42530 (N_42530,N_40038,N_41833);
xor U42531 (N_42531,N_41756,N_40240);
xnor U42532 (N_42532,N_42405,N_40969);
or U42533 (N_42533,N_42013,N_40191);
xor U42534 (N_42534,N_41969,N_41554);
xor U42535 (N_42535,N_41503,N_40672);
nand U42536 (N_42536,N_40984,N_41947);
xnor U42537 (N_42537,N_42357,N_41637);
or U42538 (N_42538,N_40461,N_40980);
and U42539 (N_42539,N_40165,N_41687);
and U42540 (N_42540,N_41881,N_41543);
and U42541 (N_42541,N_40105,N_41578);
nor U42542 (N_42542,N_40011,N_42180);
or U42543 (N_42543,N_40798,N_42153);
nor U42544 (N_42544,N_40340,N_41829);
nor U42545 (N_42545,N_41188,N_40310);
and U42546 (N_42546,N_41621,N_41000);
and U42547 (N_42547,N_40520,N_41220);
or U42548 (N_42548,N_41497,N_40385);
or U42549 (N_42549,N_40661,N_41928);
and U42550 (N_42550,N_41769,N_41338);
nor U42551 (N_42551,N_41654,N_40555);
or U42552 (N_42552,N_41852,N_40214);
nor U42553 (N_42553,N_42495,N_41345);
nor U42554 (N_42554,N_40495,N_40820);
or U42555 (N_42555,N_41206,N_41940);
nor U42556 (N_42556,N_41229,N_41111);
and U42557 (N_42557,N_40997,N_41391);
xnor U42558 (N_42558,N_42433,N_42316);
and U42559 (N_42559,N_41542,N_40311);
xor U42560 (N_42560,N_41530,N_41420);
or U42561 (N_42561,N_42334,N_41717);
xnor U42562 (N_42562,N_40329,N_40182);
xnor U42563 (N_42563,N_41789,N_40654);
xnor U42564 (N_42564,N_41923,N_40999);
xor U42565 (N_42565,N_41147,N_40230);
nand U42566 (N_42566,N_40828,N_41179);
xnor U42567 (N_42567,N_40288,N_40298);
xor U42568 (N_42568,N_42481,N_41269);
nor U42569 (N_42569,N_41252,N_41512);
nand U42570 (N_42570,N_42419,N_40700);
nand U42571 (N_42571,N_41859,N_40504);
xnor U42572 (N_42572,N_41146,N_40111);
xnor U42573 (N_42573,N_40781,N_42445);
xnor U42574 (N_42574,N_41041,N_41332);
nor U42575 (N_42575,N_40768,N_40493);
xor U42576 (N_42576,N_40979,N_41083);
nor U42577 (N_42577,N_42389,N_40481);
nor U42578 (N_42578,N_41939,N_40147);
and U42579 (N_42579,N_42290,N_42270);
and U42580 (N_42580,N_40625,N_41893);
nor U42581 (N_42581,N_41732,N_41262);
nand U42582 (N_42582,N_40838,N_41959);
nand U42583 (N_42583,N_40136,N_42003);
xnor U42584 (N_42584,N_42320,N_40894);
xor U42585 (N_42585,N_41096,N_40610);
xor U42586 (N_42586,N_42338,N_42475);
nor U42587 (N_42587,N_42403,N_40887);
nor U42588 (N_42588,N_41210,N_41130);
xnor U42589 (N_42589,N_42289,N_40062);
nor U42590 (N_42590,N_41692,N_41050);
nand U42591 (N_42591,N_40598,N_42312);
and U42592 (N_42592,N_42148,N_41815);
nand U42593 (N_42593,N_41945,N_41604);
nand U42594 (N_42594,N_42079,N_41990);
and U42595 (N_42595,N_41297,N_41168);
nor U42596 (N_42596,N_40759,N_42450);
nand U42597 (N_42597,N_41448,N_42154);
and U42598 (N_42598,N_41404,N_42129);
and U42599 (N_42599,N_41202,N_40843);
xor U42600 (N_42600,N_42123,N_42084);
nor U42601 (N_42601,N_40280,N_41460);
and U42602 (N_42602,N_40955,N_40730);
nor U42603 (N_42603,N_42023,N_41540);
or U42604 (N_42604,N_40579,N_41259);
and U42605 (N_42605,N_41753,N_40289);
and U42606 (N_42606,N_41326,N_40725);
or U42607 (N_42607,N_40534,N_42062);
or U42608 (N_42608,N_41067,N_41409);
nand U42609 (N_42609,N_41061,N_41645);
nor U42610 (N_42610,N_40553,N_40767);
xnor U42611 (N_42611,N_41548,N_40536);
xnor U42612 (N_42612,N_41248,N_40133);
nand U42613 (N_42613,N_40490,N_41697);
xor U42614 (N_42614,N_41970,N_40891);
nor U42615 (N_42615,N_40852,N_40295);
xor U42616 (N_42616,N_41555,N_41527);
nand U42617 (N_42617,N_40305,N_40751);
and U42618 (N_42618,N_42375,N_41797);
nand U42619 (N_42619,N_40988,N_41099);
nand U42620 (N_42620,N_42304,N_40548);
xor U42621 (N_42621,N_40784,N_40306);
xnor U42622 (N_42622,N_40110,N_41397);
xnor U42623 (N_42623,N_41211,N_41656);
nand U42624 (N_42624,N_40998,N_42147);
nor U42625 (N_42625,N_40965,N_41875);
xor U42626 (N_42626,N_42169,N_42071);
xor U42627 (N_42627,N_42335,N_40934);
nand U42628 (N_42628,N_42344,N_41561);
nor U42629 (N_42629,N_41136,N_40990);
nor U42630 (N_42630,N_40633,N_42234);
xor U42631 (N_42631,N_42022,N_40749);
xnor U42632 (N_42632,N_41462,N_40455);
and U42633 (N_42633,N_40694,N_40102);
nor U42634 (N_42634,N_40512,N_40791);
or U42635 (N_42635,N_42324,N_41754);
nand U42636 (N_42636,N_40713,N_40695);
nand U42637 (N_42637,N_40243,N_42039);
or U42638 (N_42638,N_42001,N_42395);
nor U42639 (N_42639,N_40617,N_42480);
nor U42640 (N_42640,N_41369,N_41268);
or U42641 (N_42641,N_40753,N_41281);
xor U42642 (N_42642,N_40100,N_41086);
xor U42643 (N_42643,N_42272,N_42257);
nor U42644 (N_42644,N_40907,N_41499);
xnor U42645 (N_42645,N_41860,N_40948);
or U42646 (N_42646,N_41325,N_40362);
and U42647 (N_42647,N_42143,N_41403);
or U42648 (N_42648,N_41105,N_42318);
or U42649 (N_42649,N_41031,N_40562);
nor U42650 (N_42650,N_42021,N_41838);
nand U42651 (N_42651,N_40411,N_42315);
and U42652 (N_42652,N_40415,N_40166);
xnor U42653 (N_42653,N_41876,N_42135);
nor U42654 (N_42654,N_41165,N_41480);
nand U42655 (N_42655,N_41337,N_40399);
or U42656 (N_42656,N_41407,N_41713);
nand U42657 (N_42657,N_41545,N_41342);
nor U42658 (N_42658,N_40971,N_42101);
nand U42659 (N_42659,N_40707,N_40012);
nor U42660 (N_42660,N_40052,N_40208);
nand U42661 (N_42661,N_41667,N_41956);
or U42662 (N_42662,N_42359,N_40912);
nor U42663 (N_42663,N_40222,N_40621);
xnor U42664 (N_42664,N_41519,N_42082);
and U42665 (N_42665,N_40279,N_40623);
xnor U42666 (N_42666,N_40373,N_40132);
nor U42667 (N_42667,N_41142,N_40454);
nor U42668 (N_42668,N_40241,N_41303);
nand U42669 (N_42669,N_41095,N_42241);
and U42670 (N_42670,N_40407,N_40920);
and U42671 (N_42671,N_42280,N_40140);
and U42672 (N_42672,N_41238,N_41377);
or U42673 (N_42673,N_42385,N_41314);
and U42674 (N_42674,N_41764,N_41446);
and U42675 (N_42675,N_42141,N_40577);
and U42676 (N_42676,N_42187,N_42461);
nor U42677 (N_42677,N_40307,N_42090);
nor U42678 (N_42678,N_42201,N_40601);
and U42679 (N_42679,N_41263,N_42009);
nor U42680 (N_42680,N_41235,N_41689);
nand U42681 (N_42681,N_42002,N_40390);
nand U42682 (N_42682,N_41176,N_40026);
xnor U42683 (N_42683,N_41057,N_40375);
and U42684 (N_42684,N_41368,N_40073);
and U42685 (N_42685,N_42031,N_41447);
or U42686 (N_42686,N_40153,N_40796);
xnor U42687 (N_42687,N_40232,N_40914);
xnor U42688 (N_42688,N_41960,N_40152);
or U42689 (N_42689,N_41971,N_40200);
xnor U42690 (N_42690,N_40845,N_41445);
nor U42691 (N_42691,N_42200,N_40365);
and U42692 (N_42692,N_41693,N_40799);
or U42693 (N_42693,N_41270,N_40322);
or U42694 (N_42694,N_41359,N_42387);
xnor U42695 (N_42695,N_42378,N_41351);
xnor U42696 (N_42696,N_41916,N_40081);
nor U42697 (N_42697,N_42107,N_42430);
xnor U42698 (N_42698,N_40699,N_40957);
nand U42699 (N_42699,N_42414,N_40650);
or U42700 (N_42700,N_41479,N_42376);
or U42701 (N_42701,N_40639,N_40058);
xnor U42702 (N_42702,N_41662,N_41094);
xnor U42703 (N_42703,N_40299,N_40134);
nand U42704 (N_42704,N_41872,N_40973);
or U42705 (N_42705,N_42469,N_41215);
nand U42706 (N_42706,N_41506,N_42228);
xor U42707 (N_42707,N_42235,N_42371);
or U42708 (N_42708,N_40148,N_41110);
and U42709 (N_42709,N_40393,N_40855);
xor U42710 (N_42710,N_40452,N_41646);
nand U42711 (N_42711,N_41257,N_41842);
and U42712 (N_42712,N_41484,N_40853);
nor U42713 (N_42713,N_42244,N_41567);
nor U42714 (N_42714,N_40413,N_40834);
nor U42715 (N_42715,N_41632,N_40457);
nor U42716 (N_42716,N_41175,N_42415);
nor U42717 (N_42717,N_41373,N_40388);
nor U42718 (N_42718,N_40320,N_40309);
nor U42719 (N_42719,N_41071,N_41085);
xnor U42720 (N_42720,N_41865,N_41596);
or U42721 (N_42721,N_40265,N_40197);
or U42722 (N_42722,N_42401,N_41465);
and U42723 (N_42723,N_40036,N_40430);
nor U42724 (N_42724,N_41247,N_41963);
xor U42725 (N_42725,N_41250,N_40439);
and U42726 (N_42726,N_42010,N_40367);
or U42727 (N_42727,N_42476,N_41158);
nor U42728 (N_42728,N_42293,N_42255);
nor U42729 (N_42729,N_41977,N_41121);
nand U42730 (N_42730,N_42331,N_41798);
or U42731 (N_42731,N_40330,N_42399);
xor U42732 (N_42732,N_40291,N_42472);
nand U42733 (N_42733,N_42170,N_41601);
and U42734 (N_42734,N_41278,N_40629);
or U42735 (N_42735,N_41261,N_41809);
and U42736 (N_42736,N_40488,N_40739);
or U42737 (N_42737,N_40316,N_42448);
nand U42738 (N_42738,N_40981,N_40364);
xnor U42739 (N_42739,N_41836,N_40652);
xnor U42740 (N_42740,N_41812,N_41221);
and U42741 (N_42741,N_41558,N_40789);
and U42742 (N_42742,N_41244,N_40764);
and U42743 (N_42743,N_41669,N_42283);
xor U42744 (N_42744,N_40016,N_41577);
nor U42745 (N_42745,N_42253,N_40875);
nand U42746 (N_42746,N_40007,N_40210);
nor U42747 (N_42747,N_42306,N_41109);
nor U42748 (N_42748,N_42150,N_41063);
nor U42749 (N_42749,N_40380,N_40785);
nand U42750 (N_42750,N_40123,N_40714);
xnor U42751 (N_42751,N_41986,N_41698);
and U42752 (N_42752,N_42033,N_41143);
or U42753 (N_42753,N_40061,N_42372);
or U42754 (N_42754,N_42432,N_41790);
and U42755 (N_42755,N_40422,N_41676);
xnor U42756 (N_42756,N_40423,N_40879);
xor U42757 (N_42757,N_40088,N_41878);
and U42758 (N_42758,N_40028,N_41120);
and U42759 (N_42759,N_41498,N_42174);
xor U42760 (N_42760,N_41395,N_41678);
or U42761 (N_42761,N_41892,N_42250);
xor U42762 (N_42762,N_41197,N_40142);
nor U42763 (N_42763,N_40508,N_41810);
xnor U42764 (N_42764,N_40670,N_42093);
nor U42765 (N_42765,N_41889,N_40389);
nor U42766 (N_42766,N_40287,N_40765);
nand U42767 (N_42767,N_42379,N_41006);
xor U42768 (N_42768,N_41207,N_42172);
nand U42769 (N_42769,N_41964,N_42287);
nand U42770 (N_42770,N_40037,N_41896);
or U42771 (N_42771,N_41438,N_41336);
nor U42772 (N_42772,N_42337,N_42043);
and U42773 (N_42773,N_41408,N_42156);
xnor U42774 (N_42774,N_41231,N_41356);
or U42775 (N_42775,N_40109,N_41767);
xnor U42776 (N_42776,N_41943,N_41440);
nor U42777 (N_42777,N_41284,N_42489);
xnor U42778 (N_42778,N_40126,N_41752);
nor U42779 (N_42779,N_42457,N_41075);
nand U42780 (N_42780,N_41826,N_42055);
xor U42781 (N_42781,N_40303,N_41774);
or U42782 (N_42782,N_42034,N_41433);
and U42783 (N_42783,N_40608,N_41937);
xor U42784 (N_42784,N_41832,N_40410);
and U42785 (N_42785,N_42299,N_40780);
nor U42786 (N_42786,N_41657,N_40545);
nand U42787 (N_42787,N_41242,N_40041);
xnor U42788 (N_42788,N_40432,N_40162);
nor U42789 (N_42789,N_41912,N_41882);
or U42790 (N_42790,N_40726,N_41449);
or U42791 (N_42791,N_42192,N_40817);
nor U42792 (N_42792,N_40778,N_40332);
nand U42793 (N_42793,N_41747,N_41877);
nor U42794 (N_42794,N_41784,N_40866);
nor U42795 (N_42795,N_41023,N_42017);
nor U42796 (N_42796,N_40966,N_40976);
xor U42797 (N_42797,N_40083,N_40368);
nor U42798 (N_42798,N_40511,N_41761);
xnor U42799 (N_42799,N_40090,N_40883);
nor U42800 (N_42800,N_41495,N_41203);
nor U42801 (N_42801,N_42451,N_41899);
and U42802 (N_42802,N_40806,N_40238);
or U42803 (N_42803,N_41988,N_40023);
nor U42804 (N_42804,N_41454,N_40675);
xnor U42805 (N_42805,N_41523,N_42203);
nor U42806 (N_42806,N_40659,N_41642);
and U42807 (N_42807,N_42046,N_40513);
and U42808 (N_42808,N_42407,N_41425);
and U42809 (N_42809,N_41212,N_40733);
nand U42810 (N_42810,N_40589,N_40290);
nor U42811 (N_42811,N_41163,N_41556);
or U42812 (N_42812,N_41995,N_40466);
or U42813 (N_42813,N_41435,N_41254);
nor U42814 (N_42814,N_41625,N_41778);
xnor U42815 (N_42815,N_41936,N_40346);
nand U42816 (N_42816,N_40547,N_40963);
nor U42817 (N_42817,N_40962,N_40906);
xnor U42818 (N_42818,N_40983,N_40760);
xnor U42819 (N_42819,N_41237,N_41196);
nor U42820 (N_42820,N_40405,N_42330);
and U42821 (N_42821,N_42163,N_40395);
nand U42822 (N_42822,N_41106,N_40438);
nor U42823 (N_42823,N_40590,N_42341);
and U42824 (N_42824,N_40952,N_40323);
or U42825 (N_42825,N_42391,N_41974);
xor U42826 (N_42826,N_41217,N_40196);
nor U42827 (N_42827,N_40927,N_41841);
nand U42828 (N_42828,N_42028,N_40130);
nand U42829 (N_42829,N_42158,N_40800);
or U42830 (N_42830,N_40215,N_41192);
nand U42831 (N_42831,N_41816,N_40262);
xnor U42832 (N_42832,N_41658,N_40544);
and U42833 (N_42833,N_41941,N_40812);
nand U42834 (N_42834,N_40762,N_41895);
and U42835 (N_42835,N_40056,N_42356);
and U42836 (N_42836,N_40462,N_40001);
nor U42837 (N_42837,N_40429,N_41887);
and U42838 (N_42838,N_41347,N_42470);
nand U42839 (N_42839,N_41660,N_41280);
and U42840 (N_42840,N_42310,N_40715);
nor U42841 (N_42841,N_40535,N_42377);
or U42842 (N_42842,N_41511,N_40304);
or U42843 (N_42843,N_41087,N_41757);
xor U42844 (N_42844,N_40522,N_41444);
and U42845 (N_42845,N_41239,N_41868);
xnor U42846 (N_42846,N_40478,N_40680);
xor U42847 (N_42847,N_42232,N_41145);
nand U42848 (N_42848,N_40050,N_41898);
xor U42849 (N_42849,N_40257,N_41502);
nor U42850 (N_42850,N_42019,N_40702);
xor U42851 (N_42851,N_40913,N_42237);
and U42852 (N_42852,N_41232,N_41216);
xnor U42853 (N_42853,N_42054,N_42417);
xor U42854 (N_42854,N_40944,N_40634);
nor U42855 (N_42855,N_41230,N_40557);
nor U42856 (N_42856,N_42057,N_40832);
xor U42857 (N_42857,N_42418,N_40592);
nor U42858 (N_42858,N_40626,N_40066);
nand U42859 (N_42859,N_41457,N_40185);
nor U42860 (N_42860,N_40977,N_41283);
nand U42861 (N_42861,N_42113,N_40941);
xnor U42862 (N_42862,N_41913,N_40638);
nand U42863 (N_42863,N_42329,N_40696);
nor U42864 (N_42864,N_41981,N_41372);
nand U42865 (N_42865,N_42268,N_42273);
nand U42866 (N_42866,N_42215,N_41437);
xor U42867 (N_42867,N_42008,N_41223);
and U42868 (N_42868,N_40527,N_40538);
or U42869 (N_42869,N_41552,N_40047);
nor U42870 (N_42870,N_41350,N_40607);
and U42871 (N_42871,N_42134,N_40537);
and U42872 (N_42872,N_40657,N_40925);
nor U42873 (N_42873,N_40246,N_41398);
nor U42874 (N_42874,N_40573,N_41950);
xor U42875 (N_42875,N_40351,N_42218);
nor U42876 (N_42876,N_42394,N_40328);
nand U42877 (N_42877,N_40961,N_41894);
xnor U42878 (N_42878,N_40575,N_40497);
nor U42879 (N_42879,N_40571,N_42178);
nor U42880 (N_42880,N_41113,N_41777);
xor U42881 (N_42881,N_40797,N_42458);
nand U42882 (N_42882,N_42313,N_40063);
nor U42883 (N_42883,N_41557,N_42284);
xnor U42884 (N_42884,N_41021,N_41818);
xor U42885 (N_42885,N_40679,N_41276);
and U42886 (N_42886,N_40744,N_41016);
xor U42887 (N_42887,N_41795,N_41133);
and U42888 (N_42888,N_40158,N_41508);
or U42889 (N_42889,N_41888,N_41516);
xor U42890 (N_42890,N_40811,N_40192);
nor U42891 (N_42891,N_40974,N_42004);
nor U42892 (N_42892,N_41354,N_41227);
or U42893 (N_42893,N_42225,N_41831);
nand U42894 (N_42894,N_41129,N_40294);
xor U42895 (N_42895,N_41027,N_40989);
nand U42896 (N_42896,N_40315,N_40342);
xor U42897 (N_42897,N_41097,N_41549);
xor U42898 (N_42898,N_40250,N_41521);
and U42899 (N_42899,N_41458,N_41694);
xor U42900 (N_42900,N_40712,N_41811);
xnor U42901 (N_42901,N_41529,N_41024);
or U42902 (N_42902,N_40688,N_41627);
or U42903 (N_42903,N_41439,N_40156);
nand U42904 (N_42904,N_40361,N_41471);
or U42905 (N_42905,N_40729,N_41664);
or U42906 (N_42906,N_40383,N_41929);
and U42907 (N_42907,N_40027,N_42285);
xnor U42908 (N_42908,N_41671,N_41200);
nor U42909 (N_42909,N_40479,N_42467);
xor U42910 (N_42910,N_42242,N_41456);
and U42911 (N_42911,N_42102,N_42085);
nand U42912 (N_42912,N_40483,N_41699);
xor U42913 (N_42913,N_40096,N_41243);
nand U42914 (N_42914,N_41101,N_41663);
xnor U42915 (N_42915,N_41029,N_41980);
nor U42916 (N_42916,N_41686,N_42142);
or U42917 (N_42917,N_42453,N_42171);
and U42918 (N_42918,N_42295,N_42104);
nor U42919 (N_42919,N_42259,N_41272);
nand U42920 (N_42920,N_41429,N_40566);
nor U42921 (N_42921,N_40521,N_40354);
or U42922 (N_42922,N_40698,N_40878);
or U42923 (N_42923,N_42067,N_41808);
xor U42924 (N_42924,N_41012,N_40543);
nand U42925 (N_42925,N_40526,N_41640);
nand U42926 (N_42926,N_40515,N_41025);
and U42927 (N_42927,N_40737,N_40379);
or U42928 (N_42928,N_42221,N_41084);
and U42929 (N_42929,N_41393,N_42230);
nor U42930 (N_42930,N_41718,N_41819);
xor U42931 (N_42931,N_42196,N_41468);
nand U42932 (N_42932,N_41910,N_41682);
or U42933 (N_42933,N_42224,N_42473);
or U42934 (N_42934,N_41450,N_41386);
nand U42935 (N_42935,N_40896,N_42262);
nor U42936 (N_42936,N_40837,N_41639);
nor U42937 (N_42937,N_40484,N_40793);
nor U42938 (N_42938,N_40568,N_42421);
or U42939 (N_42939,N_42006,N_40456);
and U42940 (N_42940,N_41022,N_40480);
or U42941 (N_42941,N_42231,N_40564);
nand U42942 (N_42942,N_41124,N_40370);
nand U42943 (N_42943,N_42011,N_41998);
and U42944 (N_42944,N_41489,N_40890);
nand U42945 (N_42945,N_40363,N_42269);
or U42946 (N_42946,N_41226,N_41944);
or U42947 (N_42947,N_40750,N_42452);
and U42948 (N_42948,N_40421,N_40256);
and U42949 (N_42949,N_40772,N_42278);
xnor U42950 (N_42950,N_40569,N_41715);
nor U42951 (N_42951,N_40779,N_41152);
and U42952 (N_42952,N_41128,N_41643);
nand U42953 (N_42953,N_42328,N_41481);
nor U42954 (N_42954,N_40155,N_41528);
nor U42955 (N_42955,N_40756,N_41201);
and U42956 (N_42956,N_41040,N_42443);
nand U42957 (N_42957,N_41043,N_42396);
or U42958 (N_42958,N_41122,N_40164);
and U42959 (N_42959,N_41559,N_40708);
or U42960 (N_42960,N_40095,N_42037);
xor U42961 (N_42961,N_40685,N_41432);
and U42962 (N_42962,N_40741,N_41349);
and U42963 (N_42963,N_41026,N_41365);
and U42964 (N_42964,N_40312,N_40195);
xor U42965 (N_42965,N_40369,N_41864);
and U42966 (N_42966,N_41423,N_42056);
xnor U42967 (N_42967,N_40078,N_40663);
nand U42968 (N_42968,N_40489,N_41731);
nand U42969 (N_42969,N_41580,N_40336);
xor U42970 (N_42970,N_41922,N_40867);
xnor U42971 (N_42971,N_41994,N_41750);
nand U42972 (N_42972,N_42199,N_42223);
nor U42973 (N_42973,N_40987,N_41474);
xor U42974 (N_42974,N_41299,N_40868);
and U42975 (N_42975,N_40417,N_41003);
nor U42976 (N_42976,N_40317,N_40337);
xor U42977 (N_42977,N_40692,N_40844);
nor U42978 (N_42978,N_40051,N_40094);
nor U42979 (N_42979,N_40030,N_42211);
and U42980 (N_42980,N_41786,N_40902);
or U42981 (N_42981,N_40851,N_42176);
and U42982 (N_42982,N_41626,N_40273);
or U42983 (N_42983,N_42348,N_41763);
and U42984 (N_42984,N_40683,N_40145);
nand U42985 (N_42985,N_41737,N_42427);
nor U42986 (N_42986,N_42247,N_41817);
xnor U42987 (N_42987,N_41488,N_41734);
nor U42988 (N_42988,N_42133,N_40179);
nor U42989 (N_42989,N_41078,N_42413);
nor U42990 (N_42990,N_41148,N_40795);
xnor U42991 (N_42991,N_41983,N_40735);
and U42992 (N_42992,N_42209,N_41848);
and U42993 (N_42993,N_40467,N_40873);
nand U42994 (N_42994,N_40384,N_40938);
or U42995 (N_42995,N_41799,N_42149);
or U42996 (N_42996,N_41695,N_40862);
nand U42997 (N_42997,N_42089,N_40400);
or U42998 (N_42998,N_42333,N_42096);
nor U42999 (N_42999,N_40602,N_41491);
and U43000 (N_43000,N_40381,N_41606);
nand U43001 (N_43001,N_40401,N_40967);
nand U43002 (N_43002,N_40341,N_40643);
nor U43003 (N_43003,N_41185,N_40766);
nor U43004 (N_43004,N_41266,N_40181);
nor U43005 (N_43005,N_41634,N_40339);
nand U43006 (N_43006,N_41614,N_41010);
nor U43007 (N_43007,N_41030,N_41037);
nand U43008 (N_43008,N_41472,N_40163);
nor U43009 (N_43009,N_40711,N_41008);
or U43010 (N_43010,N_41144,N_40161);
and U43011 (N_43011,N_40135,N_41126);
xor U43012 (N_43012,N_41953,N_41092);
nor U43013 (N_43013,N_40414,N_40946);
nor U43014 (N_43014,N_42291,N_40580);
and U43015 (N_43015,N_41909,N_41991);
nor U43016 (N_43016,N_42429,N_40217);
and U43017 (N_43017,N_41840,N_41137);
nor U43018 (N_43018,N_41153,N_42412);
xnor U43019 (N_43019,N_40464,N_42303);
xnor U43020 (N_43020,N_40187,N_41487);
nand U43021 (N_43021,N_41758,N_42179);
and U43022 (N_43022,N_42352,N_40325);
nor U43023 (N_43023,N_40949,N_41775);
nand U43024 (N_43024,N_41670,N_41166);
or U43025 (N_43025,N_41182,N_41090);
xor U43026 (N_43026,N_42297,N_40173);
xnor U43027 (N_43027,N_41644,N_41032);
or U43028 (N_43028,N_40404,N_40371);
or U43029 (N_43029,N_42436,N_41076);
xor U43030 (N_43030,N_40045,N_42298);
or U43031 (N_43031,N_40213,N_41360);
nor U43032 (N_43032,N_41004,N_41992);
xor U43033 (N_43033,N_42390,N_41015);
or U43034 (N_43034,N_40801,N_42210);
or U43035 (N_43035,N_40486,N_41089);
or U43036 (N_43036,N_41691,N_42275);
nor U43037 (N_43037,N_40529,N_40492);
or U43038 (N_43038,N_40567,N_41586);
and U43039 (N_43039,N_42212,N_40003);
nand U43040 (N_43040,N_42321,N_41961);
nand U43041 (N_43041,N_41906,N_41535);
xor U43042 (N_43042,N_40253,N_40752);
xor U43043 (N_43043,N_40706,N_40180);
nor U43044 (N_43044,N_41107,N_41419);
xnor U43045 (N_43045,N_40098,N_40002);
nor U43046 (N_43046,N_40443,N_41828);
xnor U43047 (N_43047,N_42070,N_42491);
nor U43048 (N_43048,N_40103,N_42047);
or U43049 (N_43049,N_40374,N_41531);
and U43050 (N_43050,N_41002,N_41466);
and U43051 (N_43051,N_41830,N_41599);
and U43052 (N_43052,N_42248,N_41613);
or U43053 (N_43053,N_40885,N_40546);
or U43054 (N_43054,N_40176,N_41233);
nor U43055 (N_43055,N_41127,N_41264);
or U43056 (N_43056,N_41571,N_40070);
xor U43057 (N_43057,N_40043,N_41886);
xor U43058 (N_43058,N_41515,N_42319);
nor U43059 (N_43059,N_40823,N_41453);
nand U43060 (N_43060,N_41659,N_40473);
nor U43061 (N_43061,N_40787,N_40360);
xor U43062 (N_43062,N_40556,N_41292);
or U43063 (N_43063,N_41289,N_41335);
xor U43064 (N_43064,N_41260,N_40703);
nand U43065 (N_43065,N_40034,N_41967);
and U43066 (N_43066,N_42222,N_40236);
xor U43067 (N_43067,N_42393,N_40006);
nand U43068 (N_43068,N_40604,N_41837);
and U43069 (N_43069,N_40910,N_41340);
nand U43070 (N_43070,N_42300,N_41514);
xor U43071 (N_43071,N_41405,N_40463);
or U43072 (N_43072,N_42444,N_42381);
and U43073 (N_43073,N_40681,N_41406);
or U43074 (N_43074,N_40588,N_41155);
xnor U43075 (N_43075,N_41392,N_42459);
nor U43076 (N_43076,N_40472,N_40732);
or U43077 (N_43077,N_40677,N_41170);
or U43078 (N_43078,N_41486,N_40704);
nand U43079 (N_43079,N_40578,N_42137);
xnor U43080 (N_43080,N_41620,N_41609);
or U43081 (N_43081,N_40860,N_40528);
or U43082 (N_43082,N_40506,N_40510);
nor U43083 (N_43083,N_40582,N_40500);
and U43084 (N_43084,N_42465,N_42309);
nor U43085 (N_43085,N_40260,N_41672);
and U43086 (N_43086,N_42392,N_41091);
and U43087 (N_43087,N_41186,N_40964);
nor U43088 (N_43088,N_41411,N_41884);
nor U43089 (N_43089,N_41702,N_40586);
nor U43090 (N_43090,N_40710,N_41866);
nor U43091 (N_43091,N_40449,N_41009);
xor U43092 (N_43092,N_42165,N_40835);
or U43093 (N_43093,N_41743,N_40237);
and U43094 (N_43094,N_40942,N_42214);
nand U43095 (N_43095,N_40943,N_40451);
or U43096 (N_43096,N_41582,N_40228);
xnor U43097 (N_43097,N_40445,N_40611);
or U43098 (N_43098,N_40458,N_41319);
or U43099 (N_43099,N_42435,N_41249);
or U43100 (N_43100,N_40029,N_41323);
or U43101 (N_43101,N_41275,N_41701);
nor U43102 (N_43102,N_40667,N_40183);
xnor U43103 (N_43103,N_42488,N_41017);
nor U43104 (N_43104,N_41900,N_40761);
xnor U43105 (N_43105,N_40223,N_41313);
xor U43106 (N_43106,N_42014,N_41803);
xor U43107 (N_43107,N_40723,N_41394);
xnor U43108 (N_43108,N_40446,N_41572);
and U43109 (N_43109,N_40338,N_40570);
xnor U43110 (N_43110,N_41160,N_40477);
or U43111 (N_43111,N_41375,N_41112);
nor U43112 (N_43112,N_41328,N_41905);
nand U43113 (N_43113,N_42484,N_40014);
nor U43114 (N_43114,N_42496,N_40086);
xnor U43115 (N_43115,N_41020,N_42189);
nand U43116 (N_43116,N_41534,N_41401);
nor U43117 (N_43117,N_40666,N_40242);
nor U43118 (N_43118,N_40382,N_40859);
and U43119 (N_43119,N_41417,N_41058);
or U43120 (N_43120,N_41001,N_40075);
nor U43121 (N_43121,N_42139,N_41619);
and U43122 (N_43122,N_42400,N_41927);
or U43123 (N_43123,N_41564,N_41463);
xnor U43124 (N_43124,N_40705,N_41282);
and U43125 (N_43125,N_41383,N_40300);
nand U43126 (N_43126,N_42087,N_40498);
or U43127 (N_43127,N_40372,N_41723);
and U43128 (N_43128,N_42111,N_42077);
or U43129 (N_43129,N_41539,N_41854);
nand U43130 (N_43130,N_40149,N_41933);
xor U43131 (N_43131,N_42064,N_41595);
and U43132 (N_43132,N_42190,N_41361);
and U43133 (N_43133,N_40450,N_42460);
nor U43134 (N_43134,N_41302,N_40641);
and U43135 (N_43135,N_41705,N_41611);
nor U43136 (N_43136,N_40847,N_42308);
nor U43137 (N_43137,N_40819,N_40656);
xnor U43138 (N_43138,N_42110,N_40199);
and U43139 (N_43139,N_41052,N_40565);
nor U43140 (N_43140,N_40727,N_40931);
nor U43141 (N_43141,N_40172,N_42182);
nor U43142 (N_43142,N_41926,N_41862);
and U43143 (N_43143,N_41873,N_40841);
and U43144 (N_43144,N_40539,N_40560);
or U43145 (N_43145,N_42264,N_42208);
nor U43146 (N_43146,N_41055,N_42140);
nor U43147 (N_43147,N_40335,N_42487);
or U43148 (N_43148,N_41733,N_41675);
xor U43149 (N_43149,N_41312,N_40101);
xor U43150 (N_43150,N_40089,N_40491);
and U43151 (N_43151,N_42265,N_41984);
or U43152 (N_43152,N_42184,N_41191);
nor U43153 (N_43153,N_41513,N_41858);
nand U43154 (N_43154,N_41441,N_40595);
and U43155 (N_43155,N_41745,N_42125);
and U43156 (N_43156,N_41762,N_41602);
nand U43157 (N_43157,N_41426,N_41573);
nor U43158 (N_43158,N_40392,N_40758);
and U43159 (N_43159,N_40924,N_40377);
and U43160 (N_43160,N_41844,N_40922);
nand U43161 (N_43161,N_41324,N_41309);
nand U43162 (N_43162,N_42105,N_40889);
or U43163 (N_43163,N_42065,N_40021);
nand U43164 (N_43164,N_41805,N_41685);
or U43165 (N_43165,N_40674,N_42346);
nor U43166 (N_43166,N_41712,N_42474);
or U43167 (N_43167,N_41485,N_41119);
or U43168 (N_43168,N_42027,N_40496);
xnor U43169 (N_43169,N_40755,N_42155);
xor U43170 (N_43170,N_41436,N_40171);
nor U43171 (N_43171,N_42288,N_41719);
and U43172 (N_43172,N_40420,N_42076);
nand U43173 (N_43173,N_40916,N_40426);
nand U43174 (N_43174,N_41477,N_42198);
nand U43175 (N_43175,N_41277,N_40552);
nor U43176 (N_43176,N_41307,N_40297);
nand U43177 (N_43177,N_40821,N_42339);
or U43178 (N_43178,N_42167,N_40635);
nand U43179 (N_43179,N_41355,N_40783);
and U43180 (N_43180,N_40814,N_40397);
and U43181 (N_43181,N_41857,N_41431);
and U43182 (N_43182,N_41414,N_42121);
nor U43183 (N_43183,N_42325,N_41034);
or U43184 (N_43184,N_42454,N_41794);
or U43185 (N_43185,N_41924,N_41251);
and U43186 (N_43186,N_40402,N_40160);
nand U43187 (N_43187,N_40459,N_40084);
and U43188 (N_43188,N_40015,N_41846);
nor U43189 (N_43189,N_41584,N_40594);
and U43190 (N_43190,N_40055,N_40720);
and U43191 (N_43191,N_40198,N_40637);
or U43192 (N_43192,N_40008,N_40099);
nand U43193 (N_43193,N_41298,N_42462);
nor U43194 (N_43194,N_40807,N_41853);
nand U43195 (N_43195,N_40684,N_41709);
nor U43196 (N_43196,N_41585,N_40433);
xor U43197 (N_43197,N_42332,N_41934);
and U43198 (N_43198,N_41070,N_42063);
and U43199 (N_43199,N_41346,N_41399);
nor U43200 (N_43200,N_41824,N_41274);
or U43201 (N_43201,N_41104,N_41741);
and U43202 (N_43202,N_41989,N_40849);
or U43203 (N_43203,N_41213,N_41164);
and U43204 (N_43204,N_41589,N_40782);
or U43205 (N_43205,N_40035,N_41932);
xor U43206 (N_43206,N_41744,N_40319);
nor U43207 (N_43207,N_40137,N_40991);
nor U43208 (N_43208,N_40292,N_42059);
nand U43209 (N_43209,N_40067,N_41366);
and U43210 (N_43210,N_40928,N_40040);
nor U43211 (N_43211,N_41501,N_41072);
nor U43212 (N_43212,N_40763,N_41547);
or U43213 (N_43213,N_40940,N_40091);
nand U43214 (N_43214,N_41115,N_40718);
nand U43215 (N_43215,N_41455,N_41100);
or U43216 (N_43216,N_41652,N_41150);
nand U43217 (N_43217,N_41389,N_40738);
nor U43218 (N_43218,N_41677,N_40412);
nor U43219 (N_43219,N_41975,N_40865);
nor U43220 (N_43220,N_41966,N_40082);
and U43221 (N_43221,N_42026,N_41553);
xor U43222 (N_43222,N_40271,N_41079);
or U43223 (N_43223,N_40809,N_41305);
or U43224 (N_43224,N_41522,N_40274);
xor U43225 (N_43225,N_41766,N_41721);
nor U43226 (N_43226,N_41726,N_40146);
or U43227 (N_43227,N_41132,N_40031);
nand U43228 (N_43228,N_41885,N_41167);
nand U43229 (N_43229,N_40453,N_41951);
nand U43230 (N_43230,N_40115,N_40394);
nor U43231 (N_43231,N_42226,N_40518);
xnor U43232 (N_43232,N_41972,N_40825);
xnor U43233 (N_43233,N_40398,N_42052);
nor U43234 (N_43234,N_41331,N_41633);
or U43235 (N_43235,N_40950,N_41517);
or U43236 (N_43236,N_42422,N_40836);
xor U43237 (N_43237,N_42124,N_41066);
xnor U43238 (N_43238,N_41294,N_41271);
nand U43239 (N_43239,N_40596,N_40930);
nand U43240 (N_43240,N_41018,N_40632);
and U43241 (N_43241,N_41199,N_41593);
and U43242 (N_43242,N_40519,N_41493);
nand U43243 (N_43243,N_40112,N_42490);
nor U43244 (N_43244,N_41402,N_40403);
xor U43245 (N_43245,N_41304,N_41285);
nand U43246 (N_43246,N_40048,N_41949);
xor U43247 (N_43247,N_41749,N_42267);
and U43248 (N_43248,N_40216,N_40188);
xor U43249 (N_43249,N_41382,N_40205);
nand U43250 (N_43250,N_42197,N_40827);
nand U43251 (N_43251,N_40523,N_42406);
nand U43252 (N_43252,N_41773,N_40349);
nor U43253 (N_43253,N_40059,N_40428);
xnor U43254 (N_43254,N_40959,N_41341);
xor U43255 (N_43255,N_41219,N_42471);
xor U43256 (N_43256,N_40193,N_40808);
or U43257 (N_43257,N_40754,N_40282);
and U43258 (N_43258,N_40956,N_40691);
and U43259 (N_43259,N_41204,N_42263);
nor U43260 (N_43260,N_40583,N_42109);
nand U43261 (N_43261,N_40716,N_42088);
or U43262 (N_43262,N_40118,N_40326);
and U43263 (N_43263,N_41180,N_42112);
and U43264 (N_43264,N_41938,N_42108);
or U43265 (N_43265,N_40686,N_40255);
nand U43266 (N_43266,N_42162,N_42426);
xnor U43267 (N_43267,N_40378,N_40788);
or U43268 (N_43268,N_42347,N_42195);
and U43269 (N_43269,N_41724,N_42388);
or U43270 (N_43270,N_40301,N_40167);
and U43271 (N_43271,N_42068,N_42206);
xnor U43272 (N_43272,N_40097,N_42048);
nand U43273 (N_43273,N_41570,N_41874);
nand U43274 (N_43274,N_40505,N_40640);
nand U43275 (N_43275,N_40144,N_41730);
nand U43276 (N_43276,N_42479,N_42302);
or U43277 (N_43277,N_42301,N_41357);
and U43278 (N_43278,N_41315,N_41069);
nor U43279 (N_43279,N_41310,N_40074);
and U43280 (N_43280,N_40169,N_42369);
and U43281 (N_43281,N_40709,N_40846);
xor U43282 (N_43282,N_42383,N_42249);
and U43283 (N_43283,N_41184,N_40476);
and U43284 (N_43284,N_40939,N_40017);
or U43285 (N_43285,N_41880,N_41174);
nor U43286 (N_43286,N_41739,N_42254);
xnor U43287 (N_43287,N_40921,N_42098);
nand U43288 (N_43288,N_40069,N_42317);
xnor U43289 (N_43289,N_41897,N_42365);
xnor U43290 (N_43290,N_42246,N_40436);
or U43291 (N_43291,N_40120,N_40995);
nor U43292 (N_43292,N_40668,N_41839);
nor U43293 (N_43293,N_41288,N_41635);
and U43294 (N_43294,N_41793,N_41081);
nand U43295 (N_43295,N_41827,N_40561);
nor U43296 (N_43296,N_41019,N_40313);
nor U43297 (N_43297,N_40502,N_40882);
xnor U43298 (N_43298,N_41256,N_41422);
nand U43299 (N_43299,N_41293,N_40947);
and U43300 (N_43300,N_40013,N_41234);
xnor U43301 (N_43301,N_40184,N_41563);
and U43302 (N_43302,N_40742,N_41209);
or U43303 (N_43303,N_42029,N_40917);
nor U43304 (N_43304,N_41668,N_41851);
and U43305 (N_43305,N_40869,N_42100);
or U43306 (N_43306,N_42292,N_40143);
and U43307 (N_43307,N_41987,N_42074);
nor U43308 (N_43308,N_42217,N_41843);
xnor U43309 (N_43309,N_42281,N_41946);
and U43310 (N_43310,N_42138,N_41116);
nor U43311 (N_43311,N_41255,N_40064);
xnor U43312 (N_43312,N_41380,N_40644);
and U43313 (N_43313,N_40106,N_40227);
and U43314 (N_43314,N_40159,N_40892);
nand U43315 (N_43315,N_41653,N_40524);
or U43316 (N_43316,N_41510,N_40877);
xor U43317 (N_43317,N_40252,N_40427);
or U43318 (N_43318,N_41679,N_41590);
xnor U43319 (N_43319,N_40308,N_41045);
xor U43320 (N_43320,N_41782,N_41729);
nor U43321 (N_43321,N_40968,N_42477);
nand U43322 (N_43322,N_41246,N_42349);
or U43323 (N_43323,N_41600,N_42276);
nand U43324 (N_43324,N_41655,N_41821);
nor U43325 (N_43325,N_40880,N_41236);
xor U43326 (N_43326,N_40270,N_41157);
and U43327 (N_43327,N_41690,N_40032);
or U43328 (N_43328,N_42194,N_41222);
and U43329 (N_43329,N_41028,N_42073);
xor U43330 (N_43330,N_42404,N_40444);
nand U43331 (N_43331,N_41461,N_40509);
nor U43332 (N_43332,N_40777,N_41982);
or U43333 (N_43333,N_41014,N_40079);
nand U43334 (N_43334,N_41225,N_42229);
nand U43335 (N_43335,N_40863,N_41565);
xor U43336 (N_43336,N_40175,N_41048);
nand U43337 (N_43337,N_41013,N_40826);
nor U43338 (N_43338,N_42066,N_40186);
or U43339 (N_43339,N_42350,N_41287);
or U43340 (N_43340,N_42428,N_41791);
and U43341 (N_43341,N_42038,N_42193);
or U43342 (N_43342,N_41612,N_42493);
and U43343 (N_43343,N_41708,N_42366);
or U43344 (N_43344,N_40978,N_42025);
or U43345 (N_43345,N_41060,N_40648);
and U43346 (N_43346,N_41728,N_42075);
and U43347 (N_43347,N_42363,N_40813);
nand U43348 (N_43348,N_42120,N_40350);
nor U43349 (N_43349,N_41711,N_41804);
nor U43350 (N_43350,N_40150,N_42202);
nor U43351 (N_43351,N_40333,N_42439);
nor U43352 (N_43352,N_42463,N_42420);
and U43353 (N_43353,N_40448,N_40239);
xnor U43354 (N_43354,N_41042,N_41993);
nor U43355 (N_43355,N_40769,N_40334);
nor U43356 (N_43356,N_41666,N_42083);
and U43357 (N_43357,N_41908,N_42146);
nand U43358 (N_43358,N_41781,N_41371);
and U43359 (N_43359,N_40833,N_40951);
xnor U43360 (N_43360,N_42416,N_41636);
and U43361 (N_43361,N_40551,N_41550);
and U43362 (N_43362,N_41178,N_41624);
nand U43363 (N_43363,N_40285,N_42127);
nand U43364 (N_43364,N_40658,N_40776);
nand U43365 (N_43365,N_40503,N_40487);
xnor U43366 (N_43366,N_40664,N_41615);
and U43367 (N_43367,N_41978,N_41883);
and U43368 (N_43368,N_41807,N_41258);
nand U43369 (N_43369,N_40039,N_40416);
nand U43370 (N_43370,N_40612,N_41295);
nand U43371 (N_43371,N_40249,N_41492);
and U43372 (N_43372,N_42173,N_40816);
nor U43373 (N_43373,N_42384,N_40202);
and U43374 (N_43374,N_42440,N_42456);
nor U43375 (N_43375,N_40009,N_41538);
and U43376 (N_43376,N_40220,N_40970);
nand U43377 (N_43377,N_40904,N_40550);
or U43378 (N_43378,N_40318,N_41536);
nand U43379 (N_43379,N_41088,N_40599);
nor U43380 (N_43380,N_41387,N_42130);
and U43381 (N_43381,N_41920,N_41996);
nand U43382 (N_43382,N_42012,N_42449);
and U43383 (N_43383,N_40276,N_41241);
or U43384 (N_43384,N_41759,N_40647);
nand U43385 (N_43385,N_40665,N_40154);
xor U43386 (N_43386,N_40909,N_40620);
nor U43387 (N_43387,N_40170,N_40630);
nand U43388 (N_43388,N_40722,N_40409);
nand U43389 (N_43389,N_42364,N_42342);
xnor U43390 (N_43390,N_41334,N_41451);
nor U43391 (N_43391,N_41997,N_42188);
or U43392 (N_43392,N_42423,N_40033);
nand U43393 (N_43393,N_40724,N_41193);
nor U43394 (N_43394,N_42382,N_42455);
xor U43395 (N_43395,N_40022,N_41494);
and U43396 (N_43396,N_41470,N_40572);
or U43397 (N_43397,N_40331,N_40324);
and U43398 (N_43398,N_41507,N_40121);
or U43399 (N_43399,N_40359,N_40655);
or U43400 (N_43400,N_41569,N_40391);
xnor U43401 (N_43401,N_41751,N_40020);
and U43402 (N_43402,N_40631,N_41544);
or U43403 (N_43403,N_40856,N_40746);
or U43404 (N_43404,N_41035,N_42499);
nand U43405 (N_43405,N_42438,N_41587);
nor U43406 (N_43406,N_40923,N_42468);
xnor U43407 (N_43407,N_40992,N_41748);
xnor U43408 (N_43408,N_41267,N_41149);
and U43409 (N_43409,N_41973,N_41080);
nor U43410 (N_43410,N_40771,N_41452);
nor U43411 (N_43411,N_40424,N_40076);
and U43412 (N_43412,N_42164,N_42351);
and U43413 (N_43413,N_41965,N_41651);
nand U43414 (N_43414,N_40994,N_40251);
or U43415 (N_43415,N_40616,N_41151);
nand U43416 (N_43416,N_41958,N_42398);
and U43417 (N_43417,N_41903,N_42069);
nor U43418 (N_43418,N_40786,N_41189);
nand U43419 (N_43419,N_40004,N_40201);
or U43420 (N_43420,N_41442,N_41957);
or U43421 (N_43421,N_42408,N_41140);
and U43422 (N_43422,N_42327,N_41847);
xnor U43423 (N_43423,N_41802,N_40804);
or U43424 (N_43424,N_40141,N_40221);
nand U43425 (N_43425,N_40231,N_41610);
nor U43426 (N_43426,N_40745,N_41746);
or U43427 (N_43427,N_41725,N_41478);
nand U43428 (N_43428,N_41835,N_41177);
or U43429 (N_43429,N_41064,N_40408);
xnor U43430 (N_43430,N_41190,N_40901);
nand U43431 (N_43431,N_41138,N_41575);
and U43432 (N_43432,N_40918,N_42119);
nor U43433 (N_43433,N_41183,N_41198);
or U43434 (N_43434,N_40366,N_42016);
xnor U43435 (N_43435,N_41631,N_41044);
nor U43436 (N_43436,N_42358,N_42437);
nand U43437 (N_43437,N_40794,N_40441);
and U43438 (N_43438,N_40072,N_42260);
nand U43439 (N_43439,N_40116,N_42402);
nor U43440 (N_43440,N_41722,N_41629);
or U43441 (N_43441,N_41367,N_41007);
nor U43442 (N_43442,N_40018,N_40606);
nor U43443 (N_43443,N_42126,N_41421);
or U43444 (N_43444,N_41476,N_41598);
nor U43445 (N_43445,N_41300,N_41714);
nor U43446 (N_43446,N_41532,N_41039);
and U43447 (N_43447,N_41703,N_42081);
or U43448 (N_43448,N_41684,N_41551);
nand U43449 (N_43449,N_40618,N_41378);
nor U43450 (N_43450,N_42411,N_41504);
and U43451 (N_43451,N_41822,N_41286);
xor U43452 (N_43452,N_40267,N_42060);
nor U43453 (N_43453,N_42336,N_41240);
xor U43454 (N_43454,N_41496,N_42061);
nor U43455 (N_43455,N_42266,N_40108);
nand U43456 (N_43456,N_41942,N_40554);
and U43457 (N_43457,N_42294,N_41688);
or U43458 (N_43458,N_42494,N_41459);
xnor U43459 (N_43459,N_42447,N_40049);
nor U43460 (N_43460,N_40669,N_42258);
xnor U43461 (N_43461,N_41776,N_40884);
or U43462 (N_43462,N_42478,N_40605);
nand U43463 (N_43463,N_41161,N_40905);
xor U43464 (N_43464,N_40437,N_40071);
nor U43465 (N_43465,N_40396,N_40986);
nor U43466 (N_43466,N_42106,N_41214);
nand U43467 (N_43467,N_40757,N_41291);
and U43468 (N_43468,N_40645,N_42080);
nand U43469 (N_43469,N_41603,N_40302);
nand U43470 (N_43470,N_41318,N_40721);
nand U43471 (N_43471,N_42261,N_41930);
nor U43472 (N_43472,N_40864,N_42092);
nor U43473 (N_43473,N_41135,N_41779);
and U43474 (N_43474,N_40954,N_41074);
nand U43475 (N_43475,N_42296,N_40803);
nor U43476 (N_43476,N_40541,N_40919);
nor U43477 (N_43477,N_41118,N_41385);
and U43478 (N_43478,N_42118,N_40591);
xnor U43479 (N_43479,N_41162,N_41696);
nand U43480 (N_43480,N_40000,N_41647);
nor U43481 (N_43481,N_40434,N_42256);
nand U43482 (N_43482,N_41597,N_40139);
nor U43483 (N_43483,N_42166,N_41131);
nor U43484 (N_43484,N_40321,N_41410);
or U43485 (N_43485,N_41605,N_40356);
nand U43486 (N_43486,N_41279,N_42245);
or U43487 (N_43487,N_41879,N_41738);
nor U43488 (N_43488,N_40474,N_41813);
and U43489 (N_43489,N_40435,N_40660);
nor U43490 (N_43490,N_41665,N_42103);
and U43491 (N_43491,N_40870,N_40259);
or U43492 (N_43492,N_40649,N_40603);
nor U43493 (N_43493,N_41475,N_42282);
or U43494 (N_43494,N_41056,N_42497);
nand U43495 (N_43495,N_40124,N_40127);
or U43496 (N_43496,N_40247,N_41500);
or U43497 (N_43497,N_40770,N_41891);
and U43498 (N_43498,N_41870,N_41364);
nand U43499 (N_43499,N_41082,N_42145);
or U43500 (N_43500,N_41914,N_42370);
nand U43501 (N_43501,N_42041,N_40138);
xor U43502 (N_43502,N_40719,N_40194);
xor U43503 (N_43503,N_41890,N_40662);
xnor U43504 (N_43504,N_40174,N_42049);
xor U43505 (N_43505,N_40281,N_41483);
and U43506 (N_43506,N_41526,N_42091);
and U43507 (N_43507,N_41755,N_41820);
or U43508 (N_43508,N_42116,N_41154);
or U43509 (N_43509,N_41490,N_40234);
nand U43510 (N_43510,N_40876,N_42252);
nand U43511 (N_43511,N_41467,N_40525);
nor U43512 (N_43512,N_41867,N_42035);
or U43513 (N_43513,N_41265,N_40829);
nor U43514 (N_43514,N_41443,N_41509);
or U43515 (N_43515,N_40226,N_42175);
or U43516 (N_43516,N_40516,N_42131);
nor U43517 (N_43517,N_41469,N_42409);
xnor U43518 (N_43518,N_40673,N_40810);
nor U43519 (N_43519,N_40831,N_42486);
xor U43520 (N_43520,N_40734,N_40499);
or U43521 (N_43521,N_41428,N_40805);
and U43522 (N_43522,N_41228,N_41796);
xor U43523 (N_43523,N_41921,N_42136);
and U43524 (N_43524,N_41871,N_40418);
and U43525 (N_43525,N_41901,N_41608);
nand U43526 (N_43526,N_40501,N_41792);
or U43527 (N_43527,N_42314,N_41321);
xor U43528 (N_43528,N_42036,N_40858);
and U43529 (N_43529,N_42005,N_40792);
and U43530 (N_43530,N_41505,N_41114);
nand U43531 (N_43531,N_41059,N_41785);
nand U43532 (N_43532,N_40189,N_42307);
or U43533 (N_43533,N_42030,N_42132);
or U43534 (N_43534,N_40345,N_41416);
nand U43535 (N_43535,N_40636,N_40926);
and U43536 (N_43536,N_40482,N_40646);
or U43537 (N_43537,N_40824,N_40277);
nand U43538 (N_43538,N_41850,N_40376);
and U43539 (N_43539,N_42050,N_41093);
and U43540 (N_43540,N_42360,N_42355);
nand U43541 (N_43541,N_42032,N_40286);
or U43542 (N_43542,N_41904,N_40278);
nor U43543 (N_43543,N_41770,N_40830);
nor U43544 (N_43544,N_41322,N_41915);
nor U43545 (N_43545,N_40119,N_42219);
nand U43546 (N_43546,N_40314,N_42483);
or U43547 (N_43547,N_40802,N_40125);
xor U43548 (N_43548,N_41413,N_41208);
and U43549 (N_43549,N_40268,N_41823);
or U43550 (N_43550,N_42115,N_41856);
and U43551 (N_43551,N_40687,N_41054);
nor U43552 (N_43552,N_42397,N_40209);
or U43553 (N_43553,N_40293,N_41783);
xnor U43554 (N_43554,N_42216,N_40935);
nor U43555 (N_43555,N_41053,N_41520);
nand U43556 (N_43556,N_42362,N_41765);
or U43557 (N_43557,N_40077,N_40233);
and U43558 (N_43558,N_41434,N_42425);
nor U43559 (N_43559,N_41716,N_42233);
nand U43560 (N_43560,N_41344,N_41396);
or U43561 (N_43561,N_40682,N_40615);
xor U43562 (N_43562,N_40932,N_42151);
xor U43563 (N_43563,N_42446,N_40468);
nand U43564 (N_43564,N_40893,N_41181);
xor U43565 (N_43565,N_40903,N_42094);
nor U43566 (N_43566,N_40531,N_42373);
nor U43567 (N_43567,N_42251,N_42144);
nor U43568 (N_43568,N_40790,N_40203);
or U43569 (N_43569,N_41661,N_41707);
xnor U43570 (N_43570,N_42040,N_41537);
and U43571 (N_43571,N_40857,N_40225);
nand U43572 (N_43572,N_40355,N_41581);
nand U43573 (N_43573,N_40207,N_41103);
xnor U43574 (N_43574,N_40740,N_41968);
nand U43575 (N_43575,N_40344,N_41907);
nor U43576 (N_43576,N_41700,N_41618);
and U43577 (N_43577,N_42243,N_40206);
nand U43578 (N_43578,N_41412,N_41641);
and U43579 (N_43579,N_40558,N_42441);
or U43580 (N_43580,N_40343,N_42122);
nor U43581 (N_43581,N_41194,N_41301);
xnor U43582 (N_43582,N_42354,N_41296);
and U43583 (N_43583,N_40177,N_41141);
and U43584 (N_43584,N_42239,N_41999);
or U43585 (N_43585,N_40025,N_41952);
xor U43586 (N_43586,N_40190,N_41955);
nor U43587 (N_43587,N_41560,N_40269);
nand U43588 (N_43588,N_40224,N_40542);
and U43589 (N_43589,N_41727,N_40248);
and U43590 (N_43590,N_40653,N_40848);
nor U43591 (N_43591,N_42238,N_40533);
nor U43592 (N_43592,N_40264,N_40085);
nand U43593 (N_43593,N_42205,N_41327);
xor U43594 (N_43594,N_41787,N_41005);
nand U43595 (N_43595,N_40068,N_41525);
nand U43596 (N_43596,N_41985,N_41911);
and U43597 (N_43597,N_40465,N_42053);
or U43598 (N_43598,N_41680,N_40619);
nand U43599 (N_43599,N_41681,N_40353);
nor U43600 (N_43600,N_40731,N_42353);
nor U43601 (N_43601,N_41588,N_42185);
and U43602 (N_43602,N_40850,N_40104);
xor U43603 (N_43603,N_40689,N_42322);
xor U43604 (N_43604,N_40114,N_40107);
xor U43605 (N_43605,N_40895,N_40600);
xnor U43606 (N_43606,N_40460,N_42277);
nand U43607 (N_43607,N_40485,N_40080);
or U43608 (N_43608,N_42078,N_40475);
xnor U43609 (N_43609,N_40743,N_41036);
xnor U43610 (N_43610,N_40839,N_41592);
nand U43611 (N_43611,N_42340,N_40044);
and U43612 (N_43612,N_40609,N_42159);
xor U43613 (N_43613,N_40157,N_41800);
nor U43614 (N_43614,N_40425,N_41772);
or U43615 (N_43615,N_42386,N_42498);
or U43616 (N_43616,N_41845,N_42305);
nor U43617 (N_43617,N_41424,N_41290);
nand U43618 (N_43618,N_42492,N_41801);
and U43619 (N_43619,N_40218,N_41172);
or U43620 (N_43620,N_41187,N_40275);
nand U43621 (N_43621,N_41117,N_41771);
nand U43622 (N_43622,N_41102,N_41622);
nand U43623 (N_43623,N_40593,N_40284);
or U43624 (N_43624,N_41954,N_40736);
and U43625 (N_43625,N_40431,N_40581);
or U43626 (N_43626,N_41673,N_41649);
and U43627 (N_43627,N_40697,N_41047);
xor U43628 (N_43628,N_41541,N_42128);
xnor U43629 (N_43629,N_41917,N_41224);
or U43630 (N_43630,N_40915,N_42045);
xor U43631 (N_43631,N_40559,N_40953);
nand U43632 (N_43632,N_42042,N_41594);
nor U43633 (N_43633,N_41038,N_40549);
nand U43634 (N_43634,N_41348,N_40872);
nor U43635 (N_43635,N_42361,N_40128);
nand U43636 (N_43636,N_41918,N_41849);
nand U43637 (N_43637,N_40348,N_40908);
nand U43638 (N_43638,N_41343,N_40574);
and U43639 (N_43639,N_42431,N_40678);
nand U43640 (N_43640,N_41317,N_42177);
xnor U43641 (N_43641,N_41362,N_41427);
or U43642 (N_43642,N_40219,N_40958);
xnor U43643 (N_43643,N_40933,N_41869);
nor U43644 (N_43644,N_42345,N_40168);
and U43645 (N_43645,N_42161,N_41650);
nand U43646 (N_43646,N_40024,N_41919);
and U43647 (N_43647,N_41415,N_41156);
nor U43648 (N_43648,N_40272,N_40010);
and U43649 (N_43649,N_41430,N_41253);
nand U43650 (N_43650,N_40235,N_42072);
nor U43651 (N_43651,N_41735,N_42186);
nand U43652 (N_43652,N_40587,N_42183);
nor U43653 (N_43653,N_41363,N_41740);
nand U43654 (N_43654,N_41316,N_40283);
nor U43655 (N_43655,N_40897,N_40151);
and U43656 (N_43656,N_41320,N_40540);
xnor U43657 (N_43657,N_41306,N_40818);
nor U43658 (N_43658,N_41814,N_41976);
xor U43659 (N_43659,N_40982,N_41931);
xnor U43660 (N_43660,N_41574,N_41566);
nor U43661 (N_43661,N_42343,N_41033);
nor U43662 (N_43662,N_40245,N_40386);
and U43663 (N_43663,N_41370,N_40929);
xnor U43664 (N_43664,N_41788,N_40773);
nand U43665 (N_43665,N_42220,N_40258);
and U43666 (N_43666,N_42323,N_40087);
and U43667 (N_43667,N_40747,N_42152);
nand U43668 (N_43668,N_41855,N_40092);
xor U43669 (N_43669,N_41674,N_41049);
and U43670 (N_43670,N_40129,N_41617);
nor U43671 (N_43671,N_42099,N_40975);
and U43672 (N_43672,N_40440,N_40899);
xor U43673 (N_43673,N_41011,N_42410);
or U43674 (N_43674,N_42000,N_42279);
nor U43675 (N_43675,N_41825,N_41374);
xor U43676 (N_43676,N_40840,N_40065);
nand U43677 (N_43677,N_42058,N_40945);
nand U43678 (N_43678,N_40701,N_41948);
nor U43679 (N_43679,N_41863,N_41376);
nand U43680 (N_43680,N_40254,N_41579);
and U43681 (N_43681,N_42157,N_40597);
xnor U43682 (N_43682,N_40690,N_42434);
or U43683 (N_43683,N_41902,N_40985);
xnor U43684 (N_43684,N_40584,N_40244);
or U43685 (N_43685,N_42326,N_42160);
nand U43686 (N_43686,N_40419,N_40871);
and U43687 (N_43687,N_42274,N_41125);
and U43688 (N_43688,N_42007,N_40642);
nor U43689 (N_43689,N_41339,N_42168);
or U43690 (N_43690,N_40960,N_40532);
or U43691 (N_43691,N_40671,N_40406);
nor U43692 (N_43692,N_40613,N_40113);
or U43693 (N_43693,N_41568,N_40651);
and U43694 (N_43694,N_40936,N_40996);
and U43695 (N_43695,N_41353,N_42424);
nand U43696 (N_43696,N_42485,N_42204);
xnor U43697 (N_43697,N_41352,N_40774);
xnor U43698 (N_43698,N_40053,N_40676);
and U43699 (N_43699,N_40886,N_40261);
xnor U43700 (N_43700,N_42442,N_42051);
nor U43701 (N_43701,N_41935,N_40717);
nor U43702 (N_43702,N_41134,N_42464);
nor U43703 (N_43703,N_41333,N_41607);
nor U43704 (N_43704,N_40530,N_41742);
nand U43705 (N_43705,N_41979,N_41098);
nor U43706 (N_43706,N_41720,N_40898);
nor U43707 (N_43707,N_41562,N_41533);
nand U43708 (N_43708,N_41638,N_40042);
xor U43709 (N_43709,N_41583,N_41925);
nor U43710 (N_43710,N_40442,N_42236);
nand U43711 (N_43711,N_41780,N_40212);
and U43712 (N_43712,N_40576,N_40046);
and U43713 (N_43713,N_40117,N_42240);
xor U43714 (N_43714,N_40352,N_41062);
xor U43715 (N_43715,N_40131,N_41518);
nor U43716 (N_43716,N_41171,N_41464);
nor U43717 (N_43717,N_42213,N_40054);
nand U43718 (N_43718,N_40471,N_40358);
nor U43719 (N_43719,N_40093,N_42286);
and U43720 (N_43720,N_41308,N_41390);
or U43721 (N_43721,N_40624,N_42368);
and U43722 (N_43722,N_41073,N_41195);
and U43723 (N_43723,N_41591,N_40357);
or U43724 (N_43724,N_42207,N_41806);
or U43725 (N_43725,N_42024,N_40614);
xor U43726 (N_43726,N_41139,N_40387);
xor U43727 (N_43727,N_40822,N_40266);
nand U43728 (N_43728,N_41418,N_40229);
and U43729 (N_43729,N_41834,N_40622);
nor U43730 (N_43730,N_40972,N_40881);
nand U43731 (N_43731,N_40861,N_42020);
xor U43732 (N_43732,N_42374,N_41108);
xor U43733 (N_43733,N_40842,N_41630);
or U43734 (N_43734,N_42018,N_40263);
nor U43735 (N_43735,N_42466,N_41169);
nor U43736 (N_43736,N_41388,N_41962);
nand U43737 (N_43737,N_40005,N_40585);
and U43738 (N_43738,N_41159,N_40563);
nand U43739 (N_43739,N_41379,N_41311);
and U43740 (N_43740,N_40900,N_42227);
or U43741 (N_43741,N_40517,N_42181);
or U43742 (N_43742,N_40748,N_41218);
xnor U43743 (N_43743,N_40728,N_40469);
or U43744 (N_43744,N_41330,N_41068);
nor U43745 (N_43745,N_41524,N_40693);
and U43746 (N_43746,N_40470,N_41051);
xor U43747 (N_43747,N_41077,N_40874);
or U43748 (N_43748,N_40627,N_41358);
xor U43749 (N_43749,N_40447,N_40296);
nor U43750 (N_43750,N_41410,N_41102);
and U43751 (N_43751,N_41739,N_42260);
xnor U43752 (N_43752,N_41206,N_40159);
xor U43753 (N_43753,N_42275,N_42188);
nand U43754 (N_43754,N_42024,N_40370);
xor U43755 (N_43755,N_42470,N_40074);
and U43756 (N_43756,N_41699,N_41752);
or U43757 (N_43757,N_40536,N_41764);
xor U43758 (N_43758,N_41249,N_42153);
and U43759 (N_43759,N_40782,N_40182);
nand U43760 (N_43760,N_42415,N_41879);
nor U43761 (N_43761,N_40565,N_40905);
xor U43762 (N_43762,N_40093,N_41922);
or U43763 (N_43763,N_41248,N_40264);
and U43764 (N_43764,N_40251,N_41564);
xor U43765 (N_43765,N_40970,N_41736);
xor U43766 (N_43766,N_40383,N_42391);
xor U43767 (N_43767,N_40176,N_40215);
xnor U43768 (N_43768,N_42126,N_41809);
xnor U43769 (N_43769,N_41877,N_41718);
xor U43770 (N_43770,N_40490,N_40612);
nand U43771 (N_43771,N_40348,N_41688);
nor U43772 (N_43772,N_40435,N_40599);
nand U43773 (N_43773,N_42019,N_41505);
xnor U43774 (N_43774,N_40511,N_40886);
nand U43775 (N_43775,N_40677,N_42374);
xnor U43776 (N_43776,N_42463,N_40736);
and U43777 (N_43777,N_41237,N_41944);
xnor U43778 (N_43778,N_40835,N_41390);
nand U43779 (N_43779,N_42123,N_42232);
xnor U43780 (N_43780,N_42236,N_40350);
or U43781 (N_43781,N_40527,N_42015);
nand U43782 (N_43782,N_42114,N_42081);
xnor U43783 (N_43783,N_40979,N_42459);
nand U43784 (N_43784,N_41945,N_40853);
nor U43785 (N_43785,N_41873,N_40783);
nor U43786 (N_43786,N_42069,N_41468);
xnor U43787 (N_43787,N_40391,N_40965);
nand U43788 (N_43788,N_40428,N_41350);
nand U43789 (N_43789,N_40052,N_41610);
nand U43790 (N_43790,N_41198,N_40961);
nor U43791 (N_43791,N_40983,N_40417);
or U43792 (N_43792,N_40884,N_41043);
nand U43793 (N_43793,N_40462,N_40110);
nand U43794 (N_43794,N_41718,N_40107);
xor U43795 (N_43795,N_42001,N_40190);
nor U43796 (N_43796,N_41042,N_42374);
or U43797 (N_43797,N_40567,N_41949);
nor U43798 (N_43798,N_40700,N_41051);
and U43799 (N_43799,N_42065,N_41809);
and U43800 (N_43800,N_40224,N_41214);
nor U43801 (N_43801,N_41576,N_40750);
and U43802 (N_43802,N_41466,N_41913);
or U43803 (N_43803,N_40060,N_42356);
or U43804 (N_43804,N_42053,N_40301);
or U43805 (N_43805,N_41993,N_42219);
xnor U43806 (N_43806,N_40466,N_40524);
and U43807 (N_43807,N_41925,N_40754);
xnor U43808 (N_43808,N_41631,N_42303);
xnor U43809 (N_43809,N_41373,N_41896);
and U43810 (N_43810,N_41778,N_41539);
or U43811 (N_43811,N_40858,N_40483);
xor U43812 (N_43812,N_41965,N_41180);
nand U43813 (N_43813,N_40441,N_41459);
nor U43814 (N_43814,N_41464,N_41095);
nand U43815 (N_43815,N_41108,N_41153);
or U43816 (N_43816,N_42024,N_40406);
and U43817 (N_43817,N_42455,N_40136);
nor U43818 (N_43818,N_40491,N_42291);
xnor U43819 (N_43819,N_41221,N_40812);
or U43820 (N_43820,N_42103,N_41555);
nand U43821 (N_43821,N_41176,N_40891);
nand U43822 (N_43822,N_40277,N_40440);
or U43823 (N_43823,N_41056,N_40332);
and U43824 (N_43824,N_40826,N_42057);
nand U43825 (N_43825,N_41705,N_40258);
xor U43826 (N_43826,N_41363,N_40591);
nand U43827 (N_43827,N_41559,N_41191);
and U43828 (N_43828,N_42432,N_41988);
or U43829 (N_43829,N_41962,N_42181);
nor U43830 (N_43830,N_41338,N_41027);
nand U43831 (N_43831,N_42057,N_40560);
and U43832 (N_43832,N_40927,N_40341);
nand U43833 (N_43833,N_41245,N_40482);
nand U43834 (N_43834,N_40060,N_40878);
xor U43835 (N_43835,N_41282,N_41097);
or U43836 (N_43836,N_41054,N_40825);
or U43837 (N_43837,N_40252,N_41850);
and U43838 (N_43838,N_41402,N_40595);
or U43839 (N_43839,N_40961,N_42133);
nand U43840 (N_43840,N_41900,N_41854);
nand U43841 (N_43841,N_41907,N_42117);
xnor U43842 (N_43842,N_41231,N_41427);
xnor U43843 (N_43843,N_40405,N_41875);
nor U43844 (N_43844,N_40352,N_41874);
nand U43845 (N_43845,N_41864,N_40149);
and U43846 (N_43846,N_40011,N_41783);
or U43847 (N_43847,N_41045,N_40706);
and U43848 (N_43848,N_40304,N_41457);
or U43849 (N_43849,N_41372,N_41472);
nor U43850 (N_43850,N_40030,N_41696);
nor U43851 (N_43851,N_41537,N_40250);
or U43852 (N_43852,N_40221,N_40620);
nand U43853 (N_43853,N_41834,N_40876);
xor U43854 (N_43854,N_40090,N_40745);
nor U43855 (N_43855,N_40134,N_41134);
nand U43856 (N_43856,N_40965,N_41536);
or U43857 (N_43857,N_42274,N_40077);
or U43858 (N_43858,N_41674,N_42377);
and U43859 (N_43859,N_40887,N_41299);
nand U43860 (N_43860,N_41824,N_40371);
nand U43861 (N_43861,N_41162,N_40621);
and U43862 (N_43862,N_41340,N_42238);
xnor U43863 (N_43863,N_40137,N_42349);
nand U43864 (N_43864,N_40726,N_41935);
or U43865 (N_43865,N_40839,N_40107);
xnor U43866 (N_43866,N_42346,N_40984);
xnor U43867 (N_43867,N_41357,N_41972);
or U43868 (N_43868,N_40328,N_41147);
and U43869 (N_43869,N_41126,N_40179);
xnor U43870 (N_43870,N_41557,N_42499);
nand U43871 (N_43871,N_40789,N_40346);
nor U43872 (N_43872,N_40683,N_41051);
nand U43873 (N_43873,N_41349,N_40118);
or U43874 (N_43874,N_41459,N_41958);
nand U43875 (N_43875,N_40804,N_41221);
xor U43876 (N_43876,N_41433,N_41950);
nor U43877 (N_43877,N_41038,N_42418);
and U43878 (N_43878,N_41097,N_40163);
nor U43879 (N_43879,N_41123,N_41727);
and U43880 (N_43880,N_41085,N_40520);
nand U43881 (N_43881,N_41116,N_40322);
nor U43882 (N_43882,N_41527,N_40081);
nand U43883 (N_43883,N_40920,N_41588);
or U43884 (N_43884,N_42042,N_42291);
and U43885 (N_43885,N_41313,N_41098);
nor U43886 (N_43886,N_41174,N_42121);
nand U43887 (N_43887,N_41518,N_41086);
or U43888 (N_43888,N_42160,N_40307);
nand U43889 (N_43889,N_41099,N_40504);
nand U43890 (N_43890,N_40125,N_40441);
or U43891 (N_43891,N_40563,N_41727);
or U43892 (N_43892,N_40688,N_42267);
and U43893 (N_43893,N_40776,N_40928);
nor U43894 (N_43894,N_41934,N_40467);
and U43895 (N_43895,N_41926,N_40572);
xnor U43896 (N_43896,N_41196,N_40459);
xnor U43897 (N_43897,N_41966,N_42082);
nor U43898 (N_43898,N_40163,N_42427);
or U43899 (N_43899,N_42374,N_40411);
nand U43900 (N_43900,N_40975,N_41969);
nor U43901 (N_43901,N_40580,N_41629);
and U43902 (N_43902,N_40297,N_40429);
xor U43903 (N_43903,N_40869,N_42433);
nand U43904 (N_43904,N_42479,N_40044);
nor U43905 (N_43905,N_41595,N_41169);
nor U43906 (N_43906,N_40444,N_40996);
or U43907 (N_43907,N_41538,N_40240);
xor U43908 (N_43908,N_40737,N_41611);
nand U43909 (N_43909,N_40694,N_42066);
nor U43910 (N_43910,N_41634,N_40093);
or U43911 (N_43911,N_41532,N_41695);
or U43912 (N_43912,N_42026,N_41943);
nor U43913 (N_43913,N_42077,N_40513);
nor U43914 (N_43914,N_42286,N_42401);
nand U43915 (N_43915,N_41669,N_42380);
nand U43916 (N_43916,N_41304,N_41519);
nor U43917 (N_43917,N_41293,N_40582);
nand U43918 (N_43918,N_41308,N_42240);
nor U43919 (N_43919,N_42330,N_42376);
xor U43920 (N_43920,N_41630,N_41842);
xor U43921 (N_43921,N_40966,N_40520);
xor U43922 (N_43922,N_40551,N_40916);
nand U43923 (N_43923,N_41559,N_40145);
xnor U43924 (N_43924,N_42158,N_41024);
xor U43925 (N_43925,N_41630,N_42328);
nor U43926 (N_43926,N_42227,N_40568);
nor U43927 (N_43927,N_41557,N_41313);
and U43928 (N_43928,N_40070,N_42481);
nor U43929 (N_43929,N_40962,N_41853);
xnor U43930 (N_43930,N_42208,N_42016);
nor U43931 (N_43931,N_41101,N_41777);
and U43932 (N_43932,N_41025,N_40152);
nand U43933 (N_43933,N_40246,N_40842);
nor U43934 (N_43934,N_41670,N_40702);
nand U43935 (N_43935,N_41887,N_40905);
xor U43936 (N_43936,N_42325,N_41320);
nand U43937 (N_43937,N_40627,N_41950);
nand U43938 (N_43938,N_41108,N_42236);
xor U43939 (N_43939,N_42288,N_42309);
xor U43940 (N_43940,N_41400,N_40023);
nand U43941 (N_43941,N_42045,N_41718);
or U43942 (N_43942,N_40258,N_41560);
and U43943 (N_43943,N_40036,N_40824);
and U43944 (N_43944,N_41593,N_41227);
xnor U43945 (N_43945,N_40986,N_40256);
nand U43946 (N_43946,N_41018,N_40509);
nor U43947 (N_43947,N_41781,N_41773);
or U43948 (N_43948,N_40865,N_40577);
nand U43949 (N_43949,N_40856,N_41884);
and U43950 (N_43950,N_40113,N_41117);
xor U43951 (N_43951,N_42242,N_40260);
xor U43952 (N_43952,N_40691,N_42078);
and U43953 (N_43953,N_42365,N_40261);
and U43954 (N_43954,N_40644,N_41279);
or U43955 (N_43955,N_41461,N_40589);
nor U43956 (N_43956,N_41081,N_41562);
and U43957 (N_43957,N_40891,N_42252);
xnor U43958 (N_43958,N_42231,N_41971);
and U43959 (N_43959,N_42281,N_40878);
nand U43960 (N_43960,N_40845,N_42016);
nand U43961 (N_43961,N_42422,N_41703);
and U43962 (N_43962,N_41652,N_41772);
and U43963 (N_43963,N_41458,N_41127);
xor U43964 (N_43964,N_40378,N_40416);
xor U43965 (N_43965,N_40696,N_41689);
nand U43966 (N_43966,N_42391,N_40746);
nand U43967 (N_43967,N_40257,N_41850);
xnor U43968 (N_43968,N_41971,N_40202);
xor U43969 (N_43969,N_41435,N_40113);
and U43970 (N_43970,N_40701,N_40015);
nand U43971 (N_43971,N_41965,N_42277);
and U43972 (N_43972,N_41771,N_41690);
xor U43973 (N_43973,N_41433,N_41855);
nor U43974 (N_43974,N_40738,N_40707);
xor U43975 (N_43975,N_42015,N_40666);
xnor U43976 (N_43976,N_41946,N_42280);
xnor U43977 (N_43977,N_42128,N_42121);
and U43978 (N_43978,N_41330,N_42497);
nor U43979 (N_43979,N_41518,N_41163);
nor U43980 (N_43980,N_41506,N_42353);
nand U43981 (N_43981,N_41451,N_41259);
xnor U43982 (N_43982,N_42314,N_40778);
or U43983 (N_43983,N_42260,N_40078);
nor U43984 (N_43984,N_40106,N_41906);
nand U43985 (N_43985,N_41099,N_40883);
or U43986 (N_43986,N_42026,N_41052);
nand U43987 (N_43987,N_40176,N_41871);
and U43988 (N_43988,N_42137,N_41429);
xor U43989 (N_43989,N_42169,N_41829);
nand U43990 (N_43990,N_42358,N_42392);
nand U43991 (N_43991,N_41275,N_41058);
xnor U43992 (N_43992,N_41865,N_41167);
nand U43993 (N_43993,N_41504,N_40281);
xor U43994 (N_43994,N_40979,N_41089);
and U43995 (N_43995,N_41291,N_40298);
and U43996 (N_43996,N_42213,N_41623);
xnor U43997 (N_43997,N_41771,N_40863);
nor U43998 (N_43998,N_40425,N_40951);
and U43999 (N_43999,N_40167,N_41766);
xnor U44000 (N_44000,N_40553,N_42025);
nor U44001 (N_44001,N_41991,N_41805);
and U44002 (N_44002,N_41024,N_42000);
nor U44003 (N_44003,N_40851,N_41598);
nor U44004 (N_44004,N_41874,N_40131);
nand U44005 (N_44005,N_42226,N_40823);
or U44006 (N_44006,N_41368,N_41033);
or U44007 (N_44007,N_42344,N_41881);
and U44008 (N_44008,N_42032,N_40739);
nor U44009 (N_44009,N_40789,N_40278);
and U44010 (N_44010,N_41352,N_40341);
xnor U44011 (N_44011,N_40931,N_42350);
xor U44012 (N_44012,N_41249,N_40244);
nand U44013 (N_44013,N_42028,N_41946);
xnor U44014 (N_44014,N_40484,N_41601);
and U44015 (N_44015,N_41125,N_40240);
nand U44016 (N_44016,N_42105,N_42150);
xor U44017 (N_44017,N_41307,N_42427);
nand U44018 (N_44018,N_40734,N_41419);
nand U44019 (N_44019,N_40547,N_42078);
xor U44020 (N_44020,N_40857,N_40172);
xnor U44021 (N_44021,N_40679,N_42499);
or U44022 (N_44022,N_41168,N_41058);
nand U44023 (N_44023,N_41564,N_42039);
nand U44024 (N_44024,N_41843,N_40056);
nand U44025 (N_44025,N_41793,N_40734);
or U44026 (N_44026,N_41936,N_42446);
xor U44027 (N_44027,N_41067,N_40103);
nor U44028 (N_44028,N_41711,N_40821);
nand U44029 (N_44029,N_40208,N_40228);
or U44030 (N_44030,N_41863,N_41238);
or U44031 (N_44031,N_40079,N_41651);
xor U44032 (N_44032,N_42176,N_41374);
nor U44033 (N_44033,N_41531,N_41388);
nand U44034 (N_44034,N_40948,N_40352);
or U44035 (N_44035,N_41992,N_40633);
nand U44036 (N_44036,N_41468,N_40549);
nand U44037 (N_44037,N_41111,N_40231);
xnor U44038 (N_44038,N_40341,N_40904);
nor U44039 (N_44039,N_41440,N_42112);
and U44040 (N_44040,N_40790,N_40244);
nand U44041 (N_44041,N_41238,N_41418);
xnor U44042 (N_44042,N_42188,N_41476);
nand U44043 (N_44043,N_40873,N_41076);
or U44044 (N_44044,N_40245,N_41268);
or U44045 (N_44045,N_40292,N_41701);
xnor U44046 (N_44046,N_41730,N_40242);
nor U44047 (N_44047,N_40431,N_42348);
nor U44048 (N_44048,N_40566,N_41403);
nand U44049 (N_44049,N_40034,N_42333);
xor U44050 (N_44050,N_40599,N_40794);
nor U44051 (N_44051,N_42046,N_40944);
nor U44052 (N_44052,N_42063,N_41653);
nand U44053 (N_44053,N_40551,N_41808);
or U44054 (N_44054,N_42282,N_41429);
nand U44055 (N_44055,N_41962,N_41720);
xnor U44056 (N_44056,N_42493,N_41076);
and U44057 (N_44057,N_41282,N_42134);
xor U44058 (N_44058,N_40131,N_40542);
xnor U44059 (N_44059,N_41816,N_40969);
or U44060 (N_44060,N_41799,N_41444);
nand U44061 (N_44061,N_42050,N_41411);
xnor U44062 (N_44062,N_40588,N_40517);
and U44063 (N_44063,N_41253,N_40912);
and U44064 (N_44064,N_41185,N_41772);
and U44065 (N_44065,N_41911,N_42104);
nand U44066 (N_44066,N_40279,N_42308);
nor U44067 (N_44067,N_40286,N_40198);
or U44068 (N_44068,N_42269,N_40555);
or U44069 (N_44069,N_42400,N_40684);
nor U44070 (N_44070,N_40262,N_42004);
xnor U44071 (N_44071,N_40925,N_42287);
nand U44072 (N_44072,N_41541,N_40469);
xnor U44073 (N_44073,N_40941,N_41807);
nor U44074 (N_44074,N_41617,N_41023);
nand U44075 (N_44075,N_42020,N_40531);
nor U44076 (N_44076,N_40034,N_41871);
and U44077 (N_44077,N_42347,N_41439);
or U44078 (N_44078,N_41510,N_42442);
xnor U44079 (N_44079,N_40437,N_40993);
and U44080 (N_44080,N_42191,N_41967);
and U44081 (N_44081,N_42432,N_41397);
or U44082 (N_44082,N_40601,N_42411);
xor U44083 (N_44083,N_41107,N_40457);
nand U44084 (N_44084,N_40539,N_40745);
and U44085 (N_44085,N_41466,N_40453);
or U44086 (N_44086,N_41380,N_40823);
or U44087 (N_44087,N_40373,N_40268);
xor U44088 (N_44088,N_40384,N_40901);
and U44089 (N_44089,N_41551,N_40192);
xor U44090 (N_44090,N_42272,N_41988);
or U44091 (N_44091,N_40850,N_40563);
xnor U44092 (N_44092,N_42074,N_41463);
or U44093 (N_44093,N_41125,N_42006);
nor U44094 (N_44094,N_40383,N_42487);
nor U44095 (N_44095,N_41210,N_41828);
xor U44096 (N_44096,N_41904,N_40126);
nor U44097 (N_44097,N_40715,N_40600);
nor U44098 (N_44098,N_41489,N_42054);
nor U44099 (N_44099,N_40750,N_40387);
nand U44100 (N_44100,N_40431,N_41793);
and U44101 (N_44101,N_42051,N_41817);
nor U44102 (N_44102,N_41164,N_40673);
or U44103 (N_44103,N_41851,N_42070);
xor U44104 (N_44104,N_41609,N_41901);
and U44105 (N_44105,N_40292,N_40715);
nand U44106 (N_44106,N_40645,N_42383);
nor U44107 (N_44107,N_41272,N_40539);
and U44108 (N_44108,N_42187,N_42258);
nor U44109 (N_44109,N_42007,N_40783);
or U44110 (N_44110,N_40310,N_40200);
or U44111 (N_44111,N_41293,N_40340);
or U44112 (N_44112,N_41366,N_40184);
nand U44113 (N_44113,N_42103,N_40057);
xor U44114 (N_44114,N_41604,N_40216);
xnor U44115 (N_44115,N_41687,N_42114);
nor U44116 (N_44116,N_41797,N_42233);
or U44117 (N_44117,N_40915,N_40717);
nor U44118 (N_44118,N_41282,N_40782);
and U44119 (N_44119,N_42304,N_41481);
and U44120 (N_44120,N_42328,N_41132);
nand U44121 (N_44121,N_42057,N_41738);
nand U44122 (N_44122,N_41403,N_41203);
nor U44123 (N_44123,N_40033,N_41241);
and U44124 (N_44124,N_41522,N_40496);
and U44125 (N_44125,N_41691,N_41193);
and U44126 (N_44126,N_41908,N_40528);
xnor U44127 (N_44127,N_40367,N_41502);
nor U44128 (N_44128,N_40773,N_41592);
or U44129 (N_44129,N_41875,N_40469);
xnor U44130 (N_44130,N_41513,N_42030);
and U44131 (N_44131,N_41236,N_40846);
nand U44132 (N_44132,N_41165,N_41179);
xor U44133 (N_44133,N_42019,N_40273);
nor U44134 (N_44134,N_40579,N_41639);
and U44135 (N_44135,N_40048,N_42195);
nor U44136 (N_44136,N_40821,N_41894);
and U44137 (N_44137,N_40398,N_42325);
nand U44138 (N_44138,N_40488,N_40789);
and U44139 (N_44139,N_42191,N_40312);
nand U44140 (N_44140,N_40864,N_40681);
nor U44141 (N_44141,N_40430,N_41515);
and U44142 (N_44142,N_42057,N_41332);
xnor U44143 (N_44143,N_41343,N_40125);
nor U44144 (N_44144,N_40757,N_41501);
xor U44145 (N_44145,N_40258,N_40721);
nand U44146 (N_44146,N_41805,N_41970);
or U44147 (N_44147,N_40013,N_40756);
nand U44148 (N_44148,N_41222,N_41846);
or U44149 (N_44149,N_41212,N_40024);
or U44150 (N_44150,N_40615,N_40092);
or U44151 (N_44151,N_41705,N_40699);
and U44152 (N_44152,N_40895,N_42136);
nand U44153 (N_44153,N_40300,N_42202);
and U44154 (N_44154,N_41872,N_40196);
xnor U44155 (N_44155,N_42146,N_41385);
nand U44156 (N_44156,N_41788,N_40793);
xnor U44157 (N_44157,N_40108,N_41139);
nor U44158 (N_44158,N_40552,N_41240);
and U44159 (N_44159,N_41660,N_41831);
xnor U44160 (N_44160,N_41786,N_40366);
or U44161 (N_44161,N_41828,N_41780);
nand U44162 (N_44162,N_41500,N_41562);
nand U44163 (N_44163,N_40542,N_41997);
or U44164 (N_44164,N_41379,N_40833);
nor U44165 (N_44165,N_41388,N_40419);
nand U44166 (N_44166,N_40531,N_41869);
nor U44167 (N_44167,N_40801,N_40301);
nand U44168 (N_44168,N_41176,N_40655);
or U44169 (N_44169,N_40581,N_40401);
xor U44170 (N_44170,N_41226,N_42140);
or U44171 (N_44171,N_40566,N_41141);
and U44172 (N_44172,N_40026,N_40307);
and U44173 (N_44173,N_40248,N_41698);
xor U44174 (N_44174,N_41887,N_40993);
nor U44175 (N_44175,N_40478,N_40239);
xnor U44176 (N_44176,N_40252,N_40230);
or U44177 (N_44177,N_41810,N_40104);
or U44178 (N_44178,N_42173,N_41168);
and U44179 (N_44179,N_42033,N_40873);
xor U44180 (N_44180,N_40956,N_40166);
or U44181 (N_44181,N_41327,N_41960);
nor U44182 (N_44182,N_40585,N_40137);
xnor U44183 (N_44183,N_41194,N_40026);
nor U44184 (N_44184,N_41773,N_40221);
nor U44185 (N_44185,N_40185,N_40495);
nor U44186 (N_44186,N_40134,N_40711);
or U44187 (N_44187,N_40539,N_41293);
nor U44188 (N_44188,N_40391,N_42051);
or U44189 (N_44189,N_40450,N_40694);
or U44190 (N_44190,N_40668,N_40828);
xnor U44191 (N_44191,N_42382,N_40661);
or U44192 (N_44192,N_40915,N_40932);
and U44193 (N_44193,N_40859,N_41205);
nand U44194 (N_44194,N_41961,N_41898);
or U44195 (N_44195,N_40526,N_42117);
nand U44196 (N_44196,N_40189,N_40566);
xnor U44197 (N_44197,N_41829,N_40855);
nor U44198 (N_44198,N_41702,N_40990);
and U44199 (N_44199,N_41301,N_40582);
nand U44200 (N_44200,N_42231,N_40975);
nor U44201 (N_44201,N_40961,N_40031);
xnor U44202 (N_44202,N_41315,N_42024);
nor U44203 (N_44203,N_41995,N_41405);
nand U44204 (N_44204,N_40297,N_41572);
nand U44205 (N_44205,N_40616,N_41894);
nor U44206 (N_44206,N_41848,N_40860);
or U44207 (N_44207,N_41221,N_40382);
xnor U44208 (N_44208,N_40203,N_40154);
and U44209 (N_44209,N_41841,N_41721);
nor U44210 (N_44210,N_42468,N_41839);
xor U44211 (N_44211,N_40783,N_41169);
and U44212 (N_44212,N_40044,N_41687);
or U44213 (N_44213,N_40553,N_40897);
or U44214 (N_44214,N_40551,N_40734);
nor U44215 (N_44215,N_41693,N_42449);
xor U44216 (N_44216,N_41888,N_42400);
nor U44217 (N_44217,N_40595,N_41022);
nor U44218 (N_44218,N_41689,N_41064);
nor U44219 (N_44219,N_41218,N_40907);
nand U44220 (N_44220,N_40219,N_40648);
nor U44221 (N_44221,N_42276,N_40591);
nand U44222 (N_44222,N_41194,N_40801);
or U44223 (N_44223,N_40624,N_40749);
or U44224 (N_44224,N_40933,N_41532);
nand U44225 (N_44225,N_41545,N_40666);
and U44226 (N_44226,N_41733,N_40581);
and U44227 (N_44227,N_40728,N_42110);
and U44228 (N_44228,N_40753,N_41033);
nand U44229 (N_44229,N_40991,N_41682);
xnor U44230 (N_44230,N_42185,N_41079);
nor U44231 (N_44231,N_40739,N_41102);
nand U44232 (N_44232,N_42379,N_40404);
or U44233 (N_44233,N_41270,N_40419);
xor U44234 (N_44234,N_41351,N_40523);
or U44235 (N_44235,N_40650,N_40852);
nor U44236 (N_44236,N_41933,N_42221);
and U44237 (N_44237,N_41747,N_40340);
nor U44238 (N_44238,N_40913,N_41740);
and U44239 (N_44239,N_42309,N_41217);
nand U44240 (N_44240,N_40468,N_42459);
or U44241 (N_44241,N_41763,N_41634);
and U44242 (N_44242,N_41265,N_42492);
xnor U44243 (N_44243,N_41179,N_41878);
nor U44244 (N_44244,N_42120,N_42225);
and U44245 (N_44245,N_40214,N_41896);
nor U44246 (N_44246,N_42158,N_40332);
xnor U44247 (N_44247,N_42469,N_40223);
or U44248 (N_44248,N_40625,N_41969);
nor U44249 (N_44249,N_40382,N_40391);
or U44250 (N_44250,N_40915,N_41107);
xor U44251 (N_44251,N_41015,N_40317);
and U44252 (N_44252,N_41124,N_41944);
and U44253 (N_44253,N_41569,N_41536);
or U44254 (N_44254,N_42108,N_41834);
and U44255 (N_44255,N_42354,N_40244);
nand U44256 (N_44256,N_41202,N_40163);
or U44257 (N_44257,N_40894,N_41333);
nor U44258 (N_44258,N_41546,N_40058);
nor U44259 (N_44259,N_42229,N_41134);
or U44260 (N_44260,N_40915,N_40255);
or U44261 (N_44261,N_41634,N_42267);
and U44262 (N_44262,N_42318,N_41612);
xnor U44263 (N_44263,N_40562,N_40657);
nand U44264 (N_44264,N_41560,N_41421);
and U44265 (N_44265,N_41714,N_40856);
nand U44266 (N_44266,N_41196,N_41463);
or U44267 (N_44267,N_42341,N_40200);
xnor U44268 (N_44268,N_42027,N_42015);
or U44269 (N_44269,N_41969,N_40008);
nor U44270 (N_44270,N_42072,N_41281);
or U44271 (N_44271,N_40547,N_41931);
or U44272 (N_44272,N_40348,N_40426);
and U44273 (N_44273,N_40664,N_40697);
or U44274 (N_44274,N_42173,N_41544);
xnor U44275 (N_44275,N_41537,N_40537);
or U44276 (N_44276,N_40247,N_41767);
xnor U44277 (N_44277,N_42124,N_41398);
and U44278 (N_44278,N_42430,N_41814);
nor U44279 (N_44279,N_40913,N_41571);
nor U44280 (N_44280,N_42358,N_40086);
nand U44281 (N_44281,N_41496,N_40999);
or U44282 (N_44282,N_41742,N_40698);
nand U44283 (N_44283,N_42252,N_40780);
or U44284 (N_44284,N_42282,N_40287);
and U44285 (N_44285,N_41964,N_41469);
nor U44286 (N_44286,N_41123,N_40064);
and U44287 (N_44287,N_41752,N_42386);
or U44288 (N_44288,N_40353,N_41933);
or U44289 (N_44289,N_40940,N_41467);
nand U44290 (N_44290,N_40713,N_41606);
xnor U44291 (N_44291,N_41820,N_41904);
and U44292 (N_44292,N_41965,N_42074);
and U44293 (N_44293,N_41856,N_41877);
and U44294 (N_44294,N_40695,N_41884);
nand U44295 (N_44295,N_41136,N_41336);
xnor U44296 (N_44296,N_41038,N_41763);
xnor U44297 (N_44297,N_41668,N_42308);
xor U44298 (N_44298,N_41316,N_41235);
nor U44299 (N_44299,N_41444,N_41902);
nor U44300 (N_44300,N_41590,N_40716);
and U44301 (N_44301,N_41507,N_42141);
nor U44302 (N_44302,N_41818,N_40308);
nor U44303 (N_44303,N_41819,N_41235);
xor U44304 (N_44304,N_41113,N_42470);
and U44305 (N_44305,N_41683,N_41188);
xnor U44306 (N_44306,N_41858,N_41563);
xor U44307 (N_44307,N_41005,N_41217);
or U44308 (N_44308,N_41040,N_40193);
nand U44309 (N_44309,N_40201,N_40432);
nand U44310 (N_44310,N_41950,N_41569);
xnor U44311 (N_44311,N_40535,N_40730);
and U44312 (N_44312,N_42148,N_41720);
or U44313 (N_44313,N_40908,N_40012);
nor U44314 (N_44314,N_41168,N_40596);
nor U44315 (N_44315,N_42265,N_42235);
and U44316 (N_44316,N_41458,N_41880);
xnor U44317 (N_44317,N_40546,N_40788);
or U44318 (N_44318,N_40158,N_40167);
xnor U44319 (N_44319,N_40918,N_40721);
nand U44320 (N_44320,N_42208,N_41914);
nor U44321 (N_44321,N_40039,N_41208);
nand U44322 (N_44322,N_41634,N_40437);
xor U44323 (N_44323,N_40604,N_41112);
nand U44324 (N_44324,N_42423,N_41680);
nor U44325 (N_44325,N_40595,N_42213);
nor U44326 (N_44326,N_42182,N_41363);
xnor U44327 (N_44327,N_40706,N_40230);
or U44328 (N_44328,N_42011,N_40608);
xor U44329 (N_44329,N_40168,N_41744);
nand U44330 (N_44330,N_41503,N_41126);
or U44331 (N_44331,N_40281,N_42409);
xnor U44332 (N_44332,N_40684,N_40003);
nand U44333 (N_44333,N_40952,N_41520);
and U44334 (N_44334,N_40592,N_40997);
and U44335 (N_44335,N_42494,N_40820);
or U44336 (N_44336,N_41182,N_40187);
and U44337 (N_44337,N_40404,N_41368);
and U44338 (N_44338,N_41393,N_41706);
or U44339 (N_44339,N_41907,N_40830);
nor U44340 (N_44340,N_41176,N_41103);
or U44341 (N_44341,N_41202,N_42214);
nand U44342 (N_44342,N_42334,N_40007);
xnor U44343 (N_44343,N_41606,N_41597);
xor U44344 (N_44344,N_41014,N_42399);
and U44345 (N_44345,N_42269,N_40891);
xor U44346 (N_44346,N_40498,N_42143);
nor U44347 (N_44347,N_40582,N_41644);
or U44348 (N_44348,N_40427,N_40992);
nor U44349 (N_44349,N_42240,N_41788);
nand U44350 (N_44350,N_40931,N_40342);
and U44351 (N_44351,N_40869,N_42353);
and U44352 (N_44352,N_40606,N_41353);
or U44353 (N_44353,N_40780,N_40295);
or U44354 (N_44354,N_40655,N_42074);
nor U44355 (N_44355,N_40763,N_40608);
and U44356 (N_44356,N_41861,N_40574);
xnor U44357 (N_44357,N_41184,N_40399);
xor U44358 (N_44358,N_41496,N_41411);
and U44359 (N_44359,N_42446,N_41211);
or U44360 (N_44360,N_41265,N_41132);
xnor U44361 (N_44361,N_42222,N_41164);
nor U44362 (N_44362,N_41887,N_40490);
xor U44363 (N_44363,N_41789,N_40818);
nand U44364 (N_44364,N_40044,N_40728);
or U44365 (N_44365,N_41959,N_42283);
nor U44366 (N_44366,N_40688,N_40995);
nor U44367 (N_44367,N_42230,N_41281);
or U44368 (N_44368,N_41589,N_42298);
nor U44369 (N_44369,N_40358,N_42268);
xnor U44370 (N_44370,N_40559,N_41552);
and U44371 (N_44371,N_41700,N_41873);
nand U44372 (N_44372,N_42034,N_40107);
or U44373 (N_44373,N_42097,N_41431);
and U44374 (N_44374,N_40983,N_40368);
xnor U44375 (N_44375,N_41430,N_41101);
or U44376 (N_44376,N_40195,N_41836);
nor U44377 (N_44377,N_40948,N_40457);
nor U44378 (N_44378,N_40292,N_41695);
and U44379 (N_44379,N_41827,N_42199);
and U44380 (N_44380,N_42234,N_41529);
nor U44381 (N_44381,N_42456,N_41223);
nor U44382 (N_44382,N_40237,N_42311);
xnor U44383 (N_44383,N_42230,N_40984);
and U44384 (N_44384,N_42360,N_40396);
nor U44385 (N_44385,N_40347,N_40605);
and U44386 (N_44386,N_41920,N_40065);
or U44387 (N_44387,N_41003,N_40440);
nor U44388 (N_44388,N_42378,N_41578);
nor U44389 (N_44389,N_42209,N_42371);
xnor U44390 (N_44390,N_41983,N_40737);
nand U44391 (N_44391,N_40435,N_40792);
and U44392 (N_44392,N_41867,N_41345);
or U44393 (N_44393,N_40963,N_42389);
nand U44394 (N_44394,N_41924,N_42047);
nor U44395 (N_44395,N_41262,N_40486);
or U44396 (N_44396,N_41151,N_42447);
xnor U44397 (N_44397,N_41663,N_40803);
xnor U44398 (N_44398,N_41085,N_40368);
and U44399 (N_44399,N_40343,N_40984);
xor U44400 (N_44400,N_42108,N_40655);
nor U44401 (N_44401,N_41817,N_41609);
and U44402 (N_44402,N_42409,N_41816);
and U44403 (N_44403,N_40809,N_41192);
or U44404 (N_44404,N_41570,N_42348);
nor U44405 (N_44405,N_41916,N_40338);
nor U44406 (N_44406,N_41508,N_41890);
and U44407 (N_44407,N_40324,N_41954);
and U44408 (N_44408,N_41914,N_42202);
nor U44409 (N_44409,N_41097,N_41600);
nor U44410 (N_44410,N_41085,N_41464);
nand U44411 (N_44411,N_41107,N_41125);
or U44412 (N_44412,N_41179,N_40015);
or U44413 (N_44413,N_40491,N_41210);
xor U44414 (N_44414,N_42096,N_42206);
nand U44415 (N_44415,N_40129,N_40975);
nor U44416 (N_44416,N_41926,N_42130);
nor U44417 (N_44417,N_40024,N_41856);
nand U44418 (N_44418,N_40119,N_41943);
nor U44419 (N_44419,N_42149,N_42431);
or U44420 (N_44420,N_41679,N_42213);
and U44421 (N_44421,N_42084,N_42314);
or U44422 (N_44422,N_41140,N_41707);
xnor U44423 (N_44423,N_40946,N_42210);
or U44424 (N_44424,N_41333,N_42281);
or U44425 (N_44425,N_42314,N_41688);
nand U44426 (N_44426,N_41192,N_40495);
nor U44427 (N_44427,N_42072,N_42033);
or U44428 (N_44428,N_42228,N_42350);
nand U44429 (N_44429,N_41345,N_41792);
nand U44430 (N_44430,N_41956,N_40464);
nand U44431 (N_44431,N_42333,N_42468);
nor U44432 (N_44432,N_40416,N_40974);
xnor U44433 (N_44433,N_42393,N_42214);
nand U44434 (N_44434,N_40432,N_40648);
or U44435 (N_44435,N_42261,N_41036);
or U44436 (N_44436,N_40073,N_42451);
or U44437 (N_44437,N_41124,N_40555);
xnor U44438 (N_44438,N_41009,N_41676);
xnor U44439 (N_44439,N_40992,N_40542);
or U44440 (N_44440,N_41631,N_40474);
xnor U44441 (N_44441,N_40422,N_41375);
nand U44442 (N_44442,N_40461,N_41259);
and U44443 (N_44443,N_41154,N_41545);
xor U44444 (N_44444,N_41423,N_41832);
nor U44445 (N_44445,N_42428,N_41847);
nand U44446 (N_44446,N_40269,N_41469);
or U44447 (N_44447,N_41079,N_41795);
nand U44448 (N_44448,N_40866,N_40190);
nor U44449 (N_44449,N_41962,N_40516);
and U44450 (N_44450,N_41627,N_40919);
nor U44451 (N_44451,N_40015,N_40157);
nand U44452 (N_44452,N_42084,N_40793);
nand U44453 (N_44453,N_40943,N_40330);
nor U44454 (N_44454,N_40798,N_42358);
xnor U44455 (N_44455,N_40780,N_40044);
or U44456 (N_44456,N_40083,N_40646);
or U44457 (N_44457,N_42361,N_40944);
xor U44458 (N_44458,N_41164,N_40985);
or U44459 (N_44459,N_42089,N_41198);
or U44460 (N_44460,N_41253,N_42490);
and U44461 (N_44461,N_41489,N_41430);
nand U44462 (N_44462,N_42377,N_41065);
or U44463 (N_44463,N_42228,N_41668);
nor U44464 (N_44464,N_41321,N_40078);
nor U44465 (N_44465,N_41716,N_41145);
and U44466 (N_44466,N_40347,N_42119);
nand U44467 (N_44467,N_41252,N_41894);
nor U44468 (N_44468,N_40263,N_40144);
xnor U44469 (N_44469,N_41588,N_41025);
xor U44470 (N_44470,N_41329,N_42198);
or U44471 (N_44471,N_40444,N_40395);
nor U44472 (N_44472,N_40264,N_41889);
and U44473 (N_44473,N_40600,N_40300);
and U44474 (N_44474,N_41361,N_41038);
or U44475 (N_44475,N_40658,N_41139);
or U44476 (N_44476,N_41476,N_41734);
and U44477 (N_44477,N_40160,N_42287);
xnor U44478 (N_44478,N_40291,N_41544);
or U44479 (N_44479,N_40435,N_40987);
or U44480 (N_44480,N_40302,N_41891);
xnor U44481 (N_44481,N_42294,N_41420);
nor U44482 (N_44482,N_41967,N_41443);
nor U44483 (N_44483,N_41029,N_40509);
nand U44484 (N_44484,N_40076,N_40961);
and U44485 (N_44485,N_42403,N_40733);
nand U44486 (N_44486,N_41313,N_41091);
or U44487 (N_44487,N_41692,N_41799);
or U44488 (N_44488,N_41615,N_42491);
nand U44489 (N_44489,N_41325,N_40731);
nor U44490 (N_44490,N_40269,N_41430);
nor U44491 (N_44491,N_41245,N_40004);
nand U44492 (N_44492,N_40108,N_41593);
xnor U44493 (N_44493,N_41696,N_40742);
nor U44494 (N_44494,N_42296,N_41506);
xnor U44495 (N_44495,N_42170,N_40306);
nor U44496 (N_44496,N_40118,N_41214);
and U44497 (N_44497,N_40811,N_40869);
or U44498 (N_44498,N_41660,N_41446);
and U44499 (N_44499,N_40041,N_40089);
nand U44500 (N_44500,N_41661,N_40475);
xor U44501 (N_44501,N_40597,N_40769);
nor U44502 (N_44502,N_42346,N_40582);
xor U44503 (N_44503,N_41142,N_41387);
nor U44504 (N_44504,N_41175,N_40170);
or U44505 (N_44505,N_40451,N_40494);
and U44506 (N_44506,N_40035,N_42142);
and U44507 (N_44507,N_41659,N_42371);
nor U44508 (N_44508,N_40347,N_40532);
nor U44509 (N_44509,N_40012,N_42243);
nor U44510 (N_44510,N_40714,N_40161);
or U44511 (N_44511,N_40349,N_40907);
nand U44512 (N_44512,N_42021,N_40162);
or U44513 (N_44513,N_40540,N_41700);
or U44514 (N_44514,N_40174,N_40941);
or U44515 (N_44515,N_41646,N_42204);
and U44516 (N_44516,N_42052,N_41210);
nand U44517 (N_44517,N_40024,N_40745);
nor U44518 (N_44518,N_42396,N_41526);
nand U44519 (N_44519,N_40796,N_41911);
and U44520 (N_44520,N_40027,N_40081);
xnor U44521 (N_44521,N_41559,N_41710);
nor U44522 (N_44522,N_41095,N_40351);
nand U44523 (N_44523,N_41223,N_40353);
and U44524 (N_44524,N_40834,N_41084);
or U44525 (N_44525,N_41622,N_40021);
and U44526 (N_44526,N_40497,N_40208);
xnor U44527 (N_44527,N_40233,N_40634);
nand U44528 (N_44528,N_40362,N_41961);
nor U44529 (N_44529,N_41123,N_40767);
nand U44530 (N_44530,N_40299,N_40856);
and U44531 (N_44531,N_40963,N_41262);
and U44532 (N_44532,N_41516,N_40951);
nand U44533 (N_44533,N_41944,N_42124);
nor U44534 (N_44534,N_41028,N_40181);
nor U44535 (N_44535,N_41825,N_41343);
and U44536 (N_44536,N_42323,N_42410);
xnor U44537 (N_44537,N_40168,N_41501);
nor U44538 (N_44538,N_40819,N_40358);
and U44539 (N_44539,N_40674,N_41343);
nor U44540 (N_44540,N_41691,N_42102);
and U44541 (N_44541,N_40192,N_40117);
xor U44542 (N_44542,N_40053,N_40225);
xnor U44543 (N_44543,N_41929,N_41449);
nor U44544 (N_44544,N_40370,N_40373);
nor U44545 (N_44545,N_41196,N_40780);
nor U44546 (N_44546,N_40252,N_40292);
nor U44547 (N_44547,N_40688,N_42086);
xnor U44548 (N_44548,N_42068,N_40619);
or U44549 (N_44549,N_42017,N_40452);
xor U44550 (N_44550,N_41818,N_41572);
and U44551 (N_44551,N_40069,N_41184);
and U44552 (N_44552,N_40274,N_40949);
xor U44553 (N_44553,N_42268,N_41321);
and U44554 (N_44554,N_40361,N_41894);
nor U44555 (N_44555,N_41633,N_41870);
xnor U44556 (N_44556,N_41596,N_42355);
xor U44557 (N_44557,N_41415,N_40817);
and U44558 (N_44558,N_41152,N_40623);
nand U44559 (N_44559,N_41412,N_41734);
nand U44560 (N_44560,N_40876,N_40839);
xnor U44561 (N_44561,N_40114,N_40302);
xnor U44562 (N_44562,N_40296,N_41459);
and U44563 (N_44563,N_42199,N_41069);
nand U44564 (N_44564,N_41575,N_41633);
or U44565 (N_44565,N_41571,N_40942);
xnor U44566 (N_44566,N_40672,N_41802);
or U44567 (N_44567,N_41113,N_41475);
nand U44568 (N_44568,N_40969,N_41714);
nand U44569 (N_44569,N_40838,N_41806);
xor U44570 (N_44570,N_41764,N_41392);
nor U44571 (N_44571,N_40514,N_42031);
xor U44572 (N_44572,N_42468,N_41878);
nand U44573 (N_44573,N_40739,N_40620);
nand U44574 (N_44574,N_41683,N_40933);
nand U44575 (N_44575,N_41636,N_41210);
or U44576 (N_44576,N_42165,N_40754);
or U44577 (N_44577,N_42261,N_41982);
or U44578 (N_44578,N_41041,N_41823);
nor U44579 (N_44579,N_42408,N_41240);
and U44580 (N_44580,N_40977,N_41264);
or U44581 (N_44581,N_40930,N_42030);
and U44582 (N_44582,N_40646,N_41146);
xor U44583 (N_44583,N_40720,N_42199);
and U44584 (N_44584,N_41587,N_42197);
nor U44585 (N_44585,N_41023,N_40974);
or U44586 (N_44586,N_41675,N_41410);
and U44587 (N_44587,N_41017,N_40011);
or U44588 (N_44588,N_42370,N_41979);
and U44589 (N_44589,N_41277,N_42460);
and U44590 (N_44590,N_41916,N_40688);
or U44591 (N_44591,N_40363,N_42301);
and U44592 (N_44592,N_40475,N_40960);
nor U44593 (N_44593,N_42227,N_41283);
xnor U44594 (N_44594,N_41101,N_40719);
xor U44595 (N_44595,N_42391,N_41428);
nor U44596 (N_44596,N_41821,N_40821);
and U44597 (N_44597,N_40637,N_42182);
nor U44598 (N_44598,N_41830,N_41577);
nand U44599 (N_44599,N_40257,N_42123);
nor U44600 (N_44600,N_40310,N_42037);
nor U44601 (N_44601,N_40946,N_40645);
nand U44602 (N_44602,N_41950,N_40108);
xor U44603 (N_44603,N_40884,N_41062);
xnor U44604 (N_44604,N_41922,N_42178);
nand U44605 (N_44605,N_41217,N_40261);
or U44606 (N_44606,N_40434,N_41959);
nand U44607 (N_44607,N_42384,N_41035);
xor U44608 (N_44608,N_40123,N_40647);
and U44609 (N_44609,N_42370,N_41648);
nand U44610 (N_44610,N_42455,N_40728);
xor U44611 (N_44611,N_40281,N_41487);
and U44612 (N_44612,N_40938,N_40706);
and U44613 (N_44613,N_41207,N_41576);
nand U44614 (N_44614,N_40904,N_42242);
or U44615 (N_44615,N_40561,N_42154);
or U44616 (N_44616,N_41587,N_41509);
and U44617 (N_44617,N_42424,N_42335);
or U44618 (N_44618,N_41164,N_40043);
nor U44619 (N_44619,N_41057,N_41248);
and U44620 (N_44620,N_41107,N_40606);
or U44621 (N_44621,N_40515,N_42040);
nor U44622 (N_44622,N_41225,N_41522);
nor U44623 (N_44623,N_41778,N_40069);
xnor U44624 (N_44624,N_41627,N_41699);
nand U44625 (N_44625,N_40685,N_40063);
xnor U44626 (N_44626,N_41686,N_42371);
nor U44627 (N_44627,N_40682,N_40485);
or U44628 (N_44628,N_41083,N_42071);
xor U44629 (N_44629,N_41673,N_40764);
nand U44630 (N_44630,N_42306,N_42348);
xnor U44631 (N_44631,N_41300,N_40963);
nand U44632 (N_44632,N_40425,N_41453);
xnor U44633 (N_44633,N_40849,N_42131);
or U44634 (N_44634,N_40402,N_41324);
xnor U44635 (N_44635,N_41802,N_40757);
and U44636 (N_44636,N_41173,N_40594);
or U44637 (N_44637,N_40900,N_42350);
or U44638 (N_44638,N_40028,N_40025);
and U44639 (N_44639,N_40665,N_41222);
or U44640 (N_44640,N_41272,N_41506);
and U44641 (N_44641,N_40820,N_40084);
nand U44642 (N_44642,N_40244,N_40703);
or U44643 (N_44643,N_41778,N_41617);
xor U44644 (N_44644,N_41496,N_40275);
and U44645 (N_44645,N_42055,N_42210);
nor U44646 (N_44646,N_41799,N_41252);
or U44647 (N_44647,N_41887,N_40796);
nand U44648 (N_44648,N_40237,N_42262);
and U44649 (N_44649,N_42145,N_41919);
or U44650 (N_44650,N_41180,N_42017);
and U44651 (N_44651,N_40116,N_42165);
xor U44652 (N_44652,N_40177,N_42009);
nand U44653 (N_44653,N_41969,N_41938);
nand U44654 (N_44654,N_42127,N_42422);
or U44655 (N_44655,N_41666,N_40545);
nor U44656 (N_44656,N_41219,N_41035);
and U44657 (N_44657,N_41744,N_40939);
xnor U44658 (N_44658,N_40751,N_41959);
and U44659 (N_44659,N_41101,N_41160);
and U44660 (N_44660,N_41415,N_42164);
or U44661 (N_44661,N_41001,N_40725);
and U44662 (N_44662,N_40255,N_41029);
nand U44663 (N_44663,N_41739,N_41035);
nor U44664 (N_44664,N_40292,N_41743);
and U44665 (N_44665,N_42355,N_40913);
nor U44666 (N_44666,N_41679,N_41514);
nand U44667 (N_44667,N_40188,N_41120);
and U44668 (N_44668,N_40429,N_41774);
or U44669 (N_44669,N_42258,N_40409);
or U44670 (N_44670,N_40400,N_41570);
nand U44671 (N_44671,N_40071,N_40277);
nor U44672 (N_44672,N_40674,N_42399);
nand U44673 (N_44673,N_41233,N_40562);
nor U44674 (N_44674,N_42103,N_41330);
nor U44675 (N_44675,N_41897,N_42060);
xor U44676 (N_44676,N_40963,N_41467);
or U44677 (N_44677,N_40033,N_41814);
and U44678 (N_44678,N_41679,N_40939);
xnor U44679 (N_44679,N_41620,N_40761);
and U44680 (N_44680,N_40148,N_41789);
and U44681 (N_44681,N_42478,N_42397);
nand U44682 (N_44682,N_42391,N_41628);
or U44683 (N_44683,N_42325,N_41702);
nor U44684 (N_44684,N_40585,N_41030);
nor U44685 (N_44685,N_41485,N_42349);
xnor U44686 (N_44686,N_41485,N_42093);
or U44687 (N_44687,N_41881,N_41675);
or U44688 (N_44688,N_41510,N_40029);
or U44689 (N_44689,N_40195,N_40759);
xnor U44690 (N_44690,N_42431,N_40975);
nor U44691 (N_44691,N_42491,N_40421);
and U44692 (N_44692,N_40928,N_40870);
and U44693 (N_44693,N_41608,N_42317);
and U44694 (N_44694,N_41007,N_42072);
xnor U44695 (N_44695,N_40936,N_40012);
nor U44696 (N_44696,N_40981,N_42271);
and U44697 (N_44697,N_41250,N_41271);
nor U44698 (N_44698,N_41463,N_41270);
xor U44699 (N_44699,N_40462,N_40354);
xor U44700 (N_44700,N_42448,N_40588);
and U44701 (N_44701,N_41474,N_41023);
xnor U44702 (N_44702,N_40046,N_42406);
nor U44703 (N_44703,N_41076,N_42103);
nor U44704 (N_44704,N_40722,N_40860);
xnor U44705 (N_44705,N_42146,N_40392);
nand U44706 (N_44706,N_42259,N_42014);
xnor U44707 (N_44707,N_41921,N_40107);
nand U44708 (N_44708,N_42033,N_40318);
and U44709 (N_44709,N_40191,N_41039);
xor U44710 (N_44710,N_40613,N_42211);
and U44711 (N_44711,N_41818,N_41277);
and U44712 (N_44712,N_40094,N_41673);
nor U44713 (N_44713,N_42010,N_41868);
nand U44714 (N_44714,N_42390,N_40209);
nand U44715 (N_44715,N_41640,N_41693);
nand U44716 (N_44716,N_40174,N_41201);
nor U44717 (N_44717,N_41557,N_41042);
xnor U44718 (N_44718,N_40318,N_40144);
nor U44719 (N_44719,N_40467,N_42036);
nor U44720 (N_44720,N_41009,N_41951);
nor U44721 (N_44721,N_40284,N_40523);
and U44722 (N_44722,N_41786,N_41834);
or U44723 (N_44723,N_40964,N_41258);
nand U44724 (N_44724,N_40925,N_41246);
xor U44725 (N_44725,N_41940,N_42373);
or U44726 (N_44726,N_41707,N_40643);
or U44727 (N_44727,N_41159,N_41464);
nand U44728 (N_44728,N_41398,N_41705);
or U44729 (N_44729,N_40481,N_41051);
xnor U44730 (N_44730,N_41365,N_41406);
or U44731 (N_44731,N_41084,N_40717);
nand U44732 (N_44732,N_40037,N_41220);
xor U44733 (N_44733,N_41369,N_42431);
nor U44734 (N_44734,N_41195,N_42130);
or U44735 (N_44735,N_41835,N_40966);
nor U44736 (N_44736,N_42288,N_41301);
and U44737 (N_44737,N_41990,N_40453);
and U44738 (N_44738,N_40001,N_41549);
or U44739 (N_44739,N_40329,N_40101);
or U44740 (N_44740,N_41017,N_41020);
xnor U44741 (N_44741,N_42162,N_40890);
nor U44742 (N_44742,N_42288,N_42290);
nand U44743 (N_44743,N_41721,N_40733);
xor U44744 (N_44744,N_40037,N_40222);
xor U44745 (N_44745,N_41007,N_41876);
nand U44746 (N_44746,N_40325,N_41218);
nor U44747 (N_44747,N_42335,N_42134);
or U44748 (N_44748,N_41925,N_40812);
or U44749 (N_44749,N_42215,N_42318);
or U44750 (N_44750,N_41686,N_40069);
xor U44751 (N_44751,N_40011,N_40428);
nor U44752 (N_44752,N_40930,N_40453);
nor U44753 (N_44753,N_40537,N_42151);
nand U44754 (N_44754,N_41499,N_42493);
nor U44755 (N_44755,N_41891,N_41168);
xor U44756 (N_44756,N_42112,N_41290);
and U44757 (N_44757,N_40674,N_41353);
xor U44758 (N_44758,N_40581,N_40242);
and U44759 (N_44759,N_40851,N_41231);
nand U44760 (N_44760,N_41857,N_40309);
nor U44761 (N_44761,N_40252,N_40565);
nor U44762 (N_44762,N_40322,N_40114);
and U44763 (N_44763,N_41714,N_41647);
or U44764 (N_44764,N_42194,N_40915);
nor U44765 (N_44765,N_41743,N_42006);
xor U44766 (N_44766,N_42450,N_41881);
nor U44767 (N_44767,N_40992,N_42035);
and U44768 (N_44768,N_41517,N_41101);
xnor U44769 (N_44769,N_41241,N_41136);
nor U44770 (N_44770,N_41302,N_42218);
and U44771 (N_44771,N_40011,N_41703);
nor U44772 (N_44772,N_42118,N_41490);
and U44773 (N_44773,N_41756,N_40840);
nor U44774 (N_44774,N_42204,N_41030);
and U44775 (N_44775,N_42024,N_41266);
nand U44776 (N_44776,N_40514,N_41406);
or U44777 (N_44777,N_41468,N_40492);
xnor U44778 (N_44778,N_41071,N_41131);
or U44779 (N_44779,N_40910,N_40235);
and U44780 (N_44780,N_41237,N_41850);
nand U44781 (N_44781,N_41109,N_40287);
or U44782 (N_44782,N_40109,N_41051);
xor U44783 (N_44783,N_42214,N_40618);
and U44784 (N_44784,N_41925,N_40146);
and U44785 (N_44785,N_41262,N_40820);
nor U44786 (N_44786,N_41324,N_41126);
nor U44787 (N_44787,N_41236,N_42323);
nor U44788 (N_44788,N_40916,N_40362);
xnor U44789 (N_44789,N_40897,N_41425);
nor U44790 (N_44790,N_40242,N_40315);
nor U44791 (N_44791,N_40875,N_42059);
and U44792 (N_44792,N_41058,N_40916);
or U44793 (N_44793,N_40839,N_41170);
nor U44794 (N_44794,N_41769,N_40732);
nor U44795 (N_44795,N_42018,N_42028);
xor U44796 (N_44796,N_40235,N_41338);
nand U44797 (N_44797,N_41898,N_41456);
nor U44798 (N_44798,N_41533,N_41867);
or U44799 (N_44799,N_40366,N_41381);
nand U44800 (N_44800,N_40836,N_40117);
nand U44801 (N_44801,N_41446,N_42478);
xor U44802 (N_44802,N_40890,N_41491);
nand U44803 (N_44803,N_41764,N_40983);
nand U44804 (N_44804,N_41527,N_41097);
or U44805 (N_44805,N_41418,N_42241);
nor U44806 (N_44806,N_42177,N_40450);
and U44807 (N_44807,N_40544,N_42134);
or U44808 (N_44808,N_41355,N_40496);
xor U44809 (N_44809,N_40070,N_40789);
or U44810 (N_44810,N_41940,N_41299);
nor U44811 (N_44811,N_41288,N_41973);
xor U44812 (N_44812,N_42123,N_41776);
nor U44813 (N_44813,N_40854,N_41043);
or U44814 (N_44814,N_41995,N_41353);
xnor U44815 (N_44815,N_42351,N_40503);
and U44816 (N_44816,N_41958,N_40020);
nand U44817 (N_44817,N_42321,N_40167);
xor U44818 (N_44818,N_42150,N_41188);
and U44819 (N_44819,N_42252,N_40816);
nor U44820 (N_44820,N_40111,N_40401);
nor U44821 (N_44821,N_40519,N_41516);
nor U44822 (N_44822,N_42236,N_40609);
nand U44823 (N_44823,N_40705,N_41484);
and U44824 (N_44824,N_41440,N_41758);
xnor U44825 (N_44825,N_41615,N_41626);
nand U44826 (N_44826,N_40549,N_40037);
xor U44827 (N_44827,N_41135,N_40627);
nor U44828 (N_44828,N_42027,N_41598);
and U44829 (N_44829,N_41782,N_40505);
xor U44830 (N_44830,N_41040,N_41369);
or U44831 (N_44831,N_40877,N_41630);
xor U44832 (N_44832,N_41736,N_40106);
or U44833 (N_44833,N_41602,N_41928);
xor U44834 (N_44834,N_40591,N_40029);
or U44835 (N_44835,N_41291,N_41154);
xnor U44836 (N_44836,N_41932,N_40864);
and U44837 (N_44837,N_40372,N_41331);
nor U44838 (N_44838,N_40015,N_41425);
nor U44839 (N_44839,N_40861,N_41214);
xor U44840 (N_44840,N_42230,N_40703);
nor U44841 (N_44841,N_42163,N_40102);
xor U44842 (N_44842,N_40162,N_41227);
xor U44843 (N_44843,N_41457,N_42422);
nand U44844 (N_44844,N_40184,N_42373);
or U44845 (N_44845,N_40331,N_42460);
xor U44846 (N_44846,N_40934,N_42381);
xor U44847 (N_44847,N_40863,N_41444);
or U44848 (N_44848,N_40233,N_42306);
nand U44849 (N_44849,N_40758,N_42137);
xnor U44850 (N_44850,N_40120,N_42183);
nor U44851 (N_44851,N_41347,N_42300);
nand U44852 (N_44852,N_42224,N_41490);
nor U44853 (N_44853,N_40230,N_42404);
nor U44854 (N_44854,N_41645,N_41853);
nand U44855 (N_44855,N_41568,N_41715);
xor U44856 (N_44856,N_41490,N_40392);
nand U44857 (N_44857,N_41279,N_40457);
xor U44858 (N_44858,N_41244,N_40316);
or U44859 (N_44859,N_41125,N_41303);
nor U44860 (N_44860,N_42360,N_41810);
nand U44861 (N_44861,N_40657,N_41898);
or U44862 (N_44862,N_41984,N_42198);
or U44863 (N_44863,N_41096,N_41084);
or U44864 (N_44864,N_42493,N_42172);
and U44865 (N_44865,N_41129,N_41411);
nand U44866 (N_44866,N_41164,N_40833);
xnor U44867 (N_44867,N_41078,N_40882);
nand U44868 (N_44868,N_41603,N_41333);
nand U44869 (N_44869,N_40505,N_41480);
nor U44870 (N_44870,N_41055,N_42487);
or U44871 (N_44871,N_40305,N_42427);
or U44872 (N_44872,N_41498,N_40287);
or U44873 (N_44873,N_41197,N_40287);
nor U44874 (N_44874,N_42411,N_42162);
nand U44875 (N_44875,N_41705,N_41756);
nor U44876 (N_44876,N_41895,N_41601);
xnor U44877 (N_44877,N_41539,N_40345);
nor U44878 (N_44878,N_40884,N_40776);
or U44879 (N_44879,N_42020,N_40086);
or U44880 (N_44880,N_42482,N_41629);
nor U44881 (N_44881,N_42140,N_41839);
xor U44882 (N_44882,N_40126,N_41158);
nor U44883 (N_44883,N_40803,N_40238);
nand U44884 (N_44884,N_41481,N_41519);
nor U44885 (N_44885,N_42479,N_40458);
xor U44886 (N_44886,N_40644,N_40667);
xnor U44887 (N_44887,N_40553,N_41490);
nor U44888 (N_44888,N_42447,N_42373);
and U44889 (N_44889,N_41329,N_40887);
nand U44890 (N_44890,N_42039,N_41382);
or U44891 (N_44891,N_40603,N_41978);
or U44892 (N_44892,N_41806,N_42138);
nor U44893 (N_44893,N_42148,N_41231);
xnor U44894 (N_44894,N_41161,N_40924);
and U44895 (N_44895,N_41915,N_40664);
and U44896 (N_44896,N_40135,N_40932);
nor U44897 (N_44897,N_41015,N_40859);
and U44898 (N_44898,N_41768,N_41841);
and U44899 (N_44899,N_41203,N_40434);
nor U44900 (N_44900,N_40992,N_41472);
nor U44901 (N_44901,N_40940,N_41839);
or U44902 (N_44902,N_42180,N_41036);
xnor U44903 (N_44903,N_41763,N_40897);
nor U44904 (N_44904,N_40088,N_40495);
or U44905 (N_44905,N_42146,N_42302);
and U44906 (N_44906,N_40805,N_40082);
nand U44907 (N_44907,N_41789,N_42088);
nor U44908 (N_44908,N_42085,N_41136);
or U44909 (N_44909,N_40144,N_42229);
and U44910 (N_44910,N_40130,N_41297);
nand U44911 (N_44911,N_41355,N_41026);
xnor U44912 (N_44912,N_41661,N_42367);
and U44913 (N_44913,N_40216,N_40167);
xor U44914 (N_44914,N_42131,N_40031);
and U44915 (N_44915,N_41271,N_40484);
xnor U44916 (N_44916,N_40728,N_41671);
nand U44917 (N_44917,N_41311,N_41538);
xor U44918 (N_44918,N_40460,N_42241);
and U44919 (N_44919,N_42083,N_42369);
and U44920 (N_44920,N_41199,N_41987);
and U44921 (N_44921,N_41274,N_41334);
or U44922 (N_44922,N_40147,N_42344);
or U44923 (N_44923,N_41866,N_41470);
and U44924 (N_44924,N_41155,N_40350);
xor U44925 (N_44925,N_42308,N_41687);
nor U44926 (N_44926,N_40829,N_40706);
or U44927 (N_44927,N_40068,N_41059);
or U44928 (N_44928,N_41377,N_42485);
nor U44929 (N_44929,N_41590,N_40324);
nor U44930 (N_44930,N_41000,N_40370);
nand U44931 (N_44931,N_42446,N_41818);
xnor U44932 (N_44932,N_41798,N_40635);
and U44933 (N_44933,N_40199,N_41227);
and U44934 (N_44934,N_40422,N_40393);
nand U44935 (N_44935,N_41186,N_41489);
nor U44936 (N_44936,N_40183,N_40641);
xnor U44937 (N_44937,N_40522,N_42278);
xnor U44938 (N_44938,N_41713,N_41970);
xnor U44939 (N_44939,N_42452,N_40329);
or U44940 (N_44940,N_41967,N_41635);
xor U44941 (N_44941,N_42314,N_41526);
nand U44942 (N_44942,N_40987,N_42334);
nand U44943 (N_44943,N_42388,N_41952);
xnor U44944 (N_44944,N_41280,N_42224);
and U44945 (N_44945,N_41370,N_41242);
nor U44946 (N_44946,N_41252,N_42309);
or U44947 (N_44947,N_41686,N_40007);
and U44948 (N_44948,N_42234,N_40877);
and U44949 (N_44949,N_42243,N_40037);
xnor U44950 (N_44950,N_42139,N_41700);
nand U44951 (N_44951,N_42262,N_41538);
nor U44952 (N_44952,N_42212,N_42452);
and U44953 (N_44953,N_40340,N_42499);
and U44954 (N_44954,N_41981,N_42256);
or U44955 (N_44955,N_40204,N_41109);
nand U44956 (N_44956,N_40535,N_40935);
xor U44957 (N_44957,N_42068,N_41107);
and U44958 (N_44958,N_41826,N_40872);
xor U44959 (N_44959,N_40214,N_40917);
nand U44960 (N_44960,N_42290,N_41115);
and U44961 (N_44961,N_41379,N_40726);
nor U44962 (N_44962,N_42392,N_42292);
or U44963 (N_44963,N_41639,N_41615);
nor U44964 (N_44964,N_40260,N_41853);
xnor U44965 (N_44965,N_40045,N_41650);
xnor U44966 (N_44966,N_42015,N_40569);
nand U44967 (N_44967,N_41389,N_40248);
and U44968 (N_44968,N_40129,N_40797);
nor U44969 (N_44969,N_40212,N_42190);
nor U44970 (N_44970,N_42114,N_40911);
nor U44971 (N_44971,N_40981,N_40507);
and U44972 (N_44972,N_40570,N_41905);
nand U44973 (N_44973,N_40955,N_41347);
nand U44974 (N_44974,N_40436,N_41430);
and U44975 (N_44975,N_41182,N_42310);
nand U44976 (N_44976,N_41750,N_40114);
nor U44977 (N_44977,N_40360,N_40566);
nor U44978 (N_44978,N_40123,N_42400);
nand U44979 (N_44979,N_41102,N_41971);
and U44980 (N_44980,N_40677,N_40326);
nand U44981 (N_44981,N_42115,N_40171);
nor U44982 (N_44982,N_40192,N_40855);
and U44983 (N_44983,N_40031,N_41885);
and U44984 (N_44984,N_40858,N_41674);
and U44985 (N_44985,N_42316,N_40795);
nor U44986 (N_44986,N_40309,N_41182);
or U44987 (N_44987,N_40885,N_40936);
or U44988 (N_44988,N_40327,N_41623);
or U44989 (N_44989,N_41999,N_40403);
and U44990 (N_44990,N_40928,N_40526);
nand U44991 (N_44991,N_40436,N_41968);
nand U44992 (N_44992,N_41599,N_40107);
or U44993 (N_44993,N_42464,N_41290);
nand U44994 (N_44994,N_40549,N_41783);
or U44995 (N_44995,N_40030,N_40074);
nor U44996 (N_44996,N_40191,N_40047);
nand U44997 (N_44997,N_41455,N_42412);
or U44998 (N_44998,N_41056,N_41584);
and U44999 (N_44999,N_40199,N_40870);
and U45000 (N_45000,N_44274,N_42968);
and U45001 (N_45001,N_43395,N_44534);
or U45002 (N_45002,N_44853,N_43916);
xnor U45003 (N_45003,N_43702,N_44894);
nand U45004 (N_45004,N_43477,N_43364);
and U45005 (N_45005,N_42823,N_44405);
nor U45006 (N_45006,N_43978,N_43407);
or U45007 (N_45007,N_44200,N_44602);
nand U45008 (N_45008,N_43119,N_44331);
and U45009 (N_45009,N_44151,N_43253);
or U45010 (N_45010,N_44635,N_42527);
nand U45011 (N_45011,N_44092,N_43362);
and U45012 (N_45012,N_43758,N_43274);
nor U45013 (N_45013,N_43520,N_44778);
nor U45014 (N_45014,N_44655,N_43834);
nor U45015 (N_45015,N_43228,N_42937);
nand U45016 (N_45016,N_42695,N_42628);
or U45017 (N_45017,N_42649,N_42733);
or U45018 (N_45018,N_42729,N_43366);
nand U45019 (N_45019,N_43210,N_44085);
nor U45020 (N_45020,N_44217,N_43763);
or U45021 (N_45021,N_43236,N_43280);
and U45022 (N_45022,N_44024,N_43466);
or U45023 (N_45023,N_43318,N_43083);
nor U45024 (N_45024,N_44075,N_43807);
xor U45025 (N_45025,N_44834,N_44388);
xnor U45026 (N_45026,N_43955,N_42963);
nor U45027 (N_45027,N_43115,N_43729);
nand U45028 (N_45028,N_44225,N_44559);
nand U45029 (N_45029,N_42935,N_44163);
nand U45030 (N_45030,N_43966,N_44667);
and U45031 (N_45031,N_43932,N_42533);
nor U45032 (N_45032,N_44960,N_44153);
and U45033 (N_45033,N_42718,N_42832);
or U45034 (N_45034,N_43441,N_43679);
nor U45035 (N_45035,N_43433,N_44745);
nand U45036 (N_45036,N_44913,N_44098);
xnor U45037 (N_45037,N_44901,N_43211);
or U45038 (N_45038,N_42940,N_44156);
nand U45039 (N_45039,N_42517,N_44760);
xor U45040 (N_45040,N_42711,N_44513);
xnor U45041 (N_45041,N_43390,N_43394);
or U45042 (N_45042,N_44932,N_43411);
or U45043 (N_45043,N_43335,N_43252);
nor U45044 (N_45044,N_42550,N_43560);
or U45045 (N_45045,N_44194,N_42822);
and U45046 (N_45046,N_42707,N_44143);
or U45047 (N_45047,N_43435,N_44781);
and U45048 (N_45048,N_44027,N_44251);
nand U45049 (N_45049,N_42507,N_44307);
nor U45050 (N_45050,N_44701,N_44650);
and U45051 (N_45051,N_44657,N_43842);
nor U45052 (N_45052,N_43712,N_42787);
nand U45053 (N_45053,N_43111,N_43895);
nor U45054 (N_45054,N_43731,N_44668);
nand U45055 (N_45055,N_44228,N_43569);
or U45056 (N_45056,N_44483,N_43371);
xnor U45057 (N_45057,N_43962,N_44378);
or U45058 (N_45058,N_44939,N_42900);
or U45059 (N_45059,N_43685,N_43740);
or U45060 (N_45060,N_44533,N_43457);
xor U45061 (N_45061,N_42677,N_43845);
nand U45062 (N_45062,N_44010,N_44077);
xnor U45063 (N_45063,N_43913,N_44006);
nor U45064 (N_45064,N_42613,N_44576);
xor U45065 (N_45065,N_42849,N_43891);
and U45066 (N_45066,N_42957,N_43381);
or U45067 (N_45067,N_44353,N_44541);
nand U45068 (N_45068,N_44833,N_43308);
and U45069 (N_45069,N_43596,N_44662);
nand U45070 (N_45070,N_43440,N_43225);
and U45071 (N_45071,N_43697,N_44794);
nor U45072 (N_45072,N_43444,N_44830);
and U45073 (N_45073,N_42591,N_44545);
or U45074 (N_45074,N_44881,N_44676);
or U45075 (N_45075,N_42619,N_43808);
and U45076 (N_45076,N_42709,N_43059);
xor U45077 (N_45077,N_43271,N_43859);
or U45078 (N_45078,N_44306,N_44494);
or U45079 (N_45079,N_42809,N_44066);
and U45080 (N_45080,N_44443,N_42859);
nand U45081 (N_45081,N_43028,N_42518);
xor U45082 (N_45082,N_42881,N_43741);
xor U45083 (N_45083,N_42555,N_43613);
nor U45084 (N_45084,N_43460,N_44209);
nor U45085 (N_45085,N_44614,N_44294);
or U45086 (N_45086,N_43802,N_44957);
nand U45087 (N_45087,N_43629,N_44051);
nor U45088 (N_45088,N_44882,N_44696);
xor U45089 (N_45089,N_44162,N_43076);
and U45090 (N_45090,N_44688,N_42973);
nor U45091 (N_45091,N_43705,N_44698);
xnor U45092 (N_45092,N_42567,N_44221);
or U45093 (N_45093,N_44304,N_43298);
and U45094 (N_45094,N_44604,N_44038);
xnor U45095 (N_45095,N_43197,N_44368);
and U45096 (N_45096,N_44183,N_42767);
nand U45097 (N_45097,N_42853,N_42757);
nor U45098 (N_45098,N_44507,N_42576);
xor U45099 (N_45099,N_43899,N_44815);
or U45100 (N_45100,N_44465,N_43812);
and U45101 (N_45101,N_43577,N_42717);
or U45102 (N_45102,N_44551,N_43150);
or U45103 (N_45103,N_44325,N_42728);
xnor U45104 (N_45104,N_44334,N_44827);
or U45105 (N_45105,N_43355,N_43536);
xnor U45106 (N_45106,N_44210,N_44869);
or U45107 (N_45107,N_44977,N_44768);
or U45108 (N_45108,N_43941,N_43869);
nand U45109 (N_45109,N_43148,N_42835);
xor U45110 (N_45110,N_42573,N_43296);
nor U45111 (N_45111,N_44298,N_43305);
xor U45112 (N_45112,N_44617,N_43222);
xor U45113 (N_45113,N_43114,N_44850);
xor U45114 (N_45114,N_44326,N_44980);
nor U45115 (N_45115,N_42916,N_44241);
nor U45116 (N_45116,N_43368,N_43455);
and U45117 (N_45117,N_42858,N_44192);
nand U45118 (N_45118,N_44190,N_44346);
xor U45119 (N_45119,N_44372,N_44218);
or U45120 (N_45120,N_42735,N_44376);
nand U45121 (N_45121,N_42948,N_43626);
nand U45122 (N_45122,N_44630,N_44505);
and U45123 (N_45123,N_43208,N_42755);
xor U45124 (N_45124,N_44742,N_42909);
nand U45125 (N_45125,N_44680,N_43982);
or U45126 (N_45126,N_43202,N_43074);
nor U45127 (N_45127,N_44837,N_44240);
nor U45128 (N_45128,N_43868,N_43288);
and U45129 (N_45129,N_43224,N_42821);
or U45130 (N_45130,N_43397,N_44305);
and U45131 (N_45131,N_43841,N_44057);
nor U45132 (N_45132,N_42843,N_44223);
or U45133 (N_45133,N_44040,N_42949);
xnor U45134 (N_45134,N_42596,N_43461);
and U45135 (N_45135,N_44642,N_43609);
nand U45136 (N_45136,N_43980,N_43401);
nand U45137 (N_45137,N_44076,N_44741);
or U45138 (N_45138,N_43662,N_44452);
and U45139 (N_45139,N_43557,N_44422);
nor U45140 (N_45140,N_43742,N_43940);
nor U45141 (N_45141,N_44284,N_43116);
nor U45142 (N_45142,N_44165,N_43836);
or U45143 (N_45143,N_44234,N_43176);
nand U45144 (N_45144,N_44523,N_43944);
or U45145 (N_45145,N_44003,N_43535);
and U45146 (N_45146,N_44054,N_44252);
xnor U45147 (N_45147,N_44538,N_44934);
xor U45148 (N_45148,N_43534,N_42913);
or U45149 (N_45149,N_42698,N_43948);
and U45150 (N_45150,N_43649,N_43524);
nor U45151 (N_45151,N_44945,N_44863);
xor U45152 (N_45152,N_44019,N_44640);
nand U45153 (N_45153,N_43102,N_44062);
nand U45154 (N_45154,N_43694,N_43618);
and U45155 (N_45155,N_43840,N_44787);
or U45156 (N_45156,N_43526,N_43965);
nand U45157 (N_45157,N_43277,N_43391);
xor U45158 (N_45158,N_43322,N_44170);
nand U45159 (N_45159,N_42540,N_44986);
or U45160 (N_45160,N_42522,N_44904);
or U45161 (N_45161,N_44127,N_44258);
and U45162 (N_45162,N_43934,N_42924);
and U45163 (N_45163,N_42623,N_43814);
nor U45164 (N_45164,N_43797,N_43794);
nor U45165 (N_45165,N_44785,N_42675);
nand U45166 (N_45166,N_44289,N_42632);
or U45167 (N_45167,N_44421,N_44502);
nand U45168 (N_45168,N_44395,N_44966);
or U45169 (N_45169,N_44141,N_43585);
and U45170 (N_45170,N_43929,N_43959);
or U45171 (N_45171,N_44364,N_43147);
or U45172 (N_45172,N_43857,N_42626);
nand U45173 (N_45173,N_42988,N_43961);
and U45174 (N_45174,N_43768,N_43843);
nor U45175 (N_45175,N_44261,N_43799);
xnor U45176 (N_45176,N_44048,N_43786);
nor U45177 (N_45177,N_44566,N_44964);
or U45178 (N_45178,N_42923,N_42993);
xnor U45179 (N_45179,N_43789,N_43738);
nand U45180 (N_45180,N_44029,N_44328);
and U45181 (N_45181,N_42813,N_42865);
or U45182 (N_45182,N_42722,N_43620);
or U45183 (N_45183,N_42788,N_44387);
xnor U45184 (N_45184,N_43704,N_43553);
xor U45185 (N_45185,N_42910,N_44779);
nor U45186 (N_45186,N_42726,N_44799);
nor U45187 (N_45187,N_42559,N_44755);
nand U45188 (N_45188,N_44885,N_44080);
or U45189 (N_45189,N_44990,N_44503);
and U45190 (N_45190,N_43587,N_43552);
and U45191 (N_45191,N_43903,N_43290);
and U45192 (N_45192,N_44584,N_43319);
or U45193 (N_45193,N_43402,N_44301);
nand U45194 (N_45194,N_42793,N_44256);
and U45195 (N_45195,N_42580,N_44236);
xnor U45196 (N_45196,N_44591,N_44970);
nand U45197 (N_45197,N_42724,N_43549);
nor U45198 (N_45198,N_43610,N_44825);
xor U45199 (N_45199,N_43492,N_44101);
and U45200 (N_45200,N_42955,N_43668);
or U45201 (N_45201,N_42647,N_43042);
nor U45202 (N_45202,N_43581,N_42713);
nand U45203 (N_45203,N_43498,N_42500);
and U45204 (N_45204,N_42561,N_44925);
or U45205 (N_45205,N_44540,N_42621);
xor U45206 (N_45206,N_43241,N_42674);
nor U45207 (N_45207,N_44568,N_44644);
or U45208 (N_45208,N_44453,N_44175);
xor U45209 (N_45209,N_43954,N_44809);
nor U45210 (N_45210,N_43356,N_42781);
nand U45211 (N_45211,N_43576,N_42952);
nor U45212 (N_45212,N_42702,N_43725);
nand U45213 (N_45213,N_43917,N_42504);
nand U45214 (N_45214,N_44474,N_44664);
and U45215 (N_45215,N_44302,N_44413);
or U45216 (N_45216,N_43947,N_44823);
xnor U45217 (N_45217,N_43328,N_44117);
xnor U45218 (N_45218,N_43136,N_44148);
xor U45219 (N_45219,N_42575,N_44951);
and U45220 (N_45220,N_42592,N_43212);
and U45221 (N_45221,N_43453,N_42556);
nor U45222 (N_45222,N_44435,N_43227);
and U45223 (N_45223,N_42691,N_43058);
and U45224 (N_45224,N_44738,N_44020);
or U45225 (N_45225,N_44748,N_43201);
nor U45226 (N_45226,N_44345,N_44426);
nor U45227 (N_45227,N_44341,N_44877);
nand U45228 (N_45228,N_44014,N_42523);
and U45229 (N_45229,N_44268,N_43465);
nor U45230 (N_45230,N_43816,N_42611);
nand U45231 (N_45231,N_44731,N_42503);
nor U45232 (N_45232,N_44616,N_42971);
and U45233 (N_45233,N_44628,N_44246);
nor U45234 (N_45234,N_44081,N_44828);
nand U45235 (N_45235,N_43990,N_44373);
or U45236 (N_45236,N_42866,N_44173);
or U45237 (N_45237,N_44404,N_44619);
nor U45238 (N_45238,N_44102,N_44247);
nor U45239 (N_45239,N_43527,N_42985);
nor U45240 (N_45240,N_43299,N_44466);
nand U45241 (N_45241,N_44311,N_42921);
or U45242 (N_45242,N_42954,N_44976);
nor U45243 (N_45243,N_42699,N_42583);
xor U45244 (N_45244,N_44047,N_44016);
and U45245 (N_45245,N_44734,N_42829);
nand U45246 (N_45246,N_44999,N_43693);
nand U45247 (N_45247,N_42799,N_43728);
and U45248 (N_45248,N_42740,N_43973);
xnor U45249 (N_45249,N_43025,N_44931);
and U45250 (N_45250,N_44436,N_42933);
xor U45251 (N_45251,N_42815,N_43006);
nand U45252 (N_45252,N_42844,N_44312);
nor U45253 (N_45253,N_43467,N_43017);
xor U45254 (N_45254,N_44295,N_44119);
xnor U45255 (N_45255,N_42884,N_44407);
and U45256 (N_45256,N_44536,N_43765);
nand U45257 (N_45257,N_44681,N_44758);
nor U45258 (N_45258,N_42607,N_44764);
or U45259 (N_45259,N_43777,N_42666);
nor U45260 (N_45260,N_43508,N_43332);
and U45261 (N_45261,N_44031,N_42908);
xor U45262 (N_45262,N_43021,N_43723);
or U45263 (N_45263,N_44214,N_42936);
and U45264 (N_45264,N_42593,N_44557);
xor U45265 (N_45265,N_43753,N_42743);
and U45266 (N_45266,N_43811,N_43504);
nand U45267 (N_45267,N_44692,N_44993);
or U45268 (N_45268,N_43471,N_43080);
nand U45269 (N_45269,N_43478,N_44458);
nor U45270 (N_45270,N_44535,N_43923);
nand U45271 (N_45271,N_43098,N_42552);
or U45272 (N_45272,N_44313,N_42679);
xor U45273 (N_45273,N_43281,N_44586);
nand U45274 (N_45274,N_44780,N_44233);
or U45275 (N_45275,N_43924,N_42554);
xor U45276 (N_45276,N_42801,N_42557);
or U45277 (N_45277,N_43522,N_43282);
xor U45278 (N_45278,N_42651,N_43986);
xnor U45279 (N_45279,N_44385,N_43935);
and U45280 (N_45280,N_42771,N_43583);
or U45281 (N_45281,N_42609,N_43635);
or U45282 (N_45282,N_43078,N_44457);
nand U45283 (N_45283,N_42814,N_44686);
or U45284 (N_45284,N_43315,N_42978);
xnor U45285 (N_45285,N_44903,N_44125);
nor U45286 (N_45286,N_43051,N_44866);
nand U45287 (N_45287,N_44208,N_42762);
or U45288 (N_45288,N_44929,N_44475);
nor U45289 (N_45289,N_43594,N_42779);
or U45290 (N_45290,N_43882,N_43068);
nand U45291 (N_45291,N_42848,N_44814);
and U45292 (N_45292,N_44093,N_43169);
or U45293 (N_45293,N_44273,N_44271);
nor U45294 (N_45294,N_44752,N_44079);
nor U45295 (N_45295,N_43369,N_42586);
xnor U45296 (N_45296,N_42511,N_43950);
or U45297 (N_45297,N_44154,N_43748);
xnor U45298 (N_45298,N_43687,N_42692);
nor U45299 (N_45299,N_43582,N_42579);
nor U45300 (N_45300,N_44499,N_43547);
nand U45301 (N_45301,N_43656,N_43447);
xnor U45302 (N_45302,N_43245,N_44041);
nand U45303 (N_45303,N_43974,N_42629);
or U45304 (N_45304,N_44260,N_44023);
and U45305 (N_45305,N_44266,N_43121);
and U45306 (N_45306,N_43064,N_42680);
nor U45307 (N_45307,N_44136,N_42716);
or U45308 (N_45308,N_44276,N_43854);
xnor U45309 (N_45309,N_43486,N_44878);
xor U45310 (N_45310,N_44623,N_44615);
or U45311 (N_45311,N_44107,N_43928);
nor U45312 (N_45312,N_42714,N_44918);
nor U45313 (N_45313,N_42806,N_44643);
nand U45314 (N_45314,N_43309,N_44028);
and U45315 (N_45315,N_42995,N_44105);
nand U45316 (N_45316,N_42548,N_44197);
xor U45317 (N_45317,N_42512,N_44508);
xor U45318 (N_45318,N_44442,N_43107);
nand U45319 (N_45319,N_44339,N_42927);
nand U45320 (N_45320,N_42947,N_43000);
and U45321 (N_45321,N_44609,N_44711);
or U45322 (N_45322,N_42636,N_43420);
nor U45323 (N_45323,N_43573,N_43472);
nand U45324 (N_45324,N_44606,N_42802);
xor U45325 (N_45325,N_42764,N_44033);
or U45326 (N_45326,N_43128,N_43695);
and U45327 (N_45327,N_43172,N_43353);
nor U45328 (N_45328,N_42683,N_43165);
and U45329 (N_45329,N_43427,N_43347);
xor U45330 (N_45330,N_43927,N_44174);
or U45331 (N_45331,N_44524,N_43782);
nor U45332 (N_45332,N_42574,N_43184);
and U45333 (N_45333,N_44481,N_44359);
nor U45334 (N_45334,N_44100,N_42687);
and U45335 (N_45335,N_42676,N_42950);
or U45336 (N_45336,N_43663,N_43297);
xor U45337 (N_45337,N_43769,N_43365);
xor U45338 (N_45338,N_44397,N_43654);
and U45339 (N_45339,N_43131,N_43852);
or U45340 (N_45340,N_42569,N_44791);
or U45341 (N_45341,N_43096,N_43911);
and U45342 (N_45342,N_44131,N_44230);
and U45343 (N_45343,N_43367,N_42820);
and U45344 (N_45344,N_43902,N_42519);
or U45345 (N_45345,N_44480,N_42774);
and U45346 (N_45346,N_44771,N_43181);
and U45347 (N_45347,N_44917,N_43358);
or U45348 (N_45348,N_44841,N_42706);
xnor U45349 (N_45349,N_43140,N_43396);
xor U45350 (N_45350,N_43469,N_44179);
xor U45351 (N_45351,N_42600,N_44546);
or U45352 (N_45352,N_44817,N_43788);
xnor U45353 (N_45353,N_42752,N_42833);
xor U45354 (N_45354,N_43135,N_43981);
xor U45355 (N_45355,N_43238,N_44928);
or U45356 (N_45356,N_43333,N_44467);
or U45357 (N_45357,N_43091,N_43943);
or U45358 (N_45358,N_43795,N_44050);
nor U45359 (N_45359,N_43791,N_43640);
or U45360 (N_45360,N_44892,N_42770);
xnor U45361 (N_45361,N_43832,N_43590);
and U45362 (N_45362,N_42520,N_42905);
nand U45363 (N_45363,N_42605,N_44981);
and U45364 (N_45364,N_43783,N_43592);
nand U45365 (N_45365,N_43041,N_44927);
nand U45366 (N_45366,N_44399,N_43343);
or U45367 (N_45367,N_43513,N_44042);
nand U45368 (N_45368,N_43045,N_44672);
xnor U45369 (N_45369,N_42989,N_43097);
and U45370 (N_45370,N_44155,N_44106);
nand U45371 (N_45371,N_44806,N_44821);
and U45372 (N_45372,N_43637,N_43246);
nand U45373 (N_45373,N_43256,N_44441);
and U45374 (N_45374,N_44521,N_43167);
and U45375 (N_45375,N_42610,N_43888);
xor U45376 (N_45376,N_44666,N_43776);
and U45377 (N_45377,N_43871,N_43864);
nand U45378 (N_45378,N_42922,N_44788);
or U45379 (N_45379,N_42502,N_43320);
xor U45380 (N_45380,N_43304,N_43700);
nor U45381 (N_45381,N_43523,N_44652);
nand U45382 (N_45382,N_43250,N_43105);
nor U45383 (N_45383,N_44908,N_42614);
and U45384 (N_45384,N_42654,N_44767);
nand U45385 (N_45385,N_42529,N_43951);
or U45386 (N_45386,N_43189,N_44888);
xnor U45387 (N_45387,N_44569,N_44431);
nand U45388 (N_45388,N_44001,N_44445);
nand U45389 (N_45389,N_44514,N_43410);
and U45390 (N_45390,N_43431,N_43608);
nand U45391 (N_45391,N_44451,N_43953);
or U45392 (N_45392,N_43785,N_44856);
and U45393 (N_45393,N_44425,N_42751);
nor U45394 (N_45394,N_42633,N_44510);
nand U45395 (N_45395,N_43010,N_44747);
nor U45396 (N_45396,N_44724,N_44820);
or U45397 (N_45397,N_42715,N_44542);
nand U45398 (N_45398,N_42560,N_44816);
xor U45399 (N_45399,N_43773,N_44037);
and U45400 (N_45400,N_44677,N_43039);
or U45401 (N_45401,N_42578,N_44839);
nand U45402 (N_45402,N_44718,N_42903);
nor U45403 (N_45403,N_44058,N_44570);
or U45404 (N_45404,N_43205,N_43260);
or U45405 (N_45405,N_44947,N_42773);
and U45406 (N_45406,N_43846,N_44227);
nor U45407 (N_45407,N_44789,N_43316);
xnor U45408 (N_45408,N_43813,N_42965);
nand U45409 (N_45409,N_44974,N_43050);
xnor U45410 (N_45410,N_44370,N_44801);
or U45411 (N_45411,N_44254,N_44340);
nor U45412 (N_45412,N_42791,N_44381);
xnor U45413 (N_45413,N_44206,N_44518);
or U45414 (N_45414,N_42531,N_42856);
nand U45415 (N_45415,N_42868,N_43752);
nor U45416 (N_45416,N_43511,N_44357);
or U45417 (N_45417,N_44746,N_44914);
or U45418 (N_45418,N_42759,N_44067);
nand U45419 (N_45419,N_44963,N_43889);
xnor U45420 (N_45420,N_43686,N_44418);
or U45421 (N_45421,N_43141,N_43220);
or U45422 (N_45422,N_44291,N_42765);
nor U45423 (N_45423,N_42758,N_42547);
and U45424 (N_45424,N_44184,N_42530);
xnor U45425 (N_45425,N_43601,N_43166);
and U45426 (N_45426,N_44958,N_44890);
and U45427 (N_45427,N_43484,N_44712);
or U45428 (N_45428,N_43699,N_42904);
nand U45429 (N_45429,N_43692,N_43030);
and U45430 (N_45430,N_42895,N_44257);
and U45431 (N_45431,N_43156,N_44461);
or U45432 (N_45432,N_43493,N_43805);
xor U45433 (N_45433,N_43239,N_44912);
and U45434 (N_45434,N_43920,N_43445);
or U45435 (N_45435,N_44496,N_44237);
and U45436 (N_45436,N_43602,N_44410);
xor U45437 (N_45437,N_42627,N_42543);
or U45438 (N_45438,N_42784,N_43195);
and U45439 (N_45439,N_44911,N_42741);
xnor U45440 (N_45440,N_43506,N_42671);
and U45441 (N_45441,N_43188,N_44950);
nor U45442 (N_45442,N_42710,N_43630);
or U45443 (N_45443,N_44553,N_43387);
and U45444 (N_45444,N_43247,N_44800);
nor U45445 (N_45445,N_44161,N_44953);
xor U45446 (N_45446,N_43317,N_42899);
or U45447 (N_45447,N_44498,N_44482);
nand U45448 (N_45448,N_43937,N_43866);
nand U45449 (N_45449,N_43993,N_44473);
or U45450 (N_45450,N_43338,N_44926);
nor U45451 (N_45451,N_42939,N_43894);
and U45452 (N_45452,N_43671,N_44180);
or U45453 (N_45453,N_44072,N_42945);
xor U45454 (N_45454,N_42887,N_43711);
or U45455 (N_45455,N_44025,N_44032);
xor U45456 (N_45456,N_43544,N_43625);
or U45457 (N_45457,N_44919,N_44375);
and U45458 (N_45458,N_43872,N_44978);
nor U45459 (N_45459,N_43715,N_42869);
nand U45460 (N_45460,N_43892,N_44133);
nand U45461 (N_45461,N_44279,N_43054);
and U45462 (N_45462,N_44969,N_42997);
and U45463 (N_45463,N_44068,N_44250);
or U45464 (N_45464,N_42852,N_43735);
nand U45465 (N_45465,N_43995,N_43746);
or U45466 (N_45466,N_42750,N_42977);
and U45467 (N_45467,N_42742,N_44786);
or U45468 (N_45468,N_44600,N_43830);
xor U45469 (N_45469,N_44808,N_44849);
and U45470 (N_45470,N_43254,N_42615);
and U45471 (N_45471,N_44782,N_44269);
xnor U45472 (N_45472,N_44300,N_44870);
or U45473 (N_45473,N_42516,N_43089);
or U45474 (N_45474,N_43018,N_43803);
xor U45475 (N_45475,N_43670,N_43910);
and U45476 (N_45476,N_43931,N_44398);
xnor U45477 (N_45477,N_43313,N_42652);
and U45478 (N_45478,N_44618,N_44103);
or U45479 (N_45479,N_43591,N_43144);
or U45480 (N_45480,N_43428,N_43790);
nor U45481 (N_45481,N_43767,N_44367);
or U45482 (N_45482,N_44716,N_43652);
nand U45483 (N_45483,N_42769,N_43530);
and U45484 (N_45484,N_42943,N_44198);
xor U45485 (N_45485,N_44139,N_42542);
nand U45486 (N_45486,N_44363,N_44776);
nor U45487 (N_45487,N_43209,N_44807);
or U45488 (N_45488,N_43709,N_44199);
or U45489 (N_45489,N_44959,N_43826);
nor U45490 (N_45490,N_43985,N_42775);
nor U45491 (N_45491,N_42785,N_42644);
nand U45492 (N_45492,N_44070,N_43230);
and U45493 (N_45493,N_42847,N_44308);
nand U45494 (N_45494,N_42842,N_43827);
xor U45495 (N_45495,N_44167,N_43015);
nor U45496 (N_45496,N_44558,N_42819);
or U45497 (N_45497,N_44922,N_44449);
nand U45498 (N_45498,N_43908,N_44594);
nor U45499 (N_45499,N_44211,N_44946);
or U45500 (N_45500,N_43120,N_44506);
nor U45501 (N_45501,N_44893,N_44543);
or U45502 (N_45502,N_43157,N_44641);
or U45503 (N_45503,N_42810,N_44347);
and U45504 (N_45504,N_44071,N_44561);
nor U45505 (N_45505,N_44181,N_44900);
or U45506 (N_45506,N_42812,N_44695);
and U45507 (N_45507,N_43837,N_43132);
nand U45508 (N_45508,N_44575,N_42723);
nor U45509 (N_45509,N_43645,N_42570);
or U45510 (N_45510,N_43754,N_44819);
xnor U45511 (N_45511,N_43370,N_42871);
or U45512 (N_45512,N_44396,N_44722);
xor U45513 (N_45513,N_44632,N_44725);
and U45514 (N_45514,N_42589,N_44318);
nand U45515 (N_45515,N_43339,N_44110);
nor U45516 (N_45516,N_44327,N_43858);
or U45517 (N_45517,N_44868,N_43994);
nand U45518 (N_45518,N_44477,N_43881);
xnor U45519 (N_45519,N_42883,N_43037);
nor U45520 (N_45520,N_44344,N_44203);
nand U45521 (N_45521,N_44299,N_43684);
or U45522 (N_45522,N_43405,N_44055);
nand U45523 (N_45523,N_43046,N_43286);
nor U45524 (N_45524,N_44262,N_44554);
nand U45525 (N_45525,N_43487,N_44484);
nor U45526 (N_45526,N_44061,N_43501);
nand U45527 (N_45527,N_44571,N_44560);
or U45528 (N_45528,N_44843,N_43603);
and U45529 (N_45529,N_42635,N_42890);
nand U45530 (N_45530,N_44515,N_44715);
or U45531 (N_45531,N_44259,N_42826);
nand U45532 (N_45532,N_42637,N_43792);
nand U45533 (N_45533,N_44146,N_43434);
xnor U45534 (N_45534,N_44333,N_43312);
xnor U45535 (N_45535,N_42951,N_44522);
and U45536 (N_45536,N_43716,N_44813);
nor U45537 (N_45537,N_44249,N_42896);
nor U45538 (N_45538,N_44109,N_43496);
nor U45539 (N_45539,N_44567,N_44171);
nand U45540 (N_45540,N_43106,N_43933);
nor U45541 (N_45541,N_44895,N_44035);
and U45542 (N_45542,N_44468,N_44137);
or U45543 (N_45543,N_44714,N_44287);
nor U45544 (N_45544,N_44416,N_43548);
nand U45545 (N_45545,N_43599,N_43022);
nor U45546 (N_45546,N_43632,N_43151);
nor U45547 (N_45547,N_43416,N_44842);
nand U45548 (N_45548,N_43240,N_44084);
or U45549 (N_45549,N_44777,N_44239);
and U45550 (N_45550,N_43232,N_43914);
nand U45551 (N_45551,N_44512,N_42508);
and U45552 (N_45552,N_43352,N_43867);
nand U45553 (N_45553,N_42514,N_44438);
nand U45554 (N_45554,N_44595,N_42992);
or U45555 (N_45555,N_44995,N_44090);
or U45556 (N_45556,N_43861,N_44428);
nor U45557 (N_45557,N_43023,N_43005);
and U45558 (N_45558,N_43681,N_42601);
nand U45559 (N_45559,N_44060,N_43450);
nor U45560 (N_45560,N_43052,N_44818);
nor U45561 (N_45561,N_44736,N_44665);
nor U45562 (N_45562,N_42824,N_43438);
and U45563 (N_45563,N_43988,N_43726);
xnor U45564 (N_45564,N_44226,N_43243);
nor U45565 (N_45565,N_43126,N_43464);
or U45566 (N_45566,N_43722,N_44631);
nor U45567 (N_45567,N_44574,N_43823);
and U45568 (N_45568,N_43856,N_43060);
and U45569 (N_45569,N_44380,N_44549);
xnor U45570 (N_45570,N_44625,N_44948);
nor U45571 (N_45571,N_44601,N_44988);
xnor U45572 (N_45572,N_42783,N_43113);
xor U45573 (N_45573,N_44906,N_42990);
or U45574 (N_45574,N_43302,N_44737);
and U45575 (N_45575,N_44487,N_43379);
nand U45576 (N_45576,N_43307,N_42725);
nand U45577 (N_45577,N_43701,N_43541);
nand U45578 (N_45578,N_43747,N_43730);
xor U45579 (N_45579,N_43027,N_43007);
and U45580 (N_45580,N_43512,N_42528);
or U45581 (N_45581,N_42686,N_42892);
nand U45582 (N_45582,N_43251,N_44094);
nand U45583 (N_45583,N_44573,N_44176);
and U45584 (N_45584,N_42587,N_42828);
nor U45585 (N_45585,N_43930,N_43915);
or U45586 (N_45586,N_43423,N_43456);
xnor U45587 (N_45587,N_42878,N_43031);
nor U45588 (N_45588,N_43013,N_44355);
nand U45589 (N_45589,N_44007,N_42689);
and U45590 (N_45590,N_43906,N_43714);
or U45591 (N_45591,N_42749,N_43925);
xor U45592 (N_45592,N_43226,N_43103);
nor U45593 (N_45593,N_43909,N_43997);
xnor U45594 (N_45594,N_44682,N_43154);
or U45595 (N_45595,N_43291,N_42545);
or U45596 (N_45596,N_44486,N_44952);
and U45597 (N_45597,N_44320,N_44717);
nor U45598 (N_45598,N_43070,N_42827);
nand U45599 (N_45599,N_44193,N_43886);
nand U45600 (N_45600,N_42705,N_44943);
nor U45601 (N_45601,N_43011,N_43542);
nand U45602 (N_45602,N_44243,N_43964);
and U45603 (N_45603,N_43839,N_43182);
or U45604 (N_45604,N_44915,N_44297);
nand U45605 (N_45605,N_44231,N_44743);
and U45606 (N_45606,N_44219,N_43200);
nand U45607 (N_45607,N_44649,N_43883);
nand U45608 (N_45608,N_43214,N_42792);
and U45609 (N_45609,N_44099,N_43771);
or U45610 (N_45610,N_43710,N_42846);
nand U45611 (N_45611,N_43393,N_44497);
or U45612 (N_45612,N_44059,N_44874);
xor U45613 (N_45613,N_42864,N_42982);
or U45614 (N_45614,N_43890,N_42501);
nand U45615 (N_45615,N_43720,N_44352);
and U45616 (N_45616,N_44790,N_44095);
nand U45617 (N_45617,N_43979,N_43904);
or U45618 (N_45618,N_42841,N_43960);
nand U45619 (N_45619,N_44824,N_43957);
nand U45620 (N_45620,N_43215,N_43255);
or U45621 (N_45621,N_44462,N_44675);
nand U45622 (N_45622,N_44578,N_44862);
and U45623 (N_45623,N_44708,N_44727);
or U45624 (N_45624,N_44865,N_44860);
nand U45625 (N_45625,N_43507,N_44867);
or U45626 (N_45626,N_43983,N_44845);
nor U45627 (N_45627,N_44844,N_44967);
nor U45628 (N_45628,N_44713,N_44158);
or U45629 (N_45629,N_44848,N_44610);
and U45630 (N_45630,N_44459,N_44750);
nor U45631 (N_45631,N_43556,N_44178);
nor U45632 (N_45632,N_43149,N_44884);
xor U45633 (N_45633,N_43644,N_42656);
nand U45634 (N_45634,N_42987,N_43999);
xor U45635 (N_45635,N_43533,N_44598);
or U45636 (N_45636,N_43636,N_43491);
or U45637 (N_45637,N_44621,N_43550);
or U45638 (N_45638,N_43117,N_42999);
nand U45639 (N_45639,N_44009,N_42658);
nand U45640 (N_45640,N_43554,N_44423);
nor U45641 (N_45641,N_43348,N_42776);
nand U45642 (N_45642,N_43284,N_43425);
nor U45643 (N_45643,N_44235,N_44394);
nor U45644 (N_45644,N_43651,N_44021);
xor U45645 (N_45645,N_44984,N_44377);
xor U45646 (N_45646,N_44292,N_44907);
nor U45647 (N_45647,N_43483,N_43183);
and U45648 (N_45648,N_44083,N_43806);
nand U45649 (N_45649,N_44005,N_43273);
and U45650 (N_45650,N_42855,N_44052);
nand U45651 (N_45651,N_43418,N_44773);
or U45652 (N_45652,N_44281,N_44444);
and U45653 (N_45653,N_44583,N_44648);
or U45654 (N_45654,N_43600,N_44485);
nand U45655 (N_45655,N_43584,N_44539);
nand U45656 (N_45656,N_43490,N_44086);
nand U45657 (N_45657,N_44253,N_44706);
or U45658 (N_45658,N_44429,N_42891);
nand U45659 (N_45659,N_42657,N_44303);
or U45660 (N_45660,N_43653,N_42625);
nand U45661 (N_45661,N_43760,N_43757);
nand U45662 (N_45662,N_43055,N_42551);
nand U45663 (N_45663,N_44147,N_42622);
nand U45664 (N_45664,N_43884,N_42811);
nor U45665 (N_45665,N_43939,N_44115);
nor U45666 (N_45666,N_44949,N_43546);
nand U45667 (N_45667,N_43593,N_42991);
nand U45668 (N_45668,N_43942,N_43809);
xor U45669 (N_45669,N_44729,N_44039);
xor U45670 (N_45670,N_44937,N_44403);
or U45671 (N_45671,N_42961,N_44417);
xor U45672 (N_45672,N_44470,N_43659);
or U45673 (N_45673,N_43489,N_43987);
or U45674 (N_45674,N_44599,N_43079);
nand U45675 (N_45675,N_43207,N_42660);
nor U45676 (N_45676,N_42539,N_43482);
or U45677 (N_45677,N_43623,N_44406);
and U45678 (N_45678,N_42642,N_44202);
nor U45679 (N_45679,N_43400,N_43996);
and U45680 (N_45680,N_44335,N_43505);
or U45681 (N_45681,N_42734,N_44012);
or U45682 (N_45682,N_44157,N_44871);
xnor U45683 (N_45683,N_43703,N_43706);
or U45684 (N_45684,N_44942,N_44605);
xnor U45685 (N_45685,N_43066,N_42582);
xor U45686 (N_45686,N_43887,N_44872);
nor U45687 (N_45687,N_42588,N_44548);
or U45688 (N_45688,N_44763,N_44544);
and U45689 (N_45689,N_43004,N_44899);
xnor U45690 (N_45690,N_43690,N_42796);
and U45691 (N_45691,N_43463,N_44622);
and U45692 (N_45692,N_43218,N_44620);
xor U45693 (N_45693,N_44792,N_43408);
or U45694 (N_45694,N_44354,N_44699);
nor U45695 (N_45695,N_42929,N_43870);
or U45696 (N_45696,N_43494,N_42838);
nor U45697 (N_45697,N_44011,N_42877);
and U45698 (N_45698,N_43860,N_43206);
nor U45699 (N_45699,N_44267,N_43152);
and U45700 (N_45700,N_43160,N_44213);
nor U45701 (N_45701,N_42938,N_43815);
or U45702 (N_45702,N_43991,N_43061);
and U45703 (N_45703,N_44660,N_44645);
xnor U45704 (N_45704,N_43907,N_42894);
nand U45705 (N_45705,N_44286,N_44002);
nor U45706 (N_45706,N_43604,N_44135);
nand U45707 (N_45707,N_43069,N_42672);
nand U45708 (N_45708,N_43249,N_44756);
xnor U45709 (N_45709,N_43158,N_44852);
nor U45710 (N_45710,N_44478,N_44495);
and U45711 (N_45711,N_43417,N_42874);
or U45712 (N_45712,N_43346,N_43342);
nor U45713 (N_45713,N_44069,N_44264);
nor U45714 (N_45714,N_43772,N_42782);
nand U45715 (N_45715,N_43634,N_43503);
and U45716 (N_45716,N_43952,N_43269);
or U45717 (N_45717,N_42777,N_44427);
or U45718 (N_45718,N_44189,N_44588);
nand U45719 (N_45719,N_44382,N_43674);
or U45720 (N_45720,N_43607,N_44030);
xnor U45721 (N_45721,N_44275,N_43597);
xor U45722 (N_45722,N_43231,N_43032);
nand U45723 (N_45723,N_43833,N_43191);
and U45724 (N_45724,N_42688,N_43056);
or U45725 (N_45725,N_42694,N_42685);
xnor U45726 (N_45726,N_43109,N_42831);
and U45727 (N_45727,N_44898,N_43235);
nand U45728 (N_45728,N_44700,N_44537);
nand U45729 (N_45729,N_43919,N_43545);
nand U45730 (N_45730,N_44739,N_43185);
and U45731 (N_45731,N_43561,N_43084);
or U45732 (N_45732,N_44826,N_43278);
and U45733 (N_45733,N_44805,N_43564);
nand U45734 (N_45734,N_43717,N_44684);
or U45735 (N_45735,N_44556,N_42928);
xor U45736 (N_45736,N_43646,N_44185);
xor U45737 (N_45737,N_42979,N_42648);
xnor U45738 (N_45738,N_43389,N_43421);
nor U45739 (N_45739,N_43631,N_44004);
or U45740 (N_45740,N_43458,N_43168);
xnor U45741 (N_45741,N_43330,N_44971);
or U45742 (N_45742,N_42918,N_44310);
and U45743 (N_45743,N_44940,N_44392);
or U45744 (N_45744,N_44693,N_43825);
nor U45745 (N_45745,N_44053,N_44469);
nor U45746 (N_45746,N_43268,N_42915);
nand U45747 (N_45747,N_43036,N_44348);
nand U45748 (N_45748,N_43223,N_42643);
xor U45749 (N_45749,N_43192,N_43244);
nor U45750 (N_45750,N_43012,N_42953);
nand U45751 (N_45751,N_44757,N_44994);
xor U45752 (N_45752,N_43562,N_44337);
xnor U45753 (N_45753,N_43666,N_44129);
nand U45754 (N_45754,N_43682,N_44420);
nand U45755 (N_45755,N_43436,N_42732);
or U45756 (N_45756,N_44204,N_43575);
xnor U45757 (N_45757,N_42532,N_43676);
nor U45758 (N_45758,N_43094,N_42753);
or U45759 (N_45759,N_44754,N_42960);
xor U45760 (N_45760,N_43664,N_44315);
nor U45761 (N_45761,N_42760,N_43551);
nor U45762 (N_45762,N_44683,N_43327);
and U45763 (N_45763,N_44968,N_42854);
or U45764 (N_45764,N_43350,N_42914);
xnor U45765 (N_45765,N_43331,N_42839);
nor U45766 (N_45766,N_43439,N_44338);
xor U45767 (N_45767,N_43388,N_44411);
xor U45768 (N_45768,N_44270,N_43043);
nor U45769 (N_45769,N_42983,N_42818);
nor U45770 (N_45770,N_44140,N_43779);
or U45771 (N_45771,N_44118,N_43563);
xor U45772 (N_45772,N_44530,N_43565);
nand U45773 (N_45773,N_44905,N_42684);
xnor U45774 (N_45774,N_43936,N_43009);
and U45775 (N_45775,N_44488,N_44391);
or U45776 (N_45776,N_42746,N_43409);
or U45777 (N_45777,N_43514,N_44280);
nor U45778 (N_45778,N_44879,N_43851);
or U45779 (N_45779,N_44587,N_43968);
or U45780 (N_45780,N_42521,N_43969);
xnor U45781 (N_45781,N_42739,N_44690);
nor U45782 (N_45782,N_42830,N_44552);
nand U45783 (N_45783,N_44531,N_42594);
nand U45784 (N_45784,N_43067,N_43992);
and U45785 (N_45785,N_44091,N_44638);
nor U45786 (N_45786,N_43164,N_43749);
nor U45787 (N_45787,N_44414,N_44191);
and U45788 (N_45788,N_42873,N_43171);
xor U45789 (N_45789,N_43821,N_44579);
xnor U45790 (N_45790,N_44245,N_42731);
or U45791 (N_45791,N_44244,N_44797);
or U45792 (N_45792,N_42737,N_42546);
xor U45793 (N_45793,N_44126,N_43516);
nand U45794 (N_45794,N_43901,N_43459);
nand U45795 (N_45795,N_44369,N_43784);
and U45796 (N_45796,N_44366,N_43124);
and U45797 (N_45797,N_44924,N_44324);
or U45798 (N_45798,N_43829,N_44384);
or U45799 (N_45799,N_42712,N_42704);
or U45800 (N_45800,N_42515,N_43614);
nand U45801 (N_45801,N_44329,N_43781);
xnor U45802 (N_45802,N_44113,N_44265);
nor U45803 (N_45803,N_44386,N_44705);
xnor U45804 (N_45804,N_43611,N_44150);
xor U45805 (N_45805,N_44653,N_42980);
xnor U45806 (N_45806,N_44766,N_43301);
nor U45807 (N_45807,N_42870,N_44242);
xor U45808 (N_45808,N_42640,N_43090);
and U45809 (N_45809,N_43627,N_43621);
and U45810 (N_45810,N_44350,N_43095);
or U45811 (N_45811,N_42558,N_44116);
or U45812 (N_45812,N_44547,N_42768);
xnor U45813 (N_45813,N_43326,N_44277);
or U45814 (N_45814,N_44840,N_43566);
or U45815 (N_45815,N_44972,N_42942);
xnor U45816 (N_45816,N_44679,N_44611);
nand U45817 (N_45817,N_42693,N_44238);
nand U45818 (N_45818,N_43403,N_42863);
xor U45819 (N_45819,N_44471,N_43673);
xor U45820 (N_45820,N_43835,N_44285);
nand U45821 (N_45821,N_44064,N_43270);
xnor U45822 (N_45822,N_42653,N_44400);
or U45823 (N_45823,N_42975,N_42981);
nor U45824 (N_45824,N_42837,N_44938);
nor U45825 (N_45825,N_43756,N_43828);
nand U45826 (N_45826,N_43775,N_42524);
or U45827 (N_45827,N_44582,N_43020);
xnor U45828 (N_45828,N_44634,N_43019);
xnor U45829 (N_45829,N_43125,N_43267);
nand U45830 (N_45830,N_43750,N_44463);
and U45831 (N_45831,N_42612,N_43258);
and U45832 (N_45832,N_44493,N_43572);
xor U45833 (N_45833,N_44804,N_44476);
nand U45834 (N_45834,N_44288,N_42670);
nor U45835 (N_45835,N_42825,N_44402);
and U45836 (N_45836,N_43034,N_42851);
and U45837 (N_45837,N_42595,N_43399);
or U45838 (N_45838,N_44159,N_43334);
nand U45839 (N_45839,N_42678,N_43329);
nand U45840 (N_45840,N_44319,N_43351);
xnor U45841 (N_45841,N_43497,N_43178);
and U45842 (N_45842,N_42646,N_43257);
xor U45843 (N_45843,N_43359,N_42624);
and U45844 (N_45844,N_42860,N_44026);
nand U45845 (N_45845,N_44795,N_44343);
nor U45846 (N_45846,N_44770,N_44454);
and U45847 (N_45847,N_43878,N_44783);
nor U45848 (N_45848,N_42564,N_43519);
xor U45849 (N_45849,N_43398,N_44489);
or U45850 (N_45850,N_44691,N_44751);
and U45851 (N_45851,N_43745,N_43110);
or U45852 (N_45852,N_44669,N_43574);
nand U45853 (N_45853,N_44580,N_43014);
nand U45854 (N_45854,N_42590,N_43127);
xor U45855 (N_45855,N_42850,N_44501);
nor U45856 (N_45856,N_44704,N_44603);
nand U45857 (N_45857,N_44596,N_42932);
xor U45858 (N_45858,N_42875,N_43404);
nand U45859 (N_45859,N_43377,N_42967);
nor U45860 (N_45860,N_42681,N_44448);
or U45861 (N_45861,N_44130,N_43718);
nor U45862 (N_45862,N_43129,N_42800);
xnor U45863 (N_45863,N_43155,N_43108);
and U45864 (N_45864,N_42616,N_43295);
nor U45865 (N_45865,N_42880,N_43448);
nor U45866 (N_45866,N_44613,N_44674);
and U45867 (N_45867,N_44593,N_44793);
nand U45868 (N_45868,N_44049,N_42754);
nand U45869 (N_45869,N_44362,N_43521);
or U45870 (N_45870,N_44627,N_43293);
xor U45871 (N_45871,N_44504,N_44263);
nor U45872 (N_45872,N_42766,N_43606);
nand U45873 (N_45873,N_43844,N_43972);
or U45874 (N_45874,N_43323,N_43633);
nand U45875 (N_45875,N_43605,N_43647);
nand U45876 (N_45876,N_44336,N_42525);
nor U45877 (N_45877,N_44608,N_43819);
or U45878 (N_45878,N_42650,N_43446);
nand U45879 (N_45879,N_44205,N_44719);
and U45880 (N_45880,N_43372,N_43531);
nor U45881 (N_45881,N_44342,N_44166);
or U45882 (N_45882,N_43146,N_44991);
or U45883 (N_45883,N_44108,N_44018);
or U45884 (N_45884,N_42565,N_44916);
and U45885 (N_45885,N_43719,N_44056);
nand U45886 (N_45886,N_43696,N_44654);
xnor U45887 (N_45887,N_42748,N_43893);
nor U45888 (N_45888,N_44744,N_42544);
nor U45889 (N_45889,N_43528,N_42703);
and U45890 (N_45890,N_44186,N_42912);
nor U45891 (N_45891,N_42667,N_43831);
nor U45892 (N_45892,N_43229,N_42700);
nand U45893 (N_45893,N_43595,N_43650);
nand U45894 (N_45894,N_43850,N_43029);
or U45895 (N_45895,N_43122,N_43073);
nor U45896 (N_45896,N_44753,N_43638);
and U45897 (N_45897,N_42571,N_44663);
and U45898 (N_45898,N_44015,N_44169);
nor U45899 (N_45899,N_43648,N_42645);
nand U45900 (N_45900,N_43798,N_43378);
or U45901 (N_45901,N_44733,N_42804);
or U45902 (N_45902,N_42931,N_42962);
and U45903 (N_45903,N_43509,N_43848);
and U45904 (N_45904,N_44321,N_44360);
nor U45905 (N_45905,N_43468,N_42563);
xor U45906 (N_45906,N_42719,N_44973);
and U45907 (N_45907,N_44529,N_43303);
xor U45908 (N_45908,N_44723,N_43219);
xor U45909 (N_45909,N_43495,N_42807);
nand U45910 (N_45910,N_43198,N_44216);
nand U45911 (N_45911,N_42599,N_43873);
or U45912 (N_45912,N_44356,N_44735);
or U45913 (N_45913,N_42944,N_43876);
nor U45914 (N_45914,N_44365,N_42996);
xnor U45915 (N_45915,N_42730,N_44624);
and U45916 (N_45916,N_43862,N_44168);
nor U45917 (N_45917,N_43265,N_43736);
or U45918 (N_45918,N_44525,N_42970);
or U45919 (N_45919,N_43849,N_43737);
xnor U45920 (N_45920,N_43261,N_44419);
or U45921 (N_45921,N_44432,N_43615);
and U45922 (N_45922,N_43667,N_43698);
and U45923 (N_45923,N_44811,N_42756);
or U45924 (N_45924,N_43196,N_43289);
xnor U45925 (N_45925,N_44550,N_44941);
and U45926 (N_45926,N_42876,N_42585);
nor U45927 (N_45927,N_44732,N_42534);
nand U45928 (N_45928,N_43118,N_44670);
and U45929 (N_45929,N_42797,N_43800);
or U45930 (N_45930,N_43093,N_43517);
and U45931 (N_45931,N_43003,N_44987);
nand U45932 (N_45932,N_43454,N_42617);
xor U45933 (N_45933,N_44073,N_44415);
or U45934 (N_45934,N_43071,N_44889);
or U45935 (N_45935,N_43989,N_44272);
xor U45936 (N_45936,N_43764,N_43744);
and U45937 (N_45937,N_44434,N_43689);
nand U45938 (N_45938,N_44961,N_43970);
nand U45939 (N_45939,N_42959,N_43529);
and U45940 (N_45940,N_44215,N_43161);
nand U45941 (N_45941,N_44212,N_44694);
and U45942 (N_45942,N_42745,N_43485);
nor U45943 (N_45943,N_42803,N_43442);
nor U45944 (N_45944,N_44207,N_43570);
nand U45945 (N_45945,N_43479,N_42631);
xor U45946 (N_45946,N_42697,N_44097);
nand U45947 (N_45947,N_44440,N_44673);
and U45948 (N_45948,N_44880,N_43213);
or U45949 (N_45949,N_43324,N_44702);
and U45950 (N_45950,N_43739,N_43008);
nand U45951 (N_45951,N_44316,N_44656);
nor U45952 (N_45952,N_44864,N_42630);
or U45953 (N_45953,N_43612,N_44332);
nor U45954 (N_45954,N_42690,N_43415);
nor U45955 (N_45955,N_44296,N_44659);
and U45956 (N_45956,N_42618,N_43360);
and U45957 (N_45957,N_42845,N_44720);
nand U45958 (N_45958,N_43437,N_42886);
xor U45959 (N_45959,N_43057,N_44784);
or U45960 (N_45960,N_43568,N_44962);
nor U45961 (N_45961,N_43233,N_43642);
and U45962 (N_45962,N_43540,N_42721);
xor U45963 (N_45963,N_44371,N_44887);
and U45964 (N_45964,N_43473,N_44726);
and U45965 (N_45965,N_43392,N_43145);
or U45966 (N_45966,N_44351,N_43755);
xnor U45967 (N_45967,N_44636,N_44728);
xnor U45968 (N_45968,N_43276,N_44074);
or U45969 (N_45969,N_43905,N_43162);
and U45970 (N_45970,N_43016,N_42778);
or U45971 (N_45971,N_44456,N_44172);
nor U45972 (N_45972,N_44492,N_42708);
and U45973 (N_45973,N_44152,N_43865);
xor U45974 (N_45974,N_42761,N_44846);
nand U45975 (N_45975,N_44944,N_44822);
xor U45976 (N_45976,N_44160,N_42639);
or U45977 (N_45977,N_43480,N_44661);
and U45978 (N_45978,N_43707,N_43430);
and U45979 (N_45979,N_44896,N_43921);
xor U45980 (N_45980,N_42893,N_43082);
or U45981 (N_45981,N_43657,N_44589);
xor U45982 (N_45982,N_42701,N_44857);
nand U45983 (N_45983,N_43967,N_43774);
or U45984 (N_45984,N_42946,N_44565);
xor U45985 (N_45985,N_43743,N_43159);
nand U45986 (N_45986,N_44122,N_43817);
nand U45987 (N_45987,N_43048,N_44430);
xnor U45988 (N_45988,N_44651,N_42727);
xor U45989 (N_45989,N_44248,N_44909);
xor U45990 (N_45990,N_44446,N_42572);
nand U45991 (N_45991,N_44532,N_43838);
and U45992 (N_45992,N_44920,N_44500);
nor U45993 (N_45993,N_44412,N_43539);
nand U45994 (N_45994,N_44390,N_43275);
nor U45995 (N_45995,N_44989,N_43759);
or U45996 (N_45996,N_43085,N_43658);
nor U45997 (N_45997,N_43672,N_43123);
nor U45998 (N_45998,N_44607,N_43262);
nand U45999 (N_45999,N_44526,N_43885);
nor U46000 (N_46000,N_42568,N_44293);
nand U46001 (N_46001,N_43818,N_44897);
xor U46002 (N_46002,N_43975,N_43810);
nor U46003 (N_46003,N_43855,N_43879);
nor U46004 (N_46004,N_43263,N_44282);
nand U46005 (N_46005,N_44802,N_42984);
nand U46006 (N_46006,N_44812,N_44861);
or U46007 (N_46007,N_44044,N_44612);
and U46008 (N_46008,N_42972,N_43088);
xnor U46009 (N_46009,N_44232,N_43306);
nand U46010 (N_46010,N_42620,N_44637);
and U46011 (N_46011,N_43248,N_44983);
nand U46012 (N_46012,N_43589,N_44022);
xnor U46013 (N_46013,N_43266,N_42872);
or U46014 (N_46014,N_43432,N_42505);
or U46015 (N_46015,N_43660,N_44930);
and U46016 (N_46016,N_42789,N_42906);
and U46017 (N_46017,N_43139,N_44687);
xnor U46018 (N_46018,N_43363,N_44374);
xor U46019 (N_46019,N_42911,N_44450);
or U46020 (N_46020,N_44979,N_43180);
xor U46021 (N_46021,N_43287,N_43001);
and U46022 (N_46022,N_42879,N_44401);
and U46023 (N_46023,N_43035,N_42661);
or U46024 (N_46024,N_44511,N_43385);
and U46025 (N_46025,N_42526,N_44224);
or U46026 (N_46026,N_44982,N_44838);
xnor U46027 (N_46027,N_44043,N_43525);
nor U46028 (N_46028,N_42986,N_44013);
xnor U46029 (N_46029,N_44201,N_44519);
nor U46030 (N_46030,N_43655,N_44424);
xor U46031 (N_46031,N_43532,N_43143);
nand U46032 (N_46032,N_42669,N_43543);
and U46033 (N_46033,N_44222,N_44323);
nor U46034 (N_46034,N_43134,N_42696);
nor U46035 (N_46035,N_44132,N_42744);
nand U46036 (N_46036,N_44509,N_43875);
or U46037 (N_46037,N_43279,N_42816);
or U46038 (N_46038,N_42663,N_43874);
and U46039 (N_46039,N_42974,N_43762);
xor U46040 (N_46040,N_44000,N_44383);
or U46041 (N_46041,N_44437,N_43778);
or U46042 (N_46042,N_42901,N_43414);
or U46043 (N_46043,N_43956,N_44798);
or U46044 (N_46044,N_42925,N_44078);
or U46045 (N_46045,N_43976,N_42926);
and U46046 (N_46046,N_44145,N_44516);
nor U46047 (N_46047,N_43361,N_44955);
nand U46048 (N_46048,N_42956,N_42897);
nor U46049 (N_46049,N_43880,N_43462);
nand U46050 (N_46050,N_42917,N_43053);
or U46051 (N_46051,N_44585,N_43203);
nor U46052 (N_46052,N_43337,N_44124);
xnor U46053 (N_46053,N_42958,N_42941);
or U46054 (N_46054,N_43216,N_43761);
and U46055 (N_46055,N_44309,N_44855);
nand U46056 (N_46056,N_44089,N_43040);
nand U46057 (N_46057,N_43661,N_42994);
nor U46058 (N_46058,N_44555,N_44710);
nand U46059 (N_46059,N_43515,N_44142);
nand U46060 (N_46060,N_43449,N_44965);
and U46061 (N_46061,N_43130,N_44290);
and U46062 (N_46062,N_43177,N_44647);
or U46063 (N_46063,N_43340,N_43376);
or U46064 (N_46064,N_42641,N_44490);
and U46065 (N_46065,N_43787,N_43724);
nand U46066 (N_46066,N_43087,N_43624);
nor U46067 (N_46067,N_44876,N_43510);
nor U46068 (N_46068,N_44997,N_44065);
nand U46069 (N_46069,N_43422,N_44935);
or U46070 (N_46070,N_43639,N_43187);
and U46071 (N_46071,N_44749,N_44439);
xnor U46072 (N_46072,N_43112,N_43499);
xnor U46073 (N_46073,N_44577,N_43669);
or U46074 (N_46074,N_43793,N_42606);
or U46075 (N_46075,N_42510,N_44096);
and U46076 (N_46076,N_42930,N_42763);
or U46077 (N_46077,N_42882,N_43822);
or U46078 (N_46078,N_44114,N_43946);
and U46079 (N_46079,N_43918,N_44088);
nand U46080 (N_46080,N_43217,N_43072);
or U46081 (N_46081,N_43081,N_43938);
or U46082 (N_46082,N_44597,N_44447);
xor U46083 (N_46083,N_44910,N_44590);
nor U46084 (N_46084,N_42541,N_44671);
and U46085 (N_46085,N_44358,N_44697);
and U46086 (N_46086,N_43443,N_42638);
xnor U46087 (N_46087,N_43796,N_43877);
xor U46088 (N_46088,N_43502,N_42862);
xnor U46089 (N_46089,N_43971,N_43419);
or U46090 (N_46090,N_43221,N_43863);
nor U46091 (N_46091,N_42720,N_43099);
xnor U46092 (N_46092,N_44581,N_43727);
or U46093 (N_46093,N_43044,N_44322);
xor U46094 (N_46094,N_43900,N_43683);
nor U46095 (N_46095,N_43194,N_42659);
nand U46096 (N_46096,N_44678,N_43958);
or U46097 (N_46097,N_44187,N_44633);
nand U46098 (N_46098,N_44772,N_43344);
nand U46099 (N_46099,N_43384,N_44149);
or U46100 (N_46100,N_44164,N_44873);
and U46101 (N_46101,N_42976,N_42857);
xor U46102 (N_46102,N_43678,N_42738);
xnor U46103 (N_46103,N_44528,N_44278);
nand U46104 (N_46104,N_44851,N_43922);
nand U46105 (N_46105,N_43853,N_43926);
nand U46106 (N_46106,N_44564,N_42634);
nor U46107 (N_46107,N_43579,N_43675);
xnor U46108 (N_46108,N_43896,N_42566);
or U46109 (N_46109,N_43451,N_43193);
xor U46110 (N_46110,N_44087,N_43984);
xor U46111 (N_46111,N_44527,N_43092);
nor U46112 (N_46112,N_42889,N_44803);
or U46113 (N_46113,N_43518,N_43429);
nor U46114 (N_46114,N_44036,N_43264);
nand U46115 (N_46115,N_43770,N_43578);
xor U46116 (N_46116,N_43588,N_44472);
or U46117 (N_46117,N_44646,N_43049);
nand U46118 (N_46118,N_42964,N_42902);
nand U46119 (N_46119,N_42736,N_44847);
or U46120 (N_46120,N_43500,N_43179);
nor U46121 (N_46121,N_43488,N_43153);
or U46122 (N_46122,N_44740,N_43104);
and U46123 (N_46123,N_44854,N_44709);
nand U46124 (N_46124,N_44936,N_43977);
or U46125 (N_46125,N_42898,N_42969);
nor U46126 (N_46126,N_43586,N_43382);
nor U46127 (N_46127,N_44996,N_44314);
xor U46128 (N_46128,N_42817,N_43033);
and U46129 (N_46129,N_43424,N_44658);
xor U46130 (N_46130,N_42581,N_43413);
or U46131 (N_46131,N_42786,N_44229);
nor U46132 (N_46132,N_43138,N_42867);
and U46133 (N_46133,N_42598,N_43801);
nand U46134 (N_46134,N_44762,N_43538);
xnor U46135 (N_46135,N_43945,N_43406);
and U46136 (N_46136,N_43426,N_42602);
or U46137 (N_46137,N_44975,N_44433);
and U46138 (N_46138,N_43175,N_44703);
nor U46139 (N_46139,N_43751,N_43101);
and U46140 (N_46140,N_43616,N_43002);
or U46141 (N_46141,N_44563,N_43294);
and U46142 (N_46142,N_42553,N_44188);
or U46143 (N_46143,N_43383,N_44562);
nand U46144 (N_46144,N_43475,N_42885);
nor U46145 (N_46145,N_44379,N_43847);
nor U46146 (N_46146,N_44769,N_43677);
or U46147 (N_46147,N_42861,N_44120);
nand U46148 (N_46148,N_44796,N_44045);
nor U46149 (N_46149,N_43024,N_42840);
xnor U46150 (N_46150,N_44517,N_44685);
and U46151 (N_46151,N_42888,N_42790);
xnor U46152 (N_46152,N_43998,N_42919);
nor U46153 (N_46153,N_43680,N_44765);
nand U46154 (N_46154,N_44491,N_44349);
or U46155 (N_46155,N_44832,N_43345);
or U46156 (N_46156,N_44121,N_43311);
or U46157 (N_46157,N_43285,N_44134);
or U46158 (N_46158,N_43537,N_44902);
xnor U46159 (N_46159,N_44759,N_44123);
nand U46160 (N_46160,N_42836,N_43732);
nor U46161 (N_46161,N_43373,N_43766);
and U46162 (N_46162,N_43321,N_43567);
xnor U46163 (N_46163,N_43357,N_43234);
xor U46164 (N_46164,N_43190,N_43580);
and U46165 (N_46165,N_43375,N_44361);
and U46166 (N_46166,N_43452,N_44985);
or U46167 (N_46167,N_44891,N_44034);
and U46168 (N_46168,N_43617,N_44730);
xor U46169 (N_46169,N_42780,N_43380);
and U46170 (N_46170,N_43100,N_43665);
and U46171 (N_46171,N_43733,N_42584);
and U46172 (N_46172,N_44283,N_44859);
xnor U46173 (N_46173,N_43622,N_44138);
or U46174 (N_46174,N_44389,N_42808);
or U46175 (N_46175,N_43075,N_44639);
nand U46176 (N_46176,N_43474,N_42966);
xor U46177 (N_46177,N_44810,N_43824);
nand U46178 (N_46178,N_43063,N_43949);
xnor U46179 (N_46179,N_43476,N_44017);
nand U46180 (N_46180,N_42682,N_42665);
nor U46181 (N_46181,N_42934,N_42998);
nand U46182 (N_46182,N_43292,N_43691);
xor U46183 (N_46183,N_43199,N_42798);
or U46184 (N_46184,N_44317,N_44082);
and U46185 (N_46185,N_44998,N_43470);
or U46186 (N_46186,N_44195,N_43412);
or U46187 (N_46187,N_43336,N_44592);
or U46188 (N_46188,N_44182,N_42668);
nor U46189 (N_46189,N_44063,N_42535);
and U46190 (N_46190,N_42805,N_43325);
nor U46191 (N_46191,N_42604,N_43310);
and U46192 (N_46192,N_43026,N_42513);
xnor U46193 (N_46193,N_43386,N_42603);
and U46194 (N_46194,N_44460,N_43897);
nand U46195 (N_46195,N_43077,N_43898);
or U46196 (N_46196,N_44629,N_44455);
xor U46197 (N_46197,N_43734,N_43065);
xnor U46198 (N_46198,N_44836,N_42562);
or U46199 (N_46199,N_43142,N_43963);
nor U46200 (N_46200,N_43186,N_44196);
and U46201 (N_46201,N_42577,N_44721);
nand U46202 (N_46202,N_43086,N_44921);
and U46203 (N_46203,N_42538,N_44992);
xor U46204 (N_46204,N_44858,N_43349);
and U46205 (N_46205,N_43242,N_43721);
nand U46206 (N_46206,N_43820,N_42772);
nor U46207 (N_46207,N_43641,N_44875);
xnor U46208 (N_46208,N_44707,N_43555);
or U46209 (N_46209,N_44220,N_43137);
or U46210 (N_46210,N_43237,N_42673);
xnor U46211 (N_46211,N_42537,N_44393);
or U46212 (N_46212,N_44883,N_43163);
nor U46213 (N_46213,N_42920,N_42536);
xnor U46214 (N_46214,N_43708,N_44774);
nand U46215 (N_46215,N_44112,N_43354);
and U46216 (N_46216,N_44829,N_43062);
nor U46217 (N_46217,N_43341,N_42795);
and U46218 (N_46218,N_44128,N_43300);
and U46219 (N_46219,N_44956,N_44008);
nor U46220 (N_46220,N_42834,N_43283);
and U46221 (N_46221,N_44572,N_43204);
nand U46222 (N_46222,N_42907,N_44831);
and U46223 (N_46223,N_44408,N_44255);
nand U46224 (N_46224,N_42747,N_44144);
or U46225 (N_46225,N_43259,N_43558);
or U46226 (N_46226,N_44409,N_42664);
and U46227 (N_46227,N_44835,N_43628);
nor U46228 (N_46228,N_44046,N_44330);
nand U46229 (N_46229,N_43314,N_44954);
or U46230 (N_46230,N_43912,N_44775);
and U46231 (N_46231,N_43170,N_44886);
xor U46232 (N_46232,N_43643,N_42608);
nor U46233 (N_46233,N_43571,N_44761);
xor U46234 (N_46234,N_43619,N_44177);
nand U46235 (N_46235,N_43374,N_44923);
or U46236 (N_46236,N_43038,N_43559);
xor U46237 (N_46237,N_43780,N_44520);
xnor U46238 (N_46238,N_43272,N_44626);
nor U46239 (N_46239,N_44464,N_42655);
and U46240 (N_46240,N_42662,N_42597);
and U46241 (N_46241,N_42509,N_42549);
xnor U46242 (N_46242,N_44111,N_43598);
or U46243 (N_46243,N_43133,N_43174);
xnor U46244 (N_46244,N_43804,N_43047);
and U46245 (N_46245,N_44104,N_42794);
or U46246 (N_46246,N_44933,N_43173);
or U46247 (N_46247,N_43481,N_42506);
nor U46248 (N_46248,N_44689,N_44479);
xnor U46249 (N_46249,N_43713,N_43688);
nor U46250 (N_46250,N_44858,N_43055);
or U46251 (N_46251,N_42516,N_44050);
nor U46252 (N_46252,N_44420,N_44581);
nor U46253 (N_46253,N_42924,N_44521);
nand U46254 (N_46254,N_44567,N_43357);
nand U46255 (N_46255,N_44924,N_42643);
nor U46256 (N_46256,N_44747,N_43468);
nor U46257 (N_46257,N_43132,N_44879);
or U46258 (N_46258,N_43838,N_43026);
xor U46259 (N_46259,N_42830,N_42789);
nand U46260 (N_46260,N_44481,N_42989);
nand U46261 (N_46261,N_43013,N_42693);
nand U46262 (N_46262,N_43810,N_43184);
or U46263 (N_46263,N_44862,N_44271);
xor U46264 (N_46264,N_43527,N_42658);
xor U46265 (N_46265,N_42572,N_43213);
and U46266 (N_46266,N_43872,N_43666);
nor U46267 (N_46267,N_42819,N_42941);
and U46268 (N_46268,N_43535,N_44571);
and U46269 (N_46269,N_43481,N_42837);
and U46270 (N_46270,N_43854,N_42636);
xor U46271 (N_46271,N_44645,N_44890);
xor U46272 (N_46272,N_44773,N_43126);
nand U46273 (N_46273,N_42582,N_44818);
xnor U46274 (N_46274,N_43633,N_43014);
nor U46275 (N_46275,N_42550,N_43801);
nor U46276 (N_46276,N_43712,N_42884);
and U46277 (N_46277,N_43954,N_43376);
nand U46278 (N_46278,N_43939,N_42990);
nor U46279 (N_46279,N_44725,N_43046);
and U46280 (N_46280,N_43397,N_43492);
and U46281 (N_46281,N_44842,N_42552);
or U46282 (N_46282,N_42515,N_43037);
nand U46283 (N_46283,N_44272,N_42866);
nand U46284 (N_46284,N_43941,N_44981);
or U46285 (N_46285,N_43786,N_43490);
nor U46286 (N_46286,N_42510,N_44132);
xnor U46287 (N_46287,N_44604,N_44770);
nor U46288 (N_46288,N_43710,N_43042);
nor U46289 (N_46289,N_44153,N_43008);
or U46290 (N_46290,N_42806,N_44209);
nand U46291 (N_46291,N_44735,N_44086);
and U46292 (N_46292,N_44864,N_43156);
nand U46293 (N_46293,N_42875,N_42663);
xnor U46294 (N_46294,N_43946,N_43793);
nand U46295 (N_46295,N_44185,N_43892);
or U46296 (N_46296,N_44223,N_44077);
or U46297 (N_46297,N_44426,N_42753);
or U46298 (N_46298,N_42827,N_44295);
xor U46299 (N_46299,N_43287,N_43696);
nor U46300 (N_46300,N_44184,N_44354);
nand U46301 (N_46301,N_43193,N_43377);
xor U46302 (N_46302,N_43794,N_43995);
nor U46303 (N_46303,N_43530,N_42946);
xor U46304 (N_46304,N_44794,N_43799);
nor U46305 (N_46305,N_43651,N_44541);
and U46306 (N_46306,N_42908,N_42653);
nor U46307 (N_46307,N_42999,N_44833);
and U46308 (N_46308,N_43935,N_44373);
nor U46309 (N_46309,N_43543,N_44904);
nor U46310 (N_46310,N_44940,N_43511);
xnor U46311 (N_46311,N_42827,N_44966);
and U46312 (N_46312,N_42562,N_44190);
xor U46313 (N_46313,N_43336,N_42614);
xor U46314 (N_46314,N_43980,N_42898);
xnor U46315 (N_46315,N_44812,N_44172);
nor U46316 (N_46316,N_43933,N_42918);
xor U46317 (N_46317,N_44456,N_42515);
and U46318 (N_46318,N_44609,N_42722);
nand U46319 (N_46319,N_43271,N_44081);
nor U46320 (N_46320,N_43665,N_44469);
nor U46321 (N_46321,N_43558,N_44249);
nor U46322 (N_46322,N_43861,N_42762);
nor U46323 (N_46323,N_44339,N_42773);
nor U46324 (N_46324,N_44034,N_43210);
nor U46325 (N_46325,N_44564,N_42822);
xnor U46326 (N_46326,N_44049,N_44417);
xnor U46327 (N_46327,N_42758,N_43852);
xor U46328 (N_46328,N_44320,N_43906);
and U46329 (N_46329,N_42503,N_44739);
xnor U46330 (N_46330,N_42922,N_43928);
xor U46331 (N_46331,N_42779,N_44844);
nor U46332 (N_46332,N_43338,N_43485);
or U46333 (N_46333,N_44210,N_44241);
xor U46334 (N_46334,N_44914,N_44487);
nor U46335 (N_46335,N_43501,N_44160);
or U46336 (N_46336,N_44100,N_43568);
nand U46337 (N_46337,N_43556,N_42941);
xor U46338 (N_46338,N_44558,N_42794);
xor U46339 (N_46339,N_44289,N_43294);
or U46340 (N_46340,N_44882,N_43751);
nand U46341 (N_46341,N_43690,N_44680);
nand U46342 (N_46342,N_43800,N_43883);
nand U46343 (N_46343,N_42760,N_42876);
nor U46344 (N_46344,N_43451,N_44159);
xor U46345 (N_46345,N_44924,N_43558);
xnor U46346 (N_46346,N_43890,N_44630);
nor U46347 (N_46347,N_44801,N_43111);
xor U46348 (N_46348,N_42519,N_42876);
nand U46349 (N_46349,N_42625,N_43175);
or U46350 (N_46350,N_44609,N_43111);
and U46351 (N_46351,N_43103,N_43869);
or U46352 (N_46352,N_44532,N_43269);
or U46353 (N_46353,N_42639,N_44432);
nand U46354 (N_46354,N_43552,N_43717);
xnor U46355 (N_46355,N_44287,N_44387);
nand U46356 (N_46356,N_44248,N_43551);
nand U46357 (N_46357,N_44529,N_43872);
or U46358 (N_46358,N_44877,N_44136);
nor U46359 (N_46359,N_44511,N_44717);
nand U46360 (N_46360,N_42859,N_43783);
and U46361 (N_46361,N_44217,N_44555);
or U46362 (N_46362,N_43319,N_44477);
xor U46363 (N_46363,N_43967,N_43250);
or U46364 (N_46364,N_44176,N_43092);
nand U46365 (N_46365,N_43612,N_44598);
nor U46366 (N_46366,N_43529,N_43533);
and U46367 (N_46367,N_44233,N_44777);
xor U46368 (N_46368,N_43829,N_43629);
nor U46369 (N_46369,N_42536,N_43915);
nor U46370 (N_46370,N_42806,N_43346);
xor U46371 (N_46371,N_42707,N_44893);
nor U46372 (N_46372,N_43027,N_44328);
or U46373 (N_46373,N_42842,N_43589);
or U46374 (N_46374,N_42532,N_44014);
and U46375 (N_46375,N_43330,N_44168);
nor U46376 (N_46376,N_43900,N_42700);
or U46377 (N_46377,N_43071,N_44993);
or U46378 (N_46378,N_43410,N_43497);
and U46379 (N_46379,N_44458,N_43472);
nand U46380 (N_46380,N_43538,N_44416);
nor U46381 (N_46381,N_42742,N_43491);
and U46382 (N_46382,N_43569,N_43425);
nor U46383 (N_46383,N_42507,N_44725);
or U46384 (N_46384,N_43006,N_43623);
xor U46385 (N_46385,N_44558,N_43073);
nand U46386 (N_46386,N_44101,N_44330);
or U46387 (N_46387,N_43446,N_43376);
and U46388 (N_46388,N_43868,N_42637);
nor U46389 (N_46389,N_44021,N_44878);
nand U46390 (N_46390,N_44615,N_44634);
nor U46391 (N_46391,N_44182,N_43234);
nand U46392 (N_46392,N_44543,N_43551);
nand U46393 (N_46393,N_44157,N_44862);
nand U46394 (N_46394,N_43082,N_44773);
or U46395 (N_46395,N_44897,N_42669);
nand U46396 (N_46396,N_43168,N_43204);
nor U46397 (N_46397,N_43030,N_44719);
xor U46398 (N_46398,N_42549,N_44858);
nor U46399 (N_46399,N_44359,N_43457);
or U46400 (N_46400,N_43143,N_42857);
nor U46401 (N_46401,N_44772,N_43131);
xor U46402 (N_46402,N_42557,N_42696);
nor U46403 (N_46403,N_43781,N_44762);
xor U46404 (N_46404,N_43074,N_43975);
and U46405 (N_46405,N_44645,N_42666);
nor U46406 (N_46406,N_44055,N_43155);
xnor U46407 (N_46407,N_43340,N_42777);
xnor U46408 (N_46408,N_43627,N_44189);
and U46409 (N_46409,N_44707,N_42615);
nor U46410 (N_46410,N_43488,N_43385);
and U46411 (N_46411,N_44626,N_44084);
and U46412 (N_46412,N_44763,N_43419);
nor U46413 (N_46413,N_44168,N_43085);
nand U46414 (N_46414,N_43619,N_43258);
nand U46415 (N_46415,N_42858,N_43498);
nor U46416 (N_46416,N_42529,N_42867);
and U46417 (N_46417,N_44689,N_43298);
and U46418 (N_46418,N_43731,N_44382);
and U46419 (N_46419,N_43275,N_44638);
and U46420 (N_46420,N_43177,N_44839);
nor U46421 (N_46421,N_44922,N_44443);
and U46422 (N_46422,N_43037,N_44596);
nor U46423 (N_46423,N_42805,N_43413);
and U46424 (N_46424,N_43531,N_44895);
nand U46425 (N_46425,N_43170,N_44368);
and U46426 (N_46426,N_43841,N_42957);
and U46427 (N_46427,N_44836,N_43169);
or U46428 (N_46428,N_44257,N_44276);
and U46429 (N_46429,N_44646,N_44410);
nor U46430 (N_46430,N_43886,N_42895);
xor U46431 (N_46431,N_43183,N_42930);
or U46432 (N_46432,N_43957,N_44912);
or U46433 (N_46433,N_43145,N_42985);
and U46434 (N_46434,N_43438,N_44482);
xnor U46435 (N_46435,N_44089,N_43113);
or U46436 (N_46436,N_43264,N_43625);
nor U46437 (N_46437,N_44994,N_44290);
xnor U46438 (N_46438,N_43079,N_43948);
or U46439 (N_46439,N_44279,N_44852);
nand U46440 (N_46440,N_44647,N_43692);
xnor U46441 (N_46441,N_44582,N_44387);
and U46442 (N_46442,N_42977,N_43654);
and U46443 (N_46443,N_43245,N_42717);
nand U46444 (N_46444,N_44422,N_43163);
nand U46445 (N_46445,N_44442,N_43158);
or U46446 (N_46446,N_42931,N_44056);
nor U46447 (N_46447,N_43904,N_43231);
nand U46448 (N_46448,N_44080,N_43124);
nor U46449 (N_46449,N_44181,N_42868);
xnor U46450 (N_46450,N_43698,N_42783);
nand U46451 (N_46451,N_43140,N_44206);
nor U46452 (N_46452,N_42906,N_42698);
nand U46453 (N_46453,N_44294,N_44767);
xor U46454 (N_46454,N_43656,N_42638);
or U46455 (N_46455,N_42921,N_43965);
and U46456 (N_46456,N_43396,N_44783);
nor U46457 (N_46457,N_43846,N_44752);
xor U46458 (N_46458,N_43905,N_44856);
and U46459 (N_46459,N_43582,N_44263);
or U46460 (N_46460,N_44697,N_43391);
or U46461 (N_46461,N_42618,N_44868);
xor U46462 (N_46462,N_44017,N_43255);
nand U46463 (N_46463,N_44326,N_44833);
nor U46464 (N_46464,N_44322,N_42670);
and U46465 (N_46465,N_42612,N_42603);
xor U46466 (N_46466,N_43438,N_43191);
nand U46467 (N_46467,N_44081,N_43526);
nor U46468 (N_46468,N_43940,N_44018);
nor U46469 (N_46469,N_43311,N_44588);
and U46470 (N_46470,N_43909,N_42811);
xnor U46471 (N_46471,N_44475,N_43900);
xor U46472 (N_46472,N_43068,N_43138);
nor U46473 (N_46473,N_43677,N_43702);
nor U46474 (N_46474,N_43964,N_43026);
nor U46475 (N_46475,N_44019,N_44136);
or U46476 (N_46476,N_44866,N_44366);
xor U46477 (N_46477,N_44023,N_42698);
xor U46478 (N_46478,N_44686,N_43366);
nor U46479 (N_46479,N_43601,N_43345);
and U46480 (N_46480,N_43485,N_43845);
nor U46481 (N_46481,N_43324,N_44719);
or U46482 (N_46482,N_42726,N_44780);
or U46483 (N_46483,N_43468,N_43896);
or U46484 (N_46484,N_44752,N_44071);
xor U46485 (N_46485,N_42655,N_44164);
nor U46486 (N_46486,N_44028,N_42726);
nand U46487 (N_46487,N_43224,N_43730);
and U46488 (N_46488,N_42861,N_43674);
xor U46489 (N_46489,N_43289,N_42995);
and U46490 (N_46490,N_43035,N_43819);
nand U46491 (N_46491,N_43773,N_43683);
nor U46492 (N_46492,N_43609,N_44149);
nor U46493 (N_46493,N_43809,N_42515);
nand U46494 (N_46494,N_43246,N_43942);
or U46495 (N_46495,N_43957,N_43812);
nor U46496 (N_46496,N_44013,N_42600);
and U46497 (N_46497,N_43335,N_42577);
xnor U46498 (N_46498,N_44402,N_44971);
xnor U46499 (N_46499,N_44912,N_44797);
and U46500 (N_46500,N_44987,N_43065);
or U46501 (N_46501,N_43634,N_43223);
and U46502 (N_46502,N_44491,N_43538);
and U46503 (N_46503,N_42795,N_44667);
xor U46504 (N_46504,N_44519,N_44186);
and U46505 (N_46505,N_43576,N_43213);
nor U46506 (N_46506,N_42506,N_44206);
nand U46507 (N_46507,N_44765,N_43529);
or U46508 (N_46508,N_43077,N_42767);
nand U46509 (N_46509,N_42614,N_42615);
and U46510 (N_46510,N_42687,N_43192);
or U46511 (N_46511,N_44622,N_43292);
nor U46512 (N_46512,N_44963,N_43203);
nand U46513 (N_46513,N_44612,N_43317);
nand U46514 (N_46514,N_43498,N_44511);
or U46515 (N_46515,N_44274,N_42605);
xnor U46516 (N_46516,N_44862,N_44825);
xor U46517 (N_46517,N_43598,N_42521);
xor U46518 (N_46518,N_43327,N_44470);
xor U46519 (N_46519,N_43302,N_44853);
and U46520 (N_46520,N_44820,N_42950);
and U46521 (N_46521,N_44283,N_42970);
nor U46522 (N_46522,N_42939,N_44643);
xnor U46523 (N_46523,N_43860,N_44572);
nor U46524 (N_46524,N_44034,N_42907);
nor U46525 (N_46525,N_44760,N_43894);
or U46526 (N_46526,N_43950,N_43927);
or U46527 (N_46527,N_42522,N_43403);
nand U46528 (N_46528,N_43331,N_43270);
or U46529 (N_46529,N_44710,N_43112);
or U46530 (N_46530,N_42969,N_43716);
nand U46531 (N_46531,N_42857,N_42601);
or U46532 (N_46532,N_42501,N_44048);
or U46533 (N_46533,N_44085,N_44304);
nand U46534 (N_46534,N_43950,N_42939);
or U46535 (N_46535,N_44412,N_43896);
nor U46536 (N_46536,N_42964,N_43744);
or U46537 (N_46537,N_43303,N_42954);
or U46538 (N_46538,N_43505,N_43339);
and U46539 (N_46539,N_44603,N_43072);
and U46540 (N_46540,N_42862,N_44328);
or U46541 (N_46541,N_43353,N_44437);
nand U46542 (N_46542,N_42817,N_43908);
nand U46543 (N_46543,N_44879,N_43239);
nand U46544 (N_46544,N_43343,N_43248);
or U46545 (N_46545,N_43059,N_43226);
and U46546 (N_46546,N_43699,N_42964);
and U46547 (N_46547,N_42658,N_42642);
and U46548 (N_46548,N_44064,N_43157);
and U46549 (N_46549,N_44244,N_42536);
nand U46550 (N_46550,N_43792,N_44134);
nor U46551 (N_46551,N_44612,N_43146);
xor U46552 (N_46552,N_42870,N_44457);
and U46553 (N_46553,N_42621,N_43132);
and U46554 (N_46554,N_43523,N_42796);
xor U46555 (N_46555,N_43991,N_44939);
or U46556 (N_46556,N_44035,N_43240);
or U46557 (N_46557,N_44390,N_44140);
and U46558 (N_46558,N_43637,N_44644);
or U46559 (N_46559,N_44497,N_43056);
or U46560 (N_46560,N_44240,N_42754);
xor U46561 (N_46561,N_42979,N_44806);
nor U46562 (N_46562,N_43028,N_44826);
nor U46563 (N_46563,N_43010,N_43548);
xor U46564 (N_46564,N_43459,N_44912);
or U46565 (N_46565,N_42738,N_44685);
nand U46566 (N_46566,N_42864,N_44991);
or U46567 (N_46567,N_44339,N_43768);
or U46568 (N_46568,N_44888,N_43270);
xor U46569 (N_46569,N_43526,N_43447);
xnor U46570 (N_46570,N_42590,N_44552);
nand U46571 (N_46571,N_42820,N_44944);
or U46572 (N_46572,N_42654,N_42835);
and U46573 (N_46573,N_42549,N_44975);
nor U46574 (N_46574,N_42547,N_43520);
nor U46575 (N_46575,N_43621,N_44485);
nand U46576 (N_46576,N_43888,N_43385);
nand U46577 (N_46577,N_44156,N_43899);
nand U46578 (N_46578,N_43389,N_43146);
nor U46579 (N_46579,N_43554,N_44016);
nand U46580 (N_46580,N_43413,N_42669);
nand U46581 (N_46581,N_44902,N_44384);
xor U46582 (N_46582,N_43776,N_43424);
xnor U46583 (N_46583,N_44457,N_42729);
and U46584 (N_46584,N_43060,N_42716);
nand U46585 (N_46585,N_44859,N_43462);
nand U46586 (N_46586,N_44662,N_44778);
nand U46587 (N_46587,N_44403,N_43673);
nand U46588 (N_46588,N_43488,N_43245);
nor U46589 (N_46589,N_44971,N_44867);
and U46590 (N_46590,N_44134,N_42815);
and U46591 (N_46591,N_42767,N_44494);
nor U46592 (N_46592,N_43148,N_42996);
and U46593 (N_46593,N_42735,N_43075);
nand U46594 (N_46594,N_42547,N_42505);
nand U46595 (N_46595,N_43832,N_43203);
or U46596 (N_46596,N_43665,N_44450);
and U46597 (N_46597,N_43312,N_43537);
and U46598 (N_46598,N_44285,N_43967);
or U46599 (N_46599,N_42887,N_43063);
and U46600 (N_46600,N_43620,N_43193);
nand U46601 (N_46601,N_42625,N_42673);
or U46602 (N_46602,N_43307,N_44395);
nor U46603 (N_46603,N_43500,N_44284);
nor U46604 (N_46604,N_43430,N_43149);
or U46605 (N_46605,N_43407,N_44195);
nor U46606 (N_46606,N_43909,N_43260);
xnor U46607 (N_46607,N_43070,N_42875);
nor U46608 (N_46608,N_44700,N_44801);
nor U46609 (N_46609,N_42748,N_43001);
or U46610 (N_46610,N_44396,N_43185);
and U46611 (N_46611,N_44373,N_44653);
nand U46612 (N_46612,N_44661,N_43654);
nor U46613 (N_46613,N_44279,N_44243);
nand U46614 (N_46614,N_43604,N_42961);
or U46615 (N_46615,N_42720,N_44396);
nand U46616 (N_46616,N_44626,N_43138);
nor U46617 (N_46617,N_44305,N_42538);
or U46618 (N_46618,N_43333,N_42565);
nand U46619 (N_46619,N_43084,N_44719);
nor U46620 (N_46620,N_42611,N_44351);
nor U46621 (N_46621,N_43263,N_43616);
nand U46622 (N_46622,N_44196,N_44259);
xnor U46623 (N_46623,N_43345,N_44482);
xor U46624 (N_46624,N_43528,N_42701);
and U46625 (N_46625,N_44477,N_44432);
or U46626 (N_46626,N_42754,N_44602);
xor U46627 (N_46627,N_43964,N_44028);
nand U46628 (N_46628,N_43986,N_44783);
xnor U46629 (N_46629,N_42637,N_44134);
nor U46630 (N_46630,N_43882,N_43131);
nor U46631 (N_46631,N_44538,N_44700);
nand U46632 (N_46632,N_44649,N_43180);
or U46633 (N_46633,N_44967,N_43938);
nor U46634 (N_46634,N_42847,N_42722);
and U46635 (N_46635,N_43752,N_43673);
and U46636 (N_46636,N_42647,N_42832);
nand U46637 (N_46637,N_43817,N_43296);
nor U46638 (N_46638,N_44047,N_43662);
nor U46639 (N_46639,N_43176,N_43607);
nand U46640 (N_46640,N_44491,N_42804);
xnor U46641 (N_46641,N_43686,N_44869);
nor U46642 (N_46642,N_44455,N_43438);
and U46643 (N_46643,N_43440,N_43420);
or U46644 (N_46644,N_42956,N_44964);
and U46645 (N_46645,N_43643,N_44589);
nand U46646 (N_46646,N_43391,N_42684);
and U46647 (N_46647,N_43069,N_43847);
xnor U46648 (N_46648,N_44348,N_44048);
and U46649 (N_46649,N_44211,N_44952);
nor U46650 (N_46650,N_44439,N_44584);
nand U46651 (N_46651,N_42670,N_44016);
nor U46652 (N_46652,N_43972,N_43726);
xnor U46653 (N_46653,N_43066,N_44882);
nand U46654 (N_46654,N_44228,N_44042);
or U46655 (N_46655,N_44009,N_44400);
nand U46656 (N_46656,N_44306,N_43254);
nor U46657 (N_46657,N_44342,N_42737);
nand U46658 (N_46658,N_44995,N_44018);
and U46659 (N_46659,N_42694,N_43386);
xnor U46660 (N_46660,N_44742,N_44886);
nand U46661 (N_46661,N_43524,N_44532);
nor U46662 (N_46662,N_44884,N_43378);
nor U46663 (N_46663,N_44361,N_43031);
and U46664 (N_46664,N_43066,N_44422);
xnor U46665 (N_46665,N_43923,N_42972);
nor U46666 (N_46666,N_43889,N_44763);
and U46667 (N_46667,N_43160,N_44561);
or U46668 (N_46668,N_42655,N_43060);
or U46669 (N_46669,N_44091,N_42845);
nand U46670 (N_46670,N_44999,N_43788);
nor U46671 (N_46671,N_42705,N_44312);
nand U46672 (N_46672,N_43001,N_42616);
nand U46673 (N_46673,N_44313,N_43630);
or U46674 (N_46674,N_43480,N_44757);
or U46675 (N_46675,N_44474,N_44704);
or U46676 (N_46676,N_44031,N_43320);
nor U46677 (N_46677,N_44073,N_44032);
and U46678 (N_46678,N_43358,N_44073);
or U46679 (N_46679,N_44978,N_42528);
nand U46680 (N_46680,N_43810,N_44052);
nor U46681 (N_46681,N_44961,N_43876);
xor U46682 (N_46682,N_43070,N_44509);
nor U46683 (N_46683,N_44868,N_44967);
nor U46684 (N_46684,N_42937,N_42683);
or U46685 (N_46685,N_44606,N_42904);
and U46686 (N_46686,N_43390,N_43219);
nand U46687 (N_46687,N_43635,N_43514);
nor U46688 (N_46688,N_42694,N_43437);
and U46689 (N_46689,N_44454,N_44437);
nor U46690 (N_46690,N_42790,N_43696);
nand U46691 (N_46691,N_44620,N_44791);
xor U46692 (N_46692,N_44130,N_44876);
and U46693 (N_46693,N_43441,N_44702);
nand U46694 (N_46694,N_42663,N_43436);
xor U46695 (N_46695,N_43311,N_42721);
and U46696 (N_46696,N_43427,N_43912);
nand U46697 (N_46697,N_42544,N_42903);
xor U46698 (N_46698,N_43257,N_43423);
nand U46699 (N_46699,N_43757,N_44811);
or U46700 (N_46700,N_44229,N_44708);
or U46701 (N_46701,N_42721,N_44250);
and U46702 (N_46702,N_44204,N_44379);
and U46703 (N_46703,N_43183,N_42603);
xnor U46704 (N_46704,N_44417,N_44143);
or U46705 (N_46705,N_44165,N_44571);
nor U46706 (N_46706,N_43953,N_43138);
or U46707 (N_46707,N_43702,N_44088);
xor U46708 (N_46708,N_42701,N_42502);
and U46709 (N_46709,N_43351,N_42505);
nand U46710 (N_46710,N_43844,N_44711);
xor U46711 (N_46711,N_42510,N_43504);
xnor U46712 (N_46712,N_42563,N_44189);
nand U46713 (N_46713,N_43562,N_43330);
and U46714 (N_46714,N_44752,N_44228);
nand U46715 (N_46715,N_43827,N_43296);
xor U46716 (N_46716,N_43487,N_44634);
xnor U46717 (N_46717,N_43915,N_44876);
xor U46718 (N_46718,N_44689,N_43965);
xnor U46719 (N_46719,N_42553,N_44582);
nand U46720 (N_46720,N_43070,N_43019);
and U46721 (N_46721,N_44679,N_44733);
nor U46722 (N_46722,N_42772,N_42573);
nor U46723 (N_46723,N_44055,N_44865);
nor U46724 (N_46724,N_42854,N_43053);
xnor U46725 (N_46725,N_42983,N_44901);
nand U46726 (N_46726,N_44340,N_44624);
or U46727 (N_46727,N_44876,N_42871);
nand U46728 (N_46728,N_43846,N_42569);
or U46729 (N_46729,N_43162,N_44247);
xor U46730 (N_46730,N_43201,N_43937);
and U46731 (N_46731,N_43861,N_44805);
and U46732 (N_46732,N_43454,N_43695);
nand U46733 (N_46733,N_44783,N_44808);
nand U46734 (N_46734,N_44253,N_44278);
nor U46735 (N_46735,N_44110,N_43816);
or U46736 (N_46736,N_44948,N_42802);
and U46737 (N_46737,N_44606,N_42809);
nor U46738 (N_46738,N_43734,N_43172);
xor U46739 (N_46739,N_44798,N_43694);
nand U46740 (N_46740,N_43611,N_44704);
nand U46741 (N_46741,N_43594,N_42864);
nor U46742 (N_46742,N_43948,N_44224);
nor U46743 (N_46743,N_42640,N_43053);
xnor U46744 (N_46744,N_43984,N_42684);
xnor U46745 (N_46745,N_43259,N_43542);
and U46746 (N_46746,N_43835,N_43094);
nor U46747 (N_46747,N_44918,N_43997);
nand U46748 (N_46748,N_44539,N_44459);
or U46749 (N_46749,N_43222,N_44198);
and U46750 (N_46750,N_43608,N_44624);
nand U46751 (N_46751,N_44247,N_43107);
or U46752 (N_46752,N_43456,N_42989);
xnor U46753 (N_46753,N_44701,N_44285);
nor U46754 (N_46754,N_43091,N_44957);
and U46755 (N_46755,N_43459,N_42717);
nand U46756 (N_46756,N_42734,N_43243);
xor U46757 (N_46757,N_43300,N_43340);
nand U46758 (N_46758,N_43054,N_42850);
and U46759 (N_46759,N_43280,N_43639);
and U46760 (N_46760,N_42703,N_43160);
or U46761 (N_46761,N_44781,N_43156);
xnor U46762 (N_46762,N_43607,N_44165);
or U46763 (N_46763,N_43912,N_44054);
and U46764 (N_46764,N_44405,N_43324);
nand U46765 (N_46765,N_43490,N_43224);
and U46766 (N_46766,N_43701,N_43764);
nor U46767 (N_46767,N_42696,N_42898);
and U46768 (N_46768,N_42534,N_42790);
nor U46769 (N_46769,N_44756,N_44451);
or U46770 (N_46770,N_44486,N_42902);
and U46771 (N_46771,N_43294,N_42763);
nand U46772 (N_46772,N_43713,N_44484);
and U46773 (N_46773,N_44241,N_43928);
nand U46774 (N_46774,N_44301,N_44442);
or U46775 (N_46775,N_42693,N_44143);
nand U46776 (N_46776,N_44511,N_44162);
and U46777 (N_46777,N_44009,N_44743);
nor U46778 (N_46778,N_44261,N_43717);
xor U46779 (N_46779,N_43280,N_43981);
nor U46780 (N_46780,N_43506,N_44378);
xnor U46781 (N_46781,N_43063,N_42644);
and U46782 (N_46782,N_43502,N_43835);
and U46783 (N_46783,N_42945,N_44123);
and U46784 (N_46784,N_42885,N_42938);
xor U46785 (N_46785,N_43521,N_44619);
or U46786 (N_46786,N_42621,N_42632);
xor U46787 (N_46787,N_42727,N_42518);
nor U46788 (N_46788,N_43433,N_44409);
xor U46789 (N_46789,N_44106,N_44996);
and U46790 (N_46790,N_44672,N_43098);
or U46791 (N_46791,N_42675,N_42635);
and U46792 (N_46792,N_44842,N_44657);
nand U46793 (N_46793,N_44427,N_43830);
nand U46794 (N_46794,N_43606,N_44353);
nor U46795 (N_46795,N_43797,N_43847);
or U46796 (N_46796,N_44502,N_44411);
and U46797 (N_46797,N_44316,N_42656);
and U46798 (N_46798,N_43677,N_43164);
nor U46799 (N_46799,N_44923,N_42750);
nor U46800 (N_46800,N_43571,N_42889);
and U46801 (N_46801,N_42853,N_44353);
and U46802 (N_46802,N_43858,N_44715);
or U46803 (N_46803,N_44395,N_44024);
and U46804 (N_46804,N_44981,N_44177);
and U46805 (N_46805,N_42796,N_42934);
or U46806 (N_46806,N_44052,N_43019);
nor U46807 (N_46807,N_44570,N_43130);
nor U46808 (N_46808,N_44532,N_44642);
nand U46809 (N_46809,N_42595,N_43855);
nor U46810 (N_46810,N_44821,N_43396);
and U46811 (N_46811,N_44747,N_43639);
and U46812 (N_46812,N_43014,N_44740);
nand U46813 (N_46813,N_42853,N_42907);
or U46814 (N_46814,N_43931,N_43536);
nand U46815 (N_46815,N_43752,N_42612);
nand U46816 (N_46816,N_44066,N_43829);
nor U46817 (N_46817,N_42873,N_42792);
xnor U46818 (N_46818,N_44338,N_44688);
or U46819 (N_46819,N_44926,N_44590);
nor U46820 (N_46820,N_44449,N_44954);
xnor U46821 (N_46821,N_43595,N_44375);
and U46822 (N_46822,N_44941,N_44767);
nand U46823 (N_46823,N_44759,N_43259);
nand U46824 (N_46824,N_43778,N_42854);
nor U46825 (N_46825,N_44696,N_44754);
xnor U46826 (N_46826,N_43763,N_43880);
and U46827 (N_46827,N_43867,N_44102);
xnor U46828 (N_46828,N_42671,N_43029);
nor U46829 (N_46829,N_44078,N_43753);
nand U46830 (N_46830,N_42819,N_42935);
nor U46831 (N_46831,N_43243,N_43436);
or U46832 (N_46832,N_43902,N_44101);
nand U46833 (N_46833,N_43079,N_44616);
xnor U46834 (N_46834,N_43184,N_44416);
nor U46835 (N_46835,N_44337,N_43053);
nand U46836 (N_46836,N_43391,N_44749);
and U46837 (N_46837,N_43778,N_44323);
nor U46838 (N_46838,N_43139,N_43710);
nand U46839 (N_46839,N_44008,N_44601);
xnor U46840 (N_46840,N_43531,N_43103);
xor U46841 (N_46841,N_44690,N_43882);
xor U46842 (N_46842,N_44736,N_44053);
nor U46843 (N_46843,N_44579,N_44134);
and U46844 (N_46844,N_43186,N_43820);
or U46845 (N_46845,N_42788,N_43018);
or U46846 (N_46846,N_42821,N_42981);
nor U46847 (N_46847,N_44538,N_43820);
xor U46848 (N_46848,N_42944,N_44312);
nand U46849 (N_46849,N_43281,N_44533);
nand U46850 (N_46850,N_44211,N_44364);
or U46851 (N_46851,N_44714,N_44851);
or U46852 (N_46852,N_42969,N_44447);
or U46853 (N_46853,N_44629,N_42956);
xor U46854 (N_46854,N_43721,N_43860);
or U46855 (N_46855,N_44971,N_44927);
xor U46856 (N_46856,N_43644,N_44776);
nor U46857 (N_46857,N_43941,N_44095);
or U46858 (N_46858,N_43511,N_44876);
or U46859 (N_46859,N_42854,N_43510);
nand U46860 (N_46860,N_44943,N_43950);
nor U46861 (N_46861,N_43349,N_43646);
or U46862 (N_46862,N_43222,N_42538);
nor U46863 (N_46863,N_44777,N_43332);
xor U46864 (N_46864,N_42761,N_43153);
nand U46865 (N_46865,N_43419,N_43868);
or U46866 (N_46866,N_42615,N_43150);
and U46867 (N_46867,N_42648,N_43324);
and U46868 (N_46868,N_44624,N_42575);
and U46869 (N_46869,N_44772,N_44175);
and U46870 (N_46870,N_44878,N_43703);
nand U46871 (N_46871,N_43594,N_42595);
nor U46872 (N_46872,N_43978,N_42553);
or U46873 (N_46873,N_43165,N_43967);
xor U46874 (N_46874,N_44793,N_42686);
nor U46875 (N_46875,N_44168,N_43879);
nor U46876 (N_46876,N_44767,N_44573);
or U46877 (N_46877,N_43927,N_44443);
nand U46878 (N_46878,N_43863,N_42825);
nand U46879 (N_46879,N_43071,N_44148);
nand U46880 (N_46880,N_44386,N_43620);
and U46881 (N_46881,N_43353,N_43432);
nand U46882 (N_46882,N_44322,N_43318);
and U46883 (N_46883,N_42629,N_43318);
nand U46884 (N_46884,N_44008,N_44449);
nand U46885 (N_46885,N_43450,N_44521);
xor U46886 (N_46886,N_42837,N_44446);
xnor U46887 (N_46887,N_42850,N_43665);
xor U46888 (N_46888,N_43243,N_43082);
nand U46889 (N_46889,N_43010,N_42619);
nand U46890 (N_46890,N_44782,N_42661);
nand U46891 (N_46891,N_43176,N_43354);
or U46892 (N_46892,N_43172,N_42940);
or U46893 (N_46893,N_44774,N_44013);
or U46894 (N_46894,N_43210,N_43386);
and U46895 (N_46895,N_43279,N_43019);
or U46896 (N_46896,N_44379,N_42529);
nor U46897 (N_46897,N_44861,N_43680);
and U46898 (N_46898,N_42638,N_42717);
nor U46899 (N_46899,N_43514,N_44108);
or U46900 (N_46900,N_42705,N_44254);
nand U46901 (N_46901,N_43863,N_44653);
nor U46902 (N_46902,N_44739,N_44345);
or U46903 (N_46903,N_43884,N_44189);
nand U46904 (N_46904,N_44684,N_42803);
nor U46905 (N_46905,N_44028,N_43437);
xnor U46906 (N_46906,N_43765,N_44413);
or U46907 (N_46907,N_43433,N_44561);
nand U46908 (N_46908,N_44251,N_43070);
or U46909 (N_46909,N_44062,N_43746);
nor U46910 (N_46910,N_42851,N_42812);
or U46911 (N_46911,N_43345,N_43613);
xor U46912 (N_46912,N_43929,N_43501);
nand U46913 (N_46913,N_43319,N_43662);
and U46914 (N_46914,N_43571,N_42582);
or U46915 (N_46915,N_44450,N_43489);
nor U46916 (N_46916,N_42542,N_43141);
and U46917 (N_46917,N_44053,N_44200);
nand U46918 (N_46918,N_43746,N_43628);
nand U46919 (N_46919,N_44111,N_42947);
or U46920 (N_46920,N_43152,N_42785);
xor U46921 (N_46921,N_43488,N_43758);
nor U46922 (N_46922,N_44152,N_44732);
and U46923 (N_46923,N_42720,N_42571);
nor U46924 (N_46924,N_42626,N_42607);
nor U46925 (N_46925,N_43598,N_43617);
and U46926 (N_46926,N_42738,N_43602);
or U46927 (N_46927,N_43355,N_44389);
or U46928 (N_46928,N_42753,N_42521);
xnor U46929 (N_46929,N_44717,N_44157);
or U46930 (N_46930,N_42598,N_43905);
or U46931 (N_46931,N_44608,N_44737);
nor U46932 (N_46932,N_44856,N_44356);
and U46933 (N_46933,N_44287,N_44010);
xor U46934 (N_46934,N_44598,N_43603);
and U46935 (N_46935,N_44335,N_44211);
and U46936 (N_46936,N_43188,N_42527);
and U46937 (N_46937,N_43878,N_44985);
nand U46938 (N_46938,N_42633,N_43789);
or U46939 (N_46939,N_44579,N_44250);
xor U46940 (N_46940,N_42619,N_43726);
and U46941 (N_46941,N_44019,N_44922);
nor U46942 (N_46942,N_43473,N_43534);
and U46943 (N_46943,N_44257,N_43096);
nand U46944 (N_46944,N_44554,N_42689);
nand U46945 (N_46945,N_43797,N_44893);
nand U46946 (N_46946,N_44719,N_43749);
nor U46947 (N_46947,N_43727,N_42505);
or U46948 (N_46948,N_43721,N_44418);
nor U46949 (N_46949,N_42507,N_44355);
nand U46950 (N_46950,N_44353,N_44825);
and U46951 (N_46951,N_43008,N_42804);
nor U46952 (N_46952,N_44709,N_43457);
xnor U46953 (N_46953,N_43261,N_42861);
xnor U46954 (N_46954,N_44909,N_44008);
nand U46955 (N_46955,N_43412,N_43756);
xnor U46956 (N_46956,N_43352,N_43205);
and U46957 (N_46957,N_44186,N_42660);
nand U46958 (N_46958,N_44009,N_43184);
nand U46959 (N_46959,N_44389,N_43348);
and U46960 (N_46960,N_43341,N_43757);
or U46961 (N_46961,N_43581,N_43635);
nand U46962 (N_46962,N_43539,N_44417);
nor U46963 (N_46963,N_44926,N_43684);
nor U46964 (N_46964,N_43360,N_44170);
nor U46965 (N_46965,N_42978,N_42517);
nor U46966 (N_46966,N_44558,N_43493);
xor U46967 (N_46967,N_44250,N_43119);
nor U46968 (N_46968,N_43278,N_43293);
and U46969 (N_46969,N_44231,N_42977);
nor U46970 (N_46970,N_42562,N_44960);
or U46971 (N_46971,N_43996,N_42814);
xor U46972 (N_46972,N_43338,N_42647);
nor U46973 (N_46973,N_44208,N_43344);
and U46974 (N_46974,N_42630,N_42718);
or U46975 (N_46975,N_43841,N_44748);
or U46976 (N_46976,N_44916,N_44643);
or U46977 (N_46977,N_42670,N_44217);
or U46978 (N_46978,N_43290,N_44003);
xnor U46979 (N_46979,N_43013,N_44448);
and U46980 (N_46980,N_43595,N_42579);
nor U46981 (N_46981,N_44072,N_43893);
nand U46982 (N_46982,N_44974,N_43346);
or U46983 (N_46983,N_43479,N_44622);
or U46984 (N_46984,N_42559,N_44339);
xor U46985 (N_46985,N_43210,N_42780);
nor U46986 (N_46986,N_42658,N_43871);
xnor U46987 (N_46987,N_42815,N_42645);
and U46988 (N_46988,N_43790,N_43357);
and U46989 (N_46989,N_42558,N_44061);
xor U46990 (N_46990,N_43129,N_44250);
xor U46991 (N_46991,N_42542,N_44392);
or U46992 (N_46992,N_43472,N_43377);
and U46993 (N_46993,N_43312,N_44772);
and U46994 (N_46994,N_43966,N_43086);
or U46995 (N_46995,N_43703,N_44582);
nor U46996 (N_46996,N_42892,N_44820);
nand U46997 (N_46997,N_44835,N_43394);
xor U46998 (N_46998,N_43537,N_44345);
or U46999 (N_46999,N_42888,N_43856);
nor U47000 (N_47000,N_43754,N_43296);
nand U47001 (N_47001,N_42681,N_42506);
nor U47002 (N_47002,N_43142,N_43161);
and U47003 (N_47003,N_42977,N_43855);
and U47004 (N_47004,N_43061,N_43535);
nand U47005 (N_47005,N_44058,N_43480);
or U47006 (N_47006,N_44292,N_44609);
or U47007 (N_47007,N_44056,N_42574);
and U47008 (N_47008,N_43982,N_44290);
nor U47009 (N_47009,N_42668,N_44599);
nor U47010 (N_47010,N_44815,N_43826);
and U47011 (N_47011,N_42804,N_43300);
or U47012 (N_47012,N_43211,N_42919);
nor U47013 (N_47013,N_43819,N_43181);
xnor U47014 (N_47014,N_43891,N_43389);
or U47015 (N_47015,N_43589,N_42905);
and U47016 (N_47016,N_43910,N_44338);
nor U47017 (N_47017,N_42664,N_44089);
nor U47018 (N_47018,N_43095,N_43084);
nand U47019 (N_47019,N_44017,N_44708);
nand U47020 (N_47020,N_43111,N_44918);
or U47021 (N_47021,N_44639,N_42582);
and U47022 (N_47022,N_44381,N_43152);
or U47023 (N_47023,N_44419,N_44318);
or U47024 (N_47024,N_43405,N_43051);
nand U47025 (N_47025,N_44153,N_42742);
and U47026 (N_47026,N_44102,N_43235);
xnor U47027 (N_47027,N_43334,N_43363);
nor U47028 (N_47028,N_43325,N_44681);
nor U47029 (N_47029,N_44049,N_44899);
nor U47030 (N_47030,N_43478,N_44504);
or U47031 (N_47031,N_44741,N_44991);
and U47032 (N_47032,N_43955,N_44094);
xnor U47033 (N_47033,N_44575,N_44118);
xnor U47034 (N_47034,N_43952,N_43017);
nor U47035 (N_47035,N_44468,N_43691);
or U47036 (N_47036,N_43667,N_42692);
nand U47037 (N_47037,N_43015,N_43831);
or U47038 (N_47038,N_43146,N_44903);
or U47039 (N_47039,N_42725,N_44205);
nor U47040 (N_47040,N_42702,N_43701);
xnor U47041 (N_47041,N_42618,N_44602);
or U47042 (N_47042,N_43928,N_44595);
or U47043 (N_47043,N_44745,N_42861);
and U47044 (N_47044,N_44694,N_43081);
and U47045 (N_47045,N_43062,N_43719);
nand U47046 (N_47046,N_44226,N_44716);
xnor U47047 (N_47047,N_42738,N_44866);
nand U47048 (N_47048,N_43751,N_44455);
nor U47049 (N_47049,N_43821,N_44991);
and U47050 (N_47050,N_42646,N_44934);
nand U47051 (N_47051,N_43895,N_42851);
or U47052 (N_47052,N_44169,N_42508);
nor U47053 (N_47053,N_42555,N_43450);
nor U47054 (N_47054,N_43480,N_44893);
xnor U47055 (N_47055,N_42860,N_44919);
xor U47056 (N_47056,N_42964,N_44249);
xor U47057 (N_47057,N_42638,N_43817);
and U47058 (N_47058,N_44042,N_44786);
nand U47059 (N_47059,N_44775,N_43173);
xnor U47060 (N_47060,N_43376,N_44157);
xnor U47061 (N_47061,N_44061,N_44661);
nor U47062 (N_47062,N_43626,N_44082);
or U47063 (N_47063,N_44645,N_42664);
or U47064 (N_47064,N_42678,N_42612);
nand U47065 (N_47065,N_44611,N_42665);
xor U47066 (N_47066,N_42789,N_44149);
xor U47067 (N_47067,N_43254,N_44495);
or U47068 (N_47068,N_43284,N_44914);
nor U47069 (N_47069,N_44520,N_43121);
or U47070 (N_47070,N_43345,N_42979);
and U47071 (N_47071,N_44827,N_42955);
xor U47072 (N_47072,N_43934,N_44503);
and U47073 (N_47073,N_43384,N_44566);
and U47074 (N_47074,N_42821,N_42688);
nand U47075 (N_47075,N_42645,N_44902);
or U47076 (N_47076,N_42684,N_43319);
nor U47077 (N_47077,N_43718,N_44975);
nor U47078 (N_47078,N_44143,N_43819);
xnor U47079 (N_47079,N_44323,N_44998);
nor U47080 (N_47080,N_43594,N_42875);
xor U47081 (N_47081,N_44616,N_44383);
nand U47082 (N_47082,N_43783,N_43864);
or U47083 (N_47083,N_42602,N_43918);
nor U47084 (N_47084,N_44062,N_43345);
xor U47085 (N_47085,N_44735,N_43213);
xor U47086 (N_47086,N_44168,N_42521);
and U47087 (N_47087,N_42668,N_43993);
and U47088 (N_47088,N_43338,N_44575);
and U47089 (N_47089,N_44882,N_43143);
nor U47090 (N_47090,N_44035,N_44396);
xor U47091 (N_47091,N_44323,N_43574);
and U47092 (N_47092,N_43710,N_43355);
nor U47093 (N_47093,N_44559,N_43271);
nor U47094 (N_47094,N_43407,N_42662);
and U47095 (N_47095,N_43794,N_43297);
or U47096 (N_47096,N_43854,N_43822);
nand U47097 (N_47097,N_42774,N_44540);
or U47098 (N_47098,N_42586,N_43523);
or U47099 (N_47099,N_44040,N_44882);
nor U47100 (N_47100,N_43538,N_43079);
or U47101 (N_47101,N_42937,N_44435);
nor U47102 (N_47102,N_43988,N_44771);
nor U47103 (N_47103,N_44896,N_43339);
xnor U47104 (N_47104,N_43515,N_43904);
or U47105 (N_47105,N_43360,N_43942);
and U47106 (N_47106,N_43473,N_43730);
nor U47107 (N_47107,N_43178,N_44928);
or U47108 (N_47108,N_43887,N_42984);
nand U47109 (N_47109,N_42679,N_44700);
xnor U47110 (N_47110,N_43209,N_43367);
xnor U47111 (N_47111,N_43082,N_43574);
xor U47112 (N_47112,N_42917,N_43745);
nand U47113 (N_47113,N_42656,N_44504);
nor U47114 (N_47114,N_44625,N_43119);
nor U47115 (N_47115,N_42649,N_44337);
and U47116 (N_47116,N_43244,N_43611);
xor U47117 (N_47117,N_44603,N_43305);
or U47118 (N_47118,N_42878,N_44641);
nand U47119 (N_47119,N_42921,N_44008);
nor U47120 (N_47120,N_44833,N_42540);
xnor U47121 (N_47121,N_42573,N_44965);
nand U47122 (N_47122,N_44629,N_43839);
xnor U47123 (N_47123,N_43421,N_43371);
nor U47124 (N_47124,N_43556,N_42956);
or U47125 (N_47125,N_44557,N_43812);
nor U47126 (N_47126,N_43810,N_43665);
or U47127 (N_47127,N_42735,N_43268);
nor U47128 (N_47128,N_44256,N_44791);
nor U47129 (N_47129,N_44453,N_44912);
xnor U47130 (N_47130,N_43942,N_44325);
or U47131 (N_47131,N_44776,N_43206);
nand U47132 (N_47132,N_44091,N_43647);
and U47133 (N_47133,N_44472,N_43774);
and U47134 (N_47134,N_44486,N_44473);
xnor U47135 (N_47135,N_44523,N_42826);
nor U47136 (N_47136,N_42998,N_44292);
xnor U47137 (N_47137,N_43138,N_44616);
nand U47138 (N_47138,N_44229,N_44328);
xor U47139 (N_47139,N_43176,N_43585);
and U47140 (N_47140,N_42673,N_42913);
xor U47141 (N_47141,N_42717,N_43889);
nand U47142 (N_47142,N_42788,N_42863);
nand U47143 (N_47143,N_44267,N_43445);
nand U47144 (N_47144,N_42876,N_43366);
nand U47145 (N_47145,N_43606,N_44157);
nand U47146 (N_47146,N_43472,N_44288);
or U47147 (N_47147,N_42606,N_43206);
or U47148 (N_47148,N_44934,N_44257);
nor U47149 (N_47149,N_43312,N_42611);
and U47150 (N_47150,N_44466,N_44065);
or U47151 (N_47151,N_44846,N_43251);
nor U47152 (N_47152,N_43149,N_43480);
nand U47153 (N_47153,N_44444,N_42598);
and U47154 (N_47154,N_43865,N_44558);
nor U47155 (N_47155,N_43522,N_43307);
nand U47156 (N_47156,N_43921,N_42821);
and U47157 (N_47157,N_42551,N_44952);
nor U47158 (N_47158,N_44121,N_42827);
and U47159 (N_47159,N_44294,N_43163);
xor U47160 (N_47160,N_44782,N_44995);
or U47161 (N_47161,N_42583,N_44126);
and U47162 (N_47162,N_44569,N_42785);
xnor U47163 (N_47163,N_43367,N_43172);
nand U47164 (N_47164,N_43446,N_43350);
and U47165 (N_47165,N_42763,N_43549);
nor U47166 (N_47166,N_43898,N_43009);
xor U47167 (N_47167,N_42867,N_43530);
or U47168 (N_47168,N_43402,N_44672);
xnor U47169 (N_47169,N_44980,N_44017);
and U47170 (N_47170,N_43301,N_43469);
nor U47171 (N_47171,N_43716,N_43819);
and U47172 (N_47172,N_42980,N_43481);
and U47173 (N_47173,N_43788,N_43760);
nor U47174 (N_47174,N_42512,N_44096);
xnor U47175 (N_47175,N_44647,N_42782);
nand U47176 (N_47176,N_42918,N_44213);
or U47177 (N_47177,N_43312,N_43237);
xor U47178 (N_47178,N_43728,N_42759);
nand U47179 (N_47179,N_44140,N_43624);
or U47180 (N_47180,N_43021,N_44163);
xor U47181 (N_47181,N_42967,N_43577);
and U47182 (N_47182,N_44781,N_43181);
xor U47183 (N_47183,N_44219,N_44714);
and U47184 (N_47184,N_43938,N_43459);
or U47185 (N_47185,N_42580,N_43390);
or U47186 (N_47186,N_44166,N_42898);
nor U47187 (N_47187,N_44053,N_43055);
and U47188 (N_47188,N_44139,N_44660);
and U47189 (N_47189,N_43634,N_43947);
nand U47190 (N_47190,N_43732,N_44256);
and U47191 (N_47191,N_43819,N_42600);
and U47192 (N_47192,N_44925,N_42815);
nand U47193 (N_47193,N_44389,N_44849);
or U47194 (N_47194,N_42918,N_44760);
nor U47195 (N_47195,N_44595,N_43837);
and U47196 (N_47196,N_43542,N_43248);
nor U47197 (N_47197,N_43342,N_43071);
nor U47198 (N_47198,N_43001,N_43017);
and U47199 (N_47199,N_43047,N_43928);
and U47200 (N_47200,N_44457,N_44867);
nand U47201 (N_47201,N_42913,N_44894);
xnor U47202 (N_47202,N_43971,N_44908);
or U47203 (N_47203,N_44552,N_43389);
xor U47204 (N_47204,N_43769,N_43966);
xor U47205 (N_47205,N_44995,N_44974);
nor U47206 (N_47206,N_43515,N_44782);
xnor U47207 (N_47207,N_43724,N_43095);
nand U47208 (N_47208,N_43074,N_43130);
nand U47209 (N_47209,N_43739,N_43777);
nand U47210 (N_47210,N_42988,N_42577);
nand U47211 (N_47211,N_43093,N_44914);
and U47212 (N_47212,N_43887,N_43705);
or U47213 (N_47213,N_44319,N_43447);
xor U47214 (N_47214,N_44388,N_43748);
xor U47215 (N_47215,N_43957,N_44761);
or U47216 (N_47216,N_44047,N_42907);
and U47217 (N_47217,N_43101,N_43875);
nand U47218 (N_47218,N_44324,N_43958);
nand U47219 (N_47219,N_42797,N_43645);
nor U47220 (N_47220,N_43204,N_43115);
nand U47221 (N_47221,N_43291,N_44686);
and U47222 (N_47222,N_43703,N_43713);
nand U47223 (N_47223,N_44330,N_43488);
and U47224 (N_47224,N_43779,N_42738);
xnor U47225 (N_47225,N_43343,N_43783);
and U47226 (N_47226,N_44425,N_42955);
and U47227 (N_47227,N_42682,N_44135);
xor U47228 (N_47228,N_43454,N_42748);
nor U47229 (N_47229,N_44532,N_44109);
nand U47230 (N_47230,N_43691,N_44980);
and U47231 (N_47231,N_44510,N_44981);
nor U47232 (N_47232,N_43911,N_43050);
nor U47233 (N_47233,N_44392,N_42860);
or U47234 (N_47234,N_43008,N_42718);
and U47235 (N_47235,N_44388,N_43761);
nand U47236 (N_47236,N_42926,N_44452);
or U47237 (N_47237,N_43879,N_44395);
and U47238 (N_47238,N_43945,N_44131);
nor U47239 (N_47239,N_44052,N_42932);
xnor U47240 (N_47240,N_44319,N_44938);
nand U47241 (N_47241,N_43515,N_44352);
or U47242 (N_47242,N_43613,N_43831);
nor U47243 (N_47243,N_43181,N_44216);
xnor U47244 (N_47244,N_44251,N_44906);
or U47245 (N_47245,N_44466,N_44431);
nand U47246 (N_47246,N_43752,N_44880);
or U47247 (N_47247,N_44417,N_43892);
nor U47248 (N_47248,N_42831,N_44204);
xnor U47249 (N_47249,N_44234,N_42917);
and U47250 (N_47250,N_44719,N_44458);
or U47251 (N_47251,N_44661,N_43377);
nand U47252 (N_47252,N_43696,N_42756);
nand U47253 (N_47253,N_43417,N_44490);
and U47254 (N_47254,N_43180,N_43652);
or U47255 (N_47255,N_44273,N_43703);
nand U47256 (N_47256,N_44671,N_44774);
or U47257 (N_47257,N_43480,N_44221);
and U47258 (N_47258,N_42829,N_44878);
nand U47259 (N_47259,N_43248,N_43743);
nand U47260 (N_47260,N_42692,N_44556);
xnor U47261 (N_47261,N_43213,N_44721);
nand U47262 (N_47262,N_44799,N_44837);
nor U47263 (N_47263,N_44897,N_44850);
nand U47264 (N_47264,N_44749,N_42783);
and U47265 (N_47265,N_44611,N_43794);
nand U47266 (N_47266,N_44576,N_42523);
nand U47267 (N_47267,N_44945,N_42991);
nor U47268 (N_47268,N_42861,N_42620);
or U47269 (N_47269,N_43841,N_44611);
nand U47270 (N_47270,N_42579,N_42953);
or U47271 (N_47271,N_44454,N_44146);
or U47272 (N_47272,N_44590,N_43561);
and U47273 (N_47273,N_43468,N_42599);
nor U47274 (N_47274,N_43165,N_44540);
nand U47275 (N_47275,N_43739,N_43816);
nor U47276 (N_47276,N_42625,N_44480);
and U47277 (N_47277,N_44108,N_44020);
nand U47278 (N_47278,N_44067,N_43357);
or U47279 (N_47279,N_43323,N_43144);
xnor U47280 (N_47280,N_43253,N_43404);
xnor U47281 (N_47281,N_43027,N_44344);
nand U47282 (N_47282,N_44126,N_44041);
xnor U47283 (N_47283,N_43037,N_42619);
nor U47284 (N_47284,N_44016,N_44713);
nand U47285 (N_47285,N_44957,N_44539);
nand U47286 (N_47286,N_44963,N_44838);
and U47287 (N_47287,N_43775,N_44739);
nor U47288 (N_47288,N_44727,N_44684);
nor U47289 (N_47289,N_44276,N_43437);
nand U47290 (N_47290,N_43189,N_43918);
nor U47291 (N_47291,N_44335,N_43406);
nand U47292 (N_47292,N_43930,N_44936);
xor U47293 (N_47293,N_42905,N_42829);
or U47294 (N_47294,N_43075,N_44883);
or U47295 (N_47295,N_42935,N_43613);
or U47296 (N_47296,N_43958,N_43754);
or U47297 (N_47297,N_44635,N_43397);
nor U47298 (N_47298,N_42866,N_43217);
nor U47299 (N_47299,N_42837,N_44102);
nand U47300 (N_47300,N_44444,N_43767);
nor U47301 (N_47301,N_43713,N_44713);
nand U47302 (N_47302,N_43630,N_43601);
xnor U47303 (N_47303,N_42628,N_44031);
nand U47304 (N_47304,N_43632,N_42700);
or U47305 (N_47305,N_43809,N_44632);
xor U47306 (N_47306,N_43592,N_44090);
xnor U47307 (N_47307,N_44962,N_43779);
and U47308 (N_47308,N_43127,N_43674);
and U47309 (N_47309,N_43417,N_43641);
xor U47310 (N_47310,N_43733,N_44850);
xnor U47311 (N_47311,N_44799,N_43106);
and U47312 (N_47312,N_44870,N_43642);
and U47313 (N_47313,N_42723,N_43740);
or U47314 (N_47314,N_44129,N_44219);
and U47315 (N_47315,N_42794,N_42507);
and U47316 (N_47316,N_42847,N_42863);
or U47317 (N_47317,N_44656,N_43244);
or U47318 (N_47318,N_42792,N_44292);
and U47319 (N_47319,N_43842,N_43819);
nor U47320 (N_47320,N_44710,N_43530);
nand U47321 (N_47321,N_44173,N_43797);
or U47322 (N_47322,N_44119,N_44649);
and U47323 (N_47323,N_44446,N_44130);
xor U47324 (N_47324,N_44290,N_44278);
nor U47325 (N_47325,N_44985,N_44044);
nor U47326 (N_47326,N_44563,N_44803);
and U47327 (N_47327,N_44150,N_42978);
nand U47328 (N_47328,N_42895,N_42804);
and U47329 (N_47329,N_44151,N_43667);
nand U47330 (N_47330,N_43470,N_44997);
nor U47331 (N_47331,N_43571,N_43457);
nand U47332 (N_47332,N_44094,N_44671);
or U47333 (N_47333,N_44894,N_44258);
and U47334 (N_47334,N_44545,N_43096);
nand U47335 (N_47335,N_44550,N_43952);
or U47336 (N_47336,N_44040,N_42555);
xnor U47337 (N_47337,N_43019,N_43254);
nand U47338 (N_47338,N_43626,N_43833);
and U47339 (N_47339,N_43900,N_42870);
xnor U47340 (N_47340,N_43773,N_44137);
or U47341 (N_47341,N_43409,N_44491);
xor U47342 (N_47342,N_43539,N_43722);
and U47343 (N_47343,N_43181,N_44751);
xor U47344 (N_47344,N_43831,N_43661);
and U47345 (N_47345,N_43278,N_42710);
nand U47346 (N_47346,N_44462,N_42942);
or U47347 (N_47347,N_43315,N_44105);
xnor U47348 (N_47348,N_43005,N_44256);
and U47349 (N_47349,N_42927,N_44406);
xnor U47350 (N_47350,N_42604,N_44679);
nand U47351 (N_47351,N_43463,N_42912);
nand U47352 (N_47352,N_44756,N_44953);
xnor U47353 (N_47353,N_43529,N_42843);
nor U47354 (N_47354,N_44969,N_43802);
nor U47355 (N_47355,N_44396,N_44080);
xnor U47356 (N_47356,N_42584,N_42544);
nor U47357 (N_47357,N_42792,N_44835);
nand U47358 (N_47358,N_44457,N_44869);
xnor U47359 (N_47359,N_44126,N_42945);
and U47360 (N_47360,N_43052,N_43204);
xnor U47361 (N_47361,N_43420,N_44230);
and U47362 (N_47362,N_42923,N_42560);
nor U47363 (N_47363,N_43266,N_44226);
or U47364 (N_47364,N_43105,N_42857);
nand U47365 (N_47365,N_44849,N_43126);
nor U47366 (N_47366,N_44821,N_43375);
or U47367 (N_47367,N_44303,N_42927);
or U47368 (N_47368,N_43202,N_44444);
nand U47369 (N_47369,N_43118,N_43570);
nand U47370 (N_47370,N_43713,N_44163);
or U47371 (N_47371,N_43959,N_43282);
nand U47372 (N_47372,N_44076,N_44001);
and U47373 (N_47373,N_43702,N_42822);
xor U47374 (N_47374,N_43843,N_42675);
nor U47375 (N_47375,N_44790,N_43510);
and U47376 (N_47376,N_42781,N_43539);
or U47377 (N_47377,N_43066,N_43065);
nor U47378 (N_47378,N_42601,N_42836);
and U47379 (N_47379,N_42742,N_43906);
or U47380 (N_47380,N_44377,N_44296);
xor U47381 (N_47381,N_43064,N_43118);
nor U47382 (N_47382,N_44284,N_43856);
nor U47383 (N_47383,N_43159,N_43936);
xnor U47384 (N_47384,N_43888,N_43776);
and U47385 (N_47385,N_42905,N_43030);
and U47386 (N_47386,N_44059,N_44093);
or U47387 (N_47387,N_44711,N_42969);
or U47388 (N_47388,N_44702,N_43240);
nand U47389 (N_47389,N_43162,N_43854);
or U47390 (N_47390,N_44485,N_43710);
xnor U47391 (N_47391,N_42525,N_42790);
nor U47392 (N_47392,N_43300,N_44542);
xnor U47393 (N_47393,N_43871,N_43938);
xnor U47394 (N_47394,N_43702,N_44859);
nor U47395 (N_47395,N_44573,N_44946);
nand U47396 (N_47396,N_42883,N_44536);
nor U47397 (N_47397,N_43816,N_43597);
and U47398 (N_47398,N_42939,N_44735);
or U47399 (N_47399,N_44943,N_44157);
and U47400 (N_47400,N_43610,N_44127);
nand U47401 (N_47401,N_43426,N_42924);
and U47402 (N_47402,N_42524,N_44280);
nand U47403 (N_47403,N_44740,N_44585);
xnor U47404 (N_47404,N_43402,N_44449);
and U47405 (N_47405,N_43169,N_44046);
xnor U47406 (N_47406,N_43737,N_43835);
or U47407 (N_47407,N_42796,N_43763);
or U47408 (N_47408,N_44172,N_44083);
nand U47409 (N_47409,N_44910,N_44506);
nor U47410 (N_47410,N_44998,N_44049);
or U47411 (N_47411,N_44104,N_43551);
and U47412 (N_47412,N_44387,N_44705);
xor U47413 (N_47413,N_43123,N_43378);
xor U47414 (N_47414,N_43636,N_43780);
nand U47415 (N_47415,N_44107,N_43365);
xor U47416 (N_47416,N_43844,N_43715);
nand U47417 (N_47417,N_43392,N_44131);
nand U47418 (N_47418,N_44094,N_43755);
xor U47419 (N_47419,N_43698,N_44109);
or U47420 (N_47420,N_42772,N_42712);
nor U47421 (N_47421,N_44024,N_43479);
and U47422 (N_47422,N_43228,N_43745);
and U47423 (N_47423,N_44886,N_43814);
xor U47424 (N_47424,N_44830,N_44977);
nor U47425 (N_47425,N_44669,N_44674);
and U47426 (N_47426,N_44903,N_42770);
xnor U47427 (N_47427,N_44131,N_44767);
xor U47428 (N_47428,N_43321,N_44588);
and U47429 (N_47429,N_44671,N_43529);
and U47430 (N_47430,N_42632,N_44342);
nand U47431 (N_47431,N_43534,N_44700);
or U47432 (N_47432,N_44858,N_42637);
xor U47433 (N_47433,N_42734,N_43175);
xnor U47434 (N_47434,N_43072,N_44609);
xor U47435 (N_47435,N_42930,N_42629);
and U47436 (N_47436,N_43906,N_42608);
nor U47437 (N_47437,N_42991,N_44693);
nor U47438 (N_47438,N_43208,N_44321);
and U47439 (N_47439,N_44126,N_44568);
nor U47440 (N_47440,N_44644,N_44804);
nand U47441 (N_47441,N_43498,N_43974);
and U47442 (N_47442,N_42964,N_43199);
xnor U47443 (N_47443,N_43026,N_44648);
or U47444 (N_47444,N_44083,N_43000);
or U47445 (N_47445,N_44058,N_44998);
or U47446 (N_47446,N_44410,N_44884);
nand U47447 (N_47447,N_43578,N_44334);
nor U47448 (N_47448,N_42588,N_42648);
nor U47449 (N_47449,N_42695,N_44359);
nor U47450 (N_47450,N_43355,N_44316);
xor U47451 (N_47451,N_43850,N_42510);
xnor U47452 (N_47452,N_44394,N_44648);
xor U47453 (N_47453,N_42964,N_43418);
nand U47454 (N_47454,N_42546,N_42908);
nand U47455 (N_47455,N_44293,N_44952);
xnor U47456 (N_47456,N_44167,N_43728);
nor U47457 (N_47457,N_43401,N_43735);
or U47458 (N_47458,N_44782,N_44388);
or U47459 (N_47459,N_42695,N_43648);
and U47460 (N_47460,N_44604,N_44615);
nor U47461 (N_47461,N_43281,N_43613);
nand U47462 (N_47462,N_44766,N_44443);
nand U47463 (N_47463,N_44657,N_43101);
or U47464 (N_47464,N_44159,N_42736);
xor U47465 (N_47465,N_44270,N_42782);
nand U47466 (N_47466,N_42964,N_43092);
xor U47467 (N_47467,N_44995,N_42858);
or U47468 (N_47468,N_42734,N_42983);
or U47469 (N_47469,N_43674,N_43984);
or U47470 (N_47470,N_44372,N_44417);
xnor U47471 (N_47471,N_44826,N_43066);
nand U47472 (N_47472,N_43469,N_44681);
nor U47473 (N_47473,N_43672,N_42815);
nand U47474 (N_47474,N_44440,N_43698);
and U47475 (N_47475,N_44783,N_43558);
nand U47476 (N_47476,N_43086,N_43625);
and U47477 (N_47477,N_43919,N_44763);
or U47478 (N_47478,N_44013,N_44755);
and U47479 (N_47479,N_44486,N_44857);
and U47480 (N_47480,N_43082,N_42785);
nand U47481 (N_47481,N_43664,N_44131);
and U47482 (N_47482,N_44609,N_43925);
nand U47483 (N_47483,N_43345,N_43340);
or U47484 (N_47484,N_43838,N_44659);
nor U47485 (N_47485,N_43067,N_42726);
xnor U47486 (N_47486,N_44177,N_43591);
nand U47487 (N_47487,N_43830,N_44436);
xor U47488 (N_47488,N_43559,N_42507);
nor U47489 (N_47489,N_42504,N_42817);
nand U47490 (N_47490,N_43875,N_44927);
nand U47491 (N_47491,N_43669,N_43659);
and U47492 (N_47492,N_42907,N_43444);
and U47493 (N_47493,N_44247,N_44389);
or U47494 (N_47494,N_43239,N_42826);
or U47495 (N_47495,N_44176,N_42520);
nand U47496 (N_47496,N_42722,N_43827);
and U47497 (N_47497,N_44783,N_44630);
nand U47498 (N_47498,N_42794,N_44585);
nand U47499 (N_47499,N_44537,N_43656);
or U47500 (N_47500,N_47117,N_47008);
nor U47501 (N_47501,N_45684,N_45272);
nor U47502 (N_47502,N_47384,N_45713);
xor U47503 (N_47503,N_45472,N_45154);
nand U47504 (N_47504,N_45956,N_46345);
xnor U47505 (N_47505,N_46058,N_46403);
and U47506 (N_47506,N_46883,N_45501);
nand U47507 (N_47507,N_45046,N_45774);
nor U47508 (N_47508,N_45582,N_46655);
or U47509 (N_47509,N_45425,N_46662);
and U47510 (N_47510,N_46445,N_45077);
xnor U47511 (N_47511,N_45932,N_45992);
xor U47512 (N_47512,N_47287,N_47068);
xor U47513 (N_47513,N_46247,N_46522);
or U47514 (N_47514,N_46553,N_45903);
nand U47515 (N_47515,N_47043,N_46430);
or U47516 (N_47516,N_45380,N_46674);
and U47517 (N_47517,N_46929,N_45883);
and U47518 (N_47518,N_46742,N_46242);
nor U47519 (N_47519,N_45906,N_46221);
xor U47520 (N_47520,N_46277,N_47203);
nand U47521 (N_47521,N_45726,N_47391);
and U47522 (N_47522,N_47317,N_45608);
nand U47523 (N_47523,N_47263,N_46377);
and U47524 (N_47524,N_47086,N_47021);
nor U47525 (N_47525,N_46811,N_45568);
nor U47526 (N_47526,N_46573,N_45764);
nor U47527 (N_47527,N_45329,N_45187);
and U47528 (N_47528,N_46535,N_46840);
xnor U47529 (N_47529,N_45673,N_45005);
nor U47530 (N_47530,N_47237,N_47176);
and U47531 (N_47531,N_47286,N_45523);
and U47532 (N_47532,N_46507,N_46803);
nor U47533 (N_47533,N_45240,N_45863);
and U47534 (N_47534,N_46176,N_46670);
xnor U47535 (N_47535,N_45689,N_46661);
xor U47536 (N_47536,N_45864,N_46266);
nor U47537 (N_47537,N_46005,N_46678);
xor U47538 (N_47538,N_46677,N_47249);
nor U47539 (N_47539,N_46822,N_46002);
nor U47540 (N_47540,N_46463,N_45557);
or U47541 (N_47541,N_47202,N_46303);
and U47542 (N_47542,N_46295,N_46290);
and U47543 (N_47543,N_47389,N_47268);
and U47544 (N_47544,N_45592,N_47280);
nor U47545 (N_47545,N_47294,N_47358);
xor U47546 (N_47546,N_46630,N_45550);
or U47547 (N_47547,N_47360,N_45064);
xnor U47548 (N_47548,N_46825,N_45198);
nor U47549 (N_47549,N_46877,N_46646);
or U47550 (N_47550,N_45423,N_46635);
nand U47551 (N_47551,N_47327,N_45375);
or U47552 (N_47552,N_47083,N_46019);
xnor U47553 (N_47553,N_45468,N_46419);
or U47554 (N_47554,N_46093,N_47055);
and U47555 (N_47555,N_46146,N_47073);
xnor U47556 (N_47556,N_45756,N_47072);
and U47557 (N_47557,N_46517,N_46140);
and U47558 (N_47558,N_45373,N_46565);
nand U47559 (N_47559,N_46502,N_47272);
xor U47560 (N_47560,N_45934,N_46210);
and U47561 (N_47561,N_46501,N_45929);
and U47562 (N_47562,N_45312,N_47416);
nand U47563 (N_47563,N_45014,N_46183);
xnor U47564 (N_47564,N_47433,N_47188);
nor U47565 (N_47565,N_45850,N_46013);
or U47566 (N_47566,N_46957,N_46784);
xnor U47567 (N_47567,N_45354,N_45035);
or U47568 (N_47568,N_47370,N_47463);
xor U47569 (N_47569,N_45034,N_46359);
nor U47570 (N_47570,N_47491,N_47329);
and U47571 (N_47571,N_46091,N_46293);
and U47572 (N_47572,N_45421,N_47366);
xor U47573 (N_47573,N_45660,N_47196);
and U47574 (N_47574,N_46105,N_47483);
nand U47575 (N_47575,N_46379,N_45114);
or U47576 (N_47576,N_45287,N_47446);
and U47577 (N_47577,N_45369,N_45862);
and U47578 (N_47578,N_45715,N_46961);
and U47579 (N_47579,N_46933,N_45922);
nor U47580 (N_47580,N_46753,N_45772);
or U47581 (N_47581,N_47146,N_45631);
and U47582 (N_47582,N_45600,N_45765);
nand U47583 (N_47583,N_47304,N_46941);
nand U47584 (N_47584,N_45967,N_45227);
and U47585 (N_47585,N_45442,N_46046);
nand U47586 (N_47586,N_47404,N_46203);
nor U47587 (N_47587,N_46799,N_46441);
nand U47588 (N_47588,N_45145,N_46763);
xnor U47589 (N_47589,N_46400,N_46619);
and U47590 (N_47590,N_46120,N_46275);
or U47591 (N_47591,N_47379,N_45703);
nor U47592 (N_47592,N_45693,N_47256);
nand U47593 (N_47593,N_45802,N_45984);
and U47594 (N_47594,N_46551,N_47096);
xor U47595 (N_47595,N_45271,N_45230);
nand U47596 (N_47596,N_47039,N_46059);
or U47597 (N_47597,N_47435,N_46174);
or U47598 (N_47598,N_46556,N_45820);
or U47599 (N_47599,N_47130,N_47000);
nand U47600 (N_47600,N_47092,N_47208);
and U47601 (N_47601,N_46425,N_46813);
or U47602 (N_47602,N_46890,N_45178);
and U47603 (N_47603,N_45352,N_45616);
nor U47604 (N_47604,N_46332,N_45307);
xor U47605 (N_47605,N_45951,N_47399);
nor U47606 (N_47606,N_45885,N_45790);
or U47607 (N_47607,N_46734,N_47323);
nor U47608 (N_47608,N_47177,N_46707);
nor U47609 (N_47609,N_45714,N_46084);
and U47610 (N_47610,N_47291,N_46424);
or U47611 (N_47611,N_45700,N_45471);
or U47612 (N_47612,N_46545,N_47163);
xor U47613 (N_47613,N_46166,N_46226);
nor U47614 (N_47614,N_45622,N_46284);
and U47615 (N_47615,N_46778,N_45718);
nor U47616 (N_47616,N_46469,N_46860);
or U47617 (N_47617,N_46557,N_46371);
xor U47618 (N_47618,N_46847,N_45742);
xor U47619 (N_47619,N_45514,N_45666);
xnor U47620 (N_47620,N_46008,N_46513);
nor U47621 (N_47621,N_46857,N_46603);
nor U47622 (N_47622,N_46600,N_47315);
nand U47623 (N_47623,N_47172,N_45844);
or U47624 (N_47624,N_45831,N_46334);
nand U47625 (N_47625,N_45098,N_46375);
and U47626 (N_47626,N_46363,N_46453);
and U47627 (N_47627,N_45437,N_46616);
nor U47628 (N_47628,N_45522,N_46532);
or U47629 (N_47629,N_45678,N_47236);
or U47630 (N_47630,N_45356,N_46063);
and U47631 (N_47631,N_46526,N_45265);
nor U47632 (N_47632,N_46828,N_46190);
nand U47633 (N_47633,N_45630,N_45047);
xnor U47634 (N_47634,N_46625,N_45422);
or U47635 (N_47635,N_46155,N_47178);
nor U47636 (N_47636,N_46383,N_47487);
nor U47637 (N_47637,N_47498,N_46353);
nand U47638 (N_47638,N_46801,N_45427);
nor U47639 (N_47639,N_45815,N_46267);
or U47640 (N_47640,N_45672,N_47201);
xor U47641 (N_47641,N_47023,N_47065);
nor U47642 (N_47642,N_47228,N_45734);
and U47643 (N_47643,N_46394,N_47207);
nand U47644 (N_47644,N_46924,N_45910);
nand U47645 (N_47645,N_47364,N_45394);
or U47646 (N_47646,N_45873,N_45736);
nand U47647 (N_47647,N_46444,N_45701);
or U47648 (N_47648,N_45092,N_46211);
nor U47649 (N_47649,N_47266,N_45403);
xor U47650 (N_47650,N_45599,N_47362);
and U47651 (N_47651,N_45118,N_46858);
or U47652 (N_47652,N_47441,N_47143);
and U47653 (N_47653,N_46082,N_47396);
and U47654 (N_47654,N_46824,N_46989);
or U47655 (N_47655,N_46997,N_46173);
nand U47656 (N_47656,N_45419,N_46200);
nor U47657 (N_47657,N_46918,N_46204);
nor U47658 (N_47658,N_45562,N_46885);
or U47659 (N_47659,N_47038,N_45481);
xor U47660 (N_47660,N_46239,N_45544);
or U47661 (N_47661,N_46596,N_46384);
nand U47662 (N_47662,N_45033,N_45779);
nor U47663 (N_47663,N_46324,N_46805);
and U47664 (N_47664,N_46388,N_46570);
and U47665 (N_47665,N_46669,N_46952);
or U47666 (N_47666,N_45185,N_46869);
or U47667 (N_47667,N_46834,N_47206);
and U47668 (N_47668,N_45829,N_45743);
nor U47669 (N_47669,N_45594,N_46560);
nand U47670 (N_47670,N_45325,N_47278);
nor U47671 (N_47671,N_45813,N_46968);
or U47672 (N_47672,N_45584,N_46697);
xor U47673 (N_47673,N_46389,N_47400);
xor U47674 (N_47674,N_45087,N_45502);
xor U47675 (N_47675,N_46761,N_47497);
or U47676 (N_47676,N_45331,N_45366);
xor U47677 (N_47677,N_46939,N_46902);
or U47678 (N_47678,N_47158,N_46282);
xnor U47679 (N_47679,N_46360,N_47140);
or U47680 (N_47680,N_46464,N_46065);
nand U47681 (N_47681,N_45722,N_45186);
xnor U47682 (N_47682,N_45027,N_45337);
nor U47683 (N_47683,N_46580,N_45099);
nor U47684 (N_47684,N_46546,N_45081);
xor U47685 (N_47685,N_46123,N_46548);
nand U47686 (N_47686,N_47063,N_46497);
xnor U47687 (N_47687,N_46346,N_45454);
and U47688 (N_47688,N_46696,N_46607);
xor U47689 (N_47689,N_45058,N_46523);
xor U47690 (N_47690,N_45542,N_47392);
nand U47691 (N_47691,N_47316,N_46244);
or U47692 (N_47692,N_45179,N_46196);
xnor U47693 (N_47693,N_45727,N_46895);
nor U47694 (N_47694,N_45635,N_47041);
nor U47695 (N_47695,N_47015,N_45121);
nor U47696 (N_47696,N_45129,N_45042);
or U47697 (N_47697,N_47118,N_45900);
nand U47698 (N_47698,N_45441,N_47415);
nor U47699 (N_47699,N_47253,N_46385);
or U47700 (N_47700,N_47462,N_47024);
and U47701 (N_47701,N_46485,N_46426);
and U47702 (N_47702,N_46539,N_46350);
nand U47703 (N_47703,N_46151,N_45881);
or U47704 (N_47704,N_45558,N_45593);
or U47705 (N_47705,N_47056,N_46982);
xor U47706 (N_47706,N_45143,N_46454);
xor U47707 (N_47707,N_46547,N_45504);
or U47708 (N_47708,N_47260,N_45220);
and U47709 (N_47709,N_46837,N_46102);
xnor U47710 (N_47710,N_46578,N_46404);
xor U47711 (N_47711,N_45604,N_45547);
and U47712 (N_47712,N_46709,N_47046);
nor U47713 (N_47713,N_45106,N_45770);
nand U47714 (N_47714,N_46327,N_47185);
nor U47715 (N_47715,N_46977,N_47213);
nand U47716 (N_47716,N_47074,N_45163);
xor U47717 (N_47717,N_45784,N_46722);
nor U47718 (N_47718,N_46964,N_45183);
xor U47719 (N_47719,N_47411,N_46762);
nor U47720 (N_47720,N_47070,N_45962);
and U47721 (N_47721,N_45310,N_47250);
and U47722 (N_47722,N_46496,N_46157);
or U47723 (N_47723,N_47326,N_46618);
xor U47724 (N_47724,N_46468,N_46294);
nand U47725 (N_47725,N_45258,N_46054);
xnor U47726 (N_47726,N_47339,N_45219);
nand U47727 (N_47727,N_46789,N_45102);
nand U47728 (N_47728,N_47368,N_45378);
xor U47729 (N_47729,N_46311,N_46505);
nand U47730 (N_47730,N_45182,N_47406);
nand U47731 (N_47731,N_45549,N_46126);
and U47732 (N_47732,N_46695,N_45509);
nand U47733 (N_47733,N_46279,N_45595);
nand U47734 (N_47734,N_46893,N_47468);
and U47735 (N_47735,N_46634,N_46168);
xor U47736 (N_47736,N_46369,N_45867);
and U47737 (N_47737,N_45978,N_45959);
or U47738 (N_47738,N_46410,N_45827);
nand U47739 (N_47739,N_45977,N_45308);
nand U47740 (N_47740,N_45979,N_45412);
and U47741 (N_47741,N_47331,N_47090);
and U47742 (N_47742,N_47114,N_46721);
or U47743 (N_47743,N_45398,N_45474);
and U47744 (N_47744,N_46593,N_45127);
nand U47745 (N_47745,N_46568,N_46639);
xnor U47746 (N_47746,N_46590,N_45644);
nor U47747 (N_47747,N_46955,N_45376);
and U47748 (N_47748,N_46199,N_46621);
nand U47749 (N_47749,N_47128,N_45073);
or U47750 (N_47750,N_46631,N_45424);
xnor U47751 (N_47751,N_45688,N_45926);
or U47752 (N_47752,N_45180,N_47034);
and U47753 (N_47753,N_46047,N_45548);
nand U47754 (N_47754,N_45225,N_46702);
or U47755 (N_47755,N_45912,N_45079);
xnor U47756 (N_47756,N_47171,N_47160);
nand U47757 (N_47757,N_46671,N_46182);
or U47758 (N_47758,N_46665,N_46132);
nand U47759 (N_47759,N_47014,N_45787);
or U47760 (N_47760,N_46029,N_46448);
and U47761 (N_47761,N_46122,N_46882);
xnor U47762 (N_47762,N_47381,N_45924);
nor U47763 (N_47763,N_46032,N_46238);
nand U47764 (N_47764,N_46352,N_45963);
nor U47765 (N_47765,N_45731,N_45800);
nor U47766 (N_47766,N_46544,N_45998);
and U47767 (N_47767,N_46848,N_46731);
and U47768 (N_47768,N_47452,N_45116);
or U47769 (N_47769,N_47003,N_45482);
or U47770 (N_47770,N_46412,N_45891);
xor U47771 (N_47771,N_47067,N_46959);
and U47772 (N_47772,N_46318,N_46393);
xor U47773 (N_47773,N_46508,N_46880);
xnor U47774 (N_47774,N_46344,N_45960);
xnor U47775 (N_47775,N_46569,N_46990);
xnor U47776 (N_47776,N_47194,N_45836);
xnor U47777 (N_47777,N_45839,N_45477);
nand U47778 (N_47778,N_45262,N_47397);
and U47779 (N_47779,N_45916,N_46835);
nand U47780 (N_47780,N_45538,N_45264);
xnor U47781 (N_47781,N_47245,N_46622);
nand U47782 (N_47782,N_46021,N_47393);
nand U47783 (N_47783,N_46215,N_46730);
xor U47784 (N_47784,N_47351,N_46107);
xnor U47785 (N_47785,N_47112,N_45276);
nor U47786 (N_47786,N_45364,N_45681);
nand U47787 (N_47787,N_47173,N_45101);
nor U47788 (N_47788,N_46489,N_45526);
nand U47789 (N_47789,N_45858,N_45964);
and U47790 (N_47790,N_47062,N_45711);
nand U47791 (N_47791,N_46237,N_46897);
nor U47792 (N_47792,N_46009,N_47174);
nand U47793 (N_47793,N_45685,N_45347);
xnor U47794 (N_47794,N_47141,N_46449);
xor U47795 (N_47795,N_45199,N_46610);
nand U47796 (N_47796,N_45295,N_47283);
or U47797 (N_47797,N_45024,N_45286);
nor U47798 (N_47798,N_45654,N_46398);
or U47799 (N_47799,N_46078,N_45254);
and U47800 (N_47800,N_46358,N_47279);
and U47801 (N_47801,N_46310,N_47119);
or U47802 (N_47802,N_46988,N_45339);
nand U47803 (N_47803,N_46816,N_46777);
nor U47804 (N_47804,N_45702,N_45796);
xor U47805 (N_47805,N_45221,N_45060);
or U47806 (N_47806,N_46846,N_46527);
or U47807 (N_47807,N_45747,N_47352);
xor U47808 (N_47808,N_45828,N_45357);
xor U47809 (N_47809,N_47057,N_46772);
and U47810 (N_47810,N_45346,N_47101);
xnor U47811 (N_47811,N_47239,N_45162);
or U47812 (N_47812,N_46067,N_45231);
xor U47813 (N_47813,N_45336,N_47145);
xnor U47814 (N_47814,N_45508,N_46498);
and U47815 (N_47815,N_46042,N_46160);
and U47816 (N_47816,N_45652,N_46724);
and U47817 (N_47817,N_46628,N_46475);
nor U47818 (N_47818,N_45462,N_46458);
nand U47819 (N_47819,N_47031,N_45946);
and U47820 (N_47820,N_46206,N_45218);
nand U47821 (N_47821,N_46647,N_46845);
and U47822 (N_47822,N_45755,N_45241);
xnor U47823 (N_47823,N_47144,N_45745);
xnor U47824 (N_47824,N_46866,N_46863);
nand U47825 (N_47825,N_46024,N_46104);
xnor U47826 (N_47826,N_45418,N_45123);
xnor U47827 (N_47827,N_46689,N_46372);
or U47828 (N_47828,N_46313,N_46726);
xor U47829 (N_47829,N_47269,N_46335);
nand U47830 (N_47830,N_45050,N_45100);
nor U47831 (N_47831,N_46033,N_45498);
xor U47832 (N_47832,N_46124,N_46749);
nand U47833 (N_47833,N_45506,N_45160);
nor U47834 (N_47834,N_46003,N_47225);
nor U47835 (N_47835,N_45029,N_45249);
xor U47836 (N_47836,N_45395,N_45445);
and U47837 (N_47837,N_45485,N_46719);
and U47838 (N_47838,N_45311,N_46405);
or U47839 (N_47839,N_47258,N_46187);
xnor U47840 (N_47840,N_45659,N_46438);
nand U47841 (N_47841,N_46477,N_46921);
and U47842 (N_47842,N_46336,N_45158);
or U47843 (N_47843,N_46632,N_45011);
nor U47844 (N_47844,N_46240,N_46053);
nor U47845 (N_47845,N_46283,N_45048);
nand U47846 (N_47846,N_46768,N_45222);
xnor U47847 (N_47847,N_46376,N_45546);
nand U47848 (N_47848,N_47181,N_45566);
and U47849 (N_47849,N_45792,N_45453);
nand U47850 (N_47850,N_46451,N_47182);
and U47851 (N_47851,N_45569,N_45294);
and U47852 (N_47852,N_45450,N_46080);
and U47853 (N_47853,N_46515,N_46720);
or U47854 (N_47854,N_46253,N_46069);
nand U47855 (N_47855,N_45012,N_45712);
and U47856 (N_47856,N_46121,N_45629);
xnor U47857 (N_47857,N_47087,N_46299);
and U47858 (N_47858,N_45305,N_45898);
xnor U47859 (N_47859,N_45074,N_47285);
or U47860 (N_47860,N_46759,N_45151);
nand U47861 (N_47861,N_45232,N_46272);
nand U47862 (N_47862,N_46608,N_45812);
nor U47863 (N_47863,N_46494,N_45128);
nand U47864 (N_47864,N_45013,N_45470);
nor U47865 (N_47865,N_45465,N_46434);
or U47866 (N_47866,N_46692,N_45954);
nor U47867 (N_47867,N_47156,N_47490);
nand U47868 (N_47868,N_46914,N_47482);
xor U47869 (N_47869,N_46423,N_46214);
nor U47870 (N_47870,N_45381,N_45390);
nor U47871 (N_47871,N_46432,N_47273);
xor U47872 (N_47872,N_46531,N_47098);
xor U47873 (N_47873,N_46452,N_47438);
nor U47874 (N_47874,N_46965,N_45645);
xor U47875 (N_47875,N_47407,N_47247);
nor U47876 (N_47876,N_45057,N_45658);
and U47877 (N_47877,N_45780,N_46606);
and U47878 (N_47878,N_45233,N_45068);
nand U47879 (N_47879,N_47170,N_47126);
or U47880 (N_47880,N_45191,N_46575);
and U47881 (N_47881,N_46459,N_45917);
nand U47882 (N_47882,N_46504,N_47169);
or U47883 (N_47883,N_45479,N_45444);
nand U47884 (N_47884,N_45018,N_45234);
or U47885 (N_47885,N_45638,N_45819);
or U47886 (N_47886,N_45729,N_46976);
nand U47887 (N_47887,N_45529,N_46681);
xnor U47888 (N_47888,N_46092,N_47495);
nand U47889 (N_47889,N_45786,N_46658);
nor U47890 (N_47890,N_45849,N_46338);
nor U47891 (N_47891,N_46874,N_47025);
or U47892 (N_47892,N_46506,N_45991);
and U47893 (N_47893,N_45860,N_46300);
nand U47894 (N_47894,N_45663,N_46700);
or U47895 (N_47895,N_45344,N_47318);
and U47896 (N_47896,N_47354,N_45144);
nand U47897 (N_47897,N_45795,N_46455);
nor U47898 (N_47898,N_47428,N_47451);
and U47899 (N_47899,N_46907,N_46373);
nand U47900 (N_47900,N_47499,N_46259);
xnor U47901 (N_47901,N_46577,N_46141);
and U47902 (N_47902,N_45406,N_47261);
or U47903 (N_47903,N_46650,N_47002);
and U47904 (N_47904,N_46083,N_45537);
or U47905 (N_47905,N_46483,N_47134);
nor U47906 (N_47906,N_46265,N_46035);
and U47907 (N_47907,N_46037,N_47198);
xor U47908 (N_47908,N_47100,N_45291);
nand U47909 (N_47909,N_45896,N_45319);
xnor U47910 (N_47910,N_47405,N_46747);
and U47911 (N_47911,N_46966,N_45880);
or U47912 (N_47912,N_47032,N_45065);
nand U47913 (N_47913,N_46257,N_46461);
nor U47914 (N_47914,N_45908,N_45530);
nand U47915 (N_47915,N_46552,N_46908);
and U47916 (N_47916,N_45621,N_46367);
and U47917 (N_47917,N_45999,N_47289);
or U47918 (N_47918,N_46030,N_45698);
nand U47919 (N_47919,N_46937,N_46911);
nand U47920 (N_47920,N_45022,N_45096);
or U47921 (N_47921,N_47284,N_46307);
nor U47922 (N_47922,N_45188,N_45516);
nor U47923 (N_47923,N_46827,N_46163);
nand U47924 (N_47924,N_46422,N_45067);
and U47925 (N_47925,N_47390,N_46343);
or U47926 (N_47926,N_45259,N_45174);
nor U47927 (N_47927,N_47122,N_46274);
nand U47928 (N_47928,N_46162,N_45794);
nor U47929 (N_47929,N_45746,N_45799);
and U47930 (N_47930,N_45705,N_46525);
nand U47931 (N_47931,N_45823,N_45499);
xnor U47932 (N_47932,N_46135,N_47312);
xor U47933 (N_47933,N_45785,N_45197);
xnor U47934 (N_47934,N_45733,N_45822);
or U47935 (N_47935,N_45695,N_45435);
xor U47936 (N_47936,N_46171,N_45115);
nand U47937 (N_47937,N_46727,N_45614);
nor U47938 (N_47938,N_47212,N_46550);
or U47939 (N_47939,N_47233,N_46980);
xor U47940 (N_47940,N_47219,N_47257);
nor U47941 (N_47941,N_47108,N_45195);
xor U47942 (N_47942,N_47109,N_45610);
and U47943 (N_47943,N_46390,N_46804);
or U47944 (N_47944,N_45069,N_45580);
xnor U47945 (N_47945,N_45930,N_45436);
or U47946 (N_47946,N_47183,N_45432);
nand U47947 (N_47947,N_46676,N_47467);
nand U47948 (N_47948,N_46129,N_46051);
nand U47949 (N_47949,N_46011,N_45677);
or U47950 (N_47950,N_45707,N_45203);
or U47951 (N_47951,N_47054,N_45494);
or U47952 (N_47952,N_46076,N_45476);
nor U47953 (N_47953,N_46001,N_45181);
nand U47954 (N_47954,N_45975,N_46062);
or U47955 (N_47955,N_46615,N_45285);
nand U47956 (N_47956,N_45478,N_45244);
xnor U47957 (N_47957,N_47457,N_45124);
nor U47958 (N_47958,N_45400,N_47037);
xnor U47959 (N_47959,N_45920,N_47262);
nor U47960 (N_47960,N_46280,N_47449);
or U47961 (N_47961,N_46045,N_46748);
or U47962 (N_47962,N_46641,N_45788);
xor U47963 (N_47963,N_45345,N_45870);
and U47964 (N_47964,N_45914,N_46213);
nand U47965 (N_47965,N_46698,N_47220);
and U47966 (N_47966,N_47200,N_45791);
xor U47967 (N_47967,N_45063,N_46664);
xor U47968 (N_47968,N_46179,N_46476);
nor U47969 (N_47969,N_45606,N_45613);
or U47970 (N_47970,N_46109,N_45090);
or U47971 (N_47971,N_46212,N_46708);
xor U47972 (N_47972,N_45730,N_46086);
xor U47973 (N_47973,N_46052,N_47157);
or U47974 (N_47974,N_45157,N_47322);
xor U47975 (N_47975,N_46809,N_45653);
nand U47976 (N_47976,N_46429,N_46288);
and U47977 (N_47977,N_47079,N_47064);
xnor U47978 (N_47978,N_45576,N_45149);
or U47979 (N_47979,N_45851,N_45687);
xor U47980 (N_47980,N_45327,N_47081);
or U47981 (N_47981,N_45136,N_46399);
nor U47982 (N_47982,N_47189,N_46150);
xor U47983 (N_47983,N_45300,N_47051);
or U47984 (N_47984,N_45553,N_46466);
xnor U47985 (N_47985,N_46016,N_47373);
and U47986 (N_47986,N_47026,N_46255);
xnor U47987 (N_47987,N_45389,N_46660);
and U47988 (N_47988,N_46865,N_47309);
or U47989 (N_47989,N_45958,N_46723);
xor U47990 (N_47990,N_45611,N_46998);
xor U47991 (N_47991,N_46286,N_46436);
nor U47992 (N_47992,N_45298,N_46447);
xnor U47993 (N_47993,N_46574,N_47431);
nand U47994 (N_47994,N_45490,N_45189);
and U47995 (N_47995,N_45237,N_46795);
xnor U47996 (N_47996,N_46320,N_45031);
or U47997 (N_47997,N_45560,N_45263);
or U47998 (N_47998,N_45290,N_46232);
nand U47999 (N_47999,N_47334,N_45861);
or U48000 (N_48000,N_45109,N_46354);
nand U48001 (N_48001,N_47150,N_46808);
nand U48002 (N_48002,N_45257,N_45717);
xnor U48003 (N_48003,N_45797,N_45933);
or U48004 (N_48004,N_45135,N_47420);
nand U48005 (N_48005,N_46881,N_45517);
xor U48006 (N_48006,N_47179,N_45633);
and U48007 (N_48007,N_46172,N_47013);
or U48008 (N_48008,N_46154,N_45596);
and U48009 (N_48009,N_45173,N_47363);
and U48010 (N_48010,N_46339,N_46983);
or U48011 (N_48011,N_45168,N_46831);
nor U48012 (N_48012,N_47004,N_47053);
nand U48013 (N_48013,N_46579,N_46637);
or U48014 (N_48014,N_47218,N_46319);
xnor U48015 (N_48015,N_45768,N_46186);
nor U48016 (N_48016,N_45075,N_45988);
nand U48017 (N_48017,N_46563,N_46856);
xnor U48018 (N_48018,N_45732,N_45279);
nor U48019 (N_48019,N_46217,N_46685);
nor U48020 (N_48020,N_46156,N_45094);
nand U48021 (N_48021,N_47349,N_45889);
and U48022 (N_48022,N_45210,N_45335);
xor U48023 (N_48023,N_46889,N_46958);
xnor U48024 (N_48024,N_45605,N_45405);
nand U48025 (N_48025,N_46962,N_45670);
and U48026 (N_48026,N_45000,N_47277);
nor U48027 (N_48027,N_45994,N_47342);
or U48028 (N_48028,N_45640,N_46690);
nor U48029 (N_48029,N_45296,N_46943);
nand U48030 (N_48030,N_45169,N_46224);
nand U48031 (N_48031,N_45634,N_45682);
xor U48032 (N_48032,N_47235,N_46873);
xnor U48033 (N_48033,N_46850,N_46216);
xnor U48034 (N_48034,N_47226,N_46910);
or U48035 (N_48035,N_45200,N_45434);
or U48036 (N_48036,N_47251,N_46055);
nand U48037 (N_48037,N_46934,N_46207);
nand U48038 (N_48038,N_46798,N_46871);
nand U48039 (N_48039,N_46725,N_46967);
xnor U48040 (N_48040,N_45059,N_45773);
xnor U48041 (N_48041,N_46602,N_45052);
nand U48042 (N_48042,N_45250,N_45414);
xor U48043 (N_48043,N_47238,N_45440);
xor U48044 (N_48044,N_45039,N_47296);
nor U48045 (N_48045,N_45273,N_47494);
and U48046 (N_48046,N_45541,N_47022);
nand U48047 (N_48047,N_45275,N_46758);
or U48048 (N_48048,N_46756,N_46566);
and U48049 (N_48049,N_45710,N_46442);
xor U48050 (N_48050,N_45103,N_46136);
or U48051 (N_48051,N_45825,N_45533);
xnor U48052 (N_48052,N_45781,N_47136);
xnor U48053 (N_48053,N_47310,N_47427);
or U48054 (N_48054,N_45416,N_46581);
or U48055 (N_48055,N_45856,N_46235);
nor U48056 (N_48056,N_45766,N_46843);
xnor U48057 (N_48057,N_45769,N_46119);
or U48058 (N_48058,N_45620,N_46325);
nand U48059 (N_48059,N_45561,N_45426);
nor U48060 (N_48060,N_45201,N_46942);
xor U48061 (N_48061,N_45567,N_45886);
and U48062 (N_48062,N_46012,N_46872);
and U48063 (N_48063,N_47151,N_47217);
nand U48064 (N_48064,N_45853,N_45651);
or U48065 (N_48065,N_46841,N_45388);
xor U48066 (N_48066,N_45457,N_46760);
or U48067 (N_48067,N_45334,N_46740);
xor U48068 (N_48068,N_46036,N_46096);
or U48069 (N_48069,N_45464,N_45838);
and U48070 (N_48070,N_46595,N_47107);
nor U48071 (N_48071,N_45093,N_46153);
nor U48072 (N_48072,N_45407,N_47049);
nor U48073 (N_48073,N_45527,N_45261);
nor U48074 (N_48074,N_45997,N_46859);
nand U48075 (N_48075,N_46912,N_46819);
nor U48076 (N_48076,N_45391,N_47275);
nor U48077 (N_48077,N_45783,N_45655);
or U48078 (N_48078,N_46133,N_45585);
nand U48079 (N_48079,N_45628,N_45540);
xnor U48080 (N_48080,N_47408,N_47432);
or U48081 (N_48081,N_47071,N_45669);
xor U48082 (N_48082,N_45256,N_45313);
nand U48083 (N_48083,N_45818,N_46302);
nand U48084 (N_48084,N_46064,N_47165);
or U48085 (N_48085,N_45359,N_45503);
xor U48086 (N_48086,N_45070,N_46340);
nand U48087 (N_48087,N_45306,N_45952);
and U48088 (N_48088,N_45942,N_45206);
or U48089 (N_48089,N_47149,N_47295);
or U48090 (N_48090,N_46472,N_46588);
nor U48091 (N_48091,N_45913,N_47116);
nor U48092 (N_48092,N_47093,N_47270);
xor U48093 (N_48093,N_45948,N_47292);
or U48094 (N_48094,N_46220,N_46457);
and U48095 (N_48095,N_47010,N_45449);
or U48096 (N_48096,N_46659,N_46167);
or U48097 (N_48097,N_47489,N_46528);
or U48098 (N_48098,N_46776,N_45888);
or U48099 (N_48099,N_46613,N_45646);
nor U48100 (N_48100,N_47191,N_47424);
and U48101 (N_48101,N_45512,N_47454);
xor U48102 (N_48102,N_46309,N_45155);
nand U48103 (N_48103,N_45455,N_46397);
nor U48104 (N_48104,N_46169,N_46147);
and U48105 (N_48105,N_46473,N_45415);
xnor U48106 (N_48106,N_46180,N_47448);
or U48107 (N_48107,N_45662,N_46439);
nand U48108 (N_48108,N_46718,N_46007);
and U48109 (N_48109,N_45045,N_47125);
nor U48110 (N_48110,N_46330,N_46783);
xor U48111 (N_48111,N_46479,N_45759);
nand U48112 (N_48112,N_45413,N_46741);
xnor U48113 (N_48113,N_46478,N_47298);
or U48114 (N_48114,N_46940,N_45845);
or U48115 (N_48115,N_45235,N_46868);
xnor U48116 (N_48116,N_46049,N_47180);
and U48117 (N_48117,N_46349,N_46999);
xnor U48118 (N_48118,N_47209,N_47231);
or U48119 (N_48119,N_46711,N_46842);
xnor U48120 (N_48120,N_45491,N_46886);
or U48121 (N_48121,N_46056,N_46737);
or U48122 (N_48122,N_45026,N_46095);
and U48123 (N_48123,N_47274,N_46420);
xor U48124 (N_48124,N_46950,N_45615);
xor U48125 (N_48125,N_46855,N_45082);
nor U48126 (N_48126,N_46717,N_46605);
or U48127 (N_48127,N_45358,N_46733);
nor U48128 (N_48128,N_47414,N_45379);
or U48129 (N_48129,N_47168,N_45559);
or U48130 (N_48130,N_46268,N_47131);
xnor U48131 (N_48131,N_47372,N_47036);
xnor U48132 (N_48132,N_47264,N_45053);
nand U48133 (N_48133,N_45322,N_47330);
or U48134 (N_48134,N_45475,N_45573);
xnor U48135 (N_48135,N_46567,N_45480);
xor U48136 (N_48136,N_46254,N_45431);
and U48137 (N_48137,N_46488,N_45872);
or U48138 (N_48138,N_46810,N_47005);
and U48139 (N_48139,N_46814,N_46088);
or U48140 (N_48140,N_46218,N_46571);
or U48141 (N_48141,N_47470,N_45142);
or U48142 (N_48142,N_45260,N_46139);
xor U48143 (N_48143,N_45321,N_45950);
or U48144 (N_48144,N_45384,N_46764);
or U48145 (N_48145,N_46559,N_45696);
or U48146 (N_48146,N_46108,N_46766);
nand U48147 (N_48147,N_46418,N_45854);
nor U48148 (N_48148,N_47387,N_45055);
xnor U48149 (N_48149,N_46862,N_46657);
nor U48150 (N_48150,N_45269,N_46978);
nor U48151 (N_48151,N_46048,N_47303);
or U48152 (N_48152,N_45811,N_45957);
nand U48153 (N_48153,N_47450,N_47078);
nand U48154 (N_48154,N_46903,N_46612);
nand U48155 (N_48155,N_46694,N_46735);
and U48156 (N_48156,N_46785,N_47197);
xor U48157 (N_48157,N_47375,N_45456);
and U48158 (N_48158,N_46791,N_46357);
nor U48159 (N_48159,N_45966,N_46867);
and U48160 (N_48160,N_47475,N_45761);
or U48161 (N_48161,N_45519,N_45170);
nand U48162 (N_48162,N_46624,N_45299);
nand U48163 (N_48163,N_45385,N_45875);
nand U48164 (N_48164,N_45625,N_47382);
nor U48165 (N_48165,N_45382,N_47338);
nand U48166 (N_48166,N_45571,N_46192);
or U48167 (N_48167,N_45981,N_45895);
or U48168 (N_48168,N_45641,N_46401);
and U48169 (N_48169,N_45720,N_45152);
nor U48170 (N_48170,N_45342,N_45507);
nor U48171 (N_48171,N_46757,N_45983);
or U48172 (N_48172,N_46538,N_45840);
nand U48173 (N_48173,N_46020,N_46838);
nand U48174 (N_48174,N_47230,N_45023);
or U48175 (N_48175,N_46038,N_45493);
and U48176 (N_48176,N_45111,N_46271);
xnor U48177 (N_48177,N_45226,N_47102);
xor U48178 (N_48178,N_45061,N_45944);
and U48179 (N_48179,N_46263,N_46361);
xor U48180 (N_48180,N_47030,N_45572);
nand U48181 (N_48181,N_46993,N_46482);
nor U48182 (N_48182,N_46913,N_46787);
and U48183 (N_48183,N_45289,N_46643);
xor U48184 (N_48184,N_45555,N_46301);
and U48185 (N_48185,N_46072,N_45985);
xor U48186 (N_48186,N_46896,N_46415);
xnor U48187 (N_48187,N_46039,N_46672);
and U48188 (N_48188,N_45428,N_45371);
nand U48189 (N_48189,N_46380,N_45377);
or U48190 (N_48190,N_46308,N_45824);
or U48191 (N_48191,N_46656,N_45939);
nor U48192 (N_48192,N_45458,N_46099);
and U48193 (N_48193,N_46414,N_45921);
nand U48194 (N_48194,N_46223,N_46744);
xor U48195 (N_48195,N_45500,N_46686);
nor U48196 (N_48196,N_46701,N_46100);
or U48197 (N_48197,N_47458,N_47359);
or U48198 (N_48198,N_47033,N_45270);
nand U48199 (N_48199,N_46587,N_47455);
xnor U48200 (N_48200,N_47159,N_46499);
xnor U48201 (N_48201,N_45724,N_47418);
nor U48202 (N_48202,N_47313,N_46576);
or U48203 (N_48203,N_47383,N_46894);
nor U48204 (N_48204,N_45484,N_46351);
xnor U48205 (N_48205,N_46802,N_45947);
or U48206 (N_48206,N_45617,N_46411);
nor U48207 (N_48207,N_46134,N_45165);
or U48208 (N_48208,N_46815,N_46081);
xor U48209 (N_48209,N_45545,N_47175);
nand U48210 (N_48210,N_47474,N_45597);
xnor U48211 (N_48211,N_45816,N_46374);
or U48212 (N_48212,N_47471,N_45280);
nand U48213 (N_48213,N_46985,N_47476);
xor U48214 (N_48214,N_46935,N_45528);
and U48215 (N_48215,N_45126,N_46000);
nand U48216 (N_48216,N_46514,N_45213);
xor U48217 (N_48217,N_46427,N_47110);
or U48218 (N_48218,N_45973,N_45190);
and U48219 (N_48219,N_45447,N_45513);
xor U48220 (N_48220,N_45446,N_46561);
and U48221 (N_48221,N_45601,N_47341);
nor U48222 (N_48222,N_46406,N_47137);
nand U48223 (N_48223,N_47337,N_46408);
nand U48224 (N_48224,N_47473,N_46061);
and U48225 (N_48225,N_46094,N_47293);
nor U48226 (N_48226,N_45833,N_45066);
nor U48227 (N_48227,N_45931,N_45753);
nand U48228 (N_48228,N_46460,N_45043);
and U48229 (N_48229,N_45323,N_46584);
or U48230 (N_48230,N_46923,N_46636);
nor U48231 (N_48231,N_45612,N_47161);
and U48232 (N_48232,N_45808,N_46111);
nor U48233 (N_48233,N_45438,N_46833);
xor U48234 (N_48234,N_46337,N_45876);
nor U48235 (N_48235,N_45019,N_46250);
or U48236 (N_48236,N_45164,N_46421);
and U48237 (N_48237,N_46209,N_45793);
xnor U48238 (N_48238,N_46945,N_45976);
nand U48239 (N_48239,N_46329,N_45309);
nand U48240 (N_48240,N_47216,N_46381);
nand U48241 (N_48241,N_46645,N_45524);
and U48242 (N_48242,N_47082,N_46969);
xnor U48243 (N_48243,N_46555,N_47395);
and U48244 (N_48244,N_46050,N_45211);
nor U48245 (N_48245,N_45040,N_45789);
or U48246 (N_48246,N_45238,N_46644);
xor U48247 (N_48247,N_46909,N_47139);
nor U48248 (N_48248,N_45004,N_45392);
and U48249 (N_48249,N_45316,N_46688);
xnor U48250 (N_48250,N_47164,N_45704);
or U48251 (N_48251,N_47422,N_45281);
and U48252 (N_48252,N_46066,N_45028);
nand U48253 (N_48253,N_45021,N_45147);
nand U48254 (N_48254,N_46653,N_45452);
nand U48255 (N_48255,N_46620,N_46994);
nor U48256 (N_48256,N_45832,N_45497);
or U48257 (N_48257,N_47479,N_47403);
xor U48258 (N_48258,N_45564,N_46006);
or U48259 (N_48259,N_47227,N_46278);
or U48260 (N_48260,N_46807,N_45171);
nand U48261 (N_48261,N_45980,N_46145);
nor U48262 (N_48262,N_46640,N_46142);
nor U48263 (N_48263,N_45317,N_45953);
and U48264 (N_48264,N_45552,N_46915);
xor U48265 (N_48265,N_47167,N_46710);
nand U48266 (N_48266,N_45138,N_45340);
nor U48267 (N_48267,N_45460,N_46431);
and U48268 (N_48268,N_46870,N_45806);
and U48269 (N_48269,N_45044,N_45565);
nor U48270 (N_48270,N_46564,N_46116);
xor U48271 (N_48271,N_45139,N_45284);
and U48272 (N_48272,N_46490,N_47409);
or U48273 (N_48273,N_45148,N_47244);
nand U48274 (N_48274,N_45543,N_45056);
xnor U48275 (N_48275,N_45393,N_45837);
or U48276 (N_48276,N_45563,N_45303);
nand U48277 (N_48277,N_45383,N_45972);
or U48278 (N_48278,N_45374,N_47028);
nand U48279 (N_48279,N_46471,N_46916);
and U48280 (N_48280,N_46500,N_46594);
and U48281 (N_48281,N_46888,N_45740);
and U48282 (N_48282,N_46495,N_46480);
xnor U48283 (N_48283,N_46861,N_45803);
or U48284 (N_48284,N_46298,N_47016);
nand U48285 (N_48285,N_46853,N_47232);
or U48286 (N_48286,N_45750,N_46792);
nand U48287 (N_48287,N_47027,N_45360);
xor U48288 (N_48288,N_46963,N_46754);
or U48289 (N_48289,N_46786,N_46227);
xnor U48290 (N_48290,N_45387,N_46973);
nand U48291 (N_48291,N_47300,N_47430);
and U48292 (N_48292,N_45901,N_45842);
or U48293 (N_48293,N_47429,N_46386);
nor U48294 (N_48294,N_45738,N_45278);
nor U48295 (N_48295,N_46149,N_45459);
nor U48296 (N_48296,N_46932,N_45466);
or U48297 (N_48297,N_46492,N_46470);
xnor U48298 (N_48298,N_45324,N_45899);
nand U48299 (N_48299,N_46366,N_47211);
or U48300 (N_48300,N_45015,N_45535);
and U48301 (N_48301,N_46437,N_46562);
nor U48302 (N_48302,N_45859,N_47190);
or U48303 (N_48303,N_47259,N_45776);
nand U48304 (N_48304,N_45866,N_47138);
xor U48305 (N_48305,N_47029,N_47091);
and U48306 (N_48306,N_45603,N_45302);
xor U48307 (N_48307,N_46728,N_47006);
xnor U48308 (N_48308,N_46623,N_46365);
and U48309 (N_48309,N_46751,N_47120);
nor U48310 (N_48310,N_46987,N_45062);
or U48311 (N_48311,N_45843,N_46031);
xor U48312 (N_48312,N_46705,N_45804);
xor U48313 (N_48313,N_47059,N_45120);
or U48314 (N_48314,N_47486,N_45006);
and U48315 (N_48315,N_47336,N_47045);
xnor U48316 (N_48316,N_45511,N_45996);
nor U48317 (N_48317,N_46316,N_45971);
nor U48318 (N_48318,N_46402,N_46592);
xnor U48319 (N_48319,N_45292,N_46057);
or U48320 (N_48320,N_45032,N_46112);
or U48321 (N_48321,N_46075,N_46509);
or U48322 (N_48322,N_45404,N_46905);
xnor U48323 (N_48323,N_46287,N_46407);
nand U48324 (N_48324,N_45708,N_46771);
xnor U48325 (N_48325,N_45937,N_46781);
or U48326 (N_48326,N_45821,N_46864);
nand U48327 (N_48327,N_45146,N_47413);
nand U48328 (N_48328,N_46970,N_47011);
nor U48329 (N_48329,N_45293,N_45556);
nand U48330 (N_48330,N_46714,N_45451);
and U48331 (N_48331,N_46633,N_45159);
nand U48332 (N_48332,N_47439,N_45207);
or U48333 (N_48333,N_45209,N_45401);
and U48334 (N_48334,N_47319,N_47111);
nor U48335 (N_48335,N_46830,N_45771);
xnor U48336 (N_48336,N_45362,N_45817);
xnor U48337 (N_48337,N_45248,N_45531);
nand U48338 (N_48338,N_45877,N_46900);
nor U48339 (N_48339,N_45609,N_46291);
xor U48340 (N_48340,N_45882,N_45525);
and U48341 (N_48341,N_45461,N_45719);
nor U48342 (N_48342,N_45408,N_46953);
nor U48343 (N_48343,N_45699,N_45846);
and U48344 (N_48344,N_47299,N_46598);
nor U48345 (N_48345,N_47453,N_45007);
nor U48346 (N_48346,N_47348,N_47282);
xnor U48347 (N_48347,N_47355,N_46023);
and U48348 (N_48348,N_46197,N_45038);
or U48349 (N_48349,N_47353,N_47365);
nand U48350 (N_48350,N_45598,N_45246);
nor U48351 (N_48351,N_45869,N_46981);
or U48352 (N_48352,N_45051,N_45215);
and U48353 (N_48353,N_45349,N_47367);
nor U48354 (N_48354,N_47155,N_45949);
and U48355 (N_48355,N_47255,N_46716);
and U48356 (N_48356,N_45489,N_45574);
or U48357 (N_48357,N_45282,N_45367);
nor U48358 (N_48358,N_46322,N_46312);
nor U48359 (N_48359,N_47459,N_46851);
nand U48360 (N_48360,N_47301,N_45857);
nand U48361 (N_48361,N_45807,N_45253);
nor U48362 (N_48362,N_47436,N_46926);
nand U48363 (N_48363,N_45911,N_47388);
xor U48364 (N_48364,N_45488,N_45686);
xnor U48365 (N_48365,N_45623,N_46409);
xor U48366 (N_48366,N_45874,N_47095);
nor U48367 (N_48367,N_46387,N_47445);
xnor U48368 (N_48368,N_47248,N_45835);
and U48369 (N_48369,N_45175,N_46130);
nor U48370 (N_48370,N_46854,N_45330);
nor U48371 (N_48371,N_47224,N_45855);
or U48372 (N_48372,N_45417,N_45752);
xor U48373 (N_48373,N_46917,N_47344);
nand U48374 (N_48374,N_47254,N_46178);
or U48375 (N_48375,N_46165,N_47135);
and U48376 (N_48376,N_46691,N_45961);
or U48377 (N_48377,N_45266,N_46184);
or U48378 (N_48378,N_45036,N_46629);
and U48379 (N_48379,N_45041,N_47058);
nand U48380 (N_48380,N_45632,N_46025);
xnor U48381 (N_48381,N_46416,N_47478);
or U48382 (N_48382,N_46654,N_45909);
xor U48383 (N_48383,N_46392,N_45723);
and U48384 (N_48384,N_45637,N_45767);
xnor U48385 (N_48385,N_45167,N_47195);
xor U48386 (N_48386,N_45304,N_46068);
or U48387 (N_48387,N_46101,N_47271);
xnor U48388 (N_48388,N_46326,N_46530);
nor U48389 (N_48389,N_45941,N_46693);
nor U48390 (N_48390,N_45945,N_46131);
xor U48391 (N_48391,N_46520,N_46829);
or U48392 (N_48392,N_45642,N_47018);
xnor U48393 (N_48393,N_45680,N_46638);
or U48394 (N_48394,N_46668,N_45879);
nor U48395 (N_48395,N_47044,N_47324);
nor U48396 (N_48396,N_46110,N_45496);
nor U48397 (N_48397,N_46585,N_46261);
nand U48398 (N_48398,N_47350,N_46090);
nor U48399 (N_48399,N_46826,N_45429);
xnor U48400 (N_48400,N_47113,N_45777);
or U48401 (N_48401,N_46536,N_46044);
or U48402 (N_48402,N_45010,N_47123);
or U48403 (N_48403,N_45928,N_45368);
and U48404 (N_48404,N_45341,N_47210);
nand U48405 (N_48405,N_46314,N_45868);
and U48406 (N_48406,N_45268,N_45749);
xor U48407 (N_48407,N_45865,N_46770);
nand U48408 (N_48408,N_47356,N_45691);
nor U48409 (N_48409,N_47302,N_46642);
or U48410 (N_48410,N_45037,N_46106);
nand U48411 (N_48411,N_46591,N_46651);
or U48412 (N_48412,N_45217,N_45196);
nor U48413 (N_48413,N_47246,N_46323);
nor U48414 (N_48414,N_46347,N_47496);
and U48415 (N_48415,N_45648,N_47240);
and U48416 (N_48416,N_46158,N_47378);
and U48417 (N_48417,N_45986,N_46193);
xor U48418 (N_48418,N_45647,N_46930);
or U48419 (N_48419,N_46821,N_47243);
xor U48420 (N_48420,N_45890,N_46230);
and U48421 (N_48421,N_46971,N_46878);
or U48422 (N_48422,N_45649,N_46986);
nor U48423 (N_48423,N_45386,N_45871);
nand U48424 (N_48424,N_45229,N_46481);
xnor U48425 (N_48425,N_46996,N_45624);
xor U48426 (N_48426,N_46609,N_47077);
or U48427 (N_48427,N_45676,N_45243);
nand U48428 (N_48428,N_46229,N_45923);
nand U48429 (N_48429,N_46904,N_45469);
or U48430 (N_48430,N_45758,N_47333);
xor U48431 (N_48431,N_45315,N_46769);
nor U48432 (N_48432,N_45274,N_46954);
or U48433 (N_48433,N_45333,N_47106);
nand U48434 (N_48434,N_46519,N_47019);
or U48435 (N_48435,N_46028,N_45725);
or U48436 (N_48436,N_46264,N_46849);
or U48437 (N_48437,N_47345,N_46098);
and U48438 (N_48438,N_45760,N_46248);
and U48439 (N_48439,N_47076,N_45088);
or U48440 (N_48440,N_45439,N_46260);
nand U48441 (N_48441,N_45078,N_45744);
nor U48442 (N_48442,N_47346,N_46228);
or U48443 (N_48443,N_47127,N_46925);
nor U48444 (N_48444,N_45675,N_46297);
and U48445 (N_48445,N_46680,N_47017);
nor U48446 (N_48446,N_45314,N_47488);
and U48447 (N_48447,N_46712,N_45072);
or U48448 (N_48448,N_46512,N_46125);
or U48449 (N_48449,N_46128,N_46800);
xnor U48450 (N_48450,N_45283,N_47204);
nand U48451 (N_48451,N_47321,N_47314);
nor U48452 (N_48452,N_46767,N_47040);
nor U48453 (N_48453,N_47465,N_46014);
xnor U48454 (N_48454,N_46944,N_47147);
xnor U48455 (N_48455,N_46289,N_46746);
nand U48456 (N_48456,N_45318,N_45486);
and U48457 (N_48457,N_46456,N_45927);
xnor U48458 (N_48458,N_45001,N_45355);
and U48459 (N_48459,N_45326,N_45894);
nand U48460 (N_48460,N_47007,N_46285);
nor U48461 (N_48461,N_45878,N_47481);
nand U48462 (N_48462,N_47440,N_47148);
nand U48463 (N_48463,N_46413,N_46995);
and U48464 (N_48464,N_47265,N_45430);
nor U48465 (N_48465,N_46817,N_45242);
or U48466 (N_48466,N_45521,N_45122);
nand U48467 (N_48467,N_45754,N_45097);
nand U48468 (N_48468,N_45551,N_45348);
nor U48469 (N_48469,N_45887,N_45955);
or U48470 (N_48470,N_46077,N_45626);
nor U48471 (N_48471,N_46185,N_46428);
nand U48472 (N_48472,N_46273,N_45365);
xor U48473 (N_48473,N_46920,N_47306);
xnor U48474 (N_48474,N_47048,N_47186);
or U48475 (N_48475,N_47187,N_47242);
nand U48476 (N_48476,N_46276,N_46626);
nand U48477 (N_48477,N_46901,N_45782);
nand U48478 (N_48478,N_47080,N_45581);
nand U48479 (N_48479,N_45016,N_47401);
and U48480 (N_48480,N_45826,N_46765);
and U48481 (N_48481,N_45267,N_46586);
xor U48482 (N_48482,N_45003,N_45935);
or U48483 (N_48483,N_45671,N_47485);
nand U48484 (N_48484,N_46382,N_47229);
nor U48485 (N_48485,N_45156,N_45030);
nand U48486 (N_48486,N_45995,N_46572);
nor U48487 (N_48487,N_45338,N_45668);
nand U48488 (N_48488,N_45539,N_46433);
nand U48489 (N_48489,N_46736,N_45590);
or U48490 (N_48490,N_47426,N_46305);
nor U48491 (N_48491,N_46516,N_46219);
nor U48492 (N_48492,N_46378,N_47276);
xor U48493 (N_48493,N_47009,N_45247);
or U48494 (N_48494,N_45208,N_47357);
and U48495 (N_48495,N_45575,N_46181);
or U48496 (N_48496,N_45236,N_47447);
or U48497 (N_48497,N_46673,N_45578);
nand U48498 (N_48498,N_46823,N_46315);
or U48499 (N_48499,N_45762,N_47380);
nand U48500 (N_48500,N_45589,N_45463);
xnor U48501 (N_48501,N_47084,N_46225);
xnor U48502 (N_48502,N_47132,N_45361);
xnor U48503 (N_48503,N_46589,N_46956);
or U48504 (N_48504,N_46715,N_46627);
nand U48505 (N_48505,N_47184,N_45505);
nand U48506 (N_48506,N_46884,N_46152);
and U48507 (N_48507,N_45137,N_45925);
and U48508 (N_48508,N_47320,N_47199);
or U48509 (N_48509,N_46074,N_47124);
xnor U48510 (N_48510,N_46443,N_46750);
xor U48511 (N_48511,N_45830,N_45697);
nand U48512 (N_48512,N_47423,N_46201);
or U48513 (N_48513,N_45841,N_46270);
or U48514 (N_48514,N_45411,N_45409);
xor U48515 (N_48515,N_46839,N_45706);
xnor U48516 (N_48516,N_47104,N_45134);
nand U48517 (N_48517,N_45848,N_47288);
nand U48518 (N_48518,N_45607,N_46832);
nor U48519 (N_48519,N_47410,N_45105);
nand U48520 (N_48520,N_46875,N_46487);
xor U48521 (N_48521,N_45443,N_45757);
xor U48522 (N_48522,N_47152,N_46256);
or U48523 (N_48523,N_46649,N_45089);
nand U48524 (N_48524,N_47328,N_46667);
nand U48525 (N_48525,N_45002,N_45483);
nand U48526 (N_48526,N_46599,N_45372);
and U48527 (N_48527,N_45328,N_46188);
nand U48528 (N_48528,N_47153,N_46292);
nand U48529 (N_48529,N_47047,N_47066);
or U48530 (N_48530,N_46679,N_45721);
xor U48531 (N_48531,N_47361,N_45709);
nand U48532 (N_48532,N_47222,N_45350);
or U48533 (N_48533,N_45150,N_45487);
and U48534 (N_48534,N_46148,N_46836);
or U48535 (N_48535,N_45618,N_46194);
nor U48536 (N_48536,N_45690,N_47129);
nand U48537 (N_48537,N_45554,N_46170);
nor U48538 (N_48538,N_46281,N_47085);
or U48539 (N_48539,N_45113,N_45202);
and U48540 (N_48540,N_46796,N_46243);
and U48541 (N_48541,N_45915,N_47437);
xor U48542 (N_48542,N_46554,N_47374);
xor U48543 (N_48543,N_45515,N_47484);
and U48544 (N_48544,N_46713,N_46060);
xnor U48545 (N_48545,N_45905,N_45936);
and U48546 (N_48546,N_46022,N_47394);
xnor U48547 (N_48547,N_45810,N_46960);
nand U48548 (N_48548,N_46919,N_45132);
nand U48549 (N_48549,N_46043,N_47477);
xor U48550 (N_48550,N_45674,N_45739);
and U48551 (N_48551,N_45735,N_45153);
nor U48552 (N_48552,N_46992,N_45694);
or U48553 (N_48553,N_45495,N_46614);
nor U48554 (N_48554,N_46542,N_46534);
nand U48555 (N_48555,N_47205,N_46364);
and U48556 (N_48556,N_46703,N_47371);
or U48557 (N_48557,N_45370,N_45009);
nor U48558 (N_48558,N_46205,N_45656);
and U48559 (N_48559,N_47115,N_47402);
and U48560 (N_48560,N_47461,N_46079);
xor U48561 (N_48561,N_45664,N_46745);
nand U48562 (N_48562,N_46462,N_45834);
nand U48563 (N_48563,N_47103,N_46938);
or U48564 (N_48564,N_46175,N_45214);
or U48565 (N_48565,N_45467,N_46222);
and U48566 (N_48566,N_47252,N_45176);
nor U48567 (N_48567,N_45987,N_47332);
or U48568 (N_48568,N_45602,N_45397);
and U48569 (N_48569,N_45536,N_45228);
nor U48570 (N_48570,N_47311,N_46246);
nand U48571 (N_48571,N_47069,N_45020);
or U48572 (N_48572,N_46790,N_45399);
xnor U48573 (N_48573,N_46844,N_45892);
or U48574 (N_48574,N_46143,N_47099);
xor U48575 (N_48575,N_47493,N_45619);
xnor U48576 (N_48576,N_46435,N_46446);
nand U48577 (N_48577,N_46018,N_45363);
nand U48578 (N_48578,N_46249,N_46202);
and U48579 (N_48579,N_46236,N_45990);
or U48580 (N_48580,N_47308,N_47215);
nor U48581 (N_48581,N_47335,N_46663);
and U48582 (N_48582,N_47385,N_45520);
and U48583 (N_48583,N_47492,N_46687);
nand U48584 (N_48584,N_47444,N_46652);
or U48585 (N_48585,N_45583,N_46879);
xor U48586 (N_48586,N_46684,N_47466);
nor U48587 (N_48587,N_45083,N_46341);
nor U48588 (N_48588,N_46892,N_47412);
or U48589 (N_48589,N_45402,N_47442);
and U48590 (N_48590,N_46780,N_46743);
nand U48591 (N_48591,N_47377,N_46683);
or U48592 (N_48592,N_46518,N_45071);
nand U48593 (N_48593,N_47154,N_45396);
xor U48594 (N_48594,N_46984,N_45982);
xor U48595 (N_48595,N_46529,N_47421);
xnor U48596 (N_48596,N_46321,N_47307);
or U48597 (N_48597,N_46775,N_45805);
or U48598 (N_48598,N_45277,N_45748);
nor U48599 (N_48599,N_46931,N_45814);
xnor U48600 (N_48600,N_47464,N_46234);
and U48601 (N_48601,N_46891,N_45025);
nand U48602 (N_48602,N_46356,N_46070);
and U48603 (N_48603,N_46818,N_46395);
nor U48604 (N_48604,N_46304,N_46486);
or U48605 (N_48605,N_45433,N_45591);
xor U48606 (N_48606,N_46348,N_46362);
nor U48607 (N_48607,N_45177,N_45775);
nand U48608 (N_48608,N_46144,N_45716);
or U48609 (N_48609,N_45252,N_46820);
nand U48610 (N_48610,N_46979,N_45579);
or U48611 (N_48611,N_46752,N_45847);
xor U48612 (N_48612,N_46396,N_45193);
or U48613 (N_48613,N_46541,N_45902);
or U48614 (N_48614,N_46114,N_46739);
or U48615 (N_48615,N_46991,N_46794);
or U48616 (N_48616,N_47343,N_46269);
xor U48617 (N_48617,N_46164,N_45683);
xor U48618 (N_48618,N_47234,N_47097);
nand U48619 (N_48619,N_45884,N_45650);
and U48620 (N_48620,N_47162,N_46017);
nor U48621 (N_48621,N_47376,N_47281);
or U48622 (N_48622,N_47297,N_46208);
xnor U48623 (N_48623,N_47417,N_45904);
xor U48624 (N_48624,N_46537,N_45692);
nor U48625 (N_48625,N_45968,N_46812);
and U48626 (N_48626,N_45643,N_46597);
or U48627 (N_48627,N_45216,N_46071);
or U48628 (N_48628,N_47020,N_46738);
xnor U48629 (N_48629,N_45974,N_45351);
and U48630 (N_48630,N_46417,N_46370);
xor U48631 (N_48631,N_47042,N_46503);
and U48632 (N_48632,N_46087,N_45054);
nand U48633 (N_48633,N_47386,N_45104);
and U48634 (N_48634,N_47456,N_45989);
nand U48635 (N_48635,N_46355,N_46138);
xnor U48636 (N_48636,N_47089,N_47052);
nand U48637 (N_48637,N_46097,N_45192);
or U48638 (N_48638,N_46604,N_45570);
nor U48639 (N_48639,N_47425,N_46927);
xor U48640 (N_48640,N_45661,N_45938);
xnor U48641 (N_48641,N_45125,N_46549);
nor U48642 (N_48642,N_46788,N_46161);
nand U48643 (N_48643,N_45017,N_45728);
nor U48644 (N_48644,N_46648,N_46117);
xor U48645 (N_48645,N_45737,N_46331);
nor U48646 (N_48646,N_45117,N_46706);
and U48647 (N_48647,N_46936,N_46368);
nand U48648 (N_48648,N_46085,N_47088);
xor U48649 (N_48649,N_45297,N_46027);
and U48650 (N_48650,N_47012,N_46004);
nor U48651 (N_48651,N_45897,N_45076);
nand U48652 (N_48652,N_45172,N_45251);
nand U48653 (N_48653,N_46922,N_45965);
and U48654 (N_48654,N_45110,N_46899);
xor U48655 (N_48655,N_45107,N_47472);
nor U48656 (N_48656,N_46876,N_46251);
xor U48657 (N_48657,N_46231,N_46177);
nand U48658 (N_48658,N_46041,N_45751);
nand U48659 (N_48659,N_45667,N_45130);
nand U48660 (N_48660,N_47193,N_45534);
xor U48661 (N_48661,N_45801,N_45639);
and U48662 (N_48662,N_45940,N_45080);
nor U48663 (N_48663,N_46524,N_45086);
xnor U48664 (N_48664,N_45893,N_45223);
nand U48665 (N_48665,N_45798,N_46198);
and U48666 (N_48666,N_46611,N_45112);
nor U48667 (N_48667,N_46328,N_46947);
nand U48668 (N_48668,N_46675,N_47142);
nand U48669 (N_48669,N_45586,N_45919);
xnor U48670 (N_48670,N_46391,N_47241);
or U48671 (N_48671,N_47325,N_45091);
nor U48672 (N_48672,N_46026,N_45852);
nor U48673 (N_48673,N_47133,N_46755);
or U48674 (N_48674,N_45636,N_47469);
or U48675 (N_48675,N_45627,N_45332);
xor U48676 (N_48676,N_46115,N_45239);
and U48677 (N_48677,N_45205,N_46601);
xnor U48678 (N_48678,N_47369,N_45301);
and U48679 (N_48679,N_47214,N_46245);
or U48680 (N_48680,N_47290,N_45119);
xnor U48681 (N_48681,N_45184,N_45778);
nand U48682 (N_48682,N_46782,N_47035);
nor U48683 (N_48683,N_46972,N_46797);
nand U48684 (N_48684,N_45907,N_47443);
nand U48685 (N_48685,N_45084,N_47305);
nor U48686 (N_48686,N_46262,N_46949);
nor U48687 (N_48687,N_47480,N_46306);
nand U48688 (N_48688,N_46191,N_47419);
xnor U48689 (N_48689,N_46617,N_46073);
and U48690 (N_48690,N_46465,N_46779);
nor U48691 (N_48691,N_45343,N_46946);
or U48692 (N_48692,N_46732,N_45410);
xnor U48693 (N_48693,N_45970,N_47223);
nor U48694 (N_48694,N_45763,N_45420);
and U48695 (N_48695,N_45492,N_46493);
nand U48696 (N_48696,N_45473,N_46974);
xnor U48697 (N_48697,N_45969,N_46296);
and U48698 (N_48698,N_45588,N_46103);
nor U48699 (N_48699,N_45095,N_45166);
nand U48700 (N_48700,N_46040,N_46233);
xor U48701 (N_48701,N_45212,N_46793);
nand U48702 (N_48702,N_47121,N_46699);
nand U48703 (N_48703,N_45657,N_46666);
nor U48704 (N_48704,N_45741,N_46543);
nor U48705 (N_48705,N_46533,N_45809);
xor U48706 (N_48706,N_46951,N_46159);
nand U48707 (N_48707,N_45008,N_46906);
and U48708 (N_48708,N_46928,N_46113);
nand U48709 (N_48709,N_46948,N_46704);
or U48710 (N_48710,N_45131,N_45943);
or U48711 (N_48711,N_47105,N_45532);
xnor U48712 (N_48712,N_47061,N_45049);
xor U48713 (N_48713,N_46252,N_45353);
xor U48714 (N_48714,N_46195,N_46118);
xor U48715 (N_48715,N_47166,N_47460);
xnor U48716 (N_48716,N_45108,N_45288);
xnor U48717 (N_48717,N_46034,N_47060);
xnor U48718 (N_48718,N_46806,N_46540);
or U48719 (N_48719,N_45194,N_46484);
nand U48720 (N_48720,N_45161,N_46317);
xnor U48721 (N_48721,N_45255,N_45510);
or U48722 (N_48722,N_46773,N_46127);
xnor U48723 (N_48723,N_47075,N_45665);
or U48724 (N_48724,N_45448,N_46510);
nand U48725 (N_48725,N_46450,N_46511);
nand U48726 (N_48726,N_45679,N_46342);
xnor U48727 (N_48727,N_46558,N_46975);
and U48728 (N_48728,N_46582,N_45141);
or U48729 (N_48729,N_45320,N_46015);
and U48730 (N_48730,N_45918,N_46898);
and U48731 (N_48731,N_46474,N_46729);
xnor U48732 (N_48732,N_47094,N_45993);
nor U48733 (N_48733,N_46010,N_45204);
nand U48734 (N_48734,N_46467,N_47340);
or U48735 (N_48735,N_45577,N_46887);
nand U48736 (N_48736,N_46491,N_46774);
or U48737 (N_48737,N_47001,N_46333);
or U48738 (N_48738,N_46521,N_46440);
and U48739 (N_48739,N_47050,N_45587);
xnor U48740 (N_48740,N_45140,N_47434);
xor U48741 (N_48741,N_46241,N_46258);
or U48742 (N_48742,N_46137,N_47398);
or U48743 (N_48743,N_46682,N_45085);
or U48744 (N_48744,N_46852,N_47267);
nand U48745 (N_48745,N_47221,N_46089);
or U48746 (N_48746,N_45518,N_46583);
and U48747 (N_48747,N_47192,N_46189);
and U48748 (N_48748,N_47347,N_45245);
or U48749 (N_48749,N_45224,N_45133);
or U48750 (N_48750,N_46428,N_45831);
xnor U48751 (N_48751,N_46004,N_45730);
or U48752 (N_48752,N_47083,N_45170);
or U48753 (N_48753,N_45058,N_45348);
xor U48754 (N_48754,N_45032,N_46878);
or U48755 (N_48755,N_46333,N_46891);
and U48756 (N_48756,N_45959,N_46870);
nand U48757 (N_48757,N_46251,N_46999);
and U48758 (N_48758,N_47054,N_46955);
nand U48759 (N_48759,N_47152,N_47260);
or U48760 (N_48760,N_47455,N_45179);
xnor U48761 (N_48761,N_46032,N_45437);
and U48762 (N_48762,N_45250,N_46596);
and U48763 (N_48763,N_47286,N_45925);
nor U48764 (N_48764,N_47326,N_45753);
and U48765 (N_48765,N_47470,N_45668);
nand U48766 (N_48766,N_46722,N_46769);
nor U48767 (N_48767,N_46238,N_47112);
nor U48768 (N_48768,N_46623,N_46446);
or U48769 (N_48769,N_46010,N_46932);
or U48770 (N_48770,N_46049,N_45024);
nor U48771 (N_48771,N_45392,N_46570);
nor U48772 (N_48772,N_46203,N_46528);
nor U48773 (N_48773,N_46197,N_46218);
nand U48774 (N_48774,N_45377,N_47179);
or U48775 (N_48775,N_45048,N_47120);
nor U48776 (N_48776,N_45356,N_46752);
and U48777 (N_48777,N_46553,N_46579);
xor U48778 (N_48778,N_46099,N_46164);
or U48779 (N_48779,N_45406,N_46749);
nor U48780 (N_48780,N_46226,N_46298);
nand U48781 (N_48781,N_47490,N_46837);
xor U48782 (N_48782,N_45556,N_46576);
or U48783 (N_48783,N_46185,N_45624);
or U48784 (N_48784,N_47399,N_46097);
or U48785 (N_48785,N_45172,N_46265);
nand U48786 (N_48786,N_45521,N_45974);
xor U48787 (N_48787,N_47443,N_45130);
and U48788 (N_48788,N_46040,N_47397);
nor U48789 (N_48789,N_46761,N_45163);
nor U48790 (N_48790,N_46767,N_45722);
xnor U48791 (N_48791,N_46276,N_46250);
nor U48792 (N_48792,N_46687,N_46904);
or U48793 (N_48793,N_45747,N_46369);
nand U48794 (N_48794,N_45028,N_45869);
or U48795 (N_48795,N_46379,N_47344);
or U48796 (N_48796,N_46568,N_47160);
nand U48797 (N_48797,N_46233,N_47268);
or U48798 (N_48798,N_47487,N_46833);
or U48799 (N_48799,N_45792,N_45582);
nand U48800 (N_48800,N_45908,N_46052);
nor U48801 (N_48801,N_47234,N_47103);
xnor U48802 (N_48802,N_45234,N_46248);
or U48803 (N_48803,N_45722,N_45258);
or U48804 (N_48804,N_47446,N_45561);
nor U48805 (N_48805,N_46392,N_46167);
or U48806 (N_48806,N_45984,N_47229);
nand U48807 (N_48807,N_45679,N_46786);
nand U48808 (N_48808,N_45867,N_47419);
xnor U48809 (N_48809,N_47193,N_45401);
nand U48810 (N_48810,N_47031,N_45451);
nor U48811 (N_48811,N_45208,N_46287);
or U48812 (N_48812,N_45485,N_46448);
and U48813 (N_48813,N_46477,N_45932);
xnor U48814 (N_48814,N_46733,N_45732);
nor U48815 (N_48815,N_45274,N_45289);
xor U48816 (N_48816,N_45086,N_45838);
xor U48817 (N_48817,N_46127,N_47284);
xnor U48818 (N_48818,N_46383,N_46899);
or U48819 (N_48819,N_46248,N_45205);
or U48820 (N_48820,N_47441,N_46857);
nand U48821 (N_48821,N_45130,N_47127);
nor U48822 (N_48822,N_46804,N_46550);
and U48823 (N_48823,N_46130,N_45889);
xnor U48824 (N_48824,N_45152,N_46140);
and U48825 (N_48825,N_45721,N_46107);
or U48826 (N_48826,N_46961,N_46518);
or U48827 (N_48827,N_47462,N_47219);
and U48828 (N_48828,N_46128,N_45037);
and U48829 (N_48829,N_47155,N_46352);
and U48830 (N_48830,N_45365,N_46291);
and U48831 (N_48831,N_45883,N_47309);
or U48832 (N_48832,N_46042,N_47080);
or U48833 (N_48833,N_46544,N_45260);
nor U48834 (N_48834,N_45468,N_46946);
or U48835 (N_48835,N_46531,N_46229);
and U48836 (N_48836,N_45914,N_46115);
or U48837 (N_48837,N_47064,N_45113);
and U48838 (N_48838,N_46948,N_45139);
nand U48839 (N_48839,N_45620,N_45984);
and U48840 (N_48840,N_45593,N_45258);
or U48841 (N_48841,N_47033,N_47152);
nand U48842 (N_48842,N_46490,N_45773);
and U48843 (N_48843,N_47293,N_46581);
nand U48844 (N_48844,N_46780,N_45246);
and U48845 (N_48845,N_45107,N_46407);
and U48846 (N_48846,N_45105,N_45087);
or U48847 (N_48847,N_45177,N_47166);
nand U48848 (N_48848,N_46666,N_46963);
xor U48849 (N_48849,N_45040,N_45258);
nand U48850 (N_48850,N_47140,N_45666);
xor U48851 (N_48851,N_45766,N_45902);
nand U48852 (N_48852,N_47426,N_45867);
nand U48853 (N_48853,N_45190,N_46964);
xnor U48854 (N_48854,N_46093,N_46191);
or U48855 (N_48855,N_46882,N_46797);
nor U48856 (N_48856,N_45862,N_47110);
xnor U48857 (N_48857,N_45717,N_45096);
or U48858 (N_48858,N_46335,N_47104);
xnor U48859 (N_48859,N_45320,N_46993);
or U48860 (N_48860,N_46992,N_45976);
xor U48861 (N_48861,N_47294,N_45022);
or U48862 (N_48862,N_45018,N_46873);
nor U48863 (N_48863,N_45192,N_45219);
and U48864 (N_48864,N_45462,N_47297);
and U48865 (N_48865,N_47011,N_45252);
xnor U48866 (N_48866,N_46878,N_45385);
nor U48867 (N_48867,N_46089,N_45138);
and U48868 (N_48868,N_45374,N_45053);
nor U48869 (N_48869,N_47363,N_45343);
and U48870 (N_48870,N_45108,N_45313);
and U48871 (N_48871,N_45899,N_46913);
xnor U48872 (N_48872,N_46540,N_45426);
and U48873 (N_48873,N_47105,N_45267);
xnor U48874 (N_48874,N_45486,N_45468);
nor U48875 (N_48875,N_47410,N_46834);
or U48876 (N_48876,N_47174,N_45505);
and U48877 (N_48877,N_47195,N_46720);
nand U48878 (N_48878,N_45536,N_46866);
and U48879 (N_48879,N_46001,N_46392);
nand U48880 (N_48880,N_45111,N_46660);
nor U48881 (N_48881,N_47067,N_46002);
or U48882 (N_48882,N_46962,N_45422);
nor U48883 (N_48883,N_45377,N_47254);
xor U48884 (N_48884,N_45396,N_46269);
nand U48885 (N_48885,N_45646,N_45994);
and U48886 (N_48886,N_45791,N_46907);
or U48887 (N_48887,N_46669,N_47118);
xnor U48888 (N_48888,N_45540,N_46115);
and U48889 (N_48889,N_46376,N_45708);
xnor U48890 (N_48890,N_46523,N_45071);
and U48891 (N_48891,N_45337,N_46379);
nor U48892 (N_48892,N_47091,N_46854);
nand U48893 (N_48893,N_46343,N_45050);
xor U48894 (N_48894,N_46813,N_45462);
nor U48895 (N_48895,N_45019,N_45159);
or U48896 (N_48896,N_46046,N_45898);
nor U48897 (N_48897,N_45824,N_47495);
nor U48898 (N_48898,N_45642,N_46000);
xor U48899 (N_48899,N_46626,N_45860);
or U48900 (N_48900,N_45531,N_46041);
nand U48901 (N_48901,N_45527,N_47078);
or U48902 (N_48902,N_45076,N_45239);
and U48903 (N_48903,N_45967,N_47252);
xnor U48904 (N_48904,N_45143,N_45693);
xnor U48905 (N_48905,N_46790,N_45315);
nand U48906 (N_48906,N_47290,N_47399);
and U48907 (N_48907,N_46492,N_45975);
nor U48908 (N_48908,N_47258,N_46595);
nor U48909 (N_48909,N_47421,N_46309);
xor U48910 (N_48910,N_45720,N_45177);
and U48911 (N_48911,N_47008,N_46252);
nor U48912 (N_48912,N_45909,N_46663);
xor U48913 (N_48913,N_45223,N_45336);
nor U48914 (N_48914,N_47122,N_47059);
xnor U48915 (N_48915,N_45112,N_45366);
nand U48916 (N_48916,N_45948,N_47487);
or U48917 (N_48917,N_46205,N_47291);
or U48918 (N_48918,N_46086,N_45491);
and U48919 (N_48919,N_46809,N_46697);
nor U48920 (N_48920,N_47449,N_45745);
or U48921 (N_48921,N_45955,N_47082);
xor U48922 (N_48922,N_47136,N_46803);
nand U48923 (N_48923,N_46201,N_46203);
xnor U48924 (N_48924,N_45264,N_45159);
and U48925 (N_48925,N_45034,N_45100);
xor U48926 (N_48926,N_46016,N_46735);
nand U48927 (N_48927,N_47453,N_47002);
nor U48928 (N_48928,N_45795,N_45192);
nand U48929 (N_48929,N_45601,N_45176);
xor U48930 (N_48930,N_45752,N_46239);
nand U48931 (N_48931,N_46423,N_45061);
and U48932 (N_48932,N_45557,N_46369);
nor U48933 (N_48933,N_46330,N_45870);
or U48934 (N_48934,N_45534,N_45154);
nand U48935 (N_48935,N_47401,N_45414);
nor U48936 (N_48936,N_45720,N_47246);
xor U48937 (N_48937,N_46803,N_46541);
nand U48938 (N_48938,N_47342,N_45122);
nand U48939 (N_48939,N_47026,N_45221);
xor U48940 (N_48940,N_45764,N_45722);
and U48941 (N_48941,N_47070,N_47484);
and U48942 (N_48942,N_46496,N_47468);
nand U48943 (N_48943,N_46131,N_46866);
and U48944 (N_48944,N_47368,N_47399);
nand U48945 (N_48945,N_45818,N_46703);
and U48946 (N_48946,N_45830,N_47449);
nand U48947 (N_48947,N_47330,N_47239);
and U48948 (N_48948,N_46370,N_46353);
nand U48949 (N_48949,N_47254,N_46640);
nand U48950 (N_48950,N_45602,N_45286);
nor U48951 (N_48951,N_46404,N_45140);
nand U48952 (N_48952,N_45113,N_45690);
or U48953 (N_48953,N_47242,N_46606);
nand U48954 (N_48954,N_46802,N_46432);
or U48955 (N_48955,N_45468,N_46955);
xnor U48956 (N_48956,N_45112,N_45530);
nor U48957 (N_48957,N_46166,N_46595);
xor U48958 (N_48958,N_45634,N_46620);
or U48959 (N_48959,N_45318,N_45658);
xnor U48960 (N_48960,N_47067,N_47092);
xnor U48961 (N_48961,N_47497,N_46306);
xor U48962 (N_48962,N_45607,N_47340);
nor U48963 (N_48963,N_47173,N_46830);
or U48964 (N_48964,N_46089,N_46849);
nand U48965 (N_48965,N_46804,N_45888);
and U48966 (N_48966,N_46445,N_47096);
and U48967 (N_48967,N_46117,N_45096);
xnor U48968 (N_48968,N_45891,N_46640);
or U48969 (N_48969,N_45322,N_47267);
nor U48970 (N_48970,N_46403,N_45350);
xnor U48971 (N_48971,N_46751,N_47289);
xnor U48972 (N_48972,N_46497,N_46307);
xnor U48973 (N_48973,N_45252,N_46917);
nand U48974 (N_48974,N_45519,N_45322);
xnor U48975 (N_48975,N_46410,N_47328);
xnor U48976 (N_48976,N_47322,N_46528);
and U48977 (N_48977,N_47056,N_45135);
nor U48978 (N_48978,N_47086,N_47267);
nor U48979 (N_48979,N_45681,N_45086);
and U48980 (N_48980,N_46960,N_46028);
nand U48981 (N_48981,N_46617,N_46544);
or U48982 (N_48982,N_47310,N_45961);
and U48983 (N_48983,N_46776,N_45443);
and U48984 (N_48984,N_46907,N_47093);
nand U48985 (N_48985,N_46477,N_45836);
nor U48986 (N_48986,N_45575,N_46898);
and U48987 (N_48987,N_46789,N_45258);
nand U48988 (N_48988,N_47265,N_47165);
xor U48989 (N_48989,N_46304,N_46811);
or U48990 (N_48990,N_47414,N_45301);
nand U48991 (N_48991,N_45236,N_47247);
and U48992 (N_48992,N_46434,N_46119);
nor U48993 (N_48993,N_47082,N_45176);
xnor U48994 (N_48994,N_47074,N_47344);
nand U48995 (N_48995,N_46092,N_45018);
and U48996 (N_48996,N_45346,N_45667);
or U48997 (N_48997,N_46488,N_45748);
and U48998 (N_48998,N_45269,N_46910);
and U48999 (N_48999,N_45161,N_45546);
xor U49000 (N_49000,N_46668,N_45492);
nand U49001 (N_49001,N_46594,N_45834);
nand U49002 (N_49002,N_45044,N_46799);
nor U49003 (N_49003,N_47204,N_46577);
and U49004 (N_49004,N_45323,N_45673);
and U49005 (N_49005,N_45008,N_47265);
and U49006 (N_49006,N_46608,N_46716);
nand U49007 (N_49007,N_46058,N_47017);
and U49008 (N_49008,N_46183,N_46915);
and U49009 (N_49009,N_47421,N_46175);
nor U49010 (N_49010,N_46944,N_45066);
nor U49011 (N_49011,N_46180,N_47185);
xnor U49012 (N_49012,N_47392,N_45797);
nand U49013 (N_49013,N_45614,N_45867);
nand U49014 (N_49014,N_45862,N_45189);
and U49015 (N_49015,N_46099,N_45778);
and U49016 (N_49016,N_47315,N_45164);
and U49017 (N_49017,N_45012,N_46965);
or U49018 (N_49018,N_46673,N_46573);
or U49019 (N_49019,N_45009,N_46801);
or U49020 (N_49020,N_46355,N_45332);
nor U49021 (N_49021,N_46059,N_45886);
and U49022 (N_49022,N_45649,N_45743);
xor U49023 (N_49023,N_45580,N_45085);
xor U49024 (N_49024,N_46240,N_46352);
and U49025 (N_49025,N_45046,N_47152);
or U49026 (N_49026,N_46957,N_45998);
or U49027 (N_49027,N_46354,N_45473);
and U49028 (N_49028,N_46474,N_47443);
xnor U49029 (N_49029,N_46437,N_46386);
or U49030 (N_49030,N_46183,N_46958);
nor U49031 (N_49031,N_45135,N_45248);
nor U49032 (N_49032,N_47074,N_47173);
xor U49033 (N_49033,N_47425,N_46397);
xnor U49034 (N_49034,N_46844,N_45338);
or U49035 (N_49035,N_46832,N_45769);
or U49036 (N_49036,N_46519,N_45296);
nor U49037 (N_49037,N_45524,N_46980);
or U49038 (N_49038,N_45640,N_45204);
nand U49039 (N_49039,N_47095,N_45992);
nor U49040 (N_49040,N_46445,N_46603);
nand U49041 (N_49041,N_47011,N_46979);
or U49042 (N_49042,N_45578,N_45720);
nand U49043 (N_49043,N_46729,N_46112);
nor U49044 (N_49044,N_46394,N_45070);
nor U49045 (N_49045,N_47217,N_46391);
or U49046 (N_49046,N_46476,N_46129);
or U49047 (N_49047,N_45909,N_46309);
or U49048 (N_49048,N_47374,N_45743);
or U49049 (N_49049,N_46796,N_45435);
nand U49050 (N_49050,N_46546,N_46467);
and U49051 (N_49051,N_47442,N_45217);
or U49052 (N_49052,N_47204,N_45736);
xor U49053 (N_49053,N_47239,N_47493);
or U49054 (N_49054,N_46134,N_46188);
nand U49055 (N_49055,N_46517,N_45612);
nand U49056 (N_49056,N_46460,N_45427);
and U49057 (N_49057,N_46558,N_45558);
xor U49058 (N_49058,N_45790,N_45805);
and U49059 (N_49059,N_45662,N_45986);
and U49060 (N_49060,N_47451,N_45744);
or U49061 (N_49061,N_46104,N_45679);
and U49062 (N_49062,N_47014,N_46332);
nor U49063 (N_49063,N_47432,N_47097);
and U49064 (N_49064,N_47366,N_46795);
xnor U49065 (N_49065,N_46930,N_46391);
or U49066 (N_49066,N_45322,N_46270);
and U49067 (N_49067,N_45644,N_46529);
nand U49068 (N_49068,N_45780,N_46107);
or U49069 (N_49069,N_46242,N_45419);
and U49070 (N_49070,N_45065,N_46121);
nand U49071 (N_49071,N_45464,N_45487);
nand U49072 (N_49072,N_45867,N_47256);
and U49073 (N_49073,N_45662,N_46922);
and U49074 (N_49074,N_45781,N_46829);
xnor U49075 (N_49075,N_46657,N_45066);
nand U49076 (N_49076,N_47234,N_45203);
nor U49077 (N_49077,N_46899,N_45498);
nand U49078 (N_49078,N_46543,N_46605);
or U49079 (N_49079,N_47403,N_46335);
nor U49080 (N_49080,N_45579,N_46883);
and U49081 (N_49081,N_45681,N_45993);
and U49082 (N_49082,N_45683,N_45846);
and U49083 (N_49083,N_46383,N_45249);
nor U49084 (N_49084,N_46424,N_45657);
and U49085 (N_49085,N_45189,N_46021);
xor U49086 (N_49086,N_46657,N_45356);
xnor U49087 (N_49087,N_47154,N_47132);
nor U49088 (N_49088,N_45338,N_47147);
nand U49089 (N_49089,N_46563,N_46555);
or U49090 (N_49090,N_45226,N_45428);
and U49091 (N_49091,N_46029,N_46764);
xor U49092 (N_49092,N_45608,N_47295);
or U49093 (N_49093,N_47071,N_45952);
or U49094 (N_49094,N_46252,N_45320);
nor U49095 (N_49095,N_46395,N_46180);
nor U49096 (N_49096,N_45569,N_45130);
nand U49097 (N_49097,N_45616,N_46493);
or U49098 (N_49098,N_46036,N_46218);
or U49099 (N_49099,N_47117,N_45817);
nor U49100 (N_49100,N_45395,N_46096);
nor U49101 (N_49101,N_45353,N_46398);
xnor U49102 (N_49102,N_46037,N_46767);
xor U49103 (N_49103,N_45092,N_46476);
nor U49104 (N_49104,N_45533,N_45279);
and U49105 (N_49105,N_46674,N_45544);
or U49106 (N_49106,N_46130,N_46723);
and U49107 (N_49107,N_45505,N_45358);
nor U49108 (N_49108,N_45398,N_47403);
nor U49109 (N_49109,N_45471,N_45312);
or U49110 (N_49110,N_46488,N_46518);
or U49111 (N_49111,N_46912,N_45299);
nor U49112 (N_49112,N_47399,N_46264);
nand U49113 (N_49113,N_47363,N_46161);
nor U49114 (N_49114,N_45254,N_46315);
nor U49115 (N_49115,N_46754,N_47182);
or U49116 (N_49116,N_47336,N_47298);
nor U49117 (N_49117,N_45861,N_46782);
nor U49118 (N_49118,N_45766,N_46829);
nand U49119 (N_49119,N_47359,N_47338);
nand U49120 (N_49120,N_45799,N_45770);
xor U49121 (N_49121,N_46643,N_46066);
or U49122 (N_49122,N_46079,N_47260);
or U49123 (N_49123,N_46047,N_46483);
xor U49124 (N_49124,N_47349,N_47018);
nand U49125 (N_49125,N_46025,N_47368);
nor U49126 (N_49126,N_45321,N_46309);
or U49127 (N_49127,N_46722,N_46844);
or U49128 (N_49128,N_46258,N_46304);
xnor U49129 (N_49129,N_46807,N_45935);
xnor U49130 (N_49130,N_47468,N_46427);
nand U49131 (N_49131,N_45224,N_46521);
and U49132 (N_49132,N_46680,N_47123);
and U49133 (N_49133,N_47205,N_45717);
and U49134 (N_49134,N_46212,N_46330);
nor U49135 (N_49135,N_45361,N_45090);
or U49136 (N_49136,N_47287,N_47303);
and U49137 (N_49137,N_45665,N_45350);
and U49138 (N_49138,N_45025,N_46384);
and U49139 (N_49139,N_47065,N_46811);
nand U49140 (N_49140,N_46769,N_45751);
or U49141 (N_49141,N_45479,N_46690);
xnor U49142 (N_49142,N_46536,N_45366);
and U49143 (N_49143,N_47026,N_47394);
nor U49144 (N_49144,N_45865,N_46535);
or U49145 (N_49145,N_45741,N_47118);
or U49146 (N_49146,N_47433,N_46490);
xor U49147 (N_49147,N_45667,N_47034);
nor U49148 (N_49148,N_46456,N_45115);
nand U49149 (N_49149,N_45987,N_45984);
or U49150 (N_49150,N_46025,N_47068);
nor U49151 (N_49151,N_46216,N_45470);
nor U49152 (N_49152,N_45269,N_45912);
nand U49153 (N_49153,N_47409,N_46340);
and U49154 (N_49154,N_46595,N_46421);
nand U49155 (N_49155,N_47199,N_46965);
and U49156 (N_49156,N_46545,N_45613);
nor U49157 (N_49157,N_45066,N_46430);
nor U49158 (N_49158,N_46297,N_47152);
nand U49159 (N_49159,N_45747,N_47268);
and U49160 (N_49160,N_47020,N_47001);
and U49161 (N_49161,N_45691,N_47171);
or U49162 (N_49162,N_47163,N_47113);
nor U49163 (N_49163,N_47207,N_45995);
nand U49164 (N_49164,N_47098,N_46538);
and U49165 (N_49165,N_46674,N_45133);
nor U49166 (N_49166,N_46689,N_46264);
nand U49167 (N_49167,N_46788,N_47366);
xor U49168 (N_49168,N_46255,N_45047);
nand U49169 (N_49169,N_46868,N_46370);
and U49170 (N_49170,N_45513,N_47047);
nor U49171 (N_49171,N_46655,N_45737);
nor U49172 (N_49172,N_46519,N_47257);
nand U49173 (N_49173,N_45814,N_47269);
xor U49174 (N_49174,N_46816,N_45600);
nand U49175 (N_49175,N_46739,N_47076);
nand U49176 (N_49176,N_47121,N_47119);
and U49177 (N_49177,N_45928,N_46905);
nand U49178 (N_49178,N_46987,N_46174);
or U49179 (N_49179,N_45803,N_46312);
or U49180 (N_49180,N_46276,N_45384);
or U49181 (N_49181,N_46456,N_45951);
nand U49182 (N_49182,N_46707,N_45381);
xor U49183 (N_49183,N_46991,N_46097);
xor U49184 (N_49184,N_47433,N_45769);
or U49185 (N_49185,N_45211,N_45599);
nand U49186 (N_49186,N_45404,N_45690);
and U49187 (N_49187,N_46612,N_46358);
nor U49188 (N_49188,N_46670,N_46150);
nor U49189 (N_49189,N_45539,N_47205);
or U49190 (N_49190,N_45198,N_45704);
nand U49191 (N_49191,N_47053,N_45193);
and U49192 (N_49192,N_46101,N_46730);
or U49193 (N_49193,N_46692,N_47052);
nor U49194 (N_49194,N_46249,N_45251);
nand U49195 (N_49195,N_45280,N_47410);
nor U49196 (N_49196,N_47075,N_45576);
nand U49197 (N_49197,N_45912,N_46548);
or U49198 (N_49198,N_46675,N_45143);
or U49199 (N_49199,N_45996,N_45658);
nand U49200 (N_49200,N_46465,N_45920);
or U49201 (N_49201,N_45219,N_45571);
or U49202 (N_49202,N_45469,N_45739);
and U49203 (N_49203,N_46745,N_45286);
or U49204 (N_49204,N_45937,N_46618);
or U49205 (N_49205,N_46365,N_45073);
nor U49206 (N_49206,N_46646,N_45667);
nand U49207 (N_49207,N_45709,N_45391);
nand U49208 (N_49208,N_45291,N_45557);
and U49209 (N_49209,N_45998,N_47021);
nand U49210 (N_49210,N_46463,N_46556);
and U49211 (N_49211,N_47402,N_47212);
and U49212 (N_49212,N_46193,N_46146);
xor U49213 (N_49213,N_46726,N_46897);
and U49214 (N_49214,N_46324,N_46999);
nand U49215 (N_49215,N_46489,N_45466);
and U49216 (N_49216,N_45049,N_46729);
nand U49217 (N_49217,N_46230,N_47020);
xor U49218 (N_49218,N_47033,N_47312);
xnor U49219 (N_49219,N_46823,N_46861);
and U49220 (N_49220,N_46463,N_46165);
xor U49221 (N_49221,N_45744,N_46704);
xor U49222 (N_49222,N_47123,N_46115);
or U49223 (N_49223,N_46291,N_45837);
nand U49224 (N_49224,N_46626,N_45411);
nor U49225 (N_49225,N_45582,N_47284);
xor U49226 (N_49226,N_45014,N_45310);
nand U49227 (N_49227,N_46106,N_46646);
xnor U49228 (N_49228,N_45690,N_45240);
and U49229 (N_49229,N_46473,N_45689);
nor U49230 (N_49230,N_46414,N_45938);
nor U49231 (N_49231,N_45197,N_45238);
and U49232 (N_49232,N_45626,N_45070);
nor U49233 (N_49233,N_46989,N_45229);
xor U49234 (N_49234,N_46591,N_45075);
nand U49235 (N_49235,N_47017,N_46789);
or U49236 (N_49236,N_46264,N_45748);
nor U49237 (N_49237,N_46457,N_47179);
and U49238 (N_49238,N_45404,N_47296);
or U49239 (N_49239,N_45492,N_45591);
nor U49240 (N_49240,N_46868,N_46384);
or U49241 (N_49241,N_45260,N_46203);
and U49242 (N_49242,N_46467,N_47454);
and U49243 (N_49243,N_46755,N_46961);
and U49244 (N_49244,N_45996,N_46461);
nor U49245 (N_49245,N_47035,N_45590);
or U49246 (N_49246,N_45593,N_45804);
xnor U49247 (N_49247,N_46503,N_46658);
or U49248 (N_49248,N_45545,N_45890);
nor U49249 (N_49249,N_47072,N_47063);
nand U49250 (N_49250,N_46360,N_46893);
or U49251 (N_49251,N_46804,N_45535);
and U49252 (N_49252,N_46390,N_47207);
or U49253 (N_49253,N_46886,N_45376);
and U49254 (N_49254,N_45280,N_46763);
and U49255 (N_49255,N_45958,N_45525);
or U49256 (N_49256,N_46274,N_46621);
and U49257 (N_49257,N_46505,N_46975);
xor U49258 (N_49258,N_45569,N_47366);
xnor U49259 (N_49259,N_45062,N_46611);
nor U49260 (N_49260,N_46816,N_46464);
nand U49261 (N_49261,N_47105,N_45721);
and U49262 (N_49262,N_46562,N_47375);
nand U49263 (N_49263,N_46654,N_46332);
and U49264 (N_49264,N_47191,N_46813);
nor U49265 (N_49265,N_45808,N_47409);
nand U49266 (N_49266,N_47089,N_46067);
and U49267 (N_49267,N_46261,N_46078);
xnor U49268 (N_49268,N_46515,N_47036);
or U49269 (N_49269,N_47327,N_46841);
nor U49270 (N_49270,N_45862,N_45879);
nor U49271 (N_49271,N_46814,N_46201);
and U49272 (N_49272,N_46417,N_47308);
nand U49273 (N_49273,N_46950,N_47430);
or U49274 (N_49274,N_45939,N_45923);
nor U49275 (N_49275,N_45088,N_47079);
nor U49276 (N_49276,N_45335,N_46876);
nor U49277 (N_49277,N_45426,N_46035);
nor U49278 (N_49278,N_45648,N_46304);
or U49279 (N_49279,N_45017,N_45837);
xnor U49280 (N_49280,N_46880,N_45745);
xnor U49281 (N_49281,N_46150,N_46630);
and U49282 (N_49282,N_47322,N_45877);
and U49283 (N_49283,N_47364,N_46197);
and U49284 (N_49284,N_45270,N_46017);
nor U49285 (N_49285,N_46148,N_46033);
and U49286 (N_49286,N_45106,N_47469);
nand U49287 (N_49287,N_45445,N_45985);
or U49288 (N_49288,N_45310,N_46081);
nor U49289 (N_49289,N_46380,N_46612);
and U49290 (N_49290,N_45884,N_46358);
and U49291 (N_49291,N_46713,N_45394);
xor U49292 (N_49292,N_45230,N_45850);
nand U49293 (N_49293,N_45491,N_46836);
or U49294 (N_49294,N_46292,N_46491);
nor U49295 (N_49295,N_45898,N_46435);
or U49296 (N_49296,N_47314,N_46576);
or U49297 (N_49297,N_46466,N_45202);
and U49298 (N_49298,N_45045,N_46095);
nor U49299 (N_49299,N_45784,N_45674);
or U49300 (N_49300,N_46036,N_45310);
and U49301 (N_49301,N_46154,N_46579);
nor U49302 (N_49302,N_46685,N_47400);
nand U49303 (N_49303,N_45395,N_45769);
nand U49304 (N_49304,N_47016,N_47277);
or U49305 (N_49305,N_45333,N_46400);
xor U49306 (N_49306,N_47229,N_46180);
xnor U49307 (N_49307,N_46452,N_46657);
and U49308 (N_49308,N_47461,N_46333);
and U49309 (N_49309,N_47134,N_45494);
and U49310 (N_49310,N_46870,N_45718);
xor U49311 (N_49311,N_47478,N_47160);
xnor U49312 (N_49312,N_46289,N_46229);
nor U49313 (N_49313,N_46545,N_45300);
xor U49314 (N_49314,N_45016,N_45112);
xor U49315 (N_49315,N_46972,N_45737);
nor U49316 (N_49316,N_46331,N_46543);
or U49317 (N_49317,N_45610,N_45507);
nand U49318 (N_49318,N_45293,N_47353);
xnor U49319 (N_49319,N_46701,N_45261);
xor U49320 (N_49320,N_47003,N_46325);
nor U49321 (N_49321,N_46412,N_45079);
nor U49322 (N_49322,N_47420,N_45662);
or U49323 (N_49323,N_45012,N_46978);
or U49324 (N_49324,N_46350,N_46262);
nand U49325 (N_49325,N_45664,N_46761);
or U49326 (N_49326,N_46039,N_46158);
and U49327 (N_49327,N_46202,N_46526);
or U49328 (N_49328,N_46278,N_47313);
or U49329 (N_49329,N_45228,N_47468);
xor U49330 (N_49330,N_46093,N_45798);
or U49331 (N_49331,N_45065,N_46576);
xnor U49332 (N_49332,N_46004,N_46139);
or U49333 (N_49333,N_47394,N_45131);
nor U49334 (N_49334,N_45724,N_45567);
xor U49335 (N_49335,N_46694,N_46260);
nand U49336 (N_49336,N_45707,N_47163);
nor U49337 (N_49337,N_45758,N_45456);
xnor U49338 (N_49338,N_46640,N_46328);
and U49339 (N_49339,N_46007,N_46193);
nand U49340 (N_49340,N_45002,N_46520);
nand U49341 (N_49341,N_46383,N_47173);
or U49342 (N_49342,N_47280,N_45087);
or U49343 (N_49343,N_47484,N_47307);
or U49344 (N_49344,N_45119,N_47206);
and U49345 (N_49345,N_45112,N_45297);
and U49346 (N_49346,N_47309,N_47368);
or U49347 (N_49347,N_45189,N_46435);
nor U49348 (N_49348,N_46238,N_45303);
nor U49349 (N_49349,N_45944,N_47412);
xnor U49350 (N_49350,N_45292,N_45035);
nor U49351 (N_49351,N_46214,N_47155);
or U49352 (N_49352,N_46794,N_45262);
or U49353 (N_49353,N_46891,N_47176);
or U49354 (N_49354,N_45214,N_46621);
and U49355 (N_49355,N_45081,N_47271);
xor U49356 (N_49356,N_45149,N_45480);
or U49357 (N_49357,N_46255,N_45686);
and U49358 (N_49358,N_45055,N_47301);
and U49359 (N_49359,N_47190,N_46532);
nor U49360 (N_49360,N_46393,N_47106);
nand U49361 (N_49361,N_46882,N_45694);
and U49362 (N_49362,N_45621,N_47145);
nand U49363 (N_49363,N_47463,N_47422);
or U49364 (N_49364,N_45510,N_45011);
nor U49365 (N_49365,N_45068,N_46243);
nand U49366 (N_49366,N_46778,N_45562);
xor U49367 (N_49367,N_45148,N_45165);
xnor U49368 (N_49368,N_47313,N_47486);
xnor U49369 (N_49369,N_45061,N_45855);
nand U49370 (N_49370,N_46165,N_45534);
xor U49371 (N_49371,N_45717,N_46069);
xor U49372 (N_49372,N_45398,N_46957);
and U49373 (N_49373,N_46239,N_46068);
or U49374 (N_49374,N_46966,N_45536);
nand U49375 (N_49375,N_46719,N_46827);
xor U49376 (N_49376,N_45371,N_46028);
or U49377 (N_49377,N_45731,N_45074);
and U49378 (N_49378,N_45469,N_45216);
or U49379 (N_49379,N_45438,N_46939);
or U49380 (N_49380,N_46896,N_46713);
xor U49381 (N_49381,N_46874,N_45889);
nor U49382 (N_49382,N_45524,N_46821);
or U49383 (N_49383,N_47456,N_45013);
nor U49384 (N_49384,N_46401,N_45448);
nand U49385 (N_49385,N_46593,N_47127);
xnor U49386 (N_49386,N_45125,N_46927);
nor U49387 (N_49387,N_46958,N_45355);
and U49388 (N_49388,N_46815,N_46123);
nand U49389 (N_49389,N_47084,N_47173);
xnor U49390 (N_49390,N_46203,N_45221);
or U49391 (N_49391,N_45980,N_45218);
xor U49392 (N_49392,N_46470,N_46209);
xnor U49393 (N_49393,N_45930,N_46155);
xor U49394 (N_49394,N_45524,N_45182);
and U49395 (N_49395,N_45254,N_46589);
nor U49396 (N_49396,N_46932,N_46891);
or U49397 (N_49397,N_45580,N_45094);
nor U49398 (N_49398,N_45430,N_46988);
nor U49399 (N_49399,N_45787,N_46140);
nor U49400 (N_49400,N_46033,N_46903);
and U49401 (N_49401,N_45549,N_46405);
nand U49402 (N_49402,N_46923,N_45221);
xor U49403 (N_49403,N_45791,N_46173);
nor U49404 (N_49404,N_46833,N_47105);
and U49405 (N_49405,N_45121,N_47070);
and U49406 (N_49406,N_47458,N_46050);
and U49407 (N_49407,N_46474,N_47309);
or U49408 (N_49408,N_47115,N_46862);
nand U49409 (N_49409,N_45742,N_46353);
and U49410 (N_49410,N_45092,N_46164);
or U49411 (N_49411,N_45059,N_46785);
xnor U49412 (N_49412,N_46800,N_45117);
or U49413 (N_49413,N_46371,N_47079);
and U49414 (N_49414,N_45376,N_45495);
and U49415 (N_49415,N_45369,N_46508);
nand U49416 (N_49416,N_45830,N_46143);
nand U49417 (N_49417,N_46644,N_45903);
nor U49418 (N_49418,N_46146,N_45901);
or U49419 (N_49419,N_46585,N_46030);
nand U49420 (N_49420,N_46075,N_45457);
and U49421 (N_49421,N_45151,N_46262);
or U49422 (N_49422,N_46012,N_45227);
xor U49423 (N_49423,N_45340,N_46779);
nand U49424 (N_49424,N_47161,N_46498);
or U49425 (N_49425,N_45100,N_46056);
nand U49426 (N_49426,N_47207,N_45508);
nand U49427 (N_49427,N_45097,N_45055);
nand U49428 (N_49428,N_46876,N_46101);
nor U49429 (N_49429,N_46219,N_46061);
xnor U49430 (N_49430,N_45728,N_46456);
xnor U49431 (N_49431,N_46504,N_47225);
and U49432 (N_49432,N_45437,N_45892);
nand U49433 (N_49433,N_46581,N_46733);
nand U49434 (N_49434,N_46291,N_45783);
nand U49435 (N_49435,N_46361,N_46994);
and U49436 (N_49436,N_45591,N_47273);
nor U49437 (N_49437,N_45806,N_46223);
xnor U49438 (N_49438,N_45754,N_45958);
and U49439 (N_49439,N_46151,N_46875);
and U49440 (N_49440,N_45424,N_46249);
nor U49441 (N_49441,N_45382,N_45281);
xnor U49442 (N_49442,N_47456,N_46016);
nand U49443 (N_49443,N_46393,N_45918);
and U49444 (N_49444,N_46117,N_45018);
nand U49445 (N_49445,N_45626,N_47024);
and U49446 (N_49446,N_45021,N_46200);
nor U49447 (N_49447,N_46950,N_46124);
nand U49448 (N_49448,N_45603,N_46023);
and U49449 (N_49449,N_45108,N_45151);
or U49450 (N_49450,N_45551,N_47385);
nand U49451 (N_49451,N_45593,N_46031);
nand U49452 (N_49452,N_46144,N_45951);
and U49453 (N_49453,N_46874,N_45091);
xor U49454 (N_49454,N_45921,N_47416);
or U49455 (N_49455,N_45640,N_47410);
or U49456 (N_49456,N_46275,N_45962);
nand U49457 (N_49457,N_46073,N_45839);
and U49458 (N_49458,N_45702,N_46336);
nand U49459 (N_49459,N_46227,N_45632);
nor U49460 (N_49460,N_45864,N_46171);
or U49461 (N_49461,N_46341,N_46714);
and U49462 (N_49462,N_45828,N_46277);
xnor U49463 (N_49463,N_45739,N_47233);
or U49464 (N_49464,N_46306,N_46300);
and U49465 (N_49465,N_46592,N_46096);
nor U49466 (N_49466,N_47123,N_45265);
nor U49467 (N_49467,N_45498,N_46661);
xor U49468 (N_49468,N_46636,N_45576);
nand U49469 (N_49469,N_45857,N_47033);
and U49470 (N_49470,N_47044,N_45652);
or U49471 (N_49471,N_46096,N_46684);
and U49472 (N_49472,N_47498,N_47345);
or U49473 (N_49473,N_46995,N_46055);
xnor U49474 (N_49474,N_46959,N_46821);
nand U49475 (N_49475,N_45758,N_45540);
nand U49476 (N_49476,N_45750,N_45849);
and U49477 (N_49477,N_46151,N_45079);
xnor U49478 (N_49478,N_45358,N_47351);
or U49479 (N_49479,N_45542,N_46388);
or U49480 (N_49480,N_46661,N_47055);
nand U49481 (N_49481,N_47185,N_46029);
nor U49482 (N_49482,N_46412,N_46512);
or U49483 (N_49483,N_45577,N_46813);
nor U49484 (N_49484,N_47400,N_45529);
or U49485 (N_49485,N_45519,N_46987);
xor U49486 (N_49486,N_46013,N_46000);
xor U49487 (N_49487,N_47493,N_47345);
or U49488 (N_49488,N_45220,N_46054);
nor U49489 (N_49489,N_47422,N_47018);
xor U49490 (N_49490,N_47336,N_45660);
nand U49491 (N_49491,N_46072,N_45078);
or U49492 (N_49492,N_45739,N_45031);
nand U49493 (N_49493,N_47023,N_47031);
or U49494 (N_49494,N_45750,N_47138);
nor U49495 (N_49495,N_47457,N_45292);
nor U49496 (N_49496,N_46420,N_45203);
and U49497 (N_49497,N_45209,N_47373);
nor U49498 (N_49498,N_46694,N_46525);
nand U49499 (N_49499,N_46780,N_46628);
and U49500 (N_49500,N_45890,N_46604);
or U49501 (N_49501,N_47256,N_45827);
nor U49502 (N_49502,N_45375,N_45886);
xor U49503 (N_49503,N_45340,N_46976);
xor U49504 (N_49504,N_45555,N_45696);
and U49505 (N_49505,N_45562,N_45875);
xor U49506 (N_49506,N_46768,N_46003);
and U49507 (N_49507,N_45385,N_47231);
or U49508 (N_49508,N_47475,N_46372);
xor U49509 (N_49509,N_46936,N_46466);
or U49510 (N_49510,N_45402,N_46316);
nand U49511 (N_49511,N_46559,N_46889);
xor U49512 (N_49512,N_46312,N_45385);
nand U49513 (N_49513,N_46401,N_45670);
or U49514 (N_49514,N_46888,N_46284);
and U49515 (N_49515,N_47273,N_46014);
and U49516 (N_49516,N_46209,N_46024);
and U49517 (N_49517,N_47414,N_46575);
or U49518 (N_49518,N_45881,N_46113);
nand U49519 (N_49519,N_45201,N_45433);
xnor U49520 (N_49520,N_46135,N_47243);
xnor U49521 (N_49521,N_46951,N_46650);
and U49522 (N_49522,N_47188,N_45020);
nand U49523 (N_49523,N_45518,N_46820);
and U49524 (N_49524,N_47494,N_45343);
and U49525 (N_49525,N_45552,N_47188);
nor U49526 (N_49526,N_45453,N_45173);
or U49527 (N_49527,N_46814,N_45602);
and U49528 (N_49528,N_46905,N_45439);
nand U49529 (N_49529,N_47494,N_47004);
nand U49530 (N_49530,N_45234,N_47387);
and U49531 (N_49531,N_46732,N_46783);
nor U49532 (N_49532,N_45718,N_46552);
nand U49533 (N_49533,N_45774,N_47139);
or U49534 (N_49534,N_46262,N_46986);
nor U49535 (N_49535,N_46509,N_45873);
nor U49536 (N_49536,N_46525,N_46469);
xnor U49537 (N_49537,N_45869,N_45961);
nor U49538 (N_49538,N_45586,N_47085);
or U49539 (N_49539,N_46960,N_46256);
nor U49540 (N_49540,N_46784,N_47304);
or U49541 (N_49541,N_47118,N_46158);
and U49542 (N_49542,N_47148,N_45529);
or U49543 (N_49543,N_47333,N_45674);
nor U49544 (N_49544,N_45391,N_47308);
nand U49545 (N_49545,N_45602,N_46399);
nand U49546 (N_49546,N_45754,N_46160);
nor U49547 (N_49547,N_45061,N_46456);
or U49548 (N_49548,N_47483,N_45743);
nor U49549 (N_49549,N_45579,N_46157);
or U49550 (N_49550,N_46410,N_45862);
nor U49551 (N_49551,N_45904,N_47214);
nor U49552 (N_49552,N_46081,N_45907);
xor U49553 (N_49553,N_45970,N_47421);
and U49554 (N_49554,N_46544,N_46657);
xor U49555 (N_49555,N_46455,N_47083);
nand U49556 (N_49556,N_46706,N_46786);
and U49557 (N_49557,N_47033,N_46550);
and U49558 (N_49558,N_47352,N_45328);
or U49559 (N_49559,N_45006,N_47217);
nor U49560 (N_49560,N_47309,N_46150);
nand U49561 (N_49561,N_46723,N_45159);
nor U49562 (N_49562,N_46228,N_46735);
xnor U49563 (N_49563,N_46170,N_45705);
nor U49564 (N_49564,N_47042,N_47376);
and U49565 (N_49565,N_45914,N_45358);
and U49566 (N_49566,N_45241,N_45190);
nor U49567 (N_49567,N_47433,N_47205);
nand U49568 (N_49568,N_45884,N_46991);
xnor U49569 (N_49569,N_45294,N_46264);
or U49570 (N_49570,N_46125,N_45270);
and U49571 (N_49571,N_45877,N_46300);
nor U49572 (N_49572,N_46874,N_47170);
nand U49573 (N_49573,N_47324,N_45501);
nor U49574 (N_49574,N_46848,N_46188);
or U49575 (N_49575,N_45580,N_47395);
nor U49576 (N_49576,N_45891,N_46743);
xor U49577 (N_49577,N_46771,N_45941);
xor U49578 (N_49578,N_46054,N_46578);
and U49579 (N_49579,N_45347,N_45248);
or U49580 (N_49580,N_45898,N_45092);
nor U49581 (N_49581,N_45078,N_47228);
or U49582 (N_49582,N_46037,N_46409);
nor U49583 (N_49583,N_46062,N_47459);
xnor U49584 (N_49584,N_46944,N_46559);
and U49585 (N_49585,N_45268,N_45160);
or U49586 (N_49586,N_46033,N_45091);
and U49587 (N_49587,N_45534,N_47166);
xor U49588 (N_49588,N_46122,N_45737);
nand U49589 (N_49589,N_46921,N_45022);
xnor U49590 (N_49590,N_47298,N_45869);
xnor U49591 (N_49591,N_46040,N_46385);
nand U49592 (N_49592,N_45685,N_47028);
and U49593 (N_49593,N_47011,N_46581);
and U49594 (N_49594,N_46706,N_45158);
xnor U49595 (N_49595,N_46837,N_45790);
nor U49596 (N_49596,N_46952,N_46360);
xnor U49597 (N_49597,N_46741,N_46239);
or U49598 (N_49598,N_46030,N_46101);
nor U49599 (N_49599,N_45769,N_46238);
and U49600 (N_49600,N_45659,N_45514);
or U49601 (N_49601,N_47095,N_46463);
and U49602 (N_49602,N_46043,N_46060);
nor U49603 (N_49603,N_45129,N_47143);
nor U49604 (N_49604,N_47015,N_45905);
xnor U49605 (N_49605,N_46777,N_46544);
and U49606 (N_49606,N_46394,N_46389);
or U49607 (N_49607,N_45491,N_47001);
xnor U49608 (N_49608,N_47200,N_46775);
or U49609 (N_49609,N_46320,N_45176);
nor U49610 (N_49610,N_47450,N_47250);
nor U49611 (N_49611,N_46537,N_47005);
xor U49612 (N_49612,N_46463,N_46957);
xnor U49613 (N_49613,N_45232,N_46235);
nor U49614 (N_49614,N_45232,N_45953);
nor U49615 (N_49615,N_46996,N_45539);
and U49616 (N_49616,N_46386,N_45588);
or U49617 (N_49617,N_47224,N_45363);
nand U49618 (N_49618,N_45596,N_45497);
or U49619 (N_49619,N_45086,N_45406);
or U49620 (N_49620,N_45099,N_45884);
nand U49621 (N_49621,N_47206,N_45266);
or U49622 (N_49622,N_46291,N_46503);
and U49623 (N_49623,N_45767,N_46372);
xnor U49624 (N_49624,N_47105,N_45260);
nand U49625 (N_49625,N_47263,N_46262);
nor U49626 (N_49626,N_46177,N_46178);
xor U49627 (N_49627,N_46732,N_47290);
nor U49628 (N_49628,N_45148,N_47350);
or U49629 (N_49629,N_47196,N_47095);
xnor U49630 (N_49630,N_45339,N_46613);
nor U49631 (N_49631,N_45246,N_45873);
nor U49632 (N_49632,N_46938,N_46145);
and U49633 (N_49633,N_47233,N_46560);
xnor U49634 (N_49634,N_45685,N_46834);
nand U49635 (N_49635,N_46922,N_47283);
nand U49636 (N_49636,N_45667,N_46433);
or U49637 (N_49637,N_46579,N_46053);
xnor U49638 (N_49638,N_45447,N_47419);
xor U49639 (N_49639,N_45445,N_46897);
and U49640 (N_49640,N_47322,N_45385);
and U49641 (N_49641,N_46710,N_47165);
nor U49642 (N_49642,N_45405,N_47159);
nand U49643 (N_49643,N_45050,N_46010);
or U49644 (N_49644,N_47039,N_45905);
nor U49645 (N_49645,N_45418,N_46839);
or U49646 (N_49646,N_46852,N_46948);
nand U49647 (N_49647,N_45560,N_46819);
nand U49648 (N_49648,N_47107,N_45257);
and U49649 (N_49649,N_47168,N_45846);
nand U49650 (N_49650,N_45746,N_46165);
or U49651 (N_49651,N_46687,N_45791);
or U49652 (N_49652,N_46690,N_45755);
and U49653 (N_49653,N_45751,N_46692);
nor U49654 (N_49654,N_45563,N_46258);
and U49655 (N_49655,N_46033,N_46979);
nand U49656 (N_49656,N_47236,N_45248);
or U49657 (N_49657,N_45328,N_45796);
xnor U49658 (N_49658,N_45233,N_47135);
or U49659 (N_49659,N_45726,N_46995);
nor U49660 (N_49660,N_45429,N_45688);
or U49661 (N_49661,N_45791,N_47176);
and U49662 (N_49662,N_46687,N_45715);
nor U49663 (N_49663,N_45992,N_45694);
xor U49664 (N_49664,N_47154,N_46009);
nor U49665 (N_49665,N_45830,N_47226);
nand U49666 (N_49666,N_46022,N_45706);
nor U49667 (N_49667,N_47324,N_47371);
and U49668 (N_49668,N_45640,N_46687);
xor U49669 (N_49669,N_45199,N_46547);
xnor U49670 (N_49670,N_46548,N_47252);
nor U49671 (N_49671,N_46149,N_46320);
and U49672 (N_49672,N_46949,N_45901);
xor U49673 (N_49673,N_46122,N_46904);
or U49674 (N_49674,N_46146,N_45053);
or U49675 (N_49675,N_45085,N_46497);
and U49676 (N_49676,N_46094,N_46222);
xor U49677 (N_49677,N_45074,N_47123);
nor U49678 (N_49678,N_46590,N_46906);
xnor U49679 (N_49679,N_45089,N_46712);
nand U49680 (N_49680,N_46722,N_45394);
xnor U49681 (N_49681,N_46464,N_46471);
xnor U49682 (N_49682,N_47448,N_47168);
or U49683 (N_49683,N_46447,N_47164);
nand U49684 (N_49684,N_47340,N_45977);
and U49685 (N_49685,N_46709,N_45052);
and U49686 (N_49686,N_45240,N_45689);
nand U49687 (N_49687,N_46545,N_46704);
and U49688 (N_49688,N_47086,N_46575);
nand U49689 (N_49689,N_47357,N_47472);
nand U49690 (N_49690,N_46023,N_45036);
xnor U49691 (N_49691,N_47342,N_46795);
xnor U49692 (N_49692,N_45171,N_46771);
or U49693 (N_49693,N_46125,N_46289);
xnor U49694 (N_49694,N_46105,N_46888);
or U49695 (N_49695,N_45844,N_45264);
xor U49696 (N_49696,N_46407,N_46455);
and U49697 (N_49697,N_46796,N_47169);
or U49698 (N_49698,N_47165,N_45290);
or U49699 (N_49699,N_47489,N_45527);
and U49700 (N_49700,N_47188,N_45787);
xnor U49701 (N_49701,N_46728,N_45198);
nor U49702 (N_49702,N_46683,N_45020);
xor U49703 (N_49703,N_46241,N_46139);
nor U49704 (N_49704,N_46123,N_46076);
xor U49705 (N_49705,N_45374,N_46453);
xnor U49706 (N_49706,N_47141,N_46462);
xnor U49707 (N_49707,N_45260,N_47004);
or U49708 (N_49708,N_45957,N_45378);
xnor U49709 (N_49709,N_46980,N_46784);
xnor U49710 (N_49710,N_45527,N_45444);
and U49711 (N_49711,N_46597,N_46551);
nand U49712 (N_49712,N_45355,N_45541);
nor U49713 (N_49713,N_46872,N_45291);
and U49714 (N_49714,N_46977,N_46380);
or U49715 (N_49715,N_46313,N_46432);
and U49716 (N_49716,N_45376,N_46269);
nand U49717 (N_49717,N_45992,N_45971);
and U49718 (N_49718,N_46238,N_47310);
and U49719 (N_49719,N_46564,N_47225);
nor U49720 (N_49720,N_46980,N_45381);
or U49721 (N_49721,N_47358,N_46809);
or U49722 (N_49722,N_47043,N_47269);
nor U49723 (N_49723,N_47024,N_46951);
xnor U49724 (N_49724,N_46147,N_45461);
nor U49725 (N_49725,N_46497,N_46244);
or U49726 (N_49726,N_45380,N_45109);
and U49727 (N_49727,N_47133,N_45527);
and U49728 (N_49728,N_46103,N_46167);
and U49729 (N_49729,N_45375,N_46952);
xor U49730 (N_49730,N_46009,N_45394);
and U49731 (N_49731,N_47219,N_46629);
nand U49732 (N_49732,N_45704,N_46783);
nor U49733 (N_49733,N_45071,N_45814);
xor U49734 (N_49734,N_45473,N_47255);
xor U49735 (N_49735,N_45198,N_47309);
nand U49736 (N_49736,N_45747,N_47488);
xnor U49737 (N_49737,N_46947,N_46317);
and U49738 (N_49738,N_46732,N_47368);
or U49739 (N_49739,N_45825,N_45077);
and U49740 (N_49740,N_46649,N_47167);
and U49741 (N_49741,N_45620,N_46546);
xor U49742 (N_49742,N_45768,N_45834);
nand U49743 (N_49743,N_46071,N_46832);
xnor U49744 (N_49744,N_46380,N_45158);
nand U49745 (N_49745,N_46704,N_46653);
and U49746 (N_49746,N_46430,N_45441);
xor U49747 (N_49747,N_45177,N_47391);
nand U49748 (N_49748,N_47324,N_46118);
or U49749 (N_49749,N_46165,N_46426);
nand U49750 (N_49750,N_46923,N_46484);
nor U49751 (N_49751,N_45600,N_46562);
or U49752 (N_49752,N_47375,N_46543);
or U49753 (N_49753,N_45513,N_46216);
xnor U49754 (N_49754,N_46691,N_46325);
xor U49755 (N_49755,N_45597,N_45233);
nand U49756 (N_49756,N_47239,N_47251);
nand U49757 (N_49757,N_45565,N_46690);
and U49758 (N_49758,N_45019,N_45981);
nand U49759 (N_49759,N_46987,N_47447);
and U49760 (N_49760,N_47415,N_47384);
xnor U49761 (N_49761,N_45493,N_45390);
xor U49762 (N_49762,N_45984,N_47023);
nand U49763 (N_49763,N_47176,N_46430);
nor U49764 (N_49764,N_47047,N_45920);
nor U49765 (N_49765,N_46927,N_45504);
xnor U49766 (N_49766,N_46909,N_45399);
nor U49767 (N_49767,N_46253,N_45661);
nand U49768 (N_49768,N_45306,N_46959);
xnor U49769 (N_49769,N_45961,N_45300);
nand U49770 (N_49770,N_46660,N_47281);
nand U49771 (N_49771,N_46222,N_46361);
nand U49772 (N_49772,N_45738,N_45031);
and U49773 (N_49773,N_46831,N_45407);
and U49774 (N_49774,N_47304,N_45621);
or U49775 (N_49775,N_46563,N_46640);
or U49776 (N_49776,N_46003,N_46928);
xnor U49777 (N_49777,N_45199,N_45200);
or U49778 (N_49778,N_46921,N_46369);
and U49779 (N_49779,N_45849,N_45393);
or U49780 (N_49780,N_45486,N_46387);
nand U49781 (N_49781,N_46918,N_45845);
or U49782 (N_49782,N_46001,N_46399);
nor U49783 (N_49783,N_46065,N_46323);
nand U49784 (N_49784,N_47341,N_45095);
and U49785 (N_49785,N_46101,N_46920);
or U49786 (N_49786,N_46520,N_45851);
nor U49787 (N_49787,N_45439,N_46194);
xnor U49788 (N_49788,N_47019,N_47491);
nor U49789 (N_49789,N_45786,N_45219);
nor U49790 (N_49790,N_46568,N_46892);
nand U49791 (N_49791,N_46187,N_46739);
nor U49792 (N_49792,N_47065,N_46406);
nor U49793 (N_49793,N_46147,N_47183);
and U49794 (N_49794,N_46466,N_47166);
or U49795 (N_49795,N_46334,N_45494);
nand U49796 (N_49796,N_46390,N_45895);
xnor U49797 (N_49797,N_47318,N_45544);
nor U49798 (N_49798,N_45088,N_45533);
or U49799 (N_49799,N_45919,N_45745);
or U49800 (N_49800,N_47171,N_45864);
or U49801 (N_49801,N_46287,N_45182);
nand U49802 (N_49802,N_46597,N_46862);
nor U49803 (N_49803,N_47385,N_47306);
and U49804 (N_49804,N_45659,N_47102);
nor U49805 (N_49805,N_47482,N_46753);
nor U49806 (N_49806,N_45626,N_47359);
xnor U49807 (N_49807,N_46377,N_46739);
and U49808 (N_49808,N_45522,N_45776);
nor U49809 (N_49809,N_45734,N_45059);
nor U49810 (N_49810,N_45996,N_46065);
xor U49811 (N_49811,N_47156,N_46354);
nand U49812 (N_49812,N_45974,N_47059);
or U49813 (N_49813,N_45983,N_47228);
nor U49814 (N_49814,N_46831,N_47301);
nand U49815 (N_49815,N_47282,N_45475);
xor U49816 (N_49816,N_46707,N_45990);
xor U49817 (N_49817,N_47455,N_45574);
nand U49818 (N_49818,N_46030,N_45344);
nor U49819 (N_49819,N_46355,N_47496);
and U49820 (N_49820,N_46890,N_45620);
nor U49821 (N_49821,N_46368,N_46611);
xor U49822 (N_49822,N_46868,N_45836);
nor U49823 (N_49823,N_45174,N_45587);
nor U49824 (N_49824,N_45509,N_46615);
nor U49825 (N_49825,N_45317,N_46507);
nand U49826 (N_49826,N_47273,N_45368);
or U49827 (N_49827,N_46930,N_46079);
xnor U49828 (N_49828,N_46727,N_45929);
xnor U49829 (N_49829,N_47169,N_46047);
xnor U49830 (N_49830,N_46950,N_46367);
nand U49831 (N_49831,N_46767,N_45615);
nor U49832 (N_49832,N_45354,N_47317);
nor U49833 (N_49833,N_46618,N_46899);
and U49834 (N_49834,N_47293,N_47139);
xnor U49835 (N_49835,N_45786,N_46013);
nor U49836 (N_49836,N_46177,N_45921);
xnor U49837 (N_49837,N_45109,N_45306);
xnor U49838 (N_49838,N_47099,N_45549);
and U49839 (N_49839,N_47234,N_45062);
and U49840 (N_49840,N_46965,N_45849);
nor U49841 (N_49841,N_47138,N_46063);
and U49842 (N_49842,N_45820,N_46920);
xnor U49843 (N_49843,N_45453,N_46665);
nand U49844 (N_49844,N_45402,N_47399);
or U49845 (N_49845,N_46612,N_47318);
nand U49846 (N_49846,N_46618,N_47450);
nand U49847 (N_49847,N_45257,N_45502);
xnor U49848 (N_49848,N_46702,N_45176);
xor U49849 (N_49849,N_45667,N_46427);
and U49850 (N_49850,N_47215,N_47218);
or U49851 (N_49851,N_45063,N_46813);
xnor U49852 (N_49852,N_45677,N_45519);
xnor U49853 (N_49853,N_47418,N_47119);
or U49854 (N_49854,N_45677,N_46342);
and U49855 (N_49855,N_46524,N_45489);
nor U49856 (N_49856,N_45003,N_46696);
nand U49857 (N_49857,N_47403,N_46099);
xor U49858 (N_49858,N_46524,N_46702);
nand U49859 (N_49859,N_45895,N_45965);
nand U49860 (N_49860,N_46720,N_46790);
xnor U49861 (N_49861,N_47200,N_45140);
and U49862 (N_49862,N_45840,N_46671);
or U49863 (N_49863,N_47155,N_46138);
xor U49864 (N_49864,N_45040,N_46963);
or U49865 (N_49865,N_45047,N_46278);
nand U49866 (N_49866,N_46610,N_46117);
nor U49867 (N_49867,N_47285,N_46919);
nand U49868 (N_49868,N_47311,N_45665);
xnor U49869 (N_49869,N_45366,N_46756);
nand U49870 (N_49870,N_46744,N_47238);
nand U49871 (N_49871,N_45409,N_46705);
xnor U49872 (N_49872,N_46502,N_47216);
nand U49873 (N_49873,N_45738,N_45277);
nor U49874 (N_49874,N_47414,N_47184);
or U49875 (N_49875,N_45273,N_47308);
xor U49876 (N_49876,N_46514,N_46606);
or U49877 (N_49877,N_47231,N_45882);
nor U49878 (N_49878,N_47037,N_45246);
nor U49879 (N_49879,N_46181,N_46688);
nor U49880 (N_49880,N_46344,N_45158);
xor U49881 (N_49881,N_45963,N_46737);
nand U49882 (N_49882,N_47407,N_45733);
or U49883 (N_49883,N_45400,N_46354);
and U49884 (N_49884,N_47484,N_46317);
nor U49885 (N_49885,N_46621,N_45654);
nand U49886 (N_49886,N_47388,N_46660);
nand U49887 (N_49887,N_46012,N_46944);
xnor U49888 (N_49888,N_45441,N_45605);
or U49889 (N_49889,N_46844,N_45405);
nor U49890 (N_49890,N_46522,N_47008);
and U49891 (N_49891,N_47292,N_46979);
and U49892 (N_49892,N_45426,N_47187);
or U49893 (N_49893,N_45395,N_45736);
and U49894 (N_49894,N_45073,N_46542);
or U49895 (N_49895,N_47272,N_47082);
or U49896 (N_49896,N_45060,N_46429);
or U49897 (N_49897,N_46850,N_45319);
and U49898 (N_49898,N_45036,N_46448);
nand U49899 (N_49899,N_47308,N_46554);
and U49900 (N_49900,N_45792,N_47402);
nand U49901 (N_49901,N_45751,N_45173);
xnor U49902 (N_49902,N_47168,N_45916);
nand U49903 (N_49903,N_47343,N_46507);
nand U49904 (N_49904,N_45160,N_45934);
xnor U49905 (N_49905,N_47093,N_46530);
xor U49906 (N_49906,N_46520,N_47172);
xor U49907 (N_49907,N_45121,N_46214);
and U49908 (N_49908,N_45703,N_45264);
and U49909 (N_49909,N_46585,N_46355);
xnor U49910 (N_49910,N_45869,N_45855);
and U49911 (N_49911,N_46749,N_45171);
xnor U49912 (N_49912,N_46752,N_46973);
nor U49913 (N_49913,N_45082,N_46284);
nand U49914 (N_49914,N_46096,N_46862);
nor U49915 (N_49915,N_45324,N_47127);
xnor U49916 (N_49916,N_47269,N_46867);
or U49917 (N_49917,N_45557,N_45877);
or U49918 (N_49918,N_45429,N_46724);
nand U49919 (N_49919,N_47126,N_46893);
nor U49920 (N_49920,N_45391,N_47017);
xor U49921 (N_49921,N_45741,N_45876);
or U49922 (N_49922,N_45196,N_46204);
xor U49923 (N_49923,N_46819,N_46381);
nor U49924 (N_49924,N_45561,N_46477);
and U49925 (N_49925,N_46203,N_47487);
or U49926 (N_49926,N_47481,N_46242);
nor U49927 (N_49927,N_47044,N_47295);
nand U49928 (N_49928,N_45949,N_47163);
and U49929 (N_49929,N_47290,N_47021);
and U49930 (N_49930,N_47471,N_46266);
and U49931 (N_49931,N_47419,N_47114);
nor U49932 (N_49932,N_46123,N_46087);
or U49933 (N_49933,N_45909,N_47471);
nand U49934 (N_49934,N_45125,N_45356);
or U49935 (N_49935,N_45051,N_45965);
and U49936 (N_49936,N_45779,N_46557);
nand U49937 (N_49937,N_47326,N_46634);
xnor U49938 (N_49938,N_46150,N_47134);
and U49939 (N_49939,N_46184,N_45439);
xnor U49940 (N_49940,N_46337,N_46285);
nand U49941 (N_49941,N_45475,N_46864);
xnor U49942 (N_49942,N_46416,N_45544);
or U49943 (N_49943,N_45173,N_45010);
nor U49944 (N_49944,N_45429,N_46135);
and U49945 (N_49945,N_46684,N_46278);
nand U49946 (N_49946,N_45325,N_46117);
nand U49947 (N_49947,N_45520,N_46389);
nand U49948 (N_49948,N_45474,N_46105);
or U49949 (N_49949,N_46686,N_45908);
nand U49950 (N_49950,N_45564,N_47069);
or U49951 (N_49951,N_46524,N_46803);
or U49952 (N_49952,N_45633,N_45797);
or U49953 (N_49953,N_45839,N_46218);
and U49954 (N_49954,N_46765,N_45632);
xnor U49955 (N_49955,N_47378,N_45008);
and U49956 (N_49956,N_47388,N_46555);
or U49957 (N_49957,N_46429,N_45071);
xor U49958 (N_49958,N_47240,N_45002);
nor U49959 (N_49959,N_45681,N_46013);
nand U49960 (N_49960,N_47102,N_46980);
or U49961 (N_49961,N_45306,N_46242);
nor U49962 (N_49962,N_47254,N_45789);
nand U49963 (N_49963,N_45122,N_46594);
or U49964 (N_49964,N_47281,N_45248);
xor U49965 (N_49965,N_46365,N_45788);
xnor U49966 (N_49966,N_45094,N_47318);
nor U49967 (N_49967,N_46845,N_45241);
nor U49968 (N_49968,N_45434,N_45894);
nand U49969 (N_49969,N_45848,N_46830);
xor U49970 (N_49970,N_45877,N_45886);
xnor U49971 (N_49971,N_47480,N_46464);
and U49972 (N_49972,N_47248,N_46057);
nand U49973 (N_49973,N_45028,N_45706);
and U49974 (N_49974,N_46882,N_45007);
xnor U49975 (N_49975,N_47249,N_46225);
and U49976 (N_49976,N_46231,N_47424);
or U49977 (N_49977,N_47266,N_46105);
or U49978 (N_49978,N_46395,N_47301);
xor U49979 (N_49979,N_46356,N_45038);
nor U49980 (N_49980,N_45949,N_46479);
nor U49981 (N_49981,N_46299,N_47326);
or U49982 (N_49982,N_45637,N_47221);
and U49983 (N_49983,N_45254,N_45435);
nand U49984 (N_49984,N_46639,N_46563);
nor U49985 (N_49985,N_46481,N_47332);
nand U49986 (N_49986,N_46865,N_47408);
nor U49987 (N_49987,N_46644,N_45526);
xor U49988 (N_49988,N_46858,N_46580);
nand U49989 (N_49989,N_45933,N_45690);
and U49990 (N_49990,N_46329,N_46771);
nand U49991 (N_49991,N_47240,N_47371);
xor U49992 (N_49992,N_46586,N_45729);
nand U49993 (N_49993,N_46663,N_46095);
and U49994 (N_49994,N_47299,N_45591);
and U49995 (N_49995,N_47009,N_46082);
xor U49996 (N_49996,N_46487,N_47127);
and U49997 (N_49997,N_46843,N_46656);
nor U49998 (N_49998,N_45969,N_47225);
or U49999 (N_49999,N_46556,N_46254);
or UO_0 (O_0,N_49658,N_47551);
xor UO_1 (O_1,N_49590,N_47603);
xor UO_2 (O_2,N_47627,N_49412);
nand UO_3 (O_3,N_48485,N_49870);
nand UO_4 (O_4,N_49557,N_48435);
nand UO_5 (O_5,N_49484,N_47983);
and UO_6 (O_6,N_49199,N_47820);
or UO_7 (O_7,N_49542,N_49717);
xor UO_8 (O_8,N_48202,N_48700);
xor UO_9 (O_9,N_47947,N_49513);
nor UO_10 (O_10,N_49926,N_47893);
nor UO_11 (O_11,N_47806,N_48938);
xor UO_12 (O_12,N_49980,N_48678);
nand UO_13 (O_13,N_49462,N_49411);
xor UO_14 (O_14,N_47920,N_49264);
and UO_15 (O_15,N_47928,N_49425);
nand UO_16 (O_16,N_48441,N_48904);
xnor UO_17 (O_17,N_49163,N_49794);
and UO_18 (O_18,N_47952,N_49402);
or UO_19 (O_19,N_48980,N_49197);
nor UO_20 (O_20,N_47989,N_48706);
nor UO_21 (O_21,N_47687,N_49622);
and UO_22 (O_22,N_48519,N_48614);
nor UO_23 (O_23,N_47673,N_49452);
nor UO_24 (O_24,N_49375,N_49167);
nand UO_25 (O_25,N_49181,N_47718);
and UO_26 (O_26,N_47981,N_48983);
nand UO_27 (O_27,N_48262,N_49093);
and UO_28 (O_28,N_49787,N_49827);
nor UO_29 (O_29,N_47871,N_47748);
nand UO_30 (O_30,N_48746,N_47508);
nor UO_31 (O_31,N_49797,N_49781);
and UO_32 (O_32,N_48307,N_48793);
nand UO_33 (O_33,N_49269,N_49888);
or UO_34 (O_34,N_49783,N_47783);
nor UO_35 (O_35,N_49683,N_49474);
and UO_36 (O_36,N_48826,N_49022);
xor UO_37 (O_37,N_48354,N_48752);
nor UO_38 (O_38,N_49766,N_47804);
nor UO_39 (O_39,N_48601,N_49242);
nor UO_40 (O_40,N_49747,N_47509);
xor UO_41 (O_41,N_49865,N_47714);
or UO_42 (O_42,N_49603,N_48003);
and UO_43 (O_43,N_47801,N_48438);
nor UO_44 (O_44,N_48268,N_48596);
or UO_45 (O_45,N_49171,N_49250);
xor UO_46 (O_46,N_49421,N_48658);
nand UO_47 (O_47,N_47629,N_49225);
nand UO_48 (O_48,N_49207,N_47858);
nor UO_49 (O_49,N_49089,N_49640);
xor UO_50 (O_50,N_49738,N_47639);
nand UO_51 (O_51,N_48227,N_48177);
nor UO_52 (O_52,N_47847,N_48504);
nand UO_53 (O_53,N_48871,N_49148);
nand UO_54 (O_54,N_48429,N_48317);
or UO_55 (O_55,N_47805,N_47516);
and UO_56 (O_56,N_48932,N_49252);
or UO_57 (O_57,N_47631,N_48180);
nor UO_58 (O_58,N_49443,N_48587);
xor UO_59 (O_59,N_49078,N_48577);
nand UO_60 (O_60,N_48673,N_48327);
and UO_61 (O_61,N_49313,N_48011);
and UO_62 (O_62,N_49393,N_49613);
or UO_63 (O_63,N_49025,N_48323);
and UO_64 (O_64,N_49731,N_49260);
xnor UO_65 (O_65,N_49862,N_48168);
or UO_66 (O_66,N_48946,N_49602);
and UO_67 (O_67,N_49869,N_47752);
nand UO_68 (O_68,N_48281,N_49232);
nand UO_69 (O_69,N_49380,N_49251);
or UO_70 (O_70,N_48960,N_49431);
or UO_71 (O_71,N_48810,N_49086);
xor UO_72 (O_72,N_47924,N_47534);
nor UO_73 (O_73,N_47915,N_49974);
nor UO_74 (O_74,N_48664,N_48620);
or UO_75 (O_75,N_48141,N_48459);
and UO_76 (O_76,N_47867,N_49301);
nand UO_77 (O_77,N_48757,N_49663);
nand UO_78 (O_78,N_49978,N_48543);
and UO_79 (O_79,N_49779,N_48784);
and UO_80 (O_80,N_47761,N_49570);
and UO_81 (O_81,N_47654,N_48032);
or UO_82 (O_82,N_49258,N_49071);
nand UO_83 (O_83,N_48583,N_48381);
and UO_84 (O_84,N_47930,N_49600);
nor UO_85 (O_85,N_49987,N_47927);
nand UO_86 (O_86,N_47731,N_48563);
nor UO_87 (O_87,N_49107,N_49111);
and UO_88 (O_88,N_48874,N_49520);
nand UO_89 (O_89,N_48047,N_48454);
nor UO_90 (O_90,N_49689,N_48539);
nand UO_91 (O_91,N_48056,N_47993);
xnor UO_92 (O_92,N_47555,N_47572);
or UO_93 (O_93,N_49955,N_48249);
and UO_94 (O_94,N_49563,N_48860);
and UO_95 (O_95,N_47765,N_48363);
nor UO_96 (O_96,N_49596,N_48802);
nor UO_97 (O_97,N_48285,N_48128);
xor UO_98 (O_98,N_49471,N_49399);
nor UO_99 (O_99,N_49147,N_49876);
nand UO_100 (O_100,N_49076,N_48819);
nor UO_101 (O_101,N_47736,N_49075);
nor UO_102 (O_102,N_48853,N_49810);
nor UO_103 (O_103,N_48146,N_48179);
xnor UO_104 (O_104,N_48240,N_49247);
xor UO_105 (O_105,N_48926,N_48712);
or UO_106 (O_106,N_49254,N_47630);
or UO_107 (O_107,N_48625,N_49579);
nor UO_108 (O_108,N_47942,N_48621);
or UO_109 (O_109,N_48149,N_47710);
and UO_110 (O_110,N_47987,N_47901);
and UO_111 (O_111,N_49261,N_47666);
and UO_112 (O_112,N_48592,N_49378);
xor UO_113 (O_113,N_47579,N_47699);
and UO_114 (O_114,N_49940,N_49604);
xor UO_115 (O_115,N_47829,N_48896);
and UO_116 (O_116,N_47708,N_48344);
and UO_117 (O_117,N_48713,N_48533);
nand UO_118 (O_118,N_48033,N_49326);
and UO_119 (O_119,N_47590,N_47956);
and UO_120 (O_120,N_47964,N_49495);
and UO_121 (O_121,N_49480,N_48201);
nor UO_122 (O_122,N_48869,N_49339);
and UO_123 (O_123,N_47824,N_47570);
xnor UO_124 (O_124,N_48366,N_49863);
nor UO_125 (O_125,N_49857,N_48430);
nor UO_126 (O_126,N_49959,N_49358);
and UO_127 (O_127,N_48081,N_48490);
xor UO_128 (O_128,N_49201,N_48844);
nor UO_129 (O_129,N_47713,N_47543);
nor UO_130 (O_130,N_47507,N_47971);
xor UO_131 (O_131,N_49165,N_48476);
and UO_132 (O_132,N_48412,N_48740);
xor UO_133 (O_133,N_48742,N_48073);
or UO_134 (O_134,N_47665,N_48699);
xor UO_135 (O_135,N_49861,N_48024);
nor UO_136 (O_136,N_49517,N_49759);
xor UO_137 (O_137,N_48199,N_47916);
nor UO_138 (O_138,N_49648,N_48575);
and UO_139 (O_139,N_49394,N_49638);
and UO_140 (O_140,N_47746,N_49131);
and UO_141 (O_141,N_49238,N_49776);
xnor UO_142 (O_142,N_48609,N_49934);
nand UO_143 (O_143,N_48615,N_48104);
nand UO_144 (O_144,N_48385,N_49208);
or UO_145 (O_145,N_47724,N_49917);
and UO_146 (O_146,N_49591,N_48642);
xor UO_147 (O_147,N_48992,N_48427);
nor UO_148 (O_148,N_48393,N_49577);
nand UO_149 (O_149,N_48382,N_49122);
nand UO_150 (O_150,N_48646,N_48554);
nor UO_151 (O_151,N_49479,N_48294);
nand UO_152 (O_152,N_48604,N_48100);
nor UO_153 (O_153,N_49021,N_48919);
or UO_154 (O_154,N_48808,N_48257);
and UO_155 (O_155,N_47607,N_49929);
or UO_156 (O_156,N_47548,N_48555);
nand UO_157 (O_157,N_48570,N_48502);
nand UO_158 (O_158,N_47727,N_48241);
nand UO_159 (O_159,N_49911,N_47960);
nand UO_160 (O_160,N_49527,N_47617);
nor UO_161 (O_161,N_48005,N_47685);
or UO_162 (O_162,N_49864,N_48356);
nor UO_163 (O_163,N_47796,N_49546);
xor UO_164 (O_164,N_48008,N_47592);
and UO_165 (O_165,N_49457,N_48226);
xor UO_166 (O_166,N_49703,N_48660);
xor UO_167 (O_167,N_48750,N_49005);
nand UO_168 (O_168,N_48103,N_48397);
nand UO_169 (O_169,N_48218,N_47596);
or UO_170 (O_170,N_47980,N_49829);
nor UO_171 (O_171,N_49690,N_47623);
xnor UO_172 (O_172,N_48834,N_48907);
nor UO_173 (O_173,N_48514,N_47537);
nor UO_174 (O_174,N_49305,N_49535);
nand UO_175 (O_175,N_48526,N_48197);
or UO_176 (O_176,N_49880,N_48733);
nor UO_177 (O_177,N_49704,N_48291);
nor UO_178 (O_178,N_49281,N_48522);
and UO_179 (O_179,N_48151,N_49108);
xor UO_180 (O_180,N_48260,N_48616);
and UO_181 (O_181,N_49317,N_48680);
xor UO_182 (O_182,N_49696,N_47840);
nand UO_183 (O_183,N_48816,N_49018);
or UO_184 (O_184,N_49068,N_48295);
and UO_185 (O_185,N_49332,N_49440);
nand UO_186 (O_186,N_49895,N_49373);
nand UO_187 (O_187,N_48126,N_48908);
nor UO_188 (O_188,N_48950,N_47802);
xnor UO_189 (O_189,N_49267,N_48417);
or UO_190 (O_190,N_48265,N_48556);
xor UO_191 (O_191,N_49488,N_47574);
or UO_192 (O_192,N_49672,N_48692);
nor UO_193 (O_193,N_49733,N_48086);
or UO_194 (O_194,N_47653,N_48690);
or UO_195 (O_195,N_48184,N_49545);
or UO_196 (O_196,N_48611,N_47722);
nand UO_197 (O_197,N_49407,N_49255);
xor UO_198 (O_198,N_47819,N_49042);
nor UO_199 (O_199,N_49562,N_48895);
xor UO_200 (O_200,N_49828,N_49427);
nor UO_201 (O_201,N_47931,N_48096);
nand UO_202 (O_202,N_47929,N_49298);
xor UO_203 (O_203,N_47988,N_47612);
nor UO_204 (O_204,N_49314,N_49796);
and UO_205 (O_205,N_49885,N_48753);
nand UO_206 (O_206,N_49388,N_49404);
or UO_207 (O_207,N_49259,N_48289);
nand UO_208 (O_208,N_48843,N_49291);
and UO_209 (O_209,N_48565,N_49453);
nand UO_210 (O_210,N_49253,N_49817);
or UO_211 (O_211,N_48303,N_49491);
nand UO_212 (O_212,N_49730,N_47587);
xor UO_213 (O_213,N_47975,N_47669);
nand UO_214 (O_214,N_48443,N_47904);
xor UO_215 (O_215,N_48696,N_48507);
or UO_216 (O_216,N_47759,N_48701);
and UO_217 (O_217,N_48138,N_47730);
nor UO_218 (O_218,N_47970,N_47575);
xnor UO_219 (O_219,N_48014,N_48520);
nor UO_220 (O_220,N_48255,N_48671);
nand UO_221 (O_221,N_49312,N_47506);
nand UO_222 (O_222,N_49556,N_49883);
or UO_223 (O_223,N_49415,N_47728);
or UO_224 (O_224,N_48756,N_49270);
nor UO_225 (O_225,N_49446,N_47739);
nor UO_226 (O_226,N_48549,N_49376);
or UO_227 (O_227,N_49081,N_49629);
nor UO_228 (O_228,N_49856,N_48191);
and UO_229 (O_229,N_49497,N_49614);
nand UO_230 (O_230,N_49344,N_49115);
or UO_231 (O_231,N_47568,N_48028);
and UO_232 (O_232,N_47869,N_49525);
nor UO_233 (O_233,N_49445,N_48416);
or UO_234 (O_234,N_49451,N_48117);
nor UO_235 (O_235,N_47521,N_47559);
and UO_236 (O_236,N_49578,N_47577);
nor UO_237 (O_237,N_49624,N_48057);
xor UO_238 (O_238,N_49195,N_48048);
and UO_239 (O_239,N_48591,N_48183);
or UO_240 (O_240,N_49782,N_48066);
or UO_241 (O_241,N_47810,N_48124);
nor UO_242 (O_242,N_48224,N_48253);
nand UO_243 (O_243,N_49494,N_48707);
nand UO_244 (O_244,N_48905,N_48783);
or UO_245 (O_245,N_48864,N_49475);
and UO_246 (O_246,N_48988,N_48610);
xnor UO_247 (O_247,N_48451,N_49278);
nor UO_248 (O_248,N_49942,N_49040);
and UO_249 (O_249,N_48383,N_47510);
or UO_250 (O_250,N_49240,N_48505);
and UO_251 (O_251,N_48098,N_49262);
xnor UO_252 (O_252,N_48942,N_49878);
and UO_253 (O_253,N_48854,N_48465);
nor UO_254 (O_254,N_47848,N_48959);
nor UO_255 (O_255,N_48953,N_49652);
or UO_256 (O_256,N_48148,N_48881);
and UO_257 (O_257,N_49051,N_48340);
and UO_258 (O_258,N_47674,N_47818);
and UO_259 (O_259,N_48153,N_48192);
or UO_260 (O_260,N_48947,N_49287);
or UO_261 (O_261,N_48362,N_48106);
nand UO_262 (O_262,N_48322,N_49792);
xor UO_263 (O_263,N_48858,N_48833);
xnor UO_264 (O_264,N_49849,N_48036);
nand UO_265 (O_265,N_48107,N_49583);
or UO_266 (O_266,N_48558,N_48888);
or UO_267 (O_267,N_48494,N_49561);
xnor UO_268 (O_268,N_48921,N_48923);
or UO_269 (O_269,N_49284,N_47668);
and UO_270 (O_270,N_48053,N_47776);
xor UO_271 (O_271,N_48885,N_48608);
and UO_272 (O_272,N_48324,N_49750);
and UO_273 (O_273,N_47715,N_47528);
or UO_274 (O_274,N_49334,N_49437);
nor UO_275 (O_275,N_48419,N_49571);
xnor UO_276 (O_276,N_48603,N_47624);
nor UO_277 (O_277,N_47941,N_48976);
or UO_278 (O_278,N_47831,N_49157);
nor UO_279 (O_279,N_47882,N_49085);
nand UO_280 (O_280,N_49034,N_49549);
xnor UO_281 (O_281,N_49189,N_48618);
nand UO_282 (O_282,N_49626,N_48185);
and UO_283 (O_283,N_48728,N_48434);
xnor UO_284 (O_284,N_49924,N_47567);
and UO_285 (O_285,N_48552,N_48276);
and UO_286 (O_286,N_49615,N_49104);
xor UO_287 (O_287,N_49463,N_47600);
xnor UO_288 (O_288,N_48930,N_49164);
nor UO_289 (O_289,N_48082,N_48789);
nor UO_290 (O_290,N_48205,N_48770);
or UO_291 (O_291,N_48631,N_48848);
nor UO_292 (O_292,N_49977,N_48538);
or UO_293 (O_293,N_48463,N_48862);
xor UO_294 (O_294,N_49938,N_48830);
and UO_295 (O_295,N_49582,N_49774);
xnor UO_296 (O_296,N_48914,N_48188);
nor UO_297 (O_297,N_49303,N_48299);
or UO_298 (O_298,N_48710,N_47948);
or UO_299 (O_299,N_47725,N_49594);
nor UO_300 (O_300,N_48997,N_47809);
nand UO_301 (O_301,N_48109,N_49020);
xnor UO_302 (O_302,N_48077,N_49688);
nor UO_303 (O_303,N_49180,N_49137);
nand UO_304 (O_304,N_49434,N_49190);
xnor UO_305 (O_305,N_48059,N_49082);
or UO_306 (O_306,N_49954,N_47511);
or UO_307 (O_307,N_48513,N_49971);
nand UO_308 (O_308,N_48493,N_49502);
nand UO_309 (O_309,N_49597,N_49681);
nand UO_310 (O_310,N_48803,N_48461);
nor UO_311 (O_311,N_47945,N_47588);
nand UO_312 (O_312,N_49932,N_49286);
nand UO_313 (O_313,N_47768,N_48252);
xor UO_314 (O_314,N_47524,N_48708);
and UO_315 (O_315,N_49639,N_47635);
and UO_316 (O_316,N_49468,N_48607);
or UO_317 (O_317,N_49853,N_48566);
or UO_318 (O_318,N_49067,N_49936);
nor UO_319 (O_319,N_49587,N_48590);
or UO_320 (O_320,N_48961,N_49654);
and UO_321 (O_321,N_47550,N_48308);
or UO_322 (O_322,N_49420,N_47908);
nand UO_323 (O_323,N_47702,N_48379);
and UO_324 (O_324,N_49322,N_49118);
xor UO_325 (O_325,N_47660,N_48634);
nand UO_326 (O_326,N_48846,N_49003);
xnor UO_327 (O_327,N_48993,N_47514);
nand UO_328 (O_328,N_48755,N_49699);
xor UO_329 (O_329,N_49019,N_49749);
nor UO_330 (O_330,N_48215,N_48488);
or UO_331 (O_331,N_48633,N_48851);
xor UO_332 (O_332,N_47625,N_49133);
or UO_333 (O_333,N_48841,N_48800);
and UO_334 (O_334,N_49345,N_49403);
nor UO_335 (O_335,N_48172,N_48236);
xnor UO_336 (O_336,N_49713,N_49182);
or UO_337 (O_337,N_48105,N_47839);
nand UO_338 (O_338,N_47837,N_48580);
nand UO_339 (O_339,N_49512,N_47505);
xnor UO_340 (O_340,N_49166,N_47613);
nor UO_341 (O_341,N_48916,N_49805);
nor UO_342 (O_342,N_49510,N_48922);
or UO_343 (O_343,N_48744,N_49012);
and UO_344 (O_344,N_48287,N_49396);
nand UO_345 (O_345,N_48716,N_48562);
nand UO_346 (O_346,N_49946,N_49295);
nor UO_347 (O_347,N_48279,N_49058);
or UO_348 (O_348,N_48447,N_49496);
or UO_349 (O_349,N_48531,N_48159);
or UO_350 (O_350,N_49271,N_48544);
xor UO_351 (O_351,N_47581,N_49979);
or UO_352 (O_352,N_49325,N_47878);
nand UO_353 (O_353,N_48127,N_48296);
nand UO_354 (O_354,N_49348,N_47691);
or UO_355 (O_355,N_48046,N_48043);
nand UO_356 (O_356,N_49090,N_49656);
nand UO_357 (O_357,N_47565,N_49692);
or UO_358 (O_358,N_47939,N_49554);
or UO_359 (O_359,N_48943,N_48035);
and UO_360 (O_360,N_49743,N_48817);
or UO_361 (O_361,N_48301,N_49055);
or UO_362 (O_362,N_47788,N_47573);
xor UO_363 (O_363,N_47585,N_49004);
and UO_364 (O_364,N_49473,N_49033);
and UO_365 (O_365,N_49625,N_47606);
or UO_366 (O_366,N_49331,N_49413);
nand UO_367 (O_367,N_47894,N_48766);
nor UO_368 (O_368,N_49514,N_47966);
or UO_369 (O_369,N_49037,N_49642);
nand UO_370 (O_370,N_48582,N_49184);
nor UO_371 (O_371,N_49172,N_48739);
and UO_372 (O_372,N_48492,N_49290);
and UO_373 (O_373,N_49569,N_48670);
nand UO_374 (O_374,N_48414,N_48002);
xor UO_375 (O_375,N_49646,N_49675);
nor UO_376 (O_376,N_47903,N_49657);
nor UO_377 (O_377,N_47742,N_47794);
or UO_378 (O_378,N_49237,N_48727);
or UO_379 (O_379,N_48061,N_48584);
nand UO_380 (O_380,N_47642,N_47615);
xnor UO_381 (O_381,N_48353,N_47892);
or UO_382 (O_382,N_49277,N_48790);
xnor UO_383 (O_383,N_48023,N_49891);
xnor UO_384 (O_384,N_49458,N_48189);
nand UO_385 (O_385,N_49433,N_49047);
nor UO_386 (O_386,N_47542,N_48052);
nor UO_387 (O_387,N_49472,N_49754);
xnor UO_388 (O_388,N_49050,N_47704);
and UO_389 (O_389,N_48346,N_49650);
nor UO_390 (O_390,N_48822,N_48763);
xnor UO_391 (O_391,N_47667,N_48472);
or UO_392 (O_392,N_49401,N_49564);
nand UO_393 (O_393,N_47729,N_49719);
xnor UO_394 (O_394,N_49372,N_49501);
nor UO_395 (O_395,N_48293,N_47677);
xor UO_396 (O_396,N_49212,N_49152);
or UO_397 (O_397,N_48861,N_49007);
nor UO_398 (O_398,N_48384,N_49522);
nand UO_399 (O_399,N_48683,N_48271);
nor UO_400 (O_400,N_49170,N_47735);
and UO_401 (O_401,N_49138,N_48906);
nand UO_402 (O_402,N_48087,N_47716);
xor UO_403 (O_403,N_49139,N_48457);
or UO_404 (O_404,N_48258,N_49426);
and UO_405 (O_405,N_48090,N_48659);
and UO_406 (O_406,N_48855,N_48263);
nor UO_407 (O_407,N_49310,N_49066);
or UO_408 (O_408,N_48762,N_49357);
xnor UO_409 (O_409,N_47734,N_48001);
nor UO_410 (O_410,N_48272,N_49419);
and UO_411 (O_411,N_48632,N_48169);
or UO_412 (O_412,N_48135,N_49052);
nor UO_413 (O_413,N_49724,N_48936);
nor UO_414 (O_414,N_47862,N_49002);
or UO_415 (O_415,N_47616,N_47599);
nand UO_416 (O_416,N_49540,N_48244);
and UO_417 (O_417,N_49493,N_48491);
nor UO_418 (O_418,N_48204,N_48889);
xor UO_419 (O_419,N_48624,N_49329);
nor UO_420 (O_420,N_48688,N_49406);
nor UO_421 (O_421,N_49060,N_48425);
and UO_422 (O_422,N_48280,N_47766);
and UO_423 (O_423,N_49112,N_48083);
or UO_424 (O_424,N_48067,N_47813);
nand UO_425 (O_425,N_48229,N_49142);
xnor UO_426 (O_426,N_48483,N_49839);
or UO_427 (O_427,N_48774,N_49811);
xnor UO_428 (O_428,N_48550,N_48359);
and UO_429 (O_429,N_48548,N_48154);
nor UO_430 (O_430,N_48560,N_47757);
and UO_431 (O_431,N_49350,N_48407);
or UO_432 (O_432,N_47923,N_47566);
nor UO_433 (O_433,N_49746,N_48473);
nor UO_434 (O_434,N_48791,N_48017);
and UO_435 (O_435,N_49140,N_49899);
nor UO_436 (O_436,N_48695,N_48355);
xor UO_437 (O_437,N_49872,N_49925);
nand UO_438 (O_438,N_48878,N_47905);
and UO_439 (O_439,N_48162,N_49231);
nor UO_440 (O_440,N_48836,N_49725);
nor UO_441 (O_441,N_49299,N_49756);
nand UO_442 (O_442,N_49073,N_49983);
and UO_443 (O_443,N_48623,N_48481);
xor UO_444 (O_444,N_48275,N_49523);
and UO_445 (O_445,N_48462,N_49601);
nand UO_446 (O_446,N_48421,N_48069);
or UO_447 (O_447,N_48741,N_47965);
and UO_448 (O_448,N_48242,N_49436);
xor UO_449 (O_449,N_49837,N_47773);
nor UO_450 (O_450,N_49490,N_47997);
nand UO_451 (O_451,N_48232,N_47822);
xor UO_452 (O_452,N_48337,N_47836);
nor UO_453 (O_453,N_48912,N_48958);
or UO_454 (O_454,N_48137,N_48486);
nor UO_455 (O_455,N_49636,N_49506);
and UO_456 (O_456,N_49874,N_49534);
or UO_457 (O_457,N_49875,N_48738);
nand UO_458 (O_458,N_48418,N_47517);
and UO_459 (O_459,N_48527,N_47959);
nand UO_460 (O_460,N_49257,N_49693);
and UO_461 (O_461,N_49526,N_48837);
or UO_462 (O_462,N_48403,N_49634);
or UO_463 (O_463,N_49937,N_49224);
and UO_464 (O_464,N_47620,N_49519);
nand UO_465 (O_465,N_49635,N_47891);
and UO_466 (O_466,N_48842,N_48589);
xnor UO_467 (O_467,N_47921,N_49751);
and UO_468 (O_468,N_48795,N_49644);
and UO_469 (O_469,N_48334,N_47610);
xnor UO_470 (O_470,N_48391,N_49336);
and UO_471 (O_471,N_49919,N_49844);
and UO_472 (O_472,N_49933,N_48635);
or UO_473 (O_473,N_48525,N_47670);
nor UO_474 (O_474,N_48015,N_49198);
and UO_475 (O_475,N_48798,N_47826);
or UO_476 (O_476,N_48812,N_48645);
xnor UO_477 (O_477,N_49099,N_49282);
nor UO_478 (O_478,N_49605,N_48251);
nor UO_479 (O_479,N_48377,N_49548);
or UO_480 (O_480,N_49176,N_49351);
xnor UO_481 (O_481,N_49850,N_48974);
nor UO_482 (O_482,N_48369,N_48092);
xnor UO_483 (O_483,N_48037,N_49304);
nor UO_484 (O_484,N_49843,N_47895);
nor UO_485 (O_485,N_48933,N_49720);
xnor UO_486 (O_486,N_47935,N_48897);
nand UO_487 (O_487,N_49945,N_48975);
and UO_488 (O_488,N_47541,N_49788);
xnor UO_489 (O_489,N_49913,N_49533);
or UO_490 (O_490,N_47732,N_49598);
nand UO_491 (O_491,N_48506,N_48573);
xor UO_492 (O_492,N_47961,N_49400);
xor UO_493 (O_493,N_48012,N_49387);
or UO_494 (O_494,N_47709,N_48532);
and UO_495 (O_495,N_49397,N_49341);
nor UO_496 (O_496,N_48681,N_48332);
and UO_497 (O_497,N_48734,N_47601);
nor UO_498 (O_498,N_49342,N_47876);
and UO_499 (O_499,N_48469,N_49981);
nor UO_500 (O_500,N_49680,N_48423);
or UO_501 (O_501,N_48743,N_48214);
xnor UO_502 (O_502,N_47689,N_49248);
nor UO_503 (O_503,N_49976,N_49054);
nor UO_504 (O_504,N_47851,N_49043);
and UO_505 (O_505,N_49617,N_49130);
nand UO_506 (O_506,N_47733,N_48440);
nor UO_507 (O_507,N_47621,N_49006);
or UO_508 (O_508,N_48339,N_48406);
and UO_509 (O_509,N_47540,N_48342);
or UO_510 (O_510,N_49061,N_49668);
or UO_511 (O_511,N_48787,N_47936);
nand UO_512 (O_512,N_49013,N_48927);
xor UO_513 (O_513,N_48792,N_49669);
or UO_514 (O_514,N_49481,N_49912);
nor UO_515 (O_515,N_49249,N_49778);
nand UO_516 (O_516,N_48031,N_49842);
xor UO_517 (O_517,N_47500,N_49503);
nand UO_518 (O_518,N_49588,N_49430);
and UO_519 (O_519,N_49092,N_49620);
nor UO_520 (O_520,N_47853,N_49324);
and UO_521 (O_521,N_48182,N_49110);
xor UO_522 (O_522,N_47502,N_49236);
nand UO_523 (O_523,N_48647,N_48387);
nand UO_524 (O_524,N_49323,N_49366);
nand UO_525 (O_525,N_48163,N_49560);
and UO_526 (O_526,N_47781,N_47954);
or UO_527 (O_527,N_48667,N_49990);
or UO_528 (O_528,N_48799,N_47637);
or UO_529 (O_529,N_48981,N_49083);
xnor UO_530 (O_530,N_48559,N_47763);
nand UO_531 (O_531,N_47774,N_47560);
nand UO_532 (O_532,N_48333,N_47957);
nand UO_533 (O_533,N_48298,N_48484);
nand UO_534 (O_534,N_49024,N_48831);
or UO_535 (O_535,N_49168,N_49592);
nand UO_536 (O_536,N_47815,N_47780);
and UO_537 (O_537,N_48129,N_48006);
nor UO_538 (O_538,N_49349,N_49340);
and UO_539 (O_539,N_47756,N_48725);
nand UO_540 (O_540,N_49192,N_49223);
or UO_541 (O_541,N_48721,N_49049);
nor UO_542 (O_542,N_49768,N_49294);
nand UO_543 (O_543,N_49854,N_47651);
xor UO_544 (O_544,N_47887,N_49764);
nand UO_545 (O_545,N_48963,N_47838);
nand UO_546 (O_546,N_47958,N_49347);
nand UO_547 (O_547,N_47614,N_49315);
or UO_548 (O_548,N_47569,N_49836);
nor UO_549 (O_549,N_49799,N_47890);
or UO_550 (O_550,N_48349,N_47549);
xnor UO_551 (O_551,N_47563,N_48439);
xor UO_552 (O_552,N_49802,N_47803);
xnor UO_553 (O_553,N_48654,N_48478);
nor UO_554 (O_554,N_48065,N_49023);
nor UO_555 (O_555,N_48786,N_47865);
or UO_556 (O_556,N_49200,N_48209);
and UO_557 (O_557,N_49823,N_48567);
nor UO_558 (O_558,N_47604,N_49529);
and UO_559 (O_559,N_49460,N_48150);
or UO_560 (O_560,N_49266,N_48445);
nand UO_561 (O_561,N_47650,N_48247);
or UO_562 (O_562,N_48371,N_47909);
xnor UO_563 (O_563,N_49311,N_48133);
and UO_564 (O_564,N_49359,N_49245);
and UO_565 (O_565,N_49611,N_47866);
or UO_566 (O_566,N_48345,N_47998);
xnor UO_567 (O_567,N_48920,N_47979);
nand UO_568 (O_568,N_48099,N_49742);
or UO_569 (O_569,N_49030,N_49498);
xnor UO_570 (O_570,N_49179,N_48283);
and UO_571 (O_571,N_49461,N_49539);
and UO_572 (O_572,N_48503,N_48155);
or UO_573 (O_573,N_49716,N_48026);
nor UO_574 (O_574,N_48649,N_48962);
nor UO_575 (O_575,N_48076,N_48969);
and UO_576 (O_576,N_49505,N_48140);
xor UO_577 (O_577,N_48380,N_48330);
xor UO_578 (O_578,N_48436,N_49466);
nand UO_579 (O_579,N_47527,N_47582);
nor UO_580 (O_580,N_48309,N_47833);
nor UO_581 (O_581,N_47856,N_48071);
xnor UO_582 (O_582,N_49804,N_49113);
or UO_583 (O_583,N_48320,N_48211);
xnor UO_584 (O_584,N_48745,N_49700);
nand UO_585 (O_585,N_49795,N_48111);
and UO_586 (O_586,N_49125,N_48877);
and UO_587 (O_587,N_48760,N_49220);
or UO_588 (O_588,N_47751,N_49813);
nand UO_589 (O_589,N_48428,N_48267);
nor UO_590 (O_590,N_47849,N_47772);
nand UO_591 (O_591,N_49383,N_48402);
and UO_592 (O_592,N_47754,N_48772);
xnor UO_593 (O_593,N_49706,N_48170);
nor UO_594 (O_594,N_48758,N_49621);
nor UO_595 (O_595,N_49177,N_47618);
xor UO_596 (O_596,N_47951,N_48498);
nand UO_597 (O_597,N_48778,N_49957);
xor UO_598 (O_598,N_48000,N_49053);
xor UO_599 (O_599,N_47854,N_48097);
nand UO_600 (O_600,N_47649,N_48684);
xor UO_601 (O_601,N_49059,N_48054);
or UO_602 (O_602,N_48143,N_49568);
nor UO_603 (O_603,N_49653,N_48731);
xor UO_604 (O_604,N_48452,N_49785);
nand UO_605 (O_605,N_49328,N_49586);
or UO_606 (O_606,N_48574,N_48222);
or UO_607 (O_607,N_47828,N_49408);
xor UO_608 (O_608,N_48957,N_49450);
nand UO_609 (O_609,N_49103,N_47857);
and UO_610 (O_610,N_48027,N_48292);
nor UO_611 (O_611,N_49205,N_49385);
nand UO_612 (O_612,N_49607,N_49884);
xor UO_613 (O_613,N_49074,N_49886);
xor UO_614 (O_614,N_49968,N_49963);
and UO_615 (O_615,N_49072,N_47552);
nor UO_616 (O_616,N_49612,N_49951);
nor UO_617 (O_617,N_48894,N_47798);
nor UO_618 (O_618,N_48945,N_48941);
or UO_619 (O_619,N_47745,N_48599);
or UO_620 (O_620,N_47902,N_48458);
xor UO_621 (O_621,N_48310,N_48376);
xnor UO_622 (O_622,N_49852,N_49552);
xor UO_623 (O_623,N_49222,N_49674);
nor UO_624 (O_624,N_47700,N_48887);
or UO_625 (O_625,N_48213,N_49800);
and UO_626 (O_626,N_48408,N_49559);
and UO_627 (O_627,N_48735,N_49908);
and UO_628 (O_628,N_48777,N_48325);
nand UO_629 (O_629,N_49748,N_48999);
nor UO_630 (O_630,N_47526,N_49982);
nand UO_631 (O_631,N_49643,N_48813);
xor UO_632 (O_632,N_49309,N_48044);
or UO_633 (O_633,N_48022,N_49909);
xor UO_634 (O_634,N_48719,N_48101);
and UO_635 (O_635,N_49530,N_47884);
and UO_636 (O_636,N_47932,N_49263);
and UO_637 (O_637,N_49338,N_48482);
nor UO_638 (O_638,N_49896,N_48186);
or UO_639 (O_639,N_49382,N_48536);
nor UO_640 (O_640,N_48062,N_49132);
nor UO_641 (O_641,N_49127,N_48219);
nand UO_642 (O_642,N_49469,N_49664);
xnor UO_643 (O_643,N_48693,N_48651);
xor UO_644 (O_644,N_49379,N_48277);
and UO_645 (O_645,N_48165,N_48198);
nand UO_646 (O_646,N_49293,N_47647);
nand UO_647 (O_647,N_49213,N_47812);
nor UO_648 (O_648,N_49045,N_48730);
nand UO_649 (O_649,N_49555,N_47740);
and UO_650 (O_650,N_49914,N_47817);
and UO_651 (O_651,N_47571,N_48480);
nand UO_652 (O_652,N_47519,N_49893);
nor UO_653 (O_653,N_49321,N_49685);
and UO_654 (O_654,N_48637,N_49029);
and UO_655 (O_655,N_47741,N_48305);
and UO_656 (O_656,N_48080,N_47814);
or UO_657 (O_657,N_48891,N_47872);
nand UO_658 (O_658,N_48900,N_48652);
nor UO_659 (O_659,N_48839,N_48225);
or UO_660 (O_660,N_49187,N_47787);
nand UO_661 (O_661,N_47723,N_48370);
nor UO_662 (O_662,N_48764,N_48768);
or UO_663 (O_663,N_49851,N_47832);
nand UO_664 (O_664,N_49485,N_49777);
and UO_665 (O_665,N_47864,N_49478);
or UO_666 (O_666,N_48374,N_48726);
xnor UO_667 (O_667,N_47978,N_49965);
nor UO_668 (O_668,N_48130,N_48108);
and UO_669 (O_669,N_47634,N_49824);
xor UO_670 (O_670,N_48949,N_48918);
and UO_671 (O_671,N_47744,N_49651);
nand UO_672 (O_672,N_48468,N_49819);
nor UO_673 (O_673,N_48411,N_48288);
nor UO_674 (O_674,N_48246,N_49000);
xnor UO_675 (O_675,N_49456,N_49581);
nand UO_676 (O_676,N_48866,N_49662);
nor UO_677 (O_677,N_48765,N_49755);
nor UO_678 (O_678,N_48901,N_48413);
nand UO_679 (O_679,N_49969,N_48114);
and UO_680 (O_680,N_47750,N_48759);
or UO_681 (O_681,N_49958,N_48593);
xor UO_682 (O_682,N_47515,N_47655);
or UO_683 (O_683,N_48517,N_47844);
nor UO_684 (O_684,N_49343,N_48653);
nand UO_685 (O_685,N_48016,N_48422);
or UO_686 (O_686,N_49178,N_48956);
or UO_687 (O_687,N_47529,N_47562);
xnor UO_688 (O_688,N_49010,N_49753);
and UO_689 (O_689,N_49360,N_48576);
and UO_690 (O_690,N_48487,N_47913);
nor UO_691 (O_691,N_48705,N_49016);
nand UO_692 (O_692,N_48815,N_49459);
and UO_693 (O_693,N_49056,N_48313);
xnor UO_694 (O_694,N_48347,N_49038);
nor UO_695 (O_695,N_49665,N_47544);
xor UO_696 (O_696,N_49031,N_48025);
and UO_697 (O_697,N_49953,N_48373);
nand UO_698 (O_698,N_49246,N_49337);
nand UO_699 (O_699,N_48801,N_49117);
xnor UO_700 (O_700,N_48702,N_48078);
xnor UO_701 (O_701,N_49712,N_49695);
and UO_702 (O_702,N_47580,N_48085);
xnor UO_703 (O_703,N_49833,N_48656);
nand UO_704 (O_704,N_48357,N_48496);
and UO_705 (O_705,N_49944,N_48112);
or UO_706 (O_706,N_49243,N_48395);
nand UO_707 (O_707,N_48985,N_47795);
nand UO_708 (O_708,N_47726,N_48828);
xor UO_709 (O_709,N_49678,N_49239);
nand UO_710 (O_710,N_49910,N_47737);
nor UO_711 (O_711,N_47643,N_48754);
xnor UO_712 (O_712,N_48825,N_49791);
and UO_713 (O_713,N_48674,N_49691);
and UO_714 (O_714,N_47501,N_48136);
nor UO_715 (O_715,N_49206,N_47898);
xor UO_716 (O_716,N_48358,N_48058);
nand UO_717 (O_717,N_49275,N_49028);
nand UO_718 (O_718,N_49721,N_47557);
and UO_719 (O_719,N_47707,N_48147);
and UO_720 (O_720,N_49930,N_49572);
or UO_721 (O_721,N_47940,N_48965);
or UO_722 (O_722,N_48910,N_49816);
and UO_723 (O_723,N_49927,N_48234);
and UO_724 (O_724,N_49998,N_48068);
nand UO_725 (O_725,N_49476,N_47767);
nor UO_726 (O_726,N_49422,N_49504);
nor UO_727 (O_727,N_48648,N_48158);
xor UO_728 (O_728,N_49790,N_48629);
nor UO_729 (O_729,N_47622,N_48426);
or UO_730 (O_730,N_49789,N_49989);
and UO_731 (O_731,N_48269,N_48641);
and UO_732 (O_732,N_47863,N_48329);
or UO_733 (O_733,N_48348,N_47694);
nor UO_734 (O_734,N_47842,N_49509);
nor UO_735 (O_735,N_48886,N_48038);
or UO_736 (O_736,N_48781,N_48775);
or UO_737 (O_737,N_49120,N_49288);
nand UO_738 (O_738,N_48306,N_49941);
xor UO_739 (O_739,N_48274,N_48850);
nand UO_740 (O_740,N_48898,N_49711);
nand UO_741 (O_741,N_49191,N_49470);
or UO_742 (O_742,N_49515,N_49840);
xor UO_743 (O_743,N_48818,N_47926);
nor UO_744 (O_744,N_48697,N_47712);
nand UO_745 (O_745,N_48952,N_47995);
xor UO_746 (O_746,N_48686,N_48351);
and UO_747 (O_747,N_47638,N_48578);
and UO_748 (O_748,N_49390,N_49558);
or UO_749 (O_749,N_48873,N_49825);
nor UO_750 (O_750,N_48372,N_48748);
nand UO_751 (O_751,N_49727,N_48404);
nor UO_752 (O_752,N_49538,N_47900);
nand UO_753 (O_753,N_48547,N_49900);
nor UO_754 (O_754,N_49057,N_47584);
nand UO_755 (O_755,N_48019,N_49573);
nand UO_756 (O_756,N_47984,N_49221);
nor UO_757 (O_757,N_49760,N_49831);
nand UO_758 (O_758,N_48863,N_47949);
or UO_759 (O_759,N_47671,N_48315);
xor UO_760 (O_760,N_49962,N_49499);
and UO_761 (O_761,N_49943,N_49279);
and UO_762 (O_762,N_49482,N_49173);
and UO_763 (O_763,N_49858,N_48523);
xor UO_764 (O_764,N_48840,N_49516);
nor UO_765 (O_765,N_49416,N_48511);
and UO_766 (O_766,N_49835,N_48655);
or UO_767 (O_767,N_49464,N_48715);
and UO_768 (O_768,N_49740,N_48820);
xnor UO_769 (O_769,N_49320,N_48989);
or UO_770 (O_770,N_48806,N_48110);
nor UO_771 (O_771,N_48661,N_49227);
nand UO_772 (O_772,N_48375,N_48466);
xor UO_773 (O_773,N_48075,N_48852);
and UO_774 (O_774,N_49106,N_49098);
and UO_775 (O_775,N_48157,N_49887);
or UO_776 (O_776,N_48319,N_47738);
nor UO_777 (O_777,N_48235,N_49409);
xnor UO_778 (O_778,N_49901,N_48911);
nand UO_779 (O_779,N_49044,N_47917);
xnor UO_780 (O_780,N_49449,N_48824);
nor UO_781 (O_781,N_48116,N_48094);
nor UO_782 (O_782,N_48968,N_48300);
nand UO_783 (O_783,N_49335,N_47530);
xnor UO_784 (O_784,N_47546,N_48449);
or UO_785 (O_785,N_49186,N_48729);
nor UO_786 (O_786,N_49149,N_48606);
or UO_787 (O_787,N_47697,N_48297);
nand UO_788 (O_788,N_49996,N_48256);
nor UO_789 (O_789,N_49296,N_49967);
nand UO_790 (O_790,N_48663,N_47553);
nand UO_791 (O_791,N_48771,N_48689);
nand UO_792 (O_792,N_49300,N_48829);
nor UO_793 (O_793,N_49333,N_49593);
nor UO_794 (O_794,N_48394,N_48270);
or UO_795 (O_795,N_49483,N_47874);
nor UO_796 (O_796,N_49952,N_47955);
or UO_797 (O_797,N_49435,N_49316);
nor UO_798 (O_798,N_47969,N_48442);
or UO_799 (O_799,N_49881,N_47775);
nor UO_800 (O_800,N_48409,N_49156);
or UO_801 (O_801,N_49745,N_47747);
or UO_802 (O_802,N_48883,N_49705);
nand UO_803 (O_803,N_49308,N_48029);
nand UO_804 (O_804,N_49289,N_48245);
nand UO_805 (O_805,N_48261,N_49677);
nand UO_806 (O_806,N_49162,N_49418);
nor UO_807 (O_807,N_49136,N_47518);
or UO_808 (O_808,N_48857,N_48091);
nand UO_809 (O_809,N_48541,N_47698);
xnor UO_810 (O_810,N_49209,N_48302);
nand UO_811 (O_811,N_49155,N_49134);
nor UO_812 (O_812,N_48230,N_48903);
nor UO_813 (O_813,N_48595,N_49361);
nor UO_814 (O_814,N_49920,N_49814);
nor UO_815 (O_815,N_47693,N_47764);
nand UO_816 (O_816,N_47793,N_48937);
or UO_817 (O_817,N_48156,N_47628);
nand UO_818 (O_818,N_48882,N_48004);
and UO_819 (O_819,N_48388,N_47972);
nor UO_820 (O_820,N_48703,N_47953);
xor UO_821 (O_821,N_49009,N_48331);
xor UO_822 (O_822,N_47897,N_47943);
or UO_823 (O_823,N_49492,N_49439);
and UO_824 (O_824,N_48233,N_49097);
nand UO_825 (O_825,N_49307,N_49803);
or UO_826 (O_826,N_49826,N_48769);
nand UO_827 (O_827,N_48588,N_47595);
xnor UO_828 (O_828,N_48679,N_49026);
nand UO_829 (O_829,N_49465,N_47808);
nand UO_830 (O_830,N_49661,N_49444);
nand UO_831 (O_831,N_47868,N_48464);
nor UO_832 (O_832,N_48200,N_47800);
nor UO_833 (O_833,N_49196,N_48123);
and UO_834 (O_834,N_49035,N_48535);
nand UO_835 (O_835,N_49567,N_48512);
or UO_836 (O_836,N_49080,N_49632);
nand UO_837 (O_837,N_48304,N_48939);
nor UO_838 (O_838,N_48175,N_49194);
nand UO_839 (O_839,N_49595,N_48328);
or UO_840 (O_840,N_49834,N_47996);
xnor UO_841 (O_841,N_47679,N_48934);
and UO_842 (O_842,N_48585,N_49994);
nand UO_843 (O_843,N_48460,N_49032);
xor UO_844 (O_844,N_47986,N_47790);
nand UO_845 (O_845,N_48448,N_49105);
xnor UO_846 (O_846,N_47888,N_48747);
or UO_847 (O_847,N_48990,N_49732);
xor UO_848 (O_848,N_49036,N_48827);
nor UO_849 (O_849,N_48955,N_47992);
nand UO_850 (O_850,N_49609,N_49467);
xor UO_851 (O_851,N_48924,N_48557);
and UO_852 (O_852,N_49144,N_49684);
nand UO_853 (O_853,N_48125,N_49708);
xnor UO_854 (O_854,N_49153,N_47589);
xor UO_855 (O_855,N_49455,N_48196);
xnor UO_856 (O_856,N_49432,N_47934);
and UO_857 (O_857,N_48677,N_49126);
or UO_858 (O_858,N_48030,N_49346);
and UO_859 (O_859,N_49353,N_48524);
nor UO_860 (O_860,N_48767,N_48338);
xor UO_861 (O_861,N_49922,N_49091);
xor UO_862 (O_862,N_49508,N_48569);
or UO_863 (O_863,N_47703,N_48450);
nor UO_864 (O_864,N_48084,N_48579);
xnor UO_865 (O_865,N_49011,N_48055);
xor UO_866 (O_866,N_47852,N_49637);
and UO_867 (O_867,N_47843,N_48628);
and UO_868 (O_868,N_47659,N_48899);
or UO_869 (O_869,N_49386,N_49121);
and UO_870 (O_870,N_48470,N_49273);
nor UO_871 (O_871,N_49211,N_47846);
nor UO_872 (O_872,N_49820,N_48561);
xor UO_873 (O_873,N_48132,N_48571);
nand UO_874 (O_874,N_48477,N_49550);
and UO_875 (O_875,N_48049,N_49898);
xor UO_876 (O_876,N_48290,N_48007);
xor UO_877 (O_877,N_47879,N_47678);
or UO_878 (O_878,N_49585,N_47720);
and UO_879 (O_879,N_48811,N_48336);
nor UO_880 (O_880,N_48437,N_49877);
nor UO_881 (O_881,N_48176,N_48987);
xnor UO_882 (O_882,N_48711,N_49903);
nor UO_883 (O_883,N_48737,N_48951);
and UO_884 (O_884,N_49234,N_48978);
or UO_885 (O_885,N_49616,N_47859);
or UO_886 (O_886,N_48415,N_47663);
and UO_887 (O_887,N_49218,N_48564);
xnor UO_888 (O_888,N_48694,N_48471);
nor UO_889 (O_889,N_49088,N_49547);
nor UO_890 (O_890,N_48928,N_48814);
nand UO_891 (O_891,N_49214,N_49935);
or UO_892 (O_892,N_47797,N_48724);
xor UO_893 (O_893,N_48221,N_49046);
xor UO_894 (O_894,N_48644,N_49772);
or UO_895 (O_895,N_49808,N_47605);
nor UO_896 (O_896,N_48021,N_47609);
and UO_897 (O_897,N_48849,N_49551);
xor UO_898 (O_898,N_49528,N_47648);
nand UO_899 (O_899,N_48994,N_47633);
or UO_900 (O_900,N_48121,N_48278);
nand UO_901 (O_901,N_48203,N_49916);
xnor UO_902 (O_902,N_48399,N_48216);
nand UO_903 (O_903,N_49889,N_49154);
nor UO_904 (O_904,N_49687,N_48178);
xnor UO_905 (O_905,N_47779,N_48343);
nor UO_906 (O_906,N_49758,N_48627);
nand UO_907 (O_907,N_48996,N_49363);
or UO_908 (O_908,N_49973,N_47925);
and UO_909 (O_909,N_49769,N_49511);
or UO_910 (O_910,N_48207,N_47974);
or UO_911 (O_911,N_49507,N_48847);
xor UO_912 (O_912,N_49628,N_49830);
nor UO_913 (O_913,N_47554,N_47743);
nand UO_914 (O_914,N_48401,N_48779);
or UO_915 (O_915,N_49414,N_49521);
xor UO_916 (O_916,N_48821,N_49860);
nand UO_917 (O_917,N_49217,N_47816);
and UO_918 (O_918,N_49210,N_49892);
nand UO_919 (O_919,N_49389,N_49715);
or UO_920 (O_920,N_48181,N_47547);
nor UO_921 (O_921,N_48161,N_49084);
xor UO_922 (O_922,N_49486,N_49230);
nand UO_923 (O_923,N_48410,N_49775);
or UO_924 (O_924,N_49150,N_48542);
and UO_925 (O_925,N_49580,N_49219);
xnor UO_926 (O_926,N_48944,N_49428);
nand UO_927 (O_927,N_49707,N_47912);
xor UO_928 (O_928,N_49815,N_48474);
or UO_929 (O_929,N_48282,N_47785);
or UO_930 (O_930,N_48212,N_48259);
nand UO_931 (O_931,N_49065,N_48264);
nand UO_932 (O_932,N_47593,N_48228);
nand UO_933 (O_933,N_48122,N_48018);
xor UO_934 (O_934,N_49897,N_47845);
nor UO_935 (O_935,N_48722,N_48497);
xnor UO_936 (O_936,N_49531,N_48723);
nor UO_937 (O_937,N_48467,N_47503);
and UO_938 (O_938,N_49618,N_49371);
and UO_939 (O_939,N_49215,N_49627);
or UO_940 (O_940,N_48250,N_49001);
xnor UO_941 (O_941,N_47807,N_47576);
nand UO_942 (O_942,N_48070,N_49233);
or UO_943 (O_943,N_48797,N_49285);
or UO_944 (O_944,N_48672,N_48572);
xnor UO_945 (O_945,N_48479,N_49736);
and UO_946 (O_946,N_49183,N_49894);
nand UO_947 (O_947,N_48194,N_49947);
or UO_948 (O_948,N_47778,N_49649);
or UO_949 (O_949,N_48167,N_49686);
nor UO_950 (O_950,N_47919,N_48273);
xor UO_951 (O_951,N_47692,N_49633);
or UO_952 (O_952,N_49676,N_49229);
nand UO_953 (O_953,N_49879,N_47758);
nor UO_954 (O_954,N_47658,N_49424);
or UO_955 (O_955,N_49907,N_48913);
and UO_956 (O_956,N_47770,N_48805);
or UO_957 (O_957,N_48931,N_47558);
or UO_958 (O_958,N_47538,N_48892);
nor UO_959 (O_959,N_48676,N_47602);
and UO_960 (O_960,N_47835,N_49848);
nand UO_961 (O_961,N_48243,N_49116);
xor UO_962 (O_962,N_47791,N_49762);
and UO_963 (O_963,N_48386,N_49079);
and UO_964 (O_964,N_48668,N_48284);
nor UO_965 (O_965,N_49374,N_49868);
nand UO_966 (O_966,N_49041,N_47830);
nand UO_967 (O_967,N_47933,N_47531);
xnor UO_968 (O_968,N_48368,N_49174);
or UO_969 (O_969,N_47645,N_48321);
nor UO_970 (O_970,N_48639,N_47762);
nand UO_971 (O_971,N_49931,N_49606);
or UO_972 (O_972,N_48142,N_49698);
and UO_973 (O_973,N_48195,N_47999);
nand UO_974 (O_974,N_49283,N_49838);
nor UO_975 (O_975,N_47701,N_49647);
or UO_976 (O_976,N_48613,N_48954);
nor UO_977 (O_977,N_49064,N_49070);
or UO_978 (O_978,N_47918,N_49773);
nor UO_979 (O_979,N_48720,N_48034);
and UO_980 (O_980,N_47885,N_48432);
xnor UO_981 (O_981,N_49697,N_48529);
nand UO_982 (O_982,N_47875,N_49143);
xor UO_983 (O_983,N_47855,N_48367);
nor UO_984 (O_984,N_49641,N_47937);
nand UO_985 (O_985,N_48597,N_49660);
or UO_986 (O_986,N_47591,N_47705);
and UO_987 (O_987,N_48364,N_47664);
and UO_988 (O_988,N_47611,N_49574);
nor UO_989 (O_989,N_49027,N_48424);
nor UO_990 (O_990,N_48088,N_48223);
nand UO_991 (O_991,N_48665,N_48064);
nor UO_992 (O_992,N_49327,N_49202);
nand UO_993 (O_993,N_49771,N_49921);
nor UO_994 (O_994,N_49966,N_49923);
or UO_995 (O_995,N_49306,N_48619);
nor UO_996 (O_996,N_48079,N_48510);
nor UO_997 (O_997,N_48174,N_49822);
nor UO_998 (O_998,N_47672,N_49095);
or UO_999 (O_999,N_49135,N_49993);
xnor UO_1000 (O_1000,N_47896,N_48009);
nand UO_1001 (O_1001,N_47533,N_49368);
nand UO_1002 (O_1002,N_48326,N_47967);
nor UO_1003 (O_1003,N_49985,N_48909);
and UO_1004 (O_1004,N_49241,N_49780);
nor UO_1005 (O_1005,N_48925,N_49204);
nand UO_1006 (O_1006,N_49109,N_49101);
and UO_1007 (O_1007,N_48495,N_49806);
nor UO_1008 (O_1008,N_47641,N_49536);
nand UO_1009 (O_1009,N_47968,N_48594);
nor UO_1010 (O_1010,N_49928,N_49297);
xor UO_1011 (O_1011,N_48940,N_49847);
nor UO_1012 (O_1012,N_48890,N_49161);
nand UO_1013 (O_1013,N_49905,N_47760);
nor UO_1014 (O_1014,N_49302,N_49039);
nand UO_1015 (O_1015,N_49015,N_47656);
nand UO_1016 (O_1016,N_49991,N_48431);
nand UO_1017 (O_1017,N_49722,N_47539);
or UO_1018 (O_1018,N_48131,N_49915);
and UO_1019 (O_1019,N_48915,N_49763);
xor UO_1020 (O_1020,N_47769,N_49682);
nor UO_1021 (O_1021,N_49999,N_48093);
or UO_1022 (O_1022,N_48119,N_47753);
xor UO_1023 (O_1023,N_49752,N_49997);
nand UO_1024 (O_1024,N_49956,N_47985);
xor UO_1025 (O_1025,N_49735,N_49146);
xor UO_1026 (O_1026,N_49158,N_47561);
nand UO_1027 (O_1027,N_49489,N_49679);
nor UO_1028 (O_1028,N_48780,N_49244);
or UO_1029 (O_1029,N_48518,N_49384);
and UO_1030 (O_1030,N_47608,N_49276);
xnor UO_1031 (O_1031,N_47513,N_49429);
nand UO_1032 (O_1032,N_47680,N_48794);
nor UO_1033 (O_1033,N_48217,N_49631);
nor UO_1034 (O_1034,N_49364,N_47662);
nand UO_1035 (O_1035,N_49017,N_48534);
xnor UO_1036 (O_1036,N_48238,N_49063);
nor UO_1037 (O_1037,N_49129,N_48361);
or UO_1038 (O_1038,N_48835,N_48231);
nor UO_1039 (O_1039,N_47711,N_48420);
nor UO_1040 (O_1040,N_49477,N_48360);
xor UO_1041 (O_1041,N_48352,N_47749);
and UO_1042 (O_1042,N_47676,N_47586);
nand UO_1043 (O_1043,N_49737,N_48626);
or UO_1044 (O_1044,N_47520,N_48509);
xor UO_1045 (O_1045,N_48717,N_49718);
nor UO_1046 (O_1046,N_48832,N_49845);
and UO_1047 (O_1047,N_48998,N_48489);
nor UO_1048 (O_1048,N_47870,N_47889);
nor UO_1049 (O_1049,N_48845,N_47640);
xor UO_1050 (O_1050,N_47504,N_47522);
xor UO_1051 (O_1051,N_48210,N_49949);
nand UO_1052 (O_1052,N_48040,N_49784);
and UO_1053 (O_1053,N_48598,N_48013);
nand UO_1054 (O_1054,N_49087,N_49939);
and UO_1055 (O_1055,N_49659,N_48010);
xnor UO_1056 (O_1056,N_47994,N_47632);
nor UO_1057 (O_1057,N_49330,N_48312);
or UO_1058 (O_1058,N_49014,N_49986);
nor UO_1059 (O_1059,N_47721,N_48691);
xnor UO_1060 (O_1060,N_48669,N_48736);
or UO_1061 (O_1061,N_49423,N_47535);
and UO_1062 (O_1062,N_48521,N_48967);
and UO_1063 (O_1063,N_48796,N_49599);
xor UO_1064 (O_1064,N_49185,N_48751);
or UO_1065 (O_1065,N_48050,N_47827);
and UO_1066 (O_1066,N_49123,N_47578);
and UO_1067 (O_1067,N_47644,N_49818);
or UO_1068 (O_1068,N_49807,N_48867);
xor UO_1069 (O_1069,N_48045,N_49859);
nor UO_1070 (O_1070,N_49801,N_49728);
or UO_1071 (O_1071,N_47594,N_47990);
nand UO_1072 (O_1072,N_48400,N_49950);
and UO_1073 (O_1073,N_47906,N_47910);
or UO_1074 (O_1074,N_48389,N_48095);
xnor UO_1075 (O_1075,N_49405,N_49988);
xnor UO_1076 (O_1076,N_47597,N_48685);
xnor UO_1077 (O_1077,N_48187,N_48072);
xor UO_1078 (O_1078,N_47690,N_49447);
nor UO_1079 (O_1079,N_49410,N_49377);
nor UO_1080 (O_1080,N_49500,N_47532);
or UO_1081 (O_1081,N_49356,N_49918);
or UO_1082 (O_1082,N_48809,N_49841);
nand UO_1083 (O_1083,N_49448,N_48405);
nand UO_1084 (O_1084,N_49667,N_49741);
nor UO_1085 (O_1085,N_47512,N_47686);
or UO_1086 (O_1086,N_49984,N_49268);
xor UO_1087 (O_1087,N_48638,N_48220);
xnor UO_1088 (O_1088,N_48948,N_49541);
xnor UO_1089 (O_1089,N_48982,N_49128);
and UO_1090 (O_1090,N_47950,N_49367);
nand UO_1091 (O_1091,N_47755,N_48612);
and UO_1092 (O_1092,N_49553,N_49701);
and UO_1093 (O_1093,N_48807,N_48051);
nor UO_1094 (O_1094,N_49821,N_48193);
nor UO_1095 (O_1095,N_48995,N_48605);
xnor UO_1096 (O_1096,N_49566,N_48318);
nor UO_1097 (O_1097,N_49729,N_48501);
and UO_1098 (O_1098,N_47880,N_49354);
nor UO_1099 (O_1099,N_49565,N_49114);
and UO_1100 (O_1100,N_47799,N_48872);
xnor UO_1101 (O_1101,N_49226,N_48042);
xor UO_1102 (O_1102,N_48875,N_48545);
xor UO_1103 (O_1103,N_48160,N_47636);
and UO_1104 (O_1104,N_47717,N_49694);
or UO_1105 (O_1105,N_48884,N_49734);
and UO_1106 (O_1106,N_48856,N_48917);
nor UO_1107 (O_1107,N_49906,N_47598);
xnor UO_1108 (O_1108,N_48986,N_49890);
and UO_1109 (O_1109,N_48640,N_49873);
nor UO_1110 (O_1110,N_47688,N_49524);
or UO_1111 (O_1111,N_48115,N_48528);
xor UO_1112 (O_1112,N_49871,N_48456);
and UO_1113 (O_1113,N_47682,N_49355);
and UO_1114 (O_1114,N_48039,N_48316);
nand UO_1115 (O_1115,N_48113,N_49645);
and UO_1116 (O_1116,N_49274,N_48144);
xor UO_1117 (O_1117,N_49809,N_47977);
nand UO_1118 (O_1118,N_47683,N_49454);
nor UO_1119 (O_1119,N_49228,N_48804);
xor UO_1120 (O_1120,N_47883,N_49882);
or UO_1121 (O_1121,N_48776,N_49119);
nor UO_1122 (O_1122,N_48553,N_48145);
nor UO_1123 (O_1123,N_49767,N_48617);
or UO_1124 (O_1124,N_47861,N_49714);
nand UO_1125 (O_1125,N_49995,N_49972);
and UO_1126 (O_1126,N_49159,N_48286);
nand UO_1127 (O_1127,N_48248,N_48709);
and UO_1128 (O_1128,N_47976,N_48546);
nand UO_1129 (O_1129,N_48972,N_48190);
and UO_1130 (O_1130,N_47583,N_49381);
xnor UO_1131 (O_1131,N_48390,N_49370);
nand UO_1132 (O_1132,N_48761,N_48537);
xnor UO_1133 (O_1133,N_49709,N_49442);
and UO_1134 (O_1134,N_49543,N_47777);
xor UO_1135 (O_1135,N_49970,N_48453);
nor UO_1136 (O_1136,N_48444,N_48662);
and UO_1137 (O_1137,N_47525,N_48870);
or UO_1138 (O_1138,N_48314,N_48530);
nand UO_1139 (O_1139,N_49589,N_48365);
or UO_1140 (O_1140,N_48041,N_48341);
or UO_1141 (O_1141,N_49062,N_47962);
nor UO_1142 (O_1142,N_47786,N_49160);
xor UO_1143 (O_1143,N_48964,N_49904);
or UO_1144 (O_1144,N_49077,N_48657);
and UO_1145 (O_1145,N_49623,N_47564);
xor UO_1146 (O_1146,N_48120,N_48879);
and UO_1147 (O_1147,N_49369,N_47834);
xnor UO_1148 (O_1148,N_49576,N_49702);
nor UO_1149 (O_1149,N_49391,N_48675);
xor UO_1150 (O_1150,N_48630,N_49739);
nand UO_1151 (O_1151,N_49438,N_49673);
nand UO_1152 (O_1152,N_49141,N_47860);
nand UO_1153 (O_1153,N_48970,N_49487);
nand UO_1154 (O_1154,N_48788,N_47646);
xnor UO_1155 (O_1155,N_47922,N_48398);
nand UO_1156 (O_1156,N_47652,N_49832);
and UO_1157 (O_1157,N_47695,N_48581);
nand UO_1158 (O_1158,N_47991,N_48977);
xor UO_1159 (O_1159,N_47626,N_47523);
xnor UO_1160 (O_1160,N_48732,N_49537);
nand UO_1161 (O_1161,N_48600,N_47873);
nor UO_1162 (O_1162,N_49008,N_48500);
nand UO_1163 (O_1163,N_48020,N_49812);
and UO_1164 (O_1164,N_47973,N_48838);
or UO_1165 (O_1165,N_48455,N_48499);
and UO_1166 (O_1166,N_49175,N_49960);
or UO_1167 (O_1167,N_48392,N_49726);
nand UO_1168 (O_1168,N_49723,N_49398);
nand UO_1169 (O_1169,N_48516,N_48173);
and UO_1170 (O_1170,N_48773,N_48666);
nor UO_1171 (O_1171,N_49102,N_47821);
and UO_1172 (O_1172,N_48060,N_49532);
nand UO_1173 (O_1173,N_49235,N_47914);
nand UO_1174 (O_1174,N_47661,N_49096);
nand UO_1175 (O_1175,N_49948,N_47792);
and UO_1176 (O_1176,N_48515,N_49203);
nor UO_1177 (O_1177,N_49584,N_48254);
nor UO_1178 (O_1178,N_49770,N_49866);
nor UO_1179 (O_1179,N_48971,N_48311);
and UO_1180 (O_1180,N_47899,N_49575);
nand UO_1181 (O_1181,N_49902,N_48475);
and UO_1182 (O_1182,N_49395,N_48166);
or UO_1183 (O_1183,N_48880,N_47911);
and UO_1184 (O_1184,N_48237,N_47841);
nor UO_1185 (O_1185,N_48979,N_48966);
and UO_1186 (O_1186,N_48865,N_49318);
or UO_1187 (O_1187,N_48063,N_47825);
or UO_1188 (O_1188,N_47881,N_48704);
xor UO_1189 (O_1189,N_47886,N_48350);
and UO_1190 (O_1190,N_48859,N_48714);
xor UO_1191 (O_1191,N_48378,N_47536);
and UO_1192 (O_1192,N_47907,N_49867);
and UO_1193 (O_1193,N_47696,N_49655);
or UO_1194 (O_1194,N_48551,N_48239);
xnor UO_1195 (O_1195,N_47877,N_48636);
and UO_1196 (O_1196,N_49619,N_48902);
nor UO_1197 (O_1197,N_48134,N_49417);
and UO_1198 (O_1198,N_48335,N_49793);
nand UO_1199 (O_1199,N_47938,N_49265);
nand UO_1200 (O_1200,N_49319,N_47944);
and UO_1201 (O_1201,N_48508,N_48687);
xnor UO_1202 (O_1202,N_48718,N_47782);
nand UO_1203 (O_1203,N_48206,N_48171);
or UO_1204 (O_1204,N_48991,N_47706);
or UO_1205 (O_1205,N_48164,N_48929);
xor UO_1206 (O_1206,N_49666,N_49272);
nor UO_1207 (O_1207,N_49786,N_48266);
or UO_1208 (O_1208,N_49145,N_49671);
xor UO_1209 (O_1209,N_49544,N_48650);
and UO_1210 (O_1210,N_47982,N_49365);
nand UO_1211 (O_1211,N_48102,N_49710);
nand UO_1212 (O_1212,N_48785,N_49441);
xor UO_1213 (O_1213,N_47545,N_48586);
xor UO_1214 (O_1214,N_47811,N_49761);
xnor UO_1215 (O_1215,N_48433,N_49975);
xor UO_1216 (O_1216,N_49362,N_49169);
nor UO_1217 (O_1217,N_48139,N_48446);
nor UO_1218 (O_1218,N_48540,N_47657);
nor UO_1219 (O_1219,N_49094,N_49392);
nand UO_1220 (O_1220,N_49100,N_47823);
and UO_1221 (O_1221,N_47556,N_49630);
xnor UO_1222 (O_1222,N_48973,N_47619);
xor UO_1223 (O_1223,N_49757,N_48568);
and UO_1224 (O_1224,N_48782,N_49670);
xor UO_1225 (O_1225,N_49256,N_49961);
nand UO_1226 (O_1226,N_47789,N_47784);
nand UO_1227 (O_1227,N_49151,N_49216);
xor UO_1228 (O_1228,N_49608,N_49352);
nand UO_1229 (O_1229,N_47719,N_49193);
nor UO_1230 (O_1230,N_48935,N_47684);
nand UO_1231 (O_1231,N_49124,N_49855);
nor UO_1232 (O_1232,N_48602,N_47963);
xnor UO_1233 (O_1233,N_49518,N_49188);
nand UO_1234 (O_1234,N_49048,N_48074);
or UO_1235 (O_1235,N_49992,N_49964);
nand UO_1236 (O_1236,N_49765,N_48698);
xor UO_1237 (O_1237,N_49280,N_48876);
nor UO_1238 (O_1238,N_48622,N_49798);
nor UO_1239 (O_1239,N_48152,N_48396);
and UO_1240 (O_1240,N_49292,N_49069);
nand UO_1241 (O_1241,N_47946,N_47675);
nand UO_1242 (O_1242,N_48868,N_48118);
and UO_1243 (O_1243,N_47771,N_48984);
nor UO_1244 (O_1244,N_48823,N_48893);
or UO_1245 (O_1245,N_47681,N_48749);
nand UO_1246 (O_1246,N_49846,N_47850);
nand UO_1247 (O_1247,N_49610,N_48089);
nand UO_1248 (O_1248,N_49744,N_48682);
or UO_1249 (O_1249,N_48643,N_48208);
nand UO_1250 (O_1250,N_47852,N_48575);
nor UO_1251 (O_1251,N_49736,N_48243);
or UO_1252 (O_1252,N_48266,N_49206);
xnor UO_1253 (O_1253,N_49240,N_47660);
and UO_1254 (O_1254,N_49618,N_49154);
nor UO_1255 (O_1255,N_48465,N_49967);
or UO_1256 (O_1256,N_49439,N_49455);
xnor UO_1257 (O_1257,N_47662,N_48779);
nor UO_1258 (O_1258,N_47827,N_49341);
nand UO_1259 (O_1259,N_49353,N_48757);
nor UO_1260 (O_1260,N_48954,N_47508);
or UO_1261 (O_1261,N_49460,N_49471);
xnor UO_1262 (O_1262,N_48997,N_48378);
or UO_1263 (O_1263,N_48581,N_47982);
or UO_1264 (O_1264,N_48601,N_49875);
xor UO_1265 (O_1265,N_48246,N_49634);
nor UO_1266 (O_1266,N_48206,N_48531);
and UO_1267 (O_1267,N_49273,N_48520);
nor UO_1268 (O_1268,N_48571,N_47949);
or UO_1269 (O_1269,N_49316,N_48747);
or UO_1270 (O_1270,N_47543,N_49844);
xor UO_1271 (O_1271,N_49175,N_47530);
or UO_1272 (O_1272,N_48397,N_47907);
nand UO_1273 (O_1273,N_49810,N_49634);
xnor UO_1274 (O_1274,N_49981,N_48057);
nor UO_1275 (O_1275,N_49544,N_47784);
or UO_1276 (O_1276,N_48982,N_48891);
or UO_1277 (O_1277,N_49576,N_49885);
nand UO_1278 (O_1278,N_48017,N_47726);
or UO_1279 (O_1279,N_48988,N_49671);
and UO_1280 (O_1280,N_49458,N_47620);
xor UO_1281 (O_1281,N_49082,N_47943);
and UO_1282 (O_1282,N_48855,N_49883);
xor UO_1283 (O_1283,N_49678,N_49323);
and UO_1284 (O_1284,N_49624,N_48008);
or UO_1285 (O_1285,N_48734,N_49358);
nor UO_1286 (O_1286,N_48021,N_49873);
or UO_1287 (O_1287,N_49314,N_47601);
or UO_1288 (O_1288,N_49342,N_49861);
and UO_1289 (O_1289,N_49017,N_49821);
xor UO_1290 (O_1290,N_49827,N_49614);
or UO_1291 (O_1291,N_49023,N_49004);
nand UO_1292 (O_1292,N_47595,N_47845);
nor UO_1293 (O_1293,N_48568,N_48727);
and UO_1294 (O_1294,N_48243,N_48393);
nor UO_1295 (O_1295,N_48436,N_49524);
and UO_1296 (O_1296,N_48830,N_49916);
xor UO_1297 (O_1297,N_47672,N_47873);
nand UO_1298 (O_1298,N_49231,N_49467);
and UO_1299 (O_1299,N_47669,N_48249);
xnor UO_1300 (O_1300,N_47830,N_49466);
nand UO_1301 (O_1301,N_48516,N_48545);
xnor UO_1302 (O_1302,N_49204,N_49107);
and UO_1303 (O_1303,N_48252,N_49643);
nand UO_1304 (O_1304,N_48816,N_48850);
xnor UO_1305 (O_1305,N_48762,N_48173);
or UO_1306 (O_1306,N_49497,N_49699);
nand UO_1307 (O_1307,N_48933,N_48168);
nand UO_1308 (O_1308,N_49278,N_49217);
nor UO_1309 (O_1309,N_49925,N_47619);
or UO_1310 (O_1310,N_49818,N_49088);
or UO_1311 (O_1311,N_48065,N_48217);
xnor UO_1312 (O_1312,N_49153,N_48694);
nand UO_1313 (O_1313,N_49991,N_49347);
nand UO_1314 (O_1314,N_49628,N_48766);
or UO_1315 (O_1315,N_49042,N_48849);
nand UO_1316 (O_1316,N_49353,N_48625);
and UO_1317 (O_1317,N_49000,N_48028);
xor UO_1318 (O_1318,N_48164,N_48363);
nand UO_1319 (O_1319,N_48706,N_49432);
nor UO_1320 (O_1320,N_48759,N_48319);
xnor UO_1321 (O_1321,N_49149,N_48110);
nor UO_1322 (O_1322,N_48728,N_49596);
and UO_1323 (O_1323,N_48634,N_49360);
or UO_1324 (O_1324,N_49454,N_49750);
nor UO_1325 (O_1325,N_48765,N_49187);
nor UO_1326 (O_1326,N_49004,N_48371);
nor UO_1327 (O_1327,N_48689,N_49159);
nand UO_1328 (O_1328,N_48117,N_49866);
and UO_1329 (O_1329,N_47630,N_49268);
nand UO_1330 (O_1330,N_49691,N_47582);
nand UO_1331 (O_1331,N_47713,N_49753);
nor UO_1332 (O_1332,N_47730,N_47771);
or UO_1333 (O_1333,N_49821,N_49055);
xor UO_1334 (O_1334,N_49969,N_49959);
xnor UO_1335 (O_1335,N_49796,N_49500);
or UO_1336 (O_1336,N_47896,N_48835);
and UO_1337 (O_1337,N_49561,N_48870);
nand UO_1338 (O_1338,N_47777,N_49889);
nor UO_1339 (O_1339,N_48837,N_48131);
xor UO_1340 (O_1340,N_48687,N_48087);
nor UO_1341 (O_1341,N_49760,N_49432);
xor UO_1342 (O_1342,N_49260,N_49798);
nor UO_1343 (O_1343,N_48423,N_47890);
nand UO_1344 (O_1344,N_49077,N_48368);
xor UO_1345 (O_1345,N_49347,N_48956);
nand UO_1346 (O_1346,N_48862,N_49856);
nor UO_1347 (O_1347,N_47636,N_48119);
nand UO_1348 (O_1348,N_48760,N_48490);
nand UO_1349 (O_1349,N_48374,N_48351);
and UO_1350 (O_1350,N_47508,N_49182);
or UO_1351 (O_1351,N_48192,N_48594);
nor UO_1352 (O_1352,N_48152,N_48951);
nand UO_1353 (O_1353,N_49676,N_49911);
xor UO_1354 (O_1354,N_48448,N_47844);
and UO_1355 (O_1355,N_49928,N_48525);
xor UO_1356 (O_1356,N_49456,N_49488);
nor UO_1357 (O_1357,N_48397,N_48875);
xor UO_1358 (O_1358,N_49822,N_47782);
nor UO_1359 (O_1359,N_49935,N_47538);
nand UO_1360 (O_1360,N_48918,N_48101);
and UO_1361 (O_1361,N_47631,N_49878);
and UO_1362 (O_1362,N_49621,N_48126);
nand UO_1363 (O_1363,N_48775,N_48950);
nor UO_1364 (O_1364,N_48540,N_49944);
and UO_1365 (O_1365,N_48903,N_49884);
and UO_1366 (O_1366,N_49035,N_48198);
nor UO_1367 (O_1367,N_48376,N_48083);
nand UO_1368 (O_1368,N_49655,N_49000);
nand UO_1369 (O_1369,N_49245,N_47807);
xnor UO_1370 (O_1370,N_49756,N_48531);
and UO_1371 (O_1371,N_48184,N_47702);
nor UO_1372 (O_1372,N_48476,N_49791);
xnor UO_1373 (O_1373,N_48071,N_49259);
xnor UO_1374 (O_1374,N_48148,N_49495);
and UO_1375 (O_1375,N_49888,N_48050);
nand UO_1376 (O_1376,N_47623,N_47768);
nand UO_1377 (O_1377,N_48279,N_47539);
xor UO_1378 (O_1378,N_48454,N_48184);
and UO_1379 (O_1379,N_49094,N_48865);
nor UO_1380 (O_1380,N_48782,N_49939);
and UO_1381 (O_1381,N_48070,N_48458);
nand UO_1382 (O_1382,N_48073,N_47501);
nor UO_1383 (O_1383,N_47584,N_49728);
nand UO_1384 (O_1384,N_49783,N_49541);
and UO_1385 (O_1385,N_49082,N_47606);
nor UO_1386 (O_1386,N_48618,N_47755);
nor UO_1387 (O_1387,N_48753,N_48996);
or UO_1388 (O_1388,N_49623,N_47674);
or UO_1389 (O_1389,N_48979,N_47977);
and UO_1390 (O_1390,N_48490,N_49996);
nor UO_1391 (O_1391,N_47821,N_48339);
nor UO_1392 (O_1392,N_49883,N_47877);
and UO_1393 (O_1393,N_48623,N_49522);
nor UO_1394 (O_1394,N_49833,N_47979);
nor UO_1395 (O_1395,N_49793,N_47947);
nand UO_1396 (O_1396,N_47901,N_48692);
or UO_1397 (O_1397,N_49711,N_48079);
or UO_1398 (O_1398,N_49678,N_49586);
or UO_1399 (O_1399,N_49667,N_48102);
nand UO_1400 (O_1400,N_49204,N_49337);
nand UO_1401 (O_1401,N_49046,N_48486);
and UO_1402 (O_1402,N_48834,N_48304);
xor UO_1403 (O_1403,N_47634,N_48521);
and UO_1404 (O_1404,N_48130,N_49361);
nand UO_1405 (O_1405,N_48051,N_47567);
nor UO_1406 (O_1406,N_48973,N_48043);
xor UO_1407 (O_1407,N_48496,N_48847);
xor UO_1408 (O_1408,N_49632,N_48891);
xnor UO_1409 (O_1409,N_48593,N_49211);
and UO_1410 (O_1410,N_48177,N_47877);
nand UO_1411 (O_1411,N_47622,N_49089);
nand UO_1412 (O_1412,N_49344,N_49623);
xnor UO_1413 (O_1413,N_49863,N_49113);
nand UO_1414 (O_1414,N_49329,N_47657);
or UO_1415 (O_1415,N_47948,N_47646);
xnor UO_1416 (O_1416,N_47611,N_48507);
nor UO_1417 (O_1417,N_49251,N_47546);
xnor UO_1418 (O_1418,N_48646,N_48177);
nor UO_1419 (O_1419,N_49289,N_47675);
nor UO_1420 (O_1420,N_49466,N_48933);
or UO_1421 (O_1421,N_48950,N_49537);
nor UO_1422 (O_1422,N_48224,N_47508);
nand UO_1423 (O_1423,N_49858,N_49142);
and UO_1424 (O_1424,N_49193,N_49536);
nor UO_1425 (O_1425,N_49905,N_47944);
nand UO_1426 (O_1426,N_49768,N_49607);
xor UO_1427 (O_1427,N_49781,N_49796);
nor UO_1428 (O_1428,N_47849,N_48653);
nand UO_1429 (O_1429,N_49866,N_48742);
nand UO_1430 (O_1430,N_49799,N_48500);
nand UO_1431 (O_1431,N_48128,N_49523);
xor UO_1432 (O_1432,N_49714,N_47739);
xor UO_1433 (O_1433,N_49769,N_49155);
and UO_1434 (O_1434,N_48153,N_49958);
xor UO_1435 (O_1435,N_49400,N_49752);
nor UO_1436 (O_1436,N_49130,N_49093);
nand UO_1437 (O_1437,N_48191,N_49077);
and UO_1438 (O_1438,N_47951,N_48976);
and UO_1439 (O_1439,N_49620,N_48651);
xor UO_1440 (O_1440,N_47877,N_49398);
xnor UO_1441 (O_1441,N_49511,N_49340);
xor UO_1442 (O_1442,N_49209,N_49429);
or UO_1443 (O_1443,N_47999,N_48237);
and UO_1444 (O_1444,N_48176,N_49816);
or UO_1445 (O_1445,N_49116,N_49620);
xnor UO_1446 (O_1446,N_48646,N_47770);
nand UO_1447 (O_1447,N_47594,N_48677);
nor UO_1448 (O_1448,N_48321,N_49402);
or UO_1449 (O_1449,N_48796,N_49893);
or UO_1450 (O_1450,N_49558,N_49866);
nand UO_1451 (O_1451,N_47559,N_48968);
or UO_1452 (O_1452,N_49535,N_49798);
or UO_1453 (O_1453,N_49772,N_49902);
or UO_1454 (O_1454,N_47671,N_48199);
nand UO_1455 (O_1455,N_49075,N_49267);
nand UO_1456 (O_1456,N_48887,N_49002);
nand UO_1457 (O_1457,N_48906,N_49901);
or UO_1458 (O_1458,N_47768,N_48723);
and UO_1459 (O_1459,N_48114,N_48135);
nand UO_1460 (O_1460,N_48412,N_49144);
or UO_1461 (O_1461,N_48825,N_47925);
nor UO_1462 (O_1462,N_49851,N_48036);
and UO_1463 (O_1463,N_49269,N_49453);
nor UO_1464 (O_1464,N_48366,N_48426);
nand UO_1465 (O_1465,N_47569,N_48433);
nand UO_1466 (O_1466,N_48014,N_48239);
or UO_1467 (O_1467,N_48130,N_49108);
xnor UO_1468 (O_1468,N_48617,N_49356);
and UO_1469 (O_1469,N_49671,N_48691);
nor UO_1470 (O_1470,N_48366,N_49731);
and UO_1471 (O_1471,N_48885,N_48740);
xor UO_1472 (O_1472,N_49123,N_48365);
or UO_1473 (O_1473,N_48541,N_49151);
and UO_1474 (O_1474,N_48197,N_47504);
or UO_1475 (O_1475,N_49394,N_49529);
xnor UO_1476 (O_1476,N_47652,N_48538);
and UO_1477 (O_1477,N_47791,N_49092);
nand UO_1478 (O_1478,N_48688,N_47921);
and UO_1479 (O_1479,N_48476,N_49955);
or UO_1480 (O_1480,N_49826,N_47853);
nand UO_1481 (O_1481,N_49842,N_49418);
or UO_1482 (O_1482,N_48020,N_49903);
nand UO_1483 (O_1483,N_48605,N_47845);
and UO_1484 (O_1484,N_48728,N_47733);
or UO_1485 (O_1485,N_49047,N_47842);
xnor UO_1486 (O_1486,N_47687,N_49255);
xor UO_1487 (O_1487,N_48440,N_49204);
nand UO_1488 (O_1488,N_49860,N_48255);
or UO_1489 (O_1489,N_49711,N_49187);
xor UO_1490 (O_1490,N_49428,N_49317);
nand UO_1491 (O_1491,N_48258,N_49902);
and UO_1492 (O_1492,N_48203,N_47609);
nor UO_1493 (O_1493,N_48936,N_49102);
nor UO_1494 (O_1494,N_49625,N_49364);
or UO_1495 (O_1495,N_47606,N_49444);
or UO_1496 (O_1496,N_48849,N_48970);
nand UO_1497 (O_1497,N_48431,N_47555);
xor UO_1498 (O_1498,N_49484,N_48625);
or UO_1499 (O_1499,N_48706,N_47714);
nor UO_1500 (O_1500,N_47747,N_48767);
nand UO_1501 (O_1501,N_48121,N_47689);
and UO_1502 (O_1502,N_47872,N_48220);
nor UO_1503 (O_1503,N_48778,N_48394);
or UO_1504 (O_1504,N_49544,N_47696);
or UO_1505 (O_1505,N_48116,N_48819);
and UO_1506 (O_1506,N_49418,N_49911);
nand UO_1507 (O_1507,N_48976,N_47919);
nand UO_1508 (O_1508,N_49397,N_49721);
xor UO_1509 (O_1509,N_48803,N_49439);
nor UO_1510 (O_1510,N_48418,N_48226);
or UO_1511 (O_1511,N_48071,N_47506);
xnor UO_1512 (O_1512,N_48253,N_47944);
and UO_1513 (O_1513,N_48055,N_48062);
nor UO_1514 (O_1514,N_48720,N_49976);
nor UO_1515 (O_1515,N_47802,N_48883);
or UO_1516 (O_1516,N_48975,N_49487);
xnor UO_1517 (O_1517,N_49050,N_49753);
xnor UO_1518 (O_1518,N_47542,N_49754);
xor UO_1519 (O_1519,N_48337,N_47896);
or UO_1520 (O_1520,N_48541,N_48068);
or UO_1521 (O_1521,N_49134,N_49659);
xor UO_1522 (O_1522,N_48619,N_49393);
xnor UO_1523 (O_1523,N_48501,N_48257);
nor UO_1524 (O_1524,N_47923,N_48058);
or UO_1525 (O_1525,N_49881,N_49971);
nand UO_1526 (O_1526,N_47926,N_49171);
xor UO_1527 (O_1527,N_49514,N_47606);
nor UO_1528 (O_1528,N_48933,N_49407);
or UO_1529 (O_1529,N_49556,N_48595);
or UO_1530 (O_1530,N_49018,N_47631);
nor UO_1531 (O_1531,N_49153,N_47605);
and UO_1532 (O_1532,N_47897,N_48886);
xnor UO_1533 (O_1533,N_49471,N_49083);
nor UO_1534 (O_1534,N_48451,N_48210);
or UO_1535 (O_1535,N_49129,N_48405);
xnor UO_1536 (O_1536,N_48249,N_49291);
and UO_1537 (O_1537,N_47868,N_49276);
or UO_1538 (O_1538,N_48365,N_47863);
or UO_1539 (O_1539,N_47673,N_49705);
and UO_1540 (O_1540,N_48514,N_47856);
nand UO_1541 (O_1541,N_48271,N_48952);
xor UO_1542 (O_1542,N_47558,N_48699);
xor UO_1543 (O_1543,N_49872,N_49646);
and UO_1544 (O_1544,N_48619,N_49061);
or UO_1545 (O_1545,N_48092,N_49236);
and UO_1546 (O_1546,N_48662,N_47845);
xor UO_1547 (O_1547,N_47962,N_49429);
or UO_1548 (O_1548,N_48771,N_47706);
or UO_1549 (O_1549,N_47964,N_49901);
nor UO_1550 (O_1550,N_48183,N_48971);
xnor UO_1551 (O_1551,N_49662,N_48587);
xnor UO_1552 (O_1552,N_49998,N_48560);
and UO_1553 (O_1553,N_48424,N_49736);
nand UO_1554 (O_1554,N_48690,N_49175);
nor UO_1555 (O_1555,N_49704,N_49830);
and UO_1556 (O_1556,N_49132,N_49926);
nand UO_1557 (O_1557,N_47952,N_48414);
nand UO_1558 (O_1558,N_48100,N_48677);
nand UO_1559 (O_1559,N_48904,N_48440);
xor UO_1560 (O_1560,N_49751,N_49302);
nand UO_1561 (O_1561,N_47991,N_47624);
nand UO_1562 (O_1562,N_48014,N_49625);
xor UO_1563 (O_1563,N_49807,N_48843);
or UO_1564 (O_1564,N_49713,N_49549);
nor UO_1565 (O_1565,N_49939,N_48700);
xor UO_1566 (O_1566,N_49205,N_47505);
xor UO_1567 (O_1567,N_48342,N_48003);
nand UO_1568 (O_1568,N_47749,N_48149);
and UO_1569 (O_1569,N_47820,N_49376);
nand UO_1570 (O_1570,N_47658,N_48456);
or UO_1571 (O_1571,N_48198,N_48847);
or UO_1572 (O_1572,N_48141,N_47731);
xor UO_1573 (O_1573,N_47558,N_49244);
nand UO_1574 (O_1574,N_49716,N_48827);
or UO_1575 (O_1575,N_49578,N_49058);
or UO_1576 (O_1576,N_48557,N_48976);
xor UO_1577 (O_1577,N_47575,N_49363);
and UO_1578 (O_1578,N_47865,N_49052);
or UO_1579 (O_1579,N_49667,N_47799);
xor UO_1580 (O_1580,N_47798,N_49928);
and UO_1581 (O_1581,N_48254,N_47684);
or UO_1582 (O_1582,N_47502,N_49441);
or UO_1583 (O_1583,N_48981,N_48440);
xnor UO_1584 (O_1584,N_48904,N_48101);
or UO_1585 (O_1585,N_49901,N_48202);
xnor UO_1586 (O_1586,N_47788,N_48376);
nor UO_1587 (O_1587,N_48074,N_48990);
nor UO_1588 (O_1588,N_49769,N_48940);
and UO_1589 (O_1589,N_49456,N_48225);
and UO_1590 (O_1590,N_49922,N_48164);
nand UO_1591 (O_1591,N_49907,N_47748);
nand UO_1592 (O_1592,N_48387,N_48335);
nand UO_1593 (O_1593,N_47709,N_49312);
nor UO_1594 (O_1594,N_49417,N_49134);
nor UO_1595 (O_1595,N_48578,N_47663);
nor UO_1596 (O_1596,N_47543,N_48467);
nand UO_1597 (O_1597,N_49684,N_48097);
and UO_1598 (O_1598,N_49663,N_48210);
nand UO_1599 (O_1599,N_49112,N_48343);
nor UO_1600 (O_1600,N_48584,N_48389);
nand UO_1601 (O_1601,N_48162,N_49429);
and UO_1602 (O_1602,N_49475,N_48036);
nand UO_1603 (O_1603,N_48265,N_49651);
xor UO_1604 (O_1604,N_48894,N_48788);
and UO_1605 (O_1605,N_48390,N_47822);
or UO_1606 (O_1606,N_47753,N_49962);
nand UO_1607 (O_1607,N_48364,N_47955);
nor UO_1608 (O_1608,N_49868,N_49239);
and UO_1609 (O_1609,N_48264,N_49616);
xor UO_1610 (O_1610,N_48108,N_49018);
nor UO_1611 (O_1611,N_47717,N_48121);
and UO_1612 (O_1612,N_48124,N_49806);
and UO_1613 (O_1613,N_48516,N_49538);
nand UO_1614 (O_1614,N_49631,N_49106);
xor UO_1615 (O_1615,N_48430,N_47522);
xor UO_1616 (O_1616,N_49426,N_47831);
or UO_1617 (O_1617,N_48682,N_47932);
xnor UO_1618 (O_1618,N_49401,N_49999);
and UO_1619 (O_1619,N_47705,N_49911);
nor UO_1620 (O_1620,N_48238,N_48566);
xor UO_1621 (O_1621,N_47921,N_48779);
and UO_1622 (O_1622,N_49671,N_47578);
and UO_1623 (O_1623,N_49675,N_49322);
xor UO_1624 (O_1624,N_49869,N_47520);
and UO_1625 (O_1625,N_48388,N_48872);
and UO_1626 (O_1626,N_48082,N_47918);
or UO_1627 (O_1627,N_48350,N_49860);
xor UO_1628 (O_1628,N_48181,N_48773);
and UO_1629 (O_1629,N_47621,N_48819);
and UO_1630 (O_1630,N_48635,N_48279);
nand UO_1631 (O_1631,N_49599,N_49459);
or UO_1632 (O_1632,N_48255,N_48978);
and UO_1633 (O_1633,N_48660,N_49562);
xnor UO_1634 (O_1634,N_48590,N_49134);
nor UO_1635 (O_1635,N_47892,N_47635);
and UO_1636 (O_1636,N_49918,N_48262);
and UO_1637 (O_1637,N_49323,N_47769);
nor UO_1638 (O_1638,N_49861,N_47718);
and UO_1639 (O_1639,N_49312,N_47963);
xor UO_1640 (O_1640,N_47754,N_49738);
and UO_1641 (O_1641,N_48345,N_49513);
nand UO_1642 (O_1642,N_48684,N_47524);
or UO_1643 (O_1643,N_49483,N_49786);
nor UO_1644 (O_1644,N_49330,N_49624);
nand UO_1645 (O_1645,N_49275,N_47593);
nand UO_1646 (O_1646,N_49085,N_47969);
and UO_1647 (O_1647,N_48590,N_49982);
nor UO_1648 (O_1648,N_47801,N_47949);
and UO_1649 (O_1649,N_48638,N_48986);
xor UO_1650 (O_1650,N_49490,N_48903);
xnor UO_1651 (O_1651,N_47893,N_49541);
or UO_1652 (O_1652,N_47613,N_48779);
xnor UO_1653 (O_1653,N_48234,N_49024);
nor UO_1654 (O_1654,N_49338,N_48948);
nor UO_1655 (O_1655,N_48357,N_49161);
nand UO_1656 (O_1656,N_48986,N_48428);
nor UO_1657 (O_1657,N_49693,N_48518);
xnor UO_1658 (O_1658,N_48711,N_49970);
or UO_1659 (O_1659,N_47952,N_49136);
and UO_1660 (O_1660,N_48448,N_48941);
or UO_1661 (O_1661,N_48568,N_47846);
or UO_1662 (O_1662,N_48579,N_49756);
and UO_1663 (O_1663,N_49104,N_49391);
xor UO_1664 (O_1664,N_49184,N_49791);
xor UO_1665 (O_1665,N_48547,N_48436);
nand UO_1666 (O_1666,N_49845,N_49460);
nor UO_1667 (O_1667,N_49887,N_47827);
and UO_1668 (O_1668,N_47656,N_49303);
and UO_1669 (O_1669,N_49382,N_49897);
nor UO_1670 (O_1670,N_49137,N_48379);
or UO_1671 (O_1671,N_49936,N_48430);
or UO_1672 (O_1672,N_48106,N_48868);
and UO_1673 (O_1673,N_48821,N_47528);
nand UO_1674 (O_1674,N_48642,N_48931);
and UO_1675 (O_1675,N_49771,N_49334);
nand UO_1676 (O_1676,N_49666,N_49565);
nand UO_1677 (O_1677,N_49260,N_47688);
and UO_1678 (O_1678,N_49642,N_49796);
and UO_1679 (O_1679,N_48936,N_48265);
or UO_1680 (O_1680,N_48795,N_48554);
xnor UO_1681 (O_1681,N_48621,N_48344);
nor UO_1682 (O_1682,N_47947,N_47696);
xor UO_1683 (O_1683,N_49267,N_49051);
nor UO_1684 (O_1684,N_47903,N_49132);
xor UO_1685 (O_1685,N_48122,N_49449);
or UO_1686 (O_1686,N_48845,N_48888);
or UO_1687 (O_1687,N_49174,N_48566);
nand UO_1688 (O_1688,N_49082,N_48863);
nand UO_1689 (O_1689,N_48886,N_49033);
or UO_1690 (O_1690,N_48753,N_47890);
or UO_1691 (O_1691,N_48391,N_47906);
xor UO_1692 (O_1692,N_48453,N_48062);
nand UO_1693 (O_1693,N_49253,N_49060);
nor UO_1694 (O_1694,N_47514,N_49743);
xnor UO_1695 (O_1695,N_49708,N_47624);
xnor UO_1696 (O_1696,N_48725,N_49331);
nor UO_1697 (O_1697,N_49422,N_48784);
nor UO_1698 (O_1698,N_49399,N_48888);
and UO_1699 (O_1699,N_48699,N_48310);
and UO_1700 (O_1700,N_47832,N_49307);
and UO_1701 (O_1701,N_48678,N_49431);
and UO_1702 (O_1702,N_49138,N_49191);
xnor UO_1703 (O_1703,N_49632,N_48748);
and UO_1704 (O_1704,N_48734,N_49949);
and UO_1705 (O_1705,N_48304,N_47903);
nor UO_1706 (O_1706,N_49379,N_49716);
nand UO_1707 (O_1707,N_49672,N_48866);
nand UO_1708 (O_1708,N_49131,N_49235);
or UO_1709 (O_1709,N_49072,N_49874);
or UO_1710 (O_1710,N_49463,N_48127);
or UO_1711 (O_1711,N_48796,N_49500);
or UO_1712 (O_1712,N_49974,N_48439);
or UO_1713 (O_1713,N_49329,N_49868);
nor UO_1714 (O_1714,N_48527,N_49070);
and UO_1715 (O_1715,N_49406,N_49135);
nand UO_1716 (O_1716,N_49139,N_48614);
or UO_1717 (O_1717,N_49492,N_48650);
and UO_1718 (O_1718,N_49062,N_47792);
or UO_1719 (O_1719,N_47923,N_48591);
or UO_1720 (O_1720,N_48090,N_47968);
or UO_1721 (O_1721,N_49113,N_48801);
nor UO_1722 (O_1722,N_49293,N_49036);
nor UO_1723 (O_1723,N_47742,N_48123);
nand UO_1724 (O_1724,N_47689,N_49717);
or UO_1725 (O_1725,N_48039,N_49418);
xnor UO_1726 (O_1726,N_48808,N_49288);
nand UO_1727 (O_1727,N_48994,N_48594);
xor UO_1728 (O_1728,N_49219,N_47908);
nor UO_1729 (O_1729,N_48354,N_49842);
nand UO_1730 (O_1730,N_49366,N_49839);
nand UO_1731 (O_1731,N_47786,N_48039);
or UO_1732 (O_1732,N_47554,N_48242);
xor UO_1733 (O_1733,N_49818,N_49040);
nor UO_1734 (O_1734,N_48129,N_49258);
and UO_1735 (O_1735,N_49370,N_48631);
xnor UO_1736 (O_1736,N_47835,N_48786);
xnor UO_1737 (O_1737,N_47628,N_49250);
and UO_1738 (O_1738,N_49882,N_49058);
xor UO_1739 (O_1739,N_48814,N_48321);
nor UO_1740 (O_1740,N_47671,N_47901);
xor UO_1741 (O_1741,N_47704,N_48467);
and UO_1742 (O_1742,N_49878,N_49154);
nor UO_1743 (O_1743,N_47535,N_48507);
nand UO_1744 (O_1744,N_48751,N_47658);
and UO_1745 (O_1745,N_49854,N_49631);
or UO_1746 (O_1746,N_47835,N_48699);
xnor UO_1747 (O_1747,N_49838,N_49085);
nand UO_1748 (O_1748,N_49235,N_48734);
nand UO_1749 (O_1749,N_49708,N_47730);
xor UO_1750 (O_1750,N_49682,N_49611);
or UO_1751 (O_1751,N_49659,N_49024);
xor UO_1752 (O_1752,N_49265,N_47738);
or UO_1753 (O_1753,N_49279,N_48175);
and UO_1754 (O_1754,N_48071,N_48468);
nand UO_1755 (O_1755,N_47744,N_49678);
xnor UO_1756 (O_1756,N_49570,N_48733);
nand UO_1757 (O_1757,N_48828,N_48430);
and UO_1758 (O_1758,N_49554,N_48631);
xor UO_1759 (O_1759,N_48007,N_48973);
and UO_1760 (O_1760,N_47595,N_49052);
or UO_1761 (O_1761,N_49860,N_48009);
or UO_1762 (O_1762,N_48640,N_49712);
nor UO_1763 (O_1763,N_49026,N_47518);
xor UO_1764 (O_1764,N_49994,N_47551);
and UO_1765 (O_1765,N_49053,N_47838);
or UO_1766 (O_1766,N_49669,N_49894);
nor UO_1767 (O_1767,N_48483,N_47583);
xnor UO_1768 (O_1768,N_48511,N_49626);
nor UO_1769 (O_1769,N_48781,N_47781);
nand UO_1770 (O_1770,N_49779,N_48180);
nor UO_1771 (O_1771,N_48575,N_48164);
or UO_1772 (O_1772,N_49724,N_49292);
nor UO_1773 (O_1773,N_47674,N_47736);
xnor UO_1774 (O_1774,N_48956,N_48017);
or UO_1775 (O_1775,N_48243,N_49508);
and UO_1776 (O_1776,N_47669,N_47828);
or UO_1777 (O_1777,N_49428,N_49779);
nand UO_1778 (O_1778,N_48566,N_48353);
nor UO_1779 (O_1779,N_47682,N_47833);
nor UO_1780 (O_1780,N_49151,N_48752);
xor UO_1781 (O_1781,N_48080,N_48362);
nor UO_1782 (O_1782,N_48289,N_49040);
nand UO_1783 (O_1783,N_49381,N_49545);
and UO_1784 (O_1784,N_49615,N_49925);
and UO_1785 (O_1785,N_47637,N_48825);
xnor UO_1786 (O_1786,N_48494,N_48073);
or UO_1787 (O_1787,N_48490,N_47752);
or UO_1788 (O_1788,N_47620,N_49349);
nor UO_1789 (O_1789,N_49926,N_49358);
nand UO_1790 (O_1790,N_49468,N_49667);
xnor UO_1791 (O_1791,N_49845,N_49823);
nor UO_1792 (O_1792,N_48883,N_47819);
nor UO_1793 (O_1793,N_47570,N_49613);
and UO_1794 (O_1794,N_48649,N_48738);
and UO_1795 (O_1795,N_48093,N_49650);
nand UO_1796 (O_1796,N_47790,N_49145);
xnor UO_1797 (O_1797,N_49647,N_49786);
and UO_1798 (O_1798,N_47946,N_48966);
nand UO_1799 (O_1799,N_47899,N_49069);
or UO_1800 (O_1800,N_48115,N_47623);
nor UO_1801 (O_1801,N_47822,N_49946);
or UO_1802 (O_1802,N_49266,N_49133);
nor UO_1803 (O_1803,N_49346,N_49921);
nand UO_1804 (O_1804,N_47580,N_47577);
nand UO_1805 (O_1805,N_48121,N_47687);
xor UO_1806 (O_1806,N_48974,N_47868);
xor UO_1807 (O_1807,N_48291,N_49712);
xnor UO_1808 (O_1808,N_48396,N_47630);
and UO_1809 (O_1809,N_49348,N_48320);
xnor UO_1810 (O_1810,N_49031,N_49620);
nand UO_1811 (O_1811,N_48474,N_48634);
nor UO_1812 (O_1812,N_47647,N_49042);
nor UO_1813 (O_1813,N_48034,N_48096);
and UO_1814 (O_1814,N_47926,N_49741);
nor UO_1815 (O_1815,N_48949,N_48370);
nand UO_1816 (O_1816,N_47839,N_49993);
nand UO_1817 (O_1817,N_47794,N_47708);
xor UO_1818 (O_1818,N_48945,N_48993);
and UO_1819 (O_1819,N_49326,N_49705);
nor UO_1820 (O_1820,N_49093,N_48882);
nand UO_1821 (O_1821,N_47577,N_48252);
or UO_1822 (O_1822,N_49230,N_49342);
nand UO_1823 (O_1823,N_47543,N_49621);
or UO_1824 (O_1824,N_48589,N_49142);
or UO_1825 (O_1825,N_48930,N_47578);
and UO_1826 (O_1826,N_47947,N_47999);
nand UO_1827 (O_1827,N_49457,N_49235);
nor UO_1828 (O_1828,N_49788,N_49470);
and UO_1829 (O_1829,N_49905,N_49461);
nor UO_1830 (O_1830,N_48719,N_49573);
xor UO_1831 (O_1831,N_49450,N_48578);
nand UO_1832 (O_1832,N_49607,N_49495);
nor UO_1833 (O_1833,N_49521,N_49752);
xnor UO_1834 (O_1834,N_48877,N_47592);
and UO_1835 (O_1835,N_49114,N_49175);
and UO_1836 (O_1836,N_47529,N_48493);
and UO_1837 (O_1837,N_48262,N_49497);
nor UO_1838 (O_1838,N_48318,N_48443);
or UO_1839 (O_1839,N_48528,N_48466);
nor UO_1840 (O_1840,N_49425,N_47996);
or UO_1841 (O_1841,N_47835,N_49955);
nor UO_1842 (O_1842,N_49043,N_47697);
nor UO_1843 (O_1843,N_49649,N_48049);
xnor UO_1844 (O_1844,N_49116,N_48686);
or UO_1845 (O_1845,N_48267,N_49509);
or UO_1846 (O_1846,N_49188,N_48909);
nor UO_1847 (O_1847,N_48784,N_49337);
and UO_1848 (O_1848,N_48456,N_49425);
nand UO_1849 (O_1849,N_49244,N_49930);
xor UO_1850 (O_1850,N_48052,N_48902);
or UO_1851 (O_1851,N_47636,N_47947);
or UO_1852 (O_1852,N_47854,N_47540);
and UO_1853 (O_1853,N_48912,N_49349);
xnor UO_1854 (O_1854,N_49477,N_47995);
nand UO_1855 (O_1855,N_48298,N_47688);
and UO_1856 (O_1856,N_48432,N_47851);
nor UO_1857 (O_1857,N_48432,N_47676);
or UO_1858 (O_1858,N_49170,N_49726);
nand UO_1859 (O_1859,N_49347,N_48375);
xor UO_1860 (O_1860,N_48056,N_49293);
xor UO_1861 (O_1861,N_49466,N_49402);
or UO_1862 (O_1862,N_48459,N_48060);
and UO_1863 (O_1863,N_48792,N_49003);
nand UO_1864 (O_1864,N_48504,N_48830);
nand UO_1865 (O_1865,N_48055,N_49969);
or UO_1866 (O_1866,N_48571,N_49286);
and UO_1867 (O_1867,N_47805,N_47844);
nand UO_1868 (O_1868,N_49656,N_49426);
and UO_1869 (O_1869,N_48216,N_48435);
nor UO_1870 (O_1870,N_48687,N_48776);
nor UO_1871 (O_1871,N_48409,N_49941);
xor UO_1872 (O_1872,N_49851,N_49531);
xor UO_1873 (O_1873,N_47616,N_49867);
nand UO_1874 (O_1874,N_48645,N_49442);
and UO_1875 (O_1875,N_48631,N_47587);
nor UO_1876 (O_1876,N_49260,N_48839);
nor UO_1877 (O_1877,N_48045,N_47831);
xnor UO_1878 (O_1878,N_49639,N_48917);
and UO_1879 (O_1879,N_48587,N_49125);
and UO_1880 (O_1880,N_48413,N_47518);
nor UO_1881 (O_1881,N_48213,N_49931);
xnor UO_1882 (O_1882,N_48748,N_48061);
xnor UO_1883 (O_1883,N_47560,N_48910);
or UO_1884 (O_1884,N_49713,N_49715);
and UO_1885 (O_1885,N_48376,N_48656);
nand UO_1886 (O_1886,N_49187,N_49699);
and UO_1887 (O_1887,N_48826,N_47687);
or UO_1888 (O_1888,N_49383,N_49006);
nor UO_1889 (O_1889,N_48215,N_49508);
and UO_1890 (O_1890,N_48762,N_48099);
nor UO_1891 (O_1891,N_47643,N_48454);
nor UO_1892 (O_1892,N_48544,N_49133);
xnor UO_1893 (O_1893,N_47523,N_47680);
nand UO_1894 (O_1894,N_49770,N_49241);
or UO_1895 (O_1895,N_47983,N_48236);
nand UO_1896 (O_1896,N_48470,N_47948);
nor UO_1897 (O_1897,N_48575,N_48995);
or UO_1898 (O_1898,N_47794,N_48184);
or UO_1899 (O_1899,N_48397,N_47908);
or UO_1900 (O_1900,N_49945,N_49840);
or UO_1901 (O_1901,N_48509,N_48132);
nand UO_1902 (O_1902,N_49079,N_49442);
and UO_1903 (O_1903,N_49221,N_48344);
and UO_1904 (O_1904,N_49671,N_48313);
nor UO_1905 (O_1905,N_48335,N_49365);
nand UO_1906 (O_1906,N_48183,N_48997);
xor UO_1907 (O_1907,N_49967,N_49095);
nor UO_1908 (O_1908,N_48817,N_48263);
nand UO_1909 (O_1909,N_47688,N_47590);
or UO_1910 (O_1910,N_48426,N_49629);
nand UO_1911 (O_1911,N_48255,N_48530);
or UO_1912 (O_1912,N_48805,N_47747);
and UO_1913 (O_1913,N_49051,N_48147);
nor UO_1914 (O_1914,N_49690,N_48608);
and UO_1915 (O_1915,N_48396,N_49475);
and UO_1916 (O_1916,N_49844,N_48011);
nor UO_1917 (O_1917,N_49413,N_49724);
or UO_1918 (O_1918,N_48614,N_48621);
nor UO_1919 (O_1919,N_49326,N_48453);
xor UO_1920 (O_1920,N_48994,N_48173);
and UO_1921 (O_1921,N_47823,N_49187);
xor UO_1922 (O_1922,N_48469,N_48702);
nand UO_1923 (O_1923,N_48613,N_48380);
or UO_1924 (O_1924,N_48547,N_49928);
xor UO_1925 (O_1925,N_48909,N_49013);
nor UO_1926 (O_1926,N_48668,N_48466);
nand UO_1927 (O_1927,N_47976,N_48275);
nand UO_1928 (O_1928,N_49328,N_49050);
and UO_1929 (O_1929,N_48004,N_47501);
or UO_1930 (O_1930,N_47521,N_48806);
or UO_1931 (O_1931,N_49692,N_48099);
nor UO_1932 (O_1932,N_47610,N_49943);
xnor UO_1933 (O_1933,N_49376,N_47562);
nor UO_1934 (O_1934,N_48501,N_49634);
nor UO_1935 (O_1935,N_48518,N_48708);
nand UO_1936 (O_1936,N_48434,N_49768);
and UO_1937 (O_1937,N_49645,N_47661);
nor UO_1938 (O_1938,N_49562,N_48282);
or UO_1939 (O_1939,N_49900,N_49961);
nor UO_1940 (O_1940,N_48346,N_48633);
xnor UO_1941 (O_1941,N_47592,N_47574);
nand UO_1942 (O_1942,N_49087,N_48236);
nor UO_1943 (O_1943,N_48777,N_48995);
or UO_1944 (O_1944,N_47792,N_49038);
xor UO_1945 (O_1945,N_48020,N_49196);
nand UO_1946 (O_1946,N_49998,N_48923);
xor UO_1947 (O_1947,N_49134,N_49154);
and UO_1948 (O_1948,N_49340,N_48128);
nor UO_1949 (O_1949,N_47992,N_47910);
and UO_1950 (O_1950,N_48347,N_48344);
or UO_1951 (O_1951,N_49985,N_49471);
nor UO_1952 (O_1952,N_49365,N_48463);
nor UO_1953 (O_1953,N_49187,N_48319);
nor UO_1954 (O_1954,N_47543,N_49795);
and UO_1955 (O_1955,N_49993,N_49513);
nor UO_1956 (O_1956,N_47506,N_49614);
nand UO_1957 (O_1957,N_49825,N_48767);
xnor UO_1958 (O_1958,N_48854,N_48531);
xnor UO_1959 (O_1959,N_47945,N_48028);
nor UO_1960 (O_1960,N_48113,N_49007);
and UO_1961 (O_1961,N_49120,N_47798);
or UO_1962 (O_1962,N_49011,N_47552);
and UO_1963 (O_1963,N_48799,N_49424);
or UO_1964 (O_1964,N_48720,N_49285);
nor UO_1965 (O_1965,N_48821,N_48144);
nand UO_1966 (O_1966,N_48394,N_47979);
nand UO_1967 (O_1967,N_49947,N_48545);
and UO_1968 (O_1968,N_47794,N_47610);
nor UO_1969 (O_1969,N_49060,N_49651);
xnor UO_1970 (O_1970,N_47767,N_48948);
nor UO_1971 (O_1971,N_49658,N_47801);
xnor UO_1972 (O_1972,N_49234,N_47680);
nand UO_1973 (O_1973,N_48859,N_49940);
or UO_1974 (O_1974,N_47975,N_49715);
nor UO_1975 (O_1975,N_47851,N_48689);
or UO_1976 (O_1976,N_49388,N_49047);
or UO_1977 (O_1977,N_49818,N_49077);
or UO_1978 (O_1978,N_48435,N_49825);
nand UO_1979 (O_1979,N_47790,N_47830);
xnor UO_1980 (O_1980,N_49290,N_47591);
nor UO_1981 (O_1981,N_47806,N_49034);
nor UO_1982 (O_1982,N_49285,N_49372);
nor UO_1983 (O_1983,N_48152,N_47809);
and UO_1984 (O_1984,N_49444,N_48284);
xor UO_1985 (O_1985,N_47738,N_47675);
nand UO_1986 (O_1986,N_48012,N_49157);
nand UO_1987 (O_1987,N_48631,N_48649);
and UO_1988 (O_1988,N_49031,N_49414);
nand UO_1989 (O_1989,N_48828,N_48897);
xor UO_1990 (O_1990,N_47953,N_49764);
and UO_1991 (O_1991,N_47806,N_49703);
and UO_1992 (O_1992,N_49847,N_49917);
and UO_1993 (O_1993,N_48269,N_49758);
xor UO_1994 (O_1994,N_47691,N_49908);
and UO_1995 (O_1995,N_47614,N_49417);
xnor UO_1996 (O_1996,N_49241,N_47827);
xor UO_1997 (O_1997,N_49567,N_47780);
or UO_1998 (O_1998,N_49321,N_47688);
and UO_1999 (O_1999,N_48290,N_48116);
and UO_2000 (O_2000,N_49764,N_49210);
and UO_2001 (O_2001,N_48590,N_48801);
nand UO_2002 (O_2002,N_47719,N_48003);
nor UO_2003 (O_2003,N_49384,N_49848);
xnor UO_2004 (O_2004,N_49434,N_47931);
xor UO_2005 (O_2005,N_48015,N_48888);
nor UO_2006 (O_2006,N_48062,N_48856);
nand UO_2007 (O_2007,N_49392,N_48993);
xnor UO_2008 (O_2008,N_49505,N_49187);
xnor UO_2009 (O_2009,N_47553,N_47825);
nand UO_2010 (O_2010,N_48900,N_47537);
or UO_2011 (O_2011,N_48746,N_47693);
nand UO_2012 (O_2012,N_49729,N_47567);
or UO_2013 (O_2013,N_49861,N_49994);
xor UO_2014 (O_2014,N_48763,N_48276);
nand UO_2015 (O_2015,N_49474,N_48754);
nand UO_2016 (O_2016,N_49722,N_47696);
xnor UO_2017 (O_2017,N_48314,N_48231);
nand UO_2018 (O_2018,N_49380,N_48163);
nor UO_2019 (O_2019,N_49396,N_47715);
nand UO_2020 (O_2020,N_49483,N_49209);
and UO_2021 (O_2021,N_48841,N_48090);
and UO_2022 (O_2022,N_47510,N_47702);
or UO_2023 (O_2023,N_48637,N_48423);
nor UO_2024 (O_2024,N_47580,N_47655);
and UO_2025 (O_2025,N_48743,N_48602);
nor UO_2026 (O_2026,N_48779,N_48198);
xnor UO_2027 (O_2027,N_48538,N_47895);
nand UO_2028 (O_2028,N_49453,N_47998);
or UO_2029 (O_2029,N_48973,N_47959);
or UO_2030 (O_2030,N_48657,N_48519);
nand UO_2031 (O_2031,N_48692,N_48020);
xor UO_2032 (O_2032,N_48792,N_47567);
or UO_2033 (O_2033,N_48468,N_49684);
or UO_2034 (O_2034,N_49639,N_49457);
and UO_2035 (O_2035,N_48473,N_49214);
or UO_2036 (O_2036,N_47996,N_48684);
nor UO_2037 (O_2037,N_49294,N_47856);
or UO_2038 (O_2038,N_49776,N_49756);
xor UO_2039 (O_2039,N_49039,N_49842);
xnor UO_2040 (O_2040,N_48490,N_48487);
nand UO_2041 (O_2041,N_48297,N_47825);
nand UO_2042 (O_2042,N_48292,N_47909);
and UO_2043 (O_2043,N_49315,N_48869);
and UO_2044 (O_2044,N_47559,N_47782);
nand UO_2045 (O_2045,N_48946,N_48911);
or UO_2046 (O_2046,N_48022,N_49071);
nor UO_2047 (O_2047,N_48931,N_47776);
and UO_2048 (O_2048,N_47999,N_49294);
or UO_2049 (O_2049,N_49001,N_49245);
nand UO_2050 (O_2050,N_48128,N_48164);
and UO_2051 (O_2051,N_48201,N_47870);
xor UO_2052 (O_2052,N_47546,N_49355);
xor UO_2053 (O_2053,N_47731,N_48008);
or UO_2054 (O_2054,N_48934,N_49192);
or UO_2055 (O_2055,N_47768,N_47627);
nor UO_2056 (O_2056,N_49489,N_49117);
and UO_2057 (O_2057,N_49255,N_48480);
or UO_2058 (O_2058,N_48225,N_49630);
nor UO_2059 (O_2059,N_48453,N_49214);
and UO_2060 (O_2060,N_49564,N_48031);
xnor UO_2061 (O_2061,N_48878,N_47894);
nand UO_2062 (O_2062,N_48044,N_47728);
nand UO_2063 (O_2063,N_49385,N_48295);
nor UO_2064 (O_2064,N_47529,N_49887);
or UO_2065 (O_2065,N_47668,N_47657);
nor UO_2066 (O_2066,N_49883,N_49371);
nor UO_2067 (O_2067,N_47929,N_49824);
nor UO_2068 (O_2068,N_49914,N_49423);
and UO_2069 (O_2069,N_49209,N_48150);
or UO_2070 (O_2070,N_49700,N_47721);
nor UO_2071 (O_2071,N_49132,N_49736);
nand UO_2072 (O_2072,N_49938,N_48423);
nor UO_2073 (O_2073,N_49544,N_48828);
nand UO_2074 (O_2074,N_48125,N_49492);
and UO_2075 (O_2075,N_48739,N_49989);
and UO_2076 (O_2076,N_49654,N_48866);
nand UO_2077 (O_2077,N_49923,N_49943);
nor UO_2078 (O_2078,N_48782,N_48836);
or UO_2079 (O_2079,N_49438,N_49194);
or UO_2080 (O_2080,N_49730,N_48775);
nand UO_2081 (O_2081,N_49731,N_48066);
nand UO_2082 (O_2082,N_47553,N_48544);
xor UO_2083 (O_2083,N_49054,N_48655);
or UO_2084 (O_2084,N_48522,N_48160);
xnor UO_2085 (O_2085,N_49214,N_49314);
and UO_2086 (O_2086,N_48384,N_47843);
nand UO_2087 (O_2087,N_49194,N_48591);
nand UO_2088 (O_2088,N_49256,N_49255);
or UO_2089 (O_2089,N_49623,N_49137);
xnor UO_2090 (O_2090,N_48855,N_49214);
and UO_2091 (O_2091,N_49313,N_47545);
nand UO_2092 (O_2092,N_49091,N_47992);
nor UO_2093 (O_2093,N_47611,N_48296);
nor UO_2094 (O_2094,N_49781,N_49420);
xor UO_2095 (O_2095,N_48663,N_48824);
xnor UO_2096 (O_2096,N_48514,N_48341);
or UO_2097 (O_2097,N_47518,N_48730);
xor UO_2098 (O_2098,N_48598,N_48905);
and UO_2099 (O_2099,N_48959,N_49717);
nor UO_2100 (O_2100,N_48220,N_47571);
nor UO_2101 (O_2101,N_49008,N_48064);
nor UO_2102 (O_2102,N_48154,N_49257);
or UO_2103 (O_2103,N_48440,N_49675);
nand UO_2104 (O_2104,N_49504,N_47655);
nand UO_2105 (O_2105,N_47992,N_49743);
nand UO_2106 (O_2106,N_49778,N_48142);
and UO_2107 (O_2107,N_47572,N_49559);
and UO_2108 (O_2108,N_49498,N_48510);
nand UO_2109 (O_2109,N_48086,N_48989);
nor UO_2110 (O_2110,N_49253,N_48239);
nor UO_2111 (O_2111,N_49499,N_48868);
and UO_2112 (O_2112,N_48953,N_48075);
nand UO_2113 (O_2113,N_49969,N_47602);
and UO_2114 (O_2114,N_48979,N_49125);
nor UO_2115 (O_2115,N_47525,N_48929);
nand UO_2116 (O_2116,N_49204,N_48552);
or UO_2117 (O_2117,N_49954,N_48131);
nand UO_2118 (O_2118,N_49601,N_49405);
and UO_2119 (O_2119,N_47784,N_48344);
nand UO_2120 (O_2120,N_49947,N_48933);
nor UO_2121 (O_2121,N_49766,N_48665);
and UO_2122 (O_2122,N_47692,N_47788);
nand UO_2123 (O_2123,N_49940,N_48483);
xnor UO_2124 (O_2124,N_49873,N_49324);
and UO_2125 (O_2125,N_48273,N_48326);
nand UO_2126 (O_2126,N_47820,N_49194);
nor UO_2127 (O_2127,N_48045,N_49897);
nand UO_2128 (O_2128,N_47713,N_48853);
xnor UO_2129 (O_2129,N_48533,N_48039);
nor UO_2130 (O_2130,N_47537,N_49760);
or UO_2131 (O_2131,N_47943,N_49147);
nor UO_2132 (O_2132,N_48527,N_47663);
or UO_2133 (O_2133,N_49610,N_47703);
and UO_2134 (O_2134,N_49202,N_48299);
nor UO_2135 (O_2135,N_48689,N_48303);
nand UO_2136 (O_2136,N_48748,N_49728);
or UO_2137 (O_2137,N_49791,N_47980);
nor UO_2138 (O_2138,N_49633,N_48339);
xnor UO_2139 (O_2139,N_49260,N_49780);
xor UO_2140 (O_2140,N_48583,N_48838);
or UO_2141 (O_2141,N_48921,N_47622);
xnor UO_2142 (O_2142,N_48107,N_49949);
and UO_2143 (O_2143,N_47738,N_49236);
xnor UO_2144 (O_2144,N_49680,N_49172);
nor UO_2145 (O_2145,N_49234,N_49820);
or UO_2146 (O_2146,N_48378,N_48590);
nand UO_2147 (O_2147,N_48497,N_47660);
nand UO_2148 (O_2148,N_49210,N_48526);
nand UO_2149 (O_2149,N_48439,N_47700);
and UO_2150 (O_2150,N_49267,N_49127);
and UO_2151 (O_2151,N_49322,N_49310);
and UO_2152 (O_2152,N_49772,N_47993);
nand UO_2153 (O_2153,N_49730,N_48880);
nand UO_2154 (O_2154,N_47547,N_49578);
nor UO_2155 (O_2155,N_48117,N_49469);
nor UO_2156 (O_2156,N_48896,N_48345);
nor UO_2157 (O_2157,N_47826,N_49694);
and UO_2158 (O_2158,N_49540,N_48872);
and UO_2159 (O_2159,N_48385,N_49659);
or UO_2160 (O_2160,N_49734,N_49005);
and UO_2161 (O_2161,N_49994,N_49474);
or UO_2162 (O_2162,N_49845,N_48510);
or UO_2163 (O_2163,N_49683,N_47653);
and UO_2164 (O_2164,N_48231,N_49959);
nor UO_2165 (O_2165,N_49274,N_49809);
nand UO_2166 (O_2166,N_48365,N_48271);
xnor UO_2167 (O_2167,N_49879,N_49062);
nor UO_2168 (O_2168,N_48654,N_48797);
and UO_2169 (O_2169,N_48203,N_49005);
or UO_2170 (O_2170,N_49276,N_47966);
nor UO_2171 (O_2171,N_48595,N_48976);
nand UO_2172 (O_2172,N_49405,N_49858);
and UO_2173 (O_2173,N_49347,N_49067);
xor UO_2174 (O_2174,N_48822,N_48107);
and UO_2175 (O_2175,N_49154,N_49040);
xnor UO_2176 (O_2176,N_49577,N_49982);
nor UO_2177 (O_2177,N_47569,N_47848);
or UO_2178 (O_2178,N_49145,N_49634);
nor UO_2179 (O_2179,N_48690,N_49391);
xnor UO_2180 (O_2180,N_48248,N_49634);
nor UO_2181 (O_2181,N_47659,N_49169);
and UO_2182 (O_2182,N_49536,N_48632);
nand UO_2183 (O_2183,N_49903,N_48583);
or UO_2184 (O_2184,N_49201,N_49558);
xor UO_2185 (O_2185,N_49332,N_47901);
nand UO_2186 (O_2186,N_48673,N_48913);
nand UO_2187 (O_2187,N_49725,N_49975);
or UO_2188 (O_2188,N_48129,N_49758);
and UO_2189 (O_2189,N_49407,N_48242);
xor UO_2190 (O_2190,N_48090,N_49558);
and UO_2191 (O_2191,N_48874,N_49735);
xor UO_2192 (O_2192,N_48163,N_49590);
nor UO_2193 (O_2193,N_48789,N_47717);
and UO_2194 (O_2194,N_48045,N_48109);
nand UO_2195 (O_2195,N_47808,N_48740);
xnor UO_2196 (O_2196,N_48867,N_49602);
nor UO_2197 (O_2197,N_49665,N_47844);
nor UO_2198 (O_2198,N_48703,N_48279);
xor UO_2199 (O_2199,N_48620,N_47715);
and UO_2200 (O_2200,N_48952,N_49986);
nor UO_2201 (O_2201,N_49819,N_49837);
and UO_2202 (O_2202,N_49572,N_48192);
and UO_2203 (O_2203,N_47598,N_49481);
nand UO_2204 (O_2204,N_48286,N_47611);
nand UO_2205 (O_2205,N_48647,N_49412);
nor UO_2206 (O_2206,N_49325,N_47983);
and UO_2207 (O_2207,N_47541,N_48443);
or UO_2208 (O_2208,N_49750,N_48406);
or UO_2209 (O_2209,N_49041,N_49667);
xor UO_2210 (O_2210,N_49160,N_49815);
nand UO_2211 (O_2211,N_48414,N_49937);
xor UO_2212 (O_2212,N_48493,N_49739);
or UO_2213 (O_2213,N_48509,N_48797);
xor UO_2214 (O_2214,N_49239,N_47916);
or UO_2215 (O_2215,N_49740,N_49477);
and UO_2216 (O_2216,N_49150,N_47726);
nand UO_2217 (O_2217,N_48190,N_48863);
nand UO_2218 (O_2218,N_48411,N_48857);
and UO_2219 (O_2219,N_49201,N_49917);
nor UO_2220 (O_2220,N_48916,N_49631);
nor UO_2221 (O_2221,N_49679,N_48562);
or UO_2222 (O_2222,N_49884,N_48607);
and UO_2223 (O_2223,N_49146,N_48741);
or UO_2224 (O_2224,N_49532,N_49189);
nor UO_2225 (O_2225,N_48128,N_48335);
nor UO_2226 (O_2226,N_49120,N_48768);
nand UO_2227 (O_2227,N_47590,N_48020);
nand UO_2228 (O_2228,N_48099,N_48628);
and UO_2229 (O_2229,N_47781,N_47975);
and UO_2230 (O_2230,N_48307,N_49634);
and UO_2231 (O_2231,N_47909,N_49117);
and UO_2232 (O_2232,N_49278,N_49856);
nor UO_2233 (O_2233,N_49285,N_49912);
nor UO_2234 (O_2234,N_47643,N_49594);
and UO_2235 (O_2235,N_47801,N_49736);
xor UO_2236 (O_2236,N_47902,N_49311);
or UO_2237 (O_2237,N_49236,N_49876);
xnor UO_2238 (O_2238,N_49833,N_48784);
and UO_2239 (O_2239,N_48461,N_48970);
xor UO_2240 (O_2240,N_49660,N_49722);
xor UO_2241 (O_2241,N_47851,N_49762);
or UO_2242 (O_2242,N_49701,N_49792);
xnor UO_2243 (O_2243,N_48680,N_48891);
nand UO_2244 (O_2244,N_48816,N_48578);
xor UO_2245 (O_2245,N_48739,N_49965);
nor UO_2246 (O_2246,N_48013,N_47612);
xor UO_2247 (O_2247,N_49987,N_49455);
and UO_2248 (O_2248,N_49687,N_47555);
and UO_2249 (O_2249,N_48983,N_48090);
or UO_2250 (O_2250,N_49520,N_48384);
and UO_2251 (O_2251,N_49606,N_48957);
nand UO_2252 (O_2252,N_47876,N_48328);
nor UO_2253 (O_2253,N_48179,N_48056);
and UO_2254 (O_2254,N_49276,N_49645);
nor UO_2255 (O_2255,N_48367,N_48356);
and UO_2256 (O_2256,N_49380,N_48858);
or UO_2257 (O_2257,N_48969,N_49346);
xnor UO_2258 (O_2258,N_48777,N_49198);
or UO_2259 (O_2259,N_47814,N_49870);
nand UO_2260 (O_2260,N_48814,N_48442);
nand UO_2261 (O_2261,N_49781,N_48634);
or UO_2262 (O_2262,N_48445,N_49297);
nand UO_2263 (O_2263,N_47815,N_47979);
and UO_2264 (O_2264,N_49869,N_49055);
and UO_2265 (O_2265,N_48170,N_48436);
or UO_2266 (O_2266,N_48292,N_47517);
or UO_2267 (O_2267,N_49835,N_49848);
and UO_2268 (O_2268,N_49264,N_48639);
xor UO_2269 (O_2269,N_49013,N_48181);
nand UO_2270 (O_2270,N_49260,N_49585);
xor UO_2271 (O_2271,N_49705,N_49728);
and UO_2272 (O_2272,N_49713,N_48624);
and UO_2273 (O_2273,N_48392,N_49097);
nand UO_2274 (O_2274,N_49102,N_47640);
xnor UO_2275 (O_2275,N_49599,N_49612);
or UO_2276 (O_2276,N_47865,N_48922);
or UO_2277 (O_2277,N_48455,N_48497);
xor UO_2278 (O_2278,N_49629,N_48739);
nand UO_2279 (O_2279,N_48448,N_48222);
or UO_2280 (O_2280,N_48860,N_49140);
and UO_2281 (O_2281,N_48919,N_48570);
xor UO_2282 (O_2282,N_48407,N_48616);
or UO_2283 (O_2283,N_47759,N_48192);
or UO_2284 (O_2284,N_48759,N_48539);
and UO_2285 (O_2285,N_48351,N_49972);
nor UO_2286 (O_2286,N_47769,N_48627);
xnor UO_2287 (O_2287,N_49513,N_48545);
nand UO_2288 (O_2288,N_48721,N_48464);
xnor UO_2289 (O_2289,N_49605,N_48355);
and UO_2290 (O_2290,N_47648,N_48666);
nor UO_2291 (O_2291,N_47509,N_49017);
and UO_2292 (O_2292,N_49804,N_49718);
or UO_2293 (O_2293,N_48997,N_48793);
or UO_2294 (O_2294,N_49398,N_49228);
or UO_2295 (O_2295,N_48242,N_47922);
or UO_2296 (O_2296,N_49114,N_47843);
xnor UO_2297 (O_2297,N_49068,N_49410);
xnor UO_2298 (O_2298,N_48104,N_48511);
nor UO_2299 (O_2299,N_48535,N_49161);
nor UO_2300 (O_2300,N_48986,N_49477);
xor UO_2301 (O_2301,N_48362,N_49183);
xor UO_2302 (O_2302,N_48790,N_48482);
and UO_2303 (O_2303,N_49947,N_47666);
xor UO_2304 (O_2304,N_49533,N_49293);
nand UO_2305 (O_2305,N_48264,N_48617);
xnor UO_2306 (O_2306,N_49465,N_47764);
and UO_2307 (O_2307,N_48576,N_48175);
xnor UO_2308 (O_2308,N_49667,N_49882);
nor UO_2309 (O_2309,N_47811,N_48292);
or UO_2310 (O_2310,N_49082,N_47690);
nand UO_2311 (O_2311,N_48003,N_48923);
or UO_2312 (O_2312,N_48732,N_48710);
and UO_2313 (O_2313,N_48713,N_49479);
nand UO_2314 (O_2314,N_49401,N_48623);
nor UO_2315 (O_2315,N_49322,N_48838);
xor UO_2316 (O_2316,N_49641,N_48156);
and UO_2317 (O_2317,N_47551,N_48437);
nor UO_2318 (O_2318,N_48541,N_49986);
nor UO_2319 (O_2319,N_48294,N_48345);
nand UO_2320 (O_2320,N_48373,N_48647);
nand UO_2321 (O_2321,N_48732,N_49875);
nor UO_2322 (O_2322,N_48302,N_47753);
and UO_2323 (O_2323,N_48863,N_49146);
nor UO_2324 (O_2324,N_49636,N_47886);
nand UO_2325 (O_2325,N_48069,N_48022);
nor UO_2326 (O_2326,N_48421,N_49512);
and UO_2327 (O_2327,N_49173,N_47878);
and UO_2328 (O_2328,N_49086,N_49036);
xor UO_2329 (O_2329,N_48564,N_49068);
and UO_2330 (O_2330,N_49874,N_47621);
nand UO_2331 (O_2331,N_48419,N_47737);
nand UO_2332 (O_2332,N_49495,N_49059);
nor UO_2333 (O_2333,N_48959,N_49992);
and UO_2334 (O_2334,N_49838,N_49335);
and UO_2335 (O_2335,N_49698,N_49986);
and UO_2336 (O_2336,N_49638,N_48218);
nand UO_2337 (O_2337,N_47758,N_48383);
nor UO_2338 (O_2338,N_48570,N_49072);
xor UO_2339 (O_2339,N_48516,N_48549);
nor UO_2340 (O_2340,N_49697,N_48898);
or UO_2341 (O_2341,N_48398,N_49921);
and UO_2342 (O_2342,N_49020,N_48976);
or UO_2343 (O_2343,N_48760,N_49424);
nand UO_2344 (O_2344,N_48879,N_48972);
or UO_2345 (O_2345,N_48143,N_48051);
xnor UO_2346 (O_2346,N_49608,N_49516);
and UO_2347 (O_2347,N_49150,N_47738);
nor UO_2348 (O_2348,N_49323,N_47996);
or UO_2349 (O_2349,N_48304,N_49915);
and UO_2350 (O_2350,N_48998,N_49285);
or UO_2351 (O_2351,N_47887,N_48350);
nor UO_2352 (O_2352,N_48142,N_48694);
xor UO_2353 (O_2353,N_49128,N_48919);
xnor UO_2354 (O_2354,N_47657,N_49744);
nor UO_2355 (O_2355,N_48261,N_49481);
nand UO_2356 (O_2356,N_49080,N_49304);
nor UO_2357 (O_2357,N_49097,N_48725);
or UO_2358 (O_2358,N_49843,N_49297);
and UO_2359 (O_2359,N_48005,N_47674);
xnor UO_2360 (O_2360,N_47720,N_48154);
xor UO_2361 (O_2361,N_49399,N_47656);
or UO_2362 (O_2362,N_49689,N_49383);
nand UO_2363 (O_2363,N_48095,N_48446);
nand UO_2364 (O_2364,N_48339,N_48119);
nand UO_2365 (O_2365,N_48430,N_48982);
nand UO_2366 (O_2366,N_49144,N_49087);
nand UO_2367 (O_2367,N_48056,N_49309);
xnor UO_2368 (O_2368,N_48411,N_47744);
nor UO_2369 (O_2369,N_48986,N_49970);
or UO_2370 (O_2370,N_47911,N_48079);
and UO_2371 (O_2371,N_48177,N_49488);
nor UO_2372 (O_2372,N_49337,N_47572);
and UO_2373 (O_2373,N_48911,N_49329);
nor UO_2374 (O_2374,N_49443,N_49296);
or UO_2375 (O_2375,N_48481,N_48504);
and UO_2376 (O_2376,N_49302,N_47567);
xor UO_2377 (O_2377,N_49742,N_47701);
nand UO_2378 (O_2378,N_49205,N_49806);
and UO_2379 (O_2379,N_49862,N_49027);
or UO_2380 (O_2380,N_49907,N_49091);
nor UO_2381 (O_2381,N_49515,N_47517);
nor UO_2382 (O_2382,N_49583,N_47518);
and UO_2383 (O_2383,N_47768,N_48602);
nand UO_2384 (O_2384,N_48226,N_48315);
nor UO_2385 (O_2385,N_47639,N_47952);
and UO_2386 (O_2386,N_49155,N_49311);
or UO_2387 (O_2387,N_47859,N_48038);
nand UO_2388 (O_2388,N_48984,N_49567);
nand UO_2389 (O_2389,N_48568,N_48784);
and UO_2390 (O_2390,N_48991,N_49641);
and UO_2391 (O_2391,N_49534,N_48454);
nor UO_2392 (O_2392,N_47731,N_48172);
nor UO_2393 (O_2393,N_48308,N_47860);
or UO_2394 (O_2394,N_47813,N_49120);
xor UO_2395 (O_2395,N_48090,N_49313);
nor UO_2396 (O_2396,N_49191,N_49965);
and UO_2397 (O_2397,N_49894,N_49279);
xnor UO_2398 (O_2398,N_48216,N_48287);
or UO_2399 (O_2399,N_48085,N_48028);
or UO_2400 (O_2400,N_49930,N_47597);
xnor UO_2401 (O_2401,N_48644,N_48986);
nand UO_2402 (O_2402,N_48112,N_48353);
nor UO_2403 (O_2403,N_48695,N_47613);
xnor UO_2404 (O_2404,N_48968,N_49780);
nand UO_2405 (O_2405,N_49856,N_49404);
and UO_2406 (O_2406,N_49021,N_47927);
nor UO_2407 (O_2407,N_47578,N_48171);
nand UO_2408 (O_2408,N_48820,N_48257);
nand UO_2409 (O_2409,N_49093,N_47656);
nand UO_2410 (O_2410,N_49199,N_48053);
xnor UO_2411 (O_2411,N_49893,N_49460);
nand UO_2412 (O_2412,N_49755,N_49837);
or UO_2413 (O_2413,N_47938,N_47548);
or UO_2414 (O_2414,N_48055,N_49707);
nand UO_2415 (O_2415,N_49401,N_49981);
and UO_2416 (O_2416,N_49721,N_49686);
and UO_2417 (O_2417,N_47737,N_49671);
or UO_2418 (O_2418,N_49206,N_48027);
nand UO_2419 (O_2419,N_48727,N_47877);
or UO_2420 (O_2420,N_48580,N_49370);
or UO_2421 (O_2421,N_48467,N_49019);
nand UO_2422 (O_2422,N_48974,N_47936);
nor UO_2423 (O_2423,N_48269,N_48035);
nand UO_2424 (O_2424,N_49034,N_48746);
xor UO_2425 (O_2425,N_49540,N_48817);
or UO_2426 (O_2426,N_48095,N_49875);
or UO_2427 (O_2427,N_49455,N_49048);
xnor UO_2428 (O_2428,N_48426,N_49570);
xnor UO_2429 (O_2429,N_48062,N_48363);
and UO_2430 (O_2430,N_48720,N_48103);
and UO_2431 (O_2431,N_49248,N_49112);
nand UO_2432 (O_2432,N_47794,N_49360);
nor UO_2433 (O_2433,N_48281,N_47617);
nand UO_2434 (O_2434,N_48053,N_49899);
xor UO_2435 (O_2435,N_47909,N_49654);
nor UO_2436 (O_2436,N_49668,N_47766);
or UO_2437 (O_2437,N_49572,N_49432);
nand UO_2438 (O_2438,N_47671,N_48553);
and UO_2439 (O_2439,N_47728,N_48411);
or UO_2440 (O_2440,N_48068,N_48278);
xnor UO_2441 (O_2441,N_48774,N_47543);
xnor UO_2442 (O_2442,N_49852,N_49626);
and UO_2443 (O_2443,N_49350,N_48737);
nand UO_2444 (O_2444,N_49768,N_49161);
xor UO_2445 (O_2445,N_48583,N_48313);
nand UO_2446 (O_2446,N_48450,N_49436);
nand UO_2447 (O_2447,N_48360,N_48031);
nor UO_2448 (O_2448,N_49735,N_47925);
or UO_2449 (O_2449,N_48595,N_49749);
nor UO_2450 (O_2450,N_49878,N_49911);
nand UO_2451 (O_2451,N_49617,N_48940);
nor UO_2452 (O_2452,N_49503,N_49430);
or UO_2453 (O_2453,N_48886,N_49297);
or UO_2454 (O_2454,N_49884,N_47916);
nand UO_2455 (O_2455,N_49764,N_47551);
or UO_2456 (O_2456,N_48048,N_47873);
nor UO_2457 (O_2457,N_48685,N_48402);
or UO_2458 (O_2458,N_49696,N_49189);
nand UO_2459 (O_2459,N_49803,N_48301);
nand UO_2460 (O_2460,N_49016,N_47855);
and UO_2461 (O_2461,N_48828,N_48978);
nand UO_2462 (O_2462,N_49901,N_47772);
and UO_2463 (O_2463,N_48302,N_48544);
and UO_2464 (O_2464,N_47993,N_49561);
and UO_2465 (O_2465,N_49056,N_48817);
and UO_2466 (O_2466,N_47632,N_48638);
nand UO_2467 (O_2467,N_49679,N_47521);
nand UO_2468 (O_2468,N_47631,N_47877);
xor UO_2469 (O_2469,N_48948,N_48237);
xor UO_2470 (O_2470,N_49737,N_49256);
nor UO_2471 (O_2471,N_48430,N_48095);
nand UO_2472 (O_2472,N_49529,N_47627);
xnor UO_2473 (O_2473,N_47515,N_47583);
and UO_2474 (O_2474,N_49081,N_48594);
nand UO_2475 (O_2475,N_49525,N_48387);
nand UO_2476 (O_2476,N_47685,N_49533);
xor UO_2477 (O_2477,N_48179,N_47812);
nand UO_2478 (O_2478,N_49316,N_49527);
nand UO_2479 (O_2479,N_49282,N_48707);
and UO_2480 (O_2480,N_48996,N_48654);
nand UO_2481 (O_2481,N_47736,N_49924);
and UO_2482 (O_2482,N_48117,N_47707);
nand UO_2483 (O_2483,N_48365,N_48471);
and UO_2484 (O_2484,N_49111,N_49042);
nor UO_2485 (O_2485,N_47778,N_48347);
nand UO_2486 (O_2486,N_48632,N_48938);
nor UO_2487 (O_2487,N_48292,N_47960);
nand UO_2488 (O_2488,N_48436,N_49527);
nor UO_2489 (O_2489,N_49828,N_48407);
nand UO_2490 (O_2490,N_49947,N_49007);
xnor UO_2491 (O_2491,N_48901,N_48502);
or UO_2492 (O_2492,N_49857,N_47789);
nand UO_2493 (O_2493,N_49875,N_48202);
nand UO_2494 (O_2494,N_47901,N_47529);
nand UO_2495 (O_2495,N_48444,N_48946);
and UO_2496 (O_2496,N_49504,N_49350);
nand UO_2497 (O_2497,N_48470,N_47588);
and UO_2498 (O_2498,N_49066,N_48248);
and UO_2499 (O_2499,N_48908,N_47543);
nor UO_2500 (O_2500,N_48480,N_47851);
xor UO_2501 (O_2501,N_49867,N_48790);
nor UO_2502 (O_2502,N_48965,N_48827);
xor UO_2503 (O_2503,N_49553,N_49846);
xor UO_2504 (O_2504,N_48924,N_49774);
xnor UO_2505 (O_2505,N_47852,N_48985);
xnor UO_2506 (O_2506,N_49972,N_49391);
or UO_2507 (O_2507,N_48639,N_49504);
or UO_2508 (O_2508,N_48976,N_49401);
or UO_2509 (O_2509,N_48568,N_49726);
nand UO_2510 (O_2510,N_49656,N_47867);
or UO_2511 (O_2511,N_48193,N_49479);
nand UO_2512 (O_2512,N_49036,N_49459);
and UO_2513 (O_2513,N_47595,N_47601);
or UO_2514 (O_2514,N_48044,N_47987);
nand UO_2515 (O_2515,N_49056,N_49872);
and UO_2516 (O_2516,N_49104,N_48029);
nand UO_2517 (O_2517,N_48365,N_49069);
nor UO_2518 (O_2518,N_49840,N_47784);
xnor UO_2519 (O_2519,N_48115,N_49870);
xor UO_2520 (O_2520,N_49508,N_49969);
and UO_2521 (O_2521,N_48023,N_48204);
xor UO_2522 (O_2522,N_49178,N_48526);
or UO_2523 (O_2523,N_48434,N_47934);
or UO_2524 (O_2524,N_49487,N_47910);
and UO_2525 (O_2525,N_48785,N_48717);
nor UO_2526 (O_2526,N_48694,N_48031);
xnor UO_2527 (O_2527,N_48309,N_49032);
nand UO_2528 (O_2528,N_49800,N_48416);
nor UO_2529 (O_2529,N_48927,N_49403);
xor UO_2530 (O_2530,N_49686,N_49429);
or UO_2531 (O_2531,N_47641,N_49864);
and UO_2532 (O_2532,N_49578,N_49367);
nand UO_2533 (O_2533,N_49674,N_48814);
and UO_2534 (O_2534,N_47638,N_47570);
xor UO_2535 (O_2535,N_48903,N_48119);
and UO_2536 (O_2536,N_48880,N_48111);
or UO_2537 (O_2537,N_49720,N_47620);
nand UO_2538 (O_2538,N_49528,N_48561);
nand UO_2539 (O_2539,N_47774,N_49770);
nand UO_2540 (O_2540,N_47720,N_47822);
nand UO_2541 (O_2541,N_49778,N_49420);
and UO_2542 (O_2542,N_48230,N_49487);
nor UO_2543 (O_2543,N_49285,N_48485);
xor UO_2544 (O_2544,N_48575,N_47811);
nor UO_2545 (O_2545,N_47803,N_49080);
or UO_2546 (O_2546,N_49323,N_47596);
or UO_2547 (O_2547,N_49560,N_49862);
nor UO_2548 (O_2548,N_48830,N_48166);
xor UO_2549 (O_2549,N_49360,N_48151);
nand UO_2550 (O_2550,N_48611,N_47950);
and UO_2551 (O_2551,N_47837,N_49116);
nand UO_2552 (O_2552,N_47662,N_49182);
nor UO_2553 (O_2553,N_49962,N_48614);
nand UO_2554 (O_2554,N_48473,N_49536);
and UO_2555 (O_2555,N_48499,N_47518);
xnor UO_2556 (O_2556,N_49091,N_48239);
xnor UO_2557 (O_2557,N_48203,N_47522);
nor UO_2558 (O_2558,N_49783,N_49203);
or UO_2559 (O_2559,N_48558,N_48992);
or UO_2560 (O_2560,N_49891,N_49953);
nor UO_2561 (O_2561,N_48296,N_48496);
and UO_2562 (O_2562,N_48838,N_48219);
nand UO_2563 (O_2563,N_48611,N_48256);
and UO_2564 (O_2564,N_48095,N_47772);
or UO_2565 (O_2565,N_48376,N_49973);
or UO_2566 (O_2566,N_47572,N_48113);
and UO_2567 (O_2567,N_49250,N_47938);
and UO_2568 (O_2568,N_49245,N_49815);
nand UO_2569 (O_2569,N_48869,N_47506);
and UO_2570 (O_2570,N_49534,N_47500);
xnor UO_2571 (O_2571,N_48491,N_48537);
or UO_2572 (O_2572,N_49701,N_49362);
xnor UO_2573 (O_2573,N_49465,N_49414);
nor UO_2574 (O_2574,N_48852,N_48951);
and UO_2575 (O_2575,N_49391,N_48620);
nor UO_2576 (O_2576,N_49375,N_49496);
or UO_2577 (O_2577,N_48173,N_49506);
and UO_2578 (O_2578,N_49640,N_48872);
and UO_2579 (O_2579,N_48354,N_48444);
nand UO_2580 (O_2580,N_49465,N_48189);
xnor UO_2581 (O_2581,N_49851,N_49611);
or UO_2582 (O_2582,N_49086,N_49504);
nand UO_2583 (O_2583,N_48691,N_47704);
and UO_2584 (O_2584,N_47975,N_48716);
and UO_2585 (O_2585,N_48166,N_48218);
nor UO_2586 (O_2586,N_48022,N_49429);
nand UO_2587 (O_2587,N_48372,N_49320);
and UO_2588 (O_2588,N_48129,N_47930);
nor UO_2589 (O_2589,N_48920,N_48028);
or UO_2590 (O_2590,N_49126,N_47957);
xor UO_2591 (O_2591,N_48198,N_48460);
and UO_2592 (O_2592,N_49167,N_49394);
and UO_2593 (O_2593,N_48544,N_47732);
and UO_2594 (O_2594,N_49852,N_48905);
or UO_2595 (O_2595,N_48732,N_49026);
nand UO_2596 (O_2596,N_49927,N_48465);
xor UO_2597 (O_2597,N_47962,N_48283);
nor UO_2598 (O_2598,N_49163,N_48268);
nand UO_2599 (O_2599,N_49428,N_48127);
and UO_2600 (O_2600,N_47866,N_49630);
nor UO_2601 (O_2601,N_48999,N_48543);
or UO_2602 (O_2602,N_49046,N_47609);
and UO_2603 (O_2603,N_49780,N_47844);
or UO_2604 (O_2604,N_49344,N_48325);
nand UO_2605 (O_2605,N_49191,N_49851);
nor UO_2606 (O_2606,N_49930,N_49834);
and UO_2607 (O_2607,N_47955,N_48005);
and UO_2608 (O_2608,N_48590,N_49191);
xor UO_2609 (O_2609,N_48652,N_49545);
or UO_2610 (O_2610,N_47668,N_48741);
nor UO_2611 (O_2611,N_47814,N_47790);
and UO_2612 (O_2612,N_48005,N_47654);
or UO_2613 (O_2613,N_48924,N_48803);
nand UO_2614 (O_2614,N_48041,N_48495);
nor UO_2615 (O_2615,N_49429,N_48012);
and UO_2616 (O_2616,N_49756,N_49967);
or UO_2617 (O_2617,N_48053,N_49175);
nor UO_2618 (O_2618,N_48144,N_48162);
or UO_2619 (O_2619,N_48415,N_47714);
nand UO_2620 (O_2620,N_47598,N_49059);
and UO_2621 (O_2621,N_49650,N_47567);
and UO_2622 (O_2622,N_47550,N_49032);
nand UO_2623 (O_2623,N_49001,N_48161);
xor UO_2624 (O_2624,N_49055,N_48937);
nand UO_2625 (O_2625,N_48211,N_49854);
or UO_2626 (O_2626,N_49278,N_48960);
or UO_2627 (O_2627,N_48047,N_49601);
nand UO_2628 (O_2628,N_47595,N_47549);
xor UO_2629 (O_2629,N_48549,N_48683);
xor UO_2630 (O_2630,N_48469,N_48608);
and UO_2631 (O_2631,N_47758,N_47674);
xor UO_2632 (O_2632,N_48645,N_48524);
or UO_2633 (O_2633,N_48858,N_48695);
nor UO_2634 (O_2634,N_49068,N_49964);
nand UO_2635 (O_2635,N_49819,N_48178);
and UO_2636 (O_2636,N_47796,N_48324);
xor UO_2637 (O_2637,N_48525,N_47812);
and UO_2638 (O_2638,N_49149,N_48516);
and UO_2639 (O_2639,N_49821,N_47772);
nor UO_2640 (O_2640,N_48081,N_48007);
nand UO_2641 (O_2641,N_48513,N_48091);
or UO_2642 (O_2642,N_47638,N_49608);
xor UO_2643 (O_2643,N_47568,N_48966);
xnor UO_2644 (O_2644,N_47851,N_48158);
xnor UO_2645 (O_2645,N_48503,N_47518);
nor UO_2646 (O_2646,N_48907,N_49552);
or UO_2647 (O_2647,N_49715,N_49347);
nand UO_2648 (O_2648,N_48710,N_49700);
nor UO_2649 (O_2649,N_49233,N_48847);
and UO_2650 (O_2650,N_49332,N_48480);
nand UO_2651 (O_2651,N_48272,N_48422);
nand UO_2652 (O_2652,N_49088,N_47750);
and UO_2653 (O_2653,N_47732,N_48553);
nor UO_2654 (O_2654,N_48195,N_49014);
or UO_2655 (O_2655,N_48823,N_47660);
nand UO_2656 (O_2656,N_48649,N_49701);
nand UO_2657 (O_2657,N_49052,N_49428);
nand UO_2658 (O_2658,N_49177,N_48784);
xor UO_2659 (O_2659,N_48621,N_48823);
or UO_2660 (O_2660,N_49392,N_48098);
nor UO_2661 (O_2661,N_48796,N_49077);
or UO_2662 (O_2662,N_49056,N_48806);
nand UO_2663 (O_2663,N_48188,N_47823);
or UO_2664 (O_2664,N_49883,N_48102);
xnor UO_2665 (O_2665,N_49306,N_48002);
nand UO_2666 (O_2666,N_49074,N_49308);
and UO_2667 (O_2667,N_47689,N_48286);
and UO_2668 (O_2668,N_49858,N_48872);
and UO_2669 (O_2669,N_47705,N_48869);
nand UO_2670 (O_2670,N_49753,N_48335);
and UO_2671 (O_2671,N_49903,N_48566);
nor UO_2672 (O_2672,N_48183,N_49665);
nor UO_2673 (O_2673,N_48432,N_49049);
and UO_2674 (O_2674,N_48970,N_47656);
and UO_2675 (O_2675,N_48913,N_47725);
and UO_2676 (O_2676,N_48953,N_48574);
nand UO_2677 (O_2677,N_49696,N_48631);
xnor UO_2678 (O_2678,N_48280,N_47512);
xor UO_2679 (O_2679,N_48415,N_49479);
nor UO_2680 (O_2680,N_48898,N_49249);
xnor UO_2681 (O_2681,N_48094,N_48445);
xnor UO_2682 (O_2682,N_48286,N_49818);
xnor UO_2683 (O_2683,N_47559,N_48719);
and UO_2684 (O_2684,N_49882,N_47738);
nor UO_2685 (O_2685,N_48146,N_48098);
xor UO_2686 (O_2686,N_48498,N_47606);
nor UO_2687 (O_2687,N_49755,N_49750);
nand UO_2688 (O_2688,N_48252,N_49781);
and UO_2689 (O_2689,N_47973,N_48446);
nand UO_2690 (O_2690,N_47663,N_47875);
xor UO_2691 (O_2691,N_48365,N_47570);
and UO_2692 (O_2692,N_49060,N_48317);
and UO_2693 (O_2693,N_48240,N_47882);
or UO_2694 (O_2694,N_49063,N_47675);
xor UO_2695 (O_2695,N_48416,N_48752);
and UO_2696 (O_2696,N_48713,N_47561);
or UO_2697 (O_2697,N_47541,N_47948);
and UO_2698 (O_2698,N_47573,N_48540);
or UO_2699 (O_2699,N_47926,N_49378);
xnor UO_2700 (O_2700,N_48184,N_49485);
or UO_2701 (O_2701,N_48081,N_48991);
or UO_2702 (O_2702,N_49618,N_48042);
nand UO_2703 (O_2703,N_49683,N_48101);
or UO_2704 (O_2704,N_49774,N_47746);
and UO_2705 (O_2705,N_49539,N_49101);
nand UO_2706 (O_2706,N_48343,N_48116);
nor UO_2707 (O_2707,N_49808,N_47742);
nor UO_2708 (O_2708,N_48151,N_49981);
nor UO_2709 (O_2709,N_47969,N_47740);
nor UO_2710 (O_2710,N_49042,N_47646);
nor UO_2711 (O_2711,N_49767,N_49157);
or UO_2712 (O_2712,N_49900,N_48931);
nor UO_2713 (O_2713,N_48256,N_49423);
xnor UO_2714 (O_2714,N_48428,N_49103);
nand UO_2715 (O_2715,N_49322,N_48129);
xnor UO_2716 (O_2716,N_48824,N_48650);
or UO_2717 (O_2717,N_49696,N_49377);
or UO_2718 (O_2718,N_47751,N_47988);
xnor UO_2719 (O_2719,N_49947,N_49051);
and UO_2720 (O_2720,N_49100,N_49146);
and UO_2721 (O_2721,N_48914,N_48790);
or UO_2722 (O_2722,N_48874,N_49349);
xor UO_2723 (O_2723,N_48614,N_48111);
and UO_2724 (O_2724,N_49809,N_49950);
and UO_2725 (O_2725,N_48865,N_48995);
xor UO_2726 (O_2726,N_48656,N_49973);
nand UO_2727 (O_2727,N_49320,N_49425);
nor UO_2728 (O_2728,N_48411,N_49022);
and UO_2729 (O_2729,N_48346,N_49115);
and UO_2730 (O_2730,N_47833,N_48864);
nand UO_2731 (O_2731,N_48379,N_49366);
or UO_2732 (O_2732,N_48853,N_49116);
or UO_2733 (O_2733,N_47748,N_48124);
and UO_2734 (O_2734,N_47898,N_49199);
nor UO_2735 (O_2735,N_49312,N_49284);
xor UO_2736 (O_2736,N_48697,N_48677);
or UO_2737 (O_2737,N_49450,N_49531);
or UO_2738 (O_2738,N_48782,N_48676);
or UO_2739 (O_2739,N_47638,N_48558);
nor UO_2740 (O_2740,N_48956,N_49892);
and UO_2741 (O_2741,N_47916,N_48839);
or UO_2742 (O_2742,N_49328,N_48348);
or UO_2743 (O_2743,N_48095,N_48306);
nor UO_2744 (O_2744,N_49809,N_48626);
and UO_2745 (O_2745,N_48788,N_49980);
or UO_2746 (O_2746,N_49028,N_48859);
and UO_2747 (O_2747,N_49432,N_49189);
and UO_2748 (O_2748,N_47723,N_47858);
nor UO_2749 (O_2749,N_48508,N_49354);
nor UO_2750 (O_2750,N_49578,N_49866);
xnor UO_2751 (O_2751,N_48719,N_49222);
nor UO_2752 (O_2752,N_48815,N_48916);
or UO_2753 (O_2753,N_48274,N_49064);
nand UO_2754 (O_2754,N_48701,N_48965);
and UO_2755 (O_2755,N_49405,N_48763);
xnor UO_2756 (O_2756,N_49945,N_47636);
nand UO_2757 (O_2757,N_47575,N_49450);
xnor UO_2758 (O_2758,N_48527,N_49698);
or UO_2759 (O_2759,N_47908,N_49835);
nor UO_2760 (O_2760,N_47955,N_48093);
and UO_2761 (O_2761,N_48217,N_47704);
or UO_2762 (O_2762,N_47908,N_47885);
nor UO_2763 (O_2763,N_49488,N_49727);
nor UO_2764 (O_2764,N_48466,N_48752);
xnor UO_2765 (O_2765,N_47897,N_49414);
or UO_2766 (O_2766,N_49553,N_49435);
and UO_2767 (O_2767,N_49792,N_49804);
xor UO_2768 (O_2768,N_47890,N_48483);
or UO_2769 (O_2769,N_48531,N_49989);
nand UO_2770 (O_2770,N_49105,N_48597);
xnor UO_2771 (O_2771,N_47777,N_49309);
or UO_2772 (O_2772,N_48499,N_48107);
nor UO_2773 (O_2773,N_48939,N_48924);
nand UO_2774 (O_2774,N_49708,N_48396);
and UO_2775 (O_2775,N_49489,N_48319);
and UO_2776 (O_2776,N_48279,N_49221);
xor UO_2777 (O_2777,N_48258,N_49977);
xor UO_2778 (O_2778,N_48779,N_48949);
nand UO_2779 (O_2779,N_49715,N_48994);
and UO_2780 (O_2780,N_49130,N_48619);
xor UO_2781 (O_2781,N_49707,N_47999);
nand UO_2782 (O_2782,N_49084,N_49355);
xor UO_2783 (O_2783,N_47927,N_49560);
nor UO_2784 (O_2784,N_48329,N_48867);
and UO_2785 (O_2785,N_49442,N_47532);
or UO_2786 (O_2786,N_48882,N_48293);
nand UO_2787 (O_2787,N_49750,N_47797);
nor UO_2788 (O_2788,N_47660,N_49238);
xnor UO_2789 (O_2789,N_47907,N_49226);
nor UO_2790 (O_2790,N_48584,N_49415);
and UO_2791 (O_2791,N_49957,N_48102);
xnor UO_2792 (O_2792,N_47570,N_47963);
or UO_2793 (O_2793,N_49292,N_47728);
xor UO_2794 (O_2794,N_49086,N_49368);
nand UO_2795 (O_2795,N_49457,N_48840);
xor UO_2796 (O_2796,N_47630,N_47896);
and UO_2797 (O_2797,N_47988,N_49113);
xnor UO_2798 (O_2798,N_49937,N_49566);
or UO_2799 (O_2799,N_48299,N_49313);
xnor UO_2800 (O_2800,N_49965,N_48004);
and UO_2801 (O_2801,N_49392,N_48689);
nand UO_2802 (O_2802,N_48647,N_49344);
and UO_2803 (O_2803,N_49599,N_49746);
or UO_2804 (O_2804,N_49990,N_48104);
nor UO_2805 (O_2805,N_48038,N_49881);
nor UO_2806 (O_2806,N_47667,N_48919);
and UO_2807 (O_2807,N_47602,N_49277);
xnor UO_2808 (O_2808,N_48773,N_48496);
nand UO_2809 (O_2809,N_47931,N_49043);
xor UO_2810 (O_2810,N_49885,N_49211);
and UO_2811 (O_2811,N_48478,N_47874);
nor UO_2812 (O_2812,N_48707,N_47909);
and UO_2813 (O_2813,N_48564,N_49688);
nand UO_2814 (O_2814,N_47685,N_48265);
and UO_2815 (O_2815,N_48624,N_48517);
and UO_2816 (O_2816,N_48191,N_48454);
or UO_2817 (O_2817,N_49860,N_48114);
nand UO_2818 (O_2818,N_48619,N_48082);
nor UO_2819 (O_2819,N_47608,N_49113);
nand UO_2820 (O_2820,N_48557,N_49824);
xnor UO_2821 (O_2821,N_48875,N_48826);
nor UO_2822 (O_2822,N_48104,N_48457);
or UO_2823 (O_2823,N_49671,N_48870);
nand UO_2824 (O_2824,N_47891,N_49237);
nor UO_2825 (O_2825,N_48401,N_48522);
nor UO_2826 (O_2826,N_48419,N_47838);
or UO_2827 (O_2827,N_47892,N_49445);
or UO_2828 (O_2828,N_48780,N_47840);
nand UO_2829 (O_2829,N_49314,N_48705);
nand UO_2830 (O_2830,N_48380,N_49936);
nand UO_2831 (O_2831,N_49529,N_48126);
xnor UO_2832 (O_2832,N_48731,N_48359);
nor UO_2833 (O_2833,N_48944,N_47737);
nand UO_2834 (O_2834,N_48551,N_48521);
and UO_2835 (O_2835,N_48965,N_48586);
xnor UO_2836 (O_2836,N_49487,N_49214);
and UO_2837 (O_2837,N_49051,N_48974);
nand UO_2838 (O_2838,N_47912,N_47614);
xnor UO_2839 (O_2839,N_47868,N_49791);
or UO_2840 (O_2840,N_48207,N_49631);
xor UO_2841 (O_2841,N_48512,N_49351);
or UO_2842 (O_2842,N_48104,N_47501);
and UO_2843 (O_2843,N_47779,N_48321);
xor UO_2844 (O_2844,N_48627,N_47735);
and UO_2845 (O_2845,N_49511,N_49789);
or UO_2846 (O_2846,N_49462,N_47572);
nor UO_2847 (O_2847,N_48957,N_49302);
and UO_2848 (O_2848,N_49153,N_48217);
or UO_2849 (O_2849,N_49350,N_47529);
or UO_2850 (O_2850,N_48195,N_48774);
nor UO_2851 (O_2851,N_49832,N_49166);
or UO_2852 (O_2852,N_49800,N_48484);
nor UO_2853 (O_2853,N_47950,N_49482);
nor UO_2854 (O_2854,N_48102,N_49654);
xor UO_2855 (O_2855,N_49301,N_49073);
nor UO_2856 (O_2856,N_48000,N_49586);
nand UO_2857 (O_2857,N_47824,N_48255);
xnor UO_2858 (O_2858,N_47514,N_48249);
and UO_2859 (O_2859,N_49401,N_49265);
and UO_2860 (O_2860,N_49020,N_47967);
nand UO_2861 (O_2861,N_48523,N_47874);
xor UO_2862 (O_2862,N_49462,N_48122);
nor UO_2863 (O_2863,N_48799,N_49609);
nor UO_2864 (O_2864,N_48885,N_49329);
nor UO_2865 (O_2865,N_49038,N_47972);
xnor UO_2866 (O_2866,N_49888,N_48544);
nand UO_2867 (O_2867,N_49379,N_48496);
nand UO_2868 (O_2868,N_49185,N_49304);
or UO_2869 (O_2869,N_48265,N_49491);
nand UO_2870 (O_2870,N_49994,N_49611);
and UO_2871 (O_2871,N_48763,N_49650);
or UO_2872 (O_2872,N_49211,N_49366);
or UO_2873 (O_2873,N_49245,N_49138);
or UO_2874 (O_2874,N_49929,N_48506);
and UO_2875 (O_2875,N_48746,N_47755);
nand UO_2876 (O_2876,N_49376,N_48920);
nand UO_2877 (O_2877,N_48273,N_48892);
and UO_2878 (O_2878,N_49035,N_48395);
xor UO_2879 (O_2879,N_47779,N_49305);
nand UO_2880 (O_2880,N_49963,N_47873);
or UO_2881 (O_2881,N_49023,N_48575);
and UO_2882 (O_2882,N_48904,N_48792);
and UO_2883 (O_2883,N_49753,N_49778);
xnor UO_2884 (O_2884,N_48260,N_48461);
nor UO_2885 (O_2885,N_49466,N_49544);
and UO_2886 (O_2886,N_47507,N_48912);
and UO_2887 (O_2887,N_49647,N_48160);
and UO_2888 (O_2888,N_48452,N_47529);
nor UO_2889 (O_2889,N_48634,N_47777);
or UO_2890 (O_2890,N_49317,N_48609);
xor UO_2891 (O_2891,N_49552,N_48672);
xnor UO_2892 (O_2892,N_48608,N_48906);
and UO_2893 (O_2893,N_47711,N_49816);
xnor UO_2894 (O_2894,N_49632,N_49831);
xor UO_2895 (O_2895,N_48459,N_48706);
nor UO_2896 (O_2896,N_49760,N_48764);
or UO_2897 (O_2897,N_49478,N_48958);
xnor UO_2898 (O_2898,N_49302,N_49206);
or UO_2899 (O_2899,N_49243,N_48680);
or UO_2900 (O_2900,N_48785,N_48851);
or UO_2901 (O_2901,N_48952,N_48523);
xnor UO_2902 (O_2902,N_48968,N_47567);
nor UO_2903 (O_2903,N_48444,N_48032);
and UO_2904 (O_2904,N_47759,N_48323);
or UO_2905 (O_2905,N_49039,N_48606);
nor UO_2906 (O_2906,N_49595,N_48907);
nor UO_2907 (O_2907,N_47764,N_47560);
and UO_2908 (O_2908,N_49958,N_49639);
or UO_2909 (O_2909,N_47924,N_47565);
or UO_2910 (O_2910,N_49073,N_48485);
nor UO_2911 (O_2911,N_49167,N_48030);
xor UO_2912 (O_2912,N_48924,N_49470);
or UO_2913 (O_2913,N_48943,N_47559);
nand UO_2914 (O_2914,N_49538,N_49399);
xor UO_2915 (O_2915,N_48295,N_49926);
nor UO_2916 (O_2916,N_48086,N_48186);
nand UO_2917 (O_2917,N_48760,N_49892);
nand UO_2918 (O_2918,N_48011,N_49805);
and UO_2919 (O_2919,N_49960,N_47803);
nand UO_2920 (O_2920,N_47631,N_49194);
or UO_2921 (O_2921,N_48758,N_48698);
nor UO_2922 (O_2922,N_48069,N_47527);
nor UO_2923 (O_2923,N_47816,N_48019);
xnor UO_2924 (O_2924,N_49053,N_49385);
and UO_2925 (O_2925,N_49876,N_47841);
and UO_2926 (O_2926,N_47540,N_49710);
xnor UO_2927 (O_2927,N_49962,N_49171);
nand UO_2928 (O_2928,N_48755,N_48291);
xnor UO_2929 (O_2929,N_49170,N_49862);
nor UO_2930 (O_2930,N_48777,N_49377);
or UO_2931 (O_2931,N_49033,N_48412);
xor UO_2932 (O_2932,N_48717,N_48895);
nand UO_2933 (O_2933,N_49033,N_49778);
and UO_2934 (O_2934,N_47563,N_48031);
nor UO_2935 (O_2935,N_47669,N_47879);
xnor UO_2936 (O_2936,N_47637,N_48080);
or UO_2937 (O_2937,N_49272,N_47643);
nand UO_2938 (O_2938,N_49571,N_49987);
xnor UO_2939 (O_2939,N_49751,N_49307);
or UO_2940 (O_2940,N_48469,N_48728);
nor UO_2941 (O_2941,N_48674,N_48323);
or UO_2942 (O_2942,N_48552,N_49792);
and UO_2943 (O_2943,N_48507,N_47987);
xnor UO_2944 (O_2944,N_47690,N_48797);
and UO_2945 (O_2945,N_47524,N_48498);
and UO_2946 (O_2946,N_48960,N_48371);
nand UO_2947 (O_2947,N_48094,N_47835);
nor UO_2948 (O_2948,N_48833,N_49783);
nor UO_2949 (O_2949,N_47776,N_49365);
xor UO_2950 (O_2950,N_49903,N_47673);
nor UO_2951 (O_2951,N_48286,N_49975);
xor UO_2952 (O_2952,N_49299,N_49588);
and UO_2953 (O_2953,N_49210,N_47756);
and UO_2954 (O_2954,N_47728,N_49163);
xor UO_2955 (O_2955,N_47506,N_49566);
nand UO_2956 (O_2956,N_49047,N_49787);
xnor UO_2957 (O_2957,N_48423,N_49370);
and UO_2958 (O_2958,N_49865,N_49539);
nand UO_2959 (O_2959,N_48445,N_48423);
nor UO_2960 (O_2960,N_47774,N_49800);
nor UO_2961 (O_2961,N_49092,N_48512);
xor UO_2962 (O_2962,N_49605,N_49652);
nor UO_2963 (O_2963,N_48963,N_47718);
nand UO_2964 (O_2964,N_49042,N_47813);
or UO_2965 (O_2965,N_48697,N_48856);
and UO_2966 (O_2966,N_49912,N_48310);
xor UO_2967 (O_2967,N_47792,N_49564);
xnor UO_2968 (O_2968,N_47602,N_49408);
nand UO_2969 (O_2969,N_49708,N_49615);
and UO_2970 (O_2970,N_48197,N_48005);
and UO_2971 (O_2971,N_49693,N_48125);
nand UO_2972 (O_2972,N_48996,N_49564);
xnor UO_2973 (O_2973,N_48020,N_47892);
and UO_2974 (O_2974,N_49763,N_48471);
or UO_2975 (O_2975,N_47598,N_48909);
nor UO_2976 (O_2976,N_47750,N_49772);
nor UO_2977 (O_2977,N_47880,N_49343);
and UO_2978 (O_2978,N_49812,N_49595);
and UO_2979 (O_2979,N_49196,N_48923);
nand UO_2980 (O_2980,N_48463,N_49438);
and UO_2981 (O_2981,N_49815,N_48003);
nor UO_2982 (O_2982,N_47886,N_49602);
or UO_2983 (O_2983,N_49861,N_47922);
nand UO_2984 (O_2984,N_48909,N_47512);
and UO_2985 (O_2985,N_48233,N_48301);
and UO_2986 (O_2986,N_48950,N_47759);
and UO_2987 (O_2987,N_47986,N_47615);
nand UO_2988 (O_2988,N_47513,N_49273);
nor UO_2989 (O_2989,N_47832,N_47608);
and UO_2990 (O_2990,N_48328,N_47523);
or UO_2991 (O_2991,N_48309,N_48809);
nand UO_2992 (O_2992,N_49558,N_47709);
or UO_2993 (O_2993,N_49093,N_49261);
and UO_2994 (O_2994,N_48822,N_48465);
xor UO_2995 (O_2995,N_48689,N_49154);
nand UO_2996 (O_2996,N_49966,N_49553);
nand UO_2997 (O_2997,N_48739,N_47595);
xor UO_2998 (O_2998,N_47537,N_49861);
and UO_2999 (O_2999,N_49316,N_49835);
xor UO_3000 (O_3000,N_49855,N_49645);
nand UO_3001 (O_3001,N_48721,N_48367);
nor UO_3002 (O_3002,N_48113,N_49033);
xnor UO_3003 (O_3003,N_49442,N_48565);
nand UO_3004 (O_3004,N_49699,N_49896);
or UO_3005 (O_3005,N_47511,N_49386);
or UO_3006 (O_3006,N_48532,N_47615);
nor UO_3007 (O_3007,N_49996,N_48389);
nor UO_3008 (O_3008,N_48429,N_47594);
and UO_3009 (O_3009,N_49839,N_49734);
nor UO_3010 (O_3010,N_48928,N_49336);
or UO_3011 (O_3011,N_48744,N_48892);
or UO_3012 (O_3012,N_48917,N_47859);
nand UO_3013 (O_3013,N_49825,N_48160);
nor UO_3014 (O_3014,N_47642,N_49091);
nor UO_3015 (O_3015,N_48528,N_48545);
nand UO_3016 (O_3016,N_49717,N_49994);
xor UO_3017 (O_3017,N_49010,N_49332);
or UO_3018 (O_3018,N_48099,N_48168);
nand UO_3019 (O_3019,N_49905,N_49156);
xnor UO_3020 (O_3020,N_48389,N_48813);
nor UO_3021 (O_3021,N_49326,N_48088);
or UO_3022 (O_3022,N_49103,N_48767);
xor UO_3023 (O_3023,N_48292,N_49073);
or UO_3024 (O_3024,N_49456,N_49138);
nand UO_3025 (O_3025,N_47705,N_48201);
nor UO_3026 (O_3026,N_49815,N_49906);
xor UO_3027 (O_3027,N_48693,N_47816);
nor UO_3028 (O_3028,N_48766,N_48156);
nand UO_3029 (O_3029,N_49166,N_49292);
nand UO_3030 (O_3030,N_48185,N_49855);
nor UO_3031 (O_3031,N_48221,N_49236);
xnor UO_3032 (O_3032,N_48684,N_49152);
nand UO_3033 (O_3033,N_47926,N_49567);
nor UO_3034 (O_3034,N_47839,N_49769);
xnor UO_3035 (O_3035,N_49237,N_47633);
nand UO_3036 (O_3036,N_48585,N_47981);
nor UO_3037 (O_3037,N_47545,N_49953);
xor UO_3038 (O_3038,N_49652,N_48723);
and UO_3039 (O_3039,N_49685,N_49726);
and UO_3040 (O_3040,N_48184,N_47638);
xnor UO_3041 (O_3041,N_48022,N_48655);
nand UO_3042 (O_3042,N_49574,N_48949);
and UO_3043 (O_3043,N_49433,N_49185);
nand UO_3044 (O_3044,N_48088,N_47588);
nor UO_3045 (O_3045,N_47914,N_48096);
or UO_3046 (O_3046,N_49968,N_49318);
and UO_3047 (O_3047,N_47769,N_49579);
nor UO_3048 (O_3048,N_47504,N_48247);
nor UO_3049 (O_3049,N_48646,N_49847);
or UO_3050 (O_3050,N_48275,N_48105);
nand UO_3051 (O_3051,N_47769,N_49640);
xnor UO_3052 (O_3052,N_49567,N_49922);
or UO_3053 (O_3053,N_48258,N_49325);
nand UO_3054 (O_3054,N_48492,N_47557);
nor UO_3055 (O_3055,N_49263,N_49746);
or UO_3056 (O_3056,N_48343,N_47727);
nor UO_3057 (O_3057,N_49723,N_47651);
nand UO_3058 (O_3058,N_48746,N_47572);
or UO_3059 (O_3059,N_48455,N_47551);
nor UO_3060 (O_3060,N_49259,N_48135);
xor UO_3061 (O_3061,N_48749,N_47961);
nor UO_3062 (O_3062,N_48096,N_49137);
and UO_3063 (O_3063,N_49334,N_48912);
nand UO_3064 (O_3064,N_49084,N_48599);
nand UO_3065 (O_3065,N_48916,N_47510);
xnor UO_3066 (O_3066,N_48026,N_48573);
or UO_3067 (O_3067,N_48303,N_49353);
xnor UO_3068 (O_3068,N_48368,N_47841);
nand UO_3069 (O_3069,N_48576,N_48024);
or UO_3070 (O_3070,N_47598,N_48222);
and UO_3071 (O_3071,N_48278,N_49918);
nor UO_3072 (O_3072,N_48966,N_49112);
nand UO_3073 (O_3073,N_48840,N_48772);
and UO_3074 (O_3074,N_48488,N_49377);
and UO_3075 (O_3075,N_47757,N_48508);
xor UO_3076 (O_3076,N_49188,N_49177);
nor UO_3077 (O_3077,N_47977,N_49732);
or UO_3078 (O_3078,N_47702,N_48634);
nand UO_3079 (O_3079,N_47647,N_48108);
and UO_3080 (O_3080,N_49727,N_48745);
and UO_3081 (O_3081,N_48577,N_48065);
nor UO_3082 (O_3082,N_48450,N_49014);
and UO_3083 (O_3083,N_47683,N_48895);
and UO_3084 (O_3084,N_48029,N_47537);
nand UO_3085 (O_3085,N_47683,N_48306);
and UO_3086 (O_3086,N_48641,N_49147);
nand UO_3087 (O_3087,N_49128,N_48690);
nand UO_3088 (O_3088,N_47560,N_48823);
xor UO_3089 (O_3089,N_48818,N_48677);
nor UO_3090 (O_3090,N_49651,N_48534);
or UO_3091 (O_3091,N_47617,N_48064);
xor UO_3092 (O_3092,N_49594,N_48284);
nand UO_3093 (O_3093,N_48909,N_49482);
xnor UO_3094 (O_3094,N_49491,N_47724);
nand UO_3095 (O_3095,N_49079,N_47974);
xor UO_3096 (O_3096,N_48372,N_48694);
and UO_3097 (O_3097,N_49505,N_47815);
nor UO_3098 (O_3098,N_48402,N_47540);
xor UO_3099 (O_3099,N_49174,N_48435);
and UO_3100 (O_3100,N_47819,N_48657);
nand UO_3101 (O_3101,N_49356,N_48864);
and UO_3102 (O_3102,N_48844,N_47775);
xor UO_3103 (O_3103,N_47817,N_49906);
xnor UO_3104 (O_3104,N_49637,N_49326);
and UO_3105 (O_3105,N_49009,N_47555);
nand UO_3106 (O_3106,N_49871,N_48512);
or UO_3107 (O_3107,N_48936,N_49368);
nor UO_3108 (O_3108,N_49042,N_49852);
nor UO_3109 (O_3109,N_49751,N_49240);
or UO_3110 (O_3110,N_48529,N_49655);
and UO_3111 (O_3111,N_49045,N_48970);
nand UO_3112 (O_3112,N_49182,N_49592);
nand UO_3113 (O_3113,N_47640,N_47558);
xnor UO_3114 (O_3114,N_48232,N_47608);
nor UO_3115 (O_3115,N_48428,N_49466);
xnor UO_3116 (O_3116,N_49493,N_49226);
xor UO_3117 (O_3117,N_48602,N_48854);
nand UO_3118 (O_3118,N_47997,N_48366);
nor UO_3119 (O_3119,N_49517,N_48775);
nor UO_3120 (O_3120,N_48515,N_48392);
xor UO_3121 (O_3121,N_48119,N_49193);
nand UO_3122 (O_3122,N_47802,N_48564);
xnor UO_3123 (O_3123,N_48521,N_49912);
and UO_3124 (O_3124,N_48193,N_48734);
nor UO_3125 (O_3125,N_48008,N_49370);
and UO_3126 (O_3126,N_49558,N_48935);
or UO_3127 (O_3127,N_49637,N_48691);
nand UO_3128 (O_3128,N_49129,N_48869);
and UO_3129 (O_3129,N_48297,N_47938);
or UO_3130 (O_3130,N_48627,N_48107);
nor UO_3131 (O_3131,N_47809,N_47505);
and UO_3132 (O_3132,N_49671,N_48433);
and UO_3133 (O_3133,N_49411,N_49891);
and UO_3134 (O_3134,N_49794,N_47643);
and UO_3135 (O_3135,N_49789,N_49014);
and UO_3136 (O_3136,N_47646,N_49116);
nor UO_3137 (O_3137,N_48898,N_48702);
and UO_3138 (O_3138,N_48450,N_48366);
nor UO_3139 (O_3139,N_48047,N_49250);
nand UO_3140 (O_3140,N_49192,N_49196);
nand UO_3141 (O_3141,N_47536,N_49656);
nor UO_3142 (O_3142,N_48971,N_49533);
and UO_3143 (O_3143,N_49221,N_48728);
nor UO_3144 (O_3144,N_48416,N_48244);
or UO_3145 (O_3145,N_48434,N_48312);
xor UO_3146 (O_3146,N_49394,N_49967);
and UO_3147 (O_3147,N_47618,N_47830);
nand UO_3148 (O_3148,N_49540,N_48625);
xnor UO_3149 (O_3149,N_48165,N_48279);
and UO_3150 (O_3150,N_49207,N_49388);
nand UO_3151 (O_3151,N_47724,N_48836);
nor UO_3152 (O_3152,N_47863,N_49721);
and UO_3153 (O_3153,N_49660,N_48031);
or UO_3154 (O_3154,N_47804,N_49755);
nand UO_3155 (O_3155,N_47748,N_48077);
nor UO_3156 (O_3156,N_49276,N_49950);
and UO_3157 (O_3157,N_48254,N_49460);
xor UO_3158 (O_3158,N_49918,N_47730);
nor UO_3159 (O_3159,N_48651,N_47522);
nor UO_3160 (O_3160,N_49114,N_48134);
xor UO_3161 (O_3161,N_47684,N_48766);
nand UO_3162 (O_3162,N_47667,N_49647);
nand UO_3163 (O_3163,N_49767,N_49002);
nand UO_3164 (O_3164,N_49457,N_49093);
or UO_3165 (O_3165,N_47761,N_48800);
xnor UO_3166 (O_3166,N_49983,N_49586);
and UO_3167 (O_3167,N_49979,N_48898);
xnor UO_3168 (O_3168,N_49469,N_48648);
nand UO_3169 (O_3169,N_49212,N_48839);
and UO_3170 (O_3170,N_49640,N_49653);
nand UO_3171 (O_3171,N_48629,N_48551);
and UO_3172 (O_3172,N_49954,N_48558);
xor UO_3173 (O_3173,N_49333,N_48348);
or UO_3174 (O_3174,N_48379,N_48081);
nand UO_3175 (O_3175,N_47792,N_49890);
or UO_3176 (O_3176,N_49716,N_49004);
or UO_3177 (O_3177,N_47602,N_48636);
and UO_3178 (O_3178,N_49208,N_47619);
nand UO_3179 (O_3179,N_48596,N_49387);
or UO_3180 (O_3180,N_47820,N_48086);
nand UO_3181 (O_3181,N_49353,N_48508);
xnor UO_3182 (O_3182,N_48278,N_48662);
nor UO_3183 (O_3183,N_48865,N_48806);
or UO_3184 (O_3184,N_49947,N_47645);
xnor UO_3185 (O_3185,N_48580,N_49625);
xnor UO_3186 (O_3186,N_49223,N_48317);
xor UO_3187 (O_3187,N_49654,N_49730);
and UO_3188 (O_3188,N_48558,N_48480);
nand UO_3189 (O_3189,N_47873,N_48727);
nand UO_3190 (O_3190,N_47804,N_49456);
nand UO_3191 (O_3191,N_48581,N_48209);
or UO_3192 (O_3192,N_48928,N_48163);
nor UO_3193 (O_3193,N_48306,N_49678);
or UO_3194 (O_3194,N_49724,N_49687);
and UO_3195 (O_3195,N_47924,N_48601);
and UO_3196 (O_3196,N_49934,N_47662);
or UO_3197 (O_3197,N_49083,N_49679);
nand UO_3198 (O_3198,N_49019,N_48540);
or UO_3199 (O_3199,N_48413,N_49080);
xor UO_3200 (O_3200,N_48734,N_47790);
or UO_3201 (O_3201,N_49333,N_48535);
and UO_3202 (O_3202,N_48831,N_49214);
nor UO_3203 (O_3203,N_49678,N_49643);
nor UO_3204 (O_3204,N_48522,N_48973);
nor UO_3205 (O_3205,N_49866,N_47704);
xor UO_3206 (O_3206,N_48031,N_48622);
and UO_3207 (O_3207,N_49560,N_48556);
nand UO_3208 (O_3208,N_49202,N_48275);
xnor UO_3209 (O_3209,N_48591,N_49382);
nor UO_3210 (O_3210,N_49185,N_49153);
and UO_3211 (O_3211,N_47572,N_49047);
and UO_3212 (O_3212,N_47715,N_48349);
and UO_3213 (O_3213,N_47766,N_47507);
and UO_3214 (O_3214,N_48127,N_48675);
nand UO_3215 (O_3215,N_49827,N_48470);
nand UO_3216 (O_3216,N_49731,N_47851);
nor UO_3217 (O_3217,N_48279,N_49353);
nor UO_3218 (O_3218,N_49259,N_49386);
or UO_3219 (O_3219,N_47570,N_47695);
nor UO_3220 (O_3220,N_47834,N_49791);
xor UO_3221 (O_3221,N_47821,N_48060);
nand UO_3222 (O_3222,N_49783,N_48905);
nand UO_3223 (O_3223,N_49401,N_49103);
or UO_3224 (O_3224,N_48017,N_48636);
nor UO_3225 (O_3225,N_47803,N_49502);
nor UO_3226 (O_3226,N_49861,N_48039);
xnor UO_3227 (O_3227,N_48169,N_48081);
and UO_3228 (O_3228,N_48130,N_49116);
xnor UO_3229 (O_3229,N_48961,N_47858);
nand UO_3230 (O_3230,N_49748,N_49207);
and UO_3231 (O_3231,N_49410,N_48991);
nor UO_3232 (O_3232,N_48347,N_49419);
nor UO_3233 (O_3233,N_49740,N_49249);
or UO_3234 (O_3234,N_49503,N_48264);
xor UO_3235 (O_3235,N_48423,N_49192);
xor UO_3236 (O_3236,N_48576,N_48489);
xor UO_3237 (O_3237,N_48828,N_48057);
xnor UO_3238 (O_3238,N_47641,N_48590);
xor UO_3239 (O_3239,N_49675,N_49249);
or UO_3240 (O_3240,N_47852,N_47811);
or UO_3241 (O_3241,N_49320,N_49123);
nand UO_3242 (O_3242,N_49152,N_48456);
and UO_3243 (O_3243,N_48482,N_48509);
nor UO_3244 (O_3244,N_49208,N_48682);
or UO_3245 (O_3245,N_49941,N_48768);
xor UO_3246 (O_3246,N_48717,N_49630);
and UO_3247 (O_3247,N_49114,N_47568);
nand UO_3248 (O_3248,N_48638,N_47504);
and UO_3249 (O_3249,N_49065,N_48418);
or UO_3250 (O_3250,N_48476,N_48307);
xor UO_3251 (O_3251,N_47717,N_48520);
xor UO_3252 (O_3252,N_47787,N_49838);
nand UO_3253 (O_3253,N_49943,N_48849);
nand UO_3254 (O_3254,N_48675,N_48640);
xnor UO_3255 (O_3255,N_48935,N_48938);
nor UO_3256 (O_3256,N_48296,N_49765);
and UO_3257 (O_3257,N_49544,N_48719);
nor UO_3258 (O_3258,N_48937,N_49873);
nor UO_3259 (O_3259,N_48535,N_49905);
nand UO_3260 (O_3260,N_49358,N_48201);
or UO_3261 (O_3261,N_49342,N_49059);
nand UO_3262 (O_3262,N_48683,N_48441);
xor UO_3263 (O_3263,N_48109,N_49825);
nor UO_3264 (O_3264,N_48553,N_47921);
or UO_3265 (O_3265,N_48390,N_47727);
xor UO_3266 (O_3266,N_47803,N_48359);
xnor UO_3267 (O_3267,N_49007,N_48617);
and UO_3268 (O_3268,N_49763,N_49179);
and UO_3269 (O_3269,N_47898,N_47658);
and UO_3270 (O_3270,N_47979,N_49046);
nand UO_3271 (O_3271,N_48343,N_47705);
nand UO_3272 (O_3272,N_48240,N_49135);
nand UO_3273 (O_3273,N_48334,N_48861);
nor UO_3274 (O_3274,N_49107,N_48629);
and UO_3275 (O_3275,N_48899,N_48758);
nand UO_3276 (O_3276,N_48521,N_47563);
nand UO_3277 (O_3277,N_48785,N_48337);
xnor UO_3278 (O_3278,N_49701,N_48723);
xnor UO_3279 (O_3279,N_48781,N_47769);
nand UO_3280 (O_3280,N_49494,N_49574);
or UO_3281 (O_3281,N_48430,N_49154);
xor UO_3282 (O_3282,N_49699,N_48436);
and UO_3283 (O_3283,N_49859,N_49352);
xor UO_3284 (O_3284,N_48561,N_47994);
nand UO_3285 (O_3285,N_49977,N_47904);
and UO_3286 (O_3286,N_49462,N_48154);
or UO_3287 (O_3287,N_49901,N_48614);
and UO_3288 (O_3288,N_49377,N_49891);
nand UO_3289 (O_3289,N_49592,N_47908);
nand UO_3290 (O_3290,N_49335,N_49754);
xnor UO_3291 (O_3291,N_49249,N_48455);
xnor UO_3292 (O_3292,N_49477,N_49044);
and UO_3293 (O_3293,N_48108,N_48082);
or UO_3294 (O_3294,N_48746,N_49886);
nor UO_3295 (O_3295,N_47854,N_49918);
or UO_3296 (O_3296,N_48038,N_48903);
xnor UO_3297 (O_3297,N_49732,N_49449);
nand UO_3298 (O_3298,N_48597,N_49223);
and UO_3299 (O_3299,N_49844,N_48628);
and UO_3300 (O_3300,N_48847,N_48782);
and UO_3301 (O_3301,N_48049,N_47821);
and UO_3302 (O_3302,N_49230,N_47734);
or UO_3303 (O_3303,N_49227,N_47616);
or UO_3304 (O_3304,N_47638,N_47760);
and UO_3305 (O_3305,N_47745,N_47979);
nor UO_3306 (O_3306,N_47546,N_48709);
and UO_3307 (O_3307,N_49529,N_47664);
or UO_3308 (O_3308,N_49042,N_48634);
nand UO_3309 (O_3309,N_48578,N_47907);
xnor UO_3310 (O_3310,N_48212,N_48476);
nor UO_3311 (O_3311,N_48957,N_48622);
xnor UO_3312 (O_3312,N_48704,N_48477);
nor UO_3313 (O_3313,N_49476,N_48501);
nor UO_3314 (O_3314,N_49014,N_49646);
xor UO_3315 (O_3315,N_47537,N_48470);
xor UO_3316 (O_3316,N_47854,N_49964);
and UO_3317 (O_3317,N_49792,N_47539);
and UO_3318 (O_3318,N_48505,N_48784);
and UO_3319 (O_3319,N_49094,N_48878);
nor UO_3320 (O_3320,N_49958,N_48791);
or UO_3321 (O_3321,N_49565,N_47716);
and UO_3322 (O_3322,N_49572,N_48017);
xnor UO_3323 (O_3323,N_48482,N_47541);
xnor UO_3324 (O_3324,N_47693,N_49231);
and UO_3325 (O_3325,N_48651,N_47860);
or UO_3326 (O_3326,N_48473,N_48004);
nor UO_3327 (O_3327,N_48334,N_48188);
nand UO_3328 (O_3328,N_48927,N_47755);
or UO_3329 (O_3329,N_48371,N_49575);
and UO_3330 (O_3330,N_49005,N_47680);
or UO_3331 (O_3331,N_48712,N_49080);
nand UO_3332 (O_3332,N_47890,N_48525);
nor UO_3333 (O_3333,N_47811,N_49542);
or UO_3334 (O_3334,N_47803,N_48584);
nand UO_3335 (O_3335,N_49292,N_49221);
xor UO_3336 (O_3336,N_49411,N_49863);
xnor UO_3337 (O_3337,N_49947,N_47945);
and UO_3338 (O_3338,N_48384,N_49951);
nand UO_3339 (O_3339,N_47811,N_49296);
or UO_3340 (O_3340,N_49043,N_47846);
nor UO_3341 (O_3341,N_48453,N_49313);
xnor UO_3342 (O_3342,N_47669,N_47618);
nor UO_3343 (O_3343,N_49217,N_49746);
nand UO_3344 (O_3344,N_49535,N_48064);
and UO_3345 (O_3345,N_48343,N_48913);
xor UO_3346 (O_3346,N_49816,N_48935);
and UO_3347 (O_3347,N_49911,N_47572);
nand UO_3348 (O_3348,N_47515,N_47588);
and UO_3349 (O_3349,N_49989,N_48385);
xnor UO_3350 (O_3350,N_48577,N_48879);
or UO_3351 (O_3351,N_49477,N_48704);
xnor UO_3352 (O_3352,N_49394,N_48859);
or UO_3353 (O_3353,N_47604,N_49129);
nor UO_3354 (O_3354,N_47959,N_47679);
and UO_3355 (O_3355,N_47660,N_49565);
nor UO_3356 (O_3356,N_49744,N_48732);
nor UO_3357 (O_3357,N_48424,N_49243);
xnor UO_3358 (O_3358,N_48910,N_49166);
nor UO_3359 (O_3359,N_49919,N_48276);
nand UO_3360 (O_3360,N_49390,N_48843);
xnor UO_3361 (O_3361,N_48664,N_48046);
or UO_3362 (O_3362,N_47644,N_49780);
or UO_3363 (O_3363,N_49639,N_48691);
and UO_3364 (O_3364,N_48705,N_48940);
nor UO_3365 (O_3365,N_48576,N_48319);
and UO_3366 (O_3366,N_47902,N_49145);
or UO_3367 (O_3367,N_49778,N_48546);
nor UO_3368 (O_3368,N_47861,N_49270);
xnor UO_3369 (O_3369,N_49956,N_48800);
nor UO_3370 (O_3370,N_49685,N_48795);
xor UO_3371 (O_3371,N_49350,N_49811);
xor UO_3372 (O_3372,N_49510,N_49864);
xor UO_3373 (O_3373,N_49048,N_47552);
xor UO_3374 (O_3374,N_48114,N_48903);
xor UO_3375 (O_3375,N_49911,N_49509);
xnor UO_3376 (O_3376,N_47670,N_49814);
and UO_3377 (O_3377,N_48479,N_47736);
nor UO_3378 (O_3378,N_48080,N_49263);
or UO_3379 (O_3379,N_49570,N_49113);
or UO_3380 (O_3380,N_47804,N_49312);
or UO_3381 (O_3381,N_49217,N_49252);
and UO_3382 (O_3382,N_49433,N_48422);
xor UO_3383 (O_3383,N_48127,N_49322);
or UO_3384 (O_3384,N_48660,N_49624);
or UO_3385 (O_3385,N_48450,N_48398);
nand UO_3386 (O_3386,N_48460,N_48492);
or UO_3387 (O_3387,N_49303,N_49912);
nor UO_3388 (O_3388,N_48338,N_48554);
nor UO_3389 (O_3389,N_47932,N_49949);
or UO_3390 (O_3390,N_48414,N_48691);
nand UO_3391 (O_3391,N_49262,N_47916);
nand UO_3392 (O_3392,N_49502,N_48967);
and UO_3393 (O_3393,N_47862,N_48547);
or UO_3394 (O_3394,N_49066,N_48314);
or UO_3395 (O_3395,N_47530,N_48930);
and UO_3396 (O_3396,N_49780,N_47679);
nand UO_3397 (O_3397,N_49662,N_48035);
and UO_3398 (O_3398,N_47768,N_47619);
and UO_3399 (O_3399,N_48066,N_47774);
nor UO_3400 (O_3400,N_49528,N_48690);
xor UO_3401 (O_3401,N_49281,N_49596);
or UO_3402 (O_3402,N_48834,N_49962);
and UO_3403 (O_3403,N_48205,N_49613);
nand UO_3404 (O_3404,N_49874,N_47526);
nand UO_3405 (O_3405,N_48292,N_48564);
nor UO_3406 (O_3406,N_48056,N_49011);
or UO_3407 (O_3407,N_49173,N_49092);
nand UO_3408 (O_3408,N_49165,N_49841);
and UO_3409 (O_3409,N_48373,N_47589);
or UO_3410 (O_3410,N_49984,N_48239);
or UO_3411 (O_3411,N_49832,N_47550);
and UO_3412 (O_3412,N_49567,N_47667);
nand UO_3413 (O_3413,N_47748,N_48532);
nand UO_3414 (O_3414,N_48743,N_47645);
or UO_3415 (O_3415,N_49950,N_48594);
xor UO_3416 (O_3416,N_48551,N_48164);
and UO_3417 (O_3417,N_47919,N_48486);
or UO_3418 (O_3418,N_48776,N_48194);
or UO_3419 (O_3419,N_48967,N_49190);
xnor UO_3420 (O_3420,N_48271,N_49050);
or UO_3421 (O_3421,N_48360,N_49610);
nand UO_3422 (O_3422,N_49038,N_47587);
and UO_3423 (O_3423,N_49919,N_47962);
and UO_3424 (O_3424,N_48412,N_49457);
xnor UO_3425 (O_3425,N_49839,N_48617);
xnor UO_3426 (O_3426,N_49057,N_48393);
xnor UO_3427 (O_3427,N_48700,N_49515);
nand UO_3428 (O_3428,N_49053,N_47571);
nor UO_3429 (O_3429,N_48455,N_47633);
nand UO_3430 (O_3430,N_49504,N_49496);
and UO_3431 (O_3431,N_47998,N_47630);
or UO_3432 (O_3432,N_49084,N_49790);
and UO_3433 (O_3433,N_47530,N_48926);
nor UO_3434 (O_3434,N_47524,N_49786);
and UO_3435 (O_3435,N_48941,N_47900);
nor UO_3436 (O_3436,N_47705,N_47838);
nand UO_3437 (O_3437,N_48311,N_49511);
or UO_3438 (O_3438,N_49790,N_48400);
or UO_3439 (O_3439,N_48286,N_49909);
nor UO_3440 (O_3440,N_49017,N_49531);
or UO_3441 (O_3441,N_49498,N_47672);
nor UO_3442 (O_3442,N_48245,N_49101);
nor UO_3443 (O_3443,N_48690,N_49689);
and UO_3444 (O_3444,N_49275,N_49384);
nor UO_3445 (O_3445,N_49002,N_49594);
or UO_3446 (O_3446,N_48525,N_48118);
xnor UO_3447 (O_3447,N_49176,N_49855);
and UO_3448 (O_3448,N_47527,N_49772);
or UO_3449 (O_3449,N_49616,N_49708);
nand UO_3450 (O_3450,N_49590,N_48306);
and UO_3451 (O_3451,N_48615,N_48129);
xor UO_3452 (O_3452,N_48780,N_48320);
or UO_3453 (O_3453,N_48972,N_48005);
nor UO_3454 (O_3454,N_49005,N_49018);
or UO_3455 (O_3455,N_48621,N_49670);
and UO_3456 (O_3456,N_49920,N_47977);
xor UO_3457 (O_3457,N_49441,N_49985);
nor UO_3458 (O_3458,N_48300,N_49511);
or UO_3459 (O_3459,N_47704,N_48282);
nor UO_3460 (O_3460,N_49751,N_47796);
xor UO_3461 (O_3461,N_47957,N_49297);
nand UO_3462 (O_3462,N_49828,N_48158);
nor UO_3463 (O_3463,N_47696,N_49138);
xnor UO_3464 (O_3464,N_47534,N_48332);
nand UO_3465 (O_3465,N_49549,N_48646);
nor UO_3466 (O_3466,N_49963,N_47801);
and UO_3467 (O_3467,N_47841,N_48532);
nor UO_3468 (O_3468,N_48308,N_48454);
or UO_3469 (O_3469,N_49128,N_47527);
or UO_3470 (O_3470,N_49095,N_49337);
nor UO_3471 (O_3471,N_47616,N_48847);
or UO_3472 (O_3472,N_49137,N_47805);
xnor UO_3473 (O_3473,N_48637,N_47702);
and UO_3474 (O_3474,N_49596,N_48297);
nor UO_3475 (O_3475,N_48306,N_48469);
nand UO_3476 (O_3476,N_49690,N_47570);
and UO_3477 (O_3477,N_48013,N_49399);
nor UO_3478 (O_3478,N_48319,N_49760);
nor UO_3479 (O_3479,N_49214,N_49810);
xnor UO_3480 (O_3480,N_48691,N_49068);
xor UO_3481 (O_3481,N_48666,N_48244);
nand UO_3482 (O_3482,N_48842,N_49596);
nand UO_3483 (O_3483,N_49590,N_48448);
xnor UO_3484 (O_3484,N_49702,N_49055);
and UO_3485 (O_3485,N_48110,N_48397);
or UO_3486 (O_3486,N_49592,N_49744);
nand UO_3487 (O_3487,N_49498,N_48331);
and UO_3488 (O_3488,N_48728,N_47688);
nor UO_3489 (O_3489,N_49176,N_49481);
or UO_3490 (O_3490,N_49661,N_49161);
xor UO_3491 (O_3491,N_49663,N_49432);
nand UO_3492 (O_3492,N_49709,N_48164);
or UO_3493 (O_3493,N_49752,N_49657);
and UO_3494 (O_3494,N_49249,N_48719);
and UO_3495 (O_3495,N_48629,N_48447);
and UO_3496 (O_3496,N_48136,N_48028);
nor UO_3497 (O_3497,N_48490,N_49066);
nor UO_3498 (O_3498,N_49891,N_47793);
xor UO_3499 (O_3499,N_48691,N_47879);
nand UO_3500 (O_3500,N_48005,N_48519);
nor UO_3501 (O_3501,N_49619,N_49797);
xnor UO_3502 (O_3502,N_49536,N_47873);
xor UO_3503 (O_3503,N_47707,N_49203);
nor UO_3504 (O_3504,N_48746,N_49103);
and UO_3505 (O_3505,N_49066,N_47677);
or UO_3506 (O_3506,N_49568,N_47557);
nor UO_3507 (O_3507,N_47976,N_49999);
nor UO_3508 (O_3508,N_48021,N_48793);
nor UO_3509 (O_3509,N_47548,N_49789);
nand UO_3510 (O_3510,N_49078,N_47813);
and UO_3511 (O_3511,N_47992,N_49244);
nand UO_3512 (O_3512,N_47545,N_47620);
or UO_3513 (O_3513,N_48367,N_48877);
and UO_3514 (O_3514,N_48718,N_48652);
or UO_3515 (O_3515,N_48260,N_48272);
nand UO_3516 (O_3516,N_48698,N_48258);
or UO_3517 (O_3517,N_49710,N_48291);
or UO_3518 (O_3518,N_49802,N_48845);
xor UO_3519 (O_3519,N_48535,N_48664);
and UO_3520 (O_3520,N_49325,N_48157);
xor UO_3521 (O_3521,N_48145,N_47984);
or UO_3522 (O_3522,N_49650,N_49093);
and UO_3523 (O_3523,N_48641,N_49928);
and UO_3524 (O_3524,N_49670,N_48597);
or UO_3525 (O_3525,N_49630,N_49595);
xor UO_3526 (O_3526,N_48758,N_49124);
and UO_3527 (O_3527,N_47563,N_49145);
nand UO_3528 (O_3528,N_49297,N_48170);
and UO_3529 (O_3529,N_47957,N_49542);
and UO_3530 (O_3530,N_48672,N_48644);
nor UO_3531 (O_3531,N_47528,N_49939);
nand UO_3532 (O_3532,N_48433,N_47706);
and UO_3533 (O_3533,N_48920,N_47813);
nor UO_3534 (O_3534,N_48221,N_47732);
or UO_3535 (O_3535,N_48699,N_48432);
nor UO_3536 (O_3536,N_49838,N_47914);
nor UO_3537 (O_3537,N_48866,N_49698);
nor UO_3538 (O_3538,N_49593,N_49343);
and UO_3539 (O_3539,N_49609,N_49630);
or UO_3540 (O_3540,N_48656,N_47942);
xnor UO_3541 (O_3541,N_49808,N_47924);
xnor UO_3542 (O_3542,N_48682,N_47937);
and UO_3543 (O_3543,N_49685,N_48623);
nand UO_3544 (O_3544,N_49725,N_49323);
nand UO_3545 (O_3545,N_48390,N_48125);
xnor UO_3546 (O_3546,N_47500,N_48117);
xor UO_3547 (O_3547,N_49328,N_49637);
nor UO_3548 (O_3548,N_49732,N_49020);
xor UO_3549 (O_3549,N_48546,N_48693);
or UO_3550 (O_3550,N_48424,N_49294);
xnor UO_3551 (O_3551,N_48406,N_49622);
and UO_3552 (O_3552,N_48257,N_47619);
xnor UO_3553 (O_3553,N_48246,N_48807);
nand UO_3554 (O_3554,N_48844,N_47677);
and UO_3555 (O_3555,N_49056,N_49230);
xnor UO_3556 (O_3556,N_48316,N_49750);
xor UO_3557 (O_3557,N_48117,N_48811);
xnor UO_3558 (O_3558,N_49840,N_48996);
and UO_3559 (O_3559,N_47534,N_49433);
xor UO_3560 (O_3560,N_49344,N_48874);
nand UO_3561 (O_3561,N_47581,N_47966);
nand UO_3562 (O_3562,N_49382,N_48051);
nor UO_3563 (O_3563,N_48002,N_49360);
nor UO_3564 (O_3564,N_48686,N_49259);
and UO_3565 (O_3565,N_48067,N_49851);
and UO_3566 (O_3566,N_48125,N_47593);
and UO_3567 (O_3567,N_49278,N_47702);
nand UO_3568 (O_3568,N_48647,N_49834);
or UO_3569 (O_3569,N_48617,N_49320);
nand UO_3570 (O_3570,N_48114,N_47509);
nor UO_3571 (O_3571,N_49532,N_49207);
and UO_3572 (O_3572,N_48486,N_48454);
nor UO_3573 (O_3573,N_47918,N_49435);
or UO_3574 (O_3574,N_48930,N_49568);
nand UO_3575 (O_3575,N_49197,N_49814);
xor UO_3576 (O_3576,N_47518,N_47847);
xnor UO_3577 (O_3577,N_48312,N_48895);
nand UO_3578 (O_3578,N_47678,N_49571);
xor UO_3579 (O_3579,N_49314,N_48323);
and UO_3580 (O_3580,N_48372,N_49063);
xnor UO_3581 (O_3581,N_48721,N_49225);
nor UO_3582 (O_3582,N_49158,N_48475);
xor UO_3583 (O_3583,N_49808,N_49243);
nand UO_3584 (O_3584,N_47993,N_47926);
xnor UO_3585 (O_3585,N_47558,N_48172);
and UO_3586 (O_3586,N_48210,N_49095);
and UO_3587 (O_3587,N_47597,N_48311);
and UO_3588 (O_3588,N_49843,N_47850);
nand UO_3589 (O_3589,N_47957,N_49658);
and UO_3590 (O_3590,N_48252,N_49855);
and UO_3591 (O_3591,N_47568,N_47881);
and UO_3592 (O_3592,N_49214,N_47918);
xnor UO_3593 (O_3593,N_49439,N_49393);
nor UO_3594 (O_3594,N_47525,N_49176);
xnor UO_3595 (O_3595,N_48068,N_48751);
xnor UO_3596 (O_3596,N_49434,N_49353);
and UO_3597 (O_3597,N_48926,N_49732);
xnor UO_3598 (O_3598,N_48594,N_48052);
and UO_3599 (O_3599,N_47605,N_49807);
or UO_3600 (O_3600,N_47622,N_49995);
nor UO_3601 (O_3601,N_49832,N_48753);
and UO_3602 (O_3602,N_47915,N_47963);
xnor UO_3603 (O_3603,N_49112,N_48890);
and UO_3604 (O_3604,N_48769,N_49770);
xnor UO_3605 (O_3605,N_48165,N_48308);
or UO_3606 (O_3606,N_49400,N_48141);
or UO_3607 (O_3607,N_48247,N_49275);
or UO_3608 (O_3608,N_49251,N_48874);
and UO_3609 (O_3609,N_49125,N_48361);
nor UO_3610 (O_3610,N_49408,N_49614);
nand UO_3611 (O_3611,N_49888,N_48783);
and UO_3612 (O_3612,N_48696,N_48588);
or UO_3613 (O_3613,N_48610,N_49026);
xor UO_3614 (O_3614,N_48061,N_47793);
or UO_3615 (O_3615,N_47992,N_49061);
or UO_3616 (O_3616,N_48567,N_49855);
nand UO_3617 (O_3617,N_48018,N_49541);
and UO_3618 (O_3618,N_49949,N_48846);
nand UO_3619 (O_3619,N_49081,N_48396);
or UO_3620 (O_3620,N_48780,N_47635);
nor UO_3621 (O_3621,N_48629,N_48080);
xor UO_3622 (O_3622,N_49784,N_49652);
nand UO_3623 (O_3623,N_49116,N_49624);
or UO_3624 (O_3624,N_49456,N_48968);
xor UO_3625 (O_3625,N_48152,N_49976);
or UO_3626 (O_3626,N_49290,N_48902);
or UO_3627 (O_3627,N_48898,N_49507);
nor UO_3628 (O_3628,N_49041,N_48378);
and UO_3629 (O_3629,N_48991,N_47750);
and UO_3630 (O_3630,N_48864,N_48484);
nand UO_3631 (O_3631,N_49966,N_49814);
xnor UO_3632 (O_3632,N_48603,N_49806);
or UO_3633 (O_3633,N_47535,N_48616);
nor UO_3634 (O_3634,N_48925,N_49812);
xnor UO_3635 (O_3635,N_48370,N_48549);
nor UO_3636 (O_3636,N_48241,N_48079);
xnor UO_3637 (O_3637,N_49194,N_49319);
nor UO_3638 (O_3638,N_49356,N_49237);
and UO_3639 (O_3639,N_47998,N_49314);
nor UO_3640 (O_3640,N_49450,N_49325);
nand UO_3641 (O_3641,N_49073,N_48213);
xnor UO_3642 (O_3642,N_49178,N_47950);
nand UO_3643 (O_3643,N_47941,N_48801);
xnor UO_3644 (O_3644,N_49809,N_47670);
and UO_3645 (O_3645,N_48112,N_49094);
or UO_3646 (O_3646,N_47839,N_48458);
nand UO_3647 (O_3647,N_48889,N_47603);
and UO_3648 (O_3648,N_49978,N_49461);
nand UO_3649 (O_3649,N_47544,N_49209);
nand UO_3650 (O_3650,N_48452,N_49434);
and UO_3651 (O_3651,N_47884,N_47779);
nand UO_3652 (O_3652,N_48259,N_49342);
xor UO_3653 (O_3653,N_48456,N_49328);
or UO_3654 (O_3654,N_48683,N_48827);
nor UO_3655 (O_3655,N_49910,N_48393);
nor UO_3656 (O_3656,N_48139,N_49768);
or UO_3657 (O_3657,N_49426,N_48988);
nor UO_3658 (O_3658,N_47785,N_48968);
xor UO_3659 (O_3659,N_47848,N_49854);
nor UO_3660 (O_3660,N_48316,N_48155);
or UO_3661 (O_3661,N_48661,N_48850);
nor UO_3662 (O_3662,N_47801,N_47513);
or UO_3663 (O_3663,N_49408,N_48596);
xor UO_3664 (O_3664,N_48867,N_48407);
or UO_3665 (O_3665,N_48283,N_47806);
xnor UO_3666 (O_3666,N_47961,N_47559);
xnor UO_3667 (O_3667,N_47718,N_48683);
nor UO_3668 (O_3668,N_49066,N_48359);
and UO_3669 (O_3669,N_49874,N_47958);
xnor UO_3670 (O_3670,N_48424,N_49354);
nor UO_3671 (O_3671,N_48043,N_47782);
and UO_3672 (O_3672,N_47880,N_49821);
nand UO_3673 (O_3673,N_48961,N_48291);
nand UO_3674 (O_3674,N_49336,N_48215);
nand UO_3675 (O_3675,N_48338,N_49602);
or UO_3676 (O_3676,N_49943,N_48807);
or UO_3677 (O_3677,N_48003,N_49226);
or UO_3678 (O_3678,N_47967,N_49869);
nor UO_3679 (O_3679,N_47872,N_49547);
xnor UO_3680 (O_3680,N_49475,N_49519);
and UO_3681 (O_3681,N_49166,N_48024);
nor UO_3682 (O_3682,N_48451,N_48250);
xor UO_3683 (O_3683,N_48343,N_49500);
or UO_3684 (O_3684,N_48757,N_47880);
nand UO_3685 (O_3685,N_48860,N_48599);
nor UO_3686 (O_3686,N_49848,N_49008);
or UO_3687 (O_3687,N_48266,N_48448);
nor UO_3688 (O_3688,N_49658,N_47641);
nand UO_3689 (O_3689,N_48909,N_49899);
xor UO_3690 (O_3690,N_49778,N_49422);
or UO_3691 (O_3691,N_48636,N_48282);
or UO_3692 (O_3692,N_47745,N_49303);
nor UO_3693 (O_3693,N_49140,N_48876);
nand UO_3694 (O_3694,N_48396,N_49742);
nand UO_3695 (O_3695,N_48652,N_48063);
nor UO_3696 (O_3696,N_48452,N_48329);
xor UO_3697 (O_3697,N_49414,N_48729);
or UO_3698 (O_3698,N_47576,N_48413);
or UO_3699 (O_3699,N_49340,N_47792);
xor UO_3700 (O_3700,N_48044,N_47851);
and UO_3701 (O_3701,N_48933,N_47776);
nand UO_3702 (O_3702,N_49196,N_48299);
nor UO_3703 (O_3703,N_47525,N_49440);
or UO_3704 (O_3704,N_47794,N_49999);
nand UO_3705 (O_3705,N_49053,N_48890);
nand UO_3706 (O_3706,N_49447,N_48718);
and UO_3707 (O_3707,N_48317,N_49164);
or UO_3708 (O_3708,N_48157,N_49755);
nand UO_3709 (O_3709,N_49417,N_49154);
xnor UO_3710 (O_3710,N_48567,N_47849);
or UO_3711 (O_3711,N_49508,N_48982);
nor UO_3712 (O_3712,N_48468,N_49859);
nor UO_3713 (O_3713,N_48459,N_49148);
or UO_3714 (O_3714,N_49521,N_47746);
or UO_3715 (O_3715,N_47767,N_49731);
nand UO_3716 (O_3716,N_49491,N_48698);
and UO_3717 (O_3717,N_49811,N_48066);
nor UO_3718 (O_3718,N_49118,N_49648);
and UO_3719 (O_3719,N_48384,N_48607);
or UO_3720 (O_3720,N_47989,N_48226);
nand UO_3721 (O_3721,N_49203,N_49013);
xnor UO_3722 (O_3722,N_48678,N_49794);
nor UO_3723 (O_3723,N_49348,N_48753);
and UO_3724 (O_3724,N_49440,N_48940);
or UO_3725 (O_3725,N_48137,N_47931);
nand UO_3726 (O_3726,N_48395,N_47922);
nand UO_3727 (O_3727,N_48277,N_48188);
nand UO_3728 (O_3728,N_49126,N_48960);
nor UO_3729 (O_3729,N_48380,N_49346);
or UO_3730 (O_3730,N_48695,N_49322);
and UO_3731 (O_3731,N_47671,N_48139);
nor UO_3732 (O_3732,N_49618,N_49797);
nand UO_3733 (O_3733,N_49374,N_48237);
nand UO_3734 (O_3734,N_49308,N_48640);
nor UO_3735 (O_3735,N_48138,N_49018);
or UO_3736 (O_3736,N_49689,N_49076);
nand UO_3737 (O_3737,N_49956,N_48250);
xnor UO_3738 (O_3738,N_49408,N_49469);
nand UO_3739 (O_3739,N_49679,N_49158);
or UO_3740 (O_3740,N_49997,N_48553);
and UO_3741 (O_3741,N_49857,N_48989);
nand UO_3742 (O_3742,N_48930,N_48479);
xor UO_3743 (O_3743,N_49241,N_47678);
or UO_3744 (O_3744,N_47862,N_47524);
or UO_3745 (O_3745,N_47871,N_47836);
nand UO_3746 (O_3746,N_48039,N_49479);
nor UO_3747 (O_3747,N_48876,N_49965);
or UO_3748 (O_3748,N_47949,N_48323);
nand UO_3749 (O_3749,N_47596,N_49627);
or UO_3750 (O_3750,N_47939,N_47655);
xor UO_3751 (O_3751,N_49053,N_47821);
nand UO_3752 (O_3752,N_48895,N_49095);
nor UO_3753 (O_3753,N_48344,N_47829);
xnor UO_3754 (O_3754,N_48578,N_48302);
nor UO_3755 (O_3755,N_47625,N_49324);
nor UO_3756 (O_3756,N_49627,N_49964);
or UO_3757 (O_3757,N_47922,N_48628);
or UO_3758 (O_3758,N_49219,N_49282);
xor UO_3759 (O_3759,N_48003,N_48415);
and UO_3760 (O_3760,N_47949,N_48388);
and UO_3761 (O_3761,N_49628,N_47924);
nand UO_3762 (O_3762,N_49812,N_47660);
xor UO_3763 (O_3763,N_49927,N_49425);
and UO_3764 (O_3764,N_48886,N_49763);
nand UO_3765 (O_3765,N_48714,N_48018);
and UO_3766 (O_3766,N_47945,N_49722);
nand UO_3767 (O_3767,N_49345,N_49152);
and UO_3768 (O_3768,N_48631,N_48115);
nand UO_3769 (O_3769,N_49708,N_47611);
nor UO_3770 (O_3770,N_47781,N_49768);
nor UO_3771 (O_3771,N_49444,N_49795);
xnor UO_3772 (O_3772,N_49342,N_48087);
xnor UO_3773 (O_3773,N_48653,N_48151);
xor UO_3774 (O_3774,N_47612,N_49778);
nor UO_3775 (O_3775,N_49639,N_49475);
nor UO_3776 (O_3776,N_49662,N_49609);
or UO_3777 (O_3777,N_48027,N_49761);
or UO_3778 (O_3778,N_47526,N_49393);
or UO_3779 (O_3779,N_47765,N_48217);
and UO_3780 (O_3780,N_48290,N_48518);
and UO_3781 (O_3781,N_47612,N_48877);
or UO_3782 (O_3782,N_49960,N_49799);
xor UO_3783 (O_3783,N_48402,N_48351);
and UO_3784 (O_3784,N_48391,N_48265);
or UO_3785 (O_3785,N_49475,N_49587);
xor UO_3786 (O_3786,N_47574,N_49898);
xnor UO_3787 (O_3787,N_48788,N_48423);
xnor UO_3788 (O_3788,N_48532,N_48118);
nand UO_3789 (O_3789,N_48744,N_48483);
nor UO_3790 (O_3790,N_48682,N_47810);
nand UO_3791 (O_3791,N_49187,N_47866);
and UO_3792 (O_3792,N_49685,N_49850);
and UO_3793 (O_3793,N_47649,N_48585);
nand UO_3794 (O_3794,N_47880,N_48939);
and UO_3795 (O_3795,N_49980,N_49976);
nor UO_3796 (O_3796,N_49496,N_49225);
xor UO_3797 (O_3797,N_49074,N_49405);
and UO_3798 (O_3798,N_48284,N_49918);
xor UO_3799 (O_3799,N_49235,N_49693);
or UO_3800 (O_3800,N_49261,N_47905);
xnor UO_3801 (O_3801,N_49420,N_48168);
nand UO_3802 (O_3802,N_48757,N_48245);
and UO_3803 (O_3803,N_49057,N_48081);
and UO_3804 (O_3804,N_49990,N_47764);
or UO_3805 (O_3805,N_48944,N_48932);
xnor UO_3806 (O_3806,N_47879,N_49903);
and UO_3807 (O_3807,N_48809,N_49785);
nand UO_3808 (O_3808,N_49966,N_48155);
nand UO_3809 (O_3809,N_48694,N_48305);
and UO_3810 (O_3810,N_49916,N_48965);
and UO_3811 (O_3811,N_48715,N_49560);
and UO_3812 (O_3812,N_49532,N_47581);
nor UO_3813 (O_3813,N_48179,N_49779);
or UO_3814 (O_3814,N_48937,N_48476);
nor UO_3815 (O_3815,N_48683,N_48471);
nor UO_3816 (O_3816,N_48319,N_48135);
and UO_3817 (O_3817,N_49688,N_48693);
or UO_3818 (O_3818,N_49561,N_49709);
nor UO_3819 (O_3819,N_47929,N_48946);
nand UO_3820 (O_3820,N_49107,N_48438);
or UO_3821 (O_3821,N_49220,N_48439);
xor UO_3822 (O_3822,N_49735,N_47746);
nand UO_3823 (O_3823,N_47566,N_49215);
nor UO_3824 (O_3824,N_49132,N_47749);
nor UO_3825 (O_3825,N_48247,N_49176);
and UO_3826 (O_3826,N_47615,N_48722);
nand UO_3827 (O_3827,N_49586,N_49991);
nand UO_3828 (O_3828,N_47790,N_48150);
nand UO_3829 (O_3829,N_48361,N_48577);
and UO_3830 (O_3830,N_48630,N_48240);
and UO_3831 (O_3831,N_49150,N_48046);
or UO_3832 (O_3832,N_48389,N_49064);
xnor UO_3833 (O_3833,N_48731,N_48651);
nand UO_3834 (O_3834,N_47642,N_47570);
nor UO_3835 (O_3835,N_47780,N_49142);
or UO_3836 (O_3836,N_47949,N_47796);
nor UO_3837 (O_3837,N_48121,N_49185);
nor UO_3838 (O_3838,N_47798,N_48035);
xor UO_3839 (O_3839,N_47713,N_49837);
or UO_3840 (O_3840,N_48462,N_48425);
nor UO_3841 (O_3841,N_48938,N_48395);
xor UO_3842 (O_3842,N_49765,N_49044);
xor UO_3843 (O_3843,N_47815,N_48526);
nor UO_3844 (O_3844,N_48283,N_47530);
xor UO_3845 (O_3845,N_49345,N_49091);
nand UO_3846 (O_3846,N_49595,N_48812);
nand UO_3847 (O_3847,N_47571,N_49607);
nor UO_3848 (O_3848,N_49850,N_49144);
nor UO_3849 (O_3849,N_47788,N_49186);
nor UO_3850 (O_3850,N_47707,N_49479);
and UO_3851 (O_3851,N_47881,N_48842);
nor UO_3852 (O_3852,N_49202,N_49505);
xor UO_3853 (O_3853,N_48147,N_49439);
and UO_3854 (O_3854,N_47764,N_48524);
nor UO_3855 (O_3855,N_49481,N_48798);
and UO_3856 (O_3856,N_48943,N_47914);
xor UO_3857 (O_3857,N_49824,N_49033);
and UO_3858 (O_3858,N_48108,N_48396);
nand UO_3859 (O_3859,N_49190,N_49526);
and UO_3860 (O_3860,N_49560,N_48761);
nand UO_3861 (O_3861,N_48591,N_47897);
nand UO_3862 (O_3862,N_47793,N_47663);
nor UO_3863 (O_3863,N_48201,N_48918);
or UO_3864 (O_3864,N_47954,N_48399);
xor UO_3865 (O_3865,N_48445,N_48430);
and UO_3866 (O_3866,N_47764,N_48780);
or UO_3867 (O_3867,N_48692,N_48147);
nand UO_3868 (O_3868,N_48584,N_47537);
nand UO_3869 (O_3869,N_49276,N_48088);
nor UO_3870 (O_3870,N_48750,N_49741);
nor UO_3871 (O_3871,N_49169,N_47689);
and UO_3872 (O_3872,N_49841,N_48017);
and UO_3873 (O_3873,N_48242,N_48498);
and UO_3874 (O_3874,N_48074,N_47574);
or UO_3875 (O_3875,N_49199,N_49043);
xnor UO_3876 (O_3876,N_48664,N_48862);
nand UO_3877 (O_3877,N_48030,N_49455);
or UO_3878 (O_3878,N_48059,N_49771);
nor UO_3879 (O_3879,N_48630,N_47846);
xor UO_3880 (O_3880,N_49326,N_48553);
or UO_3881 (O_3881,N_49144,N_49596);
nor UO_3882 (O_3882,N_48969,N_49661);
or UO_3883 (O_3883,N_47659,N_48452);
or UO_3884 (O_3884,N_47843,N_49472);
or UO_3885 (O_3885,N_49983,N_49917);
and UO_3886 (O_3886,N_49890,N_49192);
nor UO_3887 (O_3887,N_49195,N_49798);
and UO_3888 (O_3888,N_47713,N_49857);
nor UO_3889 (O_3889,N_49083,N_49606);
nand UO_3890 (O_3890,N_48509,N_48042);
nor UO_3891 (O_3891,N_48219,N_49448);
nand UO_3892 (O_3892,N_48377,N_47999);
nor UO_3893 (O_3893,N_48158,N_48464);
xnor UO_3894 (O_3894,N_49060,N_49845);
nand UO_3895 (O_3895,N_49400,N_47700);
nand UO_3896 (O_3896,N_47725,N_49101);
or UO_3897 (O_3897,N_47554,N_49444);
nor UO_3898 (O_3898,N_49257,N_49048);
and UO_3899 (O_3899,N_48252,N_49663);
and UO_3900 (O_3900,N_47581,N_47862);
nor UO_3901 (O_3901,N_48876,N_47649);
xnor UO_3902 (O_3902,N_48951,N_47795);
and UO_3903 (O_3903,N_48532,N_49558);
nand UO_3904 (O_3904,N_49726,N_49979);
nor UO_3905 (O_3905,N_47699,N_48412);
and UO_3906 (O_3906,N_48819,N_48552);
and UO_3907 (O_3907,N_47516,N_49914);
or UO_3908 (O_3908,N_47530,N_48024);
nand UO_3909 (O_3909,N_48324,N_48649);
or UO_3910 (O_3910,N_48203,N_47566);
nand UO_3911 (O_3911,N_49225,N_48037);
or UO_3912 (O_3912,N_47966,N_48417);
nor UO_3913 (O_3913,N_49583,N_49973);
nand UO_3914 (O_3914,N_49175,N_49967);
or UO_3915 (O_3915,N_48461,N_48264);
nor UO_3916 (O_3916,N_48066,N_49771);
and UO_3917 (O_3917,N_48859,N_48191);
and UO_3918 (O_3918,N_49181,N_48539);
and UO_3919 (O_3919,N_48663,N_48415);
xor UO_3920 (O_3920,N_47515,N_48960);
or UO_3921 (O_3921,N_48019,N_48127);
and UO_3922 (O_3922,N_49414,N_48688);
xnor UO_3923 (O_3923,N_47561,N_49400);
nand UO_3924 (O_3924,N_48142,N_47668);
or UO_3925 (O_3925,N_48493,N_49684);
and UO_3926 (O_3926,N_47525,N_49484);
or UO_3927 (O_3927,N_48070,N_49049);
nor UO_3928 (O_3928,N_48735,N_48461);
nor UO_3929 (O_3929,N_48307,N_49156);
xor UO_3930 (O_3930,N_49648,N_49307);
nor UO_3931 (O_3931,N_49764,N_49327);
and UO_3932 (O_3932,N_49153,N_48235);
and UO_3933 (O_3933,N_49270,N_49981);
xnor UO_3934 (O_3934,N_48756,N_49840);
nand UO_3935 (O_3935,N_49079,N_49191);
nand UO_3936 (O_3936,N_49946,N_48507);
xor UO_3937 (O_3937,N_49988,N_49307);
or UO_3938 (O_3938,N_48563,N_49534);
nand UO_3939 (O_3939,N_47576,N_49691);
nand UO_3940 (O_3940,N_48410,N_48112);
nand UO_3941 (O_3941,N_47836,N_47856);
nor UO_3942 (O_3942,N_49685,N_47512);
and UO_3943 (O_3943,N_47785,N_47866);
and UO_3944 (O_3944,N_49908,N_48849);
and UO_3945 (O_3945,N_49492,N_49767);
nor UO_3946 (O_3946,N_47701,N_49708);
or UO_3947 (O_3947,N_49129,N_49324);
xor UO_3948 (O_3948,N_48598,N_49199);
xor UO_3949 (O_3949,N_49256,N_48474);
and UO_3950 (O_3950,N_48255,N_49008);
and UO_3951 (O_3951,N_48925,N_49159);
xnor UO_3952 (O_3952,N_49525,N_47823);
and UO_3953 (O_3953,N_49099,N_48459);
xnor UO_3954 (O_3954,N_47955,N_49019);
xor UO_3955 (O_3955,N_48706,N_48323);
and UO_3956 (O_3956,N_49436,N_49307);
or UO_3957 (O_3957,N_48133,N_49663);
or UO_3958 (O_3958,N_49619,N_49785);
nor UO_3959 (O_3959,N_48110,N_47919);
xor UO_3960 (O_3960,N_48740,N_49723);
or UO_3961 (O_3961,N_49452,N_49291);
and UO_3962 (O_3962,N_49078,N_48791);
nor UO_3963 (O_3963,N_48978,N_47553);
nor UO_3964 (O_3964,N_49289,N_47578);
and UO_3965 (O_3965,N_49913,N_47609);
and UO_3966 (O_3966,N_49194,N_49857);
and UO_3967 (O_3967,N_47750,N_49580);
and UO_3968 (O_3968,N_49365,N_48669);
nor UO_3969 (O_3969,N_48925,N_47921);
nor UO_3970 (O_3970,N_49004,N_47821);
nand UO_3971 (O_3971,N_49602,N_48003);
nor UO_3972 (O_3972,N_48627,N_49547);
nand UO_3973 (O_3973,N_49259,N_48420);
and UO_3974 (O_3974,N_48098,N_48669);
nand UO_3975 (O_3975,N_47722,N_49580);
nand UO_3976 (O_3976,N_48494,N_49515);
nor UO_3977 (O_3977,N_48352,N_47818);
nor UO_3978 (O_3978,N_47740,N_49163);
nand UO_3979 (O_3979,N_48926,N_48518);
xnor UO_3980 (O_3980,N_47866,N_49502);
nand UO_3981 (O_3981,N_48563,N_47722);
nor UO_3982 (O_3982,N_49504,N_49564);
and UO_3983 (O_3983,N_48602,N_49788);
nor UO_3984 (O_3984,N_48634,N_49213);
and UO_3985 (O_3985,N_48179,N_48253);
and UO_3986 (O_3986,N_49578,N_48154);
and UO_3987 (O_3987,N_49114,N_48085);
or UO_3988 (O_3988,N_49547,N_49982);
nor UO_3989 (O_3989,N_47822,N_47886);
nand UO_3990 (O_3990,N_49011,N_47594);
and UO_3991 (O_3991,N_48347,N_47744);
or UO_3992 (O_3992,N_48634,N_48431);
xor UO_3993 (O_3993,N_49533,N_47667);
and UO_3994 (O_3994,N_49285,N_47968);
and UO_3995 (O_3995,N_49681,N_49850);
nand UO_3996 (O_3996,N_48417,N_49491);
xor UO_3997 (O_3997,N_49815,N_49413);
or UO_3998 (O_3998,N_48235,N_48538);
and UO_3999 (O_3999,N_48524,N_49214);
or UO_4000 (O_4000,N_47638,N_49112);
or UO_4001 (O_4001,N_49332,N_48252);
xnor UO_4002 (O_4002,N_48204,N_48070);
and UO_4003 (O_4003,N_48470,N_49856);
and UO_4004 (O_4004,N_49059,N_48185);
nor UO_4005 (O_4005,N_49867,N_49300);
nand UO_4006 (O_4006,N_47859,N_47508);
or UO_4007 (O_4007,N_49855,N_48014);
xnor UO_4008 (O_4008,N_49278,N_48206);
and UO_4009 (O_4009,N_49246,N_49868);
nand UO_4010 (O_4010,N_48303,N_49636);
nor UO_4011 (O_4011,N_48097,N_49141);
or UO_4012 (O_4012,N_48023,N_49589);
or UO_4013 (O_4013,N_49548,N_47587);
nand UO_4014 (O_4014,N_48462,N_47856);
or UO_4015 (O_4015,N_49156,N_48528);
or UO_4016 (O_4016,N_49992,N_47952);
nor UO_4017 (O_4017,N_48590,N_48197);
nand UO_4018 (O_4018,N_48313,N_48122);
or UO_4019 (O_4019,N_48223,N_49414);
or UO_4020 (O_4020,N_48400,N_48334);
nand UO_4021 (O_4021,N_48390,N_48481);
or UO_4022 (O_4022,N_49148,N_47611);
nor UO_4023 (O_4023,N_48653,N_47838);
or UO_4024 (O_4024,N_47784,N_49854);
and UO_4025 (O_4025,N_48463,N_48383);
and UO_4026 (O_4026,N_49252,N_49358);
xor UO_4027 (O_4027,N_49596,N_47769);
nor UO_4028 (O_4028,N_47516,N_49354);
nor UO_4029 (O_4029,N_48385,N_47876);
nor UO_4030 (O_4030,N_49645,N_47863);
nor UO_4031 (O_4031,N_49674,N_47956);
nor UO_4032 (O_4032,N_47583,N_47717);
xor UO_4033 (O_4033,N_47910,N_47716);
xor UO_4034 (O_4034,N_48166,N_48962);
nand UO_4035 (O_4035,N_47774,N_47840);
nand UO_4036 (O_4036,N_47851,N_48384);
xor UO_4037 (O_4037,N_49743,N_49894);
nor UO_4038 (O_4038,N_48884,N_49965);
xor UO_4039 (O_4039,N_49453,N_49160);
xor UO_4040 (O_4040,N_47880,N_49855);
nor UO_4041 (O_4041,N_49759,N_47641);
nor UO_4042 (O_4042,N_47581,N_48540);
nor UO_4043 (O_4043,N_48851,N_48060);
nor UO_4044 (O_4044,N_49490,N_49690);
xor UO_4045 (O_4045,N_48218,N_49732);
nor UO_4046 (O_4046,N_49729,N_48241);
nand UO_4047 (O_4047,N_48283,N_48983);
and UO_4048 (O_4048,N_48308,N_47709);
and UO_4049 (O_4049,N_48714,N_47636);
and UO_4050 (O_4050,N_49449,N_48206);
nor UO_4051 (O_4051,N_47603,N_48610);
or UO_4052 (O_4052,N_49520,N_47804);
nor UO_4053 (O_4053,N_48617,N_48531);
nand UO_4054 (O_4054,N_47575,N_48267);
nor UO_4055 (O_4055,N_48638,N_47967);
and UO_4056 (O_4056,N_47717,N_49055);
or UO_4057 (O_4057,N_49267,N_49772);
and UO_4058 (O_4058,N_47524,N_49012);
xnor UO_4059 (O_4059,N_48694,N_49155);
or UO_4060 (O_4060,N_48058,N_47772);
nor UO_4061 (O_4061,N_48003,N_49144);
and UO_4062 (O_4062,N_48844,N_48123);
nor UO_4063 (O_4063,N_49978,N_48848);
or UO_4064 (O_4064,N_47658,N_48644);
xnor UO_4065 (O_4065,N_49856,N_48090);
and UO_4066 (O_4066,N_48588,N_48661);
nand UO_4067 (O_4067,N_49326,N_48077);
nand UO_4068 (O_4068,N_49110,N_49850);
and UO_4069 (O_4069,N_48218,N_49756);
nand UO_4070 (O_4070,N_49047,N_48489);
or UO_4071 (O_4071,N_49478,N_49055);
nand UO_4072 (O_4072,N_48002,N_48107);
or UO_4073 (O_4073,N_49079,N_48683);
nand UO_4074 (O_4074,N_48410,N_48418);
or UO_4075 (O_4075,N_48586,N_48853);
nand UO_4076 (O_4076,N_48868,N_49307);
and UO_4077 (O_4077,N_47722,N_48319);
xnor UO_4078 (O_4078,N_49849,N_49249);
and UO_4079 (O_4079,N_49282,N_47648);
nor UO_4080 (O_4080,N_48477,N_49555);
or UO_4081 (O_4081,N_47956,N_48654);
or UO_4082 (O_4082,N_48314,N_49210);
or UO_4083 (O_4083,N_48392,N_49333);
nand UO_4084 (O_4084,N_48348,N_49341);
xor UO_4085 (O_4085,N_48946,N_49398);
xnor UO_4086 (O_4086,N_48802,N_48408);
or UO_4087 (O_4087,N_48052,N_49124);
nand UO_4088 (O_4088,N_48073,N_47890);
or UO_4089 (O_4089,N_49220,N_47924);
and UO_4090 (O_4090,N_49665,N_49870);
or UO_4091 (O_4091,N_49316,N_49272);
nand UO_4092 (O_4092,N_49439,N_49572);
xor UO_4093 (O_4093,N_48120,N_49368);
nor UO_4094 (O_4094,N_48495,N_49388);
and UO_4095 (O_4095,N_47640,N_48565);
and UO_4096 (O_4096,N_49915,N_47785);
and UO_4097 (O_4097,N_48267,N_48881);
nor UO_4098 (O_4098,N_48601,N_49931);
and UO_4099 (O_4099,N_48662,N_49035);
and UO_4100 (O_4100,N_48764,N_49462);
or UO_4101 (O_4101,N_47966,N_48814);
nor UO_4102 (O_4102,N_49961,N_49643);
and UO_4103 (O_4103,N_47789,N_48802);
or UO_4104 (O_4104,N_49754,N_49712);
nor UO_4105 (O_4105,N_48809,N_48478);
xor UO_4106 (O_4106,N_49609,N_47650);
or UO_4107 (O_4107,N_49775,N_48020);
and UO_4108 (O_4108,N_47916,N_48860);
nand UO_4109 (O_4109,N_48579,N_48461);
nor UO_4110 (O_4110,N_48614,N_47978);
or UO_4111 (O_4111,N_48646,N_49723);
and UO_4112 (O_4112,N_47633,N_48402);
and UO_4113 (O_4113,N_47616,N_47961);
xnor UO_4114 (O_4114,N_48236,N_47815);
xnor UO_4115 (O_4115,N_48928,N_49326);
and UO_4116 (O_4116,N_49762,N_48528);
xor UO_4117 (O_4117,N_49882,N_49877);
and UO_4118 (O_4118,N_49140,N_47763);
xnor UO_4119 (O_4119,N_49897,N_47696);
nor UO_4120 (O_4120,N_49695,N_49170);
or UO_4121 (O_4121,N_48504,N_49904);
xnor UO_4122 (O_4122,N_49515,N_48764);
nor UO_4123 (O_4123,N_48330,N_49182);
xor UO_4124 (O_4124,N_48469,N_48968);
or UO_4125 (O_4125,N_49024,N_49633);
nand UO_4126 (O_4126,N_47958,N_49711);
and UO_4127 (O_4127,N_47594,N_47787);
and UO_4128 (O_4128,N_48511,N_48628);
and UO_4129 (O_4129,N_49057,N_48863);
xnor UO_4130 (O_4130,N_48610,N_49700);
and UO_4131 (O_4131,N_48146,N_48500);
or UO_4132 (O_4132,N_48737,N_49772);
xor UO_4133 (O_4133,N_49199,N_49209);
or UO_4134 (O_4134,N_47963,N_48244);
and UO_4135 (O_4135,N_48146,N_47892);
nand UO_4136 (O_4136,N_49773,N_49601);
nor UO_4137 (O_4137,N_47746,N_49571);
xnor UO_4138 (O_4138,N_48128,N_48287);
and UO_4139 (O_4139,N_48035,N_49098);
or UO_4140 (O_4140,N_47702,N_48555);
xor UO_4141 (O_4141,N_48736,N_49694);
nand UO_4142 (O_4142,N_47723,N_47764);
xnor UO_4143 (O_4143,N_47559,N_48039);
nand UO_4144 (O_4144,N_48442,N_48063);
or UO_4145 (O_4145,N_47538,N_48914);
xnor UO_4146 (O_4146,N_49035,N_48970);
and UO_4147 (O_4147,N_48259,N_47766);
nand UO_4148 (O_4148,N_49607,N_49765);
or UO_4149 (O_4149,N_48414,N_48754);
xor UO_4150 (O_4150,N_47552,N_49294);
xnor UO_4151 (O_4151,N_48265,N_47518);
nand UO_4152 (O_4152,N_49862,N_49845);
and UO_4153 (O_4153,N_49407,N_48830);
nand UO_4154 (O_4154,N_48764,N_47812);
and UO_4155 (O_4155,N_49392,N_48875);
or UO_4156 (O_4156,N_49180,N_49061);
xnor UO_4157 (O_4157,N_48192,N_48396);
or UO_4158 (O_4158,N_48983,N_47825);
or UO_4159 (O_4159,N_48984,N_47882);
nor UO_4160 (O_4160,N_49718,N_48236);
nor UO_4161 (O_4161,N_48734,N_47709);
and UO_4162 (O_4162,N_49006,N_48295);
or UO_4163 (O_4163,N_48544,N_48043);
nor UO_4164 (O_4164,N_48133,N_49201);
xnor UO_4165 (O_4165,N_48848,N_47975);
and UO_4166 (O_4166,N_49452,N_47998);
nand UO_4167 (O_4167,N_48727,N_48185);
nand UO_4168 (O_4168,N_48545,N_48554);
and UO_4169 (O_4169,N_48197,N_48694);
nand UO_4170 (O_4170,N_48488,N_48694);
xor UO_4171 (O_4171,N_49902,N_49339);
nand UO_4172 (O_4172,N_49823,N_48432);
xor UO_4173 (O_4173,N_48227,N_49157);
nor UO_4174 (O_4174,N_48422,N_48402);
nand UO_4175 (O_4175,N_49730,N_48348);
nand UO_4176 (O_4176,N_49907,N_49412);
and UO_4177 (O_4177,N_48134,N_49110);
or UO_4178 (O_4178,N_47903,N_48852);
nor UO_4179 (O_4179,N_49025,N_47930);
nand UO_4180 (O_4180,N_48866,N_48587);
nor UO_4181 (O_4181,N_47940,N_49743);
nor UO_4182 (O_4182,N_49852,N_49036);
xor UO_4183 (O_4183,N_48431,N_49763);
xnor UO_4184 (O_4184,N_47817,N_48555);
xor UO_4185 (O_4185,N_48733,N_48986);
xnor UO_4186 (O_4186,N_48123,N_48228);
nand UO_4187 (O_4187,N_48501,N_49049);
and UO_4188 (O_4188,N_48562,N_49967);
nand UO_4189 (O_4189,N_47945,N_48496);
nor UO_4190 (O_4190,N_48312,N_49690);
or UO_4191 (O_4191,N_48415,N_47545);
xnor UO_4192 (O_4192,N_47674,N_49246);
xor UO_4193 (O_4193,N_49266,N_48012);
or UO_4194 (O_4194,N_48230,N_47650);
nor UO_4195 (O_4195,N_48507,N_49097);
or UO_4196 (O_4196,N_49522,N_48791);
and UO_4197 (O_4197,N_49488,N_49543);
xor UO_4198 (O_4198,N_48199,N_49702);
nor UO_4199 (O_4199,N_48741,N_48125);
nor UO_4200 (O_4200,N_48839,N_47612);
nor UO_4201 (O_4201,N_48096,N_48018);
nand UO_4202 (O_4202,N_49674,N_48728);
nand UO_4203 (O_4203,N_49830,N_49879);
xor UO_4204 (O_4204,N_47920,N_49856);
and UO_4205 (O_4205,N_48110,N_48782);
nor UO_4206 (O_4206,N_49781,N_47971);
and UO_4207 (O_4207,N_48797,N_49989);
and UO_4208 (O_4208,N_47739,N_47712);
nand UO_4209 (O_4209,N_49725,N_48621);
xnor UO_4210 (O_4210,N_47732,N_48586);
and UO_4211 (O_4211,N_49436,N_49782);
and UO_4212 (O_4212,N_48463,N_48879);
nor UO_4213 (O_4213,N_48538,N_49264);
nor UO_4214 (O_4214,N_48948,N_49727);
or UO_4215 (O_4215,N_49147,N_47509);
or UO_4216 (O_4216,N_47975,N_48706);
xor UO_4217 (O_4217,N_48085,N_47680);
nor UO_4218 (O_4218,N_49032,N_49143);
xnor UO_4219 (O_4219,N_49694,N_48414);
or UO_4220 (O_4220,N_49288,N_47790);
and UO_4221 (O_4221,N_47614,N_47984);
nand UO_4222 (O_4222,N_48314,N_48837);
and UO_4223 (O_4223,N_48471,N_48264);
or UO_4224 (O_4224,N_49047,N_49215);
nor UO_4225 (O_4225,N_48605,N_48606);
nor UO_4226 (O_4226,N_48887,N_48494);
nor UO_4227 (O_4227,N_48277,N_48543);
nor UO_4228 (O_4228,N_47906,N_49260);
nand UO_4229 (O_4229,N_49514,N_47951);
and UO_4230 (O_4230,N_47599,N_47649);
xnor UO_4231 (O_4231,N_48389,N_48847);
and UO_4232 (O_4232,N_47512,N_47809);
nand UO_4233 (O_4233,N_49039,N_47616);
nand UO_4234 (O_4234,N_49408,N_48275);
or UO_4235 (O_4235,N_49225,N_48915);
nor UO_4236 (O_4236,N_49249,N_48613);
xnor UO_4237 (O_4237,N_49080,N_48958);
xnor UO_4238 (O_4238,N_48861,N_47936);
nor UO_4239 (O_4239,N_48114,N_48935);
or UO_4240 (O_4240,N_47773,N_47925);
nor UO_4241 (O_4241,N_49124,N_48516);
xnor UO_4242 (O_4242,N_49025,N_48211);
and UO_4243 (O_4243,N_47627,N_48837);
nand UO_4244 (O_4244,N_47581,N_48408);
nand UO_4245 (O_4245,N_49340,N_49467);
and UO_4246 (O_4246,N_47867,N_47520);
xor UO_4247 (O_4247,N_49452,N_49524);
nor UO_4248 (O_4248,N_48040,N_49825);
or UO_4249 (O_4249,N_49248,N_48223);
and UO_4250 (O_4250,N_48720,N_49955);
and UO_4251 (O_4251,N_48249,N_47961);
nor UO_4252 (O_4252,N_48795,N_48293);
or UO_4253 (O_4253,N_48423,N_48260);
nand UO_4254 (O_4254,N_48428,N_48208);
xor UO_4255 (O_4255,N_48122,N_49265);
and UO_4256 (O_4256,N_48879,N_48071);
and UO_4257 (O_4257,N_49070,N_48844);
nor UO_4258 (O_4258,N_47974,N_49386);
nand UO_4259 (O_4259,N_49794,N_49434);
nor UO_4260 (O_4260,N_47931,N_48504);
or UO_4261 (O_4261,N_47866,N_49172);
or UO_4262 (O_4262,N_49187,N_49988);
nor UO_4263 (O_4263,N_49984,N_49821);
nand UO_4264 (O_4264,N_48443,N_48513);
xor UO_4265 (O_4265,N_48049,N_47707);
nand UO_4266 (O_4266,N_48117,N_49425);
nand UO_4267 (O_4267,N_49065,N_48778);
nor UO_4268 (O_4268,N_48926,N_49625);
nor UO_4269 (O_4269,N_48883,N_47565);
nand UO_4270 (O_4270,N_48863,N_47896);
and UO_4271 (O_4271,N_49377,N_48681);
and UO_4272 (O_4272,N_49066,N_47930);
and UO_4273 (O_4273,N_47929,N_49966);
and UO_4274 (O_4274,N_48911,N_49229);
xor UO_4275 (O_4275,N_47734,N_49423);
or UO_4276 (O_4276,N_47922,N_49155);
nor UO_4277 (O_4277,N_48278,N_47740);
nor UO_4278 (O_4278,N_48225,N_48393);
nand UO_4279 (O_4279,N_48982,N_49075);
and UO_4280 (O_4280,N_47741,N_48984);
and UO_4281 (O_4281,N_49594,N_48303);
or UO_4282 (O_4282,N_49970,N_48915);
nand UO_4283 (O_4283,N_49044,N_47750);
xor UO_4284 (O_4284,N_48074,N_49824);
nand UO_4285 (O_4285,N_48287,N_49412);
or UO_4286 (O_4286,N_48658,N_48328);
and UO_4287 (O_4287,N_48013,N_48839);
nor UO_4288 (O_4288,N_49592,N_49398);
or UO_4289 (O_4289,N_49046,N_48317);
or UO_4290 (O_4290,N_49470,N_48468);
nand UO_4291 (O_4291,N_48006,N_48670);
xnor UO_4292 (O_4292,N_47572,N_47605);
xnor UO_4293 (O_4293,N_47602,N_48014);
xnor UO_4294 (O_4294,N_48717,N_49441);
and UO_4295 (O_4295,N_49899,N_47753);
nand UO_4296 (O_4296,N_47741,N_48631);
nor UO_4297 (O_4297,N_49808,N_49734);
and UO_4298 (O_4298,N_49351,N_47882);
nand UO_4299 (O_4299,N_49543,N_48323);
nand UO_4300 (O_4300,N_48670,N_48220);
nand UO_4301 (O_4301,N_48409,N_48917);
nor UO_4302 (O_4302,N_49082,N_47573);
or UO_4303 (O_4303,N_48295,N_48813);
nand UO_4304 (O_4304,N_48364,N_47754);
or UO_4305 (O_4305,N_49313,N_48220);
xor UO_4306 (O_4306,N_49468,N_48030);
or UO_4307 (O_4307,N_48701,N_48280);
and UO_4308 (O_4308,N_49008,N_48090);
nand UO_4309 (O_4309,N_48163,N_48310);
nand UO_4310 (O_4310,N_49786,N_47986);
or UO_4311 (O_4311,N_49440,N_49644);
and UO_4312 (O_4312,N_48246,N_49706);
xnor UO_4313 (O_4313,N_47538,N_48061);
or UO_4314 (O_4314,N_49776,N_48840);
nand UO_4315 (O_4315,N_48072,N_47794);
or UO_4316 (O_4316,N_49036,N_48748);
nor UO_4317 (O_4317,N_49540,N_49211);
and UO_4318 (O_4318,N_48176,N_47690);
and UO_4319 (O_4319,N_48692,N_48076);
nand UO_4320 (O_4320,N_49735,N_48357);
and UO_4321 (O_4321,N_48512,N_49517);
and UO_4322 (O_4322,N_49264,N_48574);
nand UO_4323 (O_4323,N_47910,N_48829);
or UO_4324 (O_4324,N_48323,N_48956);
nor UO_4325 (O_4325,N_49948,N_49644);
nor UO_4326 (O_4326,N_47676,N_48604);
and UO_4327 (O_4327,N_48186,N_49323);
xor UO_4328 (O_4328,N_49895,N_49789);
and UO_4329 (O_4329,N_49268,N_48458);
and UO_4330 (O_4330,N_49656,N_49536);
nor UO_4331 (O_4331,N_48843,N_48181);
and UO_4332 (O_4332,N_48473,N_49742);
and UO_4333 (O_4333,N_47993,N_48176);
and UO_4334 (O_4334,N_49010,N_48034);
xor UO_4335 (O_4335,N_49302,N_47827);
nand UO_4336 (O_4336,N_49833,N_48225);
nand UO_4337 (O_4337,N_49475,N_48394);
xnor UO_4338 (O_4338,N_49211,N_48403);
xnor UO_4339 (O_4339,N_49379,N_49625);
nand UO_4340 (O_4340,N_49077,N_48678);
nor UO_4341 (O_4341,N_48281,N_48929);
xnor UO_4342 (O_4342,N_47697,N_49590);
nand UO_4343 (O_4343,N_47709,N_49451);
nor UO_4344 (O_4344,N_48044,N_48342);
nor UO_4345 (O_4345,N_48243,N_49622);
nor UO_4346 (O_4346,N_48834,N_49851);
nand UO_4347 (O_4347,N_47934,N_48398);
xnor UO_4348 (O_4348,N_48538,N_48097);
nor UO_4349 (O_4349,N_49581,N_47556);
nor UO_4350 (O_4350,N_49710,N_49986);
xor UO_4351 (O_4351,N_48437,N_49009);
nor UO_4352 (O_4352,N_49390,N_49918);
nand UO_4353 (O_4353,N_48715,N_48696);
nor UO_4354 (O_4354,N_48542,N_48733);
nand UO_4355 (O_4355,N_47836,N_49617);
nand UO_4356 (O_4356,N_47613,N_47975);
and UO_4357 (O_4357,N_49353,N_48846);
nor UO_4358 (O_4358,N_48466,N_48955);
and UO_4359 (O_4359,N_49421,N_47676);
nor UO_4360 (O_4360,N_49785,N_48594);
nand UO_4361 (O_4361,N_48070,N_48104);
xor UO_4362 (O_4362,N_49956,N_48446);
or UO_4363 (O_4363,N_48010,N_49206);
xor UO_4364 (O_4364,N_47835,N_49660);
nand UO_4365 (O_4365,N_47640,N_49837);
xnor UO_4366 (O_4366,N_47704,N_48333);
nor UO_4367 (O_4367,N_49131,N_49414);
nor UO_4368 (O_4368,N_49199,N_47533);
nand UO_4369 (O_4369,N_49493,N_48473);
or UO_4370 (O_4370,N_48495,N_49718);
nor UO_4371 (O_4371,N_47700,N_49857);
and UO_4372 (O_4372,N_47819,N_48342);
and UO_4373 (O_4373,N_48502,N_48449);
and UO_4374 (O_4374,N_48532,N_49128);
or UO_4375 (O_4375,N_48970,N_49776);
or UO_4376 (O_4376,N_48743,N_49123);
or UO_4377 (O_4377,N_49517,N_47638);
nand UO_4378 (O_4378,N_48972,N_47658);
nor UO_4379 (O_4379,N_49483,N_49450);
xnor UO_4380 (O_4380,N_48456,N_48513);
xnor UO_4381 (O_4381,N_48618,N_49649);
or UO_4382 (O_4382,N_48618,N_48294);
xor UO_4383 (O_4383,N_49984,N_49705);
xnor UO_4384 (O_4384,N_49356,N_48869);
or UO_4385 (O_4385,N_48485,N_48039);
and UO_4386 (O_4386,N_47751,N_49733);
or UO_4387 (O_4387,N_49158,N_49116);
nor UO_4388 (O_4388,N_47935,N_49872);
xnor UO_4389 (O_4389,N_48049,N_47843);
nor UO_4390 (O_4390,N_49580,N_47626);
nor UO_4391 (O_4391,N_49151,N_48527);
nor UO_4392 (O_4392,N_48271,N_49000);
or UO_4393 (O_4393,N_48813,N_47832);
or UO_4394 (O_4394,N_47528,N_48400);
nor UO_4395 (O_4395,N_49147,N_49595);
nor UO_4396 (O_4396,N_49143,N_48814);
xnor UO_4397 (O_4397,N_49827,N_48602);
nand UO_4398 (O_4398,N_47734,N_49219);
nand UO_4399 (O_4399,N_49278,N_47890);
xnor UO_4400 (O_4400,N_48330,N_47583);
and UO_4401 (O_4401,N_48993,N_47651);
or UO_4402 (O_4402,N_49128,N_48125);
nand UO_4403 (O_4403,N_47676,N_49153);
and UO_4404 (O_4404,N_48804,N_48362);
or UO_4405 (O_4405,N_48348,N_49194);
or UO_4406 (O_4406,N_49591,N_49190);
or UO_4407 (O_4407,N_48180,N_47780);
or UO_4408 (O_4408,N_49545,N_48812);
nand UO_4409 (O_4409,N_49676,N_48848);
nor UO_4410 (O_4410,N_48870,N_47550);
xnor UO_4411 (O_4411,N_49909,N_49014);
nand UO_4412 (O_4412,N_48719,N_48342);
nor UO_4413 (O_4413,N_48032,N_48764);
nor UO_4414 (O_4414,N_47714,N_48732);
xor UO_4415 (O_4415,N_47828,N_48544);
xor UO_4416 (O_4416,N_47728,N_47833);
nand UO_4417 (O_4417,N_49152,N_49565);
nor UO_4418 (O_4418,N_49002,N_47809);
xnor UO_4419 (O_4419,N_49688,N_47855);
xnor UO_4420 (O_4420,N_49120,N_48838);
nand UO_4421 (O_4421,N_48870,N_48952);
and UO_4422 (O_4422,N_48085,N_48551);
or UO_4423 (O_4423,N_48847,N_49722);
nor UO_4424 (O_4424,N_48714,N_49284);
or UO_4425 (O_4425,N_49105,N_49533);
nand UO_4426 (O_4426,N_47978,N_48976);
or UO_4427 (O_4427,N_47534,N_48530);
nor UO_4428 (O_4428,N_48483,N_47614);
nor UO_4429 (O_4429,N_49893,N_49789);
and UO_4430 (O_4430,N_49546,N_49544);
nand UO_4431 (O_4431,N_48538,N_49675);
and UO_4432 (O_4432,N_48846,N_47516);
or UO_4433 (O_4433,N_49347,N_48632);
xnor UO_4434 (O_4434,N_47944,N_49056);
nor UO_4435 (O_4435,N_49420,N_48883);
nand UO_4436 (O_4436,N_47736,N_49275);
xor UO_4437 (O_4437,N_49414,N_48538);
nor UO_4438 (O_4438,N_49809,N_47701);
nand UO_4439 (O_4439,N_47904,N_48198);
xnor UO_4440 (O_4440,N_48285,N_48570);
or UO_4441 (O_4441,N_48513,N_49484);
and UO_4442 (O_4442,N_48130,N_49374);
or UO_4443 (O_4443,N_48569,N_47737);
nor UO_4444 (O_4444,N_48672,N_47737);
nand UO_4445 (O_4445,N_48355,N_49466);
nor UO_4446 (O_4446,N_48141,N_48550);
xnor UO_4447 (O_4447,N_49584,N_49960);
nand UO_4448 (O_4448,N_49011,N_48936);
xor UO_4449 (O_4449,N_49157,N_47517);
nand UO_4450 (O_4450,N_49724,N_48946);
nor UO_4451 (O_4451,N_47636,N_49875);
nor UO_4452 (O_4452,N_49634,N_48356);
xor UO_4453 (O_4453,N_47749,N_49696);
or UO_4454 (O_4454,N_49707,N_48967);
or UO_4455 (O_4455,N_48731,N_48865);
xnor UO_4456 (O_4456,N_47948,N_47630);
nand UO_4457 (O_4457,N_48401,N_49294);
nor UO_4458 (O_4458,N_49082,N_49829);
or UO_4459 (O_4459,N_47759,N_49774);
and UO_4460 (O_4460,N_48379,N_48719);
nor UO_4461 (O_4461,N_48180,N_48702);
or UO_4462 (O_4462,N_49633,N_48398);
nand UO_4463 (O_4463,N_48829,N_48702);
and UO_4464 (O_4464,N_47677,N_47567);
or UO_4465 (O_4465,N_48535,N_48695);
and UO_4466 (O_4466,N_49213,N_48806);
xor UO_4467 (O_4467,N_47575,N_48438);
and UO_4468 (O_4468,N_49253,N_49601);
or UO_4469 (O_4469,N_47999,N_48432);
nand UO_4470 (O_4470,N_49500,N_47561);
nor UO_4471 (O_4471,N_48233,N_48790);
or UO_4472 (O_4472,N_48480,N_47991);
or UO_4473 (O_4473,N_49918,N_47619);
xor UO_4474 (O_4474,N_48622,N_49732);
xor UO_4475 (O_4475,N_49197,N_49781);
nor UO_4476 (O_4476,N_49167,N_48411);
and UO_4477 (O_4477,N_49652,N_47555);
and UO_4478 (O_4478,N_48069,N_49453);
nand UO_4479 (O_4479,N_48675,N_48922);
nand UO_4480 (O_4480,N_48057,N_47732);
nor UO_4481 (O_4481,N_49449,N_47504);
and UO_4482 (O_4482,N_48081,N_48532);
xnor UO_4483 (O_4483,N_48863,N_48956);
nor UO_4484 (O_4484,N_48136,N_48305);
and UO_4485 (O_4485,N_48957,N_49379);
and UO_4486 (O_4486,N_49753,N_49796);
xnor UO_4487 (O_4487,N_49297,N_48013);
nor UO_4488 (O_4488,N_49628,N_48570);
and UO_4489 (O_4489,N_49848,N_48167);
xor UO_4490 (O_4490,N_48084,N_47681);
nand UO_4491 (O_4491,N_48234,N_48046);
or UO_4492 (O_4492,N_48123,N_48907);
nor UO_4493 (O_4493,N_47628,N_48517);
or UO_4494 (O_4494,N_49262,N_48112);
nor UO_4495 (O_4495,N_49469,N_47690);
nand UO_4496 (O_4496,N_49602,N_48358);
nor UO_4497 (O_4497,N_49404,N_48940);
nor UO_4498 (O_4498,N_49444,N_49063);
and UO_4499 (O_4499,N_49422,N_49554);
and UO_4500 (O_4500,N_48354,N_48937);
and UO_4501 (O_4501,N_47860,N_49356);
and UO_4502 (O_4502,N_49003,N_47525);
or UO_4503 (O_4503,N_47796,N_49816);
nand UO_4504 (O_4504,N_49138,N_47902);
nor UO_4505 (O_4505,N_48651,N_48778);
nor UO_4506 (O_4506,N_48509,N_49268);
nand UO_4507 (O_4507,N_49255,N_49771);
nand UO_4508 (O_4508,N_49972,N_48449);
and UO_4509 (O_4509,N_48707,N_48419);
nand UO_4510 (O_4510,N_49666,N_47550);
or UO_4511 (O_4511,N_48197,N_49181);
or UO_4512 (O_4512,N_49698,N_49982);
nand UO_4513 (O_4513,N_47582,N_49495);
nand UO_4514 (O_4514,N_49835,N_48779);
and UO_4515 (O_4515,N_49101,N_47546);
xor UO_4516 (O_4516,N_47658,N_48389);
and UO_4517 (O_4517,N_48392,N_48850);
nor UO_4518 (O_4518,N_49339,N_48752);
and UO_4519 (O_4519,N_48011,N_48410);
and UO_4520 (O_4520,N_47795,N_47513);
xor UO_4521 (O_4521,N_48721,N_49739);
xor UO_4522 (O_4522,N_48276,N_48688);
nand UO_4523 (O_4523,N_49717,N_49583);
and UO_4524 (O_4524,N_47992,N_49991);
nand UO_4525 (O_4525,N_49345,N_49228);
nand UO_4526 (O_4526,N_47564,N_49143);
or UO_4527 (O_4527,N_48731,N_48926);
nor UO_4528 (O_4528,N_48631,N_47753);
and UO_4529 (O_4529,N_48439,N_48168);
and UO_4530 (O_4530,N_49001,N_49040);
xor UO_4531 (O_4531,N_48496,N_48781);
or UO_4532 (O_4532,N_48250,N_49057);
nor UO_4533 (O_4533,N_48382,N_48605);
or UO_4534 (O_4534,N_48822,N_49074);
nor UO_4535 (O_4535,N_48422,N_49375);
or UO_4536 (O_4536,N_48219,N_48164);
or UO_4537 (O_4537,N_49088,N_49007);
xor UO_4538 (O_4538,N_49950,N_49051);
nor UO_4539 (O_4539,N_48237,N_48584);
xnor UO_4540 (O_4540,N_49545,N_49592);
xnor UO_4541 (O_4541,N_49870,N_49513);
nor UO_4542 (O_4542,N_49060,N_48128);
or UO_4543 (O_4543,N_48784,N_48214);
or UO_4544 (O_4544,N_49982,N_48288);
nor UO_4545 (O_4545,N_49612,N_49593);
nand UO_4546 (O_4546,N_49576,N_49630);
nor UO_4547 (O_4547,N_48923,N_49501);
nand UO_4548 (O_4548,N_48529,N_49416);
or UO_4549 (O_4549,N_48452,N_49666);
nand UO_4550 (O_4550,N_49898,N_49941);
nor UO_4551 (O_4551,N_48281,N_47531);
nor UO_4552 (O_4552,N_49221,N_47805);
xnor UO_4553 (O_4553,N_49201,N_49136);
xnor UO_4554 (O_4554,N_48985,N_48850);
nand UO_4555 (O_4555,N_49161,N_49536);
and UO_4556 (O_4556,N_47542,N_49217);
nand UO_4557 (O_4557,N_49791,N_49290);
nand UO_4558 (O_4558,N_48730,N_47769);
and UO_4559 (O_4559,N_48264,N_48646);
or UO_4560 (O_4560,N_48470,N_48100);
nand UO_4561 (O_4561,N_49600,N_49988);
and UO_4562 (O_4562,N_48560,N_48767);
nand UO_4563 (O_4563,N_48688,N_48224);
or UO_4564 (O_4564,N_48141,N_49071);
and UO_4565 (O_4565,N_49242,N_48756);
nand UO_4566 (O_4566,N_47847,N_49295);
and UO_4567 (O_4567,N_47819,N_48618);
or UO_4568 (O_4568,N_49083,N_49460);
and UO_4569 (O_4569,N_48243,N_48072);
xor UO_4570 (O_4570,N_47592,N_49012);
nand UO_4571 (O_4571,N_49014,N_49411);
or UO_4572 (O_4572,N_47934,N_49749);
or UO_4573 (O_4573,N_49565,N_49405);
nand UO_4574 (O_4574,N_49258,N_49112);
or UO_4575 (O_4575,N_48098,N_48833);
and UO_4576 (O_4576,N_47825,N_47795);
and UO_4577 (O_4577,N_47838,N_49988);
or UO_4578 (O_4578,N_48796,N_49416);
and UO_4579 (O_4579,N_48760,N_47700);
xnor UO_4580 (O_4580,N_48530,N_48135);
nor UO_4581 (O_4581,N_47677,N_48817);
or UO_4582 (O_4582,N_47719,N_49851);
xor UO_4583 (O_4583,N_48867,N_49512);
and UO_4584 (O_4584,N_49203,N_47560);
xor UO_4585 (O_4585,N_47621,N_49758);
nand UO_4586 (O_4586,N_49608,N_49046);
nor UO_4587 (O_4587,N_49490,N_48796);
or UO_4588 (O_4588,N_48865,N_49511);
and UO_4589 (O_4589,N_48838,N_49999);
nor UO_4590 (O_4590,N_49850,N_49204);
and UO_4591 (O_4591,N_48724,N_47973);
nor UO_4592 (O_4592,N_48335,N_49579);
nor UO_4593 (O_4593,N_48927,N_48175);
xor UO_4594 (O_4594,N_48987,N_49857);
xor UO_4595 (O_4595,N_49204,N_49206);
nand UO_4596 (O_4596,N_48743,N_48109);
nor UO_4597 (O_4597,N_49290,N_47565);
nor UO_4598 (O_4598,N_47965,N_49794);
xnor UO_4599 (O_4599,N_48254,N_49660);
xnor UO_4600 (O_4600,N_48793,N_48414);
or UO_4601 (O_4601,N_48302,N_47980);
or UO_4602 (O_4602,N_47990,N_49666);
nor UO_4603 (O_4603,N_48369,N_49260);
and UO_4604 (O_4604,N_49441,N_49756);
nand UO_4605 (O_4605,N_48651,N_48700);
nor UO_4606 (O_4606,N_49119,N_47873);
xnor UO_4607 (O_4607,N_48644,N_48698);
and UO_4608 (O_4608,N_47529,N_47910);
xnor UO_4609 (O_4609,N_47706,N_49807);
nand UO_4610 (O_4610,N_47674,N_49629);
or UO_4611 (O_4611,N_49655,N_48548);
and UO_4612 (O_4612,N_48835,N_48761);
xnor UO_4613 (O_4613,N_47999,N_48009);
and UO_4614 (O_4614,N_47524,N_48556);
xor UO_4615 (O_4615,N_49246,N_48553);
and UO_4616 (O_4616,N_48123,N_47607);
nand UO_4617 (O_4617,N_47639,N_49022);
xnor UO_4618 (O_4618,N_47946,N_49931);
nor UO_4619 (O_4619,N_49585,N_49693);
nor UO_4620 (O_4620,N_48141,N_47982);
nor UO_4621 (O_4621,N_48606,N_48710);
nor UO_4622 (O_4622,N_47949,N_48457);
nor UO_4623 (O_4623,N_49914,N_47961);
or UO_4624 (O_4624,N_49925,N_49459);
and UO_4625 (O_4625,N_48353,N_48479);
and UO_4626 (O_4626,N_47511,N_47958);
xnor UO_4627 (O_4627,N_48402,N_48875);
or UO_4628 (O_4628,N_48360,N_48779);
nor UO_4629 (O_4629,N_48742,N_49249);
nor UO_4630 (O_4630,N_49626,N_48751);
xor UO_4631 (O_4631,N_48068,N_49484);
or UO_4632 (O_4632,N_49870,N_48435);
nor UO_4633 (O_4633,N_49771,N_48432);
or UO_4634 (O_4634,N_48657,N_48212);
and UO_4635 (O_4635,N_49960,N_49742);
and UO_4636 (O_4636,N_49734,N_47823);
or UO_4637 (O_4637,N_48022,N_48361);
or UO_4638 (O_4638,N_49834,N_48393);
nor UO_4639 (O_4639,N_49900,N_47712);
or UO_4640 (O_4640,N_48195,N_47740);
nor UO_4641 (O_4641,N_48768,N_48817);
nor UO_4642 (O_4642,N_49601,N_49369);
or UO_4643 (O_4643,N_48540,N_49551);
or UO_4644 (O_4644,N_48995,N_49003);
xor UO_4645 (O_4645,N_49860,N_48353);
xor UO_4646 (O_4646,N_49974,N_48641);
nand UO_4647 (O_4647,N_49767,N_49114);
or UO_4648 (O_4648,N_49828,N_49282);
or UO_4649 (O_4649,N_48404,N_49275);
or UO_4650 (O_4650,N_48369,N_48961);
nor UO_4651 (O_4651,N_49593,N_47997);
or UO_4652 (O_4652,N_48201,N_48639);
and UO_4653 (O_4653,N_48034,N_47884);
or UO_4654 (O_4654,N_48693,N_48060);
nand UO_4655 (O_4655,N_48861,N_48538);
nand UO_4656 (O_4656,N_49839,N_47558);
nand UO_4657 (O_4657,N_48003,N_48735);
xor UO_4658 (O_4658,N_49718,N_48187);
and UO_4659 (O_4659,N_47801,N_48580);
or UO_4660 (O_4660,N_48445,N_49255);
or UO_4661 (O_4661,N_48713,N_48734);
and UO_4662 (O_4662,N_47984,N_49287);
xnor UO_4663 (O_4663,N_49876,N_47643);
xnor UO_4664 (O_4664,N_47976,N_49562);
xor UO_4665 (O_4665,N_48760,N_49972);
nand UO_4666 (O_4666,N_47811,N_48039);
xnor UO_4667 (O_4667,N_48657,N_48367);
nand UO_4668 (O_4668,N_48695,N_49178);
nand UO_4669 (O_4669,N_49138,N_48225);
or UO_4670 (O_4670,N_49531,N_49524);
or UO_4671 (O_4671,N_48508,N_47504);
nand UO_4672 (O_4672,N_48303,N_49868);
nand UO_4673 (O_4673,N_49722,N_49238);
nand UO_4674 (O_4674,N_48951,N_48459);
nor UO_4675 (O_4675,N_47623,N_49329);
and UO_4676 (O_4676,N_49495,N_48369);
xnor UO_4677 (O_4677,N_48777,N_49079);
xor UO_4678 (O_4678,N_48610,N_49006);
or UO_4679 (O_4679,N_48597,N_49983);
or UO_4680 (O_4680,N_49590,N_47990);
nor UO_4681 (O_4681,N_48966,N_49735);
and UO_4682 (O_4682,N_49951,N_48780);
nor UO_4683 (O_4683,N_49006,N_48588);
xnor UO_4684 (O_4684,N_49576,N_49542);
xor UO_4685 (O_4685,N_47921,N_48329);
and UO_4686 (O_4686,N_48165,N_47987);
nand UO_4687 (O_4687,N_49097,N_47626);
nor UO_4688 (O_4688,N_48991,N_48978);
and UO_4689 (O_4689,N_47571,N_48579);
nor UO_4690 (O_4690,N_47867,N_48819);
or UO_4691 (O_4691,N_49304,N_48270);
nor UO_4692 (O_4692,N_47790,N_48320);
and UO_4693 (O_4693,N_48989,N_48146);
nor UO_4694 (O_4694,N_48871,N_49370);
or UO_4695 (O_4695,N_47951,N_48638);
and UO_4696 (O_4696,N_49371,N_48993);
or UO_4697 (O_4697,N_49982,N_49719);
and UO_4698 (O_4698,N_49590,N_49075);
and UO_4699 (O_4699,N_48561,N_49365);
nand UO_4700 (O_4700,N_47924,N_47876);
or UO_4701 (O_4701,N_48956,N_47673);
or UO_4702 (O_4702,N_47692,N_49331);
or UO_4703 (O_4703,N_48353,N_48755);
and UO_4704 (O_4704,N_48121,N_48991);
and UO_4705 (O_4705,N_48080,N_49033);
nand UO_4706 (O_4706,N_49417,N_47503);
nand UO_4707 (O_4707,N_48802,N_49277);
or UO_4708 (O_4708,N_48749,N_48025);
and UO_4709 (O_4709,N_49044,N_48680);
nor UO_4710 (O_4710,N_48184,N_48608);
nand UO_4711 (O_4711,N_49068,N_49537);
nor UO_4712 (O_4712,N_49363,N_49904);
nand UO_4713 (O_4713,N_47768,N_47798);
and UO_4714 (O_4714,N_49756,N_49138);
nor UO_4715 (O_4715,N_47998,N_48472);
xnor UO_4716 (O_4716,N_48405,N_48679);
nand UO_4717 (O_4717,N_49640,N_49852);
nor UO_4718 (O_4718,N_49133,N_48842);
nand UO_4719 (O_4719,N_48164,N_48872);
nand UO_4720 (O_4720,N_47755,N_48036);
nand UO_4721 (O_4721,N_49079,N_48979);
nor UO_4722 (O_4722,N_49393,N_48019);
and UO_4723 (O_4723,N_48559,N_47918);
nor UO_4724 (O_4724,N_49555,N_48090);
nor UO_4725 (O_4725,N_49881,N_49019);
nand UO_4726 (O_4726,N_47620,N_49376);
xnor UO_4727 (O_4727,N_48663,N_48769);
xnor UO_4728 (O_4728,N_49353,N_49750);
or UO_4729 (O_4729,N_49318,N_48663);
xor UO_4730 (O_4730,N_48871,N_49074);
nand UO_4731 (O_4731,N_49895,N_49338);
nor UO_4732 (O_4732,N_47757,N_47789);
xor UO_4733 (O_4733,N_49447,N_49750);
or UO_4734 (O_4734,N_48500,N_49136);
and UO_4735 (O_4735,N_48288,N_48874);
and UO_4736 (O_4736,N_49367,N_47843);
nand UO_4737 (O_4737,N_49102,N_49908);
or UO_4738 (O_4738,N_48500,N_49284);
nor UO_4739 (O_4739,N_47756,N_48654);
or UO_4740 (O_4740,N_47827,N_49959);
and UO_4741 (O_4741,N_48833,N_49083);
nor UO_4742 (O_4742,N_47931,N_48361);
xor UO_4743 (O_4743,N_48386,N_49962);
and UO_4744 (O_4744,N_49006,N_48560);
nor UO_4745 (O_4745,N_49150,N_47736);
xor UO_4746 (O_4746,N_48306,N_48076);
xnor UO_4747 (O_4747,N_49204,N_48488);
xor UO_4748 (O_4748,N_49852,N_48477);
and UO_4749 (O_4749,N_47904,N_49825);
xnor UO_4750 (O_4750,N_48008,N_49342);
nand UO_4751 (O_4751,N_47903,N_48284);
nor UO_4752 (O_4752,N_47614,N_49793);
xor UO_4753 (O_4753,N_49960,N_49592);
nor UO_4754 (O_4754,N_48575,N_49674);
nand UO_4755 (O_4755,N_48925,N_48975);
nor UO_4756 (O_4756,N_49140,N_48229);
and UO_4757 (O_4757,N_48199,N_48974);
nand UO_4758 (O_4758,N_47669,N_47627);
xnor UO_4759 (O_4759,N_49587,N_49665);
nor UO_4760 (O_4760,N_47878,N_47682);
xnor UO_4761 (O_4761,N_49331,N_48429);
and UO_4762 (O_4762,N_49055,N_49329);
or UO_4763 (O_4763,N_49895,N_48118);
xor UO_4764 (O_4764,N_48435,N_48174);
nand UO_4765 (O_4765,N_48090,N_48448);
or UO_4766 (O_4766,N_48495,N_47639);
xnor UO_4767 (O_4767,N_47971,N_48024);
xnor UO_4768 (O_4768,N_47951,N_48954);
nand UO_4769 (O_4769,N_49486,N_48911);
and UO_4770 (O_4770,N_49849,N_49566);
xnor UO_4771 (O_4771,N_49357,N_47683);
or UO_4772 (O_4772,N_47694,N_49814);
xor UO_4773 (O_4773,N_48239,N_49644);
and UO_4774 (O_4774,N_47940,N_48100);
or UO_4775 (O_4775,N_49822,N_47651);
or UO_4776 (O_4776,N_47910,N_47633);
and UO_4777 (O_4777,N_49704,N_48695);
nand UO_4778 (O_4778,N_47760,N_48220);
and UO_4779 (O_4779,N_48707,N_49110);
xnor UO_4780 (O_4780,N_47777,N_48728);
xor UO_4781 (O_4781,N_47926,N_48985);
and UO_4782 (O_4782,N_49193,N_48362);
or UO_4783 (O_4783,N_48301,N_47525);
nand UO_4784 (O_4784,N_48930,N_47680);
nor UO_4785 (O_4785,N_49384,N_48752);
and UO_4786 (O_4786,N_48938,N_48062);
or UO_4787 (O_4787,N_48190,N_47742);
nand UO_4788 (O_4788,N_49337,N_47918);
nand UO_4789 (O_4789,N_49492,N_49594);
and UO_4790 (O_4790,N_48803,N_47902);
and UO_4791 (O_4791,N_49070,N_48498);
nor UO_4792 (O_4792,N_47633,N_49583);
and UO_4793 (O_4793,N_47947,N_47602);
xnor UO_4794 (O_4794,N_48137,N_49479);
and UO_4795 (O_4795,N_48738,N_49478);
and UO_4796 (O_4796,N_48923,N_49352);
xnor UO_4797 (O_4797,N_48148,N_49662);
and UO_4798 (O_4798,N_49926,N_49543);
nand UO_4799 (O_4799,N_48505,N_49889);
and UO_4800 (O_4800,N_48066,N_48684);
or UO_4801 (O_4801,N_48310,N_48953);
or UO_4802 (O_4802,N_49032,N_48847);
xnor UO_4803 (O_4803,N_49439,N_49468);
xnor UO_4804 (O_4804,N_47939,N_49706);
and UO_4805 (O_4805,N_48521,N_48812);
xor UO_4806 (O_4806,N_49593,N_49633);
nand UO_4807 (O_4807,N_48039,N_48550);
nor UO_4808 (O_4808,N_48150,N_48257);
nand UO_4809 (O_4809,N_48185,N_49208);
nand UO_4810 (O_4810,N_49798,N_49602);
and UO_4811 (O_4811,N_48742,N_49207);
nand UO_4812 (O_4812,N_47858,N_47517);
and UO_4813 (O_4813,N_47694,N_47979);
xor UO_4814 (O_4814,N_47737,N_48797);
nand UO_4815 (O_4815,N_47922,N_47772);
xor UO_4816 (O_4816,N_48388,N_48101);
nor UO_4817 (O_4817,N_48891,N_48613);
nor UO_4818 (O_4818,N_49064,N_49269);
and UO_4819 (O_4819,N_48365,N_48077);
or UO_4820 (O_4820,N_49571,N_48756);
or UO_4821 (O_4821,N_49387,N_49488);
and UO_4822 (O_4822,N_48192,N_49650);
xor UO_4823 (O_4823,N_49824,N_47538);
nor UO_4824 (O_4824,N_47603,N_48184);
xnor UO_4825 (O_4825,N_48600,N_47503);
xnor UO_4826 (O_4826,N_48952,N_48873);
xnor UO_4827 (O_4827,N_49763,N_49397);
or UO_4828 (O_4828,N_48530,N_48471);
and UO_4829 (O_4829,N_49611,N_47622);
and UO_4830 (O_4830,N_49564,N_49947);
nor UO_4831 (O_4831,N_49622,N_49513);
nor UO_4832 (O_4832,N_47511,N_48460);
xnor UO_4833 (O_4833,N_48314,N_48190);
xor UO_4834 (O_4834,N_48667,N_49232);
nor UO_4835 (O_4835,N_49504,N_48396);
nand UO_4836 (O_4836,N_49864,N_47584);
and UO_4837 (O_4837,N_47891,N_48252);
nand UO_4838 (O_4838,N_48956,N_47985);
and UO_4839 (O_4839,N_47735,N_48005);
xnor UO_4840 (O_4840,N_47922,N_47725);
nor UO_4841 (O_4841,N_49515,N_48685);
or UO_4842 (O_4842,N_48654,N_47991);
nand UO_4843 (O_4843,N_49639,N_47964);
or UO_4844 (O_4844,N_47884,N_49718);
nand UO_4845 (O_4845,N_48650,N_48801);
xor UO_4846 (O_4846,N_49056,N_48877);
xor UO_4847 (O_4847,N_47858,N_49211);
xnor UO_4848 (O_4848,N_49754,N_49122);
nor UO_4849 (O_4849,N_48549,N_48450);
nor UO_4850 (O_4850,N_49595,N_48634);
xor UO_4851 (O_4851,N_49165,N_47799);
nor UO_4852 (O_4852,N_48281,N_48614);
or UO_4853 (O_4853,N_47583,N_49321);
nor UO_4854 (O_4854,N_49416,N_48620);
nand UO_4855 (O_4855,N_48546,N_47761);
nand UO_4856 (O_4856,N_48593,N_47519);
and UO_4857 (O_4857,N_48872,N_48611);
or UO_4858 (O_4858,N_47527,N_47560);
nand UO_4859 (O_4859,N_48428,N_48569);
and UO_4860 (O_4860,N_49797,N_49622);
or UO_4861 (O_4861,N_49704,N_47959);
nand UO_4862 (O_4862,N_48682,N_47868);
and UO_4863 (O_4863,N_49108,N_48152);
and UO_4864 (O_4864,N_49094,N_48251);
nor UO_4865 (O_4865,N_49224,N_47817);
xnor UO_4866 (O_4866,N_49391,N_49535);
and UO_4867 (O_4867,N_47898,N_49120);
nand UO_4868 (O_4868,N_49145,N_48497);
nor UO_4869 (O_4869,N_49732,N_48513);
and UO_4870 (O_4870,N_49722,N_49664);
or UO_4871 (O_4871,N_47515,N_49345);
and UO_4872 (O_4872,N_49611,N_49396);
and UO_4873 (O_4873,N_49363,N_48230);
xnor UO_4874 (O_4874,N_48640,N_49423);
nand UO_4875 (O_4875,N_49141,N_49745);
nand UO_4876 (O_4876,N_47895,N_48927);
and UO_4877 (O_4877,N_49296,N_47647);
nor UO_4878 (O_4878,N_49903,N_49705);
and UO_4879 (O_4879,N_48696,N_47534);
and UO_4880 (O_4880,N_47773,N_48579);
and UO_4881 (O_4881,N_49474,N_48111);
or UO_4882 (O_4882,N_49530,N_47744);
xnor UO_4883 (O_4883,N_49852,N_48829);
and UO_4884 (O_4884,N_48899,N_49987);
nor UO_4885 (O_4885,N_49277,N_47856);
and UO_4886 (O_4886,N_47551,N_49701);
xor UO_4887 (O_4887,N_49169,N_48820);
or UO_4888 (O_4888,N_49078,N_48214);
nor UO_4889 (O_4889,N_47979,N_48566);
nor UO_4890 (O_4890,N_47687,N_48416);
or UO_4891 (O_4891,N_47608,N_49345);
nor UO_4892 (O_4892,N_48113,N_48782);
xor UO_4893 (O_4893,N_48797,N_48903);
nand UO_4894 (O_4894,N_48548,N_48545);
nand UO_4895 (O_4895,N_49547,N_48354);
nor UO_4896 (O_4896,N_47762,N_47657);
nand UO_4897 (O_4897,N_47741,N_49618);
or UO_4898 (O_4898,N_49204,N_49144);
or UO_4899 (O_4899,N_47788,N_48442);
xor UO_4900 (O_4900,N_48055,N_47792);
nor UO_4901 (O_4901,N_49388,N_48737);
xor UO_4902 (O_4902,N_48487,N_48732);
xnor UO_4903 (O_4903,N_49690,N_47773);
nand UO_4904 (O_4904,N_47541,N_49002);
and UO_4905 (O_4905,N_48433,N_49647);
nor UO_4906 (O_4906,N_48773,N_49352);
nand UO_4907 (O_4907,N_48350,N_49945);
nor UO_4908 (O_4908,N_48001,N_48722);
xor UO_4909 (O_4909,N_49208,N_47531);
or UO_4910 (O_4910,N_48980,N_49369);
and UO_4911 (O_4911,N_48426,N_48043);
or UO_4912 (O_4912,N_48301,N_48809);
and UO_4913 (O_4913,N_49238,N_49828);
and UO_4914 (O_4914,N_47551,N_49267);
and UO_4915 (O_4915,N_48564,N_49633);
nand UO_4916 (O_4916,N_47943,N_49729);
nand UO_4917 (O_4917,N_48684,N_48880);
nor UO_4918 (O_4918,N_47898,N_49356);
or UO_4919 (O_4919,N_49683,N_49088);
or UO_4920 (O_4920,N_47596,N_49806);
nor UO_4921 (O_4921,N_48371,N_49753);
xor UO_4922 (O_4922,N_49804,N_49281);
nor UO_4923 (O_4923,N_47818,N_48422);
nand UO_4924 (O_4924,N_48972,N_48597);
xnor UO_4925 (O_4925,N_49963,N_47702);
nor UO_4926 (O_4926,N_49652,N_47584);
or UO_4927 (O_4927,N_47954,N_49933);
xnor UO_4928 (O_4928,N_48801,N_49753);
xnor UO_4929 (O_4929,N_47965,N_49306);
nand UO_4930 (O_4930,N_48520,N_48502);
and UO_4931 (O_4931,N_49235,N_47924);
or UO_4932 (O_4932,N_48475,N_47558);
or UO_4933 (O_4933,N_49784,N_49718);
xor UO_4934 (O_4934,N_47738,N_48845);
nand UO_4935 (O_4935,N_48198,N_47541);
or UO_4936 (O_4936,N_48460,N_48848);
nand UO_4937 (O_4937,N_48371,N_49266);
nor UO_4938 (O_4938,N_47649,N_48601);
or UO_4939 (O_4939,N_47998,N_48215);
xor UO_4940 (O_4940,N_48910,N_49813);
nor UO_4941 (O_4941,N_49678,N_49220);
xor UO_4942 (O_4942,N_49109,N_48612);
nand UO_4943 (O_4943,N_49665,N_47983);
nand UO_4944 (O_4944,N_49420,N_48308);
or UO_4945 (O_4945,N_48537,N_49388);
and UO_4946 (O_4946,N_48184,N_49487);
and UO_4947 (O_4947,N_49808,N_47687);
xor UO_4948 (O_4948,N_49149,N_48548);
and UO_4949 (O_4949,N_49199,N_48755);
or UO_4950 (O_4950,N_48204,N_48384);
and UO_4951 (O_4951,N_49124,N_49097);
or UO_4952 (O_4952,N_47569,N_49345);
or UO_4953 (O_4953,N_48395,N_49849);
xor UO_4954 (O_4954,N_48084,N_48523);
and UO_4955 (O_4955,N_49785,N_49129);
nand UO_4956 (O_4956,N_47996,N_49846);
nor UO_4957 (O_4957,N_49159,N_47579);
xor UO_4958 (O_4958,N_47973,N_48563);
nand UO_4959 (O_4959,N_48086,N_47770);
or UO_4960 (O_4960,N_48057,N_49091);
xnor UO_4961 (O_4961,N_49414,N_47550);
nand UO_4962 (O_4962,N_49334,N_47757);
and UO_4963 (O_4963,N_48466,N_47754);
nand UO_4964 (O_4964,N_47682,N_49384);
or UO_4965 (O_4965,N_47912,N_49533);
nor UO_4966 (O_4966,N_48085,N_48137);
nor UO_4967 (O_4967,N_48570,N_48134);
nor UO_4968 (O_4968,N_48146,N_49989);
and UO_4969 (O_4969,N_49047,N_47709);
nor UO_4970 (O_4970,N_48044,N_49265);
or UO_4971 (O_4971,N_49070,N_49237);
and UO_4972 (O_4972,N_47604,N_49319);
nor UO_4973 (O_4973,N_48095,N_48582);
nor UO_4974 (O_4974,N_48495,N_47911);
or UO_4975 (O_4975,N_48893,N_48821);
and UO_4976 (O_4976,N_47694,N_48911);
or UO_4977 (O_4977,N_48645,N_48660);
nand UO_4978 (O_4978,N_49655,N_48440);
or UO_4979 (O_4979,N_47664,N_49768);
or UO_4980 (O_4980,N_48926,N_48858);
nor UO_4981 (O_4981,N_49083,N_49041);
xnor UO_4982 (O_4982,N_48094,N_49315);
nand UO_4983 (O_4983,N_47655,N_49488);
nand UO_4984 (O_4984,N_47685,N_48755);
nand UO_4985 (O_4985,N_48142,N_47576);
xnor UO_4986 (O_4986,N_48405,N_48471);
and UO_4987 (O_4987,N_49900,N_49303);
nand UO_4988 (O_4988,N_49522,N_49109);
nor UO_4989 (O_4989,N_48154,N_48075);
xnor UO_4990 (O_4990,N_48641,N_49755);
or UO_4991 (O_4991,N_49604,N_48567);
and UO_4992 (O_4992,N_48416,N_49222);
nor UO_4993 (O_4993,N_48177,N_48190);
or UO_4994 (O_4994,N_49240,N_48499);
nand UO_4995 (O_4995,N_49773,N_48902);
and UO_4996 (O_4996,N_47911,N_49312);
xor UO_4997 (O_4997,N_48248,N_48244);
xnor UO_4998 (O_4998,N_47554,N_49030);
or UO_4999 (O_4999,N_48709,N_49005);
endmodule